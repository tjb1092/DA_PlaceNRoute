magic
tech scmos
timestamp 1555071808 
<< pdiffusion >>
rect 1 -12 7 -6
rect 8 -12 14 -6
rect 15 -12 21 -6
rect 22 -12 28 -6
rect 29 -12 35 -6
rect 36 -12 42 -6
rect 43 -12 49 -6
rect 50 -12 56 -6
rect 57 -12 63 -6
rect 64 -12 70 -6
rect 71 -12 77 -6
rect 78 -12 84 -6
rect 85 -12 91 -6
rect 92 -12 98 -6
rect 99 -12 105 -6
rect 106 -12 112 -6
rect 113 -12 119 -6
rect 120 -12 126 -6
rect 127 -12 133 -6
rect 134 -12 140 -6
rect 141 -12 147 -6
rect 148 -12 154 -6
rect 281 -12 287 -6
rect 316 -12 319 -6
rect 344 -12 347 -6
rect 351 -12 357 -6
rect 421 -12 427 -6
rect 435 -12 441 -6
rect 442 -12 445 -6
rect 449 -12 452 -6
rect 456 -12 462 -6
rect 463 -12 466 -6
rect 477 -12 483 -6
rect 505 -12 511 -6
rect 512 -12 515 -6
rect 904 -12 907 -6
rect 946 -12 952 -6
rect 988 -12 991 -6
rect 1 -31 7 -25
rect 8 -31 14 -25
rect 15 -31 21 -25
rect 22 -31 28 -25
rect 29 -31 35 -25
rect 36 -31 42 -25
rect 43 -31 49 -25
rect 50 -31 56 -25
rect 57 -31 63 -25
rect 64 -31 70 -25
rect 71 -31 77 -25
rect 78 -31 84 -25
rect 85 -31 91 -25
rect 92 -31 98 -25
rect 99 -31 105 -25
rect 106 -31 112 -25
rect 113 -31 119 -25
rect 225 -31 228 -25
rect 288 -31 291 -25
rect 302 -31 305 -25
rect 337 -31 340 -25
rect 344 -31 350 -25
rect 351 -31 354 -25
rect 358 -31 364 -25
rect 365 -31 368 -25
rect 372 -31 375 -25
rect 379 -31 382 -25
rect 386 -31 389 -25
rect 393 -31 396 -25
rect 407 -31 410 -25
rect 414 -31 420 -25
rect 421 -31 424 -25
rect 435 -31 438 -25
rect 449 -31 452 -25
rect 456 -31 459 -25
rect 463 -31 466 -25
rect 498 -31 501 -25
rect 505 -31 511 -25
rect 512 -31 515 -25
rect 519 -31 525 -25
rect 526 -31 532 -25
rect 533 -31 539 -25
rect 540 -31 543 -25
rect 547 -31 550 -25
rect 575 -31 581 -25
rect 582 -31 588 -25
rect 589 -31 592 -25
rect 596 -31 599 -25
rect 603 -31 606 -25
rect 610 -31 613 -25
rect 617 -31 623 -25
rect 624 -31 627 -25
rect 631 -31 637 -25
rect 638 -31 644 -25
rect 673 -31 676 -25
rect 890 -31 893 -25
rect 1002 -31 1005 -25
rect 1 -54 7 -48
rect 8 -54 14 -48
rect 15 -54 21 -48
rect 22 -54 28 -48
rect 29 -54 35 -48
rect 36 -54 42 -48
rect 43 -54 49 -48
rect 50 -54 56 -48
rect 57 -54 63 -48
rect 64 -54 70 -48
rect 71 -54 77 -48
rect 78 -54 84 -48
rect 85 -54 91 -48
rect 92 -54 98 -48
rect 99 -54 105 -48
rect 106 -54 112 -48
rect 218 -54 221 -48
rect 274 -54 277 -48
rect 281 -54 284 -48
rect 295 -54 301 -48
rect 302 -54 305 -48
rect 316 -54 322 -48
rect 323 -54 326 -48
rect 330 -54 333 -48
rect 337 -54 343 -48
rect 344 -54 347 -48
rect 351 -54 354 -48
rect 358 -54 361 -48
rect 365 -54 368 -48
rect 372 -54 375 -48
rect 379 -54 382 -48
rect 386 -54 392 -48
rect 393 -54 396 -48
rect 400 -54 403 -48
rect 407 -54 410 -48
rect 414 -54 417 -48
rect 421 -54 424 -48
rect 428 -54 434 -48
rect 435 -54 438 -48
rect 442 -54 445 -48
rect 449 -54 452 -48
rect 456 -54 462 -48
rect 463 -54 466 -48
rect 470 -54 473 -48
rect 484 -54 487 -48
rect 491 -54 494 -48
rect 498 -54 501 -48
rect 505 -54 508 -48
rect 519 -54 522 -48
rect 540 -54 543 -48
rect 547 -54 553 -48
rect 554 -54 557 -48
rect 561 -54 567 -48
rect 568 -54 574 -48
rect 575 -54 578 -48
rect 582 -54 585 -48
rect 589 -54 592 -48
rect 596 -54 599 -48
rect 603 -54 606 -48
rect 610 -54 616 -48
rect 617 -54 623 -48
rect 624 -54 627 -48
rect 631 -54 634 -48
rect 638 -54 641 -48
rect 652 -54 655 -48
rect 673 -54 676 -48
rect 680 -54 686 -48
rect 722 -54 725 -48
rect 729 -54 732 -48
rect 757 -54 760 -48
rect 827 -54 833 -48
rect 883 -54 886 -48
rect 1009 -54 1012 -48
rect 1 -105 7 -99
rect 8 -105 14 -99
rect 15 -105 21 -99
rect 22 -105 28 -99
rect 29 -105 35 -99
rect 36 -105 42 -99
rect 43 -105 49 -99
rect 50 -105 56 -99
rect 57 -105 63 -99
rect 64 -105 70 -99
rect 71 -105 77 -99
rect 78 -105 84 -99
rect 190 -105 193 -99
rect 204 -105 207 -99
rect 218 -105 221 -99
rect 232 -105 235 -99
rect 239 -105 245 -99
rect 246 -105 249 -99
rect 253 -105 259 -99
rect 260 -105 263 -99
rect 267 -105 273 -99
rect 274 -105 280 -99
rect 281 -105 284 -99
rect 288 -105 291 -99
rect 295 -105 301 -99
rect 302 -105 305 -99
rect 309 -105 312 -99
rect 316 -105 319 -99
rect 323 -105 326 -99
rect 330 -105 333 -99
rect 337 -105 340 -99
rect 344 -105 347 -99
rect 351 -105 354 -99
rect 358 -105 361 -99
rect 365 -105 368 -99
rect 372 -105 375 -99
rect 379 -105 385 -99
rect 386 -105 392 -99
rect 393 -105 396 -99
rect 400 -105 403 -99
rect 407 -105 410 -99
rect 414 -105 417 -99
rect 421 -105 424 -99
rect 428 -105 431 -99
rect 435 -105 438 -99
rect 442 -105 445 -99
rect 449 -105 452 -99
rect 456 -105 459 -99
rect 463 -105 466 -99
rect 470 -105 473 -99
rect 477 -105 480 -99
rect 484 -105 487 -99
rect 491 -105 494 -99
rect 498 -105 501 -99
rect 505 -105 511 -99
rect 512 -105 518 -99
rect 519 -105 525 -99
rect 526 -105 529 -99
rect 533 -105 539 -99
rect 540 -105 546 -99
rect 547 -105 550 -99
rect 554 -105 557 -99
rect 561 -105 567 -99
rect 568 -105 571 -99
rect 575 -105 578 -99
rect 582 -105 588 -99
rect 589 -105 592 -99
rect 596 -105 599 -99
rect 603 -105 606 -99
rect 610 -105 613 -99
rect 617 -105 620 -99
rect 624 -105 630 -99
rect 631 -105 634 -99
rect 638 -105 641 -99
rect 645 -105 648 -99
rect 652 -105 655 -99
rect 659 -105 662 -99
rect 666 -105 669 -99
rect 680 -105 683 -99
rect 687 -105 690 -99
rect 701 -105 704 -99
rect 708 -105 711 -99
rect 722 -105 725 -99
rect 729 -105 732 -99
rect 736 -105 739 -99
rect 778 -105 784 -99
rect 785 -105 791 -99
rect 792 -105 795 -99
rect 799 -105 805 -99
rect 806 -105 809 -99
rect 862 -105 865 -99
rect 890 -105 893 -99
rect 897 -105 900 -99
rect 1016 -105 1019 -99
rect 1 -172 7 -166
rect 8 -172 14 -166
rect 15 -172 21 -166
rect 22 -172 28 -166
rect 29 -172 35 -166
rect 36 -172 42 -166
rect 43 -172 49 -166
rect 50 -172 56 -166
rect 57 -172 63 -166
rect 64 -172 70 -166
rect 71 -172 77 -166
rect 78 -172 84 -166
rect 113 -172 116 -166
rect 120 -172 123 -166
rect 127 -172 130 -166
rect 134 -172 137 -166
rect 141 -172 144 -166
rect 148 -172 151 -166
rect 155 -172 158 -166
rect 162 -172 165 -166
rect 169 -172 172 -166
rect 176 -172 179 -166
rect 183 -172 186 -166
rect 190 -172 193 -166
rect 197 -172 200 -166
rect 204 -172 207 -166
rect 211 -172 214 -166
rect 218 -172 221 -166
rect 225 -172 231 -166
rect 232 -172 235 -166
rect 239 -172 242 -166
rect 246 -172 249 -166
rect 253 -172 256 -166
rect 260 -172 263 -166
rect 267 -172 270 -166
rect 274 -172 277 -166
rect 281 -172 284 -166
rect 288 -172 291 -166
rect 295 -172 301 -166
rect 302 -172 305 -166
rect 309 -172 312 -166
rect 316 -172 319 -166
rect 323 -172 326 -166
rect 330 -172 336 -166
rect 337 -172 340 -166
rect 344 -172 347 -166
rect 351 -172 354 -166
rect 358 -172 361 -166
rect 365 -172 371 -166
rect 372 -172 375 -166
rect 379 -172 382 -166
rect 386 -172 392 -166
rect 393 -172 396 -166
rect 400 -172 406 -166
rect 407 -172 410 -166
rect 414 -172 417 -166
rect 421 -172 424 -166
rect 428 -172 431 -166
rect 435 -172 438 -166
rect 442 -172 445 -166
rect 449 -172 455 -166
rect 456 -172 459 -166
rect 463 -172 466 -166
rect 470 -172 473 -166
rect 477 -172 480 -166
rect 484 -172 487 -166
rect 491 -172 494 -166
rect 498 -172 504 -166
rect 505 -172 508 -166
rect 512 -172 518 -166
rect 519 -172 525 -166
rect 526 -172 532 -166
rect 533 -172 536 -166
rect 540 -172 543 -166
rect 547 -172 550 -166
rect 554 -172 560 -166
rect 561 -172 564 -166
rect 568 -172 574 -166
rect 575 -172 578 -166
rect 582 -172 585 -166
rect 589 -172 595 -166
rect 596 -172 599 -166
rect 603 -172 609 -166
rect 610 -172 616 -166
rect 617 -172 620 -166
rect 624 -172 627 -166
rect 631 -172 634 -166
rect 638 -172 641 -166
rect 645 -172 648 -166
rect 652 -172 658 -166
rect 659 -172 662 -166
rect 666 -172 669 -166
rect 673 -172 676 -166
rect 680 -172 683 -166
rect 687 -172 690 -166
rect 694 -172 697 -166
rect 701 -172 704 -166
rect 708 -172 711 -166
rect 715 -172 718 -166
rect 722 -172 725 -166
rect 729 -172 735 -166
rect 736 -172 739 -166
rect 743 -172 746 -166
rect 750 -172 753 -166
rect 757 -172 760 -166
rect 764 -172 767 -166
rect 771 -172 774 -166
rect 778 -172 781 -166
rect 785 -172 788 -166
rect 792 -172 795 -166
rect 799 -172 802 -166
rect 806 -172 809 -166
rect 813 -172 816 -166
rect 820 -172 823 -166
rect 827 -172 830 -166
rect 834 -172 837 -166
rect 841 -172 844 -166
rect 848 -172 851 -166
rect 855 -172 858 -166
rect 862 -172 865 -166
rect 869 -172 872 -166
rect 876 -172 879 -166
rect 897 -172 900 -166
rect 918 -172 921 -166
rect 939 -172 942 -166
rect 1009 -172 1015 -166
rect 1023 -172 1026 -166
rect 1135 -172 1138 -166
rect 1170 -172 1173 -166
rect 1 -239 7 -233
rect 8 -239 14 -233
rect 15 -239 21 -233
rect 22 -239 28 -233
rect 29 -239 35 -233
rect 36 -239 42 -233
rect 43 -239 49 -233
rect 50 -239 56 -233
rect 57 -239 63 -233
rect 64 -239 70 -233
rect 71 -239 74 -233
rect 78 -239 81 -233
rect 85 -239 88 -233
rect 92 -239 95 -233
rect 99 -239 102 -233
rect 106 -239 109 -233
rect 113 -239 116 -233
rect 120 -239 123 -233
rect 127 -239 130 -233
rect 134 -239 137 -233
rect 141 -239 144 -233
rect 148 -239 151 -233
rect 155 -239 161 -233
rect 162 -239 165 -233
rect 169 -239 172 -233
rect 176 -239 179 -233
rect 183 -239 186 -233
rect 190 -239 193 -233
rect 197 -239 200 -233
rect 204 -239 210 -233
rect 211 -239 214 -233
rect 218 -239 224 -233
rect 225 -239 231 -233
rect 232 -239 238 -233
rect 239 -239 245 -233
rect 246 -239 249 -233
rect 253 -239 259 -233
rect 260 -239 263 -233
rect 267 -239 270 -233
rect 274 -239 277 -233
rect 281 -239 284 -233
rect 288 -239 291 -233
rect 295 -239 298 -233
rect 302 -239 305 -233
rect 309 -239 312 -233
rect 316 -239 319 -233
rect 323 -239 326 -233
rect 330 -239 333 -233
rect 337 -239 340 -233
rect 344 -239 347 -233
rect 351 -239 354 -233
rect 358 -239 361 -233
rect 365 -239 371 -233
rect 372 -239 375 -233
rect 379 -239 382 -233
rect 386 -239 389 -233
rect 393 -239 396 -233
rect 400 -239 403 -233
rect 407 -239 413 -233
rect 414 -239 417 -233
rect 421 -239 424 -233
rect 428 -239 434 -233
rect 435 -239 438 -233
rect 442 -239 448 -233
rect 449 -239 455 -233
rect 456 -239 459 -233
rect 463 -239 466 -233
rect 470 -239 473 -233
rect 477 -239 483 -233
rect 484 -239 490 -233
rect 491 -239 494 -233
rect 498 -239 504 -233
rect 505 -239 508 -233
rect 512 -239 515 -233
rect 519 -239 522 -233
rect 526 -239 529 -233
rect 533 -239 536 -233
rect 540 -239 543 -233
rect 547 -239 553 -233
rect 554 -239 557 -233
rect 561 -239 564 -233
rect 568 -239 571 -233
rect 575 -239 578 -233
rect 582 -239 585 -233
rect 589 -239 592 -233
rect 596 -239 599 -233
rect 603 -239 606 -233
rect 610 -239 616 -233
rect 617 -239 620 -233
rect 624 -239 630 -233
rect 631 -239 634 -233
rect 638 -239 641 -233
rect 645 -239 648 -233
rect 652 -239 655 -233
rect 659 -239 662 -233
rect 666 -239 669 -233
rect 673 -239 676 -233
rect 680 -239 683 -233
rect 687 -239 690 -233
rect 694 -239 697 -233
rect 701 -239 704 -233
rect 708 -239 711 -233
rect 715 -239 718 -233
rect 722 -239 725 -233
rect 729 -239 732 -233
rect 736 -239 739 -233
rect 743 -239 746 -233
rect 750 -239 756 -233
rect 757 -239 760 -233
rect 764 -239 767 -233
rect 771 -239 774 -233
rect 778 -239 781 -233
rect 785 -239 788 -233
rect 792 -239 795 -233
rect 799 -239 802 -233
rect 806 -239 809 -233
rect 813 -239 816 -233
rect 820 -239 823 -233
rect 827 -239 833 -233
rect 834 -239 837 -233
rect 841 -239 844 -233
rect 848 -239 854 -233
rect 855 -239 858 -233
rect 862 -239 865 -233
rect 869 -239 872 -233
rect 876 -239 879 -233
rect 883 -239 886 -233
rect 890 -239 893 -233
rect 897 -239 900 -233
rect 904 -239 907 -233
rect 911 -239 914 -233
rect 918 -239 921 -233
rect 925 -239 928 -233
rect 932 -239 935 -233
rect 939 -239 942 -233
rect 946 -239 949 -233
rect 953 -239 956 -233
rect 960 -239 963 -233
rect 967 -239 970 -233
rect 974 -239 977 -233
rect 981 -239 984 -233
rect 988 -239 991 -233
rect 995 -239 998 -233
rect 1002 -239 1005 -233
rect 1009 -239 1012 -233
rect 1016 -239 1019 -233
rect 1023 -239 1026 -233
rect 1037 -239 1040 -233
rect 1184 -239 1187 -233
rect 1324 -239 1327 -233
rect 1 -322 7 -316
rect 8 -322 14 -316
rect 15 -322 21 -316
rect 22 -322 28 -316
rect 29 -322 35 -316
rect 36 -322 42 -316
rect 43 -322 49 -316
rect 50 -322 56 -316
rect 57 -322 63 -316
rect 64 -322 67 -316
rect 71 -322 77 -316
rect 78 -322 81 -316
rect 85 -322 88 -316
rect 92 -322 95 -316
rect 99 -322 102 -316
rect 106 -322 109 -316
rect 113 -322 116 -316
rect 120 -322 123 -316
rect 127 -322 130 -316
rect 134 -322 140 -316
rect 141 -322 147 -316
rect 148 -322 151 -316
rect 155 -322 158 -316
rect 162 -322 165 -316
rect 169 -322 175 -316
rect 176 -322 179 -316
rect 183 -322 189 -316
rect 190 -322 193 -316
rect 197 -322 200 -316
rect 204 -322 210 -316
rect 211 -322 214 -316
rect 218 -322 221 -316
rect 225 -322 228 -316
rect 232 -322 235 -316
rect 239 -322 242 -316
rect 246 -322 249 -316
rect 253 -322 256 -316
rect 260 -322 263 -316
rect 267 -322 270 -316
rect 274 -322 277 -316
rect 281 -322 284 -316
rect 288 -322 291 -316
rect 295 -322 298 -316
rect 302 -322 305 -316
rect 309 -322 315 -316
rect 316 -322 319 -316
rect 323 -322 326 -316
rect 330 -322 333 -316
rect 337 -322 340 -316
rect 344 -322 347 -316
rect 351 -322 354 -316
rect 358 -322 361 -316
rect 365 -322 368 -316
rect 372 -322 378 -316
rect 379 -322 385 -316
rect 386 -322 392 -316
rect 393 -322 396 -316
rect 400 -322 403 -316
rect 407 -322 410 -316
rect 414 -322 417 -316
rect 421 -322 424 -316
rect 428 -322 431 -316
rect 435 -322 438 -316
rect 442 -322 448 -316
rect 449 -322 452 -316
rect 456 -322 459 -316
rect 463 -322 466 -316
rect 470 -322 473 -316
rect 477 -322 483 -316
rect 484 -322 487 -316
rect 491 -322 494 -316
rect 498 -322 501 -316
rect 505 -322 508 -316
rect 512 -322 515 -316
rect 519 -322 522 -316
rect 526 -322 529 -316
rect 533 -322 539 -316
rect 540 -322 543 -316
rect 547 -322 553 -316
rect 554 -322 557 -316
rect 561 -322 564 -316
rect 568 -322 571 -316
rect 575 -322 578 -316
rect 582 -322 585 -316
rect 589 -322 595 -316
rect 596 -322 602 -316
rect 603 -322 609 -316
rect 610 -322 613 -316
rect 617 -322 620 -316
rect 624 -322 630 -316
rect 631 -322 634 -316
rect 638 -322 641 -316
rect 645 -322 651 -316
rect 652 -322 655 -316
rect 659 -322 662 -316
rect 666 -322 672 -316
rect 673 -322 676 -316
rect 680 -322 683 -316
rect 687 -322 690 -316
rect 694 -322 700 -316
rect 701 -322 704 -316
rect 708 -322 711 -316
rect 715 -322 718 -316
rect 722 -322 725 -316
rect 729 -322 732 -316
rect 736 -322 739 -316
rect 743 -322 749 -316
rect 750 -322 753 -316
rect 757 -322 760 -316
rect 764 -322 767 -316
rect 771 -322 774 -316
rect 778 -322 781 -316
rect 785 -322 788 -316
rect 792 -322 795 -316
rect 799 -322 802 -316
rect 806 -322 809 -316
rect 813 -322 816 -316
rect 820 -322 823 -316
rect 827 -322 830 -316
rect 834 -322 837 -316
rect 841 -322 844 -316
rect 848 -322 851 -316
rect 855 -322 858 -316
rect 862 -322 865 -316
rect 869 -322 872 -316
rect 876 -322 879 -316
rect 883 -322 886 -316
rect 890 -322 893 -316
rect 897 -322 900 -316
rect 904 -322 907 -316
rect 911 -322 914 -316
rect 918 -322 921 -316
rect 925 -322 928 -316
rect 932 -322 935 -316
rect 939 -322 942 -316
rect 946 -322 949 -316
rect 953 -322 956 -316
rect 960 -322 963 -316
rect 967 -322 970 -316
rect 974 -322 977 -316
rect 981 -322 984 -316
rect 988 -322 991 -316
rect 995 -322 998 -316
rect 1002 -322 1005 -316
rect 1009 -322 1012 -316
rect 1016 -322 1019 -316
rect 1023 -322 1026 -316
rect 1030 -322 1033 -316
rect 1037 -322 1040 -316
rect 1044 -322 1047 -316
rect 1051 -322 1054 -316
rect 1058 -322 1061 -316
rect 1065 -322 1068 -316
rect 1072 -322 1075 -316
rect 1079 -322 1082 -316
rect 1086 -322 1089 -316
rect 1093 -322 1096 -316
rect 1100 -322 1103 -316
rect 1107 -322 1110 -316
rect 1114 -322 1117 -316
rect 1121 -322 1124 -316
rect 1205 -322 1208 -316
rect 1303 -322 1309 -316
rect 1380 -322 1383 -316
rect 1457 -322 1460 -316
rect 1 -421 7 -415
rect 8 -421 14 -415
rect 15 -421 21 -415
rect 22 -421 28 -415
rect 29 -421 35 -415
rect 36 -421 42 -415
rect 43 -421 49 -415
rect 50 -421 56 -415
rect 57 -421 63 -415
rect 64 -421 70 -415
rect 71 -421 74 -415
rect 78 -421 81 -415
rect 85 -421 88 -415
rect 92 -421 95 -415
rect 99 -421 102 -415
rect 106 -421 109 -415
rect 113 -421 116 -415
rect 120 -421 123 -415
rect 127 -421 130 -415
rect 134 -421 137 -415
rect 141 -421 144 -415
rect 148 -421 154 -415
rect 155 -421 158 -415
rect 162 -421 168 -415
rect 169 -421 175 -415
rect 176 -421 179 -415
rect 183 -421 189 -415
rect 190 -421 196 -415
rect 197 -421 200 -415
rect 204 -421 207 -415
rect 211 -421 214 -415
rect 218 -421 221 -415
rect 225 -421 228 -415
rect 232 -421 235 -415
rect 239 -421 242 -415
rect 246 -421 252 -415
rect 253 -421 256 -415
rect 260 -421 263 -415
rect 267 -421 270 -415
rect 274 -421 277 -415
rect 281 -421 284 -415
rect 288 -421 291 -415
rect 295 -421 298 -415
rect 302 -421 305 -415
rect 309 -421 312 -415
rect 316 -421 319 -415
rect 323 -421 326 -415
rect 330 -421 333 -415
rect 337 -421 340 -415
rect 344 -421 347 -415
rect 351 -421 354 -415
rect 358 -421 364 -415
rect 365 -421 371 -415
rect 372 -421 375 -415
rect 379 -421 385 -415
rect 386 -421 389 -415
rect 393 -421 396 -415
rect 400 -421 403 -415
rect 407 -421 410 -415
rect 414 -421 420 -415
rect 421 -421 424 -415
rect 428 -421 431 -415
rect 435 -421 438 -415
rect 442 -421 445 -415
rect 449 -421 452 -415
rect 456 -421 459 -415
rect 463 -421 466 -415
rect 470 -421 473 -415
rect 477 -421 480 -415
rect 484 -421 487 -415
rect 491 -421 497 -415
rect 498 -421 501 -415
rect 505 -421 508 -415
rect 512 -421 515 -415
rect 519 -421 522 -415
rect 526 -421 529 -415
rect 533 -421 536 -415
rect 540 -421 546 -415
rect 547 -421 550 -415
rect 554 -421 557 -415
rect 561 -421 567 -415
rect 568 -421 574 -415
rect 575 -421 578 -415
rect 582 -421 588 -415
rect 589 -421 592 -415
rect 596 -421 599 -415
rect 603 -421 606 -415
rect 610 -421 613 -415
rect 617 -421 620 -415
rect 624 -421 630 -415
rect 631 -421 637 -415
rect 638 -421 641 -415
rect 645 -421 648 -415
rect 652 -421 655 -415
rect 659 -421 662 -415
rect 666 -421 669 -415
rect 673 -421 676 -415
rect 680 -421 683 -415
rect 687 -421 693 -415
rect 694 -421 697 -415
rect 701 -421 704 -415
rect 708 -421 711 -415
rect 715 -421 721 -415
rect 722 -421 728 -415
rect 729 -421 732 -415
rect 736 -421 739 -415
rect 743 -421 746 -415
rect 750 -421 753 -415
rect 757 -421 760 -415
rect 764 -421 767 -415
rect 771 -421 774 -415
rect 778 -421 781 -415
rect 785 -421 791 -415
rect 792 -421 795 -415
rect 799 -421 802 -415
rect 806 -421 809 -415
rect 813 -421 816 -415
rect 820 -421 823 -415
rect 827 -421 830 -415
rect 834 -421 840 -415
rect 841 -421 844 -415
rect 848 -421 851 -415
rect 855 -421 858 -415
rect 862 -421 865 -415
rect 869 -421 872 -415
rect 876 -421 879 -415
rect 883 -421 886 -415
rect 890 -421 893 -415
rect 897 -421 900 -415
rect 904 -421 907 -415
rect 911 -421 914 -415
rect 918 -421 921 -415
rect 925 -421 928 -415
rect 932 -421 935 -415
rect 939 -421 942 -415
rect 946 -421 949 -415
rect 953 -421 956 -415
rect 960 -421 963 -415
rect 967 -421 970 -415
rect 974 -421 977 -415
rect 981 -421 984 -415
rect 988 -421 991 -415
rect 995 -421 998 -415
rect 1002 -421 1005 -415
rect 1009 -421 1012 -415
rect 1016 -421 1019 -415
rect 1023 -421 1026 -415
rect 1030 -421 1033 -415
rect 1037 -421 1040 -415
rect 1044 -421 1047 -415
rect 1051 -421 1054 -415
rect 1058 -421 1061 -415
rect 1065 -421 1068 -415
rect 1072 -421 1075 -415
rect 1079 -421 1082 -415
rect 1086 -421 1089 -415
rect 1093 -421 1096 -415
rect 1100 -421 1103 -415
rect 1107 -421 1110 -415
rect 1114 -421 1117 -415
rect 1121 -421 1124 -415
rect 1128 -421 1131 -415
rect 1135 -421 1138 -415
rect 1142 -421 1145 -415
rect 1149 -421 1152 -415
rect 1156 -421 1159 -415
rect 1163 -421 1166 -415
rect 1170 -421 1173 -415
rect 1177 -421 1180 -415
rect 1184 -421 1187 -415
rect 1191 -421 1194 -415
rect 1198 -421 1201 -415
rect 1205 -421 1208 -415
rect 1212 -421 1215 -415
rect 1219 -421 1225 -415
rect 1387 -421 1390 -415
rect 1408 -421 1411 -415
rect 1520 -421 1523 -415
rect 1 -510 7 -504
rect 8 -510 14 -504
rect 15 -510 21 -504
rect 22 -510 28 -504
rect 29 -510 35 -504
rect 36 -510 42 -504
rect 43 -510 49 -504
rect 50 -510 53 -504
rect 57 -510 60 -504
rect 64 -510 67 -504
rect 71 -510 74 -504
rect 78 -510 81 -504
rect 85 -510 88 -504
rect 92 -510 95 -504
rect 99 -510 102 -504
rect 106 -510 109 -504
rect 113 -510 116 -504
rect 120 -510 126 -504
rect 127 -510 130 -504
rect 134 -510 140 -504
rect 141 -510 147 -504
rect 148 -510 151 -504
rect 155 -510 158 -504
rect 162 -510 168 -504
rect 169 -510 172 -504
rect 176 -510 179 -504
rect 183 -510 186 -504
rect 190 -510 196 -504
rect 197 -510 200 -504
rect 204 -510 207 -504
rect 211 -510 214 -504
rect 218 -510 221 -504
rect 225 -510 228 -504
rect 232 -510 238 -504
rect 239 -510 242 -504
rect 246 -510 249 -504
rect 253 -510 259 -504
rect 260 -510 263 -504
rect 267 -510 270 -504
rect 274 -510 277 -504
rect 281 -510 284 -504
rect 288 -510 291 -504
rect 295 -510 301 -504
rect 302 -510 305 -504
rect 309 -510 312 -504
rect 316 -510 319 -504
rect 323 -510 326 -504
rect 330 -510 333 -504
rect 337 -510 340 -504
rect 344 -510 347 -504
rect 351 -510 354 -504
rect 358 -510 361 -504
rect 365 -510 368 -504
rect 372 -510 375 -504
rect 379 -510 382 -504
rect 386 -510 392 -504
rect 393 -510 396 -504
rect 400 -510 406 -504
rect 407 -510 410 -504
rect 414 -510 417 -504
rect 421 -510 427 -504
rect 428 -510 431 -504
rect 435 -510 438 -504
rect 442 -510 445 -504
rect 449 -510 452 -504
rect 456 -510 459 -504
rect 463 -510 469 -504
rect 470 -510 473 -504
rect 477 -510 480 -504
rect 484 -510 487 -504
rect 491 -510 494 -504
rect 498 -510 501 -504
rect 505 -510 508 -504
rect 512 -510 515 -504
rect 519 -510 522 -504
rect 526 -510 529 -504
rect 533 -510 536 -504
rect 540 -510 543 -504
rect 547 -510 553 -504
rect 554 -510 560 -504
rect 561 -510 564 -504
rect 568 -510 571 -504
rect 575 -510 578 -504
rect 582 -510 585 -504
rect 589 -510 595 -504
rect 596 -510 599 -504
rect 603 -510 606 -504
rect 610 -510 613 -504
rect 617 -510 623 -504
rect 624 -510 627 -504
rect 631 -510 634 -504
rect 638 -510 641 -504
rect 645 -510 651 -504
rect 652 -510 658 -504
rect 659 -510 665 -504
rect 666 -510 669 -504
rect 673 -510 676 -504
rect 680 -510 686 -504
rect 687 -510 690 -504
rect 694 -510 700 -504
rect 701 -510 704 -504
rect 708 -510 711 -504
rect 715 -510 718 -504
rect 722 -510 725 -504
rect 729 -510 732 -504
rect 736 -510 739 -504
rect 743 -510 746 -504
rect 750 -510 756 -504
rect 757 -510 760 -504
rect 764 -510 767 -504
rect 771 -510 774 -504
rect 778 -510 781 -504
rect 785 -510 788 -504
rect 792 -510 795 -504
rect 799 -510 802 -504
rect 806 -510 809 -504
rect 813 -510 816 -504
rect 820 -510 826 -504
rect 827 -510 830 -504
rect 834 -510 837 -504
rect 841 -510 847 -504
rect 848 -510 854 -504
rect 855 -510 858 -504
rect 862 -510 865 -504
rect 869 -510 872 -504
rect 876 -510 879 -504
rect 883 -510 886 -504
rect 890 -510 893 -504
rect 897 -510 900 -504
rect 904 -510 907 -504
rect 911 -510 914 -504
rect 918 -510 921 -504
rect 925 -510 928 -504
rect 932 -510 935 -504
rect 939 -510 942 -504
rect 946 -510 949 -504
rect 953 -510 956 -504
rect 960 -510 963 -504
rect 967 -510 970 -504
rect 974 -510 977 -504
rect 981 -510 984 -504
rect 988 -510 991 -504
rect 995 -510 998 -504
rect 1002 -510 1005 -504
rect 1009 -510 1012 -504
rect 1016 -510 1019 -504
rect 1023 -510 1026 -504
rect 1030 -510 1033 -504
rect 1037 -510 1040 -504
rect 1044 -510 1047 -504
rect 1051 -510 1054 -504
rect 1058 -510 1061 -504
rect 1065 -510 1068 -504
rect 1072 -510 1075 -504
rect 1079 -510 1082 -504
rect 1086 -510 1089 -504
rect 1093 -510 1096 -504
rect 1100 -510 1103 -504
rect 1107 -510 1110 -504
rect 1114 -510 1117 -504
rect 1121 -510 1124 -504
rect 1128 -510 1131 -504
rect 1135 -510 1138 -504
rect 1142 -510 1145 -504
rect 1149 -510 1152 -504
rect 1156 -510 1159 -504
rect 1163 -510 1166 -504
rect 1170 -510 1173 -504
rect 1177 -510 1180 -504
rect 1184 -510 1187 -504
rect 1191 -510 1194 -504
rect 1198 -510 1201 -504
rect 1205 -510 1208 -504
rect 1212 -510 1215 -504
rect 1219 -510 1225 -504
rect 1226 -510 1229 -504
rect 1233 -510 1236 -504
rect 1240 -510 1243 -504
rect 1247 -510 1253 -504
rect 1254 -510 1257 -504
rect 1429 -510 1432 -504
rect 1485 -510 1488 -504
rect 1541 -510 1544 -504
rect 1 -631 7 -625
rect 8 -631 14 -625
rect 15 -631 21 -625
rect 22 -631 28 -625
rect 29 -631 35 -625
rect 36 -631 42 -625
rect 43 -631 46 -625
rect 50 -631 53 -625
rect 57 -631 60 -625
rect 64 -631 67 -625
rect 71 -631 74 -625
rect 78 -631 84 -625
rect 85 -631 88 -625
rect 92 -631 95 -625
rect 99 -631 102 -625
rect 106 -631 112 -625
rect 113 -631 116 -625
rect 120 -631 123 -625
rect 127 -631 130 -625
rect 134 -631 137 -625
rect 141 -631 144 -625
rect 148 -631 151 -625
rect 155 -631 158 -625
rect 162 -631 165 -625
rect 169 -631 172 -625
rect 176 -631 179 -625
rect 183 -631 186 -625
rect 190 -631 193 -625
rect 197 -631 203 -625
rect 204 -631 207 -625
rect 211 -631 214 -625
rect 218 -631 221 -625
rect 225 -631 228 -625
rect 232 -631 238 -625
rect 239 -631 245 -625
rect 246 -631 249 -625
rect 253 -631 256 -625
rect 260 -631 266 -625
rect 267 -631 270 -625
rect 274 -631 277 -625
rect 281 -631 284 -625
rect 288 -631 294 -625
rect 295 -631 298 -625
rect 302 -631 305 -625
rect 309 -631 312 -625
rect 316 -631 319 -625
rect 323 -631 329 -625
rect 330 -631 333 -625
rect 337 -631 340 -625
rect 344 -631 347 -625
rect 351 -631 357 -625
rect 358 -631 361 -625
rect 365 -631 368 -625
rect 372 -631 375 -625
rect 379 -631 382 -625
rect 386 -631 392 -625
rect 393 -631 396 -625
rect 400 -631 403 -625
rect 407 -631 410 -625
rect 414 -631 417 -625
rect 421 -631 427 -625
rect 428 -631 431 -625
rect 435 -631 438 -625
rect 442 -631 445 -625
rect 449 -631 452 -625
rect 456 -631 462 -625
rect 463 -631 466 -625
rect 470 -631 473 -625
rect 477 -631 483 -625
rect 484 -631 487 -625
rect 491 -631 497 -625
rect 498 -631 501 -625
rect 505 -631 508 -625
rect 512 -631 515 -625
rect 519 -631 522 -625
rect 526 -631 529 -625
rect 533 -631 536 -625
rect 540 -631 543 -625
rect 547 -631 550 -625
rect 554 -631 557 -625
rect 561 -631 564 -625
rect 568 -631 571 -625
rect 575 -631 578 -625
rect 582 -631 585 -625
rect 589 -631 592 -625
rect 596 -631 599 -625
rect 603 -631 609 -625
rect 610 -631 613 -625
rect 617 -631 620 -625
rect 624 -631 627 -625
rect 631 -631 634 -625
rect 638 -631 644 -625
rect 645 -631 651 -625
rect 652 -631 655 -625
rect 659 -631 662 -625
rect 666 -631 669 -625
rect 673 -631 676 -625
rect 680 -631 686 -625
rect 687 -631 690 -625
rect 694 -631 700 -625
rect 701 -631 704 -625
rect 708 -631 711 -625
rect 715 -631 718 -625
rect 722 -631 725 -625
rect 729 -631 735 -625
rect 736 -631 739 -625
rect 743 -631 749 -625
rect 750 -631 753 -625
rect 757 -631 763 -625
rect 764 -631 767 -625
rect 771 -631 774 -625
rect 778 -631 781 -625
rect 785 -631 791 -625
rect 792 -631 795 -625
rect 799 -631 805 -625
rect 806 -631 809 -625
rect 813 -631 816 -625
rect 820 -631 823 -625
rect 827 -631 830 -625
rect 834 -631 837 -625
rect 841 -631 847 -625
rect 848 -631 851 -625
rect 855 -631 858 -625
rect 862 -631 865 -625
rect 869 -631 875 -625
rect 876 -631 879 -625
rect 883 -631 886 -625
rect 890 -631 893 -625
rect 897 -631 900 -625
rect 904 -631 907 -625
rect 911 -631 914 -625
rect 918 -631 921 -625
rect 925 -631 928 -625
rect 932 -631 935 -625
rect 939 -631 942 -625
rect 946 -631 949 -625
rect 953 -631 956 -625
rect 960 -631 963 -625
rect 967 -631 970 -625
rect 974 -631 977 -625
rect 981 -631 984 -625
rect 988 -631 991 -625
rect 995 -631 998 -625
rect 1002 -631 1005 -625
rect 1009 -631 1012 -625
rect 1016 -631 1022 -625
rect 1023 -631 1026 -625
rect 1030 -631 1036 -625
rect 1037 -631 1040 -625
rect 1044 -631 1047 -625
rect 1051 -631 1054 -625
rect 1058 -631 1061 -625
rect 1065 -631 1068 -625
rect 1072 -631 1075 -625
rect 1079 -631 1082 -625
rect 1086 -631 1089 -625
rect 1093 -631 1096 -625
rect 1100 -631 1103 -625
rect 1107 -631 1110 -625
rect 1114 -631 1117 -625
rect 1121 -631 1124 -625
rect 1128 -631 1131 -625
rect 1135 -631 1138 -625
rect 1142 -631 1145 -625
rect 1149 -631 1152 -625
rect 1156 -631 1159 -625
rect 1163 -631 1166 -625
rect 1170 -631 1173 -625
rect 1177 -631 1180 -625
rect 1184 -631 1187 -625
rect 1191 -631 1194 -625
rect 1198 -631 1201 -625
rect 1205 -631 1208 -625
rect 1212 -631 1215 -625
rect 1219 -631 1222 -625
rect 1226 -631 1229 -625
rect 1233 -631 1236 -625
rect 1240 -631 1243 -625
rect 1247 -631 1250 -625
rect 1254 -631 1257 -625
rect 1261 -631 1264 -625
rect 1268 -631 1271 -625
rect 1275 -631 1278 -625
rect 1282 -631 1285 -625
rect 1289 -631 1292 -625
rect 1296 -631 1299 -625
rect 1303 -631 1306 -625
rect 1310 -631 1313 -625
rect 1317 -631 1320 -625
rect 1324 -631 1327 -625
rect 1331 -631 1334 -625
rect 1338 -631 1341 -625
rect 1345 -631 1348 -625
rect 1352 -631 1355 -625
rect 1359 -631 1362 -625
rect 1366 -631 1369 -625
rect 1373 -631 1376 -625
rect 1380 -631 1383 -625
rect 1387 -631 1390 -625
rect 1394 -631 1397 -625
rect 1401 -631 1404 -625
rect 1408 -631 1411 -625
rect 1415 -631 1421 -625
rect 1422 -631 1425 -625
rect 1429 -631 1432 -625
rect 1436 -631 1439 -625
rect 1443 -631 1446 -625
rect 1450 -631 1453 -625
rect 1457 -631 1460 -625
rect 1464 -631 1467 -625
rect 1527 -631 1530 -625
rect 1548 -631 1551 -625
rect 1618 -631 1621 -625
rect 1 -764 7 -758
rect 8 -764 14 -758
rect 15 -764 21 -758
rect 22 -764 28 -758
rect 29 -764 35 -758
rect 36 -764 42 -758
rect 43 -764 46 -758
rect 50 -764 53 -758
rect 57 -764 63 -758
rect 64 -764 70 -758
rect 71 -764 74 -758
rect 78 -764 81 -758
rect 85 -764 88 -758
rect 92 -764 95 -758
rect 99 -764 102 -758
rect 106 -764 109 -758
rect 113 -764 119 -758
rect 120 -764 123 -758
rect 127 -764 130 -758
rect 134 -764 137 -758
rect 141 -764 144 -758
rect 148 -764 151 -758
rect 155 -764 161 -758
rect 162 -764 165 -758
rect 169 -764 172 -758
rect 176 -764 179 -758
rect 183 -764 186 -758
rect 190 -764 193 -758
rect 197 -764 200 -758
rect 204 -764 210 -758
rect 211 -764 214 -758
rect 218 -764 224 -758
rect 225 -764 228 -758
rect 232 -764 235 -758
rect 239 -764 242 -758
rect 246 -764 249 -758
rect 253 -764 259 -758
rect 260 -764 263 -758
rect 267 -764 270 -758
rect 274 -764 277 -758
rect 281 -764 284 -758
rect 288 -764 291 -758
rect 295 -764 298 -758
rect 302 -764 305 -758
rect 309 -764 312 -758
rect 316 -764 319 -758
rect 323 -764 326 -758
rect 330 -764 336 -758
rect 337 -764 340 -758
rect 344 -764 347 -758
rect 351 -764 354 -758
rect 358 -764 361 -758
rect 365 -764 368 -758
rect 372 -764 375 -758
rect 379 -764 382 -758
rect 386 -764 389 -758
rect 393 -764 396 -758
rect 400 -764 403 -758
rect 407 -764 410 -758
rect 414 -764 417 -758
rect 421 -764 424 -758
rect 428 -764 434 -758
rect 435 -764 438 -758
rect 442 -764 445 -758
rect 449 -764 452 -758
rect 456 -764 459 -758
rect 463 -764 469 -758
rect 470 -764 473 -758
rect 477 -764 480 -758
rect 484 -764 487 -758
rect 491 -764 497 -758
rect 498 -764 501 -758
rect 505 -764 508 -758
rect 512 -764 515 -758
rect 519 -764 525 -758
rect 526 -764 532 -758
rect 533 -764 536 -758
rect 540 -764 543 -758
rect 547 -764 550 -758
rect 554 -764 560 -758
rect 561 -764 564 -758
rect 568 -764 574 -758
rect 575 -764 578 -758
rect 582 -764 585 -758
rect 589 -764 592 -758
rect 596 -764 599 -758
rect 603 -764 609 -758
rect 610 -764 613 -758
rect 617 -764 620 -758
rect 624 -764 627 -758
rect 631 -764 637 -758
rect 638 -764 641 -758
rect 645 -764 651 -758
rect 652 -764 655 -758
rect 659 -764 662 -758
rect 666 -764 669 -758
rect 673 -764 679 -758
rect 680 -764 683 -758
rect 687 -764 693 -758
rect 694 -764 697 -758
rect 701 -764 704 -758
rect 708 -764 711 -758
rect 715 -764 721 -758
rect 722 -764 725 -758
rect 729 -764 735 -758
rect 736 -764 739 -758
rect 743 -764 746 -758
rect 750 -764 753 -758
rect 757 -764 760 -758
rect 764 -764 767 -758
rect 771 -764 774 -758
rect 778 -764 781 -758
rect 785 -764 788 -758
rect 792 -764 798 -758
rect 799 -764 805 -758
rect 806 -764 809 -758
rect 813 -764 816 -758
rect 820 -764 823 -758
rect 827 -764 833 -758
rect 834 -764 840 -758
rect 841 -764 844 -758
rect 848 -764 851 -758
rect 855 -764 858 -758
rect 862 -764 865 -758
rect 869 -764 875 -758
rect 876 -764 879 -758
rect 883 -764 886 -758
rect 890 -764 893 -758
rect 897 -764 900 -758
rect 904 -764 910 -758
rect 911 -764 914 -758
rect 918 -764 921 -758
rect 925 -764 931 -758
rect 932 -764 935 -758
rect 939 -764 942 -758
rect 946 -764 949 -758
rect 953 -764 956 -758
rect 960 -764 963 -758
rect 967 -764 970 -758
rect 974 -764 977 -758
rect 981 -764 984 -758
rect 988 -764 991 -758
rect 995 -764 998 -758
rect 1002 -764 1005 -758
rect 1009 -764 1012 -758
rect 1016 -764 1019 -758
rect 1023 -764 1029 -758
rect 1030 -764 1033 -758
rect 1037 -764 1040 -758
rect 1044 -764 1047 -758
rect 1051 -764 1054 -758
rect 1058 -764 1061 -758
rect 1065 -764 1068 -758
rect 1072 -764 1075 -758
rect 1079 -764 1082 -758
rect 1086 -764 1089 -758
rect 1093 -764 1096 -758
rect 1100 -764 1103 -758
rect 1107 -764 1110 -758
rect 1114 -764 1117 -758
rect 1121 -764 1124 -758
rect 1128 -764 1131 -758
rect 1135 -764 1138 -758
rect 1142 -764 1145 -758
rect 1149 -764 1152 -758
rect 1156 -764 1159 -758
rect 1163 -764 1166 -758
rect 1170 -764 1173 -758
rect 1177 -764 1180 -758
rect 1184 -764 1187 -758
rect 1191 -764 1194 -758
rect 1198 -764 1201 -758
rect 1205 -764 1208 -758
rect 1212 -764 1215 -758
rect 1219 -764 1222 -758
rect 1226 -764 1229 -758
rect 1233 -764 1236 -758
rect 1240 -764 1243 -758
rect 1247 -764 1250 -758
rect 1254 -764 1257 -758
rect 1261 -764 1264 -758
rect 1268 -764 1271 -758
rect 1275 -764 1278 -758
rect 1282 -764 1285 -758
rect 1289 -764 1292 -758
rect 1296 -764 1299 -758
rect 1303 -764 1306 -758
rect 1310 -764 1313 -758
rect 1317 -764 1320 -758
rect 1324 -764 1327 -758
rect 1331 -764 1334 -758
rect 1338 -764 1341 -758
rect 1345 -764 1348 -758
rect 1352 -764 1355 -758
rect 1359 -764 1362 -758
rect 1366 -764 1369 -758
rect 1373 -764 1376 -758
rect 1380 -764 1383 -758
rect 1387 -764 1390 -758
rect 1394 -764 1397 -758
rect 1401 -764 1404 -758
rect 1408 -764 1411 -758
rect 1415 -764 1418 -758
rect 1422 -764 1425 -758
rect 1429 -764 1432 -758
rect 1436 -764 1439 -758
rect 1443 -764 1446 -758
rect 1450 -764 1453 -758
rect 1457 -764 1460 -758
rect 1464 -764 1467 -758
rect 1471 -764 1474 -758
rect 1478 -764 1481 -758
rect 1485 -764 1488 -758
rect 1527 -764 1530 -758
rect 1548 -764 1551 -758
rect 1555 -764 1558 -758
rect 1695 -764 1698 -758
rect 1 -877 7 -871
rect 8 -877 14 -871
rect 15 -877 21 -871
rect 22 -877 28 -871
rect 29 -877 35 -871
rect 36 -877 39 -871
rect 43 -877 46 -871
rect 50 -877 53 -871
rect 57 -877 60 -871
rect 64 -877 67 -871
rect 71 -877 74 -871
rect 78 -877 81 -871
rect 85 -877 88 -871
rect 92 -877 95 -871
rect 99 -877 102 -871
rect 106 -877 112 -871
rect 113 -877 116 -871
rect 120 -877 126 -871
rect 127 -877 130 -871
rect 134 -877 137 -871
rect 141 -877 144 -871
rect 148 -877 154 -871
rect 155 -877 158 -871
rect 162 -877 168 -871
rect 169 -877 172 -871
rect 176 -877 179 -871
rect 183 -877 189 -871
rect 190 -877 193 -871
rect 197 -877 200 -871
rect 204 -877 210 -871
rect 211 -877 214 -871
rect 218 -877 224 -871
rect 225 -877 228 -871
rect 232 -877 235 -871
rect 239 -877 242 -871
rect 246 -877 249 -871
rect 253 -877 259 -871
rect 260 -877 263 -871
rect 267 -877 270 -871
rect 274 -877 277 -871
rect 281 -877 284 -871
rect 288 -877 291 -871
rect 295 -877 298 -871
rect 302 -877 305 -871
rect 309 -877 312 -871
rect 316 -877 319 -871
rect 323 -877 326 -871
rect 330 -877 333 -871
rect 337 -877 340 -871
rect 344 -877 347 -871
rect 351 -877 354 -871
rect 358 -877 361 -871
rect 365 -877 368 -871
rect 372 -877 375 -871
rect 379 -877 382 -871
rect 386 -877 389 -871
rect 393 -877 396 -871
rect 400 -877 403 -871
rect 407 -877 413 -871
rect 414 -877 417 -871
rect 421 -877 424 -871
rect 428 -877 431 -871
rect 435 -877 438 -871
rect 442 -877 445 -871
rect 449 -877 452 -871
rect 456 -877 459 -871
rect 463 -877 466 -871
rect 470 -877 473 -871
rect 477 -877 480 -871
rect 484 -877 487 -871
rect 491 -877 494 -871
rect 498 -877 504 -871
rect 505 -877 511 -871
rect 512 -877 515 -871
rect 519 -877 525 -871
rect 526 -877 532 -871
rect 533 -877 539 -871
rect 540 -877 543 -871
rect 547 -877 553 -871
rect 554 -877 557 -871
rect 561 -877 564 -871
rect 568 -877 571 -871
rect 575 -877 578 -871
rect 582 -877 585 -871
rect 589 -877 592 -871
rect 596 -877 599 -871
rect 603 -877 606 -871
rect 610 -877 613 -871
rect 617 -877 620 -871
rect 624 -877 630 -871
rect 631 -877 634 -871
rect 638 -877 641 -871
rect 645 -877 651 -871
rect 652 -877 655 -871
rect 659 -877 662 -871
rect 666 -877 672 -871
rect 673 -877 679 -871
rect 680 -877 686 -871
rect 687 -877 690 -871
rect 694 -877 697 -871
rect 701 -877 704 -871
rect 708 -877 711 -871
rect 715 -877 718 -871
rect 722 -877 725 -871
rect 729 -877 732 -871
rect 736 -877 739 -871
rect 743 -877 746 -871
rect 750 -877 753 -871
rect 757 -877 760 -871
rect 764 -877 767 -871
rect 771 -877 774 -871
rect 778 -877 784 -871
rect 785 -877 788 -871
rect 792 -877 795 -871
rect 799 -877 802 -871
rect 806 -877 809 -871
rect 813 -877 819 -871
rect 820 -877 823 -871
rect 827 -877 833 -871
rect 834 -877 840 -871
rect 841 -877 844 -871
rect 848 -877 851 -871
rect 855 -877 858 -871
rect 862 -877 865 -871
rect 869 -877 875 -871
rect 876 -877 882 -871
rect 883 -877 886 -871
rect 890 -877 893 -871
rect 897 -877 900 -871
rect 904 -877 907 -871
rect 911 -877 914 -871
rect 918 -877 924 -871
rect 925 -877 928 -871
rect 932 -877 935 -871
rect 939 -877 942 -871
rect 946 -877 949 -871
rect 953 -877 956 -871
rect 960 -877 966 -871
rect 967 -877 970 -871
rect 974 -877 977 -871
rect 981 -877 984 -871
rect 988 -877 991 -871
rect 995 -877 998 -871
rect 1002 -877 1005 -871
rect 1009 -877 1012 -871
rect 1016 -877 1019 -871
rect 1023 -877 1026 -871
rect 1030 -877 1033 -871
rect 1037 -877 1040 -871
rect 1044 -877 1047 -871
rect 1051 -877 1054 -871
rect 1058 -877 1061 -871
rect 1065 -877 1071 -871
rect 1072 -877 1075 -871
rect 1079 -877 1082 -871
rect 1086 -877 1089 -871
rect 1093 -877 1096 -871
rect 1100 -877 1103 -871
rect 1107 -877 1110 -871
rect 1114 -877 1117 -871
rect 1121 -877 1124 -871
rect 1128 -877 1131 -871
rect 1135 -877 1138 -871
rect 1142 -877 1145 -871
rect 1149 -877 1152 -871
rect 1156 -877 1159 -871
rect 1163 -877 1166 -871
rect 1170 -877 1173 -871
rect 1177 -877 1180 -871
rect 1184 -877 1187 -871
rect 1191 -877 1194 -871
rect 1198 -877 1201 -871
rect 1205 -877 1208 -871
rect 1212 -877 1215 -871
rect 1219 -877 1222 -871
rect 1226 -877 1229 -871
rect 1233 -877 1236 -871
rect 1240 -877 1243 -871
rect 1247 -877 1250 -871
rect 1254 -877 1257 -871
rect 1261 -877 1264 -871
rect 1268 -877 1271 -871
rect 1275 -877 1278 -871
rect 1282 -877 1285 -871
rect 1289 -877 1292 -871
rect 1296 -877 1299 -871
rect 1303 -877 1306 -871
rect 1310 -877 1313 -871
rect 1317 -877 1320 -871
rect 1324 -877 1327 -871
rect 1331 -877 1334 -871
rect 1338 -877 1341 -871
rect 1345 -877 1348 -871
rect 1352 -877 1355 -871
rect 1359 -877 1362 -871
rect 1366 -877 1369 -871
rect 1373 -877 1376 -871
rect 1380 -877 1383 -871
rect 1387 -877 1390 -871
rect 1394 -877 1397 -871
rect 1401 -877 1404 -871
rect 1408 -877 1411 -871
rect 1415 -877 1418 -871
rect 1422 -877 1425 -871
rect 1429 -877 1432 -871
rect 1436 -877 1439 -871
rect 1443 -877 1446 -871
rect 1450 -877 1453 -871
rect 1457 -877 1460 -871
rect 1464 -877 1467 -871
rect 1471 -877 1474 -871
rect 1478 -877 1481 -871
rect 1485 -877 1488 -871
rect 1492 -877 1495 -871
rect 1499 -877 1502 -871
rect 1506 -877 1509 -871
rect 1513 -877 1516 -871
rect 1520 -877 1523 -871
rect 1527 -877 1530 -871
rect 1534 -877 1537 -871
rect 1541 -877 1544 -871
rect 1548 -877 1551 -871
rect 1555 -877 1561 -871
rect 1562 -877 1568 -871
rect 1569 -877 1572 -871
rect 1576 -877 1579 -871
rect 1583 -877 1586 -871
rect 1723 -877 1726 -871
rect 1 -1004 7 -998
rect 8 -1004 14 -998
rect 15 -1004 21 -998
rect 22 -1004 28 -998
rect 29 -1004 32 -998
rect 36 -1004 39 -998
rect 43 -1004 46 -998
rect 50 -1004 53 -998
rect 57 -1004 60 -998
rect 64 -1004 67 -998
rect 71 -1004 74 -998
rect 78 -1004 84 -998
rect 85 -1004 88 -998
rect 92 -1004 95 -998
rect 99 -1004 102 -998
rect 106 -1004 109 -998
rect 113 -1004 116 -998
rect 120 -1004 123 -998
rect 127 -1004 133 -998
rect 134 -1004 140 -998
rect 141 -1004 144 -998
rect 148 -1004 154 -998
rect 155 -1004 158 -998
rect 162 -1004 165 -998
rect 169 -1004 172 -998
rect 176 -1004 179 -998
rect 183 -1004 186 -998
rect 190 -1004 193 -998
rect 197 -1004 200 -998
rect 204 -1004 207 -998
rect 211 -1004 214 -998
rect 218 -1004 221 -998
rect 225 -1004 228 -998
rect 232 -1004 235 -998
rect 239 -1004 242 -998
rect 246 -1004 252 -998
rect 253 -1004 256 -998
rect 260 -1004 263 -998
rect 267 -1004 270 -998
rect 274 -1004 277 -998
rect 281 -1004 284 -998
rect 288 -1004 291 -998
rect 295 -1004 298 -998
rect 302 -1004 305 -998
rect 309 -1004 312 -998
rect 316 -1004 319 -998
rect 323 -1004 326 -998
rect 330 -1004 333 -998
rect 337 -1004 340 -998
rect 344 -1004 347 -998
rect 351 -1004 354 -998
rect 358 -1004 361 -998
rect 365 -1004 368 -998
rect 372 -1004 375 -998
rect 379 -1004 382 -998
rect 386 -1004 389 -998
rect 393 -1004 396 -998
rect 400 -1004 403 -998
rect 407 -1004 410 -998
rect 414 -1004 417 -998
rect 421 -1004 427 -998
rect 428 -1004 431 -998
rect 435 -1004 438 -998
rect 442 -1004 448 -998
rect 449 -1004 452 -998
rect 456 -1004 459 -998
rect 463 -1004 466 -998
rect 470 -1004 473 -998
rect 477 -1004 480 -998
rect 484 -1004 487 -998
rect 491 -1004 494 -998
rect 498 -1004 504 -998
rect 505 -1004 511 -998
rect 512 -1004 515 -998
rect 519 -1004 522 -998
rect 526 -1004 529 -998
rect 533 -1004 536 -998
rect 540 -1004 543 -998
rect 547 -1004 550 -998
rect 554 -1004 557 -998
rect 561 -1004 564 -998
rect 568 -1004 571 -998
rect 575 -1004 578 -998
rect 582 -1004 588 -998
rect 589 -1004 592 -998
rect 596 -1004 599 -998
rect 603 -1004 606 -998
rect 610 -1004 613 -998
rect 617 -1004 623 -998
rect 624 -1004 627 -998
rect 631 -1004 634 -998
rect 638 -1004 644 -998
rect 645 -1004 651 -998
rect 652 -1004 658 -998
rect 659 -1004 662 -998
rect 666 -1004 669 -998
rect 673 -1004 676 -998
rect 680 -1004 686 -998
rect 687 -1004 693 -998
rect 694 -1004 700 -998
rect 701 -1004 704 -998
rect 708 -1004 711 -998
rect 715 -1004 718 -998
rect 722 -1004 725 -998
rect 729 -1004 735 -998
rect 736 -1004 739 -998
rect 743 -1004 746 -998
rect 750 -1004 753 -998
rect 757 -1004 760 -998
rect 764 -1004 770 -998
rect 771 -1004 777 -998
rect 778 -1004 781 -998
rect 785 -1004 788 -998
rect 792 -1004 795 -998
rect 799 -1004 802 -998
rect 806 -1004 809 -998
rect 813 -1004 816 -998
rect 820 -1004 823 -998
rect 827 -1004 830 -998
rect 834 -1004 837 -998
rect 841 -1004 847 -998
rect 848 -1004 851 -998
rect 855 -1004 858 -998
rect 862 -1004 865 -998
rect 869 -1004 872 -998
rect 876 -1004 879 -998
rect 883 -1004 889 -998
rect 890 -1004 893 -998
rect 897 -1004 903 -998
rect 904 -1004 907 -998
rect 911 -1004 914 -998
rect 918 -1004 921 -998
rect 925 -1004 928 -998
rect 932 -1004 935 -998
rect 939 -1004 942 -998
rect 946 -1004 949 -998
rect 953 -1004 956 -998
rect 960 -1004 966 -998
rect 967 -1004 970 -998
rect 974 -1004 980 -998
rect 981 -1004 987 -998
rect 988 -1004 994 -998
rect 995 -1004 1001 -998
rect 1002 -1004 1005 -998
rect 1009 -1004 1015 -998
rect 1016 -1004 1019 -998
rect 1023 -1004 1026 -998
rect 1030 -1004 1033 -998
rect 1037 -1004 1040 -998
rect 1044 -1004 1047 -998
rect 1051 -1004 1054 -998
rect 1058 -1004 1061 -998
rect 1065 -1004 1068 -998
rect 1072 -1004 1075 -998
rect 1079 -1004 1082 -998
rect 1086 -1004 1089 -998
rect 1093 -1004 1096 -998
rect 1100 -1004 1103 -998
rect 1107 -1004 1113 -998
rect 1114 -1004 1117 -998
rect 1121 -1004 1124 -998
rect 1128 -1004 1131 -998
rect 1135 -1004 1138 -998
rect 1142 -1004 1145 -998
rect 1149 -1004 1152 -998
rect 1156 -1004 1159 -998
rect 1163 -1004 1166 -998
rect 1170 -1004 1173 -998
rect 1177 -1004 1180 -998
rect 1184 -1004 1187 -998
rect 1191 -1004 1194 -998
rect 1198 -1004 1201 -998
rect 1205 -1004 1208 -998
rect 1212 -1004 1215 -998
rect 1219 -1004 1222 -998
rect 1226 -1004 1229 -998
rect 1233 -1004 1236 -998
rect 1240 -1004 1243 -998
rect 1247 -1004 1250 -998
rect 1254 -1004 1257 -998
rect 1261 -1004 1264 -998
rect 1268 -1004 1271 -998
rect 1275 -1004 1278 -998
rect 1282 -1004 1285 -998
rect 1289 -1004 1292 -998
rect 1296 -1004 1299 -998
rect 1303 -1004 1306 -998
rect 1310 -1004 1313 -998
rect 1317 -1004 1320 -998
rect 1324 -1004 1327 -998
rect 1331 -1004 1334 -998
rect 1338 -1004 1341 -998
rect 1345 -1004 1348 -998
rect 1352 -1004 1355 -998
rect 1359 -1004 1362 -998
rect 1366 -1004 1369 -998
rect 1373 -1004 1376 -998
rect 1380 -1004 1383 -998
rect 1387 -1004 1390 -998
rect 1394 -1004 1397 -998
rect 1401 -1004 1404 -998
rect 1408 -1004 1411 -998
rect 1415 -1004 1418 -998
rect 1422 -1004 1425 -998
rect 1429 -1004 1432 -998
rect 1436 -1004 1439 -998
rect 1443 -1004 1446 -998
rect 1450 -1004 1453 -998
rect 1457 -1004 1460 -998
rect 1464 -1004 1467 -998
rect 1471 -1004 1474 -998
rect 1478 -1004 1481 -998
rect 1485 -1004 1488 -998
rect 1492 -1004 1495 -998
rect 1499 -1004 1502 -998
rect 1506 -1004 1509 -998
rect 1513 -1004 1516 -998
rect 1520 -1004 1523 -998
rect 1527 -1004 1530 -998
rect 1534 -1004 1537 -998
rect 1541 -1004 1544 -998
rect 1548 -1004 1554 -998
rect 1555 -1004 1558 -998
rect 1562 -1004 1568 -998
rect 1569 -1004 1575 -998
rect 1576 -1004 1579 -998
rect 1583 -1004 1586 -998
rect 1590 -1004 1593 -998
rect 1597 -1004 1600 -998
rect 1604 -1004 1607 -998
rect 1611 -1004 1614 -998
rect 1618 -1004 1621 -998
rect 1625 -1004 1628 -998
rect 1632 -1004 1635 -998
rect 1737 -1004 1740 -998
rect 1 -1105 7 -1099
rect 8 -1105 14 -1099
rect 15 -1105 21 -1099
rect 22 -1105 25 -1099
rect 29 -1105 32 -1099
rect 36 -1105 42 -1099
rect 43 -1105 46 -1099
rect 50 -1105 53 -1099
rect 57 -1105 60 -1099
rect 64 -1105 67 -1099
rect 71 -1105 77 -1099
rect 78 -1105 81 -1099
rect 85 -1105 91 -1099
rect 92 -1105 95 -1099
rect 99 -1105 102 -1099
rect 106 -1105 109 -1099
rect 113 -1105 116 -1099
rect 120 -1105 123 -1099
rect 127 -1105 130 -1099
rect 134 -1105 140 -1099
rect 141 -1105 144 -1099
rect 148 -1105 151 -1099
rect 155 -1105 158 -1099
rect 162 -1105 165 -1099
rect 169 -1105 172 -1099
rect 176 -1105 179 -1099
rect 183 -1105 186 -1099
rect 190 -1105 193 -1099
rect 197 -1105 200 -1099
rect 204 -1105 207 -1099
rect 211 -1105 217 -1099
rect 218 -1105 221 -1099
rect 225 -1105 228 -1099
rect 232 -1105 238 -1099
rect 239 -1105 242 -1099
rect 246 -1105 252 -1099
rect 253 -1105 256 -1099
rect 260 -1105 266 -1099
rect 267 -1105 270 -1099
rect 274 -1105 277 -1099
rect 281 -1105 284 -1099
rect 288 -1105 291 -1099
rect 295 -1105 298 -1099
rect 302 -1105 305 -1099
rect 309 -1105 312 -1099
rect 316 -1105 319 -1099
rect 323 -1105 326 -1099
rect 330 -1105 333 -1099
rect 337 -1105 343 -1099
rect 344 -1105 347 -1099
rect 351 -1105 354 -1099
rect 358 -1105 361 -1099
rect 365 -1105 368 -1099
rect 372 -1105 375 -1099
rect 379 -1105 382 -1099
rect 386 -1105 389 -1099
rect 393 -1105 399 -1099
rect 400 -1105 403 -1099
rect 407 -1105 410 -1099
rect 414 -1105 417 -1099
rect 421 -1105 427 -1099
rect 428 -1105 431 -1099
rect 435 -1105 438 -1099
rect 442 -1105 445 -1099
rect 449 -1105 452 -1099
rect 456 -1105 459 -1099
rect 463 -1105 466 -1099
rect 470 -1105 476 -1099
rect 477 -1105 483 -1099
rect 484 -1105 487 -1099
rect 491 -1105 494 -1099
rect 498 -1105 501 -1099
rect 505 -1105 508 -1099
rect 512 -1105 518 -1099
rect 519 -1105 522 -1099
rect 526 -1105 529 -1099
rect 533 -1105 536 -1099
rect 540 -1105 543 -1099
rect 547 -1105 550 -1099
rect 554 -1105 557 -1099
rect 561 -1105 564 -1099
rect 568 -1105 571 -1099
rect 575 -1105 578 -1099
rect 582 -1105 585 -1099
rect 589 -1105 592 -1099
rect 596 -1105 599 -1099
rect 603 -1105 606 -1099
rect 610 -1105 613 -1099
rect 617 -1105 620 -1099
rect 624 -1105 630 -1099
rect 631 -1105 634 -1099
rect 638 -1105 644 -1099
rect 645 -1105 651 -1099
rect 652 -1105 655 -1099
rect 659 -1105 662 -1099
rect 666 -1105 669 -1099
rect 673 -1105 679 -1099
rect 680 -1105 683 -1099
rect 687 -1105 693 -1099
rect 694 -1105 700 -1099
rect 701 -1105 704 -1099
rect 708 -1105 711 -1099
rect 715 -1105 718 -1099
rect 722 -1105 725 -1099
rect 729 -1105 735 -1099
rect 736 -1105 739 -1099
rect 743 -1105 746 -1099
rect 750 -1105 753 -1099
rect 757 -1105 760 -1099
rect 764 -1105 767 -1099
rect 771 -1105 774 -1099
rect 778 -1105 781 -1099
rect 785 -1105 788 -1099
rect 792 -1105 795 -1099
rect 799 -1105 805 -1099
rect 806 -1105 809 -1099
rect 813 -1105 816 -1099
rect 820 -1105 823 -1099
rect 827 -1105 830 -1099
rect 834 -1105 837 -1099
rect 841 -1105 844 -1099
rect 848 -1105 851 -1099
rect 855 -1105 858 -1099
rect 862 -1105 868 -1099
rect 869 -1105 872 -1099
rect 876 -1105 882 -1099
rect 883 -1105 889 -1099
rect 890 -1105 896 -1099
rect 897 -1105 900 -1099
rect 904 -1105 907 -1099
rect 911 -1105 914 -1099
rect 918 -1105 921 -1099
rect 925 -1105 928 -1099
rect 932 -1105 935 -1099
rect 939 -1105 942 -1099
rect 946 -1105 949 -1099
rect 953 -1105 956 -1099
rect 960 -1105 963 -1099
rect 967 -1105 970 -1099
rect 974 -1105 977 -1099
rect 981 -1105 984 -1099
rect 988 -1105 991 -1099
rect 995 -1105 998 -1099
rect 1002 -1105 1008 -1099
rect 1009 -1105 1012 -1099
rect 1016 -1105 1019 -1099
rect 1023 -1105 1026 -1099
rect 1030 -1105 1033 -1099
rect 1037 -1105 1040 -1099
rect 1044 -1105 1050 -1099
rect 1051 -1105 1057 -1099
rect 1058 -1105 1061 -1099
rect 1065 -1105 1068 -1099
rect 1072 -1105 1075 -1099
rect 1079 -1105 1082 -1099
rect 1086 -1105 1092 -1099
rect 1093 -1105 1096 -1099
rect 1100 -1105 1103 -1099
rect 1107 -1105 1110 -1099
rect 1114 -1105 1117 -1099
rect 1121 -1105 1124 -1099
rect 1128 -1105 1131 -1099
rect 1135 -1105 1138 -1099
rect 1142 -1105 1145 -1099
rect 1149 -1105 1152 -1099
rect 1156 -1105 1159 -1099
rect 1163 -1105 1166 -1099
rect 1170 -1105 1173 -1099
rect 1177 -1105 1180 -1099
rect 1184 -1105 1187 -1099
rect 1191 -1105 1194 -1099
rect 1198 -1105 1201 -1099
rect 1205 -1105 1208 -1099
rect 1212 -1105 1215 -1099
rect 1219 -1105 1225 -1099
rect 1226 -1105 1229 -1099
rect 1233 -1105 1236 -1099
rect 1240 -1105 1243 -1099
rect 1247 -1105 1250 -1099
rect 1254 -1105 1257 -1099
rect 1261 -1105 1264 -1099
rect 1268 -1105 1271 -1099
rect 1275 -1105 1278 -1099
rect 1282 -1105 1285 -1099
rect 1289 -1105 1292 -1099
rect 1296 -1105 1299 -1099
rect 1303 -1105 1306 -1099
rect 1310 -1105 1313 -1099
rect 1317 -1105 1320 -1099
rect 1324 -1105 1327 -1099
rect 1331 -1105 1334 -1099
rect 1338 -1105 1341 -1099
rect 1345 -1105 1348 -1099
rect 1352 -1105 1355 -1099
rect 1359 -1105 1362 -1099
rect 1366 -1105 1369 -1099
rect 1373 -1105 1376 -1099
rect 1380 -1105 1386 -1099
rect 1387 -1105 1390 -1099
rect 1394 -1105 1397 -1099
rect 1401 -1105 1404 -1099
rect 1408 -1105 1411 -1099
rect 1415 -1105 1418 -1099
rect 1422 -1105 1425 -1099
rect 1429 -1105 1432 -1099
rect 1436 -1105 1439 -1099
rect 1443 -1105 1446 -1099
rect 1450 -1105 1456 -1099
rect 1457 -1105 1460 -1099
rect 1464 -1105 1467 -1099
rect 1471 -1105 1477 -1099
rect 1478 -1105 1481 -1099
rect 1485 -1105 1488 -1099
rect 1492 -1105 1498 -1099
rect 1499 -1105 1502 -1099
rect 1506 -1105 1509 -1099
rect 1513 -1105 1516 -1099
rect 1520 -1105 1523 -1099
rect 1527 -1105 1530 -1099
rect 1534 -1105 1537 -1099
rect 1541 -1105 1544 -1099
rect 1548 -1105 1551 -1099
rect 1555 -1105 1558 -1099
rect 1562 -1105 1565 -1099
rect 1569 -1105 1572 -1099
rect 1576 -1105 1579 -1099
rect 1583 -1105 1586 -1099
rect 1590 -1105 1593 -1099
rect 1597 -1105 1600 -1099
rect 1604 -1105 1607 -1099
rect 1611 -1105 1614 -1099
rect 1618 -1105 1621 -1099
rect 1625 -1105 1628 -1099
rect 1632 -1105 1635 -1099
rect 1639 -1105 1642 -1099
rect 1646 -1105 1649 -1099
rect 1653 -1105 1656 -1099
rect 1674 -1105 1677 -1099
rect 1681 -1105 1684 -1099
rect 1744 -1105 1747 -1099
rect 1 -1224 7 -1218
rect 8 -1224 14 -1218
rect 15 -1224 21 -1218
rect 22 -1224 25 -1218
rect 29 -1224 32 -1218
rect 36 -1224 39 -1218
rect 43 -1224 46 -1218
rect 50 -1224 53 -1218
rect 57 -1224 60 -1218
rect 64 -1224 70 -1218
rect 71 -1224 74 -1218
rect 78 -1224 81 -1218
rect 85 -1224 91 -1218
rect 92 -1224 95 -1218
rect 99 -1224 102 -1218
rect 106 -1224 112 -1218
rect 113 -1224 116 -1218
rect 120 -1224 126 -1218
rect 127 -1224 130 -1218
rect 134 -1224 137 -1218
rect 141 -1224 147 -1218
rect 148 -1224 151 -1218
rect 155 -1224 158 -1218
rect 162 -1224 165 -1218
rect 169 -1224 175 -1218
rect 176 -1224 182 -1218
rect 183 -1224 186 -1218
rect 190 -1224 193 -1218
rect 197 -1224 200 -1218
rect 204 -1224 207 -1218
rect 211 -1224 214 -1218
rect 218 -1224 221 -1218
rect 225 -1224 231 -1218
rect 232 -1224 235 -1218
rect 239 -1224 245 -1218
rect 246 -1224 249 -1218
rect 253 -1224 256 -1218
rect 260 -1224 266 -1218
rect 267 -1224 270 -1218
rect 274 -1224 277 -1218
rect 281 -1224 284 -1218
rect 288 -1224 291 -1218
rect 295 -1224 298 -1218
rect 302 -1224 305 -1218
rect 309 -1224 312 -1218
rect 316 -1224 319 -1218
rect 323 -1224 326 -1218
rect 330 -1224 333 -1218
rect 337 -1224 340 -1218
rect 344 -1224 347 -1218
rect 351 -1224 354 -1218
rect 358 -1224 361 -1218
rect 365 -1224 368 -1218
rect 372 -1224 375 -1218
rect 379 -1224 382 -1218
rect 386 -1224 389 -1218
rect 393 -1224 396 -1218
rect 400 -1224 403 -1218
rect 407 -1224 410 -1218
rect 414 -1224 417 -1218
rect 421 -1224 424 -1218
rect 428 -1224 431 -1218
rect 435 -1224 441 -1218
rect 442 -1224 445 -1218
rect 449 -1224 452 -1218
rect 456 -1224 459 -1218
rect 463 -1224 466 -1218
rect 470 -1224 473 -1218
rect 477 -1224 480 -1218
rect 484 -1224 487 -1218
rect 491 -1224 494 -1218
rect 498 -1224 501 -1218
rect 505 -1224 511 -1218
rect 512 -1224 515 -1218
rect 519 -1224 522 -1218
rect 526 -1224 529 -1218
rect 533 -1224 536 -1218
rect 540 -1224 546 -1218
rect 547 -1224 550 -1218
rect 554 -1224 557 -1218
rect 561 -1224 567 -1218
rect 568 -1224 571 -1218
rect 575 -1224 578 -1218
rect 582 -1224 585 -1218
rect 589 -1224 592 -1218
rect 596 -1224 602 -1218
rect 603 -1224 609 -1218
rect 610 -1224 613 -1218
rect 617 -1224 620 -1218
rect 624 -1224 627 -1218
rect 631 -1224 637 -1218
rect 638 -1224 641 -1218
rect 645 -1224 651 -1218
rect 652 -1224 658 -1218
rect 659 -1224 662 -1218
rect 666 -1224 669 -1218
rect 673 -1224 676 -1218
rect 680 -1224 683 -1218
rect 687 -1224 690 -1218
rect 694 -1224 700 -1218
rect 701 -1224 707 -1218
rect 708 -1224 711 -1218
rect 715 -1224 718 -1218
rect 722 -1224 725 -1218
rect 729 -1224 732 -1218
rect 736 -1224 742 -1218
rect 743 -1224 746 -1218
rect 750 -1224 753 -1218
rect 757 -1224 760 -1218
rect 764 -1224 770 -1218
rect 771 -1224 774 -1218
rect 778 -1224 781 -1218
rect 785 -1224 788 -1218
rect 792 -1224 798 -1218
rect 799 -1224 802 -1218
rect 806 -1224 809 -1218
rect 813 -1224 819 -1218
rect 820 -1224 826 -1218
rect 827 -1224 833 -1218
rect 834 -1224 837 -1218
rect 841 -1224 844 -1218
rect 848 -1224 851 -1218
rect 855 -1224 861 -1218
rect 862 -1224 865 -1218
rect 869 -1224 872 -1218
rect 876 -1224 879 -1218
rect 883 -1224 886 -1218
rect 890 -1224 896 -1218
rect 897 -1224 900 -1218
rect 904 -1224 907 -1218
rect 911 -1224 914 -1218
rect 918 -1224 921 -1218
rect 925 -1224 931 -1218
rect 932 -1224 935 -1218
rect 939 -1224 942 -1218
rect 946 -1224 952 -1218
rect 953 -1224 956 -1218
rect 960 -1224 963 -1218
rect 967 -1224 970 -1218
rect 974 -1224 977 -1218
rect 981 -1224 984 -1218
rect 988 -1224 991 -1218
rect 995 -1224 998 -1218
rect 1002 -1224 1005 -1218
rect 1009 -1224 1012 -1218
rect 1016 -1224 1019 -1218
rect 1023 -1224 1026 -1218
rect 1030 -1224 1033 -1218
rect 1037 -1224 1040 -1218
rect 1044 -1224 1047 -1218
rect 1051 -1224 1057 -1218
rect 1058 -1224 1061 -1218
rect 1065 -1224 1068 -1218
rect 1072 -1224 1075 -1218
rect 1079 -1224 1082 -1218
rect 1086 -1224 1089 -1218
rect 1093 -1224 1096 -1218
rect 1100 -1224 1103 -1218
rect 1107 -1224 1110 -1218
rect 1114 -1224 1117 -1218
rect 1121 -1224 1124 -1218
rect 1128 -1224 1131 -1218
rect 1135 -1224 1138 -1218
rect 1142 -1224 1145 -1218
rect 1149 -1224 1152 -1218
rect 1156 -1224 1159 -1218
rect 1163 -1224 1166 -1218
rect 1170 -1224 1173 -1218
rect 1177 -1224 1180 -1218
rect 1184 -1224 1187 -1218
rect 1191 -1224 1194 -1218
rect 1198 -1224 1201 -1218
rect 1205 -1224 1208 -1218
rect 1212 -1224 1215 -1218
rect 1219 -1224 1222 -1218
rect 1226 -1224 1229 -1218
rect 1233 -1224 1236 -1218
rect 1240 -1224 1243 -1218
rect 1247 -1224 1250 -1218
rect 1254 -1224 1257 -1218
rect 1261 -1224 1264 -1218
rect 1268 -1224 1271 -1218
rect 1275 -1224 1278 -1218
rect 1282 -1224 1285 -1218
rect 1289 -1224 1292 -1218
rect 1296 -1224 1299 -1218
rect 1303 -1224 1306 -1218
rect 1310 -1224 1313 -1218
rect 1317 -1224 1320 -1218
rect 1324 -1224 1327 -1218
rect 1331 -1224 1334 -1218
rect 1338 -1224 1341 -1218
rect 1345 -1224 1348 -1218
rect 1352 -1224 1355 -1218
rect 1359 -1224 1362 -1218
rect 1366 -1224 1369 -1218
rect 1373 -1224 1376 -1218
rect 1380 -1224 1383 -1218
rect 1387 -1224 1390 -1218
rect 1394 -1224 1397 -1218
rect 1401 -1224 1404 -1218
rect 1408 -1224 1411 -1218
rect 1415 -1224 1418 -1218
rect 1422 -1224 1425 -1218
rect 1429 -1224 1432 -1218
rect 1436 -1224 1439 -1218
rect 1443 -1224 1446 -1218
rect 1450 -1224 1453 -1218
rect 1457 -1224 1460 -1218
rect 1464 -1224 1467 -1218
rect 1471 -1224 1474 -1218
rect 1478 -1224 1481 -1218
rect 1485 -1224 1488 -1218
rect 1492 -1224 1495 -1218
rect 1499 -1224 1502 -1218
rect 1506 -1224 1509 -1218
rect 1513 -1224 1516 -1218
rect 1520 -1224 1523 -1218
rect 1527 -1224 1530 -1218
rect 1534 -1224 1537 -1218
rect 1541 -1224 1544 -1218
rect 1548 -1224 1551 -1218
rect 1555 -1224 1558 -1218
rect 1562 -1224 1565 -1218
rect 1569 -1224 1572 -1218
rect 1576 -1224 1579 -1218
rect 1583 -1224 1586 -1218
rect 1590 -1224 1593 -1218
rect 1597 -1224 1600 -1218
rect 1604 -1224 1607 -1218
rect 1611 -1224 1614 -1218
rect 1618 -1224 1621 -1218
rect 1625 -1224 1628 -1218
rect 1632 -1224 1635 -1218
rect 1639 -1224 1642 -1218
rect 1646 -1224 1649 -1218
rect 1653 -1224 1656 -1218
rect 1660 -1224 1663 -1218
rect 1667 -1224 1670 -1218
rect 1674 -1224 1677 -1218
rect 1681 -1224 1684 -1218
rect 1688 -1224 1691 -1218
rect 1695 -1224 1698 -1218
rect 1702 -1224 1705 -1218
rect 1709 -1224 1712 -1218
rect 1716 -1224 1719 -1218
rect 1723 -1224 1726 -1218
rect 1730 -1224 1733 -1218
rect 1737 -1224 1740 -1218
rect 1744 -1224 1750 -1218
rect 1751 -1224 1754 -1218
rect 1758 -1224 1761 -1218
rect 1765 -1224 1771 -1218
rect 1772 -1224 1778 -1218
rect 1779 -1224 1782 -1218
rect 1786 -1224 1789 -1218
rect 1 -1367 7 -1361
rect 8 -1367 14 -1361
rect 15 -1367 18 -1361
rect 22 -1367 25 -1361
rect 29 -1367 32 -1361
rect 36 -1367 42 -1361
rect 43 -1367 46 -1361
rect 50 -1367 56 -1361
rect 57 -1367 63 -1361
rect 64 -1367 67 -1361
rect 71 -1367 74 -1361
rect 78 -1367 84 -1361
rect 85 -1367 88 -1361
rect 92 -1367 95 -1361
rect 99 -1367 105 -1361
rect 106 -1367 112 -1361
rect 113 -1367 116 -1361
rect 120 -1367 123 -1361
rect 127 -1367 133 -1361
rect 134 -1367 137 -1361
rect 141 -1367 144 -1361
rect 148 -1367 151 -1361
rect 155 -1367 158 -1361
rect 162 -1367 165 -1361
rect 169 -1367 172 -1361
rect 176 -1367 179 -1361
rect 183 -1367 189 -1361
rect 190 -1367 193 -1361
rect 197 -1367 203 -1361
rect 204 -1367 210 -1361
rect 211 -1367 214 -1361
rect 218 -1367 224 -1361
rect 225 -1367 228 -1361
rect 232 -1367 235 -1361
rect 239 -1367 242 -1361
rect 246 -1367 249 -1361
rect 253 -1367 256 -1361
rect 260 -1367 263 -1361
rect 267 -1367 270 -1361
rect 274 -1367 277 -1361
rect 281 -1367 284 -1361
rect 288 -1367 294 -1361
rect 295 -1367 298 -1361
rect 302 -1367 305 -1361
rect 309 -1367 312 -1361
rect 316 -1367 319 -1361
rect 323 -1367 326 -1361
rect 330 -1367 333 -1361
rect 337 -1367 340 -1361
rect 344 -1367 347 -1361
rect 351 -1367 354 -1361
rect 358 -1367 361 -1361
rect 365 -1367 368 -1361
rect 372 -1367 375 -1361
rect 379 -1367 382 -1361
rect 386 -1367 389 -1361
rect 393 -1367 396 -1361
rect 400 -1367 403 -1361
rect 407 -1367 410 -1361
rect 414 -1367 417 -1361
rect 421 -1367 424 -1361
rect 428 -1367 431 -1361
rect 435 -1367 438 -1361
rect 442 -1367 448 -1361
rect 449 -1367 455 -1361
rect 456 -1367 459 -1361
rect 463 -1367 466 -1361
rect 470 -1367 473 -1361
rect 477 -1367 480 -1361
rect 484 -1367 487 -1361
rect 491 -1367 494 -1361
rect 498 -1367 501 -1361
rect 505 -1367 508 -1361
rect 512 -1367 515 -1361
rect 519 -1367 522 -1361
rect 526 -1367 529 -1361
rect 533 -1367 536 -1361
rect 540 -1367 543 -1361
rect 547 -1367 553 -1361
rect 554 -1367 560 -1361
rect 561 -1367 567 -1361
rect 568 -1367 574 -1361
rect 575 -1367 578 -1361
rect 582 -1367 585 -1361
rect 589 -1367 592 -1361
rect 596 -1367 602 -1361
rect 603 -1367 606 -1361
rect 610 -1367 613 -1361
rect 617 -1367 620 -1361
rect 624 -1367 627 -1361
rect 631 -1367 634 -1361
rect 638 -1367 641 -1361
rect 645 -1367 648 -1361
rect 652 -1367 655 -1361
rect 659 -1367 662 -1361
rect 666 -1367 669 -1361
rect 673 -1367 676 -1361
rect 680 -1367 683 -1361
rect 687 -1367 690 -1361
rect 694 -1367 697 -1361
rect 701 -1367 704 -1361
rect 708 -1367 711 -1361
rect 715 -1367 718 -1361
rect 722 -1367 725 -1361
rect 729 -1367 732 -1361
rect 736 -1367 742 -1361
rect 743 -1367 746 -1361
rect 750 -1367 756 -1361
rect 757 -1367 760 -1361
rect 764 -1367 767 -1361
rect 771 -1367 774 -1361
rect 778 -1367 781 -1361
rect 785 -1367 791 -1361
rect 792 -1367 795 -1361
rect 799 -1367 802 -1361
rect 806 -1367 809 -1361
rect 813 -1367 819 -1361
rect 820 -1367 826 -1361
rect 827 -1367 833 -1361
rect 834 -1367 837 -1361
rect 841 -1367 844 -1361
rect 848 -1367 854 -1361
rect 855 -1367 858 -1361
rect 862 -1367 865 -1361
rect 869 -1367 872 -1361
rect 876 -1367 879 -1361
rect 883 -1367 886 -1361
rect 890 -1367 893 -1361
rect 897 -1367 900 -1361
rect 904 -1367 907 -1361
rect 911 -1367 914 -1361
rect 918 -1367 924 -1361
rect 925 -1367 928 -1361
rect 932 -1367 938 -1361
rect 939 -1367 942 -1361
rect 946 -1367 952 -1361
rect 953 -1367 956 -1361
rect 960 -1367 963 -1361
rect 967 -1367 970 -1361
rect 974 -1367 977 -1361
rect 981 -1367 987 -1361
rect 988 -1367 991 -1361
rect 995 -1367 998 -1361
rect 1002 -1367 1008 -1361
rect 1009 -1367 1012 -1361
rect 1016 -1367 1022 -1361
rect 1023 -1367 1026 -1361
rect 1030 -1367 1033 -1361
rect 1037 -1367 1040 -1361
rect 1044 -1367 1047 -1361
rect 1051 -1367 1054 -1361
rect 1058 -1367 1061 -1361
rect 1065 -1367 1068 -1361
rect 1072 -1367 1075 -1361
rect 1079 -1367 1082 -1361
rect 1086 -1367 1089 -1361
rect 1093 -1367 1096 -1361
rect 1100 -1367 1106 -1361
rect 1107 -1367 1110 -1361
rect 1114 -1367 1117 -1361
rect 1121 -1367 1124 -1361
rect 1128 -1367 1131 -1361
rect 1135 -1367 1138 -1361
rect 1142 -1367 1148 -1361
rect 1149 -1367 1152 -1361
rect 1156 -1367 1159 -1361
rect 1163 -1367 1166 -1361
rect 1170 -1367 1173 -1361
rect 1177 -1367 1180 -1361
rect 1184 -1367 1187 -1361
rect 1191 -1367 1194 -1361
rect 1198 -1367 1204 -1361
rect 1205 -1367 1208 -1361
rect 1212 -1367 1218 -1361
rect 1219 -1367 1222 -1361
rect 1226 -1367 1229 -1361
rect 1233 -1367 1236 -1361
rect 1240 -1367 1243 -1361
rect 1247 -1367 1250 -1361
rect 1254 -1367 1257 -1361
rect 1261 -1367 1264 -1361
rect 1268 -1367 1271 -1361
rect 1275 -1367 1278 -1361
rect 1282 -1367 1285 -1361
rect 1289 -1367 1292 -1361
rect 1296 -1367 1299 -1361
rect 1303 -1367 1306 -1361
rect 1310 -1367 1313 -1361
rect 1317 -1367 1320 -1361
rect 1324 -1367 1327 -1361
rect 1331 -1367 1334 -1361
rect 1338 -1367 1341 -1361
rect 1345 -1367 1348 -1361
rect 1352 -1367 1355 -1361
rect 1359 -1367 1362 -1361
rect 1366 -1367 1369 -1361
rect 1373 -1367 1376 -1361
rect 1380 -1367 1383 -1361
rect 1387 -1367 1390 -1361
rect 1394 -1367 1397 -1361
rect 1401 -1367 1404 -1361
rect 1408 -1367 1411 -1361
rect 1415 -1367 1418 -1361
rect 1422 -1367 1425 -1361
rect 1429 -1367 1432 -1361
rect 1436 -1367 1439 -1361
rect 1443 -1367 1446 -1361
rect 1450 -1367 1453 -1361
rect 1457 -1367 1460 -1361
rect 1464 -1367 1467 -1361
rect 1471 -1367 1474 -1361
rect 1478 -1367 1481 -1361
rect 1485 -1367 1488 -1361
rect 1492 -1367 1495 -1361
rect 1499 -1367 1502 -1361
rect 1506 -1367 1509 -1361
rect 1513 -1367 1516 -1361
rect 1520 -1367 1523 -1361
rect 1527 -1367 1530 -1361
rect 1534 -1367 1537 -1361
rect 1541 -1367 1544 -1361
rect 1548 -1367 1551 -1361
rect 1555 -1367 1558 -1361
rect 1562 -1367 1565 -1361
rect 1569 -1367 1572 -1361
rect 1576 -1367 1579 -1361
rect 1583 -1367 1586 -1361
rect 1590 -1367 1593 -1361
rect 1597 -1367 1600 -1361
rect 1604 -1367 1607 -1361
rect 1611 -1367 1614 -1361
rect 1618 -1367 1621 -1361
rect 1625 -1367 1628 -1361
rect 1632 -1367 1635 -1361
rect 1639 -1367 1642 -1361
rect 1646 -1367 1649 -1361
rect 1653 -1367 1656 -1361
rect 1660 -1367 1663 -1361
rect 1667 -1367 1670 -1361
rect 1674 -1367 1677 -1361
rect 1681 -1367 1684 -1361
rect 1688 -1367 1691 -1361
rect 1695 -1367 1698 -1361
rect 1702 -1367 1705 -1361
rect 1709 -1367 1712 -1361
rect 1716 -1367 1719 -1361
rect 1723 -1367 1726 -1361
rect 1730 -1367 1733 -1361
rect 1737 -1367 1740 -1361
rect 1744 -1367 1747 -1361
rect 1751 -1367 1754 -1361
rect 1 -1508 7 -1502
rect 8 -1508 14 -1502
rect 15 -1508 21 -1502
rect 22 -1508 25 -1502
rect 29 -1508 32 -1502
rect 36 -1508 39 -1502
rect 43 -1508 46 -1502
rect 50 -1508 53 -1502
rect 57 -1508 60 -1502
rect 64 -1508 70 -1502
rect 71 -1508 74 -1502
rect 78 -1508 81 -1502
rect 85 -1508 88 -1502
rect 92 -1508 95 -1502
rect 99 -1508 102 -1502
rect 106 -1508 109 -1502
rect 113 -1508 116 -1502
rect 120 -1508 126 -1502
rect 127 -1508 133 -1502
rect 134 -1508 137 -1502
rect 141 -1508 144 -1502
rect 148 -1508 151 -1502
rect 155 -1508 161 -1502
rect 162 -1508 165 -1502
rect 169 -1508 172 -1502
rect 176 -1508 179 -1502
rect 183 -1508 189 -1502
rect 190 -1508 196 -1502
rect 197 -1508 200 -1502
rect 204 -1508 207 -1502
rect 211 -1508 217 -1502
rect 218 -1508 221 -1502
rect 225 -1508 231 -1502
rect 232 -1508 235 -1502
rect 239 -1508 242 -1502
rect 246 -1508 249 -1502
rect 253 -1508 259 -1502
rect 260 -1508 263 -1502
rect 267 -1508 270 -1502
rect 274 -1508 277 -1502
rect 281 -1508 284 -1502
rect 288 -1508 291 -1502
rect 295 -1508 298 -1502
rect 302 -1508 305 -1502
rect 309 -1508 312 -1502
rect 316 -1508 322 -1502
rect 323 -1508 326 -1502
rect 330 -1508 333 -1502
rect 337 -1508 340 -1502
rect 344 -1508 347 -1502
rect 351 -1508 354 -1502
rect 358 -1508 361 -1502
rect 365 -1508 368 -1502
rect 372 -1508 375 -1502
rect 379 -1508 382 -1502
rect 386 -1508 389 -1502
rect 393 -1508 396 -1502
rect 400 -1508 403 -1502
rect 407 -1508 410 -1502
rect 414 -1508 420 -1502
rect 421 -1508 424 -1502
rect 428 -1508 431 -1502
rect 435 -1508 438 -1502
rect 442 -1508 445 -1502
rect 449 -1508 452 -1502
rect 456 -1508 462 -1502
rect 463 -1508 466 -1502
rect 470 -1508 473 -1502
rect 477 -1508 483 -1502
rect 484 -1508 487 -1502
rect 491 -1508 494 -1502
rect 498 -1508 501 -1502
rect 505 -1508 508 -1502
rect 512 -1508 518 -1502
rect 519 -1508 522 -1502
rect 526 -1508 529 -1502
rect 533 -1508 536 -1502
rect 540 -1508 543 -1502
rect 547 -1508 550 -1502
rect 554 -1508 557 -1502
rect 561 -1508 564 -1502
rect 568 -1508 571 -1502
rect 575 -1508 578 -1502
rect 582 -1508 585 -1502
rect 589 -1508 592 -1502
rect 596 -1508 599 -1502
rect 603 -1508 606 -1502
rect 610 -1508 613 -1502
rect 617 -1508 620 -1502
rect 624 -1508 630 -1502
rect 631 -1508 634 -1502
rect 638 -1508 641 -1502
rect 645 -1508 648 -1502
rect 652 -1508 658 -1502
rect 659 -1508 662 -1502
rect 666 -1508 672 -1502
rect 673 -1508 676 -1502
rect 680 -1508 683 -1502
rect 687 -1508 690 -1502
rect 694 -1508 697 -1502
rect 701 -1508 704 -1502
rect 708 -1508 711 -1502
rect 715 -1508 721 -1502
rect 722 -1508 728 -1502
rect 729 -1508 732 -1502
rect 736 -1508 742 -1502
rect 743 -1508 746 -1502
rect 750 -1508 753 -1502
rect 757 -1508 763 -1502
rect 764 -1508 767 -1502
rect 771 -1508 774 -1502
rect 778 -1508 781 -1502
rect 785 -1508 791 -1502
rect 792 -1508 795 -1502
rect 799 -1508 802 -1502
rect 806 -1508 809 -1502
rect 813 -1508 816 -1502
rect 820 -1508 826 -1502
rect 827 -1508 833 -1502
rect 834 -1508 837 -1502
rect 841 -1508 844 -1502
rect 848 -1508 851 -1502
rect 855 -1508 858 -1502
rect 862 -1508 868 -1502
rect 869 -1508 872 -1502
rect 876 -1508 879 -1502
rect 883 -1508 886 -1502
rect 890 -1508 893 -1502
rect 897 -1508 900 -1502
rect 904 -1508 907 -1502
rect 911 -1508 914 -1502
rect 918 -1508 921 -1502
rect 925 -1508 928 -1502
rect 932 -1508 938 -1502
rect 939 -1508 942 -1502
rect 946 -1508 952 -1502
rect 953 -1508 956 -1502
rect 960 -1508 963 -1502
rect 967 -1508 970 -1502
rect 974 -1508 980 -1502
rect 981 -1508 984 -1502
rect 988 -1508 991 -1502
rect 995 -1508 998 -1502
rect 1002 -1508 1005 -1502
rect 1009 -1508 1012 -1502
rect 1016 -1508 1019 -1502
rect 1023 -1508 1026 -1502
rect 1030 -1508 1036 -1502
rect 1037 -1508 1040 -1502
rect 1044 -1508 1050 -1502
rect 1051 -1508 1054 -1502
rect 1058 -1508 1061 -1502
rect 1065 -1508 1068 -1502
rect 1072 -1508 1075 -1502
rect 1079 -1508 1082 -1502
rect 1086 -1508 1089 -1502
rect 1093 -1508 1096 -1502
rect 1100 -1508 1103 -1502
rect 1107 -1508 1110 -1502
rect 1114 -1508 1117 -1502
rect 1121 -1508 1124 -1502
rect 1128 -1508 1131 -1502
rect 1135 -1508 1138 -1502
rect 1142 -1508 1145 -1502
rect 1149 -1508 1152 -1502
rect 1156 -1508 1159 -1502
rect 1163 -1508 1166 -1502
rect 1170 -1508 1173 -1502
rect 1177 -1508 1180 -1502
rect 1184 -1508 1187 -1502
rect 1191 -1508 1194 -1502
rect 1198 -1508 1201 -1502
rect 1205 -1508 1208 -1502
rect 1212 -1508 1215 -1502
rect 1219 -1508 1222 -1502
rect 1226 -1508 1229 -1502
rect 1233 -1508 1236 -1502
rect 1240 -1508 1243 -1502
rect 1247 -1508 1250 -1502
rect 1254 -1508 1257 -1502
rect 1261 -1508 1264 -1502
rect 1268 -1508 1271 -1502
rect 1275 -1508 1278 -1502
rect 1282 -1508 1285 -1502
rect 1289 -1508 1292 -1502
rect 1296 -1508 1299 -1502
rect 1303 -1508 1306 -1502
rect 1310 -1508 1313 -1502
rect 1317 -1508 1320 -1502
rect 1324 -1508 1327 -1502
rect 1331 -1508 1334 -1502
rect 1338 -1508 1341 -1502
rect 1345 -1508 1348 -1502
rect 1352 -1508 1355 -1502
rect 1359 -1508 1362 -1502
rect 1366 -1508 1369 -1502
rect 1373 -1508 1376 -1502
rect 1380 -1508 1383 -1502
rect 1387 -1508 1390 -1502
rect 1394 -1508 1397 -1502
rect 1401 -1508 1404 -1502
rect 1408 -1508 1411 -1502
rect 1415 -1508 1418 -1502
rect 1422 -1508 1425 -1502
rect 1429 -1508 1432 -1502
rect 1436 -1508 1439 -1502
rect 1443 -1508 1446 -1502
rect 1450 -1508 1453 -1502
rect 1457 -1508 1460 -1502
rect 1464 -1508 1467 -1502
rect 1471 -1508 1474 -1502
rect 1478 -1508 1481 -1502
rect 1485 -1508 1488 -1502
rect 1492 -1508 1495 -1502
rect 1499 -1508 1502 -1502
rect 1506 -1508 1509 -1502
rect 1513 -1508 1516 -1502
rect 1520 -1508 1523 -1502
rect 1527 -1508 1530 -1502
rect 1534 -1508 1540 -1502
rect 1541 -1508 1544 -1502
rect 1548 -1508 1554 -1502
rect 1555 -1508 1558 -1502
rect 1562 -1508 1565 -1502
rect 1569 -1508 1572 -1502
rect 1576 -1508 1579 -1502
rect 1583 -1508 1589 -1502
rect 1590 -1508 1593 -1502
rect 1597 -1508 1600 -1502
rect 1604 -1508 1610 -1502
rect 1611 -1508 1614 -1502
rect 1618 -1508 1621 -1502
rect 1625 -1508 1628 -1502
rect 1632 -1508 1635 -1502
rect 1639 -1508 1645 -1502
rect 1646 -1508 1649 -1502
rect 1653 -1508 1656 -1502
rect 1660 -1508 1663 -1502
rect 1667 -1508 1670 -1502
rect 1674 -1508 1677 -1502
rect 1681 -1508 1684 -1502
rect 1688 -1508 1691 -1502
rect 1695 -1508 1698 -1502
rect 1702 -1508 1705 -1502
rect 1709 -1508 1712 -1502
rect 1716 -1508 1719 -1502
rect 1723 -1508 1726 -1502
rect 1730 -1508 1733 -1502
rect 1800 -1508 1803 -1502
rect 1 -1643 7 -1637
rect 8 -1643 14 -1637
rect 15 -1643 21 -1637
rect 22 -1643 25 -1637
rect 29 -1643 32 -1637
rect 36 -1643 39 -1637
rect 43 -1643 46 -1637
rect 50 -1643 53 -1637
rect 57 -1643 63 -1637
rect 64 -1643 67 -1637
rect 71 -1643 74 -1637
rect 78 -1643 81 -1637
rect 85 -1643 88 -1637
rect 92 -1643 95 -1637
rect 99 -1643 102 -1637
rect 106 -1643 109 -1637
rect 113 -1643 116 -1637
rect 120 -1643 126 -1637
rect 127 -1643 130 -1637
rect 134 -1643 137 -1637
rect 141 -1643 144 -1637
rect 148 -1643 151 -1637
rect 155 -1643 158 -1637
rect 162 -1643 168 -1637
rect 169 -1643 172 -1637
rect 176 -1643 179 -1637
rect 183 -1643 189 -1637
rect 190 -1643 193 -1637
rect 197 -1643 200 -1637
rect 204 -1643 207 -1637
rect 211 -1643 214 -1637
rect 218 -1643 224 -1637
rect 225 -1643 228 -1637
rect 232 -1643 235 -1637
rect 239 -1643 242 -1637
rect 246 -1643 249 -1637
rect 253 -1643 256 -1637
rect 260 -1643 266 -1637
rect 267 -1643 270 -1637
rect 274 -1643 277 -1637
rect 281 -1643 284 -1637
rect 288 -1643 291 -1637
rect 295 -1643 298 -1637
rect 302 -1643 305 -1637
rect 309 -1643 315 -1637
rect 316 -1643 319 -1637
rect 323 -1643 326 -1637
rect 330 -1643 333 -1637
rect 337 -1643 340 -1637
rect 344 -1643 347 -1637
rect 351 -1643 354 -1637
rect 358 -1643 361 -1637
rect 365 -1643 368 -1637
rect 372 -1643 375 -1637
rect 379 -1643 382 -1637
rect 386 -1643 389 -1637
rect 393 -1643 396 -1637
rect 400 -1643 403 -1637
rect 407 -1643 410 -1637
rect 414 -1643 417 -1637
rect 421 -1643 424 -1637
rect 428 -1643 431 -1637
rect 435 -1643 438 -1637
rect 442 -1643 448 -1637
rect 449 -1643 455 -1637
rect 456 -1643 459 -1637
rect 463 -1643 466 -1637
rect 470 -1643 473 -1637
rect 477 -1643 480 -1637
rect 484 -1643 487 -1637
rect 491 -1643 494 -1637
rect 498 -1643 501 -1637
rect 505 -1643 508 -1637
rect 512 -1643 515 -1637
rect 519 -1643 522 -1637
rect 526 -1643 529 -1637
rect 533 -1643 536 -1637
rect 540 -1643 546 -1637
rect 547 -1643 553 -1637
rect 554 -1643 557 -1637
rect 561 -1643 564 -1637
rect 568 -1643 571 -1637
rect 575 -1643 578 -1637
rect 582 -1643 585 -1637
rect 589 -1643 592 -1637
rect 596 -1643 599 -1637
rect 603 -1643 609 -1637
rect 610 -1643 613 -1637
rect 617 -1643 620 -1637
rect 624 -1643 627 -1637
rect 631 -1643 634 -1637
rect 638 -1643 641 -1637
rect 645 -1643 648 -1637
rect 652 -1643 655 -1637
rect 659 -1643 662 -1637
rect 666 -1643 669 -1637
rect 673 -1643 676 -1637
rect 680 -1643 683 -1637
rect 687 -1643 690 -1637
rect 694 -1643 697 -1637
rect 701 -1643 704 -1637
rect 708 -1643 711 -1637
rect 715 -1643 718 -1637
rect 722 -1643 728 -1637
rect 729 -1643 735 -1637
rect 736 -1643 739 -1637
rect 743 -1643 749 -1637
rect 750 -1643 756 -1637
rect 757 -1643 760 -1637
rect 764 -1643 767 -1637
rect 771 -1643 774 -1637
rect 778 -1643 781 -1637
rect 785 -1643 788 -1637
rect 792 -1643 795 -1637
rect 799 -1643 802 -1637
rect 806 -1643 809 -1637
rect 813 -1643 819 -1637
rect 820 -1643 826 -1637
rect 827 -1643 830 -1637
rect 834 -1643 837 -1637
rect 841 -1643 844 -1637
rect 848 -1643 851 -1637
rect 855 -1643 861 -1637
rect 862 -1643 868 -1637
rect 869 -1643 872 -1637
rect 876 -1643 882 -1637
rect 883 -1643 886 -1637
rect 890 -1643 896 -1637
rect 897 -1643 900 -1637
rect 904 -1643 907 -1637
rect 911 -1643 914 -1637
rect 918 -1643 921 -1637
rect 925 -1643 928 -1637
rect 932 -1643 935 -1637
rect 939 -1643 942 -1637
rect 946 -1643 949 -1637
rect 953 -1643 959 -1637
rect 960 -1643 963 -1637
rect 967 -1643 970 -1637
rect 974 -1643 977 -1637
rect 981 -1643 984 -1637
rect 988 -1643 991 -1637
rect 995 -1643 998 -1637
rect 1002 -1643 1008 -1637
rect 1009 -1643 1012 -1637
rect 1016 -1643 1022 -1637
rect 1023 -1643 1026 -1637
rect 1030 -1643 1033 -1637
rect 1037 -1643 1040 -1637
rect 1044 -1643 1047 -1637
rect 1051 -1643 1054 -1637
rect 1058 -1643 1064 -1637
rect 1065 -1643 1068 -1637
rect 1072 -1643 1075 -1637
rect 1079 -1643 1085 -1637
rect 1086 -1643 1089 -1637
rect 1093 -1643 1096 -1637
rect 1100 -1643 1103 -1637
rect 1107 -1643 1113 -1637
rect 1114 -1643 1117 -1637
rect 1121 -1643 1127 -1637
rect 1128 -1643 1131 -1637
rect 1135 -1643 1138 -1637
rect 1142 -1643 1145 -1637
rect 1149 -1643 1152 -1637
rect 1156 -1643 1159 -1637
rect 1163 -1643 1166 -1637
rect 1170 -1643 1173 -1637
rect 1177 -1643 1180 -1637
rect 1184 -1643 1190 -1637
rect 1191 -1643 1194 -1637
rect 1198 -1643 1201 -1637
rect 1205 -1643 1211 -1637
rect 1212 -1643 1215 -1637
rect 1219 -1643 1222 -1637
rect 1226 -1643 1229 -1637
rect 1233 -1643 1236 -1637
rect 1240 -1643 1243 -1637
rect 1247 -1643 1250 -1637
rect 1254 -1643 1257 -1637
rect 1261 -1643 1264 -1637
rect 1268 -1643 1271 -1637
rect 1275 -1643 1278 -1637
rect 1282 -1643 1285 -1637
rect 1289 -1643 1292 -1637
rect 1296 -1643 1302 -1637
rect 1303 -1643 1306 -1637
rect 1310 -1643 1313 -1637
rect 1317 -1643 1320 -1637
rect 1324 -1643 1327 -1637
rect 1331 -1643 1334 -1637
rect 1338 -1643 1341 -1637
rect 1345 -1643 1348 -1637
rect 1352 -1643 1355 -1637
rect 1359 -1643 1362 -1637
rect 1366 -1643 1369 -1637
rect 1373 -1643 1376 -1637
rect 1380 -1643 1383 -1637
rect 1387 -1643 1390 -1637
rect 1394 -1643 1397 -1637
rect 1401 -1643 1404 -1637
rect 1408 -1643 1411 -1637
rect 1415 -1643 1418 -1637
rect 1422 -1643 1425 -1637
rect 1429 -1643 1432 -1637
rect 1436 -1643 1439 -1637
rect 1443 -1643 1446 -1637
rect 1450 -1643 1453 -1637
rect 1457 -1643 1460 -1637
rect 1464 -1643 1467 -1637
rect 1471 -1643 1474 -1637
rect 1478 -1643 1481 -1637
rect 1485 -1643 1488 -1637
rect 1492 -1643 1495 -1637
rect 1499 -1643 1502 -1637
rect 1506 -1643 1509 -1637
rect 1513 -1643 1516 -1637
rect 1520 -1643 1523 -1637
rect 1527 -1643 1530 -1637
rect 1534 -1643 1537 -1637
rect 1541 -1643 1544 -1637
rect 1548 -1643 1551 -1637
rect 1555 -1643 1558 -1637
rect 1562 -1643 1565 -1637
rect 1569 -1643 1572 -1637
rect 1576 -1643 1579 -1637
rect 1583 -1643 1586 -1637
rect 1590 -1643 1593 -1637
rect 1597 -1643 1600 -1637
rect 1604 -1643 1607 -1637
rect 1611 -1643 1614 -1637
rect 1618 -1643 1621 -1637
rect 1625 -1643 1628 -1637
rect 1632 -1643 1635 -1637
rect 1639 -1643 1642 -1637
rect 1646 -1643 1652 -1637
rect 1653 -1643 1656 -1637
rect 1660 -1643 1663 -1637
rect 1667 -1643 1670 -1637
rect 1674 -1643 1677 -1637
rect 1681 -1643 1687 -1637
rect 1688 -1643 1691 -1637
rect 1695 -1643 1698 -1637
rect 1702 -1643 1708 -1637
rect 1709 -1643 1712 -1637
rect 1716 -1643 1719 -1637
rect 1723 -1643 1726 -1637
rect 1821 -1643 1824 -1637
rect 1 -1790 7 -1784
rect 8 -1790 14 -1784
rect 15 -1790 21 -1784
rect 22 -1790 25 -1784
rect 29 -1790 32 -1784
rect 36 -1790 39 -1784
rect 43 -1790 46 -1784
rect 50 -1790 53 -1784
rect 57 -1790 60 -1784
rect 64 -1790 67 -1784
rect 71 -1790 77 -1784
rect 78 -1790 81 -1784
rect 85 -1790 91 -1784
rect 92 -1790 95 -1784
rect 99 -1790 102 -1784
rect 106 -1790 109 -1784
rect 113 -1790 119 -1784
rect 120 -1790 123 -1784
rect 127 -1790 130 -1784
rect 134 -1790 137 -1784
rect 141 -1790 147 -1784
rect 148 -1790 151 -1784
rect 155 -1790 161 -1784
rect 162 -1790 165 -1784
rect 169 -1790 172 -1784
rect 176 -1790 179 -1784
rect 183 -1790 186 -1784
rect 190 -1790 193 -1784
rect 197 -1790 200 -1784
rect 204 -1790 207 -1784
rect 211 -1790 214 -1784
rect 218 -1790 224 -1784
rect 225 -1790 228 -1784
rect 232 -1790 238 -1784
rect 239 -1790 242 -1784
rect 246 -1790 249 -1784
rect 253 -1790 256 -1784
rect 260 -1790 266 -1784
rect 267 -1790 270 -1784
rect 274 -1790 277 -1784
rect 281 -1790 284 -1784
rect 288 -1790 291 -1784
rect 295 -1790 298 -1784
rect 302 -1790 305 -1784
rect 309 -1790 312 -1784
rect 316 -1790 319 -1784
rect 323 -1790 326 -1784
rect 330 -1790 333 -1784
rect 337 -1790 340 -1784
rect 344 -1790 347 -1784
rect 351 -1790 354 -1784
rect 358 -1790 364 -1784
rect 365 -1790 368 -1784
rect 372 -1790 375 -1784
rect 379 -1790 385 -1784
rect 386 -1790 389 -1784
rect 393 -1790 396 -1784
rect 400 -1790 403 -1784
rect 407 -1790 410 -1784
rect 414 -1790 417 -1784
rect 421 -1790 424 -1784
rect 428 -1790 431 -1784
rect 435 -1790 438 -1784
rect 442 -1790 445 -1784
rect 449 -1790 452 -1784
rect 456 -1790 459 -1784
rect 463 -1790 466 -1784
rect 470 -1790 473 -1784
rect 477 -1790 480 -1784
rect 484 -1790 487 -1784
rect 491 -1790 494 -1784
rect 498 -1790 504 -1784
rect 505 -1790 508 -1784
rect 512 -1790 515 -1784
rect 519 -1790 522 -1784
rect 526 -1790 529 -1784
rect 533 -1790 539 -1784
rect 540 -1790 546 -1784
rect 547 -1790 553 -1784
rect 554 -1790 557 -1784
rect 561 -1790 564 -1784
rect 568 -1790 571 -1784
rect 575 -1790 581 -1784
rect 582 -1790 588 -1784
rect 589 -1790 595 -1784
rect 596 -1790 599 -1784
rect 603 -1790 606 -1784
rect 610 -1790 613 -1784
rect 617 -1790 620 -1784
rect 624 -1790 627 -1784
rect 631 -1790 637 -1784
rect 638 -1790 641 -1784
rect 645 -1790 648 -1784
rect 652 -1790 655 -1784
rect 659 -1790 662 -1784
rect 666 -1790 669 -1784
rect 673 -1790 679 -1784
rect 680 -1790 683 -1784
rect 687 -1790 690 -1784
rect 694 -1790 697 -1784
rect 701 -1790 707 -1784
rect 708 -1790 711 -1784
rect 715 -1790 721 -1784
rect 722 -1790 728 -1784
rect 729 -1790 735 -1784
rect 736 -1790 739 -1784
rect 743 -1790 746 -1784
rect 750 -1790 753 -1784
rect 757 -1790 760 -1784
rect 764 -1790 767 -1784
rect 771 -1790 774 -1784
rect 778 -1790 784 -1784
rect 785 -1790 791 -1784
rect 792 -1790 795 -1784
rect 799 -1790 802 -1784
rect 806 -1790 809 -1784
rect 813 -1790 816 -1784
rect 820 -1790 826 -1784
rect 827 -1790 830 -1784
rect 834 -1790 837 -1784
rect 841 -1790 844 -1784
rect 848 -1790 851 -1784
rect 855 -1790 858 -1784
rect 862 -1790 865 -1784
rect 869 -1790 872 -1784
rect 876 -1790 879 -1784
rect 883 -1790 889 -1784
rect 890 -1790 893 -1784
rect 897 -1790 903 -1784
rect 904 -1790 907 -1784
rect 911 -1790 914 -1784
rect 918 -1790 921 -1784
rect 925 -1790 928 -1784
rect 932 -1790 935 -1784
rect 939 -1790 942 -1784
rect 946 -1790 952 -1784
rect 953 -1790 956 -1784
rect 960 -1790 963 -1784
rect 967 -1790 970 -1784
rect 974 -1790 980 -1784
rect 981 -1790 984 -1784
rect 988 -1790 991 -1784
rect 995 -1790 998 -1784
rect 1002 -1790 1005 -1784
rect 1009 -1790 1012 -1784
rect 1016 -1790 1019 -1784
rect 1023 -1790 1029 -1784
rect 1030 -1790 1033 -1784
rect 1037 -1790 1040 -1784
rect 1044 -1790 1047 -1784
rect 1051 -1790 1057 -1784
rect 1058 -1790 1061 -1784
rect 1065 -1790 1068 -1784
rect 1072 -1790 1075 -1784
rect 1079 -1790 1082 -1784
rect 1086 -1790 1089 -1784
rect 1093 -1790 1096 -1784
rect 1100 -1790 1103 -1784
rect 1107 -1790 1110 -1784
rect 1114 -1790 1117 -1784
rect 1121 -1790 1124 -1784
rect 1128 -1790 1131 -1784
rect 1135 -1790 1138 -1784
rect 1142 -1790 1148 -1784
rect 1149 -1790 1152 -1784
rect 1156 -1790 1159 -1784
rect 1163 -1790 1166 -1784
rect 1170 -1790 1173 -1784
rect 1177 -1790 1180 -1784
rect 1184 -1790 1187 -1784
rect 1191 -1790 1194 -1784
rect 1198 -1790 1201 -1784
rect 1205 -1790 1208 -1784
rect 1212 -1790 1215 -1784
rect 1219 -1790 1222 -1784
rect 1226 -1790 1229 -1784
rect 1233 -1790 1236 -1784
rect 1240 -1790 1243 -1784
rect 1247 -1790 1250 -1784
rect 1254 -1790 1257 -1784
rect 1261 -1790 1264 -1784
rect 1268 -1790 1271 -1784
rect 1275 -1790 1278 -1784
rect 1282 -1790 1285 -1784
rect 1289 -1790 1295 -1784
rect 1296 -1790 1299 -1784
rect 1303 -1790 1306 -1784
rect 1310 -1790 1313 -1784
rect 1317 -1790 1320 -1784
rect 1324 -1790 1327 -1784
rect 1331 -1790 1334 -1784
rect 1338 -1790 1341 -1784
rect 1345 -1790 1348 -1784
rect 1352 -1790 1355 -1784
rect 1359 -1790 1362 -1784
rect 1366 -1790 1369 -1784
rect 1373 -1790 1376 -1784
rect 1380 -1790 1383 -1784
rect 1387 -1790 1390 -1784
rect 1394 -1790 1397 -1784
rect 1401 -1790 1404 -1784
rect 1408 -1790 1411 -1784
rect 1415 -1790 1418 -1784
rect 1422 -1790 1425 -1784
rect 1429 -1790 1432 -1784
rect 1436 -1790 1439 -1784
rect 1443 -1790 1446 -1784
rect 1450 -1790 1453 -1784
rect 1457 -1790 1460 -1784
rect 1464 -1790 1467 -1784
rect 1471 -1790 1474 -1784
rect 1478 -1790 1481 -1784
rect 1485 -1790 1488 -1784
rect 1492 -1790 1495 -1784
rect 1499 -1790 1502 -1784
rect 1506 -1790 1509 -1784
rect 1513 -1790 1516 -1784
rect 1520 -1790 1523 -1784
rect 1527 -1790 1530 -1784
rect 1534 -1790 1537 -1784
rect 1541 -1790 1544 -1784
rect 1548 -1790 1551 -1784
rect 1555 -1790 1558 -1784
rect 1562 -1790 1565 -1784
rect 1569 -1790 1572 -1784
rect 1576 -1790 1579 -1784
rect 1583 -1790 1586 -1784
rect 1590 -1790 1593 -1784
rect 1597 -1790 1600 -1784
rect 1604 -1790 1607 -1784
rect 1611 -1790 1614 -1784
rect 1618 -1790 1621 -1784
rect 1625 -1790 1628 -1784
rect 1632 -1790 1635 -1784
rect 1639 -1790 1642 -1784
rect 1646 -1790 1649 -1784
rect 1653 -1790 1656 -1784
rect 1660 -1790 1663 -1784
rect 1667 -1790 1670 -1784
rect 1674 -1790 1677 -1784
rect 1681 -1790 1684 -1784
rect 1688 -1790 1691 -1784
rect 1695 -1790 1698 -1784
rect 1702 -1790 1705 -1784
rect 1709 -1790 1712 -1784
rect 1716 -1790 1719 -1784
rect 1723 -1790 1726 -1784
rect 1730 -1790 1733 -1784
rect 1737 -1790 1740 -1784
rect 1744 -1790 1747 -1784
rect 1751 -1790 1754 -1784
rect 1758 -1790 1761 -1784
rect 1765 -1790 1768 -1784
rect 1772 -1790 1775 -1784
rect 1779 -1790 1782 -1784
rect 1786 -1790 1789 -1784
rect 1793 -1790 1796 -1784
rect 1800 -1790 1803 -1784
rect 1807 -1790 1810 -1784
rect 1814 -1790 1817 -1784
rect 1821 -1790 1824 -1784
rect 1828 -1790 1831 -1784
rect 1835 -1790 1841 -1784
rect 1 -1929 7 -1923
rect 8 -1929 14 -1923
rect 15 -1929 21 -1923
rect 22 -1929 28 -1923
rect 29 -1929 32 -1923
rect 36 -1929 39 -1923
rect 43 -1929 46 -1923
rect 50 -1929 53 -1923
rect 57 -1929 63 -1923
rect 64 -1929 70 -1923
rect 71 -1929 74 -1923
rect 78 -1929 81 -1923
rect 85 -1929 88 -1923
rect 92 -1929 95 -1923
rect 99 -1929 102 -1923
rect 106 -1929 112 -1923
rect 113 -1929 116 -1923
rect 120 -1929 123 -1923
rect 127 -1929 130 -1923
rect 134 -1929 137 -1923
rect 141 -1929 144 -1923
rect 148 -1929 151 -1923
rect 155 -1929 158 -1923
rect 162 -1929 165 -1923
rect 169 -1929 175 -1923
rect 176 -1929 179 -1923
rect 183 -1929 186 -1923
rect 190 -1929 193 -1923
rect 197 -1929 200 -1923
rect 204 -1929 207 -1923
rect 211 -1929 214 -1923
rect 218 -1929 224 -1923
rect 225 -1929 231 -1923
rect 232 -1929 235 -1923
rect 239 -1929 245 -1923
rect 246 -1929 252 -1923
rect 253 -1929 256 -1923
rect 260 -1929 263 -1923
rect 267 -1929 270 -1923
rect 274 -1929 277 -1923
rect 281 -1929 284 -1923
rect 288 -1929 291 -1923
rect 295 -1929 298 -1923
rect 302 -1929 305 -1923
rect 309 -1929 312 -1923
rect 316 -1929 319 -1923
rect 323 -1929 326 -1923
rect 330 -1929 333 -1923
rect 337 -1929 343 -1923
rect 344 -1929 347 -1923
rect 351 -1929 354 -1923
rect 358 -1929 361 -1923
rect 365 -1929 368 -1923
rect 372 -1929 375 -1923
rect 379 -1929 382 -1923
rect 386 -1929 389 -1923
rect 393 -1929 396 -1923
rect 400 -1929 406 -1923
rect 407 -1929 410 -1923
rect 414 -1929 417 -1923
rect 421 -1929 424 -1923
rect 428 -1929 434 -1923
rect 435 -1929 438 -1923
rect 442 -1929 445 -1923
rect 449 -1929 452 -1923
rect 456 -1929 459 -1923
rect 463 -1929 466 -1923
rect 470 -1929 473 -1923
rect 477 -1929 480 -1923
rect 484 -1929 487 -1923
rect 491 -1929 494 -1923
rect 498 -1929 501 -1923
rect 505 -1929 508 -1923
rect 512 -1929 515 -1923
rect 519 -1929 522 -1923
rect 526 -1929 532 -1923
rect 533 -1929 536 -1923
rect 540 -1929 543 -1923
rect 547 -1929 550 -1923
rect 554 -1929 557 -1923
rect 561 -1929 564 -1923
rect 568 -1929 571 -1923
rect 575 -1929 578 -1923
rect 582 -1929 585 -1923
rect 589 -1929 595 -1923
rect 596 -1929 599 -1923
rect 603 -1929 606 -1923
rect 610 -1929 613 -1923
rect 617 -1929 623 -1923
rect 624 -1929 627 -1923
rect 631 -1929 634 -1923
rect 638 -1929 641 -1923
rect 645 -1929 648 -1923
rect 652 -1929 658 -1923
rect 659 -1929 662 -1923
rect 666 -1929 672 -1923
rect 673 -1929 676 -1923
rect 680 -1929 686 -1923
rect 687 -1929 690 -1923
rect 694 -1929 697 -1923
rect 701 -1929 704 -1923
rect 708 -1929 711 -1923
rect 715 -1929 718 -1923
rect 722 -1929 728 -1923
rect 729 -1929 732 -1923
rect 736 -1929 739 -1923
rect 743 -1929 746 -1923
rect 750 -1929 753 -1923
rect 757 -1929 760 -1923
rect 764 -1929 767 -1923
rect 771 -1929 777 -1923
rect 778 -1929 781 -1923
rect 785 -1929 791 -1923
rect 792 -1929 795 -1923
rect 799 -1929 802 -1923
rect 806 -1929 812 -1923
rect 813 -1929 816 -1923
rect 820 -1929 823 -1923
rect 827 -1929 833 -1923
rect 834 -1929 837 -1923
rect 841 -1929 844 -1923
rect 848 -1929 854 -1923
rect 855 -1929 858 -1923
rect 862 -1929 865 -1923
rect 869 -1929 875 -1923
rect 876 -1929 879 -1923
rect 883 -1929 886 -1923
rect 890 -1929 893 -1923
rect 897 -1929 900 -1923
rect 904 -1929 907 -1923
rect 911 -1929 917 -1923
rect 918 -1929 921 -1923
rect 925 -1929 928 -1923
rect 932 -1929 935 -1923
rect 939 -1929 942 -1923
rect 946 -1929 949 -1923
rect 953 -1929 956 -1923
rect 960 -1929 963 -1923
rect 967 -1929 970 -1923
rect 974 -1929 977 -1923
rect 981 -1929 987 -1923
rect 988 -1929 994 -1923
rect 995 -1929 998 -1923
rect 1002 -1929 1005 -1923
rect 1009 -1929 1012 -1923
rect 1016 -1929 1019 -1923
rect 1023 -1929 1026 -1923
rect 1030 -1929 1033 -1923
rect 1037 -1929 1040 -1923
rect 1044 -1929 1047 -1923
rect 1051 -1929 1054 -1923
rect 1058 -1929 1061 -1923
rect 1065 -1929 1068 -1923
rect 1072 -1929 1075 -1923
rect 1079 -1929 1082 -1923
rect 1086 -1929 1089 -1923
rect 1093 -1929 1099 -1923
rect 1100 -1929 1103 -1923
rect 1107 -1929 1110 -1923
rect 1114 -1929 1117 -1923
rect 1121 -1929 1127 -1923
rect 1128 -1929 1131 -1923
rect 1135 -1929 1138 -1923
rect 1142 -1929 1145 -1923
rect 1149 -1929 1152 -1923
rect 1156 -1929 1162 -1923
rect 1163 -1929 1169 -1923
rect 1170 -1929 1173 -1923
rect 1177 -1929 1180 -1923
rect 1184 -1929 1187 -1923
rect 1191 -1929 1194 -1923
rect 1198 -1929 1201 -1923
rect 1205 -1929 1208 -1923
rect 1212 -1929 1215 -1923
rect 1219 -1929 1222 -1923
rect 1226 -1929 1232 -1923
rect 1233 -1929 1236 -1923
rect 1240 -1929 1243 -1923
rect 1247 -1929 1250 -1923
rect 1254 -1929 1257 -1923
rect 1261 -1929 1264 -1923
rect 1268 -1929 1271 -1923
rect 1275 -1929 1278 -1923
rect 1282 -1929 1285 -1923
rect 1289 -1929 1292 -1923
rect 1296 -1929 1299 -1923
rect 1303 -1929 1306 -1923
rect 1310 -1929 1313 -1923
rect 1317 -1929 1320 -1923
rect 1324 -1929 1327 -1923
rect 1331 -1929 1334 -1923
rect 1338 -1929 1341 -1923
rect 1345 -1929 1348 -1923
rect 1352 -1929 1355 -1923
rect 1359 -1929 1362 -1923
rect 1366 -1929 1369 -1923
rect 1373 -1929 1376 -1923
rect 1380 -1929 1386 -1923
rect 1387 -1929 1390 -1923
rect 1394 -1929 1397 -1923
rect 1401 -1929 1404 -1923
rect 1408 -1929 1411 -1923
rect 1415 -1929 1418 -1923
rect 1422 -1929 1425 -1923
rect 1429 -1929 1432 -1923
rect 1436 -1929 1439 -1923
rect 1443 -1929 1446 -1923
rect 1450 -1929 1453 -1923
rect 1457 -1929 1460 -1923
rect 1464 -1929 1467 -1923
rect 1471 -1929 1474 -1923
rect 1478 -1929 1481 -1923
rect 1485 -1929 1488 -1923
rect 1492 -1929 1495 -1923
rect 1499 -1929 1502 -1923
rect 1506 -1929 1509 -1923
rect 1513 -1929 1516 -1923
rect 1520 -1929 1523 -1923
rect 1527 -1929 1530 -1923
rect 1534 -1929 1537 -1923
rect 1541 -1929 1544 -1923
rect 1548 -1929 1551 -1923
rect 1555 -1929 1558 -1923
rect 1562 -1929 1565 -1923
rect 1569 -1929 1572 -1923
rect 1576 -1929 1579 -1923
rect 1583 -1929 1586 -1923
rect 1590 -1929 1593 -1923
rect 1597 -1929 1600 -1923
rect 1604 -1929 1607 -1923
rect 1611 -1929 1614 -1923
rect 1618 -1929 1621 -1923
rect 1625 -1929 1628 -1923
rect 1632 -1929 1635 -1923
rect 1639 -1929 1642 -1923
rect 1646 -1929 1649 -1923
rect 1653 -1929 1656 -1923
rect 1660 -1929 1663 -1923
rect 1667 -1929 1670 -1923
rect 1674 -1929 1677 -1923
rect 1681 -1929 1684 -1923
rect 1688 -1929 1691 -1923
rect 1695 -1929 1698 -1923
rect 1702 -1929 1705 -1923
rect 1709 -1929 1712 -1923
rect 1716 -1929 1719 -1923
rect 1723 -1929 1726 -1923
rect 1730 -1929 1733 -1923
rect 1737 -1929 1740 -1923
rect 1744 -1929 1747 -1923
rect 1751 -1929 1757 -1923
rect 1758 -1929 1761 -1923
rect 1765 -1929 1768 -1923
rect 1793 -1929 1796 -1923
rect 1 -2056 7 -2050
rect 8 -2056 14 -2050
rect 15 -2056 21 -2050
rect 22 -2056 25 -2050
rect 29 -2056 35 -2050
rect 36 -2056 39 -2050
rect 43 -2056 46 -2050
rect 50 -2056 53 -2050
rect 57 -2056 60 -2050
rect 64 -2056 67 -2050
rect 71 -2056 74 -2050
rect 78 -2056 81 -2050
rect 85 -2056 88 -2050
rect 92 -2056 95 -2050
rect 99 -2056 102 -2050
rect 106 -2056 112 -2050
rect 113 -2056 119 -2050
rect 120 -2056 123 -2050
rect 127 -2056 133 -2050
rect 134 -2056 140 -2050
rect 141 -2056 144 -2050
rect 148 -2056 151 -2050
rect 155 -2056 161 -2050
rect 162 -2056 168 -2050
rect 169 -2056 172 -2050
rect 176 -2056 179 -2050
rect 183 -2056 186 -2050
rect 190 -2056 193 -2050
rect 197 -2056 200 -2050
rect 204 -2056 210 -2050
rect 211 -2056 214 -2050
rect 218 -2056 221 -2050
rect 225 -2056 228 -2050
rect 232 -2056 235 -2050
rect 239 -2056 242 -2050
rect 246 -2056 249 -2050
rect 253 -2056 256 -2050
rect 260 -2056 263 -2050
rect 267 -2056 270 -2050
rect 274 -2056 277 -2050
rect 281 -2056 284 -2050
rect 288 -2056 291 -2050
rect 295 -2056 298 -2050
rect 302 -2056 305 -2050
rect 309 -2056 312 -2050
rect 316 -2056 319 -2050
rect 323 -2056 326 -2050
rect 330 -2056 333 -2050
rect 337 -2056 340 -2050
rect 344 -2056 347 -2050
rect 351 -2056 354 -2050
rect 358 -2056 361 -2050
rect 365 -2056 371 -2050
rect 372 -2056 375 -2050
rect 379 -2056 382 -2050
rect 386 -2056 389 -2050
rect 393 -2056 396 -2050
rect 400 -2056 403 -2050
rect 407 -2056 410 -2050
rect 414 -2056 417 -2050
rect 421 -2056 424 -2050
rect 428 -2056 431 -2050
rect 435 -2056 438 -2050
rect 442 -2056 445 -2050
rect 449 -2056 452 -2050
rect 456 -2056 459 -2050
rect 463 -2056 466 -2050
rect 470 -2056 473 -2050
rect 477 -2056 480 -2050
rect 484 -2056 487 -2050
rect 491 -2056 494 -2050
rect 498 -2056 501 -2050
rect 505 -2056 508 -2050
rect 512 -2056 515 -2050
rect 519 -2056 522 -2050
rect 526 -2056 532 -2050
rect 533 -2056 536 -2050
rect 540 -2056 543 -2050
rect 547 -2056 550 -2050
rect 554 -2056 557 -2050
rect 561 -2056 564 -2050
rect 568 -2056 571 -2050
rect 575 -2056 578 -2050
rect 582 -2056 585 -2050
rect 589 -2056 595 -2050
rect 596 -2056 602 -2050
rect 603 -2056 609 -2050
rect 610 -2056 613 -2050
rect 617 -2056 623 -2050
rect 624 -2056 627 -2050
rect 631 -2056 637 -2050
rect 638 -2056 641 -2050
rect 645 -2056 648 -2050
rect 652 -2056 655 -2050
rect 659 -2056 665 -2050
rect 666 -2056 672 -2050
rect 673 -2056 676 -2050
rect 680 -2056 683 -2050
rect 687 -2056 693 -2050
rect 694 -2056 697 -2050
rect 701 -2056 704 -2050
rect 708 -2056 711 -2050
rect 715 -2056 718 -2050
rect 722 -2056 725 -2050
rect 729 -2056 732 -2050
rect 736 -2056 739 -2050
rect 743 -2056 746 -2050
rect 750 -2056 756 -2050
rect 757 -2056 760 -2050
rect 764 -2056 770 -2050
rect 771 -2056 774 -2050
rect 778 -2056 784 -2050
rect 785 -2056 788 -2050
rect 792 -2056 795 -2050
rect 799 -2056 805 -2050
rect 806 -2056 809 -2050
rect 813 -2056 819 -2050
rect 820 -2056 823 -2050
rect 827 -2056 830 -2050
rect 834 -2056 837 -2050
rect 841 -2056 844 -2050
rect 848 -2056 851 -2050
rect 855 -2056 858 -2050
rect 862 -2056 865 -2050
rect 869 -2056 872 -2050
rect 876 -2056 879 -2050
rect 883 -2056 886 -2050
rect 890 -2056 893 -2050
rect 897 -2056 900 -2050
rect 904 -2056 910 -2050
rect 911 -2056 914 -2050
rect 918 -2056 921 -2050
rect 925 -2056 931 -2050
rect 932 -2056 938 -2050
rect 939 -2056 942 -2050
rect 946 -2056 952 -2050
rect 953 -2056 956 -2050
rect 960 -2056 963 -2050
rect 967 -2056 970 -2050
rect 974 -2056 977 -2050
rect 981 -2056 987 -2050
rect 988 -2056 991 -2050
rect 995 -2056 998 -2050
rect 1002 -2056 1005 -2050
rect 1009 -2056 1012 -2050
rect 1016 -2056 1022 -2050
rect 1023 -2056 1026 -2050
rect 1030 -2056 1033 -2050
rect 1037 -2056 1040 -2050
rect 1044 -2056 1047 -2050
rect 1051 -2056 1054 -2050
rect 1058 -2056 1061 -2050
rect 1065 -2056 1068 -2050
rect 1072 -2056 1075 -2050
rect 1079 -2056 1082 -2050
rect 1086 -2056 1092 -2050
rect 1093 -2056 1096 -2050
rect 1100 -2056 1103 -2050
rect 1107 -2056 1110 -2050
rect 1114 -2056 1117 -2050
rect 1121 -2056 1124 -2050
rect 1128 -2056 1131 -2050
rect 1135 -2056 1138 -2050
rect 1142 -2056 1145 -2050
rect 1149 -2056 1152 -2050
rect 1156 -2056 1159 -2050
rect 1163 -2056 1166 -2050
rect 1170 -2056 1173 -2050
rect 1177 -2056 1180 -2050
rect 1184 -2056 1187 -2050
rect 1191 -2056 1194 -2050
rect 1198 -2056 1201 -2050
rect 1205 -2056 1208 -2050
rect 1212 -2056 1215 -2050
rect 1219 -2056 1222 -2050
rect 1226 -2056 1229 -2050
rect 1233 -2056 1236 -2050
rect 1240 -2056 1243 -2050
rect 1247 -2056 1250 -2050
rect 1254 -2056 1260 -2050
rect 1261 -2056 1264 -2050
rect 1268 -2056 1271 -2050
rect 1275 -2056 1278 -2050
rect 1282 -2056 1285 -2050
rect 1289 -2056 1292 -2050
rect 1296 -2056 1299 -2050
rect 1303 -2056 1306 -2050
rect 1310 -2056 1313 -2050
rect 1317 -2056 1320 -2050
rect 1324 -2056 1327 -2050
rect 1331 -2056 1334 -2050
rect 1338 -2056 1341 -2050
rect 1345 -2056 1348 -2050
rect 1352 -2056 1355 -2050
rect 1359 -2056 1362 -2050
rect 1366 -2056 1369 -2050
rect 1373 -2056 1376 -2050
rect 1380 -2056 1383 -2050
rect 1387 -2056 1390 -2050
rect 1394 -2056 1397 -2050
rect 1401 -2056 1404 -2050
rect 1408 -2056 1411 -2050
rect 1415 -2056 1418 -2050
rect 1422 -2056 1425 -2050
rect 1429 -2056 1432 -2050
rect 1436 -2056 1439 -2050
rect 1443 -2056 1446 -2050
rect 1450 -2056 1456 -2050
rect 1457 -2056 1460 -2050
rect 1464 -2056 1467 -2050
rect 1471 -2056 1474 -2050
rect 1478 -2056 1481 -2050
rect 1485 -2056 1488 -2050
rect 1492 -2056 1495 -2050
rect 1499 -2056 1502 -2050
rect 1506 -2056 1509 -2050
rect 1513 -2056 1516 -2050
rect 1520 -2056 1523 -2050
rect 1527 -2056 1530 -2050
rect 1534 -2056 1537 -2050
rect 1541 -2056 1544 -2050
rect 1548 -2056 1551 -2050
rect 1555 -2056 1558 -2050
rect 1562 -2056 1565 -2050
rect 1569 -2056 1572 -2050
rect 1576 -2056 1579 -2050
rect 1583 -2056 1586 -2050
rect 1590 -2056 1593 -2050
rect 1597 -2056 1600 -2050
rect 1604 -2056 1607 -2050
rect 1611 -2056 1614 -2050
rect 1618 -2056 1621 -2050
rect 1625 -2056 1628 -2050
rect 1632 -2056 1635 -2050
rect 1639 -2056 1642 -2050
rect 1646 -2056 1649 -2050
rect 1653 -2056 1656 -2050
rect 1660 -2056 1663 -2050
rect 1667 -2056 1670 -2050
rect 1674 -2056 1677 -2050
rect 1681 -2056 1684 -2050
rect 1688 -2056 1691 -2050
rect 1695 -2056 1698 -2050
rect 1702 -2056 1705 -2050
rect 1709 -2056 1712 -2050
rect 1716 -2056 1719 -2050
rect 1723 -2056 1726 -2050
rect 1730 -2056 1733 -2050
rect 1737 -2056 1740 -2050
rect 1744 -2056 1750 -2050
rect 1751 -2056 1757 -2050
rect 1758 -2056 1764 -2050
rect 1765 -2056 1768 -2050
rect 1772 -2056 1775 -2050
rect 1 -2195 7 -2189
rect 8 -2195 14 -2189
rect 15 -2195 21 -2189
rect 22 -2195 28 -2189
rect 29 -2195 32 -2189
rect 36 -2195 42 -2189
rect 43 -2195 49 -2189
rect 50 -2195 56 -2189
rect 57 -2195 60 -2189
rect 64 -2195 70 -2189
rect 71 -2195 74 -2189
rect 78 -2195 81 -2189
rect 85 -2195 91 -2189
rect 92 -2195 98 -2189
rect 99 -2195 102 -2189
rect 106 -2195 109 -2189
rect 113 -2195 116 -2189
rect 120 -2195 123 -2189
rect 127 -2195 133 -2189
rect 134 -2195 137 -2189
rect 141 -2195 144 -2189
rect 148 -2195 154 -2189
rect 155 -2195 158 -2189
rect 162 -2195 165 -2189
rect 169 -2195 175 -2189
rect 176 -2195 179 -2189
rect 183 -2195 186 -2189
rect 190 -2195 193 -2189
rect 197 -2195 200 -2189
rect 204 -2195 207 -2189
rect 211 -2195 214 -2189
rect 218 -2195 221 -2189
rect 225 -2195 231 -2189
rect 232 -2195 235 -2189
rect 239 -2195 242 -2189
rect 246 -2195 249 -2189
rect 253 -2195 256 -2189
rect 260 -2195 263 -2189
rect 267 -2195 273 -2189
rect 274 -2195 277 -2189
rect 281 -2195 284 -2189
rect 288 -2195 291 -2189
rect 295 -2195 298 -2189
rect 302 -2195 305 -2189
rect 309 -2195 312 -2189
rect 316 -2195 319 -2189
rect 323 -2195 326 -2189
rect 330 -2195 333 -2189
rect 337 -2195 340 -2189
rect 344 -2195 347 -2189
rect 351 -2195 354 -2189
rect 358 -2195 364 -2189
rect 365 -2195 368 -2189
rect 372 -2195 375 -2189
rect 379 -2195 382 -2189
rect 386 -2195 389 -2189
rect 393 -2195 396 -2189
rect 400 -2195 403 -2189
rect 407 -2195 413 -2189
rect 414 -2195 417 -2189
rect 421 -2195 424 -2189
rect 428 -2195 431 -2189
rect 435 -2195 438 -2189
rect 442 -2195 445 -2189
rect 449 -2195 455 -2189
rect 456 -2195 459 -2189
rect 463 -2195 466 -2189
rect 470 -2195 473 -2189
rect 477 -2195 480 -2189
rect 484 -2195 487 -2189
rect 491 -2195 494 -2189
rect 498 -2195 501 -2189
rect 505 -2195 508 -2189
rect 512 -2195 515 -2189
rect 519 -2195 525 -2189
rect 526 -2195 529 -2189
rect 533 -2195 536 -2189
rect 540 -2195 543 -2189
rect 547 -2195 550 -2189
rect 554 -2195 557 -2189
rect 561 -2195 564 -2189
rect 568 -2195 571 -2189
rect 575 -2195 578 -2189
rect 582 -2195 585 -2189
rect 589 -2195 592 -2189
rect 596 -2195 599 -2189
rect 603 -2195 609 -2189
rect 610 -2195 613 -2189
rect 617 -2195 623 -2189
rect 624 -2195 627 -2189
rect 631 -2195 634 -2189
rect 638 -2195 641 -2189
rect 645 -2195 648 -2189
rect 652 -2195 655 -2189
rect 659 -2195 662 -2189
rect 666 -2195 669 -2189
rect 673 -2195 676 -2189
rect 680 -2195 683 -2189
rect 687 -2195 690 -2189
rect 694 -2195 697 -2189
rect 701 -2195 707 -2189
rect 708 -2195 711 -2189
rect 715 -2195 718 -2189
rect 722 -2195 728 -2189
rect 729 -2195 735 -2189
rect 736 -2195 739 -2189
rect 743 -2195 749 -2189
rect 750 -2195 753 -2189
rect 757 -2195 763 -2189
rect 764 -2195 767 -2189
rect 771 -2195 777 -2189
rect 778 -2195 781 -2189
rect 785 -2195 788 -2189
rect 792 -2195 798 -2189
rect 799 -2195 802 -2189
rect 806 -2195 809 -2189
rect 813 -2195 819 -2189
rect 820 -2195 823 -2189
rect 827 -2195 833 -2189
rect 834 -2195 837 -2189
rect 841 -2195 844 -2189
rect 848 -2195 851 -2189
rect 855 -2195 858 -2189
rect 862 -2195 865 -2189
rect 869 -2195 875 -2189
rect 876 -2195 879 -2189
rect 883 -2195 886 -2189
rect 890 -2195 893 -2189
rect 897 -2195 900 -2189
rect 904 -2195 907 -2189
rect 911 -2195 914 -2189
rect 918 -2195 921 -2189
rect 925 -2195 928 -2189
rect 932 -2195 938 -2189
rect 939 -2195 942 -2189
rect 946 -2195 949 -2189
rect 953 -2195 956 -2189
rect 960 -2195 963 -2189
rect 967 -2195 970 -2189
rect 974 -2195 980 -2189
rect 981 -2195 984 -2189
rect 988 -2195 991 -2189
rect 995 -2195 1001 -2189
rect 1002 -2195 1005 -2189
rect 1009 -2195 1015 -2189
rect 1016 -2195 1019 -2189
rect 1023 -2195 1026 -2189
rect 1030 -2195 1033 -2189
rect 1037 -2195 1040 -2189
rect 1044 -2195 1047 -2189
rect 1051 -2195 1054 -2189
rect 1058 -2195 1061 -2189
rect 1065 -2195 1068 -2189
rect 1072 -2195 1075 -2189
rect 1079 -2195 1082 -2189
rect 1086 -2195 1089 -2189
rect 1093 -2195 1096 -2189
rect 1100 -2195 1106 -2189
rect 1107 -2195 1110 -2189
rect 1114 -2195 1120 -2189
rect 1121 -2195 1124 -2189
rect 1128 -2195 1131 -2189
rect 1135 -2195 1138 -2189
rect 1142 -2195 1145 -2189
rect 1149 -2195 1152 -2189
rect 1156 -2195 1159 -2189
rect 1163 -2195 1166 -2189
rect 1170 -2195 1173 -2189
rect 1177 -2195 1180 -2189
rect 1184 -2195 1187 -2189
rect 1191 -2195 1194 -2189
rect 1198 -2195 1201 -2189
rect 1205 -2195 1208 -2189
rect 1212 -2195 1215 -2189
rect 1219 -2195 1222 -2189
rect 1226 -2195 1229 -2189
rect 1233 -2195 1236 -2189
rect 1240 -2195 1243 -2189
rect 1247 -2195 1250 -2189
rect 1254 -2195 1257 -2189
rect 1261 -2195 1264 -2189
rect 1268 -2195 1271 -2189
rect 1275 -2195 1278 -2189
rect 1282 -2195 1285 -2189
rect 1289 -2195 1292 -2189
rect 1296 -2195 1299 -2189
rect 1303 -2195 1306 -2189
rect 1310 -2195 1313 -2189
rect 1317 -2195 1320 -2189
rect 1324 -2195 1327 -2189
rect 1331 -2195 1334 -2189
rect 1338 -2195 1341 -2189
rect 1345 -2195 1348 -2189
rect 1352 -2195 1355 -2189
rect 1359 -2195 1362 -2189
rect 1366 -2195 1369 -2189
rect 1373 -2195 1376 -2189
rect 1380 -2195 1383 -2189
rect 1387 -2195 1390 -2189
rect 1394 -2195 1397 -2189
rect 1401 -2195 1404 -2189
rect 1408 -2195 1411 -2189
rect 1415 -2195 1418 -2189
rect 1422 -2195 1425 -2189
rect 1429 -2195 1432 -2189
rect 1436 -2195 1439 -2189
rect 1443 -2195 1446 -2189
rect 1450 -2195 1453 -2189
rect 1457 -2195 1460 -2189
rect 1464 -2195 1467 -2189
rect 1471 -2195 1474 -2189
rect 1478 -2195 1481 -2189
rect 1485 -2195 1488 -2189
rect 1492 -2195 1495 -2189
rect 1499 -2195 1502 -2189
rect 1506 -2195 1509 -2189
rect 1513 -2195 1516 -2189
rect 1520 -2195 1523 -2189
rect 1527 -2195 1530 -2189
rect 1534 -2195 1537 -2189
rect 1541 -2195 1544 -2189
rect 1548 -2195 1551 -2189
rect 1555 -2195 1558 -2189
rect 1562 -2195 1565 -2189
rect 1569 -2195 1572 -2189
rect 1576 -2195 1579 -2189
rect 1583 -2195 1586 -2189
rect 1590 -2195 1593 -2189
rect 1597 -2195 1600 -2189
rect 1604 -2195 1607 -2189
rect 1611 -2195 1614 -2189
rect 1618 -2195 1621 -2189
rect 1625 -2195 1628 -2189
rect 1632 -2195 1635 -2189
rect 1639 -2195 1642 -2189
rect 1646 -2195 1649 -2189
rect 1653 -2195 1656 -2189
rect 1660 -2195 1663 -2189
rect 1667 -2195 1670 -2189
rect 1674 -2195 1677 -2189
rect 1681 -2195 1684 -2189
rect 1688 -2195 1691 -2189
rect 1695 -2195 1698 -2189
rect 1702 -2195 1705 -2189
rect 1709 -2195 1712 -2189
rect 1716 -2195 1719 -2189
rect 1723 -2195 1726 -2189
rect 1730 -2195 1733 -2189
rect 1737 -2195 1740 -2189
rect 1744 -2195 1747 -2189
rect 1751 -2195 1757 -2189
rect 1758 -2195 1761 -2189
rect 1765 -2195 1768 -2189
rect 1 -2330 7 -2324
rect 8 -2330 14 -2324
rect 15 -2330 21 -2324
rect 22 -2330 28 -2324
rect 29 -2330 35 -2324
rect 36 -2330 42 -2324
rect 43 -2330 46 -2324
rect 50 -2330 53 -2324
rect 57 -2330 60 -2324
rect 64 -2330 67 -2324
rect 71 -2330 74 -2324
rect 78 -2330 81 -2324
rect 85 -2330 91 -2324
rect 92 -2330 98 -2324
rect 99 -2330 102 -2324
rect 106 -2330 109 -2324
rect 113 -2330 119 -2324
rect 120 -2330 123 -2324
rect 127 -2330 130 -2324
rect 134 -2330 140 -2324
rect 141 -2330 144 -2324
rect 148 -2330 151 -2324
rect 155 -2330 158 -2324
rect 162 -2330 165 -2324
rect 169 -2330 175 -2324
rect 176 -2330 179 -2324
rect 183 -2330 186 -2324
rect 190 -2330 193 -2324
rect 197 -2330 200 -2324
rect 204 -2330 207 -2324
rect 211 -2330 217 -2324
rect 218 -2330 221 -2324
rect 225 -2330 228 -2324
rect 232 -2330 238 -2324
rect 239 -2330 242 -2324
rect 246 -2330 249 -2324
rect 253 -2330 256 -2324
rect 260 -2330 263 -2324
rect 267 -2330 270 -2324
rect 274 -2330 277 -2324
rect 281 -2330 284 -2324
rect 288 -2330 291 -2324
rect 295 -2330 298 -2324
rect 302 -2330 305 -2324
rect 309 -2330 312 -2324
rect 316 -2330 319 -2324
rect 323 -2330 326 -2324
rect 330 -2330 333 -2324
rect 337 -2330 340 -2324
rect 344 -2330 347 -2324
rect 351 -2330 354 -2324
rect 358 -2330 361 -2324
rect 365 -2330 368 -2324
rect 372 -2330 375 -2324
rect 379 -2330 382 -2324
rect 386 -2330 389 -2324
rect 393 -2330 396 -2324
rect 400 -2330 403 -2324
rect 407 -2330 410 -2324
rect 414 -2330 417 -2324
rect 421 -2330 424 -2324
rect 428 -2330 431 -2324
rect 435 -2330 438 -2324
rect 442 -2330 445 -2324
rect 449 -2330 452 -2324
rect 456 -2330 459 -2324
rect 463 -2330 466 -2324
rect 470 -2330 473 -2324
rect 477 -2330 480 -2324
rect 484 -2330 487 -2324
rect 491 -2330 494 -2324
rect 498 -2330 501 -2324
rect 505 -2330 508 -2324
rect 512 -2330 515 -2324
rect 519 -2330 522 -2324
rect 526 -2330 529 -2324
rect 533 -2330 539 -2324
rect 540 -2330 543 -2324
rect 547 -2330 550 -2324
rect 554 -2330 557 -2324
rect 561 -2330 564 -2324
rect 568 -2330 571 -2324
rect 575 -2330 578 -2324
rect 582 -2330 588 -2324
rect 589 -2330 592 -2324
rect 596 -2330 599 -2324
rect 603 -2330 606 -2324
rect 610 -2330 613 -2324
rect 617 -2330 620 -2324
rect 624 -2330 627 -2324
rect 631 -2330 634 -2324
rect 638 -2330 644 -2324
rect 645 -2330 648 -2324
rect 652 -2330 658 -2324
rect 659 -2330 662 -2324
rect 666 -2330 669 -2324
rect 673 -2330 676 -2324
rect 680 -2330 683 -2324
rect 687 -2330 693 -2324
rect 694 -2330 697 -2324
rect 701 -2330 707 -2324
rect 708 -2330 711 -2324
rect 715 -2330 718 -2324
rect 722 -2330 725 -2324
rect 729 -2330 735 -2324
rect 736 -2330 739 -2324
rect 743 -2330 749 -2324
rect 750 -2330 753 -2324
rect 757 -2330 760 -2324
rect 764 -2330 767 -2324
rect 771 -2330 777 -2324
rect 778 -2330 781 -2324
rect 785 -2330 788 -2324
rect 792 -2330 795 -2324
rect 799 -2330 802 -2324
rect 806 -2330 809 -2324
rect 813 -2330 816 -2324
rect 820 -2330 823 -2324
rect 827 -2330 830 -2324
rect 834 -2330 837 -2324
rect 841 -2330 844 -2324
rect 848 -2330 854 -2324
rect 855 -2330 858 -2324
rect 862 -2330 865 -2324
rect 869 -2330 875 -2324
rect 876 -2330 879 -2324
rect 883 -2330 886 -2324
rect 890 -2330 893 -2324
rect 897 -2330 903 -2324
rect 904 -2330 907 -2324
rect 911 -2330 914 -2324
rect 918 -2330 921 -2324
rect 925 -2330 928 -2324
rect 932 -2330 935 -2324
rect 939 -2330 942 -2324
rect 946 -2330 949 -2324
rect 953 -2330 959 -2324
rect 960 -2330 963 -2324
rect 967 -2330 973 -2324
rect 974 -2330 977 -2324
rect 981 -2330 984 -2324
rect 988 -2330 991 -2324
rect 995 -2330 1001 -2324
rect 1002 -2330 1005 -2324
rect 1009 -2330 1012 -2324
rect 1016 -2330 1019 -2324
rect 1023 -2330 1026 -2324
rect 1030 -2330 1033 -2324
rect 1037 -2330 1040 -2324
rect 1044 -2330 1047 -2324
rect 1051 -2330 1054 -2324
rect 1058 -2330 1061 -2324
rect 1065 -2330 1068 -2324
rect 1072 -2330 1075 -2324
rect 1079 -2330 1085 -2324
rect 1086 -2330 1089 -2324
rect 1093 -2330 1099 -2324
rect 1100 -2330 1103 -2324
rect 1107 -2330 1110 -2324
rect 1114 -2330 1117 -2324
rect 1121 -2330 1127 -2324
rect 1128 -2330 1131 -2324
rect 1135 -2330 1138 -2324
rect 1142 -2330 1148 -2324
rect 1149 -2330 1152 -2324
rect 1156 -2330 1159 -2324
rect 1163 -2330 1166 -2324
rect 1170 -2330 1176 -2324
rect 1177 -2330 1180 -2324
rect 1184 -2330 1187 -2324
rect 1191 -2330 1194 -2324
rect 1198 -2330 1201 -2324
rect 1205 -2330 1208 -2324
rect 1212 -2330 1215 -2324
rect 1219 -2330 1222 -2324
rect 1226 -2330 1229 -2324
rect 1233 -2330 1239 -2324
rect 1240 -2330 1243 -2324
rect 1247 -2330 1250 -2324
rect 1254 -2330 1257 -2324
rect 1261 -2330 1264 -2324
rect 1268 -2330 1271 -2324
rect 1275 -2330 1278 -2324
rect 1282 -2330 1285 -2324
rect 1289 -2330 1292 -2324
rect 1296 -2330 1299 -2324
rect 1303 -2330 1309 -2324
rect 1310 -2330 1313 -2324
rect 1317 -2330 1320 -2324
rect 1324 -2330 1327 -2324
rect 1331 -2330 1337 -2324
rect 1338 -2330 1341 -2324
rect 1345 -2330 1348 -2324
rect 1352 -2330 1355 -2324
rect 1359 -2330 1362 -2324
rect 1366 -2330 1369 -2324
rect 1373 -2330 1376 -2324
rect 1380 -2330 1383 -2324
rect 1387 -2330 1390 -2324
rect 1394 -2330 1397 -2324
rect 1401 -2330 1404 -2324
rect 1408 -2330 1411 -2324
rect 1415 -2330 1418 -2324
rect 1422 -2330 1425 -2324
rect 1429 -2330 1432 -2324
rect 1436 -2330 1439 -2324
rect 1443 -2330 1446 -2324
rect 1450 -2330 1453 -2324
rect 1457 -2330 1460 -2324
rect 1464 -2330 1467 -2324
rect 1471 -2330 1474 -2324
rect 1478 -2330 1481 -2324
rect 1485 -2330 1488 -2324
rect 1492 -2330 1495 -2324
rect 1499 -2330 1502 -2324
rect 1506 -2330 1509 -2324
rect 1513 -2330 1516 -2324
rect 1520 -2330 1523 -2324
rect 1527 -2330 1530 -2324
rect 1534 -2330 1537 -2324
rect 1541 -2330 1544 -2324
rect 1548 -2330 1551 -2324
rect 1555 -2330 1558 -2324
rect 1562 -2330 1565 -2324
rect 1569 -2330 1572 -2324
rect 1576 -2330 1579 -2324
rect 1583 -2330 1586 -2324
rect 1590 -2330 1593 -2324
rect 1597 -2330 1600 -2324
rect 1604 -2330 1607 -2324
rect 1611 -2330 1614 -2324
rect 1618 -2330 1621 -2324
rect 1625 -2330 1628 -2324
rect 1632 -2330 1635 -2324
rect 1639 -2330 1642 -2324
rect 1646 -2330 1649 -2324
rect 1653 -2330 1656 -2324
rect 1660 -2330 1663 -2324
rect 1667 -2330 1670 -2324
rect 1674 -2330 1677 -2324
rect 1681 -2330 1684 -2324
rect 1688 -2330 1691 -2324
rect 1695 -2330 1698 -2324
rect 1702 -2330 1708 -2324
rect 1709 -2330 1715 -2324
rect 1716 -2330 1719 -2324
rect 1723 -2330 1726 -2324
rect 1730 -2330 1733 -2324
rect 1737 -2330 1740 -2324
rect 1 -2445 7 -2439
rect 8 -2445 14 -2439
rect 15 -2445 21 -2439
rect 22 -2445 28 -2439
rect 29 -2445 35 -2439
rect 50 -2445 53 -2439
rect 57 -2445 60 -2439
rect 64 -2445 67 -2439
rect 71 -2445 74 -2439
rect 78 -2445 81 -2439
rect 85 -2445 88 -2439
rect 92 -2445 95 -2439
rect 99 -2445 102 -2439
rect 106 -2445 109 -2439
rect 113 -2445 116 -2439
rect 120 -2445 123 -2439
rect 127 -2445 130 -2439
rect 134 -2445 137 -2439
rect 141 -2445 144 -2439
rect 148 -2445 151 -2439
rect 155 -2445 158 -2439
rect 162 -2445 165 -2439
rect 169 -2445 172 -2439
rect 176 -2445 182 -2439
rect 183 -2445 186 -2439
rect 190 -2445 193 -2439
rect 197 -2445 200 -2439
rect 204 -2445 207 -2439
rect 211 -2445 217 -2439
rect 218 -2445 221 -2439
rect 225 -2445 228 -2439
rect 232 -2445 235 -2439
rect 239 -2445 242 -2439
rect 246 -2445 249 -2439
rect 253 -2445 259 -2439
rect 260 -2445 263 -2439
rect 267 -2445 270 -2439
rect 274 -2445 277 -2439
rect 281 -2445 284 -2439
rect 288 -2445 291 -2439
rect 295 -2445 298 -2439
rect 302 -2445 305 -2439
rect 309 -2445 315 -2439
rect 316 -2445 319 -2439
rect 323 -2445 326 -2439
rect 330 -2445 333 -2439
rect 337 -2445 340 -2439
rect 344 -2445 347 -2439
rect 351 -2445 354 -2439
rect 358 -2445 361 -2439
rect 365 -2445 368 -2439
rect 372 -2445 375 -2439
rect 379 -2445 382 -2439
rect 386 -2445 389 -2439
rect 393 -2445 396 -2439
rect 400 -2445 403 -2439
rect 407 -2445 410 -2439
rect 414 -2445 417 -2439
rect 421 -2445 424 -2439
rect 428 -2445 434 -2439
rect 435 -2445 438 -2439
rect 442 -2445 445 -2439
rect 449 -2445 452 -2439
rect 456 -2445 459 -2439
rect 463 -2445 466 -2439
rect 470 -2445 476 -2439
rect 477 -2445 480 -2439
rect 484 -2445 487 -2439
rect 491 -2445 494 -2439
rect 498 -2445 504 -2439
rect 505 -2445 508 -2439
rect 512 -2445 515 -2439
rect 519 -2445 522 -2439
rect 526 -2445 532 -2439
rect 533 -2445 536 -2439
rect 540 -2445 546 -2439
rect 547 -2445 550 -2439
rect 554 -2445 557 -2439
rect 561 -2445 564 -2439
rect 568 -2445 571 -2439
rect 575 -2445 578 -2439
rect 582 -2445 585 -2439
rect 589 -2445 592 -2439
rect 596 -2445 599 -2439
rect 603 -2445 606 -2439
rect 610 -2445 616 -2439
rect 617 -2445 620 -2439
rect 624 -2445 627 -2439
rect 631 -2445 634 -2439
rect 638 -2445 644 -2439
rect 645 -2445 648 -2439
rect 652 -2445 655 -2439
rect 659 -2445 662 -2439
rect 666 -2445 669 -2439
rect 673 -2445 679 -2439
rect 680 -2445 686 -2439
rect 687 -2445 690 -2439
rect 694 -2445 697 -2439
rect 701 -2445 707 -2439
rect 708 -2445 711 -2439
rect 715 -2445 718 -2439
rect 722 -2445 725 -2439
rect 729 -2445 735 -2439
rect 736 -2445 739 -2439
rect 743 -2445 749 -2439
rect 750 -2445 753 -2439
rect 757 -2445 760 -2439
rect 764 -2445 767 -2439
rect 771 -2445 774 -2439
rect 778 -2445 781 -2439
rect 785 -2445 788 -2439
rect 792 -2445 795 -2439
rect 799 -2445 802 -2439
rect 806 -2445 812 -2439
rect 813 -2445 816 -2439
rect 820 -2445 826 -2439
rect 827 -2445 830 -2439
rect 834 -2445 837 -2439
rect 841 -2445 847 -2439
rect 848 -2445 854 -2439
rect 855 -2445 861 -2439
rect 862 -2445 865 -2439
rect 869 -2445 872 -2439
rect 876 -2445 879 -2439
rect 883 -2445 886 -2439
rect 890 -2445 896 -2439
rect 897 -2445 903 -2439
rect 904 -2445 907 -2439
rect 911 -2445 914 -2439
rect 918 -2445 921 -2439
rect 925 -2445 928 -2439
rect 932 -2445 935 -2439
rect 939 -2445 942 -2439
rect 946 -2445 949 -2439
rect 953 -2445 956 -2439
rect 960 -2445 963 -2439
rect 967 -2445 973 -2439
rect 974 -2445 977 -2439
rect 981 -2445 984 -2439
rect 988 -2445 991 -2439
rect 995 -2445 998 -2439
rect 1002 -2445 1005 -2439
rect 1009 -2445 1012 -2439
rect 1016 -2445 1019 -2439
rect 1023 -2445 1026 -2439
rect 1030 -2445 1033 -2439
rect 1037 -2445 1040 -2439
rect 1044 -2445 1047 -2439
rect 1051 -2445 1054 -2439
rect 1058 -2445 1061 -2439
rect 1065 -2445 1068 -2439
rect 1072 -2445 1078 -2439
rect 1079 -2445 1082 -2439
rect 1086 -2445 1089 -2439
rect 1093 -2445 1096 -2439
rect 1100 -2445 1103 -2439
rect 1107 -2445 1110 -2439
rect 1114 -2445 1117 -2439
rect 1121 -2445 1124 -2439
rect 1128 -2445 1131 -2439
rect 1135 -2445 1138 -2439
rect 1142 -2445 1145 -2439
rect 1149 -2445 1152 -2439
rect 1156 -2445 1159 -2439
rect 1163 -2445 1166 -2439
rect 1170 -2445 1173 -2439
rect 1177 -2445 1180 -2439
rect 1184 -2445 1187 -2439
rect 1191 -2445 1197 -2439
rect 1198 -2445 1201 -2439
rect 1205 -2445 1211 -2439
rect 1212 -2445 1215 -2439
rect 1219 -2445 1222 -2439
rect 1226 -2445 1229 -2439
rect 1233 -2445 1236 -2439
rect 1240 -2445 1246 -2439
rect 1247 -2445 1250 -2439
rect 1254 -2445 1257 -2439
rect 1261 -2445 1264 -2439
rect 1268 -2445 1271 -2439
rect 1275 -2445 1278 -2439
rect 1282 -2445 1285 -2439
rect 1289 -2445 1292 -2439
rect 1296 -2445 1302 -2439
rect 1303 -2445 1306 -2439
rect 1310 -2445 1316 -2439
rect 1317 -2445 1320 -2439
rect 1324 -2445 1327 -2439
rect 1331 -2445 1334 -2439
rect 1338 -2445 1341 -2439
rect 1345 -2445 1348 -2439
rect 1352 -2445 1355 -2439
rect 1359 -2445 1362 -2439
rect 1366 -2445 1369 -2439
rect 1373 -2445 1376 -2439
rect 1380 -2445 1386 -2439
rect 1387 -2445 1390 -2439
rect 1394 -2445 1397 -2439
rect 1401 -2445 1404 -2439
rect 1408 -2445 1411 -2439
rect 1415 -2445 1418 -2439
rect 1422 -2445 1425 -2439
rect 1429 -2445 1432 -2439
rect 1436 -2445 1439 -2439
rect 1443 -2445 1446 -2439
rect 1450 -2445 1453 -2439
rect 1457 -2445 1460 -2439
rect 1464 -2445 1467 -2439
rect 1471 -2445 1474 -2439
rect 1478 -2445 1481 -2439
rect 1485 -2445 1488 -2439
rect 1492 -2445 1495 -2439
rect 1499 -2445 1502 -2439
rect 1506 -2445 1509 -2439
rect 1513 -2445 1516 -2439
rect 1520 -2445 1523 -2439
rect 1527 -2445 1530 -2439
rect 1534 -2445 1540 -2439
rect 1541 -2445 1544 -2439
rect 1548 -2445 1551 -2439
rect 1555 -2445 1558 -2439
rect 1562 -2445 1565 -2439
rect 1569 -2445 1572 -2439
rect 1576 -2445 1582 -2439
rect 1583 -2445 1586 -2439
rect 1590 -2445 1593 -2439
rect 1597 -2445 1600 -2439
rect 1604 -2445 1607 -2439
rect 1674 -2445 1677 -2439
rect 1 -2562 7 -2556
rect 8 -2562 14 -2556
rect 15 -2562 21 -2556
rect 22 -2562 28 -2556
rect 29 -2562 35 -2556
rect 36 -2562 42 -2556
rect 43 -2562 46 -2556
rect 50 -2562 53 -2556
rect 57 -2562 60 -2556
rect 64 -2562 70 -2556
rect 71 -2562 77 -2556
rect 78 -2562 81 -2556
rect 85 -2562 88 -2556
rect 92 -2562 95 -2556
rect 99 -2562 105 -2556
rect 106 -2562 109 -2556
rect 113 -2562 116 -2556
rect 120 -2562 123 -2556
rect 127 -2562 130 -2556
rect 134 -2562 137 -2556
rect 141 -2562 144 -2556
rect 148 -2562 154 -2556
rect 155 -2562 158 -2556
rect 162 -2562 168 -2556
rect 169 -2562 175 -2556
rect 176 -2562 179 -2556
rect 183 -2562 186 -2556
rect 190 -2562 193 -2556
rect 197 -2562 200 -2556
rect 204 -2562 207 -2556
rect 211 -2562 214 -2556
rect 218 -2562 221 -2556
rect 225 -2562 228 -2556
rect 232 -2562 235 -2556
rect 239 -2562 242 -2556
rect 246 -2562 249 -2556
rect 253 -2562 259 -2556
rect 260 -2562 263 -2556
rect 267 -2562 270 -2556
rect 274 -2562 277 -2556
rect 281 -2562 284 -2556
rect 288 -2562 291 -2556
rect 295 -2562 298 -2556
rect 302 -2562 305 -2556
rect 309 -2562 312 -2556
rect 316 -2562 319 -2556
rect 323 -2562 326 -2556
rect 330 -2562 333 -2556
rect 337 -2562 340 -2556
rect 344 -2562 347 -2556
rect 351 -2562 354 -2556
rect 358 -2562 361 -2556
rect 365 -2562 368 -2556
rect 372 -2562 375 -2556
rect 379 -2562 382 -2556
rect 386 -2562 389 -2556
rect 393 -2562 396 -2556
rect 400 -2562 403 -2556
rect 407 -2562 413 -2556
rect 414 -2562 417 -2556
rect 421 -2562 424 -2556
rect 428 -2562 434 -2556
rect 435 -2562 438 -2556
rect 442 -2562 448 -2556
rect 449 -2562 452 -2556
rect 456 -2562 459 -2556
rect 463 -2562 466 -2556
rect 470 -2562 473 -2556
rect 477 -2562 480 -2556
rect 484 -2562 487 -2556
rect 491 -2562 494 -2556
rect 498 -2562 501 -2556
rect 505 -2562 508 -2556
rect 512 -2562 515 -2556
rect 519 -2562 522 -2556
rect 526 -2562 529 -2556
rect 533 -2562 536 -2556
rect 540 -2562 543 -2556
rect 547 -2562 553 -2556
rect 554 -2562 557 -2556
rect 561 -2562 564 -2556
rect 568 -2562 571 -2556
rect 575 -2562 578 -2556
rect 582 -2562 585 -2556
rect 589 -2562 595 -2556
rect 596 -2562 599 -2556
rect 603 -2562 606 -2556
rect 610 -2562 613 -2556
rect 617 -2562 620 -2556
rect 624 -2562 630 -2556
rect 631 -2562 634 -2556
rect 638 -2562 641 -2556
rect 645 -2562 651 -2556
rect 652 -2562 655 -2556
rect 659 -2562 665 -2556
rect 666 -2562 669 -2556
rect 673 -2562 676 -2556
rect 680 -2562 683 -2556
rect 687 -2562 690 -2556
rect 694 -2562 697 -2556
rect 701 -2562 704 -2556
rect 708 -2562 711 -2556
rect 715 -2562 718 -2556
rect 722 -2562 725 -2556
rect 729 -2562 735 -2556
rect 736 -2562 742 -2556
rect 743 -2562 749 -2556
rect 750 -2562 756 -2556
rect 757 -2562 760 -2556
rect 764 -2562 767 -2556
rect 771 -2562 774 -2556
rect 778 -2562 781 -2556
rect 785 -2562 791 -2556
rect 792 -2562 795 -2556
rect 799 -2562 802 -2556
rect 806 -2562 809 -2556
rect 813 -2562 816 -2556
rect 820 -2562 826 -2556
rect 827 -2562 830 -2556
rect 834 -2562 837 -2556
rect 841 -2562 844 -2556
rect 848 -2562 851 -2556
rect 855 -2562 858 -2556
rect 862 -2562 865 -2556
rect 869 -2562 875 -2556
rect 876 -2562 879 -2556
rect 883 -2562 886 -2556
rect 890 -2562 893 -2556
rect 897 -2562 900 -2556
rect 904 -2562 907 -2556
rect 911 -2562 914 -2556
rect 918 -2562 921 -2556
rect 925 -2562 931 -2556
rect 932 -2562 935 -2556
rect 939 -2562 942 -2556
rect 946 -2562 949 -2556
rect 953 -2562 959 -2556
rect 960 -2562 963 -2556
rect 967 -2562 970 -2556
rect 974 -2562 977 -2556
rect 981 -2562 984 -2556
rect 988 -2562 991 -2556
rect 995 -2562 998 -2556
rect 1002 -2562 1005 -2556
rect 1009 -2562 1012 -2556
rect 1016 -2562 1019 -2556
rect 1023 -2562 1026 -2556
rect 1030 -2562 1033 -2556
rect 1037 -2562 1040 -2556
rect 1044 -2562 1047 -2556
rect 1051 -2562 1054 -2556
rect 1058 -2562 1064 -2556
rect 1065 -2562 1068 -2556
rect 1072 -2562 1075 -2556
rect 1079 -2562 1085 -2556
rect 1086 -2562 1092 -2556
rect 1093 -2562 1096 -2556
rect 1100 -2562 1103 -2556
rect 1107 -2562 1110 -2556
rect 1114 -2562 1117 -2556
rect 1121 -2562 1124 -2556
rect 1128 -2562 1131 -2556
rect 1135 -2562 1138 -2556
rect 1142 -2562 1145 -2556
rect 1149 -2562 1152 -2556
rect 1156 -2562 1159 -2556
rect 1163 -2562 1169 -2556
rect 1170 -2562 1173 -2556
rect 1177 -2562 1180 -2556
rect 1184 -2562 1190 -2556
rect 1191 -2562 1194 -2556
rect 1198 -2562 1201 -2556
rect 1205 -2562 1208 -2556
rect 1212 -2562 1215 -2556
rect 1219 -2562 1222 -2556
rect 1226 -2562 1229 -2556
rect 1233 -2562 1236 -2556
rect 1240 -2562 1243 -2556
rect 1247 -2562 1250 -2556
rect 1254 -2562 1257 -2556
rect 1261 -2562 1264 -2556
rect 1268 -2562 1271 -2556
rect 1275 -2562 1278 -2556
rect 1282 -2562 1285 -2556
rect 1289 -2562 1292 -2556
rect 1296 -2562 1299 -2556
rect 1303 -2562 1306 -2556
rect 1310 -2562 1313 -2556
rect 1317 -2562 1320 -2556
rect 1324 -2562 1327 -2556
rect 1331 -2562 1334 -2556
rect 1338 -2562 1341 -2556
rect 1345 -2562 1348 -2556
rect 1352 -2562 1355 -2556
rect 1359 -2562 1362 -2556
rect 1366 -2562 1369 -2556
rect 1373 -2562 1376 -2556
rect 1380 -2562 1383 -2556
rect 1387 -2562 1390 -2556
rect 1394 -2562 1397 -2556
rect 1401 -2562 1404 -2556
rect 1408 -2562 1411 -2556
rect 1415 -2562 1418 -2556
rect 1422 -2562 1425 -2556
rect 1429 -2562 1432 -2556
rect 1436 -2562 1439 -2556
rect 1443 -2562 1446 -2556
rect 1450 -2562 1453 -2556
rect 1457 -2562 1460 -2556
rect 1464 -2562 1467 -2556
rect 1471 -2562 1474 -2556
rect 1478 -2562 1481 -2556
rect 1485 -2562 1488 -2556
rect 1492 -2562 1495 -2556
rect 1499 -2562 1502 -2556
rect 1506 -2562 1509 -2556
rect 1513 -2562 1516 -2556
rect 1520 -2562 1523 -2556
rect 1527 -2562 1530 -2556
rect 1534 -2562 1537 -2556
rect 1541 -2562 1544 -2556
rect 1548 -2562 1551 -2556
rect 1555 -2562 1558 -2556
rect 1562 -2562 1565 -2556
rect 1569 -2562 1572 -2556
rect 1576 -2562 1579 -2556
rect 1583 -2562 1586 -2556
rect 1590 -2562 1593 -2556
rect 1597 -2562 1600 -2556
rect 1604 -2562 1607 -2556
rect 1611 -2562 1614 -2556
rect 1618 -2562 1621 -2556
rect 1625 -2562 1628 -2556
rect 1632 -2562 1635 -2556
rect 1639 -2562 1642 -2556
rect 1646 -2562 1649 -2556
rect 1653 -2562 1656 -2556
rect 1660 -2562 1663 -2556
rect 1667 -2562 1670 -2556
rect 1674 -2562 1680 -2556
rect 1681 -2562 1684 -2556
rect 1688 -2562 1691 -2556
rect 1695 -2562 1698 -2556
rect 1702 -2562 1708 -2556
rect 1709 -2562 1712 -2556
rect 1716 -2562 1719 -2556
rect 1723 -2562 1726 -2556
rect 1730 -2562 1733 -2556
rect 1737 -2562 1740 -2556
rect 1 -2691 7 -2685
rect 8 -2691 14 -2685
rect 15 -2691 21 -2685
rect 22 -2691 28 -2685
rect 29 -2691 35 -2685
rect 36 -2691 42 -2685
rect 43 -2691 46 -2685
rect 50 -2691 53 -2685
rect 57 -2691 60 -2685
rect 64 -2691 70 -2685
rect 71 -2691 74 -2685
rect 78 -2691 84 -2685
rect 85 -2691 91 -2685
rect 92 -2691 95 -2685
rect 99 -2691 102 -2685
rect 106 -2691 109 -2685
rect 113 -2691 119 -2685
rect 120 -2691 123 -2685
rect 127 -2691 130 -2685
rect 134 -2691 137 -2685
rect 141 -2691 144 -2685
rect 148 -2691 151 -2685
rect 155 -2691 158 -2685
rect 162 -2691 168 -2685
rect 169 -2691 172 -2685
rect 176 -2691 179 -2685
rect 183 -2691 186 -2685
rect 190 -2691 193 -2685
rect 197 -2691 203 -2685
rect 204 -2691 207 -2685
rect 211 -2691 214 -2685
rect 218 -2691 221 -2685
rect 225 -2691 228 -2685
rect 232 -2691 235 -2685
rect 239 -2691 242 -2685
rect 246 -2691 252 -2685
rect 253 -2691 256 -2685
rect 260 -2691 263 -2685
rect 267 -2691 270 -2685
rect 274 -2691 277 -2685
rect 281 -2691 284 -2685
rect 288 -2691 291 -2685
rect 295 -2691 298 -2685
rect 302 -2691 305 -2685
rect 309 -2691 312 -2685
rect 316 -2691 319 -2685
rect 323 -2691 326 -2685
rect 330 -2691 333 -2685
rect 337 -2691 340 -2685
rect 344 -2691 347 -2685
rect 351 -2691 354 -2685
rect 358 -2691 361 -2685
rect 365 -2691 368 -2685
rect 372 -2691 375 -2685
rect 379 -2691 382 -2685
rect 386 -2691 389 -2685
rect 393 -2691 396 -2685
rect 400 -2691 403 -2685
rect 407 -2691 413 -2685
rect 414 -2691 420 -2685
rect 421 -2691 424 -2685
rect 428 -2691 431 -2685
rect 435 -2691 438 -2685
rect 442 -2691 445 -2685
rect 449 -2691 455 -2685
rect 456 -2691 462 -2685
rect 463 -2691 469 -2685
rect 470 -2691 473 -2685
rect 477 -2691 483 -2685
rect 484 -2691 487 -2685
rect 491 -2691 494 -2685
rect 498 -2691 501 -2685
rect 505 -2691 508 -2685
rect 512 -2691 515 -2685
rect 519 -2691 522 -2685
rect 526 -2691 529 -2685
rect 533 -2691 536 -2685
rect 540 -2691 543 -2685
rect 547 -2691 550 -2685
rect 554 -2691 557 -2685
rect 561 -2691 564 -2685
rect 568 -2691 571 -2685
rect 575 -2691 581 -2685
rect 582 -2691 585 -2685
rect 589 -2691 592 -2685
rect 596 -2691 602 -2685
rect 603 -2691 606 -2685
rect 610 -2691 613 -2685
rect 617 -2691 620 -2685
rect 624 -2691 630 -2685
rect 631 -2691 634 -2685
rect 638 -2691 641 -2685
rect 645 -2691 648 -2685
rect 652 -2691 655 -2685
rect 659 -2691 662 -2685
rect 666 -2691 672 -2685
rect 673 -2691 679 -2685
rect 680 -2691 683 -2685
rect 687 -2691 693 -2685
rect 694 -2691 697 -2685
rect 701 -2691 704 -2685
rect 708 -2691 711 -2685
rect 715 -2691 718 -2685
rect 722 -2691 725 -2685
rect 729 -2691 735 -2685
rect 736 -2691 739 -2685
rect 743 -2691 746 -2685
rect 750 -2691 756 -2685
rect 757 -2691 760 -2685
rect 764 -2691 770 -2685
rect 771 -2691 774 -2685
rect 778 -2691 781 -2685
rect 785 -2691 788 -2685
rect 792 -2691 795 -2685
rect 799 -2691 805 -2685
rect 806 -2691 809 -2685
rect 813 -2691 816 -2685
rect 820 -2691 823 -2685
rect 827 -2691 830 -2685
rect 834 -2691 840 -2685
rect 841 -2691 847 -2685
rect 848 -2691 851 -2685
rect 855 -2691 858 -2685
rect 862 -2691 865 -2685
rect 869 -2691 875 -2685
rect 876 -2691 879 -2685
rect 883 -2691 886 -2685
rect 890 -2691 896 -2685
rect 897 -2691 900 -2685
rect 904 -2691 907 -2685
rect 911 -2691 914 -2685
rect 918 -2691 921 -2685
rect 925 -2691 928 -2685
rect 932 -2691 935 -2685
rect 939 -2691 942 -2685
rect 946 -2691 949 -2685
rect 953 -2691 959 -2685
rect 960 -2691 963 -2685
rect 967 -2691 970 -2685
rect 974 -2691 977 -2685
rect 981 -2691 984 -2685
rect 988 -2691 994 -2685
rect 995 -2691 998 -2685
rect 1002 -2691 1005 -2685
rect 1009 -2691 1012 -2685
rect 1016 -2691 1019 -2685
rect 1023 -2691 1026 -2685
rect 1030 -2691 1036 -2685
rect 1037 -2691 1040 -2685
rect 1044 -2691 1047 -2685
rect 1051 -2691 1054 -2685
rect 1058 -2691 1061 -2685
rect 1065 -2691 1068 -2685
rect 1072 -2691 1075 -2685
rect 1079 -2691 1082 -2685
rect 1086 -2691 1089 -2685
rect 1093 -2691 1099 -2685
rect 1100 -2691 1103 -2685
rect 1107 -2691 1110 -2685
rect 1114 -2691 1117 -2685
rect 1121 -2691 1124 -2685
rect 1128 -2691 1131 -2685
rect 1135 -2691 1138 -2685
rect 1142 -2691 1145 -2685
rect 1149 -2691 1152 -2685
rect 1156 -2691 1159 -2685
rect 1163 -2691 1166 -2685
rect 1170 -2691 1173 -2685
rect 1177 -2691 1180 -2685
rect 1184 -2691 1187 -2685
rect 1191 -2691 1194 -2685
rect 1198 -2691 1201 -2685
rect 1205 -2691 1208 -2685
rect 1212 -2691 1215 -2685
rect 1219 -2691 1222 -2685
rect 1226 -2691 1229 -2685
rect 1233 -2691 1236 -2685
rect 1240 -2691 1243 -2685
rect 1247 -2691 1250 -2685
rect 1254 -2691 1257 -2685
rect 1261 -2691 1264 -2685
rect 1268 -2691 1271 -2685
rect 1275 -2691 1278 -2685
rect 1282 -2691 1285 -2685
rect 1289 -2691 1292 -2685
rect 1296 -2691 1299 -2685
rect 1303 -2691 1306 -2685
rect 1310 -2691 1313 -2685
rect 1317 -2691 1320 -2685
rect 1324 -2691 1327 -2685
rect 1331 -2691 1334 -2685
rect 1338 -2691 1341 -2685
rect 1345 -2691 1348 -2685
rect 1352 -2691 1355 -2685
rect 1359 -2691 1362 -2685
rect 1366 -2691 1369 -2685
rect 1373 -2691 1376 -2685
rect 1380 -2691 1383 -2685
rect 1387 -2691 1390 -2685
rect 1394 -2691 1397 -2685
rect 1401 -2691 1404 -2685
rect 1408 -2691 1411 -2685
rect 1415 -2691 1418 -2685
rect 1422 -2691 1425 -2685
rect 1429 -2691 1432 -2685
rect 1436 -2691 1439 -2685
rect 1443 -2691 1446 -2685
rect 1450 -2691 1453 -2685
rect 1457 -2691 1460 -2685
rect 1464 -2691 1467 -2685
rect 1471 -2691 1474 -2685
rect 1478 -2691 1481 -2685
rect 1485 -2691 1488 -2685
rect 1492 -2691 1495 -2685
rect 1499 -2691 1502 -2685
rect 1506 -2691 1509 -2685
rect 1513 -2691 1516 -2685
rect 1520 -2691 1523 -2685
rect 1527 -2691 1530 -2685
rect 1534 -2691 1537 -2685
rect 1541 -2691 1544 -2685
rect 1548 -2691 1551 -2685
rect 1555 -2691 1558 -2685
rect 1562 -2691 1565 -2685
rect 1569 -2691 1572 -2685
rect 1576 -2691 1579 -2685
rect 1583 -2691 1586 -2685
rect 1590 -2691 1593 -2685
rect 1597 -2691 1600 -2685
rect 1604 -2691 1607 -2685
rect 1611 -2691 1614 -2685
rect 1618 -2691 1621 -2685
rect 1625 -2691 1628 -2685
rect 1632 -2691 1635 -2685
rect 1639 -2691 1642 -2685
rect 1646 -2691 1649 -2685
rect 1653 -2691 1656 -2685
rect 1660 -2691 1663 -2685
rect 1667 -2691 1670 -2685
rect 1674 -2691 1677 -2685
rect 1681 -2691 1684 -2685
rect 1688 -2691 1691 -2685
rect 1695 -2691 1698 -2685
rect 1702 -2691 1705 -2685
rect 1 -2840 7 -2834
rect 8 -2840 14 -2834
rect 15 -2840 21 -2834
rect 22 -2840 28 -2834
rect 29 -2840 35 -2834
rect 36 -2840 39 -2834
rect 43 -2840 46 -2834
rect 50 -2840 53 -2834
rect 57 -2840 60 -2834
rect 64 -2840 67 -2834
rect 71 -2840 74 -2834
rect 78 -2840 81 -2834
rect 85 -2840 91 -2834
rect 92 -2840 98 -2834
rect 99 -2840 102 -2834
rect 106 -2840 112 -2834
rect 113 -2840 116 -2834
rect 120 -2840 123 -2834
rect 127 -2840 133 -2834
rect 134 -2840 137 -2834
rect 141 -2840 144 -2834
rect 148 -2840 151 -2834
rect 155 -2840 158 -2834
rect 162 -2840 168 -2834
rect 169 -2840 172 -2834
rect 176 -2840 182 -2834
rect 183 -2840 186 -2834
rect 190 -2840 193 -2834
rect 197 -2840 200 -2834
rect 204 -2840 207 -2834
rect 211 -2840 214 -2834
rect 218 -2840 221 -2834
rect 225 -2840 231 -2834
rect 232 -2840 235 -2834
rect 239 -2840 242 -2834
rect 246 -2840 252 -2834
rect 253 -2840 256 -2834
rect 260 -2840 263 -2834
rect 267 -2840 270 -2834
rect 274 -2840 277 -2834
rect 281 -2840 284 -2834
rect 288 -2840 291 -2834
rect 295 -2840 298 -2834
rect 302 -2840 305 -2834
rect 309 -2840 312 -2834
rect 316 -2840 319 -2834
rect 323 -2840 326 -2834
rect 330 -2840 333 -2834
rect 337 -2840 340 -2834
rect 344 -2840 347 -2834
rect 351 -2840 354 -2834
rect 358 -2840 361 -2834
rect 365 -2840 368 -2834
rect 372 -2840 375 -2834
rect 379 -2840 385 -2834
rect 386 -2840 389 -2834
rect 393 -2840 396 -2834
rect 400 -2840 403 -2834
rect 407 -2840 410 -2834
rect 414 -2840 417 -2834
rect 421 -2840 424 -2834
rect 428 -2840 431 -2834
rect 435 -2840 438 -2834
rect 442 -2840 445 -2834
rect 449 -2840 455 -2834
rect 456 -2840 459 -2834
rect 463 -2840 466 -2834
rect 470 -2840 473 -2834
rect 477 -2840 480 -2834
rect 484 -2840 487 -2834
rect 491 -2840 494 -2834
rect 498 -2840 501 -2834
rect 505 -2840 508 -2834
rect 512 -2840 515 -2834
rect 519 -2840 525 -2834
rect 526 -2840 529 -2834
rect 533 -2840 536 -2834
rect 540 -2840 543 -2834
rect 547 -2840 550 -2834
rect 554 -2840 557 -2834
rect 561 -2840 564 -2834
rect 568 -2840 571 -2834
rect 575 -2840 578 -2834
rect 582 -2840 585 -2834
rect 589 -2840 595 -2834
rect 596 -2840 599 -2834
rect 603 -2840 606 -2834
rect 610 -2840 613 -2834
rect 617 -2840 620 -2834
rect 624 -2840 627 -2834
rect 631 -2840 634 -2834
rect 638 -2840 641 -2834
rect 645 -2840 651 -2834
rect 652 -2840 658 -2834
rect 659 -2840 662 -2834
rect 666 -2840 669 -2834
rect 673 -2840 676 -2834
rect 680 -2840 686 -2834
rect 687 -2840 690 -2834
rect 694 -2840 697 -2834
rect 701 -2840 704 -2834
rect 708 -2840 711 -2834
rect 715 -2840 718 -2834
rect 722 -2840 725 -2834
rect 729 -2840 732 -2834
rect 736 -2840 739 -2834
rect 743 -2840 746 -2834
rect 750 -2840 753 -2834
rect 757 -2840 763 -2834
rect 764 -2840 770 -2834
rect 771 -2840 777 -2834
rect 778 -2840 781 -2834
rect 785 -2840 788 -2834
rect 792 -2840 795 -2834
rect 799 -2840 805 -2834
rect 806 -2840 809 -2834
rect 813 -2840 816 -2834
rect 820 -2840 823 -2834
rect 827 -2840 830 -2834
rect 834 -2840 837 -2834
rect 841 -2840 844 -2834
rect 848 -2840 851 -2834
rect 855 -2840 858 -2834
rect 862 -2840 865 -2834
rect 869 -2840 872 -2834
rect 876 -2840 879 -2834
rect 883 -2840 889 -2834
rect 890 -2840 896 -2834
rect 897 -2840 903 -2834
rect 904 -2840 907 -2834
rect 911 -2840 914 -2834
rect 918 -2840 921 -2834
rect 925 -2840 928 -2834
rect 932 -2840 935 -2834
rect 939 -2840 942 -2834
rect 946 -2840 949 -2834
rect 953 -2840 956 -2834
rect 960 -2840 963 -2834
rect 967 -2840 970 -2834
rect 974 -2840 977 -2834
rect 981 -2840 987 -2834
rect 988 -2840 991 -2834
rect 995 -2840 1001 -2834
rect 1002 -2840 1005 -2834
rect 1009 -2840 1012 -2834
rect 1016 -2840 1019 -2834
rect 1023 -2840 1026 -2834
rect 1030 -2840 1033 -2834
rect 1037 -2840 1040 -2834
rect 1044 -2840 1050 -2834
rect 1051 -2840 1054 -2834
rect 1058 -2840 1061 -2834
rect 1065 -2840 1068 -2834
rect 1072 -2840 1075 -2834
rect 1079 -2840 1082 -2834
rect 1086 -2840 1089 -2834
rect 1093 -2840 1099 -2834
rect 1100 -2840 1103 -2834
rect 1107 -2840 1110 -2834
rect 1114 -2840 1120 -2834
rect 1121 -2840 1124 -2834
rect 1128 -2840 1131 -2834
rect 1135 -2840 1138 -2834
rect 1142 -2840 1145 -2834
rect 1149 -2840 1152 -2834
rect 1156 -2840 1159 -2834
rect 1163 -2840 1166 -2834
rect 1170 -2840 1173 -2834
rect 1177 -2840 1180 -2834
rect 1184 -2840 1190 -2834
rect 1191 -2840 1194 -2834
rect 1198 -2840 1201 -2834
rect 1205 -2840 1208 -2834
rect 1212 -2840 1215 -2834
rect 1219 -2840 1222 -2834
rect 1226 -2840 1229 -2834
rect 1233 -2840 1236 -2834
rect 1240 -2840 1243 -2834
rect 1247 -2840 1250 -2834
rect 1254 -2840 1257 -2834
rect 1261 -2840 1264 -2834
rect 1268 -2840 1271 -2834
rect 1275 -2840 1281 -2834
rect 1282 -2840 1285 -2834
rect 1289 -2840 1292 -2834
rect 1296 -2840 1299 -2834
rect 1303 -2840 1306 -2834
rect 1310 -2840 1313 -2834
rect 1317 -2840 1320 -2834
rect 1324 -2840 1327 -2834
rect 1331 -2840 1334 -2834
rect 1338 -2840 1341 -2834
rect 1345 -2840 1348 -2834
rect 1352 -2840 1355 -2834
rect 1359 -2840 1362 -2834
rect 1366 -2840 1369 -2834
rect 1373 -2840 1376 -2834
rect 1380 -2840 1383 -2834
rect 1387 -2840 1390 -2834
rect 1394 -2840 1397 -2834
rect 1401 -2840 1404 -2834
rect 1408 -2840 1411 -2834
rect 1415 -2840 1418 -2834
rect 1422 -2840 1425 -2834
rect 1429 -2840 1432 -2834
rect 1436 -2840 1439 -2834
rect 1443 -2840 1446 -2834
rect 1450 -2840 1453 -2834
rect 1457 -2840 1460 -2834
rect 1464 -2840 1467 -2834
rect 1471 -2840 1474 -2834
rect 1478 -2840 1481 -2834
rect 1485 -2840 1488 -2834
rect 1492 -2840 1495 -2834
rect 1499 -2840 1502 -2834
rect 1506 -2840 1512 -2834
rect 1513 -2840 1519 -2834
rect 1520 -2840 1523 -2834
rect 1527 -2840 1530 -2834
rect 1534 -2840 1537 -2834
rect 1541 -2840 1544 -2834
rect 1548 -2840 1551 -2834
rect 1555 -2840 1558 -2834
rect 1 -2951 7 -2945
rect 8 -2951 14 -2945
rect 15 -2951 21 -2945
rect 22 -2951 28 -2945
rect 29 -2951 32 -2945
rect 36 -2951 39 -2945
rect 43 -2951 46 -2945
rect 50 -2951 53 -2945
rect 57 -2951 60 -2945
rect 64 -2951 67 -2945
rect 71 -2951 77 -2945
rect 78 -2951 81 -2945
rect 85 -2951 88 -2945
rect 92 -2951 95 -2945
rect 99 -2951 102 -2945
rect 106 -2951 109 -2945
rect 113 -2951 119 -2945
rect 120 -2951 123 -2945
rect 127 -2951 130 -2945
rect 134 -2951 137 -2945
rect 141 -2951 144 -2945
rect 148 -2951 151 -2945
rect 155 -2951 161 -2945
rect 162 -2951 165 -2945
rect 169 -2951 172 -2945
rect 176 -2951 182 -2945
rect 183 -2951 186 -2945
rect 190 -2951 193 -2945
rect 197 -2951 200 -2945
rect 204 -2951 207 -2945
rect 211 -2951 214 -2945
rect 218 -2951 221 -2945
rect 225 -2951 228 -2945
rect 232 -2951 235 -2945
rect 239 -2951 242 -2945
rect 246 -2951 252 -2945
rect 253 -2951 259 -2945
rect 260 -2951 266 -2945
rect 267 -2951 270 -2945
rect 274 -2951 277 -2945
rect 281 -2951 284 -2945
rect 288 -2951 291 -2945
rect 295 -2951 298 -2945
rect 302 -2951 305 -2945
rect 309 -2951 312 -2945
rect 316 -2951 319 -2945
rect 323 -2951 326 -2945
rect 330 -2951 333 -2945
rect 337 -2951 340 -2945
rect 344 -2951 347 -2945
rect 351 -2951 354 -2945
rect 358 -2951 361 -2945
rect 365 -2951 368 -2945
rect 372 -2951 378 -2945
rect 379 -2951 382 -2945
rect 386 -2951 389 -2945
rect 393 -2951 396 -2945
rect 400 -2951 406 -2945
rect 407 -2951 413 -2945
rect 414 -2951 417 -2945
rect 421 -2951 424 -2945
rect 428 -2951 431 -2945
rect 435 -2951 438 -2945
rect 442 -2951 445 -2945
rect 449 -2951 452 -2945
rect 456 -2951 459 -2945
rect 463 -2951 466 -2945
rect 470 -2951 476 -2945
rect 477 -2951 483 -2945
rect 484 -2951 487 -2945
rect 491 -2951 494 -2945
rect 498 -2951 504 -2945
rect 505 -2951 508 -2945
rect 512 -2951 515 -2945
rect 519 -2951 522 -2945
rect 526 -2951 529 -2945
rect 533 -2951 536 -2945
rect 540 -2951 543 -2945
rect 547 -2951 550 -2945
rect 554 -2951 557 -2945
rect 561 -2951 567 -2945
rect 568 -2951 571 -2945
rect 575 -2951 578 -2945
rect 582 -2951 585 -2945
rect 589 -2951 592 -2945
rect 596 -2951 599 -2945
rect 603 -2951 609 -2945
rect 610 -2951 613 -2945
rect 617 -2951 620 -2945
rect 624 -2951 627 -2945
rect 631 -2951 637 -2945
rect 638 -2951 641 -2945
rect 645 -2951 648 -2945
rect 652 -2951 655 -2945
rect 659 -2951 662 -2945
rect 666 -2951 672 -2945
rect 673 -2951 676 -2945
rect 680 -2951 683 -2945
rect 687 -2951 693 -2945
rect 694 -2951 697 -2945
rect 701 -2951 707 -2945
rect 708 -2951 711 -2945
rect 715 -2951 718 -2945
rect 722 -2951 725 -2945
rect 729 -2951 735 -2945
rect 736 -2951 739 -2945
rect 743 -2951 746 -2945
rect 750 -2951 753 -2945
rect 757 -2951 763 -2945
rect 764 -2951 767 -2945
rect 771 -2951 774 -2945
rect 778 -2951 781 -2945
rect 785 -2951 788 -2945
rect 792 -2951 795 -2945
rect 799 -2951 802 -2945
rect 806 -2951 809 -2945
rect 813 -2951 816 -2945
rect 820 -2951 823 -2945
rect 827 -2951 830 -2945
rect 834 -2951 837 -2945
rect 841 -2951 844 -2945
rect 848 -2951 851 -2945
rect 855 -2951 858 -2945
rect 862 -2951 868 -2945
rect 869 -2951 872 -2945
rect 876 -2951 879 -2945
rect 883 -2951 886 -2945
rect 890 -2951 893 -2945
rect 897 -2951 900 -2945
rect 904 -2951 907 -2945
rect 911 -2951 917 -2945
rect 918 -2951 921 -2945
rect 925 -2951 931 -2945
rect 932 -2951 938 -2945
rect 939 -2951 942 -2945
rect 946 -2951 949 -2945
rect 953 -2951 956 -2945
rect 960 -2951 963 -2945
rect 967 -2951 970 -2945
rect 974 -2951 977 -2945
rect 981 -2951 984 -2945
rect 988 -2951 991 -2945
rect 995 -2951 1001 -2945
rect 1002 -2951 1005 -2945
rect 1009 -2951 1012 -2945
rect 1016 -2951 1022 -2945
rect 1023 -2951 1029 -2945
rect 1030 -2951 1033 -2945
rect 1037 -2951 1040 -2945
rect 1044 -2951 1047 -2945
rect 1051 -2951 1054 -2945
rect 1058 -2951 1061 -2945
rect 1065 -2951 1068 -2945
rect 1072 -2951 1075 -2945
rect 1079 -2951 1082 -2945
rect 1086 -2951 1089 -2945
rect 1093 -2951 1096 -2945
rect 1100 -2951 1103 -2945
rect 1107 -2951 1110 -2945
rect 1114 -2951 1117 -2945
rect 1121 -2951 1124 -2945
rect 1128 -2951 1131 -2945
rect 1135 -2951 1138 -2945
rect 1142 -2951 1145 -2945
rect 1149 -2951 1152 -2945
rect 1156 -2951 1159 -2945
rect 1163 -2951 1166 -2945
rect 1170 -2951 1173 -2945
rect 1177 -2951 1180 -2945
rect 1184 -2951 1187 -2945
rect 1191 -2951 1194 -2945
rect 1198 -2951 1204 -2945
rect 1205 -2951 1208 -2945
rect 1212 -2951 1215 -2945
rect 1219 -2951 1222 -2945
rect 1226 -2951 1229 -2945
rect 1233 -2951 1236 -2945
rect 1240 -2951 1243 -2945
rect 1247 -2951 1250 -2945
rect 1254 -2951 1257 -2945
rect 1261 -2951 1264 -2945
rect 1268 -2951 1271 -2945
rect 1275 -2951 1278 -2945
rect 1282 -2951 1285 -2945
rect 1289 -2951 1292 -2945
rect 1296 -2951 1299 -2945
rect 1303 -2951 1306 -2945
rect 1310 -2951 1313 -2945
rect 1317 -2951 1320 -2945
rect 1324 -2951 1327 -2945
rect 1331 -2951 1334 -2945
rect 1338 -2951 1341 -2945
rect 1345 -2951 1348 -2945
rect 1352 -2951 1355 -2945
rect 1359 -2951 1362 -2945
rect 1366 -2951 1369 -2945
rect 1373 -2951 1376 -2945
rect 1380 -2951 1383 -2945
rect 1387 -2951 1390 -2945
rect 1394 -2951 1397 -2945
rect 1401 -2951 1404 -2945
rect 1408 -2951 1411 -2945
rect 1415 -2951 1418 -2945
rect 1422 -2951 1425 -2945
rect 1429 -2951 1432 -2945
rect 1436 -2951 1439 -2945
rect 1443 -2951 1449 -2945
rect 1450 -2951 1453 -2945
rect 1457 -2951 1460 -2945
rect 1464 -2951 1467 -2945
rect 1478 -2951 1481 -2945
rect 1485 -2951 1488 -2945
rect 1492 -2951 1495 -2945
rect 1499 -2951 1502 -2945
rect 1 -3070 7 -3064
rect 8 -3070 14 -3064
rect 15 -3070 21 -3064
rect 36 -3070 39 -3064
rect 43 -3070 46 -3064
rect 50 -3070 53 -3064
rect 57 -3070 60 -3064
rect 64 -3070 67 -3064
rect 71 -3070 74 -3064
rect 78 -3070 81 -3064
rect 85 -3070 88 -3064
rect 92 -3070 98 -3064
rect 99 -3070 102 -3064
rect 106 -3070 109 -3064
rect 113 -3070 116 -3064
rect 120 -3070 126 -3064
rect 127 -3070 130 -3064
rect 134 -3070 137 -3064
rect 141 -3070 144 -3064
rect 148 -3070 151 -3064
rect 155 -3070 158 -3064
rect 162 -3070 165 -3064
rect 169 -3070 172 -3064
rect 176 -3070 182 -3064
rect 183 -3070 186 -3064
rect 190 -3070 193 -3064
rect 197 -3070 203 -3064
rect 204 -3070 207 -3064
rect 211 -3070 214 -3064
rect 218 -3070 224 -3064
rect 225 -3070 228 -3064
rect 232 -3070 235 -3064
rect 239 -3070 245 -3064
rect 246 -3070 252 -3064
rect 253 -3070 256 -3064
rect 260 -3070 266 -3064
rect 267 -3070 270 -3064
rect 274 -3070 277 -3064
rect 281 -3070 284 -3064
rect 288 -3070 291 -3064
rect 295 -3070 301 -3064
rect 302 -3070 305 -3064
rect 309 -3070 312 -3064
rect 316 -3070 319 -3064
rect 323 -3070 326 -3064
rect 330 -3070 333 -3064
rect 337 -3070 340 -3064
rect 344 -3070 347 -3064
rect 351 -3070 357 -3064
rect 358 -3070 361 -3064
rect 365 -3070 368 -3064
rect 372 -3070 375 -3064
rect 379 -3070 382 -3064
rect 386 -3070 389 -3064
rect 393 -3070 396 -3064
rect 400 -3070 403 -3064
rect 407 -3070 413 -3064
rect 414 -3070 417 -3064
rect 421 -3070 424 -3064
rect 428 -3070 431 -3064
rect 435 -3070 438 -3064
rect 442 -3070 445 -3064
rect 449 -3070 452 -3064
rect 456 -3070 459 -3064
rect 463 -3070 466 -3064
rect 470 -3070 473 -3064
rect 477 -3070 480 -3064
rect 484 -3070 487 -3064
rect 491 -3070 494 -3064
rect 498 -3070 501 -3064
rect 505 -3070 508 -3064
rect 512 -3070 515 -3064
rect 519 -3070 525 -3064
rect 526 -3070 529 -3064
rect 533 -3070 536 -3064
rect 540 -3070 543 -3064
rect 547 -3070 550 -3064
rect 554 -3070 557 -3064
rect 561 -3070 564 -3064
rect 568 -3070 571 -3064
rect 575 -3070 578 -3064
rect 582 -3070 585 -3064
rect 589 -3070 592 -3064
rect 596 -3070 599 -3064
rect 603 -3070 609 -3064
rect 610 -3070 613 -3064
rect 617 -3070 623 -3064
rect 624 -3070 627 -3064
rect 631 -3070 634 -3064
rect 638 -3070 644 -3064
rect 645 -3070 648 -3064
rect 652 -3070 655 -3064
rect 659 -3070 662 -3064
rect 666 -3070 669 -3064
rect 673 -3070 676 -3064
rect 680 -3070 686 -3064
rect 687 -3070 690 -3064
rect 694 -3070 697 -3064
rect 701 -3070 707 -3064
rect 708 -3070 711 -3064
rect 715 -3070 718 -3064
rect 722 -3070 725 -3064
rect 729 -3070 732 -3064
rect 736 -3070 742 -3064
rect 743 -3070 746 -3064
rect 750 -3070 753 -3064
rect 757 -3070 760 -3064
rect 764 -3070 767 -3064
rect 771 -3070 774 -3064
rect 778 -3070 781 -3064
rect 785 -3070 788 -3064
rect 792 -3070 798 -3064
rect 799 -3070 802 -3064
rect 806 -3070 809 -3064
rect 813 -3070 816 -3064
rect 820 -3070 823 -3064
rect 827 -3070 830 -3064
rect 834 -3070 837 -3064
rect 841 -3070 844 -3064
rect 848 -3070 854 -3064
rect 855 -3070 858 -3064
rect 862 -3070 865 -3064
rect 869 -3070 875 -3064
rect 876 -3070 879 -3064
rect 883 -3070 886 -3064
rect 890 -3070 893 -3064
rect 897 -3070 900 -3064
rect 904 -3070 907 -3064
rect 911 -3070 914 -3064
rect 918 -3070 924 -3064
rect 925 -3070 931 -3064
rect 932 -3070 935 -3064
rect 939 -3070 942 -3064
rect 946 -3070 949 -3064
rect 953 -3070 956 -3064
rect 960 -3070 966 -3064
rect 967 -3070 970 -3064
rect 974 -3070 977 -3064
rect 981 -3070 984 -3064
rect 988 -3070 991 -3064
rect 995 -3070 1001 -3064
rect 1002 -3070 1005 -3064
rect 1009 -3070 1012 -3064
rect 1016 -3070 1019 -3064
rect 1023 -3070 1026 -3064
rect 1030 -3070 1033 -3064
rect 1037 -3070 1040 -3064
rect 1044 -3070 1047 -3064
rect 1051 -3070 1054 -3064
rect 1058 -3070 1064 -3064
rect 1065 -3070 1068 -3064
rect 1072 -3070 1075 -3064
rect 1079 -3070 1082 -3064
rect 1086 -3070 1092 -3064
rect 1093 -3070 1096 -3064
rect 1100 -3070 1103 -3064
rect 1107 -3070 1110 -3064
rect 1114 -3070 1117 -3064
rect 1121 -3070 1124 -3064
rect 1128 -3070 1131 -3064
rect 1135 -3070 1138 -3064
rect 1142 -3070 1145 -3064
rect 1149 -3070 1152 -3064
rect 1156 -3070 1159 -3064
rect 1163 -3070 1166 -3064
rect 1170 -3070 1173 -3064
rect 1177 -3070 1180 -3064
rect 1184 -3070 1187 -3064
rect 1191 -3070 1194 -3064
rect 1198 -3070 1201 -3064
rect 1205 -3070 1208 -3064
rect 1212 -3070 1215 -3064
rect 1219 -3070 1225 -3064
rect 1226 -3070 1229 -3064
rect 1233 -3070 1236 -3064
rect 1240 -3070 1243 -3064
rect 1247 -3070 1250 -3064
rect 1254 -3070 1257 -3064
rect 1261 -3070 1264 -3064
rect 1268 -3070 1271 -3064
rect 1275 -3070 1278 -3064
rect 1282 -3070 1288 -3064
rect 1289 -3070 1292 -3064
rect 1296 -3070 1299 -3064
rect 1303 -3070 1306 -3064
rect 1310 -3070 1313 -3064
rect 1317 -3070 1320 -3064
rect 1324 -3070 1327 -3064
rect 1331 -3070 1334 -3064
rect 1338 -3070 1341 -3064
rect 1345 -3070 1348 -3064
rect 1373 -3070 1376 -3064
rect 1380 -3070 1383 -3064
rect 1415 -3070 1418 -3064
rect 1457 -3070 1460 -3064
rect 1464 -3070 1467 -3064
rect 1471 -3070 1474 -3064
rect 1 -3159 7 -3153
rect 8 -3159 14 -3153
rect 78 -3159 81 -3153
rect 85 -3159 88 -3153
rect 92 -3159 95 -3153
rect 99 -3159 102 -3153
rect 106 -3159 109 -3153
rect 113 -3159 116 -3153
rect 120 -3159 123 -3153
rect 127 -3159 130 -3153
rect 134 -3159 137 -3153
rect 141 -3159 144 -3153
rect 148 -3159 151 -3153
rect 155 -3159 158 -3153
rect 162 -3159 165 -3153
rect 169 -3159 172 -3153
rect 176 -3159 179 -3153
rect 183 -3159 189 -3153
rect 190 -3159 193 -3153
rect 197 -3159 200 -3153
rect 204 -3159 207 -3153
rect 211 -3159 217 -3153
rect 218 -3159 224 -3153
rect 225 -3159 228 -3153
rect 232 -3159 235 -3153
rect 239 -3159 242 -3153
rect 246 -3159 249 -3153
rect 253 -3159 256 -3153
rect 260 -3159 263 -3153
rect 267 -3159 270 -3153
rect 274 -3159 277 -3153
rect 281 -3159 284 -3153
rect 288 -3159 291 -3153
rect 295 -3159 298 -3153
rect 302 -3159 308 -3153
rect 309 -3159 312 -3153
rect 316 -3159 319 -3153
rect 323 -3159 326 -3153
rect 330 -3159 333 -3153
rect 337 -3159 340 -3153
rect 344 -3159 347 -3153
rect 351 -3159 354 -3153
rect 358 -3159 364 -3153
rect 365 -3159 368 -3153
rect 372 -3159 375 -3153
rect 379 -3159 382 -3153
rect 386 -3159 389 -3153
rect 393 -3159 396 -3153
rect 400 -3159 403 -3153
rect 407 -3159 410 -3153
rect 414 -3159 417 -3153
rect 421 -3159 424 -3153
rect 428 -3159 434 -3153
rect 435 -3159 438 -3153
rect 442 -3159 445 -3153
rect 449 -3159 452 -3153
rect 456 -3159 459 -3153
rect 463 -3159 466 -3153
rect 470 -3159 473 -3153
rect 477 -3159 480 -3153
rect 484 -3159 487 -3153
rect 491 -3159 494 -3153
rect 498 -3159 501 -3153
rect 505 -3159 508 -3153
rect 512 -3159 515 -3153
rect 519 -3159 522 -3153
rect 526 -3159 529 -3153
rect 533 -3159 536 -3153
rect 540 -3159 543 -3153
rect 547 -3159 550 -3153
rect 554 -3159 557 -3153
rect 561 -3159 564 -3153
rect 568 -3159 571 -3153
rect 575 -3159 581 -3153
rect 582 -3159 585 -3153
rect 589 -3159 592 -3153
rect 596 -3159 599 -3153
rect 603 -3159 609 -3153
rect 610 -3159 613 -3153
rect 617 -3159 623 -3153
rect 624 -3159 627 -3153
rect 631 -3159 637 -3153
rect 638 -3159 641 -3153
rect 645 -3159 648 -3153
rect 652 -3159 658 -3153
rect 659 -3159 665 -3153
rect 666 -3159 669 -3153
rect 673 -3159 676 -3153
rect 680 -3159 683 -3153
rect 687 -3159 693 -3153
rect 694 -3159 697 -3153
rect 701 -3159 707 -3153
rect 708 -3159 711 -3153
rect 715 -3159 718 -3153
rect 722 -3159 725 -3153
rect 729 -3159 735 -3153
rect 736 -3159 739 -3153
rect 743 -3159 746 -3153
rect 750 -3159 753 -3153
rect 757 -3159 760 -3153
rect 764 -3159 767 -3153
rect 771 -3159 777 -3153
rect 778 -3159 784 -3153
rect 785 -3159 788 -3153
rect 792 -3159 795 -3153
rect 799 -3159 802 -3153
rect 806 -3159 809 -3153
rect 813 -3159 816 -3153
rect 820 -3159 823 -3153
rect 827 -3159 830 -3153
rect 834 -3159 837 -3153
rect 841 -3159 847 -3153
rect 848 -3159 851 -3153
rect 855 -3159 861 -3153
rect 862 -3159 865 -3153
rect 869 -3159 872 -3153
rect 876 -3159 882 -3153
rect 883 -3159 886 -3153
rect 890 -3159 893 -3153
rect 897 -3159 900 -3153
rect 904 -3159 907 -3153
rect 911 -3159 914 -3153
rect 918 -3159 921 -3153
rect 925 -3159 928 -3153
rect 932 -3159 935 -3153
rect 939 -3159 942 -3153
rect 946 -3159 949 -3153
rect 953 -3159 956 -3153
rect 960 -3159 966 -3153
rect 967 -3159 970 -3153
rect 974 -3159 977 -3153
rect 981 -3159 984 -3153
rect 988 -3159 991 -3153
rect 995 -3159 1001 -3153
rect 1002 -3159 1005 -3153
rect 1009 -3159 1012 -3153
rect 1016 -3159 1019 -3153
rect 1023 -3159 1026 -3153
rect 1030 -3159 1033 -3153
rect 1037 -3159 1040 -3153
rect 1044 -3159 1047 -3153
rect 1051 -3159 1054 -3153
rect 1058 -3159 1061 -3153
rect 1065 -3159 1068 -3153
rect 1072 -3159 1075 -3153
rect 1079 -3159 1082 -3153
rect 1086 -3159 1092 -3153
rect 1093 -3159 1096 -3153
rect 1100 -3159 1103 -3153
rect 1107 -3159 1110 -3153
rect 1114 -3159 1117 -3153
rect 1121 -3159 1124 -3153
rect 1128 -3159 1131 -3153
rect 1135 -3159 1138 -3153
rect 1142 -3159 1145 -3153
rect 1149 -3159 1152 -3153
rect 1156 -3159 1159 -3153
rect 1163 -3159 1166 -3153
rect 1170 -3159 1173 -3153
rect 1177 -3159 1180 -3153
rect 1184 -3159 1190 -3153
rect 1191 -3159 1194 -3153
rect 1198 -3159 1201 -3153
rect 1205 -3159 1208 -3153
rect 1212 -3159 1215 -3153
rect 1219 -3159 1222 -3153
rect 1226 -3159 1232 -3153
rect 1233 -3159 1239 -3153
rect 1240 -3159 1246 -3153
rect 1261 -3159 1264 -3153
rect 1275 -3159 1278 -3153
rect 1289 -3159 1295 -3153
rect 1345 -3159 1348 -3153
rect 1352 -3159 1355 -3153
rect 1366 -3159 1369 -3153
rect 1408 -3159 1411 -3153
rect 1450 -3159 1453 -3153
rect 1457 -3159 1460 -3153
rect 1464 -3159 1467 -3153
rect 1 -3220 7 -3214
rect 57 -3220 60 -3214
rect 64 -3220 67 -3214
rect 71 -3220 74 -3214
rect 78 -3220 81 -3214
rect 85 -3220 88 -3214
rect 92 -3220 95 -3214
rect 99 -3220 102 -3214
rect 106 -3220 109 -3214
rect 113 -3220 119 -3214
rect 120 -3220 123 -3214
rect 127 -3220 133 -3214
rect 134 -3220 137 -3214
rect 141 -3220 147 -3214
rect 148 -3220 154 -3214
rect 155 -3220 158 -3214
rect 162 -3220 165 -3214
rect 169 -3220 175 -3214
rect 176 -3220 182 -3214
rect 183 -3220 186 -3214
rect 190 -3220 196 -3214
rect 197 -3220 203 -3214
rect 204 -3220 210 -3214
rect 211 -3220 214 -3214
rect 218 -3220 221 -3214
rect 225 -3220 228 -3214
rect 232 -3220 235 -3214
rect 239 -3220 242 -3214
rect 246 -3220 252 -3214
rect 253 -3220 256 -3214
rect 260 -3220 266 -3214
rect 267 -3220 270 -3214
rect 274 -3220 277 -3214
rect 281 -3220 284 -3214
rect 288 -3220 291 -3214
rect 295 -3220 298 -3214
rect 302 -3220 305 -3214
rect 309 -3220 312 -3214
rect 316 -3220 319 -3214
rect 323 -3220 329 -3214
rect 330 -3220 333 -3214
rect 337 -3220 340 -3214
rect 344 -3220 347 -3214
rect 351 -3220 354 -3214
rect 358 -3220 361 -3214
rect 365 -3220 368 -3214
rect 372 -3220 375 -3214
rect 379 -3220 382 -3214
rect 386 -3220 389 -3214
rect 393 -3220 396 -3214
rect 400 -3220 403 -3214
rect 407 -3220 410 -3214
rect 414 -3220 417 -3214
rect 421 -3220 424 -3214
rect 428 -3220 431 -3214
rect 435 -3220 438 -3214
rect 442 -3220 445 -3214
rect 449 -3220 452 -3214
rect 456 -3220 459 -3214
rect 463 -3220 466 -3214
rect 470 -3220 473 -3214
rect 477 -3220 480 -3214
rect 484 -3220 487 -3214
rect 491 -3220 494 -3214
rect 498 -3220 501 -3214
rect 505 -3220 508 -3214
rect 512 -3220 515 -3214
rect 519 -3220 522 -3214
rect 526 -3220 529 -3214
rect 533 -3220 536 -3214
rect 540 -3220 543 -3214
rect 547 -3220 550 -3214
rect 554 -3220 560 -3214
rect 561 -3220 564 -3214
rect 568 -3220 571 -3214
rect 575 -3220 581 -3214
rect 582 -3220 585 -3214
rect 589 -3220 592 -3214
rect 596 -3220 599 -3214
rect 603 -3220 609 -3214
rect 610 -3220 613 -3214
rect 617 -3220 620 -3214
rect 624 -3220 630 -3214
rect 631 -3220 637 -3214
rect 638 -3220 641 -3214
rect 645 -3220 648 -3214
rect 652 -3220 655 -3214
rect 659 -3220 665 -3214
rect 666 -3220 669 -3214
rect 673 -3220 676 -3214
rect 680 -3220 683 -3214
rect 687 -3220 690 -3214
rect 694 -3220 697 -3214
rect 701 -3220 704 -3214
rect 708 -3220 711 -3214
rect 715 -3220 718 -3214
rect 722 -3220 725 -3214
rect 729 -3220 732 -3214
rect 736 -3220 739 -3214
rect 743 -3220 746 -3214
rect 750 -3220 753 -3214
rect 757 -3220 763 -3214
rect 764 -3220 767 -3214
rect 771 -3220 774 -3214
rect 778 -3220 781 -3214
rect 785 -3220 788 -3214
rect 792 -3220 795 -3214
rect 799 -3220 802 -3214
rect 806 -3220 809 -3214
rect 813 -3220 816 -3214
rect 820 -3220 823 -3214
rect 827 -3220 830 -3214
rect 834 -3220 837 -3214
rect 841 -3220 844 -3214
rect 848 -3220 851 -3214
rect 855 -3220 858 -3214
rect 862 -3220 868 -3214
rect 869 -3220 872 -3214
rect 876 -3220 879 -3214
rect 883 -3220 886 -3214
rect 890 -3220 893 -3214
rect 897 -3220 900 -3214
rect 904 -3220 907 -3214
rect 911 -3220 914 -3214
rect 918 -3220 921 -3214
rect 925 -3220 928 -3214
rect 932 -3220 935 -3214
rect 939 -3220 942 -3214
rect 946 -3220 949 -3214
rect 953 -3220 956 -3214
rect 960 -3220 963 -3214
rect 967 -3220 970 -3214
rect 974 -3220 977 -3214
rect 981 -3220 987 -3214
rect 988 -3220 991 -3214
rect 995 -3220 998 -3214
rect 1002 -3220 1008 -3214
rect 1009 -3220 1012 -3214
rect 1016 -3220 1019 -3214
rect 1023 -3220 1026 -3214
rect 1030 -3220 1033 -3214
rect 1037 -3220 1040 -3214
rect 1044 -3220 1047 -3214
rect 1051 -3220 1054 -3214
rect 1058 -3220 1064 -3214
rect 1072 -3220 1075 -3214
rect 1079 -3220 1082 -3214
rect 1086 -3220 1089 -3214
rect 1093 -3220 1096 -3214
rect 1100 -3220 1103 -3214
rect 1107 -3220 1113 -3214
rect 1114 -3220 1117 -3214
rect 1121 -3220 1124 -3214
rect 1128 -3220 1131 -3214
rect 1135 -3220 1138 -3214
rect 1142 -3220 1145 -3214
rect 1149 -3220 1152 -3214
rect 1156 -3220 1162 -3214
rect 1163 -3220 1169 -3214
rect 1170 -3220 1173 -3214
rect 1184 -3220 1187 -3214
rect 1191 -3220 1194 -3214
rect 1198 -3220 1201 -3214
rect 1205 -3220 1208 -3214
rect 1212 -3220 1215 -3214
rect 1233 -3220 1236 -3214
rect 1331 -3220 1334 -3214
rect 1359 -3220 1362 -3214
rect 1366 -3220 1369 -3214
rect 1408 -3220 1411 -3214
rect 1450 -3220 1453 -3214
rect 1457 -3220 1460 -3214
rect 1464 -3220 1467 -3214
rect 155 -3275 158 -3269
rect 162 -3275 165 -3269
rect 169 -3275 172 -3269
rect 176 -3275 179 -3269
rect 183 -3275 189 -3269
rect 190 -3275 193 -3269
rect 197 -3275 200 -3269
rect 204 -3275 210 -3269
rect 211 -3275 214 -3269
rect 218 -3275 221 -3269
rect 225 -3275 228 -3269
rect 232 -3275 235 -3269
rect 239 -3275 245 -3269
rect 246 -3275 252 -3269
rect 253 -3275 256 -3269
rect 260 -3275 266 -3269
rect 267 -3275 270 -3269
rect 274 -3275 277 -3269
rect 281 -3275 284 -3269
rect 288 -3275 291 -3269
rect 295 -3275 298 -3269
rect 302 -3275 305 -3269
rect 309 -3275 312 -3269
rect 316 -3275 319 -3269
rect 323 -3275 326 -3269
rect 330 -3275 333 -3269
rect 337 -3275 340 -3269
rect 344 -3275 347 -3269
rect 351 -3275 354 -3269
rect 358 -3275 361 -3269
rect 365 -3275 368 -3269
rect 372 -3275 375 -3269
rect 379 -3275 382 -3269
rect 386 -3275 389 -3269
rect 393 -3275 399 -3269
rect 400 -3275 406 -3269
rect 407 -3275 410 -3269
rect 414 -3275 417 -3269
rect 421 -3275 424 -3269
rect 428 -3275 431 -3269
rect 435 -3275 438 -3269
rect 442 -3275 445 -3269
rect 449 -3275 452 -3269
rect 456 -3275 459 -3269
rect 463 -3275 466 -3269
rect 470 -3275 476 -3269
rect 477 -3275 480 -3269
rect 484 -3275 490 -3269
rect 491 -3275 494 -3269
rect 498 -3275 501 -3269
rect 505 -3275 508 -3269
rect 512 -3275 515 -3269
rect 519 -3275 522 -3269
rect 526 -3275 529 -3269
rect 533 -3275 536 -3269
rect 540 -3275 543 -3269
rect 547 -3275 550 -3269
rect 554 -3275 557 -3269
rect 561 -3275 564 -3269
rect 568 -3275 571 -3269
rect 575 -3275 578 -3269
rect 582 -3275 585 -3269
rect 589 -3275 595 -3269
rect 596 -3275 599 -3269
rect 603 -3275 606 -3269
rect 610 -3275 613 -3269
rect 617 -3275 620 -3269
rect 624 -3275 627 -3269
rect 631 -3275 637 -3269
rect 638 -3275 641 -3269
rect 645 -3275 648 -3269
rect 652 -3275 655 -3269
rect 659 -3275 662 -3269
rect 666 -3275 669 -3269
rect 673 -3275 676 -3269
rect 680 -3275 683 -3269
rect 687 -3275 690 -3269
rect 694 -3275 697 -3269
rect 701 -3275 704 -3269
rect 708 -3275 711 -3269
rect 715 -3275 718 -3269
rect 722 -3275 728 -3269
rect 729 -3275 735 -3269
rect 736 -3275 739 -3269
rect 743 -3275 746 -3269
rect 750 -3275 753 -3269
rect 757 -3275 760 -3269
rect 764 -3275 767 -3269
rect 771 -3275 774 -3269
rect 778 -3275 784 -3269
rect 785 -3275 788 -3269
rect 792 -3275 795 -3269
rect 799 -3275 802 -3269
rect 806 -3275 809 -3269
rect 813 -3275 816 -3269
rect 820 -3275 823 -3269
rect 827 -3275 830 -3269
rect 841 -3275 844 -3269
rect 869 -3275 872 -3269
rect 876 -3275 882 -3269
rect 883 -3275 886 -3269
rect 890 -3275 893 -3269
rect 897 -3275 900 -3269
rect 904 -3275 907 -3269
rect 911 -3275 914 -3269
rect 918 -3275 921 -3269
rect 925 -3275 928 -3269
rect 932 -3275 935 -3269
rect 939 -3275 942 -3269
rect 946 -3275 949 -3269
rect 953 -3275 956 -3269
rect 960 -3275 963 -3269
rect 981 -3275 984 -3269
rect 988 -3275 994 -3269
rect 995 -3275 998 -3269
rect 1002 -3275 1005 -3269
rect 1065 -3275 1068 -3269
rect 1072 -3275 1075 -3269
rect 1079 -3275 1082 -3269
rect 1093 -3275 1096 -3269
rect 1100 -3275 1103 -3269
rect 1107 -3275 1110 -3269
rect 1121 -3275 1127 -3269
rect 1128 -3275 1131 -3269
rect 1135 -3275 1138 -3269
rect 1142 -3275 1145 -3269
rect 1149 -3275 1152 -3269
rect 1156 -3275 1162 -3269
rect 1163 -3275 1166 -3269
rect 1170 -3275 1173 -3269
rect 1184 -3275 1190 -3269
rect 1205 -3275 1208 -3269
rect 1212 -3275 1218 -3269
rect 1219 -3275 1222 -3269
rect 1233 -3275 1239 -3269
rect 1247 -3275 1253 -3269
rect 1289 -3275 1292 -3269
rect 1324 -3275 1330 -3269
rect 1359 -3275 1362 -3269
rect 1366 -3275 1369 -3269
rect 1408 -3275 1411 -3269
rect 1450 -3275 1453 -3269
rect 1457 -3275 1463 -3269
rect 1464 -3275 1467 -3269
rect 176 -3338 179 -3332
rect 183 -3338 186 -3332
rect 190 -3338 193 -3332
rect 197 -3338 200 -3332
rect 204 -3338 207 -3332
rect 211 -3338 214 -3332
rect 218 -3338 221 -3332
rect 225 -3338 231 -3332
rect 232 -3338 235 -3332
rect 239 -3338 242 -3332
rect 246 -3338 249 -3332
rect 253 -3338 256 -3332
rect 260 -3338 266 -3332
rect 267 -3338 270 -3332
rect 274 -3338 277 -3332
rect 281 -3338 284 -3332
rect 288 -3338 291 -3332
rect 295 -3338 298 -3332
rect 302 -3338 305 -3332
rect 309 -3338 312 -3332
rect 316 -3338 319 -3332
rect 323 -3338 326 -3332
rect 330 -3338 333 -3332
rect 337 -3338 340 -3332
rect 344 -3338 347 -3332
rect 351 -3338 354 -3332
rect 358 -3338 361 -3332
rect 365 -3338 368 -3332
rect 372 -3338 375 -3332
rect 379 -3338 385 -3332
rect 386 -3338 389 -3332
rect 393 -3338 396 -3332
rect 400 -3338 403 -3332
rect 407 -3338 413 -3332
rect 414 -3338 417 -3332
rect 421 -3338 424 -3332
rect 428 -3338 431 -3332
rect 435 -3338 438 -3332
rect 442 -3338 448 -3332
rect 449 -3338 452 -3332
rect 456 -3338 459 -3332
rect 463 -3338 469 -3332
rect 470 -3338 473 -3332
rect 477 -3338 480 -3332
rect 484 -3338 487 -3332
rect 491 -3338 494 -3332
rect 498 -3338 501 -3332
rect 505 -3338 508 -3332
rect 512 -3338 515 -3332
rect 519 -3338 522 -3332
rect 526 -3338 529 -3332
rect 533 -3338 536 -3332
rect 540 -3338 546 -3332
rect 547 -3338 550 -3332
rect 554 -3338 557 -3332
rect 561 -3338 564 -3332
rect 568 -3338 574 -3332
rect 575 -3338 578 -3332
rect 582 -3338 585 -3332
rect 589 -3338 595 -3332
rect 596 -3338 599 -3332
rect 603 -3338 606 -3332
rect 610 -3338 613 -3332
rect 617 -3338 623 -3332
rect 624 -3338 627 -3332
rect 631 -3338 634 -3332
rect 638 -3338 641 -3332
rect 645 -3338 648 -3332
rect 652 -3338 655 -3332
rect 659 -3338 662 -3332
rect 666 -3338 672 -3332
rect 673 -3338 676 -3332
rect 680 -3338 686 -3332
rect 687 -3338 690 -3332
rect 694 -3338 697 -3332
rect 701 -3338 704 -3332
rect 708 -3338 714 -3332
rect 715 -3338 718 -3332
rect 722 -3338 725 -3332
rect 729 -3338 732 -3332
rect 736 -3338 742 -3332
rect 743 -3338 746 -3332
rect 750 -3338 753 -3332
rect 757 -3338 760 -3332
rect 764 -3338 767 -3332
rect 771 -3338 774 -3332
rect 778 -3338 781 -3332
rect 785 -3338 788 -3332
rect 792 -3338 795 -3332
rect 799 -3338 802 -3332
rect 806 -3338 809 -3332
rect 813 -3338 816 -3332
rect 820 -3338 823 -3332
rect 827 -3338 830 -3332
rect 834 -3338 840 -3332
rect 841 -3338 847 -3332
rect 848 -3338 851 -3332
rect 855 -3338 858 -3332
rect 862 -3338 865 -3332
rect 869 -3338 872 -3332
rect 876 -3338 879 -3332
rect 883 -3338 886 -3332
rect 890 -3338 893 -3332
rect 897 -3338 900 -3332
rect 904 -3338 907 -3332
rect 911 -3338 914 -3332
rect 918 -3338 921 -3332
rect 925 -3338 928 -3332
rect 932 -3338 938 -3332
rect 939 -3338 942 -3332
rect 946 -3338 952 -3332
rect 953 -3338 956 -3332
rect 960 -3338 963 -3332
rect 974 -3338 977 -3332
rect 988 -3338 991 -3332
rect 1058 -3338 1064 -3332
rect 1065 -3338 1068 -3332
rect 1072 -3338 1075 -3332
rect 1079 -3338 1082 -3332
rect 1093 -3338 1099 -3332
rect 1107 -3338 1110 -3332
rect 1114 -3338 1117 -3332
rect 1135 -3338 1141 -3332
rect 1142 -3338 1145 -3332
rect 1212 -3338 1215 -3332
rect 1289 -3338 1292 -3332
rect 1359 -3338 1362 -3332
rect 1366 -3338 1369 -3332
rect 1408 -3338 1411 -3332
rect 176 -3403 179 -3397
rect 183 -3403 186 -3397
rect 190 -3403 193 -3397
rect 197 -3403 200 -3397
rect 204 -3403 207 -3397
rect 211 -3403 214 -3397
rect 218 -3403 221 -3397
rect 225 -3403 231 -3397
rect 232 -3403 235 -3397
rect 239 -3403 242 -3397
rect 246 -3403 249 -3397
rect 253 -3403 256 -3397
rect 260 -3403 263 -3397
rect 267 -3403 270 -3397
rect 274 -3403 277 -3397
rect 281 -3403 284 -3397
rect 288 -3403 291 -3397
rect 295 -3403 298 -3397
rect 302 -3403 305 -3397
rect 309 -3403 312 -3397
rect 316 -3403 319 -3397
rect 323 -3403 326 -3397
rect 330 -3403 333 -3397
rect 337 -3403 343 -3397
rect 344 -3403 347 -3397
rect 351 -3403 357 -3397
rect 358 -3403 361 -3397
rect 365 -3403 368 -3397
rect 372 -3403 375 -3397
rect 379 -3403 385 -3397
rect 386 -3403 389 -3397
rect 393 -3403 399 -3397
rect 400 -3403 403 -3397
rect 407 -3403 410 -3397
rect 414 -3403 417 -3397
rect 421 -3403 424 -3397
rect 428 -3403 431 -3397
rect 435 -3403 438 -3397
rect 442 -3403 445 -3397
rect 449 -3403 452 -3397
rect 456 -3403 459 -3397
rect 463 -3403 469 -3397
rect 470 -3403 473 -3397
rect 477 -3403 480 -3397
rect 484 -3403 490 -3397
rect 491 -3403 497 -3397
rect 498 -3403 501 -3397
rect 505 -3403 511 -3397
rect 512 -3403 515 -3397
rect 519 -3403 522 -3397
rect 526 -3403 529 -3397
rect 533 -3403 539 -3397
rect 540 -3403 546 -3397
rect 547 -3403 550 -3397
rect 554 -3403 560 -3397
rect 561 -3403 564 -3397
rect 568 -3403 571 -3397
rect 575 -3403 581 -3397
rect 582 -3403 585 -3397
rect 589 -3403 592 -3397
rect 596 -3403 599 -3397
rect 603 -3403 606 -3397
rect 610 -3403 613 -3397
rect 617 -3403 620 -3397
rect 624 -3403 627 -3397
rect 631 -3403 634 -3397
rect 638 -3403 641 -3397
rect 645 -3403 648 -3397
rect 652 -3403 655 -3397
rect 659 -3403 662 -3397
rect 666 -3403 669 -3397
rect 673 -3403 676 -3397
rect 680 -3403 683 -3397
rect 687 -3403 690 -3397
rect 694 -3403 697 -3397
rect 701 -3403 707 -3397
rect 708 -3403 711 -3397
rect 715 -3403 718 -3397
rect 722 -3403 725 -3397
rect 729 -3403 732 -3397
rect 736 -3403 739 -3397
rect 743 -3403 746 -3397
rect 750 -3403 753 -3397
rect 757 -3403 760 -3397
rect 764 -3403 767 -3397
rect 771 -3403 777 -3397
rect 778 -3403 781 -3397
rect 813 -3403 816 -3397
rect 820 -3403 823 -3397
rect 827 -3403 833 -3397
rect 834 -3403 837 -3397
rect 841 -3403 847 -3397
rect 848 -3403 851 -3397
rect 855 -3403 858 -3397
rect 862 -3403 868 -3397
rect 869 -3403 872 -3397
rect 876 -3403 879 -3397
rect 883 -3403 886 -3397
rect 890 -3403 896 -3397
rect 904 -3403 907 -3397
rect 911 -3403 914 -3397
rect 918 -3403 921 -3397
rect 925 -3403 928 -3397
rect 939 -3403 942 -3397
rect 988 -3403 991 -3397
rect 995 -3403 998 -3397
rect 1072 -3403 1075 -3397
rect 1114 -3403 1117 -3397
rect 1121 -3403 1124 -3397
rect 1212 -3403 1215 -3397
rect 1352 -3403 1355 -3397
rect 1359 -3403 1362 -3397
rect 1366 -3403 1369 -3397
rect 1408 -3403 1411 -3397
rect 218 -3446 224 -3440
rect 239 -3446 242 -3440
rect 253 -3446 256 -3440
rect 260 -3446 266 -3440
rect 267 -3446 270 -3440
rect 274 -3446 277 -3440
rect 281 -3446 284 -3440
rect 288 -3446 294 -3440
rect 295 -3446 298 -3440
rect 302 -3446 308 -3440
rect 309 -3446 312 -3440
rect 316 -3446 319 -3440
rect 323 -3446 329 -3440
rect 337 -3446 343 -3440
rect 344 -3446 347 -3440
rect 351 -3446 354 -3440
rect 358 -3446 361 -3440
rect 372 -3446 375 -3440
rect 386 -3446 389 -3440
rect 393 -3446 396 -3440
rect 400 -3446 403 -3440
rect 407 -3446 410 -3440
rect 421 -3446 424 -3440
rect 428 -3446 431 -3440
rect 435 -3446 438 -3440
rect 442 -3446 445 -3440
rect 449 -3446 452 -3440
rect 470 -3446 473 -3440
rect 484 -3446 487 -3440
rect 491 -3446 494 -3440
rect 498 -3446 504 -3440
rect 533 -3446 536 -3440
rect 540 -3446 543 -3440
rect 547 -3446 550 -3440
rect 554 -3446 557 -3440
rect 561 -3446 564 -3440
rect 568 -3446 574 -3440
rect 575 -3446 578 -3440
rect 582 -3446 585 -3440
rect 596 -3446 599 -3440
rect 624 -3446 627 -3440
rect 631 -3446 634 -3440
rect 638 -3446 644 -3440
rect 645 -3446 648 -3440
rect 652 -3446 655 -3440
rect 659 -3446 662 -3440
rect 666 -3446 669 -3440
rect 673 -3446 676 -3440
rect 680 -3446 683 -3440
rect 687 -3446 690 -3440
rect 694 -3446 697 -3440
rect 701 -3446 704 -3440
rect 708 -3446 711 -3440
rect 715 -3446 721 -3440
rect 722 -3446 728 -3440
rect 729 -3446 732 -3440
rect 736 -3446 742 -3440
rect 743 -3446 746 -3440
rect 750 -3446 753 -3440
rect 757 -3446 760 -3440
rect 764 -3446 767 -3440
rect 771 -3446 777 -3440
rect 778 -3446 784 -3440
rect 820 -3446 823 -3440
rect 827 -3446 833 -3440
rect 834 -3446 837 -3440
rect 841 -3446 844 -3440
rect 848 -3446 851 -3440
rect 855 -3446 858 -3440
rect 862 -3446 865 -3440
rect 869 -3446 872 -3440
rect 883 -3446 886 -3440
rect 911 -3446 914 -3440
rect 918 -3446 921 -3440
rect 925 -3446 928 -3440
rect 939 -3446 942 -3440
rect 946 -3446 949 -3440
rect 953 -3446 959 -3440
rect 960 -3446 966 -3440
rect 967 -3446 970 -3440
rect 974 -3446 980 -3440
rect 981 -3446 984 -3440
rect 988 -3446 991 -3440
rect 995 -3446 998 -3440
rect 1009 -3446 1012 -3440
rect 1072 -3446 1075 -3440
rect 1093 -3446 1096 -3440
rect 1114 -3446 1117 -3440
rect 1121 -3446 1124 -3440
rect 1212 -3446 1215 -3440
rect 1352 -3446 1355 -3440
rect 1359 -3446 1362 -3440
rect 1394 -3446 1397 -3440
rect 1408 -3446 1411 -3440
rect 253 -3473 256 -3467
rect 260 -3473 263 -3467
rect 302 -3473 305 -3467
rect 316 -3473 319 -3467
rect 323 -3473 329 -3467
rect 330 -3473 333 -3467
rect 337 -3473 340 -3467
rect 351 -3473 354 -3467
rect 358 -3473 361 -3467
rect 379 -3473 382 -3467
rect 393 -3473 396 -3467
rect 400 -3473 403 -3467
rect 407 -3473 413 -3467
rect 414 -3473 417 -3467
rect 421 -3473 427 -3467
rect 428 -3473 431 -3467
rect 435 -3473 441 -3467
rect 442 -3473 445 -3467
rect 456 -3473 462 -3467
rect 463 -3473 469 -3467
rect 470 -3473 476 -3467
rect 477 -3473 480 -3467
rect 484 -3473 487 -3467
rect 491 -3473 494 -3467
rect 498 -3473 504 -3467
rect 505 -3473 508 -3467
rect 512 -3473 518 -3467
rect 519 -3473 522 -3467
rect 540 -3473 543 -3467
rect 547 -3473 550 -3467
rect 554 -3473 557 -3467
rect 561 -3473 564 -3467
rect 568 -3473 571 -3467
rect 575 -3473 578 -3467
rect 582 -3473 585 -3467
rect 603 -3473 606 -3467
rect 610 -3473 616 -3467
rect 617 -3473 623 -3467
rect 624 -3473 627 -3467
rect 645 -3473 648 -3467
rect 652 -3473 655 -3467
rect 659 -3473 662 -3467
rect 673 -3473 676 -3467
rect 680 -3473 683 -3467
rect 687 -3473 693 -3467
rect 694 -3473 700 -3467
rect 708 -3473 711 -3467
rect 736 -3473 739 -3467
rect 757 -3473 760 -3467
rect 820 -3473 826 -3467
rect 834 -3473 837 -3467
rect 841 -3473 844 -3467
rect 848 -3473 854 -3467
rect 855 -3473 858 -3467
rect 869 -3473 872 -3467
rect 883 -3473 886 -3467
rect 890 -3473 893 -3467
rect 911 -3473 914 -3467
rect 918 -3473 921 -3467
rect 925 -3473 928 -3467
rect 932 -3473 935 -3467
rect 939 -3473 942 -3467
rect 988 -3473 991 -3467
rect 995 -3473 998 -3467
rect 1065 -3473 1068 -3467
rect 1072 -3473 1078 -3467
rect 1114 -3473 1117 -3467
rect 1121 -3473 1124 -3467
rect 1212 -3473 1215 -3467
rect 1219 -3473 1225 -3467
rect 1226 -3473 1229 -3467
rect 1352 -3473 1355 -3467
rect 1359 -3473 1362 -3467
rect 1408 -3473 1411 -3467
rect 1415 -3473 1418 -3467
rect 260 -3496 263 -3490
rect 267 -3496 270 -3490
rect 309 -3496 312 -3490
rect 330 -3496 333 -3490
rect 337 -3496 340 -3490
rect 344 -3496 350 -3490
rect 351 -3496 354 -3490
rect 407 -3496 410 -3490
rect 414 -3496 420 -3490
rect 428 -3496 434 -3490
rect 435 -3496 438 -3490
rect 477 -3496 480 -3490
rect 540 -3496 543 -3490
rect 547 -3496 550 -3490
rect 554 -3496 557 -3490
rect 568 -3496 571 -3490
rect 575 -3496 578 -3490
rect 582 -3496 585 -3490
rect 589 -3496 592 -3490
rect 596 -3496 602 -3490
rect 645 -3496 651 -3490
rect 652 -3496 655 -3490
rect 659 -3496 662 -3490
rect 680 -3496 683 -3490
rect 687 -3496 690 -3490
rect 715 -3496 718 -3490
rect 722 -3496 728 -3490
rect 827 -3496 830 -3490
rect 834 -3496 837 -3490
rect 841 -3496 847 -3490
rect 848 -3496 851 -3490
rect 876 -3496 879 -3490
rect 883 -3496 889 -3490
rect 897 -3496 903 -3490
rect 904 -3496 907 -3490
rect 911 -3496 914 -3490
rect 918 -3496 921 -3490
rect 925 -3496 928 -3490
rect 939 -3496 942 -3490
rect 946 -3496 952 -3490
rect 988 -3496 994 -3490
rect 995 -3496 998 -3490
rect 1093 -3496 1096 -3490
rect 1114 -3496 1120 -3490
rect 1121 -3496 1124 -3490
rect 1219 -3496 1225 -3490
rect 1352 -3496 1355 -3490
rect 1359 -3496 1362 -3490
rect 1408 -3496 1414 -3490
rect 1415 -3496 1418 -3490
rect 267 -3511 273 -3505
rect 274 -3511 277 -3505
rect 323 -3511 329 -3505
rect 330 -3511 333 -3505
rect 351 -3511 357 -3505
rect 358 -3511 361 -3505
rect 540 -3511 543 -3505
rect 547 -3511 553 -3505
rect 554 -3511 560 -3505
rect 561 -3511 567 -3505
rect 568 -3511 571 -3505
rect 575 -3511 581 -3505
rect 582 -3511 585 -3505
rect 659 -3511 665 -3505
rect 666 -3511 669 -3505
rect 687 -3511 693 -3505
rect 855 -3511 861 -3505
rect 869 -3511 872 -3505
rect 876 -3511 879 -3505
rect 911 -3511 917 -3505
rect 918 -3511 924 -3505
rect 1352 -3511 1355 -3505
rect 1359 -3511 1365 -3505
rect 1366 -3511 1369 -3505
<< polysilicon >>
rect 282 -7 283 -5
rect 285 -13 286 -11
rect 317 -7 318 -5
rect 317 -13 318 -11
rect 345 -7 346 -5
rect 345 -13 346 -11
rect 352 -7 353 -5
rect 352 -13 353 -11
rect 425 -7 426 -5
rect 425 -13 426 -11
rect 436 -7 437 -5
rect 436 -13 437 -11
rect 443 -7 444 -5
rect 443 -13 444 -11
rect 450 -7 451 -5
rect 450 -13 451 -11
rect 457 -7 458 -5
rect 460 -13 461 -11
rect 464 -7 465 -5
rect 464 -13 465 -11
rect 478 -7 479 -5
rect 478 -13 479 -11
rect 506 -13 507 -11
rect 509 -13 510 -11
rect 513 -7 514 -5
rect 513 -13 514 -11
rect 905 -7 906 -5
rect 905 -13 906 -11
rect 947 -7 948 -5
rect 950 -7 951 -5
rect 989 -7 990 -5
rect 989 -13 990 -11
rect 226 -26 227 -24
rect 226 -32 227 -30
rect 289 -26 290 -24
rect 289 -32 290 -30
rect 303 -26 304 -24
rect 303 -32 304 -30
rect 338 -26 339 -24
rect 338 -32 339 -30
rect 345 -26 346 -24
rect 348 -26 349 -24
rect 352 -26 353 -24
rect 352 -32 353 -30
rect 359 -26 360 -24
rect 362 -26 363 -24
rect 366 -26 367 -24
rect 366 -32 367 -30
rect 373 -26 374 -24
rect 373 -32 374 -30
rect 380 -26 381 -24
rect 380 -32 381 -30
rect 387 -26 388 -24
rect 387 -32 388 -30
rect 394 -26 395 -24
rect 394 -32 395 -30
rect 408 -26 409 -24
rect 408 -32 409 -30
rect 418 -26 419 -24
rect 418 -32 419 -30
rect 422 -26 423 -24
rect 422 -32 423 -30
rect 436 -26 437 -24
rect 436 -32 437 -30
rect 450 -26 451 -24
rect 450 -32 451 -30
rect 457 -26 458 -24
rect 457 -32 458 -30
rect 464 -26 465 -24
rect 464 -32 465 -30
rect 499 -26 500 -24
rect 499 -32 500 -30
rect 509 -26 510 -24
rect 506 -32 507 -30
rect 513 -26 514 -24
rect 513 -32 514 -30
rect 520 -32 521 -30
rect 523 -32 524 -30
rect 527 -26 528 -24
rect 527 -32 528 -30
rect 537 -26 538 -24
rect 537 -32 538 -30
rect 541 -26 542 -24
rect 541 -32 542 -30
rect 548 -26 549 -24
rect 548 -32 549 -30
rect 579 -26 580 -24
rect 583 -26 584 -24
rect 590 -26 591 -24
rect 590 -32 591 -30
rect 597 -26 598 -24
rect 597 -32 598 -30
rect 604 -26 605 -24
rect 604 -32 605 -30
rect 611 -26 612 -24
rect 611 -32 612 -30
rect 618 -26 619 -24
rect 625 -26 626 -24
rect 625 -32 626 -30
rect 635 -32 636 -30
rect 639 -26 640 -24
rect 639 -32 640 -30
rect 674 -26 675 -24
rect 674 -32 675 -30
rect 891 -26 892 -24
rect 891 -32 892 -30
rect 1003 -26 1004 -24
rect 1003 -32 1004 -30
rect 219 -49 220 -47
rect 219 -55 220 -53
rect 275 -49 276 -47
rect 275 -55 276 -53
rect 282 -49 283 -47
rect 282 -55 283 -53
rect 296 -49 297 -47
rect 299 -55 300 -53
rect 303 -49 304 -47
rect 303 -55 304 -53
rect 320 -55 321 -53
rect 324 -49 325 -47
rect 324 -55 325 -53
rect 331 -49 332 -47
rect 331 -55 332 -53
rect 338 -49 339 -47
rect 341 -49 342 -47
rect 338 -55 339 -53
rect 341 -55 342 -53
rect 345 -49 346 -47
rect 345 -55 346 -53
rect 352 -49 353 -47
rect 352 -55 353 -53
rect 359 -49 360 -47
rect 359 -55 360 -53
rect 366 -49 367 -47
rect 366 -55 367 -53
rect 373 -49 374 -47
rect 373 -55 374 -53
rect 380 -49 381 -47
rect 380 -55 381 -53
rect 387 -49 388 -47
rect 390 -55 391 -53
rect 394 -49 395 -47
rect 394 -55 395 -53
rect 401 -49 402 -47
rect 401 -55 402 -53
rect 408 -49 409 -47
rect 408 -55 409 -53
rect 415 -49 416 -47
rect 415 -55 416 -53
rect 422 -49 423 -47
rect 422 -55 423 -53
rect 429 -49 430 -47
rect 432 -49 433 -47
rect 429 -55 430 -53
rect 436 -49 437 -47
rect 436 -55 437 -53
rect 443 -49 444 -47
rect 443 -55 444 -53
rect 450 -49 451 -47
rect 450 -55 451 -53
rect 457 -49 458 -47
rect 457 -55 458 -53
rect 464 -49 465 -47
rect 464 -55 465 -53
rect 471 -49 472 -47
rect 471 -55 472 -53
rect 485 -49 486 -47
rect 485 -55 486 -53
rect 492 -49 493 -47
rect 492 -55 493 -53
rect 499 -49 500 -47
rect 499 -55 500 -53
rect 506 -49 507 -47
rect 506 -55 507 -53
rect 520 -49 521 -47
rect 520 -55 521 -53
rect 541 -49 542 -47
rect 541 -55 542 -53
rect 551 -49 552 -47
rect 548 -55 549 -53
rect 555 -49 556 -47
rect 555 -55 556 -53
rect 565 -49 566 -47
rect 562 -55 563 -53
rect 569 -55 570 -53
rect 572 -55 573 -53
rect 576 -49 577 -47
rect 576 -55 577 -53
rect 583 -49 584 -47
rect 583 -55 584 -53
rect 590 -49 591 -47
rect 590 -55 591 -53
rect 597 -49 598 -47
rect 597 -55 598 -53
rect 604 -49 605 -47
rect 604 -55 605 -53
rect 611 -55 612 -53
rect 614 -55 615 -53
rect 621 -49 622 -47
rect 621 -55 622 -53
rect 625 -49 626 -47
rect 625 -55 626 -53
rect 632 -49 633 -47
rect 632 -55 633 -53
rect 639 -49 640 -47
rect 639 -55 640 -53
rect 653 -49 654 -47
rect 653 -55 654 -53
rect 674 -49 675 -47
rect 674 -55 675 -53
rect 681 -49 682 -47
rect 681 -55 682 -53
rect 723 -49 724 -47
rect 723 -55 724 -53
rect 730 -49 731 -47
rect 730 -55 731 -53
rect 758 -49 759 -47
rect 758 -55 759 -53
rect 828 -49 829 -47
rect 828 -55 829 -53
rect 884 -49 885 -47
rect 884 -55 885 -53
rect 1010 -49 1011 -47
rect 1010 -55 1011 -53
rect 191 -100 192 -98
rect 191 -106 192 -104
rect 205 -100 206 -98
rect 205 -106 206 -104
rect 219 -100 220 -98
rect 219 -106 220 -104
rect 233 -100 234 -98
rect 233 -106 234 -104
rect 240 -100 241 -98
rect 243 -100 244 -98
rect 247 -100 248 -98
rect 247 -106 248 -104
rect 254 -100 255 -98
rect 254 -106 255 -104
rect 257 -106 258 -104
rect 261 -100 262 -98
rect 261 -106 262 -104
rect 271 -106 272 -104
rect 275 -100 276 -98
rect 278 -100 279 -98
rect 275 -106 276 -104
rect 282 -100 283 -98
rect 282 -106 283 -104
rect 289 -100 290 -98
rect 289 -106 290 -104
rect 296 -100 297 -98
rect 299 -100 300 -98
rect 299 -106 300 -104
rect 303 -100 304 -98
rect 303 -106 304 -104
rect 310 -100 311 -98
rect 310 -106 311 -104
rect 317 -100 318 -98
rect 317 -106 318 -104
rect 324 -100 325 -98
rect 324 -106 325 -104
rect 331 -100 332 -98
rect 331 -106 332 -104
rect 338 -100 339 -98
rect 338 -106 339 -104
rect 345 -100 346 -98
rect 345 -106 346 -104
rect 352 -100 353 -98
rect 352 -106 353 -104
rect 359 -100 360 -98
rect 359 -106 360 -104
rect 366 -100 367 -98
rect 366 -106 367 -104
rect 373 -100 374 -98
rect 373 -106 374 -104
rect 380 -100 381 -98
rect 383 -100 384 -98
rect 383 -106 384 -104
rect 390 -100 391 -98
rect 387 -106 388 -104
rect 390 -106 391 -104
rect 394 -100 395 -98
rect 394 -106 395 -104
rect 401 -100 402 -98
rect 401 -106 402 -104
rect 408 -100 409 -98
rect 408 -106 409 -104
rect 415 -100 416 -98
rect 415 -106 416 -104
rect 422 -100 423 -98
rect 422 -106 423 -104
rect 429 -100 430 -98
rect 429 -106 430 -104
rect 436 -100 437 -98
rect 436 -106 437 -104
rect 443 -100 444 -98
rect 443 -106 444 -104
rect 450 -100 451 -98
rect 450 -106 451 -104
rect 457 -100 458 -98
rect 457 -106 458 -104
rect 464 -100 465 -98
rect 464 -106 465 -104
rect 471 -100 472 -98
rect 471 -106 472 -104
rect 478 -100 479 -98
rect 478 -106 479 -104
rect 485 -100 486 -98
rect 485 -106 486 -104
rect 492 -100 493 -98
rect 492 -106 493 -104
rect 499 -100 500 -98
rect 499 -106 500 -104
rect 509 -100 510 -98
rect 506 -106 507 -104
rect 509 -106 510 -104
rect 513 -100 514 -98
rect 516 -100 517 -98
rect 513 -106 514 -104
rect 516 -106 517 -104
rect 520 -100 521 -98
rect 523 -100 524 -98
rect 520 -106 521 -104
rect 527 -100 528 -98
rect 527 -106 528 -104
rect 534 -100 535 -98
rect 537 -106 538 -104
rect 541 -106 542 -104
rect 548 -100 549 -98
rect 548 -106 549 -104
rect 555 -100 556 -98
rect 555 -106 556 -104
rect 562 -106 563 -104
rect 565 -106 566 -104
rect 569 -100 570 -98
rect 569 -106 570 -104
rect 576 -100 577 -98
rect 576 -106 577 -104
rect 586 -100 587 -98
rect 583 -106 584 -104
rect 586 -106 587 -104
rect 590 -100 591 -98
rect 590 -106 591 -104
rect 597 -100 598 -98
rect 597 -106 598 -104
rect 604 -100 605 -98
rect 604 -106 605 -104
rect 611 -100 612 -98
rect 611 -106 612 -104
rect 618 -100 619 -98
rect 618 -106 619 -104
rect 628 -100 629 -98
rect 625 -106 626 -104
rect 628 -106 629 -104
rect 632 -100 633 -98
rect 632 -106 633 -104
rect 639 -100 640 -98
rect 639 -106 640 -104
rect 646 -100 647 -98
rect 646 -106 647 -104
rect 653 -100 654 -98
rect 653 -106 654 -104
rect 660 -100 661 -98
rect 660 -106 661 -104
rect 667 -100 668 -98
rect 667 -106 668 -104
rect 681 -100 682 -98
rect 681 -106 682 -104
rect 688 -100 689 -98
rect 688 -106 689 -104
rect 702 -100 703 -98
rect 702 -106 703 -104
rect 709 -100 710 -98
rect 709 -106 710 -104
rect 723 -100 724 -98
rect 723 -106 724 -104
rect 730 -100 731 -98
rect 730 -106 731 -104
rect 737 -100 738 -98
rect 737 -106 738 -104
rect 779 -100 780 -98
rect 782 -100 783 -98
rect 782 -106 783 -104
rect 789 -100 790 -98
rect 786 -106 787 -104
rect 793 -100 794 -98
rect 793 -106 794 -104
rect 800 -100 801 -98
rect 800 -106 801 -104
rect 807 -100 808 -98
rect 807 -106 808 -104
rect 863 -100 864 -98
rect 863 -106 864 -104
rect 891 -100 892 -98
rect 891 -106 892 -104
rect 898 -100 899 -98
rect 898 -106 899 -104
rect 1017 -100 1018 -98
rect 1017 -106 1018 -104
rect 114 -167 115 -165
rect 114 -173 115 -171
rect 121 -167 122 -165
rect 121 -173 122 -171
rect 128 -167 129 -165
rect 128 -173 129 -171
rect 135 -167 136 -165
rect 135 -173 136 -171
rect 142 -167 143 -165
rect 142 -173 143 -171
rect 149 -167 150 -165
rect 149 -173 150 -171
rect 156 -167 157 -165
rect 156 -173 157 -171
rect 163 -167 164 -165
rect 163 -173 164 -171
rect 170 -167 171 -165
rect 170 -173 171 -171
rect 177 -167 178 -165
rect 177 -173 178 -171
rect 184 -167 185 -165
rect 184 -173 185 -171
rect 191 -167 192 -165
rect 191 -173 192 -171
rect 198 -167 199 -165
rect 198 -173 199 -171
rect 205 -167 206 -165
rect 205 -173 206 -171
rect 212 -167 213 -165
rect 212 -173 213 -171
rect 219 -167 220 -165
rect 219 -173 220 -171
rect 226 -167 227 -165
rect 229 -167 230 -165
rect 226 -173 227 -171
rect 233 -167 234 -165
rect 233 -173 234 -171
rect 240 -167 241 -165
rect 240 -173 241 -171
rect 247 -167 248 -165
rect 247 -173 248 -171
rect 254 -167 255 -165
rect 254 -173 255 -171
rect 261 -167 262 -165
rect 261 -173 262 -171
rect 268 -167 269 -165
rect 268 -173 269 -171
rect 275 -167 276 -165
rect 275 -173 276 -171
rect 282 -167 283 -165
rect 282 -173 283 -171
rect 289 -167 290 -165
rect 289 -173 290 -171
rect 296 -167 297 -165
rect 299 -167 300 -165
rect 296 -173 297 -171
rect 303 -167 304 -165
rect 303 -173 304 -171
rect 310 -167 311 -165
rect 310 -173 311 -171
rect 317 -167 318 -165
rect 317 -173 318 -171
rect 324 -167 325 -165
rect 324 -173 325 -171
rect 331 -167 332 -165
rect 334 -167 335 -165
rect 331 -173 332 -171
rect 334 -173 335 -171
rect 338 -167 339 -165
rect 338 -173 339 -171
rect 345 -167 346 -165
rect 345 -173 346 -171
rect 352 -167 353 -165
rect 352 -173 353 -171
rect 359 -167 360 -165
rect 359 -173 360 -171
rect 366 -167 367 -165
rect 369 -167 370 -165
rect 369 -173 370 -171
rect 373 -167 374 -165
rect 373 -173 374 -171
rect 380 -167 381 -165
rect 380 -173 381 -171
rect 390 -167 391 -165
rect 387 -173 388 -171
rect 390 -173 391 -171
rect 394 -167 395 -165
rect 394 -173 395 -171
rect 401 -167 402 -165
rect 401 -173 402 -171
rect 404 -173 405 -171
rect 408 -167 409 -165
rect 408 -173 409 -171
rect 415 -167 416 -165
rect 415 -173 416 -171
rect 422 -167 423 -165
rect 422 -173 423 -171
rect 429 -167 430 -165
rect 429 -173 430 -171
rect 436 -167 437 -165
rect 436 -173 437 -171
rect 443 -167 444 -165
rect 443 -173 444 -171
rect 450 -167 451 -165
rect 453 -167 454 -165
rect 450 -173 451 -171
rect 457 -167 458 -165
rect 457 -173 458 -171
rect 464 -167 465 -165
rect 464 -173 465 -171
rect 471 -167 472 -165
rect 471 -173 472 -171
rect 478 -167 479 -165
rect 478 -173 479 -171
rect 485 -167 486 -165
rect 485 -173 486 -171
rect 492 -167 493 -165
rect 492 -173 493 -171
rect 499 -167 500 -165
rect 502 -167 503 -165
rect 499 -173 500 -171
rect 506 -167 507 -165
rect 506 -173 507 -171
rect 513 -167 514 -165
rect 516 -167 517 -165
rect 513 -173 514 -171
rect 523 -167 524 -165
rect 520 -173 521 -171
rect 523 -173 524 -171
rect 527 -167 528 -165
rect 530 -167 531 -165
rect 530 -173 531 -171
rect 534 -167 535 -165
rect 534 -173 535 -171
rect 541 -167 542 -165
rect 541 -173 542 -171
rect 548 -167 549 -165
rect 548 -173 549 -171
rect 555 -167 556 -165
rect 558 -167 559 -165
rect 558 -173 559 -171
rect 562 -167 563 -165
rect 562 -173 563 -171
rect 569 -167 570 -165
rect 572 -167 573 -165
rect 569 -173 570 -171
rect 576 -167 577 -165
rect 576 -173 577 -171
rect 583 -167 584 -165
rect 583 -173 584 -171
rect 593 -167 594 -165
rect 593 -173 594 -171
rect 597 -167 598 -165
rect 597 -173 598 -171
rect 604 -167 605 -165
rect 607 -173 608 -171
rect 611 -167 612 -165
rect 614 -167 615 -165
rect 611 -173 612 -171
rect 618 -167 619 -165
rect 618 -173 619 -171
rect 625 -167 626 -165
rect 625 -173 626 -171
rect 632 -167 633 -165
rect 632 -173 633 -171
rect 639 -167 640 -165
rect 639 -173 640 -171
rect 646 -167 647 -165
rect 646 -173 647 -171
rect 653 -167 654 -165
rect 656 -167 657 -165
rect 656 -173 657 -171
rect 660 -167 661 -165
rect 660 -173 661 -171
rect 667 -167 668 -165
rect 667 -173 668 -171
rect 674 -167 675 -165
rect 674 -173 675 -171
rect 681 -167 682 -165
rect 681 -173 682 -171
rect 688 -167 689 -165
rect 688 -173 689 -171
rect 695 -167 696 -165
rect 695 -173 696 -171
rect 702 -167 703 -165
rect 702 -173 703 -171
rect 709 -167 710 -165
rect 709 -173 710 -171
rect 716 -167 717 -165
rect 716 -173 717 -171
rect 723 -167 724 -165
rect 723 -173 724 -171
rect 730 -167 731 -165
rect 737 -167 738 -165
rect 737 -173 738 -171
rect 744 -167 745 -165
rect 744 -173 745 -171
rect 751 -167 752 -165
rect 751 -173 752 -171
rect 758 -167 759 -165
rect 758 -173 759 -171
rect 765 -167 766 -165
rect 765 -173 766 -171
rect 772 -167 773 -165
rect 772 -173 773 -171
rect 779 -167 780 -165
rect 779 -173 780 -171
rect 786 -167 787 -165
rect 786 -173 787 -171
rect 793 -167 794 -165
rect 793 -173 794 -171
rect 800 -167 801 -165
rect 800 -173 801 -171
rect 807 -167 808 -165
rect 807 -173 808 -171
rect 814 -167 815 -165
rect 814 -173 815 -171
rect 821 -167 822 -165
rect 821 -173 822 -171
rect 828 -167 829 -165
rect 828 -173 829 -171
rect 835 -167 836 -165
rect 835 -173 836 -171
rect 842 -167 843 -165
rect 842 -173 843 -171
rect 849 -167 850 -165
rect 849 -173 850 -171
rect 856 -167 857 -165
rect 856 -173 857 -171
rect 863 -167 864 -165
rect 863 -173 864 -171
rect 870 -167 871 -165
rect 870 -173 871 -171
rect 877 -167 878 -165
rect 877 -173 878 -171
rect 898 -167 899 -165
rect 898 -173 899 -171
rect 919 -167 920 -165
rect 919 -173 920 -171
rect 940 -167 941 -165
rect 940 -173 941 -171
rect 1010 -167 1011 -165
rect 1013 -167 1014 -165
rect 1024 -167 1025 -165
rect 1024 -173 1025 -171
rect 1136 -167 1137 -165
rect 1136 -173 1137 -171
rect 1171 -167 1172 -165
rect 1171 -173 1172 -171
rect 72 -234 73 -232
rect 72 -240 73 -238
rect 79 -234 80 -232
rect 79 -240 80 -238
rect 86 -234 87 -232
rect 86 -240 87 -238
rect 93 -234 94 -232
rect 93 -240 94 -238
rect 100 -234 101 -232
rect 100 -240 101 -238
rect 107 -234 108 -232
rect 107 -240 108 -238
rect 114 -234 115 -232
rect 114 -240 115 -238
rect 121 -234 122 -232
rect 121 -240 122 -238
rect 128 -234 129 -232
rect 128 -240 129 -238
rect 135 -234 136 -232
rect 135 -240 136 -238
rect 142 -234 143 -232
rect 142 -240 143 -238
rect 149 -234 150 -232
rect 149 -240 150 -238
rect 156 -240 157 -238
rect 159 -240 160 -238
rect 163 -234 164 -232
rect 163 -240 164 -238
rect 170 -234 171 -232
rect 170 -240 171 -238
rect 177 -234 178 -232
rect 177 -240 178 -238
rect 184 -234 185 -232
rect 184 -240 185 -238
rect 191 -234 192 -232
rect 191 -240 192 -238
rect 198 -234 199 -232
rect 198 -240 199 -238
rect 205 -234 206 -232
rect 208 -234 209 -232
rect 205 -240 206 -238
rect 208 -240 209 -238
rect 212 -234 213 -232
rect 212 -240 213 -238
rect 219 -234 220 -232
rect 222 -234 223 -232
rect 219 -240 220 -238
rect 229 -234 230 -232
rect 226 -240 227 -238
rect 233 -234 234 -232
rect 236 -234 237 -232
rect 236 -240 237 -238
rect 243 -234 244 -232
rect 243 -240 244 -238
rect 247 -234 248 -232
rect 247 -240 248 -238
rect 254 -234 255 -232
rect 254 -240 255 -238
rect 257 -240 258 -238
rect 261 -234 262 -232
rect 261 -240 262 -238
rect 268 -234 269 -232
rect 268 -240 269 -238
rect 275 -234 276 -232
rect 275 -240 276 -238
rect 282 -234 283 -232
rect 282 -240 283 -238
rect 289 -234 290 -232
rect 289 -240 290 -238
rect 296 -234 297 -232
rect 296 -240 297 -238
rect 303 -234 304 -232
rect 303 -240 304 -238
rect 310 -234 311 -232
rect 310 -240 311 -238
rect 317 -234 318 -232
rect 317 -240 318 -238
rect 324 -234 325 -232
rect 324 -240 325 -238
rect 331 -234 332 -232
rect 331 -240 332 -238
rect 338 -234 339 -232
rect 338 -240 339 -238
rect 345 -234 346 -232
rect 345 -240 346 -238
rect 352 -234 353 -232
rect 352 -240 353 -238
rect 359 -234 360 -232
rect 359 -240 360 -238
rect 366 -234 367 -232
rect 366 -240 367 -238
rect 369 -240 370 -238
rect 373 -234 374 -232
rect 373 -240 374 -238
rect 380 -234 381 -232
rect 380 -240 381 -238
rect 387 -234 388 -232
rect 387 -240 388 -238
rect 394 -234 395 -232
rect 394 -240 395 -238
rect 401 -234 402 -232
rect 401 -240 402 -238
rect 408 -234 409 -232
rect 411 -240 412 -238
rect 415 -234 416 -232
rect 415 -240 416 -238
rect 422 -234 423 -232
rect 422 -240 423 -238
rect 429 -234 430 -232
rect 432 -234 433 -232
rect 429 -240 430 -238
rect 436 -234 437 -232
rect 436 -240 437 -238
rect 443 -234 444 -232
rect 446 -234 447 -232
rect 446 -240 447 -238
rect 450 -234 451 -232
rect 453 -234 454 -232
rect 450 -240 451 -238
rect 453 -240 454 -238
rect 457 -234 458 -232
rect 457 -240 458 -238
rect 464 -234 465 -232
rect 464 -240 465 -238
rect 471 -234 472 -232
rect 471 -240 472 -238
rect 478 -234 479 -232
rect 478 -240 479 -238
rect 481 -240 482 -238
rect 485 -234 486 -232
rect 485 -240 486 -238
rect 488 -240 489 -238
rect 492 -234 493 -232
rect 492 -240 493 -238
rect 499 -234 500 -232
rect 499 -240 500 -238
rect 502 -240 503 -238
rect 506 -234 507 -232
rect 506 -240 507 -238
rect 513 -234 514 -232
rect 513 -240 514 -238
rect 520 -234 521 -232
rect 520 -240 521 -238
rect 527 -234 528 -232
rect 527 -240 528 -238
rect 534 -234 535 -232
rect 534 -240 535 -238
rect 541 -234 542 -232
rect 541 -240 542 -238
rect 551 -234 552 -232
rect 551 -240 552 -238
rect 555 -234 556 -232
rect 555 -240 556 -238
rect 562 -234 563 -232
rect 562 -240 563 -238
rect 569 -234 570 -232
rect 569 -240 570 -238
rect 576 -234 577 -232
rect 576 -240 577 -238
rect 583 -234 584 -232
rect 583 -240 584 -238
rect 590 -234 591 -232
rect 590 -240 591 -238
rect 597 -234 598 -232
rect 597 -240 598 -238
rect 604 -234 605 -232
rect 604 -240 605 -238
rect 611 -234 612 -232
rect 614 -234 615 -232
rect 611 -240 612 -238
rect 618 -234 619 -232
rect 618 -240 619 -238
rect 625 -234 626 -232
rect 628 -234 629 -232
rect 628 -240 629 -238
rect 632 -234 633 -232
rect 632 -240 633 -238
rect 639 -234 640 -232
rect 639 -240 640 -238
rect 646 -234 647 -232
rect 646 -240 647 -238
rect 653 -234 654 -232
rect 653 -240 654 -238
rect 660 -234 661 -232
rect 660 -240 661 -238
rect 667 -234 668 -232
rect 667 -240 668 -238
rect 674 -234 675 -232
rect 674 -240 675 -238
rect 681 -234 682 -232
rect 681 -240 682 -238
rect 688 -234 689 -232
rect 688 -240 689 -238
rect 695 -234 696 -232
rect 695 -240 696 -238
rect 702 -234 703 -232
rect 702 -240 703 -238
rect 709 -234 710 -232
rect 709 -240 710 -238
rect 716 -234 717 -232
rect 716 -240 717 -238
rect 723 -234 724 -232
rect 723 -240 724 -238
rect 730 -234 731 -232
rect 730 -240 731 -238
rect 737 -234 738 -232
rect 737 -240 738 -238
rect 744 -234 745 -232
rect 744 -240 745 -238
rect 751 -234 752 -232
rect 754 -240 755 -238
rect 758 -234 759 -232
rect 758 -240 759 -238
rect 765 -234 766 -232
rect 765 -240 766 -238
rect 772 -234 773 -232
rect 772 -240 773 -238
rect 779 -234 780 -232
rect 779 -240 780 -238
rect 786 -234 787 -232
rect 786 -240 787 -238
rect 793 -234 794 -232
rect 793 -240 794 -238
rect 800 -234 801 -232
rect 800 -240 801 -238
rect 807 -234 808 -232
rect 807 -240 808 -238
rect 814 -234 815 -232
rect 814 -240 815 -238
rect 821 -234 822 -232
rect 821 -240 822 -238
rect 831 -234 832 -232
rect 828 -240 829 -238
rect 835 -234 836 -232
rect 835 -240 836 -238
rect 842 -234 843 -232
rect 842 -240 843 -238
rect 849 -234 850 -232
rect 849 -240 850 -238
rect 856 -234 857 -232
rect 856 -240 857 -238
rect 863 -234 864 -232
rect 863 -240 864 -238
rect 870 -234 871 -232
rect 870 -240 871 -238
rect 877 -234 878 -232
rect 877 -240 878 -238
rect 884 -234 885 -232
rect 884 -240 885 -238
rect 891 -234 892 -232
rect 891 -240 892 -238
rect 898 -234 899 -232
rect 898 -240 899 -238
rect 905 -234 906 -232
rect 905 -240 906 -238
rect 912 -234 913 -232
rect 912 -240 913 -238
rect 919 -234 920 -232
rect 919 -240 920 -238
rect 926 -234 927 -232
rect 926 -240 927 -238
rect 933 -234 934 -232
rect 933 -240 934 -238
rect 940 -234 941 -232
rect 940 -240 941 -238
rect 947 -234 948 -232
rect 947 -240 948 -238
rect 954 -234 955 -232
rect 954 -240 955 -238
rect 961 -234 962 -232
rect 961 -240 962 -238
rect 968 -234 969 -232
rect 968 -240 969 -238
rect 975 -234 976 -232
rect 975 -240 976 -238
rect 982 -234 983 -232
rect 982 -240 983 -238
rect 989 -234 990 -232
rect 989 -240 990 -238
rect 996 -234 997 -232
rect 996 -240 997 -238
rect 1003 -234 1004 -232
rect 1003 -240 1004 -238
rect 1010 -234 1011 -232
rect 1010 -240 1011 -238
rect 1017 -234 1018 -232
rect 1017 -240 1018 -238
rect 1024 -234 1025 -232
rect 1024 -240 1025 -238
rect 1038 -234 1039 -232
rect 1038 -240 1039 -238
rect 1185 -234 1186 -232
rect 1185 -240 1186 -238
rect 1325 -234 1326 -232
rect 1325 -240 1326 -238
rect 65 -317 66 -315
rect 65 -323 66 -321
rect 72 -317 73 -315
rect 72 -323 73 -321
rect 79 -317 80 -315
rect 79 -323 80 -321
rect 86 -317 87 -315
rect 86 -323 87 -321
rect 93 -317 94 -315
rect 93 -323 94 -321
rect 100 -317 101 -315
rect 100 -323 101 -321
rect 107 -317 108 -315
rect 107 -323 108 -321
rect 114 -317 115 -315
rect 114 -323 115 -321
rect 121 -317 122 -315
rect 121 -323 122 -321
rect 128 -317 129 -315
rect 128 -323 129 -321
rect 138 -317 139 -315
rect 138 -323 139 -321
rect 142 -317 143 -315
rect 145 -317 146 -315
rect 142 -323 143 -321
rect 149 -317 150 -315
rect 149 -323 150 -321
rect 156 -317 157 -315
rect 156 -323 157 -321
rect 163 -317 164 -315
rect 163 -323 164 -321
rect 170 -317 171 -315
rect 173 -317 174 -315
rect 170 -323 171 -321
rect 173 -323 174 -321
rect 177 -317 178 -315
rect 177 -323 178 -321
rect 184 -317 185 -315
rect 187 -317 188 -315
rect 184 -323 185 -321
rect 187 -323 188 -321
rect 191 -317 192 -315
rect 191 -323 192 -321
rect 198 -317 199 -315
rect 198 -323 199 -321
rect 208 -317 209 -315
rect 205 -323 206 -321
rect 208 -323 209 -321
rect 212 -317 213 -315
rect 212 -323 213 -321
rect 219 -317 220 -315
rect 219 -323 220 -321
rect 226 -317 227 -315
rect 226 -323 227 -321
rect 233 -317 234 -315
rect 233 -323 234 -321
rect 240 -317 241 -315
rect 240 -323 241 -321
rect 247 -317 248 -315
rect 247 -323 248 -321
rect 254 -317 255 -315
rect 254 -323 255 -321
rect 261 -317 262 -315
rect 261 -323 262 -321
rect 268 -317 269 -315
rect 268 -323 269 -321
rect 275 -317 276 -315
rect 275 -323 276 -321
rect 282 -317 283 -315
rect 282 -323 283 -321
rect 289 -317 290 -315
rect 289 -323 290 -321
rect 296 -317 297 -315
rect 296 -323 297 -321
rect 303 -317 304 -315
rect 303 -323 304 -321
rect 310 -317 311 -315
rect 310 -323 311 -321
rect 313 -323 314 -321
rect 317 -317 318 -315
rect 317 -323 318 -321
rect 324 -317 325 -315
rect 324 -323 325 -321
rect 331 -317 332 -315
rect 331 -323 332 -321
rect 338 -317 339 -315
rect 338 -323 339 -321
rect 345 -317 346 -315
rect 345 -323 346 -321
rect 352 -317 353 -315
rect 352 -323 353 -321
rect 359 -317 360 -315
rect 359 -323 360 -321
rect 366 -317 367 -315
rect 366 -323 367 -321
rect 373 -317 374 -315
rect 376 -317 377 -315
rect 376 -323 377 -321
rect 380 -317 381 -315
rect 383 -317 384 -315
rect 383 -323 384 -321
rect 387 -317 388 -315
rect 390 -317 391 -315
rect 387 -323 388 -321
rect 390 -323 391 -321
rect 394 -317 395 -315
rect 394 -323 395 -321
rect 401 -317 402 -315
rect 401 -323 402 -321
rect 408 -317 409 -315
rect 408 -323 409 -321
rect 415 -317 416 -315
rect 415 -323 416 -321
rect 422 -317 423 -315
rect 422 -323 423 -321
rect 429 -317 430 -315
rect 429 -323 430 -321
rect 436 -317 437 -315
rect 436 -323 437 -321
rect 443 -317 444 -315
rect 446 -317 447 -315
rect 443 -323 444 -321
rect 446 -323 447 -321
rect 450 -317 451 -315
rect 450 -323 451 -321
rect 457 -317 458 -315
rect 457 -323 458 -321
rect 464 -317 465 -315
rect 464 -323 465 -321
rect 471 -317 472 -315
rect 471 -323 472 -321
rect 478 -317 479 -315
rect 481 -323 482 -321
rect 485 -317 486 -315
rect 485 -323 486 -321
rect 492 -317 493 -315
rect 492 -323 493 -321
rect 499 -317 500 -315
rect 499 -323 500 -321
rect 506 -317 507 -315
rect 506 -323 507 -321
rect 513 -317 514 -315
rect 513 -323 514 -321
rect 520 -317 521 -315
rect 520 -323 521 -321
rect 527 -317 528 -315
rect 527 -323 528 -321
rect 534 -317 535 -315
rect 537 -317 538 -315
rect 534 -323 535 -321
rect 537 -323 538 -321
rect 541 -317 542 -315
rect 541 -323 542 -321
rect 548 -317 549 -315
rect 551 -317 552 -315
rect 548 -323 549 -321
rect 551 -323 552 -321
rect 555 -317 556 -315
rect 555 -323 556 -321
rect 562 -317 563 -315
rect 562 -323 563 -321
rect 569 -317 570 -315
rect 569 -323 570 -321
rect 576 -317 577 -315
rect 576 -323 577 -321
rect 583 -317 584 -315
rect 583 -323 584 -321
rect 590 -317 591 -315
rect 590 -323 591 -321
rect 593 -323 594 -321
rect 597 -317 598 -315
rect 600 -317 601 -315
rect 597 -323 598 -321
rect 600 -323 601 -321
rect 604 -317 605 -315
rect 607 -317 608 -315
rect 604 -323 605 -321
rect 611 -317 612 -315
rect 611 -323 612 -321
rect 618 -317 619 -315
rect 618 -323 619 -321
rect 625 -317 626 -315
rect 628 -317 629 -315
rect 625 -323 626 -321
rect 628 -323 629 -321
rect 632 -317 633 -315
rect 632 -323 633 -321
rect 639 -317 640 -315
rect 639 -323 640 -321
rect 646 -317 647 -315
rect 649 -323 650 -321
rect 653 -317 654 -315
rect 653 -323 654 -321
rect 660 -317 661 -315
rect 660 -323 661 -321
rect 667 -317 668 -315
rect 670 -317 671 -315
rect 670 -323 671 -321
rect 674 -317 675 -315
rect 674 -323 675 -321
rect 681 -317 682 -315
rect 681 -323 682 -321
rect 688 -317 689 -315
rect 688 -323 689 -321
rect 695 -317 696 -315
rect 695 -323 696 -321
rect 702 -317 703 -315
rect 702 -323 703 -321
rect 709 -317 710 -315
rect 709 -323 710 -321
rect 716 -317 717 -315
rect 716 -323 717 -321
rect 723 -317 724 -315
rect 723 -323 724 -321
rect 730 -317 731 -315
rect 730 -323 731 -321
rect 737 -317 738 -315
rect 737 -323 738 -321
rect 744 -317 745 -315
rect 747 -317 748 -315
rect 747 -323 748 -321
rect 751 -317 752 -315
rect 751 -323 752 -321
rect 758 -317 759 -315
rect 758 -323 759 -321
rect 765 -317 766 -315
rect 765 -323 766 -321
rect 772 -317 773 -315
rect 772 -323 773 -321
rect 779 -317 780 -315
rect 779 -323 780 -321
rect 786 -317 787 -315
rect 786 -323 787 -321
rect 793 -317 794 -315
rect 793 -323 794 -321
rect 800 -317 801 -315
rect 800 -323 801 -321
rect 807 -317 808 -315
rect 807 -323 808 -321
rect 814 -317 815 -315
rect 814 -323 815 -321
rect 821 -317 822 -315
rect 821 -323 822 -321
rect 828 -317 829 -315
rect 828 -323 829 -321
rect 835 -317 836 -315
rect 835 -323 836 -321
rect 842 -317 843 -315
rect 842 -323 843 -321
rect 849 -317 850 -315
rect 849 -323 850 -321
rect 856 -317 857 -315
rect 856 -323 857 -321
rect 863 -317 864 -315
rect 863 -323 864 -321
rect 870 -317 871 -315
rect 870 -323 871 -321
rect 877 -317 878 -315
rect 877 -323 878 -321
rect 884 -317 885 -315
rect 884 -323 885 -321
rect 891 -317 892 -315
rect 891 -323 892 -321
rect 898 -317 899 -315
rect 898 -323 899 -321
rect 905 -317 906 -315
rect 905 -323 906 -321
rect 912 -317 913 -315
rect 912 -323 913 -321
rect 919 -317 920 -315
rect 919 -323 920 -321
rect 926 -317 927 -315
rect 926 -323 927 -321
rect 933 -317 934 -315
rect 933 -323 934 -321
rect 940 -317 941 -315
rect 940 -323 941 -321
rect 947 -317 948 -315
rect 947 -323 948 -321
rect 954 -317 955 -315
rect 954 -323 955 -321
rect 961 -317 962 -315
rect 961 -323 962 -321
rect 968 -317 969 -315
rect 968 -323 969 -321
rect 975 -317 976 -315
rect 975 -323 976 -321
rect 982 -317 983 -315
rect 982 -323 983 -321
rect 989 -317 990 -315
rect 989 -323 990 -321
rect 996 -317 997 -315
rect 996 -323 997 -321
rect 1003 -317 1004 -315
rect 1003 -323 1004 -321
rect 1010 -317 1011 -315
rect 1010 -323 1011 -321
rect 1017 -317 1018 -315
rect 1017 -323 1018 -321
rect 1024 -317 1025 -315
rect 1024 -323 1025 -321
rect 1031 -317 1032 -315
rect 1031 -323 1032 -321
rect 1038 -317 1039 -315
rect 1038 -323 1039 -321
rect 1045 -317 1046 -315
rect 1045 -323 1046 -321
rect 1052 -317 1053 -315
rect 1052 -323 1053 -321
rect 1059 -317 1060 -315
rect 1059 -323 1060 -321
rect 1066 -317 1067 -315
rect 1066 -323 1067 -321
rect 1073 -317 1074 -315
rect 1073 -323 1074 -321
rect 1080 -317 1081 -315
rect 1080 -323 1081 -321
rect 1087 -317 1088 -315
rect 1087 -323 1088 -321
rect 1094 -317 1095 -315
rect 1094 -323 1095 -321
rect 1101 -317 1102 -315
rect 1101 -323 1102 -321
rect 1108 -317 1109 -315
rect 1108 -323 1109 -321
rect 1115 -317 1116 -315
rect 1115 -323 1116 -321
rect 1122 -317 1123 -315
rect 1122 -323 1123 -321
rect 1206 -317 1207 -315
rect 1206 -323 1207 -321
rect 1307 -317 1308 -315
rect 1307 -323 1308 -321
rect 1381 -317 1382 -315
rect 1381 -323 1382 -321
rect 1458 -317 1459 -315
rect 1458 -323 1459 -321
rect 58 -416 59 -414
rect 72 -416 73 -414
rect 72 -422 73 -420
rect 79 -416 80 -414
rect 79 -422 80 -420
rect 86 -416 87 -414
rect 86 -422 87 -420
rect 93 -416 94 -414
rect 93 -422 94 -420
rect 100 -416 101 -414
rect 100 -422 101 -420
rect 107 -416 108 -414
rect 107 -422 108 -420
rect 114 -416 115 -414
rect 114 -422 115 -420
rect 121 -416 122 -414
rect 121 -422 122 -420
rect 128 -416 129 -414
rect 128 -422 129 -420
rect 135 -416 136 -414
rect 135 -422 136 -420
rect 142 -416 143 -414
rect 142 -422 143 -420
rect 149 -416 150 -414
rect 149 -422 150 -420
rect 152 -422 153 -420
rect 156 -416 157 -414
rect 156 -422 157 -420
rect 166 -416 167 -414
rect 163 -422 164 -420
rect 166 -422 167 -420
rect 173 -416 174 -414
rect 173 -422 174 -420
rect 177 -416 178 -414
rect 177 -422 178 -420
rect 184 -416 185 -414
rect 187 -416 188 -414
rect 187 -422 188 -420
rect 194 -416 195 -414
rect 191 -422 192 -420
rect 194 -422 195 -420
rect 198 -416 199 -414
rect 198 -422 199 -420
rect 205 -416 206 -414
rect 205 -422 206 -420
rect 212 -416 213 -414
rect 212 -422 213 -420
rect 219 -416 220 -414
rect 219 -422 220 -420
rect 226 -416 227 -414
rect 226 -422 227 -420
rect 233 -416 234 -414
rect 233 -422 234 -420
rect 240 -416 241 -414
rect 240 -422 241 -420
rect 247 -416 248 -414
rect 250 -416 251 -414
rect 247 -422 248 -420
rect 250 -422 251 -420
rect 254 -416 255 -414
rect 254 -422 255 -420
rect 261 -416 262 -414
rect 261 -422 262 -420
rect 268 -416 269 -414
rect 268 -422 269 -420
rect 275 -416 276 -414
rect 275 -422 276 -420
rect 282 -416 283 -414
rect 282 -422 283 -420
rect 289 -416 290 -414
rect 289 -422 290 -420
rect 296 -416 297 -414
rect 296 -422 297 -420
rect 303 -416 304 -414
rect 303 -422 304 -420
rect 310 -416 311 -414
rect 310 -422 311 -420
rect 317 -416 318 -414
rect 317 -422 318 -420
rect 324 -416 325 -414
rect 324 -422 325 -420
rect 331 -416 332 -414
rect 331 -422 332 -420
rect 338 -416 339 -414
rect 338 -422 339 -420
rect 345 -416 346 -414
rect 345 -422 346 -420
rect 352 -416 353 -414
rect 352 -422 353 -420
rect 362 -416 363 -414
rect 359 -422 360 -420
rect 362 -422 363 -420
rect 369 -416 370 -414
rect 366 -422 367 -420
rect 369 -422 370 -420
rect 373 -416 374 -414
rect 373 -422 374 -420
rect 380 -416 381 -414
rect 383 -416 384 -414
rect 380 -422 381 -420
rect 383 -422 384 -420
rect 387 -416 388 -414
rect 387 -422 388 -420
rect 394 -416 395 -414
rect 394 -422 395 -420
rect 401 -416 402 -414
rect 401 -422 402 -420
rect 408 -416 409 -414
rect 408 -422 409 -420
rect 415 -416 416 -414
rect 418 -416 419 -414
rect 415 -422 416 -420
rect 418 -422 419 -420
rect 422 -416 423 -414
rect 422 -422 423 -420
rect 429 -416 430 -414
rect 429 -422 430 -420
rect 436 -416 437 -414
rect 436 -422 437 -420
rect 443 -416 444 -414
rect 443 -422 444 -420
rect 450 -416 451 -414
rect 450 -422 451 -420
rect 457 -416 458 -414
rect 457 -422 458 -420
rect 464 -416 465 -414
rect 464 -422 465 -420
rect 471 -416 472 -414
rect 471 -422 472 -420
rect 478 -416 479 -414
rect 478 -422 479 -420
rect 485 -416 486 -414
rect 485 -422 486 -420
rect 492 -416 493 -414
rect 495 -416 496 -414
rect 495 -422 496 -420
rect 499 -416 500 -414
rect 499 -422 500 -420
rect 506 -416 507 -414
rect 506 -422 507 -420
rect 513 -416 514 -414
rect 513 -422 514 -420
rect 520 -416 521 -414
rect 520 -422 521 -420
rect 527 -416 528 -414
rect 527 -422 528 -420
rect 534 -416 535 -414
rect 534 -422 535 -420
rect 541 -416 542 -414
rect 541 -422 542 -420
rect 544 -422 545 -420
rect 548 -416 549 -414
rect 548 -422 549 -420
rect 555 -416 556 -414
rect 555 -422 556 -420
rect 565 -416 566 -414
rect 562 -422 563 -420
rect 569 -416 570 -414
rect 572 -416 573 -414
rect 569 -422 570 -420
rect 572 -422 573 -420
rect 576 -416 577 -414
rect 576 -422 577 -420
rect 583 -416 584 -414
rect 586 -416 587 -414
rect 583 -422 584 -420
rect 586 -422 587 -420
rect 590 -416 591 -414
rect 590 -422 591 -420
rect 597 -416 598 -414
rect 597 -422 598 -420
rect 604 -416 605 -414
rect 604 -422 605 -420
rect 611 -416 612 -414
rect 611 -422 612 -420
rect 618 -416 619 -414
rect 618 -422 619 -420
rect 625 -416 626 -414
rect 625 -422 626 -420
rect 628 -422 629 -420
rect 632 -416 633 -414
rect 635 -416 636 -414
rect 632 -422 633 -420
rect 639 -416 640 -414
rect 639 -422 640 -420
rect 646 -416 647 -414
rect 646 -422 647 -420
rect 653 -416 654 -414
rect 653 -422 654 -420
rect 660 -416 661 -414
rect 660 -422 661 -420
rect 667 -416 668 -414
rect 667 -422 668 -420
rect 674 -416 675 -414
rect 674 -422 675 -420
rect 681 -416 682 -414
rect 681 -422 682 -420
rect 688 -416 689 -414
rect 691 -416 692 -414
rect 688 -422 689 -420
rect 691 -422 692 -420
rect 695 -416 696 -414
rect 695 -422 696 -420
rect 702 -416 703 -414
rect 702 -422 703 -420
rect 709 -416 710 -414
rect 709 -422 710 -420
rect 716 -416 717 -414
rect 719 -422 720 -420
rect 723 -416 724 -414
rect 723 -422 724 -420
rect 726 -422 727 -420
rect 730 -416 731 -414
rect 730 -422 731 -420
rect 737 -416 738 -414
rect 737 -422 738 -420
rect 744 -416 745 -414
rect 744 -422 745 -420
rect 751 -416 752 -414
rect 751 -422 752 -420
rect 758 -416 759 -414
rect 758 -422 759 -420
rect 765 -416 766 -414
rect 765 -422 766 -420
rect 772 -416 773 -414
rect 772 -422 773 -420
rect 779 -416 780 -414
rect 779 -422 780 -420
rect 786 -416 787 -414
rect 789 -416 790 -414
rect 789 -422 790 -420
rect 793 -416 794 -414
rect 793 -422 794 -420
rect 800 -416 801 -414
rect 800 -422 801 -420
rect 807 -416 808 -414
rect 807 -422 808 -420
rect 814 -416 815 -414
rect 814 -422 815 -420
rect 821 -416 822 -414
rect 821 -422 822 -420
rect 828 -416 829 -414
rect 828 -422 829 -420
rect 835 -416 836 -414
rect 835 -422 836 -420
rect 838 -422 839 -420
rect 842 -416 843 -414
rect 842 -422 843 -420
rect 849 -416 850 -414
rect 849 -422 850 -420
rect 856 -416 857 -414
rect 856 -422 857 -420
rect 863 -416 864 -414
rect 863 -422 864 -420
rect 870 -416 871 -414
rect 870 -422 871 -420
rect 877 -416 878 -414
rect 877 -422 878 -420
rect 884 -416 885 -414
rect 884 -422 885 -420
rect 891 -416 892 -414
rect 891 -422 892 -420
rect 898 -416 899 -414
rect 898 -422 899 -420
rect 905 -416 906 -414
rect 905 -422 906 -420
rect 912 -416 913 -414
rect 912 -422 913 -420
rect 919 -416 920 -414
rect 919 -422 920 -420
rect 926 -416 927 -414
rect 926 -422 927 -420
rect 933 -416 934 -414
rect 933 -422 934 -420
rect 940 -416 941 -414
rect 940 -422 941 -420
rect 947 -416 948 -414
rect 947 -422 948 -420
rect 954 -416 955 -414
rect 954 -422 955 -420
rect 961 -416 962 -414
rect 961 -422 962 -420
rect 968 -416 969 -414
rect 968 -422 969 -420
rect 975 -416 976 -414
rect 975 -422 976 -420
rect 982 -416 983 -414
rect 982 -422 983 -420
rect 989 -416 990 -414
rect 989 -422 990 -420
rect 996 -416 997 -414
rect 996 -422 997 -420
rect 1003 -416 1004 -414
rect 1003 -422 1004 -420
rect 1010 -416 1011 -414
rect 1010 -422 1011 -420
rect 1017 -416 1018 -414
rect 1017 -422 1018 -420
rect 1024 -416 1025 -414
rect 1024 -422 1025 -420
rect 1031 -416 1032 -414
rect 1031 -422 1032 -420
rect 1038 -416 1039 -414
rect 1038 -422 1039 -420
rect 1045 -416 1046 -414
rect 1045 -422 1046 -420
rect 1052 -416 1053 -414
rect 1052 -422 1053 -420
rect 1059 -416 1060 -414
rect 1059 -422 1060 -420
rect 1066 -416 1067 -414
rect 1066 -422 1067 -420
rect 1073 -416 1074 -414
rect 1073 -422 1074 -420
rect 1080 -416 1081 -414
rect 1080 -422 1081 -420
rect 1087 -416 1088 -414
rect 1087 -422 1088 -420
rect 1094 -416 1095 -414
rect 1094 -422 1095 -420
rect 1101 -416 1102 -414
rect 1101 -422 1102 -420
rect 1108 -416 1109 -414
rect 1108 -422 1109 -420
rect 1115 -416 1116 -414
rect 1115 -422 1116 -420
rect 1122 -416 1123 -414
rect 1122 -422 1123 -420
rect 1129 -416 1130 -414
rect 1129 -422 1130 -420
rect 1136 -416 1137 -414
rect 1136 -422 1137 -420
rect 1143 -416 1144 -414
rect 1143 -422 1144 -420
rect 1150 -416 1151 -414
rect 1150 -422 1151 -420
rect 1157 -416 1158 -414
rect 1157 -422 1158 -420
rect 1164 -416 1165 -414
rect 1164 -422 1165 -420
rect 1171 -416 1172 -414
rect 1171 -422 1172 -420
rect 1178 -416 1179 -414
rect 1178 -422 1179 -420
rect 1185 -416 1186 -414
rect 1185 -422 1186 -420
rect 1192 -416 1193 -414
rect 1192 -422 1193 -420
rect 1199 -416 1200 -414
rect 1199 -422 1200 -420
rect 1206 -416 1207 -414
rect 1206 -422 1207 -420
rect 1213 -416 1214 -414
rect 1213 -422 1214 -420
rect 1223 -416 1224 -414
rect 1220 -422 1221 -420
rect 1223 -422 1224 -420
rect 1388 -416 1389 -414
rect 1388 -422 1389 -420
rect 1409 -416 1410 -414
rect 1409 -422 1410 -420
rect 1521 -416 1522 -414
rect 1521 -422 1522 -420
rect 51 -505 52 -503
rect 51 -511 52 -509
rect 58 -505 59 -503
rect 58 -511 59 -509
rect 65 -505 66 -503
rect 65 -511 66 -509
rect 72 -505 73 -503
rect 72 -511 73 -509
rect 79 -505 80 -503
rect 79 -511 80 -509
rect 86 -505 87 -503
rect 86 -511 87 -509
rect 93 -505 94 -503
rect 93 -511 94 -509
rect 100 -505 101 -503
rect 100 -511 101 -509
rect 107 -505 108 -503
rect 107 -511 108 -509
rect 114 -505 115 -503
rect 114 -511 115 -509
rect 121 -505 122 -503
rect 124 -505 125 -503
rect 124 -511 125 -509
rect 128 -505 129 -503
rect 128 -511 129 -509
rect 135 -505 136 -503
rect 138 -505 139 -503
rect 142 -505 143 -503
rect 145 -505 146 -503
rect 142 -511 143 -509
rect 145 -511 146 -509
rect 149 -505 150 -503
rect 149 -511 150 -509
rect 156 -505 157 -503
rect 156 -511 157 -509
rect 163 -505 164 -503
rect 166 -505 167 -503
rect 163 -511 164 -509
rect 166 -511 167 -509
rect 170 -505 171 -503
rect 170 -511 171 -509
rect 177 -505 178 -503
rect 177 -511 178 -509
rect 184 -505 185 -503
rect 184 -511 185 -509
rect 191 -505 192 -503
rect 194 -505 195 -503
rect 191 -511 192 -509
rect 194 -511 195 -509
rect 198 -505 199 -503
rect 198 -511 199 -509
rect 205 -505 206 -503
rect 205 -511 206 -509
rect 212 -505 213 -503
rect 212 -511 213 -509
rect 219 -505 220 -503
rect 219 -511 220 -509
rect 226 -505 227 -503
rect 226 -511 227 -509
rect 233 -511 234 -509
rect 240 -505 241 -503
rect 240 -511 241 -509
rect 247 -505 248 -503
rect 247 -511 248 -509
rect 254 -505 255 -503
rect 257 -505 258 -503
rect 261 -505 262 -503
rect 261 -511 262 -509
rect 268 -505 269 -503
rect 268 -511 269 -509
rect 275 -505 276 -503
rect 275 -511 276 -509
rect 282 -505 283 -503
rect 282 -511 283 -509
rect 289 -505 290 -503
rect 289 -511 290 -509
rect 296 -505 297 -503
rect 299 -505 300 -503
rect 296 -511 297 -509
rect 299 -511 300 -509
rect 303 -505 304 -503
rect 303 -511 304 -509
rect 310 -505 311 -503
rect 310 -511 311 -509
rect 317 -505 318 -503
rect 317 -511 318 -509
rect 324 -505 325 -503
rect 324 -511 325 -509
rect 331 -505 332 -503
rect 331 -511 332 -509
rect 338 -505 339 -503
rect 338 -511 339 -509
rect 345 -505 346 -503
rect 345 -511 346 -509
rect 352 -505 353 -503
rect 352 -511 353 -509
rect 359 -505 360 -503
rect 359 -511 360 -509
rect 366 -505 367 -503
rect 366 -511 367 -509
rect 373 -505 374 -503
rect 373 -511 374 -509
rect 380 -505 381 -503
rect 380 -511 381 -509
rect 387 -505 388 -503
rect 390 -505 391 -503
rect 387 -511 388 -509
rect 390 -511 391 -509
rect 394 -505 395 -503
rect 394 -511 395 -509
rect 404 -505 405 -503
rect 404 -511 405 -509
rect 408 -505 409 -503
rect 408 -511 409 -509
rect 415 -505 416 -503
rect 415 -511 416 -509
rect 422 -505 423 -503
rect 425 -505 426 -503
rect 422 -511 423 -509
rect 425 -511 426 -509
rect 429 -505 430 -503
rect 429 -511 430 -509
rect 436 -505 437 -503
rect 436 -511 437 -509
rect 443 -505 444 -503
rect 443 -511 444 -509
rect 450 -505 451 -503
rect 450 -511 451 -509
rect 457 -505 458 -503
rect 457 -511 458 -509
rect 464 -505 465 -503
rect 467 -505 468 -503
rect 464 -511 465 -509
rect 467 -511 468 -509
rect 471 -505 472 -503
rect 471 -511 472 -509
rect 478 -505 479 -503
rect 478 -511 479 -509
rect 485 -505 486 -503
rect 485 -511 486 -509
rect 492 -505 493 -503
rect 492 -511 493 -509
rect 499 -505 500 -503
rect 499 -511 500 -509
rect 506 -505 507 -503
rect 506 -511 507 -509
rect 513 -505 514 -503
rect 513 -511 514 -509
rect 520 -505 521 -503
rect 520 -511 521 -509
rect 527 -505 528 -503
rect 527 -511 528 -509
rect 534 -505 535 -503
rect 534 -511 535 -509
rect 541 -505 542 -503
rect 541 -511 542 -509
rect 548 -505 549 -503
rect 551 -505 552 -503
rect 555 -505 556 -503
rect 558 -505 559 -503
rect 555 -511 556 -509
rect 562 -505 563 -503
rect 562 -511 563 -509
rect 569 -505 570 -503
rect 569 -511 570 -509
rect 576 -505 577 -503
rect 576 -511 577 -509
rect 583 -505 584 -503
rect 583 -511 584 -509
rect 590 -505 591 -503
rect 593 -505 594 -503
rect 590 -511 591 -509
rect 593 -511 594 -509
rect 597 -505 598 -503
rect 597 -511 598 -509
rect 604 -505 605 -503
rect 604 -511 605 -509
rect 611 -505 612 -503
rect 611 -511 612 -509
rect 618 -505 619 -503
rect 621 -505 622 -503
rect 618 -511 619 -509
rect 621 -511 622 -509
rect 625 -505 626 -503
rect 625 -511 626 -509
rect 632 -505 633 -503
rect 632 -511 633 -509
rect 639 -505 640 -503
rect 639 -511 640 -509
rect 649 -505 650 -503
rect 646 -511 647 -509
rect 649 -511 650 -509
rect 653 -505 654 -503
rect 656 -505 657 -503
rect 653 -511 654 -509
rect 656 -511 657 -509
rect 663 -505 664 -503
rect 660 -511 661 -509
rect 663 -511 664 -509
rect 667 -505 668 -503
rect 667 -511 668 -509
rect 674 -505 675 -503
rect 674 -511 675 -509
rect 681 -505 682 -503
rect 684 -505 685 -503
rect 684 -511 685 -509
rect 688 -505 689 -503
rect 688 -511 689 -509
rect 698 -505 699 -503
rect 695 -511 696 -509
rect 698 -511 699 -509
rect 702 -505 703 -503
rect 702 -511 703 -509
rect 709 -505 710 -503
rect 709 -511 710 -509
rect 716 -505 717 -503
rect 716 -511 717 -509
rect 723 -505 724 -503
rect 723 -511 724 -509
rect 730 -505 731 -503
rect 730 -511 731 -509
rect 737 -505 738 -503
rect 737 -511 738 -509
rect 744 -505 745 -503
rect 744 -511 745 -509
rect 751 -505 752 -503
rect 754 -505 755 -503
rect 751 -511 752 -509
rect 754 -511 755 -509
rect 758 -505 759 -503
rect 758 -511 759 -509
rect 765 -505 766 -503
rect 765 -511 766 -509
rect 772 -505 773 -503
rect 772 -511 773 -509
rect 779 -505 780 -503
rect 779 -511 780 -509
rect 786 -505 787 -503
rect 786 -511 787 -509
rect 793 -505 794 -503
rect 793 -511 794 -509
rect 800 -505 801 -503
rect 800 -511 801 -509
rect 807 -505 808 -503
rect 807 -511 808 -509
rect 814 -505 815 -503
rect 814 -511 815 -509
rect 821 -505 822 -503
rect 824 -505 825 -503
rect 821 -511 822 -509
rect 824 -511 825 -509
rect 828 -505 829 -503
rect 828 -511 829 -509
rect 835 -505 836 -503
rect 835 -511 836 -509
rect 845 -505 846 -503
rect 842 -511 843 -509
rect 845 -511 846 -509
rect 852 -505 853 -503
rect 852 -511 853 -509
rect 856 -505 857 -503
rect 856 -511 857 -509
rect 863 -505 864 -503
rect 863 -511 864 -509
rect 870 -505 871 -503
rect 870 -511 871 -509
rect 877 -505 878 -503
rect 877 -511 878 -509
rect 884 -505 885 -503
rect 884 -511 885 -509
rect 891 -505 892 -503
rect 891 -511 892 -509
rect 898 -505 899 -503
rect 898 -511 899 -509
rect 905 -505 906 -503
rect 905 -511 906 -509
rect 912 -505 913 -503
rect 912 -511 913 -509
rect 919 -505 920 -503
rect 919 -511 920 -509
rect 926 -505 927 -503
rect 926 -511 927 -509
rect 933 -505 934 -503
rect 933 -511 934 -509
rect 940 -505 941 -503
rect 940 -511 941 -509
rect 947 -505 948 -503
rect 947 -511 948 -509
rect 954 -505 955 -503
rect 954 -511 955 -509
rect 961 -505 962 -503
rect 961 -511 962 -509
rect 968 -505 969 -503
rect 968 -511 969 -509
rect 975 -505 976 -503
rect 975 -511 976 -509
rect 982 -505 983 -503
rect 982 -511 983 -509
rect 989 -505 990 -503
rect 989 -511 990 -509
rect 996 -505 997 -503
rect 996 -511 997 -509
rect 1003 -505 1004 -503
rect 1003 -511 1004 -509
rect 1010 -505 1011 -503
rect 1010 -511 1011 -509
rect 1017 -505 1018 -503
rect 1017 -511 1018 -509
rect 1024 -505 1025 -503
rect 1024 -511 1025 -509
rect 1031 -505 1032 -503
rect 1031 -511 1032 -509
rect 1038 -505 1039 -503
rect 1038 -511 1039 -509
rect 1045 -505 1046 -503
rect 1045 -511 1046 -509
rect 1052 -505 1053 -503
rect 1052 -511 1053 -509
rect 1059 -505 1060 -503
rect 1059 -511 1060 -509
rect 1066 -505 1067 -503
rect 1066 -511 1067 -509
rect 1073 -505 1074 -503
rect 1073 -511 1074 -509
rect 1080 -505 1081 -503
rect 1080 -511 1081 -509
rect 1087 -505 1088 -503
rect 1087 -511 1088 -509
rect 1094 -505 1095 -503
rect 1094 -511 1095 -509
rect 1101 -505 1102 -503
rect 1101 -511 1102 -509
rect 1108 -505 1109 -503
rect 1108 -511 1109 -509
rect 1115 -505 1116 -503
rect 1115 -511 1116 -509
rect 1122 -505 1123 -503
rect 1122 -511 1123 -509
rect 1129 -505 1130 -503
rect 1129 -511 1130 -509
rect 1136 -505 1137 -503
rect 1136 -511 1137 -509
rect 1143 -505 1144 -503
rect 1143 -511 1144 -509
rect 1150 -505 1151 -503
rect 1150 -511 1151 -509
rect 1157 -505 1158 -503
rect 1157 -511 1158 -509
rect 1164 -505 1165 -503
rect 1164 -511 1165 -509
rect 1171 -505 1172 -503
rect 1171 -511 1172 -509
rect 1178 -505 1179 -503
rect 1178 -511 1179 -509
rect 1185 -505 1186 -503
rect 1185 -511 1186 -509
rect 1192 -505 1193 -503
rect 1192 -511 1193 -509
rect 1199 -505 1200 -503
rect 1199 -511 1200 -509
rect 1206 -505 1207 -503
rect 1206 -511 1207 -509
rect 1213 -505 1214 -503
rect 1213 -511 1214 -509
rect 1223 -511 1224 -509
rect 1227 -505 1228 -503
rect 1227 -511 1228 -509
rect 1234 -505 1235 -503
rect 1234 -511 1235 -509
rect 1241 -505 1242 -503
rect 1241 -511 1242 -509
rect 1251 -505 1252 -503
rect 1251 -511 1252 -509
rect 1255 -505 1256 -503
rect 1255 -511 1256 -509
rect 1430 -505 1431 -503
rect 1430 -511 1431 -509
rect 1486 -505 1487 -503
rect 1486 -511 1487 -509
rect 1542 -505 1543 -503
rect 1542 -511 1543 -509
rect 44 -626 45 -624
rect 44 -632 45 -630
rect 51 -626 52 -624
rect 51 -632 52 -630
rect 58 -626 59 -624
rect 58 -632 59 -630
rect 65 -626 66 -624
rect 65 -632 66 -630
rect 72 -626 73 -624
rect 72 -632 73 -630
rect 79 -626 80 -624
rect 79 -632 80 -630
rect 86 -626 87 -624
rect 86 -632 87 -630
rect 93 -626 94 -624
rect 93 -632 94 -630
rect 100 -626 101 -624
rect 100 -632 101 -630
rect 107 -626 108 -624
rect 110 -626 111 -624
rect 107 -632 108 -630
rect 114 -626 115 -624
rect 114 -632 115 -630
rect 121 -626 122 -624
rect 121 -632 122 -630
rect 128 -626 129 -624
rect 128 -632 129 -630
rect 135 -626 136 -624
rect 135 -632 136 -630
rect 142 -626 143 -624
rect 142 -632 143 -630
rect 149 -626 150 -624
rect 149 -632 150 -630
rect 156 -626 157 -624
rect 156 -632 157 -630
rect 163 -626 164 -624
rect 163 -632 164 -630
rect 170 -626 171 -624
rect 170 -632 171 -630
rect 177 -626 178 -624
rect 177 -632 178 -630
rect 184 -626 185 -624
rect 184 -632 185 -630
rect 191 -626 192 -624
rect 191 -632 192 -630
rect 198 -626 199 -624
rect 198 -632 199 -630
rect 201 -632 202 -630
rect 205 -626 206 -624
rect 205 -632 206 -630
rect 212 -626 213 -624
rect 212 -632 213 -630
rect 219 -626 220 -624
rect 219 -632 220 -630
rect 226 -626 227 -624
rect 226 -632 227 -630
rect 233 -626 234 -624
rect 236 -626 237 -624
rect 233 -632 234 -630
rect 240 -626 241 -624
rect 240 -632 241 -630
rect 243 -632 244 -630
rect 247 -626 248 -624
rect 247 -632 248 -630
rect 254 -626 255 -624
rect 254 -632 255 -630
rect 261 -626 262 -624
rect 264 -626 265 -624
rect 261 -632 262 -630
rect 264 -632 265 -630
rect 268 -626 269 -624
rect 268 -632 269 -630
rect 275 -626 276 -624
rect 275 -632 276 -630
rect 282 -626 283 -624
rect 282 -632 283 -630
rect 289 -626 290 -624
rect 292 -626 293 -624
rect 289 -632 290 -630
rect 296 -626 297 -624
rect 296 -632 297 -630
rect 303 -626 304 -624
rect 303 -632 304 -630
rect 310 -626 311 -624
rect 310 -632 311 -630
rect 317 -626 318 -624
rect 317 -632 318 -630
rect 324 -626 325 -624
rect 327 -626 328 -624
rect 324 -632 325 -630
rect 327 -632 328 -630
rect 331 -626 332 -624
rect 331 -632 332 -630
rect 338 -626 339 -624
rect 338 -632 339 -630
rect 345 -626 346 -624
rect 345 -632 346 -630
rect 352 -626 353 -624
rect 355 -626 356 -624
rect 352 -632 353 -630
rect 355 -632 356 -630
rect 359 -626 360 -624
rect 359 -632 360 -630
rect 366 -626 367 -624
rect 366 -632 367 -630
rect 373 -626 374 -624
rect 373 -632 374 -630
rect 380 -626 381 -624
rect 380 -632 381 -630
rect 387 -626 388 -624
rect 390 -626 391 -624
rect 387 -632 388 -630
rect 394 -626 395 -624
rect 394 -632 395 -630
rect 401 -626 402 -624
rect 401 -632 402 -630
rect 408 -626 409 -624
rect 408 -632 409 -630
rect 415 -626 416 -624
rect 415 -632 416 -630
rect 422 -626 423 -624
rect 425 -626 426 -624
rect 422 -632 423 -630
rect 425 -632 426 -630
rect 429 -626 430 -624
rect 429 -632 430 -630
rect 436 -626 437 -624
rect 436 -632 437 -630
rect 443 -626 444 -624
rect 443 -632 444 -630
rect 450 -626 451 -624
rect 450 -632 451 -630
rect 457 -626 458 -624
rect 460 -626 461 -624
rect 457 -632 458 -630
rect 460 -632 461 -630
rect 464 -626 465 -624
rect 464 -632 465 -630
rect 471 -626 472 -624
rect 471 -632 472 -630
rect 478 -626 479 -624
rect 481 -626 482 -624
rect 478 -632 479 -630
rect 481 -632 482 -630
rect 485 -626 486 -624
rect 485 -632 486 -630
rect 492 -626 493 -624
rect 495 -626 496 -624
rect 492 -632 493 -630
rect 499 -626 500 -624
rect 499 -632 500 -630
rect 506 -626 507 -624
rect 506 -632 507 -630
rect 513 -626 514 -624
rect 513 -632 514 -630
rect 520 -626 521 -624
rect 520 -632 521 -630
rect 527 -626 528 -624
rect 527 -632 528 -630
rect 534 -626 535 -624
rect 534 -632 535 -630
rect 541 -626 542 -624
rect 541 -632 542 -630
rect 548 -626 549 -624
rect 548 -632 549 -630
rect 555 -626 556 -624
rect 555 -632 556 -630
rect 562 -626 563 -624
rect 562 -632 563 -630
rect 569 -626 570 -624
rect 569 -632 570 -630
rect 576 -626 577 -624
rect 576 -632 577 -630
rect 583 -626 584 -624
rect 583 -632 584 -630
rect 590 -626 591 -624
rect 590 -632 591 -630
rect 597 -626 598 -624
rect 597 -632 598 -630
rect 604 -626 605 -624
rect 607 -626 608 -624
rect 604 -632 605 -630
rect 607 -632 608 -630
rect 611 -626 612 -624
rect 611 -632 612 -630
rect 618 -626 619 -624
rect 618 -632 619 -630
rect 625 -626 626 -624
rect 625 -632 626 -630
rect 632 -626 633 -624
rect 632 -632 633 -630
rect 639 -626 640 -624
rect 642 -626 643 -624
rect 642 -632 643 -630
rect 646 -626 647 -624
rect 649 -626 650 -624
rect 653 -626 654 -624
rect 653 -632 654 -630
rect 660 -626 661 -624
rect 660 -632 661 -630
rect 667 -626 668 -624
rect 667 -632 668 -630
rect 674 -626 675 -624
rect 674 -632 675 -630
rect 681 -626 682 -624
rect 684 -626 685 -624
rect 681 -632 682 -630
rect 684 -632 685 -630
rect 688 -626 689 -624
rect 688 -632 689 -630
rect 695 -626 696 -624
rect 698 -626 699 -624
rect 698 -632 699 -630
rect 702 -626 703 -624
rect 702 -632 703 -630
rect 709 -626 710 -624
rect 709 -632 710 -630
rect 716 -626 717 -624
rect 716 -632 717 -630
rect 723 -626 724 -624
rect 723 -632 724 -630
rect 730 -632 731 -630
rect 733 -632 734 -630
rect 737 -626 738 -624
rect 737 -632 738 -630
rect 744 -626 745 -624
rect 747 -626 748 -624
rect 744 -632 745 -630
rect 751 -626 752 -624
rect 751 -632 752 -630
rect 758 -626 759 -624
rect 761 -626 762 -624
rect 758 -632 759 -630
rect 761 -632 762 -630
rect 765 -626 766 -624
rect 765 -632 766 -630
rect 772 -626 773 -624
rect 772 -632 773 -630
rect 779 -626 780 -624
rect 779 -632 780 -630
rect 789 -626 790 -624
rect 786 -632 787 -630
rect 789 -632 790 -630
rect 793 -626 794 -624
rect 793 -632 794 -630
rect 803 -626 804 -624
rect 800 -632 801 -630
rect 807 -626 808 -624
rect 807 -632 808 -630
rect 814 -626 815 -624
rect 814 -632 815 -630
rect 821 -626 822 -624
rect 821 -632 822 -630
rect 828 -626 829 -624
rect 828 -632 829 -630
rect 835 -626 836 -624
rect 835 -632 836 -630
rect 845 -626 846 -624
rect 842 -632 843 -630
rect 845 -632 846 -630
rect 849 -626 850 -624
rect 849 -632 850 -630
rect 856 -626 857 -624
rect 856 -632 857 -630
rect 863 -626 864 -624
rect 863 -632 864 -630
rect 870 -626 871 -624
rect 873 -626 874 -624
rect 873 -632 874 -630
rect 877 -626 878 -624
rect 877 -632 878 -630
rect 884 -626 885 -624
rect 884 -632 885 -630
rect 891 -626 892 -624
rect 891 -632 892 -630
rect 898 -626 899 -624
rect 898 -632 899 -630
rect 905 -626 906 -624
rect 905 -632 906 -630
rect 912 -626 913 -624
rect 912 -632 913 -630
rect 919 -626 920 -624
rect 919 -632 920 -630
rect 926 -626 927 -624
rect 926 -632 927 -630
rect 933 -626 934 -624
rect 933 -632 934 -630
rect 940 -626 941 -624
rect 940 -632 941 -630
rect 947 -626 948 -624
rect 947 -632 948 -630
rect 954 -626 955 -624
rect 954 -632 955 -630
rect 961 -626 962 -624
rect 961 -632 962 -630
rect 968 -626 969 -624
rect 968 -632 969 -630
rect 975 -626 976 -624
rect 975 -632 976 -630
rect 982 -626 983 -624
rect 982 -632 983 -630
rect 989 -626 990 -624
rect 989 -632 990 -630
rect 996 -626 997 -624
rect 996 -632 997 -630
rect 1003 -626 1004 -624
rect 1003 -632 1004 -630
rect 1010 -626 1011 -624
rect 1010 -632 1011 -630
rect 1017 -626 1018 -624
rect 1017 -632 1018 -630
rect 1020 -632 1021 -630
rect 1024 -626 1025 -624
rect 1024 -632 1025 -630
rect 1034 -626 1035 -624
rect 1038 -626 1039 -624
rect 1038 -632 1039 -630
rect 1045 -626 1046 -624
rect 1045 -632 1046 -630
rect 1052 -626 1053 -624
rect 1052 -632 1053 -630
rect 1059 -626 1060 -624
rect 1059 -632 1060 -630
rect 1066 -626 1067 -624
rect 1066 -632 1067 -630
rect 1073 -626 1074 -624
rect 1073 -632 1074 -630
rect 1080 -626 1081 -624
rect 1080 -632 1081 -630
rect 1087 -626 1088 -624
rect 1087 -632 1088 -630
rect 1094 -626 1095 -624
rect 1094 -632 1095 -630
rect 1101 -626 1102 -624
rect 1101 -632 1102 -630
rect 1108 -626 1109 -624
rect 1108 -632 1109 -630
rect 1115 -626 1116 -624
rect 1115 -632 1116 -630
rect 1122 -626 1123 -624
rect 1122 -632 1123 -630
rect 1129 -626 1130 -624
rect 1129 -632 1130 -630
rect 1136 -626 1137 -624
rect 1136 -632 1137 -630
rect 1143 -626 1144 -624
rect 1143 -632 1144 -630
rect 1150 -626 1151 -624
rect 1150 -632 1151 -630
rect 1157 -626 1158 -624
rect 1157 -632 1158 -630
rect 1164 -626 1165 -624
rect 1164 -632 1165 -630
rect 1171 -626 1172 -624
rect 1171 -632 1172 -630
rect 1178 -626 1179 -624
rect 1178 -632 1179 -630
rect 1185 -626 1186 -624
rect 1185 -632 1186 -630
rect 1192 -626 1193 -624
rect 1192 -632 1193 -630
rect 1199 -626 1200 -624
rect 1199 -632 1200 -630
rect 1206 -626 1207 -624
rect 1206 -632 1207 -630
rect 1213 -626 1214 -624
rect 1213 -632 1214 -630
rect 1220 -626 1221 -624
rect 1220 -632 1221 -630
rect 1227 -626 1228 -624
rect 1227 -632 1228 -630
rect 1234 -626 1235 -624
rect 1234 -632 1235 -630
rect 1241 -626 1242 -624
rect 1241 -632 1242 -630
rect 1248 -626 1249 -624
rect 1248 -632 1249 -630
rect 1255 -626 1256 -624
rect 1255 -632 1256 -630
rect 1262 -626 1263 -624
rect 1262 -632 1263 -630
rect 1269 -626 1270 -624
rect 1269 -632 1270 -630
rect 1276 -626 1277 -624
rect 1276 -632 1277 -630
rect 1283 -626 1284 -624
rect 1283 -632 1284 -630
rect 1290 -626 1291 -624
rect 1290 -632 1291 -630
rect 1297 -626 1298 -624
rect 1297 -632 1298 -630
rect 1304 -626 1305 -624
rect 1304 -632 1305 -630
rect 1311 -626 1312 -624
rect 1311 -632 1312 -630
rect 1318 -626 1319 -624
rect 1318 -632 1319 -630
rect 1325 -626 1326 -624
rect 1325 -632 1326 -630
rect 1332 -626 1333 -624
rect 1332 -632 1333 -630
rect 1339 -626 1340 -624
rect 1339 -632 1340 -630
rect 1346 -626 1347 -624
rect 1346 -632 1347 -630
rect 1353 -626 1354 -624
rect 1353 -632 1354 -630
rect 1360 -626 1361 -624
rect 1360 -632 1361 -630
rect 1367 -626 1368 -624
rect 1367 -632 1368 -630
rect 1374 -626 1375 -624
rect 1374 -632 1375 -630
rect 1381 -626 1382 -624
rect 1381 -632 1382 -630
rect 1388 -626 1389 -624
rect 1388 -632 1389 -630
rect 1395 -626 1396 -624
rect 1395 -632 1396 -630
rect 1402 -626 1403 -624
rect 1402 -632 1403 -630
rect 1409 -626 1410 -624
rect 1409 -632 1410 -630
rect 1419 -626 1420 -624
rect 1416 -632 1417 -630
rect 1419 -632 1420 -630
rect 1423 -626 1424 -624
rect 1423 -632 1424 -630
rect 1430 -626 1431 -624
rect 1430 -632 1431 -630
rect 1437 -626 1438 -624
rect 1437 -632 1438 -630
rect 1444 -626 1445 -624
rect 1444 -632 1445 -630
rect 1451 -626 1452 -624
rect 1451 -632 1452 -630
rect 1458 -626 1459 -624
rect 1458 -632 1459 -630
rect 1465 -626 1466 -624
rect 1465 -632 1466 -630
rect 1528 -626 1529 -624
rect 1528 -632 1529 -630
rect 1549 -626 1550 -624
rect 1549 -632 1550 -630
rect 1619 -626 1620 -624
rect 1619 -632 1620 -630
rect 44 -759 45 -757
rect 44 -765 45 -763
rect 51 -759 52 -757
rect 51 -765 52 -763
rect 58 -759 59 -757
rect 61 -765 62 -763
rect 68 -759 69 -757
rect 65 -765 66 -763
rect 72 -759 73 -757
rect 72 -765 73 -763
rect 79 -759 80 -757
rect 79 -765 80 -763
rect 86 -759 87 -757
rect 86 -765 87 -763
rect 93 -759 94 -757
rect 93 -765 94 -763
rect 100 -759 101 -757
rect 100 -765 101 -763
rect 107 -759 108 -757
rect 107 -765 108 -763
rect 114 -759 115 -757
rect 117 -759 118 -757
rect 117 -765 118 -763
rect 121 -759 122 -757
rect 121 -765 122 -763
rect 128 -759 129 -757
rect 128 -765 129 -763
rect 135 -759 136 -757
rect 135 -765 136 -763
rect 142 -759 143 -757
rect 142 -765 143 -763
rect 149 -759 150 -757
rect 149 -765 150 -763
rect 156 -759 157 -757
rect 159 -759 160 -757
rect 156 -765 157 -763
rect 159 -765 160 -763
rect 163 -759 164 -757
rect 163 -765 164 -763
rect 170 -759 171 -757
rect 170 -765 171 -763
rect 177 -759 178 -757
rect 177 -765 178 -763
rect 184 -759 185 -757
rect 184 -765 185 -763
rect 191 -759 192 -757
rect 191 -765 192 -763
rect 198 -759 199 -757
rect 198 -765 199 -763
rect 205 -759 206 -757
rect 205 -765 206 -763
rect 208 -765 209 -763
rect 212 -759 213 -757
rect 212 -765 213 -763
rect 219 -759 220 -757
rect 222 -759 223 -757
rect 226 -759 227 -757
rect 226 -765 227 -763
rect 233 -759 234 -757
rect 233 -765 234 -763
rect 240 -759 241 -757
rect 240 -765 241 -763
rect 247 -759 248 -757
rect 247 -765 248 -763
rect 254 -759 255 -757
rect 257 -759 258 -757
rect 261 -759 262 -757
rect 261 -765 262 -763
rect 268 -759 269 -757
rect 268 -765 269 -763
rect 275 -759 276 -757
rect 275 -765 276 -763
rect 282 -759 283 -757
rect 282 -765 283 -763
rect 289 -759 290 -757
rect 289 -765 290 -763
rect 296 -759 297 -757
rect 296 -765 297 -763
rect 303 -759 304 -757
rect 303 -765 304 -763
rect 310 -759 311 -757
rect 310 -765 311 -763
rect 317 -759 318 -757
rect 317 -765 318 -763
rect 324 -759 325 -757
rect 324 -765 325 -763
rect 331 -759 332 -757
rect 334 -759 335 -757
rect 331 -765 332 -763
rect 338 -759 339 -757
rect 338 -765 339 -763
rect 345 -759 346 -757
rect 345 -765 346 -763
rect 352 -759 353 -757
rect 352 -765 353 -763
rect 359 -759 360 -757
rect 359 -765 360 -763
rect 366 -759 367 -757
rect 366 -765 367 -763
rect 373 -759 374 -757
rect 373 -765 374 -763
rect 380 -759 381 -757
rect 380 -765 381 -763
rect 387 -759 388 -757
rect 387 -765 388 -763
rect 394 -759 395 -757
rect 394 -765 395 -763
rect 401 -759 402 -757
rect 401 -765 402 -763
rect 408 -759 409 -757
rect 408 -765 409 -763
rect 415 -759 416 -757
rect 415 -765 416 -763
rect 422 -759 423 -757
rect 422 -765 423 -763
rect 429 -759 430 -757
rect 432 -759 433 -757
rect 429 -765 430 -763
rect 432 -765 433 -763
rect 436 -759 437 -757
rect 436 -765 437 -763
rect 443 -759 444 -757
rect 443 -765 444 -763
rect 450 -759 451 -757
rect 450 -765 451 -763
rect 457 -759 458 -757
rect 457 -765 458 -763
rect 464 -759 465 -757
rect 467 -759 468 -757
rect 464 -765 465 -763
rect 471 -759 472 -757
rect 471 -765 472 -763
rect 478 -759 479 -757
rect 478 -765 479 -763
rect 485 -759 486 -757
rect 485 -765 486 -763
rect 492 -759 493 -757
rect 495 -759 496 -757
rect 492 -765 493 -763
rect 499 -759 500 -757
rect 499 -765 500 -763
rect 506 -759 507 -757
rect 506 -765 507 -763
rect 513 -759 514 -757
rect 513 -765 514 -763
rect 523 -759 524 -757
rect 520 -765 521 -763
rect 523 -765 524 -763
rect 527 -759 528 -757
rect 530 -759 531 -757
rect 527 -765 528 -763
rect 530 -765 531 -763
rect 534 -759 535 -757
rect 534 -765 535 -763
rect 541 -759 542 -757
rect 541 -765 542 -763
rect 548 -759 549 -757
rect 548 -765 549 -763
rect 555 -759 556 -757
rect 558 -759 559 -757
rect 555 -765 556 -763
rect 558 -765 559 -763
rect 562 -759 563 -757
rect 562 -765 563 -763
rect 569 -759 570 -757
rect 572 -759 573 -757
rect 572 -765 573 -763
rect 576 -759 577 -757
rect 576 -765 577 -763
rect 583 -759 584 -757
rect 583 -765 584 -763
rect 590 -759 591 -757
rect 590 -765 591 -763
rect 597 -759 598 -757
rect 597 -765 598 -763
rect 604 -759 605 -757
rect 607 -759 608 -757
rect 604 -765 605 -763
rect 607 -765 608 -763
rect 611 -759 612 -757
rect 611 -765 612 -763
rect 618 -759 619 -757
rect 618 -765 619 -763
rect 625 -759 626 -757
rect 625 -765 626 -763
rect 632 -759 633 -757
rect 635 -759 636 -757
rect 635 -765 636 -763
rect 639 -759 640 -757
rect 639 -765 640 -763
rect 646 -759 647 -757
rect 649 -759 650 -757
rect 646 -765 647 -763
rect 649 -765 650 -763
rect 653 -759 654 -757
rect 653 -765 654 -763
rect 660 -759 661 -757
rect 660 -765 661 -763
rect 667 -759 668 -757
rect 667 -765 668 -763
rect 674 -759 675 -757
rect 677 -759 678 -757
rect 674 -765 675 -763
rect 677 -765 678 -763
rect 681 -759 682 -757
rect 681 -765 682 -763
rect 691 -759 692 -757
rect 688 -765 689 -763
rect 691 -765 692 -763
rect 695 -759 696 -757
rect 695 -765 696 -763
rect 702 -759 703 -757
rect 702 -765 703 -763
rect 709 -759 710 -757
rect 709 -765 710 -763
rect 716 -759 717 -757
rect 719 -759 720 -757
rect 716 -765 717 -763
rect 719 -765 720 -763
rect 723 -759 724 -757
rect 723 -765 724 -763
rect 733 -759 734 -757
rect 730 -765 731 -763
rect 737 -759 738 -757
rect 737 -765 738 -763
rect 744 -759 745 -757
rect 744 -765 745 -763
rect 751 -759 752 -757
rect 751 -765 752 -763
rect 758 -759 759 -757
rect 758 -765 759 -763
rect 765 -759 766 -757
rect 765 -765 766 -763
rect 772 -759 773 -757
rect 772 -765 773 -763
rect 779 -759 780 -757
rect 779 -765 780 -763
rect 786 -759 787 -757
rect 786 -765 787 -763
rect 796 -759 797 -757
rect 793 -765 794 -763
rect 796 -765 797 -763
rect 800 -759 801 -757
rect 803 -759 804 -757
rect 800 -765 801 -763
rect 807 -759 808 -757
rect 807 -765 808 -763
rect 814 -759 815 -757
rect 814 -765 815 -763
rect 821 -759 822 -757
rect 821 -765 822 -763
rect 828 -759 829 -757
rect 831 -759 832 -757
rect 828 -765 829 -763
rect 831 -765 832 -763
rect 835 -759 836 -757
rect 838 -759 839 -757
rect 835 -765 836 -763
rect 838 -765 839 -763
rect 842 -759 843 -757
rect 842 -765 843 -763
rect 849 -759 850 -757
rect 849 -765 850 -763
rect 856 -759 857 -757
rect 856 -765 857 -763
rect 863 -759 864 -757
rect 863 -765 864 -763
rect 870 -759 871 -757
rect 870 -765 871 -763
rect 873 -765 874 -763
rect 877 -759 878 -757
rect 877 -765 878 -763
rect 884 -759 885 -757
rect 884 -765 885 -763
rect 891 -759 892 -757
rect 891 -765 892 -763
rect 898 -759 899 -757
rect 898 -765 899 -763
rect 905 -759 906 -757
rect 908 -759 909 -757
rect 905 -765 906 -763
rect 908 -765 909 -763
rect 912 -759 913 -757
rect 912 -765 913 -763
rect 919 -759 920 -757
rect 919 -765 920 -763
rect 929 -759 930 -757
rect 926 -765 927 -763
rect 929 -765 930 -763
rect 933 -759 934 -757
rect 933 -765 934 -763
rect 940 -759 941 -757
rect 940 -765 941 -763
rect 947 -759 948 -757
rect 947 -765 948 -763
rect 954 -759 955 -757
rect 954 -765 955 -763
rect 961 -759 962 -757
rect 961 -765 962 -763
rect 968 -759 969 -757
rect 968 -765 969 -763
rect 975 -759 976 -757
rect 975 -765 976 -763
rect 982 -759 983 -757
rect 982 -765 983 -763
rect 989 -759 990 -757
rect 989 -765 990 -763
rect 996 -759 997 -757
rect 996 -765 997 -763
rect 1003 -759 1004 -757
rect 1003 -765 1004 -763
rect 1010 -759 1011 -757
rect 1010 -765 1011 -763
rect 1017 -759 1018 -757
rect 1017 -765 1018 -763
rect 1024 -759 1025 -757
rect 1024 -765 1025 -763
rect 1027 -765 1028 -763
rect 1031 -759 1032 -757
rect 1031 -765 1032 -763
rect 1038 -759 1039 -757
rect 1038 -765 1039 -763
rect 1045 -759 1046 -757
rect 1045 -765 1046 -763
rect 1052 -759 1053 -757
rect 1052 -765 1053 -763
rect 1059 -759 1060 -757
rect 1059 -765 1060 -763
rect 1066 -759 1067 -757
rect 1066 -765 1067 -763
rect 1073 -759 1074 -757
rect 1073 -765 1074 -763
rect 1080 -759 1081 -757
rect 1080 -765 1081 -763
rect 1087 -759 1088 -757
rect 1087 -765 1088 -763
rect 1094 -759 1095 -757
rect 1094 -765 1095 -763
rect 1101 -759 1102 -757
rect 1101 -765 1102 -763
rect 1108 -759 1109 -757
rect 1108 -765 1109 -763
rect 1115 -759 1116 -757
rect 1115 -765 1116 -763
rect 1122 -759 1123 -757
rect 1122 -765 1123 -763
rect 1129 -759 1130 -757
rect 1129 -765 1130 -763
rect 1136 -759 1137 -757
rect 1136 -765 1137 -763
rect 1143 -759 1144 -757
rect 1143 -765 1144 -763
rect 1150 -759 1151 -757
rect 1150 -765 1151 -763
rect 1157 -759 1158 -757
rect 1157 -765 1158 -763
rect 1164 -759 1165 -757
rect 1164 -765 1165 -763
rect 1171 -759 1172 -757
rect 1171 -765 1172 -763
rect 1178 -759 1179 -757
rect 1178 -765 1179 -763
rect 1185 -759 1186 -757
rect 1185 -765 1186 -763
rect 1192 -759 1193 -757
rect 1192 -765 1193 -763
rect 1199 -759 1200 -757
rect 1199 -765 1200 -763
rect 1206 -759 1207 -757
rect 1206 -765 1207 -763
rect 1213 -759 1214 -757
rect 1213 -765 1214 -763
rect 1220 -759 1221 -757
rect 1220 -765 1221 -763
rect 1227 -759 1228 -757
rect 1227 -765 1228 -763
rect 1234 -759 1235 -757
rect 1234 -765 1235 -763
rect 1241 -759 1242 -757
rect 1241 -765 1242 -763
rect 1248 -759 1249 -757
rect 1248 -765 1249 -763
rect 1255 -759 1256 -757
rect 1255 -765 1256 -763
rect 1262 -759 1263 -757
rect 1262 -765 1263 -763
rect 1269 -759 1270 -757
rect 1269 -765 1270 -763
rect 1276 -759 1277 -757
rect 1276 -765 1277 -763
rect 1283 -759 1284 -757
rect 1283 -765 1284 -763
rect 1290 -759 1291 -757
rect 1290 -765 1291 -763
rect 1297 -759 1298 -757
rect 1297 -765 1298 -763
rect 1304 -759 1305 -757
rect 1304 -765 1305 -763
rect 1311 -759 1312 -757
rect 1311 -765 1312 -763
rect 1318 -759 1319 -757
rect 1318 -765 1319 -763
rect 1325 -759 1326 -757
rect 1325 -765 1326 -763
rect 1332 -759 1333 -757
rect 1332 -765 1333 -763
rect 1339 -759 1340 -757
rect 1339 -765 1340 -763
rect 1346 -759 1347 -757
rect 1346 -765 1347 -763
rect 1353 -759 1354 -757
rect 1353 -765 1354 -763
rect 1360 -759 1361 -757
rect 1360 -765 1361 -763
rect 1367 -759 1368 -757
rect 1367 -765 1368 -763
rect 1374 -759 1375 -757
rect 1374 -765 1375 -763
rect 1381 -759 1382 -757
rect 1381 -765 1382 -763
rect 1388 -759 1389 -757
rect 1388 -765 1389 -763
rect 1395 -759 1396 -757
rect 1395 -765 1396 -763
rect 1402 -759 1403 -757
rect 1402 -765 1403 -763
rect 1409 -759 1410 -757
rect 1409 -765 1410 -763
rect 1416 -759 1417 -757
rect 1416 -765 1417 -763
rect 1423 -759 1424 -757
rect 1423 -765 1424 -763
rect 1430 -759 1431 -757
rect 1430 -765 1431 -763
rect 1437 -759 1438 -757
rect 1437 -765 1438 -763
rect 1444 -759 1445 -757
rect 1444 -765 1445 -763
rect 1451 -759 1452 -757
rect 1451 -765 1452 -763
rect 1458 -759 1459 -757
rect 1458 -765 1459 -763
rect 1465 -759 1466 -757
rect 1465 -765 1466 -763
rect 1472 -759 1473 -757
rect 1472 -765 1473 -763
rect 1479 -759 1480 -757
rect 1479 -765 1480 -763
rect 1486 -759 1487 -757
rect 1486 -765 1487 -763
rect 1528 -759 1529 -757
rect 1528 -765 1529 -763
rect 1549 -759 1550 -757
rect 1549 -765 1550 -763
rect 1556 -759 1557 -757
rect 1556 -765 1557 -763
rect 1696 -759 1697 -757
rect 1696 -765 1697 -763
rect 37 -872 38 -870
rect 37 -878 38 -876
rect 44 -872 45 -870
rect 44 -878 45 -876
rect 51 -872 52 -870
rect 51 -878 52 -876
rect 58 -872 59 -870
rect 58 -878 59 -876
rect 65 -872 66 -870
rect 65 -878 66 -876
rect 72 -872 73 -870
rect 72 -878 73 -876
rect 79 -872 80 -870
rect 79 -878 80 -876
rect 86 -872 87 -870
rect 86 -878 87 -876
rect 93 -872 94 -870
rect 93 -878 94 -876
rect 100 -872 101 -870
rect 100 -878 101 -876
rect 107 -872 108 -870
rect 107 -878 108 -876
rect 110 -878 111 -876
rect 114 -872 115 -870
rect 114 -878 115 -876
rect 121 -872 122 -870
rect 124 -872 125 -870
rect 121 -878 122 -876
rect 124 -878 125 -876
rect 128 -872 129 -870
rect 128 -878 129 -876
rect 135 -872 136 -870
rect 135 -878 136 -876
rect 142 -872 143 -870
rect 142 -878 143 -876
rect 149 -872 150 -870
rect 152 -872 153 -870
rect 149 -878 150 -876
rect 156 -872 157 -870
rect 156 -878 157 -876
rect 163 -872 164 -870
rect 166 -872 167 -870
rect 163 -878 164 -876
rect 166 -878 167 -876
rect 170 -872 171 -870
rect 170 -878 171 -876
rect 177 -872 178 -870
rect 177 -878 178 -876
rect 184 -872 185 -870
rect 187 -872 188 -870
rect 184 -878 185 -876
rect 191 -872 192 -870
rect 191 -878 192 -876
rect 198 -872 199 -870
rect 198 -878 199 -876
rect 205 -872 206 -870
rect 208 -872 209 -870
rect 205 -878 206 -876
rect 208 -878 209 -876
rect 212 -872 213 -870
rect 212 -878 213 -876
rect 222 -878 223 -876
rect 226 -872 227 -870
rect 226 -878 227 -876
rect 233 -872 234 -870
rect 233 -878 234 -876
rect 240 -872 241 -870
rect 240 -878 241 -876
rect 247 -872 248 -870
rect 247 -878 248 -876
rect 254 -872 255 -870
rect 254 -878 255 -876
rect 257 -878 258 -876
rect 261 -872 262 -870
rect 261 -878 262 -876
rect 268 -872 269 -870
rect 268 -878 269 -876
rect 275 -872 276 -870
rect 275 -878 276 -876
rect 282 -872 283 -870
rect 282 -878 283 -876
rect 289 -872 290 -870
rect 289 -878 290 -876
rect 296 -872 297 -870
rect 296 -878 297 -876
rect 303 -872 304 -870
rect 303 -878 304 -876
rect 310 -872 311 -870
rect 310 -878 311 -876
rect 317 -872 318 -870
rect 317 -878 318 -876
rect 324 -872 325 -870
rect 331 -872 332 -870
rect 331 -878 332 -876
rect 338 -872 339 -870
rect 338 -878 339 -876
rect 345 -872 346 -870
rect 345 -878 346 -876
rect 352 -872 353 -870
rect 352 -878 353 -876
rect 359 -872 360 -870
rect 359 -878 360 -876
rect 366 -872 367 -870
rect 366 -878 367 -876
rect 373 -872 374 -870
rect 373 -878 374 -876
rect 380 -872 381 -870
rect 380 -878 381 -876
rect 387 -872 388 -870
rect 387 -878 388 -876
rect 394 -872 395 -870
rect 394 -878 395 -876
rect 401 -872 402 -870
rect 401 -878 402 -876
rect 411 -872 412 -870
rect 408 -878 409 -876
rect 411 -878 412 -876
rect 415 -872 416 -870
rect 415 -878 416 -876
rect 422 -872 423 -870
rect 422 -878 423 -876
rect 429 -872 430 -870
rect 429 -878 430 -876
rect 436 -872 437 -870
rect 436 -878 437 -876
rect 443 -872 444 -870
rect 443 -878 444 -876
rect 450 -872 451 -870
rect 450 -878 451 -876
rect 457 -872 458 -870
rect 457 -878 458 -876
rect 464 -872 465 -870
rect 464 -878 465 -876
rect 471 -872 472 -870
rect 471 -878 472 -876
rect 478 -872 479 -870
rect 478 -878 479 -876
rect 485 -872 486 -870
rect 485 -878 486 -876
rect 492 -872 493 -870
rect 492 -878 493 -876
rect 499 -872 500 -870
rect 499 -878 500 -876
rect 502 -878 503 -876
rect 506 -872 507 -870
rect 509 -872 510 -870
rect 506 -878 507 -876
rect 509 -878 510 -876
rect 513 -872 514 -870
rect 513 -878 514 -876
rect 520 -872 521 -870
rect 523 -872 524 -870
rect 520 -878 521 -876
rect 523 -878 524 -876
rect 527 -872 528 -870
rect 530 -872 531 -870
rect 527 -878 528 -876
rect 530 -878 531 -876
rect 534 -872 535 -870
rect 534 -878 535 -876
rect 537 -878 538 -876
rect 541 -872 542 -870
rect 541 -878 542 -876
rect 548 -872 549 -870
rect 551 -872 552 -870
rect 548 -878 549 -876
rect 551 -878 552 -876
rect 555 -872 556 -870
rect 555 -878 556 -876
rect 562 -872 563 -870
rect 562 -878 563 -876
rect 569 -872 570 -870
rect 569 -878 570 -876
rect 576 -872 577 -870
rect 576 -878 577 -876
rect 583 -872 584 -870
rect 583 -878 584 -876
rect 590 -872 591 -870
rect 590 -878 591 -876
rect 597 -872 598 -870
rect 597 -878 598 -876
rect 604 -872 605 -870
rect 604 -878 605 -876
rect 611 -872 612 -870
rect 611 -878 612 -876
rect 618 -872 619 -870
rect 618 -878 619 -876
rect 625 -878 626 -876
rect 628 -878 629 -876
rect 632 -872 633 -870
rect 632 -878 633 -876
rect 639 -872 640 -870
rect 639 -878 640 -876
rect 646 -872 647 -870
rect 649 -872 650 -870
rect 646 -878 647 -876
rect 649 -878 650 -876
rect 653 -872 654 -870
rect 653 -878 654 -876
rect 660 -872 661 -870
rect 660 -878 661 -876
rect 667 -872 668 -870
rect 667 -878 668 -876
rect 670 -878 671 -876
rect 674 -872 675 -870
rect 674 -878 675 -876
rect 677 -878 678 -876
rect 681 -872 682 -870
rect 684 -872 685 -870
rect 681 -878 682 -876
rect 684 -878 685 -876
rect 688 -872 689 -870
rect 688 -878 689 -876
rect 695 -872 696 -870
rect 695 -878 696 -876
rect 702 -872 703 -870
rect 702 -878 703 -876
rect 709 -872 710 -870
rect 709 -878 710 -876
rect 716 -872 717 -870
rect 716 -878 717 -876
rect 723 -872 724 -870
rect 723 -878 724 -876
rect 730 -872 731 -870
rect 730 -878 731 -876
rect 737 -872 738 -870
rect 737 -878 738 -876
rect 744 -872 745 -870
rect 744 -878 745 -876
rect 751 -872 752 -870
rect 751 -878 752 -876
rect 758 -872 759 -870
rect 758 -878 759 -876
rect 765 -872 766 -870
rect 765 -878 766 -876
rect 772 -872 773 -870
rect 772 -878 773 -876
rect 779 -872 780 -870
rect 782 -872 783 -870
rect 782 -878 783 -876
rect 786 -872 787 -870
rect 786 -878 787 -876
rect 793 -872 794 -870
rect 793 -878 794 -876
rect 800 -872 801 -870
rect 800 -878 801 -876
rect 807 -872 808 -870
rect 807 -878 808 -876
rect 814 -872 815 -870
rect 814 -878 815 -876
rect 821 -872 822 -870
rect 821 -878 822 -876
rect 828 -872 829 -870
rect 831 -872 832 -870
rect 828 -878 829 -876
rect 831 -878 832 -876
rect 835 -872 836 -870
rect 838 -872 839 -870
rect 835 -878 836 -876
rect 838 -878 839 -876
rect 842 -872 843 -870
rect 842 -878 843 -876
rect 849 -872 850 -870
rect 849 -878 850 -876
rect 856 -872 857 -870
rect 856 -878 857 -876
rect 863 -872 864 -870
rect 863 -878 864 -876
rect 870 -872 871 -870
rect 873 -872 874 -870
rect 870 -878 871 -876
rect 873 -878 874 -876
rect 877 -872 878 -870
rect 880 -872 881 -870
rect 877 -878 878 -876
rect 880 -878 881 -876
rect 884 -872 885 -870
rect 884 -878 885 -876
rect 891 -872 892 -870
rect 891 -878 892 -876
rect 898 -872 899 -870
rect 898 -878 899 -876
rect 905 -872 906 -870
rect 905 -878 906 -876
rect 912 -872 913 -870
rect 912 -878 913 -876
rect 919 -872 920 -870
rect 922 -872 923 -870
rect 919 -878 920 -876
rect 922 -878 923 -876
rect 926 -872 927 -870
rect 926 -878 927 -876
rect 929 -878 930 -876
rect 933 -872 934 -870
rect 933 -878 934 -876
rect 940 -872 941 -870
rect 940 -878 941 -876
rect 947 -872 948 -870
rect 947 -878 948 -876
rect 954 -872 955 -870
rect 954 -878 955 -876
rect 961 -872 962 -870
rect 964 -872 965 -870
rect 964 -878 965 -876
rect 968 -872 969 -870
rect 968 -878 969 -876
rect 975 -872 976 -870
rect 975 -878 976 -876
rect 982 -872 983 -870
rect 982 -878 983 -876
rect 989 -872 990 -870
rect 989 -878 990 -876
rect 996 -872 997 -870
rect 996 -878 997 -876
rect 1003 -872 1004 -870
rect 1003 -878 1004 -876
rect 1010 -872 1011 -870
rect 1010 -878 1011 -876
rect 1017 -872 1018 -870
rect 1017 -878 1018 -876
rect 1024 -872 1025 -870
rect 1024 -878 1025 -876
rect 1031 -872 1032 -870
rect 1031 -878 1032 -876
rect 1038 -872 1039 -870
rect 1038 -878 1039 -876
rect 1045 -872 1046 -870
rect 1045 -878 1046 -876
rect 1052 -872 1053 -870
rect 1052 -878 1053 -876
rect 1059 -872 1060 -870
rect 1059 -878 1060 -876
rect 1066 -872 1067 -870
rect 1066 -878 1067 -876
rect 1069 -878 1070 -876
rect 1073 -872 1074 -870
rect 1073 -878 1074 -876
rect 1080 -872 1081 -870
rect 1080 -878 1081 -876
rect 1087 -872 1088 -870
rect 1087 -878 1088 -876
rect 1094 -872 1095 -870
rect 1094 -878 1095 -876
rect 1101 -872 1102 -870
rect 1101 -878 1102 -876
rect 1108 -872 1109 -870
rect 1108 -878 1109 -876
rect 1115 -872 1116 -870
rect 1115 -878 1116 -876
rect 1122 -872 1123 -870
rect 1122 -878 1123 -876
rect 1129 -872 1130 -870
rect 1129 -878 1130 -876
rect 1136 -872 1137 -870
rect 1136 -878 1137 -876
rect 1143 -872 1144 -870
rect 1143 -878 1144 -876
rect 1150 -872 1151 -870
rect 1150 -878 1151 -876
rect 1157 -872 1158 -870
rect 1157 -878 1158 -876
rect 1164 -872 1165 -870
rect 1164 -878 1165 -876
rect 1171 -872 1172 -870
rect 1171 -878 1172 -876
rect 1178 -872 1179 -870
rect 1178 -878 1179 -876
rect 1185 -872 1186 -870
rect 1185 -878 1186 -876
rect 1192 -872 1193 -870
rect 1192 -878 1193 -876
rect 1199 -872 1200 -870
rect 1199 -878 1200 -876
rect 1206 -872 1207 -870
rect 1206 -878 1207 -876
rect 1213 -872 1214 -870
rect 1213 -878 1214 -876
rect 1220 -872 1221 -870
rect 1220 -878 1221 -876
rect 1227 -872 1228 -870
rect 1227 -878 1228 -876
rect 1234 -872 1235 -870
rect 1234 -878 1235 -876
rect 1241 -872 1242 -870
rect 1241 -878 1242 -876
rect 1248 -872 1249 -870
rect 1248 -878 1249 -876
rect 1255 -872 1256 -870
rect 1255 -878 1256 -876
rect 1262 -872 1263 -870
rect 1262 -878 1263 -876
rect 1269 -872 1270 -870
rect 1269 -878 1270 -876
rect 1276 -872 1277 -870
rect 1276 -878 1277 -876
rect 1283 -872 1284 -870
rect 1283 -878 1284 -876
rect 1290 -872 1291 -870
rect 1290 -878 1291 -876
rect 1297 -872 1298 -870
rect 1297 -878 1298 -876
rect 1304 -872 1305 -870
rect 1304 -878 1305 -876
rect 1311 -872 1312 -870
rect 1311 -878 1312 -876
rect 1318 -872 1319 -870
rect 1318 -878 1319 -876
rect 1325 -872 1326 -870
rect 1325 -878 1326 -876
rect 1332 -872 1333 -870
rect 1332 -878 1333 -876
rect 1339 -872 1340 -870
rect 1339 -878 1340 -876
rect 1346 -872 1347 -870
rect 1346 -878 1347 -876
rect 1353 -872 1354 -870
rect 1353 -878 1354 -876
rect 1360 -872 1361 -870
rect 1360 -878 1361 -876
rect 1367 -872 1368 -870
rect 1367 -878 1368 -876
rect 1374 -872 1375 -870
rect 1374 -878 1375 -876
rect 1381 -872 1382 -870
rect 1381 -878 1382 -876
rect 1388 -872 1389 -870
rect 1388 -878 1389 -876
rect 1395 -872 1396 -870
rect 1395 -878 1396 -876
rect 1402 -872 1403 -870
rect 1402 -878 1403 -876
rect 1409 -872 1410 -870
rect 1409 -878 1410 -876
rect 1416 -872 1417 -870
rect 1416 -878 1417 -876
rect 1423 -872 1424 -870
rect 1423 -878 1424 -876
rect 1430 -872 1431 -870
rect 1430 -878 1431 -876
rect 1437 -872 1438 -870
rect 1437 -878 1438 -876
rect 1444 -872 1445 -870
rect 1444 -878 1445 -876
rect 1451 -872 1452 -870
rect 1451 -878 1452 -876
rect 1458 -872 1459 -870
rect 1458 -878 1459 -876
rect 1465 -872 1466 -870
rect 1465 -878 1466 -876
rect 1472 -872 1473 -870
rect 1472 -878 1473 -876
rect 1479 -872 1480 -870
rect 1479 -878 1480 -876
rect 1486 -872 1487 -870
rect 1486 -878 1487 -876
rect 1493 -872 1494 -870
rect 1493 -878 1494 -876
rect 1500 -872 1501 -870
rect 1500 -878 1501 -876
rect 1507 -872 1508 -870
rect 1507 -878 1508 -876
rect 1514 -872 1515 -870
rect 1514 -878 1515 -876
rect 1521 -872 1522 -870
rect 1521 -878 1522 -876
rect 1528 -872 1529 -870
rect 1528 -878 1529 -876
rect 1535 -872 1536 -870
rect 1535 -878 1536 -876
rect 1542 -872 1543 -870
rect 1542 -878 1543 -876
rect 1549 -872 1550 -870
rect 1549 -878 1550 -876
rect 1556 -872 1557 -870
rect 1559 -872 1560 -870
rect 1556 -878 1557 -876
rect 1563 -878 1564 -876
rect 1570 -872 1571 -870
rect 1570 -878 1571 -876
rect 1577 -872 1578 -870
rect 1577 -878 1578 -876
rect 1584 -872 1585 -870
rect 1584 -878 1585 -876
rect 1724 -872 1725 -870
rect 1724 -878 1725 -876
rect 30 -999 31 -997
rect 30 -1005 31 -1003
rect 37 -999 38 -997
rect 37 -1005 38 -1003
rect 44 -999 45 -997
rect 44 -1005 45 -1003
rect 51 -999 52 -997
rect 51 -1005 52 -1003
rect 58 -999 59 -997
rect 58 -1005 59 -1003
rect 65 -999 66 -997
rect 72 -999 73 -997
rect 72 -1005 73 -1003
rect 79 -999 80 -997
rect 82 -999 83 -997
rect 79 -1005 80 -1003
rect 82 -1005 83 -1003
rect 86 -999 87 -997
rect 86 -1005 87 -1003
rect 93 -999 94 -997
rect 93 -1005 94 -1003
rect 100 -999 101 -997
rect 100 -1005 101 -1003
rect 107 -999 108 -997
rect 107 -1005 108 -1003
rect 114 -999 115 -997
rect 114 -1005 115 -1003
rect 121 -999 122 -997
rect 121 -1005 122 -1003
rect 128 -999 129 -997
rect 128 -1005 129 -1003
rect 131 -1005 132 -1003
rect 135 -999 136 -997
rect 138 -999 139 -997
rect 138 -1005 139 -1003
rect 142 -999 143 -997
rect 142 -1005 143 -1003
rect 149 -999 150 -997
rect 152 -999 153 -997
rect 156 -999 157 -997
rect 156 -1005 157 -1003
rect 163 -999 164 -997
rect 163 -1005 164 -1003
rect 170 -999 171 -997
rect 170 -1005 171 -1003
rect 177 -999 178 -997
rect 177 -1005 178 -1003
rect 184 -999 185 -997
rect 184 -1005 185 -1003
rect 191 -999 192 -997
rect 191 -1005 192 -1003
rect 198 -999 199 -997
rect 198 -1005 199 -1003
rect 205 -999 206 -997
rect 205 -1005 206 -1003
rect 212 -999 213 -997
rect 212 -1005 213 -1003
rect 219 -999 220 -997
rect 219 -1005 220 -1003
rect 226 -999 227 -997
rect 226 -1005 227 -1003
rect 233 -999 234 -997
rect 233 -1005 234 -1003
rect 240 -999 241 -997
rect 250 -999 251 -997
rect 250 -1005 251 -1003
rect 254 -999 255 -997
rect 254 -1005 255 -1003
rect 261 -999 262 -997
rect 261 -1005 262 -1003
rect 268 -999 269 -997
rect 268 -1005 269 -1003
rect 275 -999 276 -997
rect 275 -1005 276 -1003
rect 282 -999 283 -997
rect 282 -1005 283 -1003
rect 289 -999 290 -997
rect 289 -1005 290 -1003
rect 296 -999 297 -997
rect 296 -1005 297 -1003
rect 303 -999 304 -997
rect 303 -1005 304 -1003
rect 310 -999 311 -997
rect 310 -1005 311 -1003
rect 317 -999 318 -997
rect 317 -1005 318 -1003
rect 324 -1005 325 -1003
rect 331 -999 332 -997
rect 331 -1005 332 -1003
rect 338 -999 339 -997
rect 338 -1005 339 -1003
rect 345 -999 346 -997
rect 345 -1005 346 -1003
rect 352 -999 353 -997
rect 352 -1005 353 -1003
rect 359 -999 360 -997
rect 359 -1005 360 -1003
rect 366 -999 367 -997
rect 366 -1005 367 -1003
rect 373 -999 374 -997
rect 373 -1005 374 -1003
rect 380 -999 381 -997
rect 380 -1005 381 -1003
rect 387 -999 388 -997
rect 387 -1005 388 -1003
rect 394 -999 395 -997
rect 394 -1005 395 -1003
rect 401 -999 402 -997
rect 401 -1005 402 -1003
rect 408 -999 409 -997
rect 408 -1005 409 -1003
rect 415 -999 416 -997
rect 415 -1005 416 -1003
rect 422 -999 423 -997
rect 425 -999 426 -997
rect 422 -1005 423 -1003
rect 425 -1005 426 -1003
rect 429 -999 430 -997
rect 429 -1005 430 -1003
rect 436 -999 437 -997
rect 436 -1005 437 -1003
rect 443 -999 444 -997
rect 446 -999 447 -997
rect 443 -1005 444 -1003
rect 446 -1005 447 -1003
rect 450 -999 451 -997
rect 450 -1005 451 -1003
rect 457 -999 458 -997
rect 457 -1005 458 -1003
rect 464 -999 465 -997
rect 464 -1005 465 -1003
rect 471 -999 472 -997
rect 471 -1005 472 -1003
rect 478 -999 479 -997
rect 478 -1005 479 -1003
rect 485 -999 486 -997
rect 485 -1005 486 -1003
rect 492 -999 493 -997
rect 492 -1005 493 -1003
rect 499 -999 500 -997
rect 502 -999 503 -997
rect 499 -1005 500 -1003
rect 502 -1005 503 -1003
rect 506 -999 507 -997
rect 509 -999 510 -997
rect 506 -1005 507 -1003
rect 509 -1005 510 -1003
rect 513 -999 514 -997
rect 513 -1005 514 -1003
rect 520 -999 521 -997
rect 520 -1005 521 -1003
rect 527 -999 528 -997
rect 527 -1005 528 -1003
rect 534 -999 535 -997
rect 534 -1005 535 -1003
rect 541 -999 542 -997
rect 541 -1005 542 -1003
rect 548 -999 549 -997
rect 548 -1005 549 -1003
rect 555 -999 556 -997
rect 555 -1005 556 -1003
rect 562 -999 563 -997
rect 562 -1005 563 -1003
rect 569 -999 570 -997
rect 569 -1005 570 -1003
rect 576 -999 577 -997
rect 576 -1005 577 -1003
rect 583 -999 584 -997
rect 586 -999 587 -997
rect 583 -1005 584 -1003
rect 586 -1005 587 -1003
rect 590 -999 591 -997
rect 590 -1005 591 -1003
rect 597 -999 598 -997
rect 597 -1005 598 -1003
rect 604 -999 605 -997
rect 604 -1005 605 -1003
rect 611 -999 612 -997
rect 611 -1005 612 -1003
rect 618 -1005 619 -1003
rect 621 -1005 622 -1003
rect 625 -999 626 -997
rect 625 -1005 626 -1003
rect 632 -999 633 -997
rect 632 -1005 633 -1003
rect 639 -999 640 -997
rect 642 -999 643 -997
rect 639 -1005 640 -1003
rect 646 -999 647 -997
rect 649 -999 650 -997
rect 646 -1005 647 -1003
rect 649 -1005 650 -1003
rect 653 -999 654 -997
rect 656 -999 657 -997
rect 653 -1005 654 -1003
rect 656 -1005 657 -1003
rect 660 -999 661 -997
rect 660 -1005 661 -1003
rect 667 -999 668 -997
rect 667 -1005 668 -1003
rect 674 -999 675 -997
rect 674 -1005 675 -1003
rect 681 -999 682 -997
rect 684 -999 685 -997
rect 681 -1005 682 -1003
rect 684 -1005 685 -1003
rect 688 -999 689 -997
rect 691 -1005 692 -1003
rect 695 -999 696 -997
rect 698 -999 699 -997
rect 695 -1005 696 -1003
rect 698 -1005 699 -1003
rect 702 -999 703 -997
rect 702 -1005 703 -1003
rect 709 -999 710 -997
rect 709 -1005 710 -1003
rect 716 -999 717 -997
rect 716 -1005 717 -1003
rect 723 -999 724 -997
rect 723 -1005 724 -1003
rect 730 -999 731 -997
rect 733 -999 734 -997
rect 730 -1005 731 -1003
rect 733 -1005 734 -1003
rect 737 -999 738 -997
rect 737 -1005 738 -1003
rect 744 -999 745 -997
rect 744 -1005 745 -1003
rect 751 -999 752 -997
rect 751 -1005 752 -1003
rect 758 -999 759 -997
rect 758 -1005 759 -1003
rect 765 -999 766 -997
rect 768 -999 769 -997
rect 765 -1005 766 -1003
rect 768 -1005 769 -1003
rect 772 -999 773 -997
rect 775 -999 776 -997
rect 775 -1005 776 -1003
rect 779 -999 780 -997
rect 779 -1005 780 -1003
rect 786 -999 787 -997
rect 786 -1005 787 -1003
rect 793 -999 794 -997
rect 793 -1005 794 -1003
rect 800 -999 801 -997
rect 800 -1005 801 -1003
rect 807 -999 808 -997
rect 807 -1005 808 -1003
rect 814 -999 815 -997
rect 814 -1005 815 -1003
rect 821 -999 822 -997
rect 821 -1005 822 -1003
rect 828 -999 829 -997
rect 828 -1005 829 -1003
rect 835 -999 836 -997
rect 835 -1005 836 -1003
rect 842 -999 843 -997
rect 845 -999 846 -997
rect 842 -1005 843 -1003
rect 845 -1005 846 -1003
rect 849 -999 850 -997
rect 849 -1005 850 -1003
rect 856 -999 857 -997
rect 856 -1005 857 -1003
rect 863 -999 864 -997
rect 863 -1005 864 -1003
rect 870 -999 871 -997
rect 870 -1005 871 -1003
rect 877 -999 878 -997
rect 877 -1005 878 -1003
rect 884 -999 885 -997
rect 887 -1005 888 -1003
rect 891 -999 892 -997
rect 891 -1005 892 -1003
rect 898 -999 899 -997
rect 901 -999 902 -997
rect 898 -1005 899 -1003
rect 901 -1005 902 -1003
rect 905 -999 906 -997
rect 905 -1005 906 -1003
rect 912 -999 913 -997
rect 912 -1005 913 -1003
rect 919 -999 920 -997
rect 919 -1005 920 -1003
rect 926 -999 927 -997
rect 929 -999 930 -997
rect 926 -1005 927 -1003
rect 933 -999 934 -997
rect 933 -1005 934 -1003
rect 940 -999 941 -997
rect 940 -1005 941 -1003
rect 947 -999 948 -997
rect 947 -1005 948 -1003
rect 954 -999 955 -997
rect 954 -1005 955 -1003
rect 961 -999 962 -997
rect 964 -999 965 -997
rect 961 -1005 962 -1003
rect 968 -999 969 -997
rect 968 -1005 969 -1003
rect 975 -999 976 -997
rect 978 -999 979 -997
rect 978 -1005 979 -1003
rect 982 -999 983 -997
rect 985 -999 986 -997
rect 982 -1005 983 -1003
rect 985 -1005 986 -1003
rect 992 -999 993 -997
rect 989 -1005 990 -1003
rect 992 -1005 993 -1003
rect 996 -999 997 -997
rect 999 -999 1000 -997
rect 996 -1005 997 -1003
rect 999 -1005 1000 -1003
rect 1003 -999 1004 -997
rect 1003 -1005 1004 -1003
rect 1010 -999 1011 -997
rect 1010 -1005 1011 -1003
rect 1013 -1005 1014 -1003
rect 1017 -999 1018 -997
rect 1017 -1005 1018 -1003
rect 1024 -999 1025 -997
rect 1024 -1005 1025 -1003
rect 1027 -1005 1028 -1003
rect 1031 -999 1032 -997
rect 1031 -1005 1032 -1003
rect 1038 -999 1039 -997
rect 1038 -1005 1039 -1003
rect 1045 -999 1046 -997
rect 1045 -1005 1046 -1003
rect 1052 -999 1053 -997
rect 1052 -1005 1053 -1003
rect 1059 -999 1060 -997
rect 1059 -1005 1060 -1003
rect 1066 -999 1067 -997
rect 1066 -1005 1067 -1003
rect 1073 -999 1074 -997
rect 1073 -1005 1074 -1003
rect 1080 -999 1081 -997
rect 1080 -1005 1081 -1003
rect 1087 -999 1088 -997
rect 1087 -1005 1088 -1003
rect 1094 -999 1095 -997
rect 1094 -1005 1095 -1003
rect 1101 -999 1102 -997
rect 1101 -1005 1102 -1003
rect 1111 -999 1112 -997
rect 1108 -1005 1109 -1003
rect 1111 -1005 1112 -1003
rect 1115 -999 1116 -997
rect 1115 -1005 1116 -1003
rect 1122 -999 1123 -997
rect 1122 -1005 1123 -1003
rect 1129 -999 1130 -997
rect 1129 -1005 1130 -1003
rect 1132 -1005 1133 -1003
rect 1136 -999 1137 -997
rect 1136 -1005 1137 -1003
rect 1143 -999 1144 -997
rect 1143 -1005 1144 -1003
rect 1150 -999 1151 -997
rect 1150 -1005 1151 -1003
rect 1157 -999 1158 -997
rect 1157 -1005 1158 -1003
rect 1164 -999 1165 -997
rect 1164 -1005 1165 -1003
rect 1171 -999 1172 -997
rect 1171 -1005 1172 -1003
rect 1178 -999 1179 -997
rect 1178 -1005 1179 -1003
rect 1185 -999 1186 -997
rect 1185 -1005 1186 -1003
rect 1192 -999 1193 -997
rect 1192 -1005 1193 -1003
rect 1199 -999 1200 -997
rect 1199 -1005 1200 -1003
rect 1206 -999 1207 -997
rect 1206 -1005 1207 -1003
rect 1213 -999 1214 -997
rect 1213 -1005 1214 -1003
rect 1220 -999 1221 -997
rect 1220 -1005 1221 -1003
rect 1227 -999 1228 -997
rect 1227 -1005 1228 -1003
rect 1234 -999 1235 -997
rect 1234 -1005 1235 -1003
rect 1241 -999 1242 -997
rect 1241 -1005 1242 -1003
rect 1248 -999 1249 -997
rect 1248 -1005 1249 -1003
rect 1255 -999 1256 -997
rect 1255 -1005 1256 -1003
rect 1262 -999 1263 -997
rect 1262 -1005 1263 -1003
rect 1269 -999 1270 -997
rect 1269 -1005 1270 -1003
rect 1276 -999 1277 -997
rect 1276 -1005 1277 -1003
rect 1283 -999 1284 -997
rect 1283 -1005 1284 -1003
rect 1290 -999 1291 -997
rect 1290 -1005 1291 -1003
rect 1297 -999 1298 -997
rect 1297 -1005 1298 -1003
rect 1304 -999 1305 -997
rect 1304 -1005 1305 -1003
rect 1311 -999 1312 -997
rect 1311 -1005 1312 -1003
rect 1318 -999 1319 -997
rect 1318 -1005 1319 -1003
rect 1325 -999 1326 -997
rect 1325 -1005 1326 -1003
rect 1332 -999 1333 -997
rect 1332 -1005 1333 -1003
rect 1339 -999 1340 -997
rect 1339 -1005 1340 -1003
rect 1346 -999 1347 -997
rect 1346 -1005 1347 -1003
rect 1353 -999 1354 -997
rect 1353 -1005 1354 -1003
rect 1360 -999 1361 -997
rect 1360 -1005 1361 -1003
rect 1367 -999 1368 -997
rect 1367 -1005 1368 -1003
rect 1374 -999 1375 -997
rect 1374 -1005 1375 -1003
rect 1381 -999 1382 -997
rect 1381 -1005 1382 -1003
rect 1388 -999 1389 -997
rect 1388 -1005 1389 -1003
rect 1395 -999 1396 -997
rect 1395 -1005 1396 -1003
rect 1402 -999 1403 -997
rect 1402 -1005 1403 -1003
rect 1409 -999 1410 -997
rect 1409 -1005 1410 -1003
rect 1416 -999 1417 -997
rect 1416 -1005 1417 -1003
rect 1423 -999 1424 -997
rect 1423 -1005 1424 -1003
rect 1430 -999 1431 -997
rect 1430 -1005 1431 -1003
rect 1437 -999 1438 -997
rect 1437 -1005 1438 -1003
rect 1444 -999 1445 -997
rect 1444 -1005 1445 -1003
rect 1451 -999 1452 -997
rect 1451 -1005 1452 -1003
rect 1458 -999 1459 -997
rect 1458 -1005 1459 -1003
rect 1465 -999 1466 -997
rect 1465 -1005 1466 -1003
rect 1472 -999 1473 -997
rect 1472 -1005 1473 -1003
rect 1479 -999 1480 -997
rect 1479 -1005 1480 -1003
rect 1486 -999 1487 -997
rect 1486 -1005 1487 -1003
rect 1493 -999 1494 -997
rect 1493 -1005 1494 -1003
rect 1500 -999 1501 -997
rect 1500 -1005 1501 -1003
rect 1507 -999 1508 -997
rect 1507 -1005 1508 -1003
rect 1514 -999 1515 -997
rect 1514 -1005 1515 -1003
rect 1521 -999 1522 -997
rect 1521 -1005 1522 -1003
rect 1528 -999 1529 -997
rect 1528 -1005 1529 -1003
rect 1535 -999 1536 -997
rect 1535 -1005 1536 -1003
rect 1542 -999 1543 -997
rect 1542 -1005 1543 -1003
rect 1549 -999 1550 -997
rect 1549 -1005 1550 -1003
rect 1552 -1005 1553 -1003
rect 1556 -999 1557 -997
rect 1556 -1005 1557 -1003
rect 1563 -999 1564 -997
rect 1566 -999 1567 -997
rect 1563 -1005 1564 -1003
rect 1566 -1005 1567 -1003
rect 1570 -999 1571 -997
rect 1573 -999 1574 -997
rect 1570 -1005 1571 -1003
rect 1577 -999 1578 -997
rect 1577 -1005 1578 -1003
rect 1584 -999 1585 -997
rect 1584 -1005 1585 -1003
rect 1591 -999 1592 -997
rect 1591 -1005 1592 -1003
rect 1598 -999 1599 -997
rect 1598 -1005 1599 -1003
rect 1605 -999 1606 -997
rect 1605 -1005 1606 -1003
rect 1612 -999 1613 -997
rect 1612 -1005 1613 -1003
rect 1619 -999 1620 -997
rect 1619 -1005 1620 -1003
rect 1626 -999 1627 -997
rect 1626 -1005 1627 -1003
rect 1633 -999 1634 -997
rect 1633 -1005 1634 -1003
rect 1738 -999 1739 -997
rect 1738 -1005 1739 -1003
rect 23 -1100 24 -1098
rect 23 -1106 24 -1104
rect 30 -1100 31 -1098
rect 30 -1106 31 -1104
rect 44 -1100 45 -1098
rect 44 -1106 45 -1104
rect 51 -1100 52 -1098
rect 51 -1106 52 -1104
rect 58 -1100 59 -1098
rect 58 -1106 59 -1104
rect 65 -1106 66 -1104
rect 72 -1100 73 -1098
rect 75 -1100 76 -1098
rect 75 -1106 76 -1104
rect 79 -1100 80 -1098
rect 79 -1106 80 -1104
rect 86 -1100 87 -1098
rect 89 -1100 90 -1098
rect 86 -1106 87 -1104
rect 89 -1106 90 -1104
rect 93 -1100 94 -1098
rect 93 -1106 94 -1104
rect 100 -1100 101 -1098
rect 100 -1106 101 -1104
rect 107 -1100 108 -1098
rect 107 -1106 108 -1104
rect 114 -1100 115 -1098
rect 114 -1106 115 -1104
rect 121 -1100 122 -1098
rect 121 -1106 122 -1104
rect 128 -1100 129 -1098
rect 128 -1106 129 -1104
rect 135 -1100 136 -1098
rect 138 -1100 139 -1098
rect 138 -1106 139 -1104
rect 142 -1100 143 -1098
rect 142 -1106 143 -1104
rect 149 -1100 150 -1098
rect 149 -1106 150 -1104
rect 156 -1100 157 -1098
rect 156 -1106 157 -1104
rect 163 -1100 164 -1098
rect 163 -1106 164 -1104
rect 170 -1100 171 -1098
rect 170 -1106 171 -1104
rect 177 -1100 178 -1098
rect 177 -1106 178 -1104
rect 184 -1100 185 -1098
rect 184 -1106 185 -1104
rect 191 -1100 192 -1098
rect 191 -1106 192 -1104
rect 198 -1100 199 -1098
rect 198 -1106 199 -1104
rect 205 -1100 206 -1098
rect 205 -1106 206 -1104
rect 212 -1100 213 -1098
rect 215 -1100 216 -1098
rect 212 -1106 213 -1104
rect 219 -1100 220 -1098
rect 219 -1106 220 -1104
rect 226 -1100 227 -1098
rect 226 -1106 227 -1104
rect 236 -1100 237 -1098
rect 233 -1106 234 -1104
rect 236 -1106 237 -1104
rect 240 -1106 241 -1104
rect 250 -1100 251 -1098
rect 247 -1106 248 -1104
rect 250 -1106 251 -1104
rect 254 -1100 255 -1098
rect 254 -1106 255 -1104
rect 261 -1106 262 -1104
rect 268 -1100 269 -1098
rect 268 -1106 269 -1104
rect 275 -1100 276 -1098
rect 275 -1106 276 -1104
rect 282 -1100 283 -1098
rect 282 -1106 283 -1104
rect 289 -1100 290 -1098
rect 289 -1106 290 -1104
rect 296 -1100 297 -1098
rect 296 -1106 297 -1104
rect 303 -1100 304 -1098
rect 303 -1106 304 -1104
rect 310 -1100 311 -1098
rect 310 -1106 311 -1104
rect 317 -1100 318 -1098
rect 317 -1106 318 -1104
rect 324 -1100 325 -1098
rect 324 -1106 325 -1104
rect 331 -1100 332 -1098
rect 331 -1106 332 -1104
rect 338 -1100 339 -1098
rect 338 -1106 339 -1104
rect 341 -1106 342 -1104
rect 345 -1100 346 -1098
rect 345 -1106 346 -1104
rect 352 -1100 353 -1098
rect 352 -1106 353 -1104
rect 359 -1100 360 -1098
rect 359 -1106 360 -1104
rect 366 -1100 367 -1098
rect 366 -1106 367 -1104
rect 373 -1100 374 -1098
rect 373 -1106 374 -1104
rect 380 -1100 381 -1098
rect 380 -1106 381 -1104
rect 387 -1100 388 -1098
rect 387 -1106 388 -1104
rect 394 -1100 395 -1098
rect 397 -1100 398 -1098
rect 394 -1106 395 -1104
rect 397 -1106 398 -1104
rect 401 -1100 402 -1098
rect 401 -1106 402 -1104
rect 408 -1100 409 -1098
rect 408 -1106 409 -1104
rect 415 -1100 416 -1098
rect 415 -1106 416 -1104
rect 425 -1106 426 -1104
rect 429 -1100 430 -1098
rect 429 -1106 430 -1104
rect 436 -1100 437 -1098
rect 436 -1106 437 -1104
rect 443 -1100 444 -1098
rect 443 -1106 444 -1104
rect 450 -1100 451 -1098
rect 450 -1106 451 -1104
rect 457 -1100 458 -1098
rect 457 -1106 458 -1104
rect 464 -1100 465 -1098
rect 464 -1106 465 -1104
rect 471 -1100 472 -1098
rect 471 -1106 472 -1104
rect 481 -1100 482 -1098
rect 481 -1106 482 -1104
rect 485 -1100 486 -1098
rect 485 -1106 486 -1104
rect 492 -1100 493 -1098
rect 492 -1106 493 -1104
rect 499 -1100 500 -1098
rect 499 -1106 500 -1104
rect 506 -1100 507 -1098
rect 506 -1106 507 -1104
rect 513 -1100 514 -1098
rect 516 -1100 517 -1098
rect 516 -1106 517 -1104
rect 520 -1100 521 -1098
rect 520 -1106 521 -1104
rect 527 -1100 528 -1098
rect 527 -1106 528 -1104
rect 534 -1100 535 -1098
rect 534 -1106 535 -1104
rect 541 -1100 542 -1098
rect 541 -1106 542 -1104
rect 548 -1100 549 -1098
rect 548 -1106 549 -1104
rect 555 -1100 556 -1098
rect 555 -1106 556 -1104
rect 562 -1100 563 -1098
rect 562 -1106 563 -1104
rect 569 -1100 570 -1098
rect 569 -1106 570 -1104
rect 576 -1100 577 -1098
rect 576 -1106 577 -1104
rect 583 -1100 584 -1098
rect 583 -1106 584 -1104
rect 590 -1100 591 -1098
rect 590 -1106 591 -1104
rect 597 -1100 598 -1098
rect 597 -1106 598 -1104
rect 604 -1100 605 -1098
rect 604 -1106 605 -1104
rect 611 -1100 612 -1098
rect 611 -1106 612 -1104
rect 618 -1100 619 -1098
rect 618 -1106 619 -1104
rect 625 -1100 626 -1098
rect 628 -1100 629 -1098
rect 625 -1106 626 -1104
rect 632 -1100 633 -1098
rect 632 -1106 633 -1104
rect 639 -1100 640 -1098
rect 642 -1100 643 -1098
rect 639 -1106 640 -1104
rect 646 -1100 647 -1098
rect 649 -1100 650 -1098
rect 649 -1106 650 -1104
rect 653 -1100 654 -1098
rect 653 -1106 654 -1104
rect 660 -1100 661 -1098
rect 660 -1106 661 -1104
rect 667 -1100 668 -1098
rect 667 -1106 668 -1104
rect 674 -1100 675 -1098
rect 677 -1100 678 -1098
rect 674 -1106 675 -1104
rect 677 -1106 678 -1104
rect 681 -1100 682 -1098
rect 681 -1106 682 -1104
rect 688 -1100 689 -1098
rect 688 -1106 689 -1104
rect 691 -1106 692 -1104
rect 695 -1100 696 -1098
rect 698 -1100 699 -1098
rect 695 -1106 696 -1104
rect 698 -1106 699 -1104
rect 702 -1100 703 -1098
rect 702 -1106 703 -1104
rect 709 -1100 710 -1098
rect 709 -1106 710 -1104
rect 716 -1100 717 -1098
rect 716 -1106 717 -1104
rect 723 -1100 724 -1098
rect 723 -1106 724 -1104
rect 730 -1100 731 -1098
rect 733 -1100 734 -1098
rect 730 -1106 731 -1104
rect 733 -1106 734 -1104
rect 737 -1100 738 -1098
rect 737 -1106 738 -1104
rect 744 -1100 745 -1098
rect 744 -1106 745 -1104
rect 751 -1100 752 -1098
rect 751 -1106 752 -1104
rect 758 -1100 759 -1098
rect 758 -1106 759 -1104
rect 765 -1100 766 -1098
rect 765 -1106 766 -1104
rect 772 -1100 773 -1098
rect 772 -1106 773 -1104
rect 779 -1100 780 -1098
rect 779 -1106 780 -1104
rect 786 -1100 787 -1098
rect 786 -1106 787 -1104
rect 793 -1100 794 -1098
rect 793 -1106 794 -1104
rect 800 -1100 801 -1098
rect 803 -1100 804 -1098
rect 803 -1106 804 -1104
rect 807 -1100 808 -1098
rect 807 -1106 808 -1104
rect 814 -1100 815 -1098
rect 814 -1106 815 -1104
rect 821 -1100 822 -1098
rect 821 -1106 822 -1104
rect 828 -1100 829 -1098
rect 828 -1106 829 -1104
rect 835 -1100 836 -1098
rect 835 -1106 836 -1104
rect 842 -1100 843 -1098
rect 842 -1106 843 -1104
rect 849 -1100 850 -1098
rect 849 -1106 850 -1104
rect 856 -1100 857 -1098
rect 856 -1106 857 -1104
rect 863 -1100 864 -1098
rect 866 -1100 867 -1098
rect 863 -1106 864 -1104
rect 866 -1106 867 -1104
rect 870 -1100 871 -1098
rect 870 -1106 871 -1104
rect 877 -1100 878 -1098
rect 880 -1100 881 -1098
rect 877 -1106 878 -1104
rect 880 -1106 881 -1104
rect 884 -1100 885 -1098
rect 887 -1100 888 -1098
rect 887 -1106 888 -1104
rect 891 -1100 892 -1098
rect 894 -1100 895 -1098
rect 891 -1106 892 -1104
rect 894 -1106 895 -1104
rect 898 -1100 899 -1098
rect 898 -1106 899 -1104
rect 905 -1100 906 -1098
rect 905 -1106 906 -1104
rect 912 -1100 913 -1098
rect 912 -1106 913 -1104
rect 919 -1100 920 -1098
rect 919 -1106 920 -1104
rect 926 -1100 927 -1098
rect 926 -1106 927 -1104
rect 933 -1100 934 -1098
rect 933 -1106 934 -1104
rect 940 -1100 941 -1098
rect 940 -1106 941 -1104
rect 947 -1100 948 -1098
rect 947 -1106 948 -1104
rect 954 -1100 955 -1098
rect 954 -1106 955 -1104
rect 961 -1100 962 -1098
rect 961 -1106 962 -1104
rect 968 -1100 969 -1098
rect 968 -1106 969 -1104
rect 975 -1100 976 -1098
rect 975 -1106 976 -1104
rect 982 -1100 983 -1098
rect 982 -1106 983 -1104
rect 989 -1100 990 -1098
rect 989 -1106 990 -1104
rect 996 -1100 997 -1098
rect 996 -1106 997 -1104
rect 1003 -1100 1004 -1098
rect 1006 -1100 1007 -1098
rect 1003 -1106 1004 -1104
rect 1010 -1100 1011 -1098
rect 1010 -1106 1011 -1104
rect 1017 -1100 1018 -1098
rect 1017 -1106 1018 -1104
rect 1024 -1100 1025 -1098
rect 1027 -1100 1028 -1098
rect 1024 -1106 1025 -1104
rect 1031 -1100 1032 -1098
rect 1031 -1106 1032 -1104
rect 1038 -1100 1039 -1098
rect 1038 -1106 1039 -1104
rect 1045 -1100 1046 -1098
rect 1045 -1106 1046 -1104
rect 1048 -1106 1049 -1104
rect 1055 -1100 1056 -1098
rect 1052 -1106 1053 -1104
rect 1055 -1106 1056 -1104
rect 1059 -1100 1060 -1098
rect 1059 -1106 1060 -1104
rect 1066 -1100 1067 -1098
rect 1066 -1106 1067 -1104
rect 1073 -1100 1074 -1098
rect 1073 -1106 1074 -1104
rect 1080 -1100 1081 -1098
rect 1080 -1106 1081 -1104
rect 1087 -1100 1088 -1098
rect 1090 -1100 1091 -1098
rect 1087 -1106 1088 -1104
rect 1094 -1100 1095 -1098
rect 1094 -1106 1095 -1104
rect 1101 -1100 1102 -1098
rect 1101 -1106 1102 -1104
rect 1108 -1100 1109 -1098
rect 1108 -1106 1109 -1104
rect 1115 -1100 1116 -1098
rect 1115 -1106 1116 -1104
rect 1122 -1100 1123 -1098
rect 1122 -1106 1123 -1104
rect 1129 -1100 1130 -1098
rect 1132 -1100 1133 -1098
rect 1129 -1106 1130 -1104
rect 1136 -1100 1137 -1098
rect 1136 -1106 1137 -1104
rect 1143 -1100 1144 -1098
rect 1143 -1106 1144 -1104
rect 1150 -1100 1151 -1098
rect 1150 -1106 1151 -1104
rect 1157 -1100 1158 -1098
rect 1157 -1106 1158 -1104
rect 1164 -1100 1165 -1098
rect 1164 -1106 1165 -1104
rect 1171 -1100 1172 -1098
rect 1171 -1106 1172 -1104
rect 1178 -1100 1179 -1098
rect 1178 -1106 1179 -1104
rect 1185 -1100 1186 -1098
rect 1185 -1106 1186 -1104
rect 1192 -1100 1193 -1098
rect 1192 -1106 1193 -1104
rect 1199 -1100 1200 -1098
rect 1199 -1106 1200 -1104
rect 1206 -1100 1207 -1098
rect 1206 -1106 1207 -1104
rect 1213 -1100 1214 -1098
rect 1213 -1106 1214 -1104
rect 1220 -1100 1221 -1098
rect 1220 -1106 1221 -1104
rect 1227 -1100 1228 -1098
rect 1227 -1106 1228 -1104
rect 1234 -1100 1235 -1098
rect 1234 -1106 1235 -1104
rect 1241 -1100 1242 -1098
rect 1241 -1106 1242 -1104
rect 1248 -1100 1249 -1098
rect 1248 -1106 1249 -1104
rect 1255 -1100 1256 -1098
rect 1255 -1106 1256 -1104
rect 1262 -1100 1263 -1098
rect 1262 -1106 1263 -1104
rect 1269 -1100 1270 -1098
rect 1269 -1106 1270 -1104
rect 1276 -1100 1277 -1098
rect 1276 -1106 1277 -1104
rect 1283 -1100 1284 -1098
rect 1283 -1106 1284 -1104
rect 1290 -1100 1291 -1098
rect 1290 -1106 1291 -1104
rect 1297 -1100 1298 -1098
rect 1297 -1106 1298 -1104
rect 1304 -1100 1305 -1098
rect 1304 -1106 1305 -1104
rect 1311 -1100 1312 -1098
rect 1311 -1106 1312 -1104
rect 1318 -1100 1319 -1098
rect 1318 -1106 1319 -1104
rect 1325 -1100 1326 -1098
rect 1325 -1106 1326 -1104
rect 1332 -1100 1333 -1098
rect 1332 -1106 1333 -1104
rect 1339 -1100 1340 -1098
rect 1339 -1106 1340 -1104
rect 1346 -1100 1347 -1098
rect 1346 -1106 1347 -1104
rect 1353 -1100 1354 -1098
rect 1353 -1106 1354 -1104
rect 1360 -1100 1361 -1098
rect 1360 -1106 1361 -1104
rect 1367 -1100 1368 -1098
rect 1367 -1106 1368 -1104
rect 1374 -1100 1375 -1098
rect 1374 -1106 1375 -1104
rect 1381 -1100 1382 -1098
rect 1384 -1100 1385 -1098
rect 1381 -1106 1382 -1104
rect 1384 -1106 1385 -1104
rect 1388 -1100 1389 -1098
rect 1388 -1106 1389 -1104
rect 1395 -1100 1396 -1098
rect 1395 -1106 1396 -1104
rect 1402 -1100 1403 -1098
rect 1402 -1106 1403 -1104
rect 1409 -1100 1410 -1098
rect 1409 -1106 1410 -1104
rect 1416 -1100 1417 -1098
rect 1416 -1106 1417 -1104
rect 1423 -1100 1424 -1098
rect 1423 -1106 1424 -1104
rect 1430 -1100 1431 -1098
rect 1430 -1106 1431 -1104
rect 1437 -1100 1438 -1098
rect 1437 -1106 1438 -1104
rect 1444 -1100 1445 -1098
rect 1444 -1106 1445 -1104
rect 1451 -1100 1452 -1098
rect 1451 -1106 1452 -1104
rect 1454 -1106 1455 -1104
rect 1458 -1100 1459 -1098
rect 1458 -1106 1459 -1104
rect 1465 -1100 1466 -1098
rect 1465 -1106 1466 -1104
rect 1472 -1100 1473 -1098
rect 1475 -1100 1476 -1098
rect 1475 -1106 1476 -1104
rect 1479 -1100 1480 -1098
rect 1479 -1106 1480 -1104
rect 1486 -1100 1487 -1098
rect 1486 -1106 1487 -1104
rect 1493 -1100 1494 -1098
rect 1493 -1106 1494 -1104
rect 1496 -1106 1497 -1104
rect 1500 -1100 1501 -1098
rect 1500 -1106 1501 -1104
rect 1507 -1100 1508 -1098
rect 1507 -1106 1508 -1104
rect 1514 -1100 1515 -1098
rect 1514 -1106 1515 -1104
rect 1521 -1100 1522 -1098
rect 1521 -1106 1522 -1104
rect 1528 -1100 1529 -1098
rect 1528 -1106 1529 -1104
rect 1535 -1100 1536 -1098
rect 1535 -1106 1536 -1104
rect 1542 -1100 1543 -1098
rect 1542 -1106 1543 -1104
rect 1549 -1100 1550 -1098
rect 1549 -1106 1550 -1104
rect 1556 -1100 1557 -1098
rect 1556 -1106 1557 -1104
rect 1563 -1100 1564 -1098
rect 1563 -1106 1564 -1104
rect 1570 -1100 1571 -1098
rect 1570 -1106 1571 -1104
rect 1577 -1100 1578 -1098
rect 1577 -1106 1578 -1104
rect 1584 -1100 1585 -1098
rect 1584 -1106 1585 -1104
rect 1591 -1100 1592 -1098
rect 1591 -1106 1592 -1104
rect 1598 -1100 1599 -1098
rect 1598 -1106 1599 -1104
rect 1605 -1100 1606 -1098
rect 1605 -1106 1606 -1104
rect 1612 -1100 1613 -1098
rect 1612 -1106 1613 -1104
rect 1619 -1100 1620 -1098
rect 1619 -1106 1620 -1104
rect 1626 -1100 1627 -1098
rect 1626 -1106 1627 -1104
rect 1633 -1100 1634 -1098
rect 1633 -1106 1634 -1104
rect 1640 -1100 1641 -1098
rect 1640 -1106 1641 -1104
rect 1647 -1100 1648 -1098
rect 1647 -1106 1648 -1104
rect 1654 -1100 1655 -1098
rect 1654 -1106 1655 -1104
rect 1675 -1100 1676 -1098
rect 1675 -1106 1676 -1104
rect 1682 -1100 1683 -1098
rect 1682 -1106 1683 -1104
rect 1745 -1100 1746 -1098
rect 1745 -1106 1746 -1104
rect 23 -1219 24 -1217
rect 23 -1225 24 -1223
rect 30 -1219 31 -1217
rect 30 -1225 31 -1223
rect 37 -1219 38 -1217
rect 37 -1225 38 -1223
rect 44 -1219 45 -1217
rect 44 -1225 45 -1223
rect 51 -1219 52 -1217
rect 51 -1225 52 -1223
rect 58 -1219 59 -1217
rect 58 -1225 59 -1223
rect 65 -1219 66 -1217
rect 68 -1219 69 -1217
rect 65 -1225 66 -1223
rect 68 -1225 69 -1223
rect 72 -1219 73 -1217
rect 72 -1225 73 -1223
rect 79 -1219 80 -1217
rect 79 -1225 80 -1223
rect 86 -1219 87 -1217
rect 89 -1219 90 -1217
rect 86 -1225 87 -1223
rect 89 -1225 90 -1223
rect 93 -1219 94 -1217
rect 93 -1225 94 -1223
rect 100 -1219 101 -1217
rect 100 -1225 101 -1223
rect 110 -1219 111 -1217
rect 107 -1225 108 -1223
rect 110 -1225 111 -1223
rect 114 -1219 115 -1217
rect 114 -1225 115 -1223
rect 121 -1219 122 -1217
rect 124 -1219 125 -1217
rect 121 -1225 122 -1223
rect 124 -1225 125 -1223
rect 128 -1219 129 -1217
rect 128 -1225 129 -1223
rect 135 -1219 136 -1217
rect 135 -1225 136 -1223
rect 142 -1219 143 -1217
rect 145 -1219 146 -1217
rect 142 -1225 143 -1223
rect 145 -1225 146 -1223
rect 149 -1219 150 -1217
rect 149 -1225 150 -1223
rect 156 -1219 157 -1217
rect 156 -1225 157 -1223
rect 163 -1219 164 -1217
rect 163 -1225 164 -1223
rect 170 -1219 171 -1217
rect 173 -1219 174 -1217
rect 170 -1225 171 -1223
rect 173 -1225 174 -1223
rect 177 -1219 178 -1217
rect 180 -1219 181 -1217
rect 177 -1225 178 -1223
rect 180 -1225 181 -1223
rect 184 -1219 185 -1217
rect 184 -1225 185 -1223
rect 191 -1219 192 -1217
rect 191 -1225 192 -1223
rect 198 -1219 199 -1217
rect 198 -1225 199 -1223
rect 205 -1219 206 -1217
rect 205 -1225 206 -1223
rect 212 -1219 213 -1217
rect 212 -1225 213 -1223
rect 219 -1219 220 -1217
rect 219 -1225 220 -1223
rect 226 -1219 227 -1217
rect 229 -1219 230 -1217
rect 226 -1225 227 -1223
rect 233 -1219 234 -1217
rect 233 -1225 234 -1223
rect 240 -1219 241 -1217
rect 243 -1219 244 -1217
rect 243 -1225 244 -1223
rect 247 -1219 248 -1217
rect 247 -1225 248 -1223
rect 254 -1219 255 -1217
rect 254 -1225 255 -1223
rect 264 -1219 265 -1217
rect 264 -1225 265 -1223
rect 268 -1219 269 -1217
rect 268 -1225 269 -1223
rect 275 -1219 276 -1217
rect 275 -1225 276 -1223
rect 282 -1219 283 -1217
rect 282 -1225 283 -1223
rect 289 -1219 290 -1217
rect 289 -1225 290 -1223
rect 296 -1219 297 -1217
rect 296 -1225 297 -1223
rect 303 -1219 304 -1217
rect 303 -1225 304 -1223
rect 310 -1219 311 -1217
rect 310 -1225 311 -1223
rect 317 -1219 318 -1217
rect 317 -1225 318 -1223
rect 324 -1219 325 -1217
rect 324 -1225 325 -1223
rect 331 -1219 332 -1217
rect 331 -1225 332 -1223
rect 338 -1219 339 -1217
rect 338 -1225 339 -1223
rect 345 -1219 346 -1217
rect 345 -1225 346 -1223
rect 352 -1219 353 -1217
rect 352 -1225 353 -1223
rect 359 -1219 360 -1217
rect 359 -1225 360 -1223
rect 366 -1219 367 -1217
rect 366 -1225 367 -1223
rect 373 -1219 374 -1217
rect 373 -1225 374 -1223
rect 380 -1219 381 -1217
rect 380 -1225 381 -1223
rect 387 -1219 388 -1217
rect 387 -1225 388 -1223
rect 394 -1219 395 -1217
rect 394 -1225 395 -1223
rect 401 -1219 402 -1217
rect 401 -1225 402 -1223
rect 408 -1219 409 -1217
rect 408 -1225 409 -1223
rect 415 -1219 416 -1217
rect 415 -1225 416 -1223
rect 422 -1219 423 -1217
rect 422 -1225 423 -1223
rect 429 -1219 430 -1217
rect 429 -1225 430 -1223
rect 436 -1219 437 -1217
rect 439 -1219 440 -1217
rect 436 -1225 437 -1223
rect 443 -1219 444 -1217
rect 443 -1225 444 -1223
rect 450 -1219 451 -1217
rect 450 -1225 451 -1223
rect 457 -1219 458 -1217
rect 457 -1225 458 -1223
rect 464 -1219 465 -1217
rect 464 -1225 465 -1223
rect 471 -1219 472 -1217
rect 471 -1225 472 -1223
rect 478 -1219 479 -1217
rect 478 -1225 479 -1223
rect 485 -1219 486 -1217
rect 485 -1225 486 -1223
rect 492 -1219 493 -1217
rect 492 -1225 493 -1223
rect 499 -1219 500 -1217
rect 499 -1225 500 -1223
rect 506 -1225 507 -1223
rect 509 -1225 510 -1223
rect 513 -1219 514 -1217
rect 513 -1225 514 -1223
rect 520 -1219 521 -1217
rect 520 -1225 521 -1223
rect 527 -1219 528 -1217
rect 527 -1225 528 -1223
rect 534 -1219 535 -1217
rect 534 -1225 535 -1223
rect 541 -1219 542 -1217
rect 544 -1219 545 -1217
rect 541 -1225 542 -1223
rect 548 -1219 549 -1217
rect 548 -1225 549 -1223
rect 555 -1219 556 -1217
rect 555 -1225 556 -1223
rect 562 -1219 563 -1217
rect 562 -1225 563 -1223
rect 565 -1225 566 -1223
rect 569 -1219 570 -1217
rect 569 -1225 570 -1223
rect 576 -1219 577 -1217
rect 576 -1225 577 -1223
rect 583 -1219 584 -1217
rect 583 -1225 584 -1223
rect 590 -1219 591 -1217
rect 590 -1225 591 -1223
rect 597 -1219 598 -1217
rect 597 -1225 598 -1223
rect 604 -1219 605 -1217
rect 604 -1225 605 -1223
rect 607 -1225 608 -1223
rect 611 -1219 612 -1217
rect 611 -1225 612 -1223
rect 618 -1219 619 -1217
rect 618 -1225 619 -1223
rect 625 -1219 626 -1217
rect 625 -1225 626 -1223
rect 635 -1219 636 -1217
rect 632 -1225 633 -1223
rect 635 -1225 636 -1223
rect 639 -1219 640 -1217
rect 639 -1225 640 -1223
rect 646 -1219 647 -1217
rect 649 -1219 650 -1217
rect 656 -1219 657 -1217
rect 656 -1225 657 -1223
rect 660 -1219 661 -1217
rect 660 -1225 661 -1223
rect 667 -1219 668 -1217
rect 667 -1225 668 -1223
rect 674 -1219 675 -1217
rect 674 -1225 675 -1223
rect 681 -1219 682 -1217
rect 681 -1225 682 -1223
rect 688 -1219 689 -1217
rect 688 -1225 689 -1223
rect 695 -1219 696 -1217
rect 698 -1219 699 -1217
rect 695 -1225 696 -1223
rect 698 -1225 699 -1223
rect 702 -1219 703 -1217
rect 702 -1225 703 -1223
rect 705 -1225 706 -1223
rect 709 -1219 710 -1217
rect 709 -1225 710 -1223
rect 716 -1219 717 -1217
rect 716 -1225 717 -1223
rect 723 -1219 724 -1217
rect 723 -1225 724 -1223
rect 730 -1219 731 -1217
rect 730 -1225 731 -1223
rect 737 -1219 738 -1217
rect 740 -1219 741 -1217
rect 737 -1225 738 -1223
rect 740 -1225 741 -1223
rect 744 -1219 745 -1217
rect 744 -1225 745 -1223
rect 751 -1219 752 -1217
rect 751 -1225 752 -1223
rect 758 -1219 759 -1217
rect 758 -1225 759 -1223
rect 765 -1219 766 -1217
rect 768 -1219 769 -1217
rect 768 -1225 769 -1223
rect 772 -1219 773 -1217
rect 772 -1225 773 -1223
rect 779 -1219 780 -1217
rect 779 -1225 780 -1223
rect 786 -1219 787 -1217
rect 786 -1225 787 -1223
rect 793 -1219 794 -1217
rect 796 -1219 797 -1217
rect 793 -1225 794 -1223
rect 796 -1225 797 -1223
rect 800 -1219 801 -1217
rect 800 -1225 801 -1223
rect 807 -1219 808 -1217
rect 807 -1225 808 -1223
rect 814 -1219 815 -1217
rect 817 -1219 818 -1217
rect 814 -1225 815 -1223
rect 817 -1225 818 -1223
rect 821 -1219 822 -1217
rect 824 -1219 825 -1217
rect 821 -1225 822 -1223
rect 828 -1219 829 -1217
rect 831 -1219 832 -1217
rect 828 -1225 829 -1223
rect 831 -1225 832 -1223
rect 835 -1219 836 -1217
rect 835 -1225 836 -1223
rect 842 -1219 843 -1217
rect 842 -1225 843 -1223
rect 849 -1219 850 -1217
rect 849 -1225 850 -1223
rect 856 -1219 857 -1217
rect 859 -1219 860 -1217
rect 856 -1225 857 -1223
rect 859 -1225 860 -1223
rect 863 -1219 864 -1217
rect 863 -1225 864 -1223
rect 870 -1219 871 -1217
rect 870 -1225 871 -1223
rect 877 -1219 878 -1217
rect 877 -1225 878 -1223
rect 884 -1219 885 -1217
rect 884 -1225 885 -1223
rect 891 -1219 892 -1217
rect 894 -1219 895 -1217
rect 891 -1225 892 -1223
rect 894 -1225 895 -1223
rect 898 -1219 899 -1217
rect 898 -1225 899 -1223
rect 905 -1219 906 -1217
rect 905 -1225 906 -1223
rect 912 -1219 913 -1217
rect 912 -1225 913 -1223
rect 919 -1219 920 -1217
rect 919 -1225 920 -1223
rect 926 -1219 927 -1217
rect 929 -1219 930 -1217
rect 926 -1225 927 -1223
rect 929 -1225 930 -1223
rect 933 -1219 934 -1217
rect 933 -1225 934 -1223
rect 940 -1219 941 -1217
rect 940 -1225 941 -1223
rect 947 -1219 948 -1217
rect 950 -1219 951 -1217
rect 950 -1225 951 -1223
rect 954 -1219 955 -1217
rect 954 -1225 955 -1223
rect 961 -1219 962 -1217
rect 961 -1225 962 -1223
rect 968 -1219 969 -1217
rect 968 -1225 969 -1223
rect 975 -1219 976 -1217
rect 975 -1225 976 -1223
rect 982 -1219 983 -1217
rect 982 -1225 983 -1223
rect 989 -1219 990 -1217
rect 989 -1225 990 -1223
rect 996 -1219 997 -1217
rect 996 -1225 997 -1223
rect 1003 -1219 1004 -1217
rect 1003 -1225 1004 -1223
rect 1010 -1219 1011 -1217
rect 1010 -1225 1011 -1223
rect 1017 -1219 1018 -1217
rect 1017 -1225 1018 -1223
rect 1024 -1219 1025 -1217
rect 1024 -1225 1025 -1223
rect 1031 -1219 1032 -1217
rect 1031 -1225 1032 -1223
rect 1038 -1219 1039 -1217
rect 1038 -1225 1039 -1223
rect 1045 -1219 1046 -1217
rect 1045 -1225 1046 -1223
rect 1055 -1219 1056 -1217
rect 1052 -1225 1053 -1223
rect 1055 -1225 1056 -1223
rect 1059 -1219 1060 -1217
rect 1059 -1225 1060 -1223
rect 1066 -1219 1067 -1217
rect 1066 -1225 1067 -1223
rect 1073 -1219 1074 -1217
rect 1073 -1225 1074 -1223
rect 1080 -1219 1081 -1217
rect 1080 -1225 1081 -1223
rect 1087 -1219 1088 -1217
rect 1087 -1225 1088 -1223
rect 1094 -1219 1095 -1217
rect 1094 -1225 1095 -1223
rect 1101 -1219 1102 -1217
rect 1101 -1225 1102 -1223
rect 1108 -1219 1109 -1217
rect 1108 -1225 1109 -1223
rect 1115 -1219 1116 -1217
rect 1115 -1225 1116 -1223
rect 1122 -1219 1123 -1217
rect 1122 -1225 1123 -1223
rect 1129 -1219 1130 -1217
rect 1129 -1225 1130 -1223
rect 1136 -1219 1137 -1217
rect 1136 -1225 1137 -1223
rect 1143 -1219 1144 -1217
rect 1143 -1225 1144 -1223
rect 1150 -1219 1151 -1217
rect 1150 -1225 1151 -1223
rect 1157 -1219 1158 -1217
rect 1157 -1225 1158 -1223
rect 1164 -1219 1165 -1217
rect 1164 -1225 1165 -1223
rect 1171 -1219 1172 -1217
rect 1171 -1225 1172 -1223
rect 1178 -1219 1179 -1217
rect 1178 -1225 1179 -1223
rect 1185 -1219 1186 -1217
rect 1185 -1225 1186 -1223
rect 1192 -1219 1193 -1217
rect 1192 -1225 1193 -1223
rect 1199 -1219 1200 -1217
rect 1199 -1225 1200 -1223
rect 1206 -1219 1207 -1217
rect 1206 -1225 1207 -1223
rect 1213 -1219 1214 -1217
rect 1213 -1225 1214 -1223
rect 1220 -1219 1221 -1217
rect 1220 -1225 1221 -1223
rect 1227 -1219 1228 -1217
rect 1227 -1225 1228 -1223
rect 1234 -1219 1235 -1217
rect 1234 -1225 1235 -1223
rect 1241 -1219 1242 -1217
rect 1241 -1225 1242 -1223
rect 1248 -1219 1249 -1217
rect 1248 -1225 1249 -1223
rect 1255 -1219 1256 -1217
rect 1255 -1225 1256 -1223
rect 1262 -1219 1263 -1217
rect 1262 -1225 1263 -1223
rect 1269 -1219 1270 -1217
rect 1269 -1225 1270 -1223
rect 1276 -1219 1277 -1217
rect 1276 -1225 1277 -1223
rect 1283 -1219 1284 -1217
rect 1283 -1225 1284 -1223
rect 1290 -1219 1291 -1217
rect 1290 -1225 1291 -1223
rect 1297 -1219 1298 -1217
rect 1297 -1225 1298 -1223
rect 1304 -1219 1305 -1217
rect 1311 -1219 1312 -1217
rect 1311 -1225 1312 -1223
rect 1314 -1225 1315 -1223
rect 1318 -1219 1319 -1217
rect 1318 -1225 1319 -1223
rect 1325 -1219 1326 -1217
rect 1325 -1225 1326 -1223
rect 1332 -1219 1333 -1217
rect 1332 -1225 1333 -1223
rect 1339 -1219 1340 -1217
rect 1339 -1225 1340 -1223
rect 1346 -1219 1347 -1217
rect 1346 -1225 1347 -1223
rect 1353 -1219 1354 -1217
rect 1353 -1225 1354 -1223
rect 1360 -1219 1361 -1217
rect 1360 -1225 1361 -1223
rect 1367 -1219 1368 -1217
rect 1367 -1225 1368 -1223
rect 1374 -1219 1375 -1217
rect 1374 -1225 1375 -1223
rect 1381 -1219 1382 -1217
rect 1381 -1225 1382 -1223
rect 1388 -1219 1389 -1217
rect 1388 -1225 1389 -1223
rect 1395 -1219 1396 -1217
rect 1395 -1225 1396 -1223
rect 1402 -1219 1403 -1217
rect 1402 -1225 1403 -1223
rect 1409 -1219 1410 -1217
rect 1409 -1225 1410 -1223
rect 1416 -1219 1417 -1217
rect 1416 -1225 1417 -1223
rect 1423 -1219 1424 -1217
rect 1423 -1225 1424 -1223
rect 1430 -1219 1431 -1217
rect 1430 -1225 1431 -1223
rect 1437 -1219 1438 -1217
rect 1437 -1225 1438 -1223
rect 1444 -1219 1445 -1217
rect 1444 -1225 1445 -1223
rect 1451 -1219 1452 -1217
rect 1451 -1225 1452 -1223
rect 1458 -1219 1459 -1217
rect 1458 -1225 1459 -1223
rect 1465 -1219 1466 -1217
rect 1465 -1225 1466 -1223
rect 1472 -1219 1473 -1217
rect 1472 -1225 1473 -1223
rect 1479 -1219 1480 -1217
rect 1479 -1225 1480 -1223
rect 1486 -1219 1487 -1217
rect 1486 -1225 1487 -1223
rect 1493 -1219 1494 -1217
rect 1493 -1225 1494 -1223
rect 1500 -1219 1501 -1217
rect 1500 -1225 1501 -1223
rect 1507 -1219 1508 -1217
rect 1507 -1225 1508 -1223
rect 1514 -1219 1515 -1217
rect 1514 -1225 1515 -1223
rect 1521 -1219 1522 -1217
rect 1521 -1225 1522 -1223
rect 1528 -1219 1529 -1217
rect 1528 -1225 1529 -1223
rect 1535 -1219 1536 -1217
rect 1535 -1225 1536 -1223
rect 1542 -1219 1543 -1217
rect 1542 -1225 1543 -1223
rect 1549 -1219 1550 -1217
rect 1549 -1225 1550 -1223
rect 1556 -1219 1557 -1217
rect 1556 -1225 1557 -1223
rect 1563 -1219 1564 -1217
rect 1563 -1225 1564 -1223
rect 1570 -1219 1571 -1217
rect 1570 -1225 1571 -1223
rect 1577 -1219 1578 -1217
rect 1577 -1225 1578 -1223
rect 1584 -1219 1585 -1217
rect 1584 -1225 1585 -1223
rect 1591 -1219 1592 -1217
rect 1591 -1225 1592 -1223
rect 1598 -1219 1599 -1217
rect 1598 -1225 1599 -1223
rect 1605 -1219 1606 -1217
rect 1605 -1225 1606 -1223
rect 1612 -1219 1613 -1217
rect 1612 -1225 1613 -1223
rect 1619 -1219 1620 -1217
rect 1619 -1225 1620 -1223
rect 1626 -1219 1627 -1217
rect 1626 -1225 1627 -1223
rect 1633 -1219 1634 -1217
rect 1633 -1225 1634 -1223
rect 1640 -1219 1641 -1217
rect 1640 -1225 1641 -1223
rect 1647 -1219 1648 -1217
rect 1647 -1225 1648 -1223
rect 1654 -1219 1655 -1217
rect 1654 -1225 1655 -1223
rect 1661 -1219 1662 -1217
rect 1661 -1225 1662 -1223
rect 1668 -1219 1669 -1217
rect 1668 -1225 1669 -1223
rect 1675 -1219 1676 -1217
rect 1675 -1225 1676 -1223
rect 1682 -1219 1683 -1217
rect 1682 -1225 1683 -1223
rect 1689 -1219 1690 -1217
rect 1689 -1225 1690 -1223
rect 1696 -1219 1697 -1217
rect 1696 -1225 1697 -1223
rect 1703 -1219 1704 -1217
rect 1703 -1225 1704 -1223
rect 1710 -1219 1711 -1217
rect 1710 -1225 1711 -1223
rect 1717 -1219 1718 -1217
rect 1717 -1225 1718 -1223
rect 1724 -1219 1725 -1217
rect 1724 -1225 1725 -1223
rect 1731 -1219 1732 -1217
rect 1731 -1225 1732 -1223
rect 1738 -1219 1739 -1217
rect 1738 -1225 1739 -1223
rect 1745 -1219 1746 -1217
rect 1748 -1219 1749 -1217
rect 1745 -1225 1746 -1223
rect 1748 -1225 1749 -1223
rect 1752 -1219 1753 -1217
rect 1752 -1225 1753 -1223
rect 1759 -1219 1760 -1217
rect 1759 -1225 1760 -1223
rect 1766 -1219 1767 -1217
rect 1769 -1219 1770 -1217
rect 1766 -1225 1767 -1223
rect 1769 -1225 1770 -1223
rect 1776 -1225 1777 -1223
rect 1780 -1219 1781 -1217
rect 1780 -1225 1781 -1223
rect 1787 -1219 1788 -1217
rect 1787 -1225 1788 -1223
rect 16 -1362 17 -1360
rect 16 -1368 17 -1366
rect 23 -1362 24 -1360
rect 23 -1368 24 -1366
rect 30 -1362 31 -1360
rect 30 -1368 31 -1366
rect 44 -1362 45 -1360
rect 44 -1368 45 -1366
rect 54 -1362 55 -1360
rect 51 -1368 52 -1366
rect 54 -1368 55 -1366
rect 58 -1362 59 -1360
rect 61 -1362 62 -1360
rect 61 -1368 62 -1366
rect 65 -1362 66 -1360
rect 65 -1368 66 -1366
rect 72 -1362 73 -1360
rect 72 -1368 73 -1366
rect 82 -1362 83 -1360
rect 79 -1368 80 -1366
rect 82 -1368 83 -1366
rect 86 -1362 87 -1360
rect 86 -1368 87 -1366
rect 93 -1362 94 -1360
rect 93 -1368 94 -1366
rect 100 -1362 101 -1360
rect 103 -1362 104 -1360
rect 100 -1368 101 -1366
rect 103 -1368 104 -1366
rect 110 -1368 111 -1366
rect 114 -1362 115 -1360
rect 114 -1368 115 -1366
rect 121 -1362 122 -1360
rect 121 -1368 122 -1366
rect 128 -1368 129 -1366
rect 131 -1368 132 -1366
rect 135 -1362 136 -1360
rect 135 -1368 136 -1366
rect 142 -1362 143 -1360
rect 142 -1368 143 -1366
rect 149 -1362 150 -1360
rect 149 -1368 150 -1366
rect 156 -1362 157 -1360
rect 156 -1368 157 -1366
rect 163 -1362 164 -1360
rect 163 -1368 164 -1366
rect 170 -1362 171 -1360
rect 170 -1368 171 -1366
rect 177 -1362 178 -1360
rect 177 -1368 178 -1366
rect 184 -1362 185 -1360
rect 187 -1362 188 -1360
rect 191 -1362 192 -1360
rect 191 -1368 192 -1366
rect 198 -1362 199 -1360
rect 198 -1368 199 -1366
rect 201 -1368 202 -1366
rect 205 -1362 206 -1360
rect 208 -1362 209 -1360
rect 205 -1368 206 -1366
rect 208 -1368 209 -1366
rect 212 -1362 213 -1360
rect 212 -1368 213 -1366
rect 222 -1362 223 -1360
rect 219 -1368 220 -1366
rect 222 -1368 223 -1366
rect 226 -1362 227 -1360
rect 226 -1368 227 -1366
rect 233 -1362 234 -1360
rect 233 -1368 234 -1366
rect 240 -1362 241 -1360
rect 240 -1368 241 -1366
rect 247 -1362 248 -1360
rect 247 -1368 248 -1366
rect 254 -1362 255 -1360
rect 254 -1368 255 -1366
rect 261 -1362 262 -1360
rect 261 -1368 262 -1366
rect 268 -1362 269 -1360
rect 268 -1368 269 -1366
rect 275 -1362 276 -1360
rect 275 -1368 276 -1366
rect 282 -1362 283 -1360
rect 282 -1368 283 -1366
rect 292 -1362 293 -1360
rect 292 -1368 293 -1366
rect 296 -1362 297 -1360
rect 296 -1368 297 -1366
rect 303 -1362 304 -1360
rect 303 -1368 304 -1366
rect 310 -1362 311 -1360
rect 310 -1368 311 -1366
rect 317 -1362 318 -1360
rect 317 -1368 318 -1366
rect 324 -1362 325 -1360
rect 324 -1368 325 -1366
rect 331 -1362 332 -1360
rect 331 -1368 332 -1366
rect 338 -1362 339 -1360
rect 338 -1368 339 -1366
rect 345 -1362 346 -1360
rect 345 -1368 346 -1366
rect 352 -1362 353 -1360
rect 352 -1368 353 -1366
rect 359 -1362 360 -1360
rect 359 -1368 360 -1366
rect 366 -1362 367 -1360
rect 366 -1368 367 -1366
rect 373 -1362 374 -1360
rect 373 -1368 374 -1366
rect 380 -1362 381 -1360
rect 380 -1368 381 -1366
rect 387 -1362 388 -1360
rect 387 -1368 388 -1366
rect 394 -1362 395 -1360
rect 394 -1368 395 -1366
rect 401 -1362 402 -1360
rect 401 -1368 402 -1366
rect 408 -1362 409 -1360
rect 408 -1368 409 -1366
rect 415 -1362 416 -1360
rect 415 -1368 416 -1366
rect 422 -1362 423 -1360
rect 422 -1368 423 -1366
rect 429 -1362 430 -1360
rect 429 -1368 430 -1366
rect 436 -1362 437 -1360
rect 436 -1368 437 -1366
rect 446 -1362 447 -1360
rect 443 -1368 444 -1366
rect 450 -1362 451 -1360
rect 453 -1362 454 -1360
rect 453 -1368 454 -1366
rect 457 -1362 458 -1360
rect 457 -1368 458 -1366
rect 464 -1362 465 -1360
rect 464 -1368 465 -1366
rect 471 -1362 472 -1360
rect 471 -1368 472 -1366
rect 478 -1362 479 -1360
rect 478 -1368 479 -1366
rect 485 -1362 486 -1360
rect 485 -1368 486 -1366
rect 492 -1362 493 -1360
rect 492 -1368 493 -1366
rect 499 -1362 500 -1360
rect 499 -1368 500 -1366
rect 506 -1362 507 -1360
rect 506 -1368 507 -1366
rect 513 -1362 514 -1360
rect 513 -1368 514 -1366
rect 520 -1362 521 -1360
rect 520 -1368 521 -1366
rect 527 -1362 528 -1360
rect 527 -1368 528 -1366
rect 534 -1362 535 -1360
rect 534 -1368 535 -1366
rect 541 -1362 542 -1360
rect 541 -1368 542 -1366
rect 548 -1362 549 -1360
rect 551 -1362 552 -1360
rect 548 -1368 549 -1366
rect 551 -1368 552 -1366
rect 555 -1362 556 -1360
rect 558 -1362 559 -1360
rect 555 -1368 556 -1366
rect 558 -1368 559 -1366
rect 562 -1362 563 -1360
rect 565 -1362 566 -1360
rect 562 -1368 563 -1366
rect 569 -1362 570 -1360
rect 572 -1362 573 -1360
rect 569 -1368 570 -1366
rect 572 -1368 573 -1366
rect 576 -1362 577 -1360
rect 576 -1368 577 -1366
rect 583 -1362 584 -1360
rect 583 -1368 584 -1366
rect 590 -1362 591 -1360
rect 590 -1368 591 -1366
rect 597 -1362 598 -1360
rect 600 -1362 601 -1360
rect 597 -1368 598 -1366
rect 604 -1362 605 -1360
rect 604 -1368 605 -1366
rect 611 -1362 612 -1360
rect 611 -1368 612 -1366
rect 618 -1362 619 -1360
rect 618 -1368 619 -1366
rect 625 -1362 626 -1360
rect 625 -1368 626 -1366
rect 632 -1362 633 -1360
rect 632 -1368 633 -1366
rect 639 -1362 640 -1360
rect 639 -1368 640 -1366
rect 646 -1362 647 -1360
rect 646 -1368 647 -1366
rect 653 -1362 654 -1360
rect 653 -1368 654 -1366
rect 660 -1362 661 -1360
rect 660 -1368 661 -1366
rect 667 -1362 668 -1360
rect 667 -1368 668 -1366
rect 674 -1362 675 -1360
rect 674 -1368 675 -1366
rect 681 -1362 682 -1360
rect 681 -1368 682 -1366
rect 688 -1362 689 -1360
rect 688 -1368 689 -1366
rect 695 -1362 696 -1360
rect 695 -1368 696 -1366
rect 702 -1362 703 -1360
rect 702 -1368 703 -1366
rect 709 -1362 710 -1360
rect 709 -1368 710 -1366
rect 716 -1362 717 -1360
rect 716 -1368 717 -1366
rect 723 -1362 724 -1360
rect 723 -1368 724 -1366
rect 730 -1362 731 -1360
rect 730 -1368 731 -1366
rect 737 -1362 738 -1360
rect 740 -1362 741 -1360
rect 737 -1368 738 -1366
rect 740 -1368 741 -1366
rect 744 -1362 745 -1360
rect 744 -1368 745 -1366
rect 751 -1362 752 -1360
rect 754 -1362 755 -1360
rect 751 -1368 752 -1366
rect 754 -1368 755 -1366
rect 758 -1362 759 -1360
rect 758 -1368 759 -1366
rect 765 -1362 766 -1360
rect 765 -1368 766 -1366
rect 772 -1362 773 -1360
rect 772 -1368 773 -1366
rect 779 -1362 780 -1360
rect 779 -1368 780 -1366
rect 786 -1362 787 -1360
rect 789 -1362 790 -1360
rect 789 -1368 790 -1366
rect 793 -1362 794 -1360
rect 793 -1368 794 -1366
rect 800 -1362 801 -1360
rect 800 -1368 801 -1366
rect 807 -1362 808 -1360
rect 807 -1368 808 -1366
rect 814 -1362 815 -1360
rect 817 -1362 818 -1360
rect 814 -1368 815 -1366
rect 817 -1368 818 -1366
rect 821 -1362 822 -1360
rect 824 -1362 825 -1360
rect 824 -1368 825 -1366
rect 831 -1362 832 -1360
rect 828 -1368 829 -1366
rect 835 -1362 836 -1360
rect 835 -1368 836 -1366
rect 842 -1362 843 -1360
rect 842 -1368 843 -1366
rect 849 -1362 850 -1360
rect 852 -1362 853 -1360
rect 849 -1368 850 -1366
rect 852 -1368 853 -1366
rect 856 -1362 857 -1360
rect 856 -1368 857 -1366
rect 863 -1362 864 -1360
rect 863 -1368 864 -1366
rect 870 -1362 871 -1360
rect 870 -1368 871 -1366
rect 877 -1362 878 -1360
rect 877 -1368 878 -1366
rect 884 -1362 885 -1360
rect 884 -1368 885 -1366
rect 891 -1362 892 -1360
rect 891 -1368 892 -1366
rect 898 -1362 899 -1360
rect 898 -1368 899 -1366
rect 905 -1362 906 -1360
rect 905 -1368 906 -1366
rect 912 -1362 913 -1360
rect 912 -1368 913 -1366
rect 922 -1362 923 -1360
rect 919 -1368 920 -1366
rect 922 -1368 923 -1366
rect 926 -1362 927 -1360
rect 926 -1368 927 -1366
rect 933 -1362 934 -1360
rect 936 -1362 937 -1360
rect 933 -1368 934 -1366
rect 936 -1368 937 -1366
rect 940 -1362 941 -1360
rect 940 -1368 941 -1366
rect 947 -1362 948 -1360
rect 950 -1362 951 -1360
rect 947 -1368 948 -1366
rect 950 -1368 951 -1366
rect 954 -1362 955 -1360
rect 954 -1368 955 -1366
rect 961 -1362 962 -1360
rect 961 -1368 962 -1366
rect 968 -1362 969 -1360
rect 968 -1368 969 -1366
rect 975 -1362 976 -1360
rect 975 -1368 976 -1366
rect 982 -1362 983 -1360
rect 982 -1368 983 -1366
rect 985 -1368 986 -1366
rect 989 -1362 990 -1360
rect 989 -1368 990 -1366
rect 996 -1362 997 -1360
rect 996 -1368 997 -1366
rect 1003 -1362 1004 -1360
rect 1006 -1362 1007 -1360
rect 1006 -1368 1007 -1366
rect 1010 -1362 1011 -1360
rect 1010 -1368 1011 -1366
rect 1020 -1362 1021 -1360
rect 1017 -1368 1018 -1366
rect 1020 -1368 1021 -1366
rect 1024 -1362 1025 -1360
rect 1024 -1368 1025 -1366
rect 1031 -1362 1032 -1360
rect 1031 -1368 1032 -1366
rect 1038 -1362 1039 -1360
rect 1038 -1368 1039 -1366
rect 1045 -1362 1046 -1360
rect 1045 -1368 1046 -1366
rect 1052 -1362 1053 -1360
rect 1052 -1368 1053 -1366
rect 1059 -1362 1060 -1360
rect 1059 -1368 1060 -1366
rect 1066 -1362 1067 -1360
rect 1066 -1368 1067 -1366
rect 1073 -1362 1074 -1360
rect 1073 -1368 1074 -1366
rect 1080 -1362 1081 -1360
rect 1080 -1368 1081 -1366
rect 1087 -1362 1088 -1360
rect 1087 -1368 1088 -1366
rect 1094 -1362 1095 -1360
rect 1094 -1368 1095 -1366
rect 1101 -1362 1102 -1360
rect 1104 -1362 1105 -1360
rect 1101 -1368 1102 -1366
rect 1104 -1368 1105 -1366
rect 1108 -1362 1109 -1360
rect 1108 -1368 1109 -1366
rect 1115 -1362 1116 -1360
rect 1115 -1368 1116 -1366
rect 1122 -1362 1123 -1360
rect 1122 -1368 1123 -1366
rect 1129 -1362 1130 -1360
rect 1129 -1368 1130 -1366
rect 1136 -1362 1137 -1360
rect 1136 -1368 1137 -1366
rect 1146 -1362 1147 -1360
rect 1143 -1368 1144 -1366
rect 1146 -1368 1147 -1366
rect 1150 -1362 1151 -1360
rect 1150 -1368 1151 -1366
rect 1157 -1362 1158 -1360
rect 1157 -1368 1158 -1366
rect 1164 -1362 1165 -1360
rect 1164 -1368 1165 -1366
rect 1171 -1362 1172 -1360
rect 1171 -1368 1172 -1366
rect 1178 -1362 1179 -1360
rect 1178 -1368 1179 -1366
rect 1185 -1362 1186 -1360
rect 1185 -1368 1186 -1366
rect 1192 -1362 1193 -1360
rect 1192 -1368 1193 -1366
rect 1199 -1362 1200 -1360
rect 1202 -1362 1203 -1360
rect 1202 -1368 1203 -1366
rect 1206 -1362 1207 -1360
rect 1206 -1368 1207 -1366
rect 1213 -1362 1214 -1360
rect 1213 -1368 1214 -1366
rect 1216 -1368 1217 -1366
rect 1220 -1362 1221 -1360
rect 1220 -1368 1221 -1366
rect 1227 -1362 1228 -1360
rect 1227 -1368 1228 -1366
rect 1234 -1362 1235 -1360
rect 1234 -1368 1235 -1366
rect 1241 -1362 1242 -1360
rect 1241 -1368 1242 -1366
rect 1248 -1362 1249 -1360
rect 1248 -1368 1249 -1366
rect 1255 -1362 1256 -1360
rect 1255 -1368 1256 -1366
rect 1262 -1362 1263 -1360
rect 1262 -1368 1263 -1366
rect 1269 -1362 1270 -1360
rect 1269 -1368 1270 -1366
rect 1276 -1362 1277 -1360
rect 1276 -1368 1277 -1366
rect 1283 -1362 1284 -1360
rect 1283 -1368 1284 -1366
rect 1290 -1362 1291 -1360
rect 1290 -1368 1291 -1366
rect 1297 -1362 1298 -1360
rect 1297 -1368 1298 -1366
rect 1304 -1368 1305 -1366
rect 1311 -1362 1312 -1360
rect 1314 -1362 1315 -1360
rect 1311 -1368 1312 -1366
rect 1318 -1362 1319 -1360
rect 1318 -1368 1319 -1366
rect 1325 -1362 1326 -1360
rect 1325 -1368 1326 -1366
rect 1332 -1362 1333 -1360
rect 1332 -1368 1333 -1366
rect 1339 -1362 1340 -1360
rect 1339 -1368 1340 -1366
rect 1346 -1362 1347 -1360
rect 1346 -1368 1347 -1366
rect 1353 -1362 1354 -1360
rect 1353 -1368 1354 -1366
rect 1360 -1362 1361 -1360
rect 1360 -1368 1361 -1366
rect 1367 -1362 1368 -1360
rect 1367 -1368 1368 -1366
rect 1374 -1362 1375 -1360
rect 1374 -1368 1375 -1366
rect 1381 -1362 1382 -1360
rect 1381 -1368 1382 -1366
rect 1388 -1362 1389 -1360
rect 1388 -1368 1389 -1366
rect 1395 -1362 1396 -1360
rect 1395 -1368 1396 -1366
rect 1402 -1362 1403 -1360
rect 1402 -1368 1403 -1366
rect 1409 -1362 1410 -1360
rect 1409 -1368 1410 -1366
rect 1416 -1362 1417 -1360
rect 1416 -1368 1417 -1366
rect 1423 -1362 1424 -1360
rect 1423 -1368 1424 -1366
rect 1430 -1362 1431 -1360
rect 1430 -1368 1431 -1366
rect 1437 -1362 1438 -1360
rect 1437 -1368 1438 -1366
rect 1444 -1362 1445 -1360
rect 1444 -1368 1445 -1366
rect 1451 -1362 1452 -1360
rect 1451 -1368 1452 -1366
rect 1458 -1362 1459 -1360
rect 1458 -1368 1459 -1366
rect 1465 -1362 1466 -1360
rect 1465 -1368 1466 -1366
rect 1472 -1362 1473 -1360
rect 1472 -1368 1473 -1366
rect 1479 -1362 1480 -1360
rect 1479 -1368 1480 -1366
rect 1486 -1362 1487 -1360
rect 1486 -1368 1487 -1366
rect 1493 -1362 1494 -1360
rect 1493 -1368 1494 -1366
rect 1500 -1362 1501 -1360
rect 1500 -1368 1501 -1366
rect 1507 -1362 1508 -1360
rect 1507 -1368 1508 -1366
rect 1514 -1362 1515 -1360
rect 1514 -1368 1515 -1366
rect 1521 -1362 1522 -1360
rect 1521 -1368 1522 -1366
rect 1528 -1362 1529 -1360
rect 1528 -1368 1529 -1366
rect 1535 -1362 1536 -1360
rect 1535 -1368 1536 -1366
rect 1542 -1362 1543 -1360
rect 1542 -1368 1543 -1366
rect 1549 -1362 1550 -1360
rect 1549 -1368 1550 -1366
rect 1556 -1362 1557 -1360
rect 1556 -1368 1557 -1366
rect 1563 -1362 1564 -1360
rect 1563 -1368 1564 -1366
rect 1570 -1362 1571 -1360
rect 1570 -1368 1571 -1366
rect 1577 -1362 1578 -1360
rect 1577 -1368 1578 -1366
rect 1584 -1362 1585 -1360
rect 1584 -1368 1585 -1366
rect 1591 -1362 1592 -1360
rect 1591 -1368 1592 -1366
rect 1598 -1362 1599 -1360
rect 1598 -1368 1599 -1366
rect 1605 -1362 1606 -1360
rect 1605 -1368 1606 -1366
rect 1612 -1362 1613 -1360
rect 1612 -1368 1613 -1366
rect 1619 -1362 1620 -1360
rect 1619 -1368 1620 -1366
rect 1626 -1362 1627 -1360
rect 1626 -1368 1627 -1366
rect 1633 -1362 1634 -1360
rect 1633 -1368 1634 -1366
rect 1640 -1362 1641 -1360
rect 1640 -1368 1641 -1366
rect 1647 -1362 1648 -1360
rect 1647 -1368 1648 -1366
rect 1654 -1362 1655 -1360
rect 1654 -1368 1655 -1366
rect 1661 -1362 1662 -1360
rect 1661 -1368 1662 -1366
rect 1668 -1362 1669 -1360
rect 1668 -1368 1669 -1366
rect 1675 -1362 1676 -1360
rect 1675 -1368 1676 -1366
rect 1682 -1362 1683 -1360
rect 1682 -1368 1683 -1366
rect 1689 -1362 1690 -1360
rect 1689 -1368 1690 -1366
rect 1696 -1362 1697 -1360
rect 1696 -1368 1697 -1366
rect 1703 -1362 1704 -1360
rect 1703 -1368 1704 -1366
rect 1710 -1362 1711 -1360
rect 1710 -1368 1711 -1366
rect 1717 -1362 1718 -1360
rect 1717 -1368 1718 -1366
rect 1724 -1362 1725 -1360
rect 1724 -1368 1725 -1366
rect 1731 -1362 1732 -1360
rect 1731 -1368 1732 -1366
rect 1738 -1362 1739 -1360
rect 1738 -1368 1739 -1366
rect 1745 -1362 1746 -1360
rect 1745 -1368 1746 -1366
rect 1752 -1362 1753 -1360
rect 1752 -1368 1753 -1366
rect 23 -1503 24 -1501
rect 23 -1509 24 -1507
rect 30 -1503 31 -1501
rect 30 -1509 31 -1507
rect 37 -1503 38 -1501
rect 37 -1509 38 -1507
rect 44 -1503 45 -1501
rect 44 -1509 45 -1507
rect 51 -1503 52 -1501
rect 51 -1509 52 -1507
rect 58 -1503 59 -1501
rect 58 -1509 59 -1507
rect 65 -1509 66 -1507
rect 68 -1509 69 -1507
rect 72 -1503 73 -1501
rect 72 -1509 73 -1507
rect 79 -1503 80 -1501
rect 79 -1509 80 -1507
rect 86 -1503 87 -1501
rect 86 -1509 87 -1507
rect 93 -1503 94 -1501
rect 93 -1509 94 -1507
rect 100 -1503 101 -1501
rect 100 -1509 101 -1507
rect 107 -1503 108 -1501
rect 107 -1509 108 -1507
rect 114 -1503 115 -1501
rect 114 -1509 115 -1507
rect 124 -1503 125 -1501
rect 121 -1509 122 -1507
rect 124 -1509 125 -1507
rect 128 -1503 129 -1501
rect 131 -1503 132 -1501
rect 128 -1509 129 -1507
rect 131 -1509 132 -1507
rect 135 -1503 136 -1501
rect 135 -1509 136 -1507
rect 142 -1503 143 -1501
rect 142 -1509 143 -1507
rect 149 -1503 150 -1501
rect 149 -1509 150 -1507
rect 156 -1503 157 -1501
rect 159 -1503 160 -1501
rect 156 -1509 157 -1507
rect 159 -1509 160 -1507
rect 163 -1503 164 -1501
rect 163 -1509 164 -1507
rect 170 -1503 171 -1501
rect 170 -1509 171 -1507
rect 177 -1503 178 -1501
rect 177 -1509 178 -1507
rect 184 -1503 185 -1501
rect 187 -1503 188 -1501
rect 184 -1509 185 -1507
rect 191 -1503 192 -1501
rect 194 -1503 195 -1501
rect 191 -1509 192 -1507
rect 194 -1509 195 -1507
rect 198 -1503 199 -1501
rect 198 -1509 199 -1507
rect 205 -1503 206 -1501
rect 205 -1509 206 -1507
rect 212 -1503 213 -1501
rect 215 -1503 216 -1501
rect 212 -1509 213 -1507
rect 215 -1509 216 -1507
rect 219 -1503 220 -1501
rect 219 -1509 220 -1507
rect 226 -1503 227 -1501
rect 229 -1503 230 -1501
rect 226 -1509 227 -1507
rect 229 -1509 230 -1507
rect 233 -1503 234 -1501
rect 233 -1509 234 -1507
rect 240 -1503 241 -1501
rect 240 -1509 241 -1507
rect 247 -1503 248 -1501
rect 247 -1509 248 -1507
rect 254 -1503 255 -1501
rect 257 -1503 258 -1501
rect 254 -1509 255 -1507
rect 261 -1503 262 -1501
rect 261 -1509 262 -1507
rect 268 -1503 269 -1501
rect 268 -1509 269 -1507
rect 275 -1503 276 -1501
rect 275 -1509 276 -1507
rect 282 -1503 283 -1501
rect 282 -1509 283 -1507
rect 289 -1503 290 -1501
rect 289 -1509 290 -1507
rect 296 -1503 297 -1501
rect 296 -1509 297 -1507
rect 303 -1503 304 -1501
rect 303 -1509 304 -1507
rect 310 -1503 311 -1501
rect 310 -1509 311 -1507
rect 320 -1509 321 -1507
rect 324 -1503 325 -1501
rect 324 -1509 325 -1507
rect 331 -1503 332 -1501
rect 331 -1509 332 -1507
rect 338 -1503 339 -1501
rect 338 -1509 339 -1507
rect 345 -1503 346 -1501
rect 345 -1509 346 -1507
rect 352 -1503 353 -1501
rect 352 -1509 353 -1507
rect 359 -1503 360 -1501
rect 359 -1509 360 -1507
rect 366 -1503 367 -1501
rect 366 -1509 367 -1507
rect 373 -1503 374 -1501
rect 373 -1509 374 -1507
rect 380 -1503 381 -1501
rect 380 -1509 381 -1507
rect 387 -1503 388 -1501
rect 387 -1509 388 -1507
rect 394 -1503 395 -1501
rect 394 -1509 395 -1507
rect 401 -1503 402 -1501
rect 401 -1509 402 -1507
rect 408 -1503 409 -1501
rect 408 -1509 409 -1507
rect 415 -1503 416 -1501
rect 415 -1509 416 -1507
rect 418 -1509 419 -1507
rect 422 -1503 423 -1501
rect 422 -1509 423 -1507
rect 429 -1503 430 -1501
rect 429 -1509 430 -1507
rect 436 -1503 437 -1501
rect 436 -1509 437 -1507
rect 443 -1503 444 -1501
rect 443 -1509 444 -1507
rect 450 -1503 451 -1501
rect 450 -1509 451 -1507
rect 457 -1503 458 -1501
rect 460 -1503 461 -1501
rect 457 -1509 458 -1507
rect 460 -1509 461 -1507
rect 464 -1503 465 -1501
rect 464 -1509 465 -1507
rect 471 -1503 472 -1501
rect 471 -1509 472 -1507
rect 478 -1503 479 -1501
rect 481 -1503 482 -1501
rect 478 -1509 479 -1507
rect 481 -1509 482 -1507
rect 485 -1503 486 -1501
rect 492 -1503 493 -1501
rect 492 -1509 493 -1507
rect 499 -1503 500 -1501
rect 499 -1509 500 -1507
rect 506 -1503 507 -1501
rect 506 -1509 507 -1507
rect 513 -1503 514 -1501
rect 516 -1503 517 -1501
rect 513 -1509 514 -1507
rect 520 -1503 521 -1501
rect 520 -1509 521 -1507
rect 527 -1503 528 -1501
rect 527 -1509 528 -1507
rect 534 -1503 535 -1501
rect 534 -1509 535 -1507
rect 541 -1503 542 -1501
rect 541 -1509 542 -1507
rect 548 -1503 549 -1501
rect 548 -1509 549 -1507
rect 555 -1503 556 -1501
rect 555 -1509 556 -1507
rect 562 -1503 563 -1501
rect 562 -1509 563 -1507
rect 569 -1503 570 -1501
rect 569 -1509 570 -1507
rect 576 -1503 577 -1501
rect 576 -1509 577 -1507
rect 583 -1503 584 -1501
rect 583 -1509 584 -1507
rect 590 -1503 591 -1501
rect 590 -1509 591 -1507
rect 597 -1503 598 -1501
rect 597 -1509 598 -1507
rect 604 -1503 605 -1501
rect 604 -1509 605 -1507
rect 611 -1503 612 -1501
rect 611 -1509 612 -1507
rect 618 -1503 619 -1501
rect 618 -1509 619 -1507
rect 625 -1509 626 -1507
rect 628 -1509 629 -1507
rect 632 -1503 633 -1501
rect 632 -1509 633 -1507
rect 639 -1503 640 -1501
rect 639 -1509 640 -1507
rect 646 -1503 647 -1501
rect 646 -1509 647 -1507
rect 653 -1503 654 -1501
rect 653 -1509 654 -1507
rect 656 -1509 657 -1507
rect 660 -1503 661 -1501
rect 660 -1509 661 -1507
rect 670 -1503 671 -1501
rect 667 -1509 668 -1507
rect 670 -1509 671 -1507
rect 674 -1503 675 -1501
rect 674 -1509 675 -1507
rect 681 -1503 682 -1501
rect 681 -1509 682 -1507
rect 688 -1503 689 -1501
rect 688 -1509 689 -1507
rect 695 -1503 696 -1501
rect 695 -1509 696 -1507
rect 702 -1503 703 -1501
rect 702 -1509 703 -1507
rect 709 -1503 710 -1501
rect 709 -1509 710 -1507
rect 716 -1503 717 -1501
rect 719 -1503 720 -1501
rect 716 -1509 717 -1507
rect 726 -1503 727 -1501
rect 726 -1509 727 -1507
rect 730 -1503 731 -1501
rect 730 -1509 731 -1507
rect 737 -1503 738 -1501
rect 740 -1503 741 -1501
rect 737 -1509 738 -1507
rect 740 -1509 741 -1507
rect 744 -1503 745 -1501
rect 744 -1509 745 -1507
rect 751 -1503 752 -1501
rect 751 -1509 752 -1507
rect 758 -1503 759 -1501
rect 761 -1503 762 -1501
rect 758 -1509 759 -1507
rect 761 -1509 762 -1507
rect 765 -1503 766 -1501
rect 765 -1509 766 -1507
rect 772 -1503 773 -1501
rect 772 -1509 773 -1507
rect 779 -1503 780 -1501
rect 779 -1509 780 -1507
rect 786 -1503 787 -1501
rect 786 -1509 787 -1507
rect 789 -1509 790 -1507
rect 793 -1503 794 -1501
rect 793 -1509 794 -1507
rect 800 -1503 801 -1501
rect 800 -1509 801 -1507
rect 807 -1503 808 -1501
rect 807 -1509 808 -1507
rect 814 -1503 815 -1501
rect 814 -1509 815 -1507
rect 821 -1503 822 -1501
rect 824 -1503 825 -1501
rect 821 -1509 822 -1507
rect 824 -1509 825 -1507
rect 828 -1503 829 -1501
rect 831 -1503 832 -1501
rect 831 -1509 832 -1507
rect 835 -1503 836 -1501
rect 835 -1509 836 -1507
rect 842 -1503 843 -1501
rect 842 -1509 843 -1507
rect 849 -1503 850 -1501
rect 849 -1509 850 -1507
rect 856 -1503 857 -1501
rect 856 -1509 857 -1507
rect 863 -1503 864 -1501
rect 866 -1503 867 -1501
rect 863 -1509 864 -1507
rect 866 -1509 867 -1507
rect 870 -1503 871 -1501
rect 870 -1509 871 -1507
rect 877 -1503 878 -1501
rect 877 -1509 878 -1507
rect 884 -1503 885 -1501
rect 884 -1509 885 -1507
rect 891 -1503 892 -1501
rect 891 -1509 892 -1507
rect 898 -1503 899 -1501
rect 898 -1509 899 -1507
rect 905 -1503 906 -1501
rect 905 -1509 906 -1507
rect 912 -1503 913 -1501
rect 912 -1509 913 -1507
rect 919 -1503 920 -1501
rect 919 -1509 920 -1507
rect 926 -1503 927 -1501
rect 926 -1509 927 -1507
rect 933 -1503 934 -1501
rect 936 -1503 937 -1501
rect 933 -1509 934 -1507
rect 936 -1509 937 -1507
rect 940 -1503 941 -1501
rect 940 -1509 941 -1507
rect 947 -1503 948 -1501
rect 950 -1503 951 -1501
rect 947 -1509 948 -1507
rect 950 -1509 951 -1507
rect 954 -1503 955 -1501
rect 954 -1509 955 -1507
rect 961 -1503 962 -1501
rect 961 -1509 962 -1507
rect 968 -1503 969 -1501
rect 968 -1509 969 -1507
rect 978 -1503 979 -1501
rect 975 -1509 976 -1507
rect 978 -1509 979 -1507
rect 982 -1503 983 -1501
rect 982 -1509 983 -1507
rect 989 -1503 990 -1501
rect 989 -1509 990 -1507
rect 996 -1503 997 -1501
rect 996 -1509 997 -1507
rect 1003 -1503 1004 -1501
rect 1003 -1509 1004 -1507
rect 1010 -1503 1011 -1501
rect 1010 -1509 1011 -1507
rect 1017 -1503 1018 -1501
rect 1017 -1509 1018 -1507
rect 1024 -1503 1025 -1501
rect 1024 -1509 1025 -1507
rect 1031 -1503 1032 -1501
rect 1034 -1503 1035 -1501
rect 1031 -1509 1032 -1507
rect 1034 -1509 1035 -1507
rect 1038 -1503 1039 -1501
rect 1038 -1509 1039 -1507
rect 1045 -1503 1046 -1501
rect 1048 -1503 1049 -1501
rect 1048 -1509 1049 -1507
rect 1052 -1503 1053 -1501
rect 1052 -1509 1053 -1507
rect 1059 -1503 1060 -1501
rect 1059 -1509 1060 -1507
rect 1066 -1503 1067 -1501
rect 1066 -1509 1067 -1507
rect 1073 -1503 1074 -1501
rect 1073 -1509 1074 -1507
rect 1080 -1503 1081 -1501
rect 1080 -1509 1081 -1507
rect 1087 -1503 1088 -1501
rect 1087 -1509 1088 -1507
rect 1094 -1503 1095 -1501
rect 1094 -1509 1095 -1507
rect 1101 -1503 1102 -1501
rect 1101 -1509 1102 -1507
rect 1108 -1503 1109 -1501
rect 1108 -1509 1109 -1507
rect 1115 -1503 1116 -1501
rect 1115 -1509 1116 -1507
rect 1122 -1503 1123 -1501
rect 1122 -1509 1123 -1507
rect 1129 -1503 1130 -1501
rect 1129 -1509 1130 -1507
rect 1136 -1503 1137 -1501
rect 1136 -1509 1137 -1507
rect 1143 -1503 1144 -1501
rect 1143 -1509 1144 -1507
rect 1150 -1503 1151 -1501
rect 1150 -1509 1151 -1507
rect 1157 -1503 1158 -1501
rect 1157 -1509 1158 -1507
rect 1164 -1503 1165 -1501
rect 1164 -1509 1165 -1507
rect 1171 -1503 1172 -1501
rect 1171 -1509 1172 -1507
rect 1178 -1503 1179 -1501
rect 1178 -1509 1179 -1507
rect 1185 -1503 1186 -1501
rect 1185 -1509 1186 -1507
rect 1192 -1503 1193 -1501
rect 1192 -1509 1193 -1507
rect 1199 -1503 1200 -1501
rect 1199 -1509 1200 -1507
rect 1206 -1503 1207 -1501
rect 1206 -1509 1207 -1507
rect 1213 -1503 1214 -1501
rect 1213 -1509 1214 -1507
rect 1220 -1503 1221 -1501
rect 1220 -1509 1221 -1507
rect 1227 -1503 1228 -1501
rect 1227 -1509 1228 -1507
rect 1234 -1503 1235 -1501
rect 1234 -1509 1235 -1507
rect 1241 -1503 1242 -1501
rect 1241 -1509 1242 -1507
rect 1248 -1503 1249 -1501
rect 1248 -1509 1249 -1507
rect 1255 -1503 1256 -1501
rect 1255 -1509 1256 -1507
rect 1262 -1503 1263 -1501
rect 1262 -1509 1263 -1507
rect 1269 -1503 1270 -1501
rect 1269 -1509 1270 -1507
rect 1276 -1503 1277 -1501
rect 1276 -1509 1277 -1507
rect 1283 -1503 1284 -1501
rect 1283 -1509 1284 -1507
rect 1290 -1503 1291 -1501
rect 1290 -1509 1291 -1507
rect 1297 -1503 1298 -1501
rect 1297 -1509 1298 -1507
rect 1304 -1503 1305 -1501
rect 1304 -1509 1305 -1507
rect 1311 -1503 1312 -1501
rect 1311 -1509 1312 -1507
rect 1318 -1503 1319 -1501
rect 1318 -1509 1319 -1507
rect 1325 -1503 1326 -1501
rect 1325 -1509 1326 -1507
rect 1332 -1503 1333 -1501
rect 1332 -1509 1333 -1507
rect 1339 -1503 1340 -1501
rect 1339 -1509 1340 -1507
rect 1346 -1503 1347 -1501
rect 1346 -1509 1347 -1507
rect 1353 -1503 1354 -1501
rect 1353 -1509 1354 -1507
rect 1360 -1503 1361 -1501
rect 1360 -1509 1361 -1507
rect 1367 -1503 1368 -1501
rect 1367 -1509 1368 -1507
rect 1374 -1503 1375 -1501
rect 1374 -1509 1375 -1507
rect 1381 -1503 1382 -1501
rect 1381 -1509 1382 -1507
rect 1388 -1503 1389 -1501
rect 1388 -1509 1389 -1507
rect 1395 -1503 1396 -1501
rect 1395 -1509 1396 -1507
rect 1402 -1503 1403 -1501
rect 1402 -1509 1403 -1507
rect 1409 -1503 1410 -1501
rect 1409 -1509 1410 -1507
rect 1416 -1503 1417 -1501
rect 1416 -1509 1417 -1507
rect 1423 -1503 1424 -1501
rect 1423 -1509 1424 -1507
rect 1430 -1503 1431 -1501
rect 1430 -1509 1431 -1507
rect 1437 -1503 1438 -1501
rect 1437 -1509 1438 -1507
rect 1444 -1503 1445 -1501
rect 1444 -1509 1445 -1507
rect 1451 -1503 1452 -1501
rect 1451 -1509 1452 -1507
rect 1454 -1509 1455 -1507
rect 1458 -1503 1459 -1501
rect 1458 -1509 1459 -1507
rect 1465 -1503 1466 -1501
rect 1465 -1509 1466 -1507
rect 1472 -1503 1473 -1501
rect 1472 -1509 1473 -1507
rect 1479 -1503 1480 -1501
rect 1479 -1509 1480 -1507
rect 1486 -1503 1487 -1501
rect 1486 -1509 1487 -1507
rect 1493 -1503 1494 -1501
rect 1493 -1509 1494 -1507
rect 1500 -1503 1501 -1501
rect 1500 -1509 1501 -1507
rect 1507 -1503 1508 -1501
rect 1507 -1509 1508 -1507
rect 1514 -1503 1515 -1501
rect 1514 -1509 1515 -1507
rect 1521 -1503 1522 -1501
rect 1521 -1509 1522 -1507
rect 1528 -1503 1529 -1501
rect 1528 -1509 1529 -1507
rect 1535 -1503 1536 -1501
rect 1538 -1503 1539 -1501
rect 1535 -1509 1536 -1507
rect 1538 -1509 1539 -1507
rect 1542 -1503 1543 -1501
rect 1542 -1509 1543 -1507
rect 1549 -1503 1550 -1501
rect 1552 -1503 1553 -1501
rect 1549 -1509 1550 -1507
rect 1556 -1503 1557 -1501
rect 1556 -1509 1557 -1507
rect 1563 -1503 1564 -1501
rect 1563 -1509 1564 -1507
rect 1570 -1503 1571 -1501
rect 1570 -1509 1571 -1507
rect 1577 -1503 1578 -1501
rect 1577 -1509 1578 -1507
rect 1584 -1503 1585 -1501
rect 1587 -1503 1588 -1501
rect 1584 -1509 1585 -1507
rect 1591 -1503 1592 -1501
rect 1591 -1509 1592 -1507
rect 1598 -1503 1599 -1501
rect 1598 -1509 1599 -1507
rect 1605 -1503 1606 -1501
rect 1608 -1503 1609 -1501
rect 1605 -1509 1606 -1507
rect 1608 -1509 1609 -1507
rect 1612 -1503 1613 -1501
rect 1612 -1509 1613 -1507
rect 1619 -1503 1620 -1501
rect 1619 -1509 1620 -1507
rect 1626 -1503 1627 -1501
rect 1626 -1509 1627 -1507
rect 1633 -1503 1634 -1501
rect 1633 -1509 1634 -1507
rect 1643 -1503 1644 -1501
rect 1640 -1509 1641 -1507
rect 1643 -1509 1644 -1507
rect 1647 -1503 1648 -1501
rect 1647 -1509 1648 -1507
rect 1654 -1503 1655 -1501
rect 1654 -1509 1655 -1507
rect 1661 -1503 1662 -1501
rect 1661 -1509 1662 -1507
rect 1668 -1503 1669 -1501
rect 1668 -1509 1669 -1507
rect 1675 -1503 1676 -1501
rect 1675 -1509 1676 -1507
rect 1682 -1503 1683 -1501
rect 1682 -1509 1683 -1507
rect 1689 -1503 1690 -1501
rect 1689 -1509 1690 -1507
rect 1696 -1503 1697 -1501
rect 1696 -1509 1697 -1507
rect 1703 -1503 1704 -1501
rect 1703 -1509 1704 -1507
rect 1710 -1503 1711 -1501
rect 1710 -1509 1711 -1507
rect 1717 -1503 1718 -1501
rect 1717 -1509 1718 -1507
rect 1724 -1503 1725 -1501
rect 1724 -1509 1725 -1507
rect 1731 -1503 1732 -1501
rect 1731 -1509 1732 -1507
rect 1801 -1503 1802 -1501
rect 1801 -1509 1802 -1507
rect 23 -1638 24 -1636
rect 23 -1644 24 -1642
rect 30 -1638 31 -1636
rect 30 -1644 31 -1642
rect 37 -1638 38 -1636
rect 37 -1644 38 -1642
rect 44 -1638 45 -1636
rect 44 -1644 45 -1642
rect 51 -1638 52 -1636
rect 51 -1644 52 -1642
rect 61 -1638 62 -1636
rect 65 -1638 66 -1636
rect 65 -1644 66 -1642
rect 72 -1638 73 -1636
rect 72 -1644 73 -1642
rect 79 -1638 80 -1636
rect 79 -1644 80 -1642
rect 86 -1638 87 -1636
rect 86 -1644 87 -1642
rect 93 -1638 94 -1636
rect 93 -1644 94 -1642
rect 100 -1638 101 -1636
rect 100 -1644 101 -1642
rect 107 -1638 108 -1636
rect 107 -1644 108 -1642
rect 114 -1638 115 -1636
rect 114 -1644 115 -1642
rect 121 -1638 122 -1636
rect 124 -1638 125 -1636
rect 121 -1644 122 -1642
rect 124 -1644 125 -1642
rect 128 -1638 129 -1636
rect 128 -1644 129 -1642
rect 135 -1638 136 -1636
rect 135 -1644 136 -1642
rect 142 -1638 143 -1636
rect 142 -1644 143 -1642
rect 149 -1638 150 -1636
rect 149 -1644 150 -1642
rect 156 -1638 157 -1636
rect 156 -1644 157 -1642
rect 163 -1638 164 -1636
rect 166 -1638 167 -1636
rect 163 -1644 164 -1642
rect 170 -1638 171 -1636
rect 170 -1644 171 -1642
rect 177 -1638 178 -1636
rect 177 -1644 178 -1642
rect 184 -1638 185 -1636
rect 187 -1638 188 -1636
rect 184 -1644 185 -1642
rect 187 -1644 188 -1642
rect 191 -1638 192 -1636
rect 191 -1644 192 -1642
rect 198 -1638 199 -1636
rect 198 -1644 199 -1642
rect 205 -1638 206 -1636
rect 205 -1644 206 -1642
rect 212 -1638 213 -1636
rect 212 -1644 213 -1642
rect 219 -1638 220 -1636
rect 222 -1638 223 -1636
rect 219 -1644 220 -1642
rect 222 -1644 223 -1642
rect 226 -1638 227 -1636
rect 226 -1644 227 -1642
rect 233 -1638 234 -1636
rect 233 -1644 234 -1642
rect 240 -1638 241 -1636
rect 240 -1644 241 -1642
rect 247 -1638 248 -1636
rect 247 -1644 248 -1642
rect 254 -1638 255 -1636
rect 254 -1644 255 -1642
rect 264 -1638 265 -1636
rect 261 -1644 262 -1642
rect 268 -1638 269 -1636
rect 268 -1644 269 -1642
rect 275 -1638 276 -1636
rect 275 -1644 276 -1642
rect 282 -1638 283 -1636
rect 282 -1644 283 -1642
rect 289 -1638 290 -1636
rect 289 -1644 290 -1642
rect 296 -1638 297 -1636
rect 296 -1644 297 -1642
rect 303 -1638 304 -1636
rect 303 -1644 304 -1642
rect 310 -1638 311 -1636
rect 313 -1638 314 -1636
rect 310 -1644 311 -1642
rect 317 -1638 318 -1636
rect 317 -1644 318 -1642
rect 324 -1638 325 -1636
rect 324 -1644 325 -1642
rect 331 -1638 332 -1636
rect 331 -1644 332 -1642
rect 338 -1638 339 -1636
rect 338 -1644 339 -1642
rect 345 -1638 346 -1636
rect 345 -1644 346 -1642
rect 352 -1638 353 -1636
rect 352 -1644 353 -1642
rect 359 -1638 360 -1636
rect 359 -1644 360 -1642
rect 366 -1638 367 -1636
rect 366 -1644 367 -1642
rect 373 -1638 374 -1636
rect 373 -1644 374 -1642
rect 380 -1638 381 -1636
rect 380 -1644 381 -1642
rect 387 -1638 388 -1636
rect 387 -1644 388 -1642
rect 394 -1638 395 -1636
rect 394 -1644 395 -1642
rect 401 -1638 402 -1636
rect 401 -1644 402 -1642
rect 408 -1638 409 -1636
rect 408 -1644 409 -1642
rect 415 -1638 416 -1636
rect 415 -1644 416 -1642
rect 422 -1638 423 -1636
rect 422 -1644 423 -1642
rect 429 -1638 430 -1636
rect 429 -1644 430 -1642
rect 436 -1638 437 -1636
rect 436 -1644 437 -1642
rect 443 -1638 444 -1636
rect 446 -1638 447 -1636
rect 443 -1644 444 -1642
rect 446 -1644 447 -1642
rect 450 -1638 451 -1636
rect 450 -1644 451 -1642
rect 453 -1644 454 -1642
rect 457 -1638 458 -1636
rect 457 -1644 458 -1642
rect 464 -1638 465 -1636
rect 464 -1644 465 -1642
rect 471 -1638 472 -1636
rect 471 -1644 472 -1642
rect 478 -1638 479 -1636
rect 478 -1644 479 -1642
rect 485 -1644 486 -1642
rect 492 -1638 493 -1636
rect 492 -1644 493 -1642
rect 499 -1638 500 -1636
rect 499 -1644 500 -1642
rect 506 -1638 507 -1636
rect 506 -1644 507 -1642
rect 513 -1638 514 -1636
rect 513 -1644 514 -1642
rect 520 -1638 521 -1636
rect 520 -1644 521 -1642
rect 527 -1638 528 -1636
rect 527 -1644 528 -1642
rect 534 -1638 535 -1636
rect 534 -1644 535 -1642
rect 541 -1638 542 -1636
rect 544 -1638 545 -1636
rect 541 -1644 542 -1642
rect 544 -1644 545 -1642
rect 548 -1638 549 -1636
rect 551 -1638 552 -1636
rect 548 -1644 549 -1642
rect 551 -1644 552 -1642
rect 555 -1638 556 -1636
rect 555 -1644 556 -1642
rect 562 -1638 563 -1636
rect 562 -1644 563 -1642
rect 569 -1638 570 -1636
rect 569 -1644 570 -1642
rect 576 -1638 577 -1636
rect 576 -1644 577 -1642
rect 583 -1638 584 -1636
rect 583 -1644 584 -1642
rect 590 -1638 591 -1636
rect 590 -1644 591 -1642
rect 597 -1638 598 -1636
rect 597 -1644 598 -1642
rect 604 -1638 605 -1636
rect 607 -1638 608 -1636
rect 607 -1644 608 -1642
rect 611 -1638 612 -1636
rect 611 -1644 612 -1642
rect 618 -1638 619 -1636
rect 618 -1644 619 -1642
rect 625 -1638 626 -1636
rect 625 -1644 626 -1642
rect 632 -1638 633 -1636
rect 632 -1644 633 -1642
rect 639 -1638 640 -1636
rect 639 -1644 640 -1642
rect 646 -1638 647 -1636
rect 646 -1644 647 -1642
rect 653 -1638 654 -1636
rect 653 -1644 654 -1642
rect 660 -1638 661 -1636
rect 660 -1644 661 -1642
rect 667 -1638 668 -1636
rect 667 -1644 668 -1642
rect 674 -1638 675 -1636
rect 674 -1644 675 -1642
rect 681 -1638 682 -1636
rect 681 -1644 682 -1642
rect 688 -1638 689 -1636
rect 688 -1644 689 -1642
rect 695 -1638 696 -1636
rect 695 -1644 696 -1642
rect 702 -1638 703 -1636
rect 702 -1644 703 -1642
rect 709 -1638 710 -1636
rect 709 -1644 710 -1642
rect 716 -1638 717 -1636
rect 716 -1644 717 -1642
rect 723 -1638 724 -1636
rect 726 -1638 727 -1636
rect 726 -1644 727 -1642
rect 730 -1638 731 -1636
rect 733 -1638 734 -1636
rect 730 -1644 731 -1642
rect 733 -1644 734 -1642
rect 737 -1638 738 -1636
rect 737 -1644 738 -1642
rect 747 -1638 748 -1636
rect 744 -1644 745 -1642
rect 747 -1644 748 -1642
rect 751 -1638 752 -1636
rect 754 -1638 755 -1636
rect 751 -1644 752 -1642
rect 754 -1644 755 -1642
rect 758 -1638 759 -1636
rect 758 -1644 759 -1642
rect 765 -1638 766 -1636
rect 765 -1644 766 -1642
rect 772 -1638 773 -1636
rect 772 -1644 773 -1642
rect 779 -1638 780 -1636
rect 779 -1644 780 -1642
rect 786 -1638 787 -1636
rect 786 -1644 787 -1642
rect 793 -1638 794 -1636
rect 793 -1644 794 -1642
rect 800 -1638 801 -1636
rect 800 -1644 801 -1642
rect 807 -1638 808 -1636
rect 807 -1644 808 -1642
rect 814 -1638 815 -1636
rect 817 -1638 818 -1636
rect 814 -1644 815 -1642
rect 817 -1644 818 -1642
rect 821 -1638 822 -1636
rect 824 -1638 825 -1636
rect 824 -1644 825 -1642
rect 828 -1638 829 -1636
rect 828 -1644 829 -1642
rect 835 -1638 836 -1636
rect 835 -1644 836 -1642
rect 842 -1638 843 -1636
rect 842 -1644 843 -1642
rect 849 -1638 850 -1636
rect 849 -1644 850 -1642
rect 859 -1644 860 -1642
rect 863 -1638 864 -1636
rect 866 -1638 867 -1636
rect 863 -1644 864 -1642
rect 866 -1644 867 -1642
rect 870 -1638 871 -1636
rect 870 -1644 871 -1642
rect 877 -1638 878 -1636
rect 880 -1638 881 -1636
rect 877 -1644 878 -1642
rect 880 -1644 881 -1642
rect 884 -1638 885 -1636
rect 884 -1644 885 -1642
rect 891 -1638 892 -1636
rect 894 -1638 895 -1636
rect 891 -1644 892 -1642
rect 898 -1638 899 -1636
rect 898 -1644 899 -1642
rect 905 -1638 906 -1636
rect 905 -1644 906 -1642
rect 912 -1638 913 -1636
rect 912 -1644 913 -1642
rect 919 -1638 920 -1636
rect 919 -1644 920 -1642
rect 926 -1638 927 -1636
rect 926 -1644 927 -1642
rect 933 -1638 934 -1636
rect 933 -1644 934 -1642
rect 940 -1638 941 -1636
rect 940 -1644 941 -1642
rect 947 -1638 948 -1636
rect 947 -1644 948 -1642
rect 954 -1638 955 -1636
rect 957 -1638 958 -1636
rect 957 -1644 958 -1642
rect 961 -1638 962 -1636
rect 961 -1644 962 -1642
rect 968 -1638 969 -1636
rect 968 -1644 969 -1642
rect 975 -1638 976 -1636
rect 975 -1644 976 -1642
rect 982 -1638 983 -1636
rect 982 -1644 983 -1642
rect 989 -1638 990 -1636
rect 989 -1644 990 -1642
rect 996 -1638 997 -1636
rect 996 -1644 997 -1642
rect 1003 -1638 1004 -1636
rect 1006 -1638 1007 -1636
rect 1003 -1644 1004 -1642
rect 1006 -1644 1007 -1642
rect 1010 -1638 1011 -1636
rect 1010 -1644 1011 -1642
rect 1017 -1638 1018 -1636
rect 1020 -1638 1021 -1636
rect 1017 -1644 1018 -1642
rect 1020 -1644 1021 -1642
rect 1024 -1638 1025 -1636
rect 1024 -1644 1025 -1642
rect 1031 -1638 1032 -1636
rect 1031 -1644 1032 -1642
rect 1038 -1638 1039 -1636
rect 1038 -1644 1039 -1642
rect 1045 -1638 1046 -1636
rect 1045 -1644 1046 -1642
rect 1052 -1638 1053 -1636
rect 1052 -1644 1053 -1642
rect 1062 -1638 1063 -1636
rect 1059 -1644 1060 -1642
rect 1062 -1644 1063 -1642
rect 1066 -1638 1067 -1636
rect 1066 -1644 1067 -1642
rect 1073 -1638 1074 -1636
rect 1073 -1644 1074 -1642
rect 1080 -1638 1081 -1636
rect 1080 -1644 1081 -1642
rect 1083 -1644 1084 -1642
rect 1087 -1638 1088 -1636
rect 1087 -1644 1088 -1642
rect 1094 -1638 1095 -1636
rect 1094 -1644 1095 -1642
rect 1101 -1638 1102 -1636
rect 1101 -1644 1102 -1642
rect 1108 -1644 1109 -1642
rect 1111 -1644 1112 -1642
rect 1115 -1638 1116 -1636
rect 1115 -1644 1116 -1642
rect 1122 -1638 1123 -1636
rect 1125 -1638 1126 -1636
rect 1122 -1644 1123 -1642
rect 1125 -1644 1126 -1642
rect 1129 -1638 1130 -1636
rect 1129 -1644 1130 -1642
rect 1136 -1638 1137 -1636
rect 1136 -1644 1137 -1642
rect 1143 -1638 1144 -1636
rect 1143 -1644 1144 -1642
rect 1150 -1638 1151 -1636
rect 1150 -1644 1151 -1642
rect 1157 -1638 1158 -1636
rect 1157 -1644 1158 -1642
rect 1164 -1638 1165 -1636
rect 1164 -1644 1165 -1642
rect 1171 -1638 1172 -1636
rect 1171 -1644 1172 -1642
rect 1178 -1638 1179 -1636
rect 1178 -1644 1179 -1642
rect 1185 -1638 1186 -1636
rect 1188 -1638 1189 -1636
rect 1185 -1644 1186 -1642
rect 1192 -1638 1193 -1636
rect 1192 -1644 1193 -1642
rect 1199 -1638 1200 -1636
rect 1199 -1644 1200 -1642
rect 1206 -1638 1207 -1636
rect 1206 -1644 1207 -1642
rect 1209 -1644 1210 -1642
rect 1213 -1638 1214 -1636
rect 1213 -1644 1214 -1642
rect 1220 -1638 1221 -1636
rect 1220 -1644 1221 -1642
rect 1227 -1638 1228 -1636
rect 1227 -1644 1228 -1642
rect 1234 -1638 1235 -1636
rect 1234 -1644 1235 -1642
rect 1241 -1638 1242 -1636
rect 1241 -1644 1242 -1642
rect 1248 -1638 1249 -1636
rect 1248 -1644 1249 -1642
rect 1255 -1638 1256 -1636
rect 1255 -1644 1256 -1642
rect 1262 -1638 1263 -1636
rect 1262 -1644 1263 -1642
rect 1269 -1638 1270 -1636
rect 1269 -1644 1270 -1642
rect 1276 -1638 1277 -1636
rect 1276 -1644 1277 -1642
rect 1283 -1638 1284 -1636
rect 1283 -1644 1284 -1642
rect 1290 -1638 1291 -1636
rect 1290 -1644 1291 -1642
rect 1297 -1638 1298 -1636
rect 1300 -1644 1301 -1642
rect 1304 -1638 1305 -1636
rect 1304 -1644 1305 -1642
rect 1311 -1638 1312 -1636
rect 1311 -1644 1312 -1642
rect 1318 -1638 1319 -1636
rect 1318 -1644 1319 -1642
rect 1325 -1638 1326 -1636
rect 1325 -1644 1326 -1642
rect 1332 -1638 1333 -1636
rect 1332 -1644 1333 -1642
rect 1339 -1638 1340 -1636
rect 1339 -1644 1340 -1642
rect 1346 -1638 1347 -1636
rect 1346 -1644 1347 -1642
rect 1353 -1638 1354 -1636
rect 1353 -1644 1354 -1642
rect 1360 -1638 1361 -1636
rect 1360 -1644 1361 -1642
rect 1367 -1638 1368 -1636
rect 1367 -1644 1368 -1642
rect 1374 -1638 1375 -1636
rect 1374 -1644 1375 -1642
rect 1381 -1638 1382 -1636
rect 1381 -1644 1382 -1642
rect 1388 -1638 1389 -1636
rect 1388 -1644 1389 -1642
rect 1395 -1638 1396 -1636
rect 1395 -1644 1396 -1642
rect 1402 -1638 1403 -1636
rect 1402 -1644 1403 -1642
rect 1409 -1638 1410 -1636
rect 1409 -1644 1410 -1642
rect 1416 -1638 1417 -1636
rect 1416 -1644 1417 -1642
rect 1423 -1638 1424 -1636
rect 1423 -1644 1424 -1642
rect 1430 -1638 1431 -1636
rect 1430 -1644 1431 -1642
rect 1437 -1638 1438 -1636
rect 1437 -1644 1438 -1642
rect 1444 -1638 1445 -1636
rect 1444 -1644 1445 -1642
rect 1451 -1638 1452 -1636
rect 1454 -1638 1455 -1636
rect 1451 -1644 1452 -1642
rect 1458 -1638 1459 -1636
rect 1458 -1644 1459 -1642
rect 1465 -1638 1466 -1636
rect 1465 -1644 1466 -1642
rect 1472 -1638 1473 -1636
rect 1472 -1644 1473 -1642
rect 1479 -1638 1480 -1636
rect 1479 -1644 1480 -1642
rect 1486 -1638 1487 -1636
rect 1486 -1644 1487 -1642
rect 1493 -1638 1494 -1636
rect 1493 -1644 1494 -1642
rect 1500 -1638 1501 -1636
rect 1500 -1644 1501 -1642
rect 1507 -1638 1508 -1636
rect 1507 -1644 1508 -1642
rect 1514 -1638 1515 -1636
rect 1514 -1644 1515 -1642
rect 1521 -1638 1522 -1636
rect 1521 -1644 1522 -1642
rect 1528 -1638 1529 -1636
rect 1528 -1644 1529 -1642
rect 1535 -1638 1536 -1636
rect 1535 -1644 1536 -1642
rect 1542 -1638 1543 -1636
rect 1542 -1644 1543 -1642
rect 1549 -1638 1550 -1636
rect 1549 -1644 1550 -1642
rect 1556 -1638 1557 -1636
rect 1556 -1644 1557 -1642
rect 1563 -1638 1564 -1636
rect 1563 -1644 1564 -1642
rect 1570 -1638 1571 -1636
rect 1570 -1644 1571 -1642
rect 1577 -1638 1578 -1636
rect 1577 -1644 1578 -1642
rect 1584 -1638 1585 -1636
rect 1584 -1644 1585 -1642
rect 1591 -1638 1592 -1636
rect 1591 -1644 1592 -1642
rect 1598 -1638 1599 -1636
rect 1598 -1644 1599 -1642
rect 1605 -1638 1606 -1636
rect 1605 -1644 1606 -1642
rect 1612 -1638 1613 -1636
rect 1612 -1644 1613 -1642
rect 1619 -1638 1620 -1636
rect 1619 -1644 1620 -1642
rect 1626 -1638 1627 -1636
rect 1626 -1644 1627 -1642
rect 1633 -1638 1634 -1636
rect 1633 -1644 1634 -1642
rect 1640 -1638 1641 -1636
rect 1640 -1644 1641 -1642
rect 1647 -1638 1648 -1636
rect 1650 -1638 1651 -1636
rect 1647 -1644 1648 -1642
rect 1650 -1644 1651 -1642
rect 1654 -1638 1655 -1636
rect 1654 -1644 1655 -1642
rect 1661 -1638 1662 -1636
rect 1661 -1644 1662 -1642
rect 1668 -1638 1669 -1636
rect 1668 -1644 1669 -1642
rect 1675 -1638 1676 -1636
rect 1675 -1644 1676 -1642
rect 1682 -1638 1683 -1636
rect 1685 -1638 1686 -1636
rect 1682 -1644 1683 -1642
rect 1685 -1644 1686 -1642
rect 1689 -1638 1690 -1636
rect 1689 -1644 1690 -1642
rect 1696 -1638 1697 -1636
rect 1696 -1644 1697 -1642
rect 1706 -1638 1707 -1636
rect 1710 -1638 1711 -1636
rect 1710 -1644 1711 -1642
rect 1717 -1638 1718 -1636
rect 1717 -1644 1718 -1642
rect 1724 -1638 1725 -1636
rect 1724 -1644 1725 -1642
rect 1822 -1638 1823 -1636
rect 1822 -1644 1823 -1642
rect 23 -1785 24 -1783
rect 23 -1791 24 -1789
rect 30 -1785 31 -1783
rect 30 -1791 31 -1789
rect 37 -1785 38 -1783
rect 37 -1791 38 -1789
rect 44 -1785 45 -1783
rect 44 -1791 45 -1789
rect 51 -1785 52 -1783
rect 51 -1791 52 -1789
rect 58 -1785 59 -1783
rect 58 -1791 59 -1789
rect 65 -1785 66 -1783
rect 65 -1791 66 -1789
rect 72 -1785 73 -1783
rect 72 -1791 73 -1789
rect 75 -1791 76 -1789
rect 79 -1785 80 -1783
rect 79 -1791 80 -1789
rect 86 -1785 87 -1783
rect 89 -1785 90 -1783
rect 86 -1791 87 -1789
rect 89 -1791 90 -1789
rect 93 -1785 94 -1783
rect 93 -1791 94 -1789
rect 100 -1785 101 -1783
rect 100 -1791 101 -1789
rect 107 -1785 108 -1783
rect 107 -1791 108 -1789
rect 114 -1785 115 -1783
rect 117 -1791 118 -1789
rect 121 -1785 122 -1783
rect 121 -1791 122 -1789
rect 128 -1785 129 -1783
rect 128 -1791 129 -1789
rect 135 -1785 136 -1783
rect 135 -1791 136 -1789
rect 145 -1785 146 -1783
rect 145 -1791 146 -1789
rect 149 -1785 150 -1783
rect 149 -1791 150 -1789
rect 156 -1785 157 -1783
rect 159 -1785 160 -1783
rect 156 -1791 157 -1789
rect 159 -1791 160 -1789
rect 163 -1785 164 -1783
rect 163 -1791 164 -1789
rect 170 -1785 171 -1783
rect 170 -1791 171 -1789
rect 177 -1785 178 -1783
rect 177 -1791 178 -1789
rect 184 -1785 185 -1783
rect 184 -1791 185 -1789
rect 191 -1785 192 -1783
rect 191 -1791 192 -1789
rect 198 -1785 199 -1783
rect 198 -1791 199 -1789
rect 205 -1785 206 -1783
rect 205 -1791 206 -1789
rect 212 -1785 213 -1783
rect 219 -1785 220 -1783
rect 222 -1785 223 -1783
rect 219 -1791 220 -1789
rect 222 -1791 223 -1789
rect 226 -1785 227 -1783
rect 226 -1791 227 -1789
rect 236 -1785 237 -1783
rect 233 -1791 234 -1789
rect 236 -1791 237 -1789
rect 240 -1785 241 -1783
rect 240 -1791 241 -1789
rect 247 -1785 248 -1783
rect 247 -1791 248 -1789
rect 254 -1785 255 -1783
rect 254 -1791 255 -1789
rect 261 -1791 262 -1789
rect 264 -1791 265 -1789
rect 268 -1785 269 -1783
rect 268 -1791 269 -1789
rect 275 -1785 276 -1783
rect 275 -1791 276 -1789
rect 282 -1785 283 -1783
rect 282 -1791 283 -1789
rect 289 -1785 290 -1783
rect 289 -1791 290 -1789
rect 296 -1785 297 -1783
rect 296 -1791 297 -1789
rect 303 -1785 304 -1783
rect 303 -1791 304 -1789
rect 310 -1785 311 -1783
rect 310 -1791 311 -1789
rect 317 -1785 318 -1783
rect 317 -1791 318 -1789
rect 324 -1785 325 -1783
rect 324 -1791 325 -1789
rect 331 -1785 332 -1783
rect 331 -1791 332 -1789
rect 338 -1785 339 -1783
rect 338 -1791 339 -1789
rect 345 -1785 346 -1783
rect 345 -1791 346 -1789
rect 352 -1785 353 -1783
rect 352 -1791 353 -1789
rect 362 -1785 363 -1783
rect 359 -1791 360 -1789
rect 362 -1791 363 -1789
rect 366 -1785 367 -1783
rect 366 -1791 367 -1789
rect 373 -1785 374 -1783
rect 373 -1791 374 -1789
rect 383 -1785 384 -1783
rect 380 -1791 381 -1789
rect 383 -1791 384 -1789
rect 387 -1785 388 -1783
rect 387 -1791 388 -1789
rect 394 -1785 395 -1783
rect 394 -1791 395 -1789
rect 401 -1785 402 -1783
rect 401 -1791 402 -1789
rect 408 -1785 409 -1783
rect 408 -1791 409 -1789
rect 415 -1785 416 -1783
rect 415 -1791 416 -1789
rect 422 -1785 423 -1783
rect 422 -1791 423 -1789
rect 429 -1785 430 -1783
rect 429 -1791 430 -1789
rect 436 -1785 437 -1783
rect 436 -1791 437 -1789
rect 443 -1785 444 -1783
rect 443 -1791 444 -1789
rect 450 -1785 451 -1783
rect 450 -1791 451 -1789
rect 457 -1785 458 -1783
rect 457 -1791 458 -1789
rect 464 -1785 465 -1783
rect 464 -1791 465 -1789
rect 471 -1785 472 -1783
rect 471 -1791 472 -1789
rect 478 -1785 479 -1783
rect 478 -1791 479 -1789
rect 485 -1785 486 -1783
rect 485 -1791 486 -1789
rect 492 -1785 493 -1783
rect 492 -1791 493 -1789
rect 499 -1785 500 -1783
rect 502 -1785 503 -1783
rect 499 -1791 500 -1789
rect 502 -1791 503 -1789
rect 506 -1785 507 -1783
rect 506 -1791 507 -1789
rect 513 -1785 514 -1783
rect 513 -1791 514 -1789
rect 520 -1785 521 -1783
rect 520 -1791 521 -1789
rect 527 -1785 528 -1783
rect 527 -1791 528 -1789
rect 534 -1785 535 -1783
rect 537 -1785 538 -1783
rect 534 -1791 535 -1789
rect 537 -1791 538 -1789
rect 541 -1785 542 -1783
rect 544 -1785 545 -1783
rect 544 -1791 545 -1789
rect 548 -1785 549 -1783
rect 551 -1785 552 -1783
rect 548 -1791 549 -1789
rect 551 -1791 552 -1789
rect 555 -1785 556 -1783
rect 555 -1791 556 -1789
rect 562 -1785 563 -1783
rect 562 -1791 563 -1789
rect 569 -1785 570 -1783
rect 569 -1791 570 -1789
rect 576 -1785 577 -1783
rect 579 -1785 580 -1783
rect 579 -1791 580 -1789
rect 583 -1785 584 -1783
rect 583 -1791 584 -1789
rect 593 -1785 594 -1783
rect 590 -1791 591 -1789
rect 593 -1791 594 -1789
rect 597 -1785 598 -1783
rect 597 -1791 598 -1789
rect 604 -1785 605 -1783
rect 604 -1791 605 -1789
rect 611 -1785 612 -1783
rect 611 -1791 612 -1789
rect 618 -1785 619 -1783
rect 618 -1791 619 -1789
rect 625 -1785 626 -1783
rect 625 -1791 626 -1789
rect 635 -1785 636 -1783
rect 632 -1791 633 -1789
rect 635 -1791 636 -1789
rect 639 -1785 640 -1783
rect 639 -1791 640 -1789
rect 646 -1785 647 -1783
rect 646 -1791 647 -1789
rect 653 -1785 654 -1783
rect 653 -1791 654 -1789
rect 660 -1785 661 -1783
rect 660 -1791 661 -1789
rect 667 -1785 668 -1783
rect 667 -1791 668 -1789
rect 674 -1785 675 -1783
rect 677 -1785 678 -1783
rect 674 -1791 675 -1789
rect 677 -1791 678 -1789
rect 681 -1785 682 -1783
rect 681 -1791 682 -1789
rect 688 -1785 689 -1783
rect 688 -1791 689 -1789
rect 695 -1785 696 -1783
rect 695 -1791 696 -1789
rect 702 -1785 703 -1783
rect 705 -1785 706 -1783
rect 702 -1791 703 -1789
rect 709 -1785 710 -1783
rect 709 -1791 710 -1789
rect 716 -1785 717 -1783
rect 719 -1785 720 -1783
rect 716 -1791 717 -1789
rect 719 -1791 720 -1789
rect 723 -1785 724 -1783
rect 726 -1785 727 -1783
rect 726 -1791 727 -1789
rect 730 -1785 731 -1783
rect 733 -1791 734 -1789
rect 737 -1785 738 -1783
rect 737 -1791 738 -1789
rect 744 -1785 745 -1783
rect 744 -1791 745 -1789
rect 751 -1785 752 -1783
rect 751 -1791 752 -1789
rect 758 -1785 759 -1783
rect 758 -1791 759 -1789
rect 765 -1785 766 -1783
rect 765 -1791 766 -1789
rect 772 -1785 773 -1783
rect 772 -1791 773 -1789
rect 779 -1785 780 -1783
rect 782 -1785 783 -1783
rect 779 -1791 780 -1789
rect 782 -1791 783 -1789
rect 786 -1785 787 -1783
rect 789 -1785 790 -1783
rect 786 -1791 787 -1789
rect 789 -1791 790 -1789
rect 793 -1785 794 -1783
rect 793 -1791 794 -1789
rect 800 -1785 801 -1783
rect 800 -1791 801 -1789
rect 807 -1785 808 -1783
rect 807 -1791 808 -1789
rect 814 -1785 815 -1783
rect 814 -1791 815 -1789
rect 824 -1785 825 -1783
rect 821 -1791 822 -1789
rect 824 -1791 825 -1789
rect 828 -1785 829 -1783
rect 828 -1791 829 -1789
rect 835 -1785 836 -1783
rect 835 -1791 836 -1789
rect 842 -1785 843 -1783
rect 842 -1791 843 -1789
rect 849 -1785 850 -1783
rect 849 -1791 850 -1789
rect 856 -1785 857 -1783
rect 856 -1791 857 -1789
rect 863 -1785 864 -1783
rect 863 -1791 864 -1789
rect 870 -1785 871 -1783
rect 870 -1791 871 -1789
rect 877 -1785 878 -1783
rect 877 -1791 878 -1789
rect 884 -1785 885 -1783
rect 887 -1785 888 -1783
rect 884 -1791 885 -1789
rect 887 -1791 888 -1789
rect 891 -1785 892 -1783
rect 891 -1791 892 -1789
rect 898 -1785 899 -1783
rect 901 -1785 902 -1783
rect 898 -1791 899 -1789
rect 901 -1791 902 -1789
rect 905 -1785 906 -1783
rect 905 -1791 906 -1789
rect 912 -1785 913 -1783
rect 912 -1791 913 -1789
rect 919 -1785 920 -1783
rect 919 -1791 920 -1789
rect 926 -1785 927 -1783
rect 926 -1791 927 -1789
rect 933 -1785 934 -1783
rect 933 -1791 934 -1789
rect 940 -1785 941 -1783
rect 940 -1791 941 -1789
rect 947 -1785 948 -1783
rect 950 -1785 951 -1783
rect 947 -1791 948 -1789
rect 954 -1785 955 -1783
rect 954 -1791 955 -1789
rect 961 -1785 962 -1783
rect 961 -1791 962 -1789
rect 968 -1785 969 -1783
rect 968 -1791 969 -1789
rect 978 -1785 979 -1783
rect 975 -1791 976 -1789
rect 978 -1791 979 -1789
rect 982 -1785 983 -1783
rect 982 -1791 983 -1789
rect 989 -1785 990 -1783
rect 989 -1791 990 -1789
rect 996 -1785 997 -1783
rect 996 -1791 997 -1789
rect 1003 -1785 1004 -1783
rect 1003 -1791 1004 -1789
rect 1010 -1785 1011 -1783
rect 1010 -1791 1011 -1789
rect 1017 -1785 1018 -1783
rect 1017 -1791 1018 -1789
rect 1024 -1785 1025 -1783
rect 1027 -1785 1028 -1783
rect 1024 -1791 1025 -1789
rect 1027 -1791 1028 -1789
rect 1031 -1785 1032 -1783
rect 1031 -1791 1032 -1789
rect 1038 -1785 1039 -1783
rect 1038 -1791 1039 -1789
rect 1045 -1785 1046 -1783
rect 1045 -1791 1046 -1789
rect 1052 -1785 1053 -1783
rect 1055 -1785 1056 -1783
rect 1052 -1791 1053 -1789
rect 1059 -1785 1060 -1783
rect 1059 -1791 1060 -1789
rect 1066 -1785 1067 -1783
rect 1066 -1791 1067 -1789
rect 1073 -1785 1074 -1783
rect 1073 -1791 1074 -1789
rect 1080 -1785 1081 -1783
rect 1080 -1791 1081 -1789
rect 1087 -1785 1088 -1783
rect 1087 -1791 1088 -1789
rect 1094 -1785 1095 -1783
rect 1094 -1791 1095 -1789
rect 1101 -1785 1102 -1783
rect 1101 -1791 1102 -1789
rect 1108 -1785 1109 -1783
rect 1108 -1791 1109 -1789
rect 1115 -1785 1116 -1783
rect 1115 -1791 1116 -1789
rect 1122 -1785 1123 -1783
rect 1122 -1791 1123 -1789
rect 1129 -1785 1130 -1783
rect 1129 -1791 1130 -1789
rect 1136 -1785 1137 -1783
rect 1136 -1791 1137 -1789
rect 1143 -1785 1144 -1783
rect 1146 -1785 1147 -1783
rect 1146 -1791 1147 -1789
rect 1150 -1785 1151 -1783
rect 1150 -1791 1151 -1789
rect 1157 -1785 1158 -1783
rect 1157 -1791 1158 -1789
rect 1164 -1785 1165 -1783
rect 1164 -1791 1165 -1789
rect 1171 -1785 1172 -1783
rect 1171 -1791 1172 -1789
rect 1178 -1785 1179 -1783
rect 1178 -1791 1179 -1789
rect 1185 -1785 1186 -1783
rect 1185 -1791 1186 -1789
rect 1192 -1785 1193 -1783
rect 1192 -1791 1193 -1789
rect 1199 -1785 1200 -1783
rect 1199 -1791 1200 -1789
rect 1206 -1785 1207 -1783
rect 1206 -1791 1207 -1789
rect 1213 -1785 1214 -1783
rect 1213 -1791 1214 -1789
rect 1220 -1785 1221 -1783
rect 1220 -1791 1221 -1789
rect 1227 -1785 1228 -1783
rect 1227 -1791 1228 -1789
rect 1234 -1785 1235 -1783
rect 1234 -1791 1235 -1789
rect 1241 -1785 1242 -1783
rect 1241 -1791 1242 -1789
rect 1248 -1785 1249 -1783
rect 1248 -1791 1249 -1789
rect 1255 -1785 1256 -1783
rect 1255 -1791 1256 -1789
rect 1262 -1785 1263 -1783
rect 1262 -1791 1263 -1789
rect 1269 -1785 1270 -1783
rect 1269 -1791 1270 -1789
rect 1276 -1785 1277 -1783
rect 1276 -1791 1277 -1789
rect 1283 -1785 1284 -1783
rect 1283 -1791 1284 -1789
rect 1290 -1791 1291 -1789
rect 1293 -1791 1294 -1789
rect 1297 -1785 1298 -1783
rect 1297 -1791 1298 -1789
rect 1304 -1785 1305 -1783
rect 1304 -1791 1305 -1789
rect 1311 -1785 1312 -1783
rect 1311 -1791 1312 -1789
rect 1318 -1785 1319 -1783
rect 1318 -1791 1319 -1789
rect 1325 -1785 1326 -1783
rect 1325 -1791 1326 -1789
rect 1332 -1785 1333 -1783
rect 1332 -1791 1333 -1789
rect 1339 -1785 1340 -1783
rect 1339 -1791 1340 -1789
rect 1346 -1785 1347 -1783
rect 1346 -1791 1347 -1789
rect 1353 -1785 1354 -1783
rect 1353 -1791 1354 -1789
rect 1360 -1785 1361 -1783
rect 1360 -1791 1361 -1789
rect 1367 -1785 1368 -1783
rect 1367 -1791 1368 -1789
rect 1374 -1785 1375 -1783
rect 1374 -1791 1375 -1789
rect 1381 -1785 1382 -1783
rect 1381 -1791 1382 -1789
rect 1388 -1785 1389 -1783
rect 1388 -1791 1389 -1789
rect 1395 -1785 1396 -1783
rect 1395 -1791 1396 -1789
rect 1402 -1785 1403 -1783
rect 1402 -1791 1403 -1789
rect 1409 -1785 1410 -1783
rect 1409 -1791 1410 -1789
rect 1416 -1785 1417 -1783
rect 1416 -1791 1417 -1789
rect 1423 -1785 1424 -1783
rect 1423 -1791 1424 -1789
rect 1426 -1791 1427 -1789
rect 1430 -1785 1431 -1783
rect 1430 -1791 1431 -1789
rect 1437 -1785 1438 -1783
rect 1437 -1791 1438 -1789
rect 1444 -1785 1445 -1783
rect 1444 -1791 1445 -1789
rect 1451 -1785 1452 -1783
rect 1451 -1791 1452 -1789
rect 1458 -1785 1459 -1783
rect 1458 -1791 1459 -1789
rect 1465 -1785 1466 -1783
rect 1465 -1791 1466 -1789
rect 1472 -1785 1473 -1783
rect 1472 -1791 1473 -1789
rect 1479 -1785 1480 -1783
rect 1479 -1791 1480 -1789
rect 1486 -1785 1487 -1783
rect 1486 -1791 1487 -1789
rect 1493 -1785 1494 -1783
rect 1493 -1791 1494 -1789
rect 1500 -1785 1501 -1783
rect 1500 -1791 1501 -1789
rect 1507 -1785 1508 -1783
rect 1507 -1791 1508 -1789
rect 1514 -1785 1515 -1783
rect 1514 -1791 1515 -1789
rect 1521 -1785 1522 -1783
rect 1521 -1791 1522 -1789
rect 1528 -1785 1529 -1783
rect 1528 -1791 1529 -1789
rect 1535 -1785 1536 -1783
rect 1535 -1791 1536 -1789
rect 1542 -1785 1543 -1783
rect 1542 -1791 1543 -1789
rect 1549 -1785 1550 -1783
rect 1549 -1791 1550 -1789
rect 1556 -1785 1557 -1783
rect 1556 -1791 1557 -1789
rect 1563 -1785 1564 -1783
rect 1563 -1791 1564 -1789
rect 1570 -1785 1571 -1783
rect 1570 -1791 1571 -1789
rect 1577 -1785 1578 -1783
rect 1577 -1791 1578 -1789
rect 1584 -1785 1585 -1783
rect 1584 -1791 1585 -1789
rect 1591 -1785 1592 -1783
rect 1591 -1791 1592 -1789
rect 1598 -1785 1599 -1783
rect 1598 -1791 1599 -1789
rect 1605 -1785 1606 -1783
rect 1605 -1791 1606 -1789
rect 1612 -1785 1613 -1783
rect 1612 -1791 1613 -1789
rect 1619 -1785 1620 -1783
rect 1619 -1791 1620 -1789
rect 1626 -1785 1627 -1783
rect 1626 -1791 1627 -1789
rect 1633 -1785 1634 -1783
rect 1633 -1791 1634 -1789
rect 1640 -1785 1641 -1783
rect 1640 -1791 1641 -1789
rect 1647 -1785 1648 -1783
rect 1647 -1791 1648 -1789
rect 1654 -1785 1655 -1783
rect 1654 -1791 1655 -1789
rect 1661 -1785 1662 -1783
rect 1661 -1791 1662 -1789
rect 1668 -1785 1669 -1783
rect 1668 -1791 1669 -1789
rect 1675 -1785 1676 -1783
rect 1675 -1791 1676 -1789
rect 1682 -1785 1683 -1783
rect 1682 -1791 1683 -1789
rect 1689 -1785 1690 -1783
rect 1689 -1791 1690 -1789
rect 1696 -1785 1697 -1783
rect 1696 -1791 1697 -1789
rect 1703 -1785 1704 -1783
rect 1703 -1791 1704 -1789
rect 1710 -1785 1711 -1783
rect 1710 -1791 1711 -1789
rect 1717 -1785 1718 -1783
rect 1717 -1791 1718 -1789
rect 1724 -1785 1725 -1783
rect 1724 -1791 1725 -1789
rect 1731 -1785 1732 -1783
rect 1731 -1791 1732 -1789
rect 1738 -1785 1739 -1783
rect 1738 -1791 1739 -1789
rect 1745 -1785 1746 -1783
rect 1745 -1791 1746 -1789
rect 1752 -1785 1753 -1783
rect 1752 -1791 1753 -1789
rect 1759 -1785 1760 -1783
rect 1759 -1791 1760 -1789
rect 1766 -1785 1767 -1783
rect 1766 -1791 1767 -1789
rect 1773 -1785 1774 -1783
rect 1773 -1791 1774 -1789
rect 1780 -1785 1781 -1783
rect 1780 -1791 1781 -1789
rect 1787 -1785 1788 -1783
rect 1787 -1791 1788 -1789
rect 1794 -1785 1795 -1783
rect 1794 -1791 1795 -1789
rect 1801 -1785 1802 -1783
rect 1801 -1791 1802 -1789
rect 1808 -1785 1809 -1783
rect 1808 -1791 1809 -1789
rect 1815 -1785 1816 -1783
rect 1815 -1791 1816 -1789
rect 1822 -1785 1823 -1783
rect 1822 -1791 1823 -1789
rect 1829 -1785 1830 -1783
rect 1829 -1791 1830 -1789
rect 1836 -1785 1837 -1783
rect 1839 -1785 1840 -1783
rect 1836 -1791 1837 -1789
rect 1839 -1791 1840 -1789
rect 30 -1924 31 -1922
rect 30 -1930 31 -1928
rect 37 -1924 38 -1922
rect 37 -1930 38 -1928
rect 44 -1924 45 -1922
rect 44 -1930 45 -1928
rect 51 -1924 52 -1922
rect 51 -1930 52 -1928
rect 58 -1924 59 -1922
rect 61 -1924 62 -1922
rect 61 -1930 62 -1928
rect 68 -1924 69 -1922
rect 65 -1930 66 -1928
rect 68 -1930 69 -1928
rect 72 -1924 73 -1922
rect 72 -1930 73 -1928
rect 79 -1924 80 -1922
rect 79 -1930 80 -1928
rect 86 -1924 87 -1922
rect 86 -1930 87 -1928
rect 93 -1924 94 -1922
rect 93 -1930 94 -1928
rect 100 -1924 101 -1922
rect 100 -1930 101 -1928
rect 107 -1924 108 -1922
rect 110 -1924 111 -1922
rect 107 -1930 108 -1928
rect 114 -1924 115 -1922
rect 114 -1930 115 -1928
rect 121 -1924 122 -1922
rect 121 -1930 122 -1928
rect 128 -1924 129 -1922
rect 128 -1930 129 -1928
rect 135 -1924 136 -1922
rect 135 -1930 136 -1928
rect 142 -1924 143 -1922
rect 142 -1930 143 -1928
rect 149 -1924 150 -1922
rect 149 -1930 150 -1928
rect 156 -1924 157 -1922
rect 156 -1930 157 -1928
rect 163 -1924 164 -1922
rect 163 -1930 164 -1928
rect 173 -1924 174 -1922
rect 170 -1930 171 -1928
rect 173 -1930 174 -1928
rect 177 -1924 178 -1922
rect 177 -1930 178 -1928
rect 184 -1924 185 -1922
rect 184 -1930 185 -1928
rect 191 -1924 192 -1922
rect 191 -1930 192 -1928
rect 198 -1924 199 -1922
rect 198 -1930 199 -1928
rect 205 -1924 206 -1922
rect 205 -1930 206 -1928
rect 212 -1930 213 -1928
rect 219 -1924 220 -1922
rect 222 -1924 223 -1922
rect 219 -1930 220 -1928
rect 226 -1924 227 -1922
rect 226 -1930 227 -1928
rect 229 -1930 230 -1928
rect 233 -1924 234 -1922
rect 233 -1930 234 -1928
rect 243 -1924 244 -1922
rect 240 -1930 241 -1928
rect 243 -1930 244 -1928
rect 250 -1924 251 -1922
rect 247 -1930 248 -1928
rect 250 -1930 251 -1928
rect 254 -1924 255 -1922
rect 254 -1930 255 -1928
rect 261 -1924 262 -1922
rect 261 -1930 262 -1928
rect 268 -1924 269 -1922
rect 268 -1930 269 -1928
rect 275 -1924 276 -1922
rect 275 -1930 276 -1928
rect 282 -1924 283 -1922
rect 282 -1930 283 -1928
rect 289 -1924 290 -1922
rect 289 -1930 290 -1928
rect 296 -1924 297 -1922
rect 296 -1930 297 -1928
rect 303 -1924 304 -1922
rect 303 -1930 304 -1928
rect 310 -1924 311 -1922
rect 310 -1930 311 -1928
rect 317 -1924 318 -1922
rect 317 -1930 318 -1928
rect 324 -1924 325 -1922
rect 324 -1930 325 -1928
rect 331 -1924 332 -1922
rect 331 -1930 332 -1928
rect 338 -1924 339 -1922
rect 341 -1924 342 -1922
rect 338 -1930 339 -1928
rect 345 -1924 346 -1922
rect 345 -1930 346 -1928
rect 352 -1924 353 -1922
rect 352 -1930 353 -1928
rect 359 -1924 360 -1922
rect 359 -1930 360 -1928
rect 366 -1924 367 -1922
rect 366 -1930 367 -1928
rect 373 -1924 374 -1922
rect 373 -1930 374 -1928
rect 380 -1924 381 -1922
rect 380 -1930 381 -1928
rect 387 -1924 388 -1922
rect 387 -1930 388 -1928
rect 394 -1924 395 -1922
rect 394 -1930 395 -1928
rect 401 -1924 402 -1922
rect 404 -1924 405 -1922
rect 401 -1930 402 -1928
rect 404 -1930 405 -1928
rect 408 -1924 409 -1922
rect 408 -1930 409 -1928
rect 415 -1924 416 -1922
rect 415 -1930 416 -1928
rect 422 -1924 423 -1922
rect 422 -1930 423 -1928
rect 432 -1924 433 -1922
rect 429 -1930 430 -1928
rect 432 -1930 433 -1928
rect 436 -1924 437 -1922
rect 436 -1930 437 -1928
rect 443 -1924 444 -1922
rect 443 -1930 444 -1928
rect 450 -1924 451 -1922
rect 450 -1930 451 -1928
rect 457 -1924 458 -1922
rect 457 -1930 458 -1928
rect 464 -1924 465 -1922
rect 464 -1930 465 -1928
rect 471 -1924 472 -1922
rect 471 -1930 472 -1928
rect 478 -1924 479 -1922
rect 478 -1930 479 -1928
rect 485 -1924 486 -1922
rect 485 -1930 486 -1928
rect 492 -1924 493 -1922
rect 492 -1930 493 -1928
rect 499 -1924 500 -1922
rect 499 -1930 500 -1928
rect 506 -1924 507 -1922
rect 506 -1930 507 -1928
rect 513 -1924 514 -1922
rect 513 -1930 514 -1928
rect 520 -1924 521 -1922
rect 520 -1930 521 -1928
rect 527 -1924 528 -1922
rect 527 -1930 528 -1928
rect 530 -1930 531 -1928
rect 534 -1924 535 -1922
rect 534 -1930 535 -1928
rect 541 -1924 542 -1922
rect 541 -1930 542 -1928
rect 548 -1924 549 -1922
rect 548 -1930 549 -1928
rect 555 -1924 556 -1922
rect 555 -1930 556 -1928
rect 562 -1924 563 -1922
rect 562 -1930 563 -1928
rect 569 -1924 570 -1922
rect 569 -1930 570 -1928
rect 576 -1924 577 -1922
rect 576 -1930 577 -1928
rect 583 -1924 584 -1922
rect 583 -1930 584 -1928
rect 590 -1924 591 -1922
rect 593 -1924 594 -1922
rect 590 -1930 591 -1928
rect 593 -1930 594 -1928
rect 597 -1924 598 -1922
rect 597 -1930 598 -1928
rect 604 -1924 605 -1922
rect 604 -1930 605 -1928
rect 611 -1924 612 -1922
rect 611 -1930 612 -1928
rect 618 -1924 619 -1922
rect 621 -1924 622 -1922
rect 618 -1930 619 -1928
rect 621 -1930 622 -1928
rect 625 -1924 626 -1922
rect 625 -1930 626 -1928
rect 632 -1924 633 -1922
rect 632 -1930 633 -1928
rect 639 -1924 640 -1922
rect 639 -1930 640 -1928
rect 646 -1924 647 -1922
rect 646 -1930 647 -1928
rect 653 -1924 654 -1922
rect 656 -1924 657 -1922
rect 653 -1930 654 -1928
rect 656 -1930 657 -1928
rect 660 -1924 661 -1922
rect 660 -1930 661 -1928
rect 670 -1924 671 -1922
rect 667 -1930 668 -1928
rect 670 -1930 671 -1928
rect 674 -1924 675 -1922
rect 674 -1930 675 -1928
rect 681 -1924 682 -1922
rect 684 -1924 685 -1922
rect 681 -1930 682 -1928
rect 684 -1930 685 -1928
rect 688 -1924 689 -1922
rect 688 -1930 689 -1928
rect 695 -1924 696 -1922
rect 695 -1930 696 -1928
rect 702 -1924 703 -1922
rect 702 -1930 703 -1928
rect 709 -1924 710 -1922
rect 709 -1930 710 -1928
rect 716 -1924 717 -1922
rect 716 -1930 717 -1928
rect 723 -1924 724 -1922
rect 726 -1924 727 -1922
rect 726 -1930 727 -1928
rect 730 -1924 731 -1922
rect 730 -1930 731 -1928
rect 737 -1924 738 -1922
rect 737 -1930 738 -1928
rect 744 -1924 745 -1922
rect 744 -1930 745 -1928
rect 751 -1924 752 -1922
rect 751 -1930 752 -1928
rect 758 -1924 759 -1922
rect 758 -1930 759 -1928
rect 765 -1924 766 -1922
rect 765 -1930 766 -1928
rect 772 -1924 773 -1922
rect 772 -1930 773 -1928
rect 779 -1924 780 -1922
rect 779 -1930 780 -1928
rect 786 -1924 787 -1922
rect 789 -1924 790 -1922
rect 786 -1930 787 -1928
rect 789 -1930 790 -1928
rect 793 -1924 794 -1922
rect 793 -1930 794 -1928
rect 800 -1924 801 -1922
rect 800 -1930 801 -1928
rect 807 -1924 808 -1922
rect 810 -1924 811 -1922
rect 807 -1930 808 -1928
rect 810 -1930 811 -1928
rect 814 -1924 815 -1922
rect 814 -1930 815 -1928
rect 821 -1924 822 -1922
rect 821 -1930 822 -1928
rect 828 -1924 829 -1922
rect 831 -1924 832 -1922
rect 828 -1930 829 -1928
rect 835 -1924 836 -1922
rect 835 -1930 836 -1928
rect 842 -1924 843 -1922
rect 842 -1930 843 -1928
rect 849 -1924 850 -1922
rect 856 -1924 857 -1922
rect 856 -1930 857 -1928
rect 863 -1924 864 -1922
rect 863 -1930 864 -1928
rect 870 -1924 871 -1922
rect 870 -1930 871 -1928
rect 873 -1930 874 -1928
rect 877 -1924 878 -1922
rect 877 -1930 878 -1928
rect 884 -1924 885 -1922
rect 884 -1930 885 -1928
rect 891 -1924 892 -1922
rect 891 -1930 892 -1928
rect 898 -1924 899 -1922
rect 898 -1930 899 -1928
rect 905 -1924 906 -1922
rect 905 -1930 906 -1928
rect 912 -1924 913 -1922
rect 915 -1924 916 -1922
rect 912 -1930 913 -1928
rect 915 -1930 916 -1928
rect 919 -1924 920 -1922
rect 919 -1930 920 -1928
rect 926 -1924 927 -1922
rect 926 -1930 927 -1928
rect 933 -1924 934 -1922
rect 933 -1930 934 -1928
rect 940 -1924 941 -1922
rect 940 -1930 941 -1928
rect 947 -1924 948 -1922
rect 947 -1930 948 -1928
rect 954 -1924 955 -1922
rect 954 -1930 955 -1928
rect 961 -1924 962 -1922
rect 961 -1930 962 -1928
rect 968 -1924 969 -1922
rect 968 -1930 969 -1928
rect 975 -1924 976 -1922
rect 975 -1930 976 -1928
rect 985 -1924 986 -1922
rect 982 -1930 983 -1928
rect 985 -1930 986 -1928
rect 989 -1924 990 -1922
rect 992 -1924 993 -1922
rect 989 -1930 990 -1928
rect 996 -1924 997 -1922
rect 996 -1930 997 -1928
rect 1003 -1924 1004 -1922
rect 1003 -1930 1004 -1928
rect 1010 -1924 1011 -1922
rect 1010 -1930 1011 -1928
rect 1017 -1924 1018 -1922
rect 1017 -1930 1018 -1928
rect 1024 -1924 1025 -1922
rect 1024 -1930 1025 -1928
rect 1031 -1924 1032 -1922
rect 1031 -1930 1032 -1928
rect 1038 -1924 1039 -1922
rect 1038 -1930 1039 -1928
rect 1045 -1924 1046 -1922
rect 1045 -1930 1046 -1928
rect 1052 -1924 1053 -1922
rect 1052 -1930 1053 -1928
rect 1059 -1924 1060 -1922
rect 1059 -1930 1060 -1928
rect 1066 -1924 1067 -1922
rect 1066 -1930 1067 -1928
rect 1073 -1924 1074 -1922
rect 1073 -1930 1074 -1928
rect 1080 -1924 1081 -1922
rect 1080 -1930 1081 -1928
rect 1087 -1924 1088 -1922
rect 1087 -1930 1088 -1928
rect 1094 -1924 1095 -1922
rect 1097 -1924 1098 -1922
rect 1094 -1930 1095 -1928
rect 1097 -1930 1098 -1928
rect 1101 -1924 1102 -1922
rect 1101 -1930 1102 -1928
rect 1108 -1924 1109 -1922
rect 1108 -1930 1109 -1928
rect 1115 -1924 1116 -1922
rect 1115 -1930 1116 -1928
rect 1125 -1924 1126 -1922
rect 1122 -1930 1123 -1928
rect 1125 -1930 1126 -1928
rect 1129 -1924 1130 -1922
rect 1129 -1930 1130 -1928
rect 1136 -1924 1137 -1922
rect 1136 -1930 1137 -1928
rect 1143 -1924 1144 -1922
rect 1143 -1930 1144 -1928
rect 1150 -1924 1151 -1922
rect 1150 -1930 1151 -1928
rect 1157 -1924 1158 -1922
rect 1160 -1924 1161 -1922
rect 1157 -1930 1158 -1928
rect 1160 -1930 1161 -1928
rect 1164 -1924 1165 -1922
rect 1167 -1924 1168 -1922
rect 1164 -1930 1165 -1928
rect 1167 -1930 1168 -1928
rect 1171 -1924 1172 -1922
rect 1171 -1930 1172 -1928
rect 1178 -1924 1179 -1922
rect 1178 -1930 1179 -1928
rect 1185 -1924 1186 -1922
rect 1185 -1930 1186 -1928
rect 1192 -1924 1193 -1922
rect 1192 -1930 1193 -1928
rect 1199 -1924 1200 -1922
rect 1199 -1930 1200 -1928
rect 1206 -1924 1207 -1922
rect 1206 -1930 1207 -1928
rect 1213 -1924 1214 -1922
rect 1213 -1930 1214 -1928
rect 1220 -1924 1221 -1922
rect 1220 -1930 1221 -1928
rect 1227 -1924 1228 -1922
rect 1230 -1924 1231 -1922
rect 1227 -1930 1228 -1928
rect 1230 -1930 1231 -1928
rect 1234 -1924 1235 -1922
rect 1234 -1930 1235 -1928
rect 1241 -1924 1242 -1922
rect 1241 -1930 1242 -1928
rect 1248 -1924 1249 -1922
rect 1248 -1930 1249 -1928
rect 1255 -1924 1256 -1922
rect 1255 -1930 1256 -1928
rect 1262 -1924 1263 -1922
rect 1262 -1930 1263 -1928
rect 1269 -1924 1270 -1922
rect 1269 -1930 1270 -1928
rect 1276 -1924 1277 -1922
rect 1276 -1930 1277 -1928
rect 1283 -1924 1284 -1922
rect 1283 -1930 1284 -1928
rect 1290 -1924 1291 -1922
rect 1290 -1930 1291 -1928
rect 1297 -1924 1298 -1922
rect 1297 -1930 1298 -1928
rect 1304 -1924 1305 -1922
rect 1304 -1930 1305 -1928
rect 1311 -1924 1312 -1922
rect 1311 -1930 1312 -1928
rect 1318 -1924 1319 -1922
rect 1318 -1930 1319 -1928
rect 1325 -1924 1326 -1922
rect 1325 -1930 1326 -1928
rect 1332 -1924 1333 -1922
rect 1332 -1930 1333 -1928
rect 1339 -1924 1340 -1922
rect 1339 -1930 1340 -1928
rect 1346 -1924 1347 -1922
rect 1346 -1930 1347 -1928
rect 1353 -1924 1354 -1922
rect 1353 -1930 1354 -1928
rect 1360 -1924 1361 -1922
rect 1360 -1930 1361 -1928
rect 1367 -1924 1368 -1922
rect 1367 -1930 1368 -1928
rect 1374 -1924 1375 -1922
rect 1374 -1930 1375 -1928
rect 1381 -1924 1382 -1922
rect 1384 -1924 1385 -1922
rect 1381 -1930 1382 -1928
rect 1384 -1930 1385 -1928
rect 1388 -1924 1389 -1922
rect 1388 -1930 1389 -1928
rect 1395 -1924 1396 -1922
rect 1395 -1930 1396 -1928
rect 1402 -1924 1403 -1922
rect 1402 -1930 1403 -1928
rect 1409 -1924 1410 -1922
rect 1409 -1930 1410 -1928
rect 1416 -1924 1417 -1922
rect 1416 -1930 1417 -1928
rect 1423 -1924 1424 -1922
rect 1426 -1924 1427 -1922
rect 1423 -1930 1424 -1928
rect 1430 -1924 1431 -1922
rect 1430 -1930 1431 -1928
rect 1437 -1924 1438 -1922
rect 1437 -1930 1438 -1928
rect 1444 -1924 1445 -1922
rect 1444 -1930 1445 -1928
rect 1451 -1924 1452 -1922
rect 1451 -1930 1452 -1928
rect 1458 -1924 1459 -1922
rect 1458 -1930 1459 -1928
rect 1465 -1924 1466 -1922
rect 1465 -1930 1466 -1928
rect 1472 -1924 1473 -1922
rect 1472 -1930 1473 -1928
rect 1479 -1924 1480 -1922
rect 1479 -1930 1480 -1928
rect 1486 -1924 1487 -1922
rect 1486 -1930 1487 -1928
rect 1493 -1924 1494 -1922
rect 1493 -1930 1494 -1928
rect 1500 -1924 1501 -1922
rect 1500 -1930 1501 -1928
rect 1507 -1924 1508 -1922
rect 1507 -1930 1508 -1928
rect 1514 -1924 1515 -1922
rect 1514 -1930 1515 -1928
rect 1521 -1924 1522 -1922
rect 1521 -1930 1522 -1928
rect 1528 -1924 1529 -1922
rect 1528 -1930 1529 -1928
rect 1535 -1924 1536 -1922
rect 1535 -1930 1536 -1928
rect 1542 -1924 1543 -1922
rect 1542 -1930 1543 -1928
rect 1549 -1924 1550 -1922
rect 1549 -1930 1550 -1928
rect 1556 -1924 1557 -1922
rect 1556 -1930 1557 -1928
rect 1563 -1924 1564 -1922
rect 1563 -1930 1564 -1928
rect 1570 -1924 1571 -1922
rect 1570 -1930 1571 -1928
rect 1577 -1924 1578 -1922
rect 1577 -1930 1578 -1928
rect 1584 -1924 1585 -1922
rect 1584 -1930 1585 -1928
rect 1591 -1924 1592 -1922
rect 1591 -1930 1592 -1928
rect 1598 -1924 1599 -1922
rect 1598 -1930 1599 -1928
rect 1605 -1924 1606 -1922
rect 1605 -1930 1606 -1928
rect 1612 -1924 1613 -1922
rect 1612 -1930 1613 -1928
rect 1619 -1924 1620 -1922
rect 1619 -1930 1620 -1928
rect 1626 -1924 1627 -1922
rect 1626 -1930 1627 -1928
rect 1633 -1924 1634 -1922
rect 1633 -1930 1634 -1928
rect 1640 -1924 1641 -1922
rect 1640 -1930 1641 -1928
rect 1647 -1924 1648 -1922
rect 1647 -1930 1648 -1928
rect 1654 -1924 1655 -1922
rect 1654 -1930 1655 -1928
rect 1661 -1924 1662 -1922
rect 1661 -1930 1662 -1928
rect 1668 -1924 1669 -1922
rect 1668 -1930 1669 -1928
rect 1675 -1924 1676 -1922
rect 1675 -1930 1676 -1928
rect 1682 -1924 1683 -1922
rect 1682 -1930 1683 -1928
rect 1689 -1924 1690 -1922
rect 1689 -1930 1690 -1928
rect 1696 -1924 1697 -1922
rect 1696 -1930 1697 -1928
rect 1703 -1924 1704 -1922
rect 1703 -1930 1704 -1928
rect 1710 -1924 1711 -1922
rect 1710 -1930 1711 -1928
rect 1717 -1924 1718 -1922
rect 1717 -1930 1718 -1928
rect 1724 -1924 1725 -1922
rect 1724 -1930 1725 -1928
rect 1731 -1924 1732 -1922
rect 1731 -1930 1732 -1928
rect 1738 -1924 1739 -1922
rect 1738 -1930 1739 -1928
rect 1745 -1924 1746 -1922
rect 1745 -1930 1746 -1928
rect 1755 -1924 1756 -1922
rect 1759 -1924 1760 -1922
rect 1759 -1930 1760 -1928
rect 1766 -1924 1767 -1922
rect 1766 -1930 1767 -1928
rect 1794 -1924 1795 -1922
rect 1794 -1930 1795 -1928
rect 23 -2051 24 -2049
rect 23 -2057 24 -2055
rect 37 -2051 38 -2049
rect 37 -2057 38 -2055
rect 44 -2051 45 -2049
rect 44 -2057 45 -2055
rect 51 -2051 52 -2049
rect 51 -2057 52 -2055
rect 58 -2051 59 -2049
rect 58 -2057 59 -2055
rect 65 -2051 66 -2049
rect 65 -2057 66 -2055
rect 72 -2051 73 -2049
rect 72 -2057 73 -2055
rect 79 -2051 80 -2049
rect 79 -2057 80 -2055
rect 86 -2051 87 -2049
rect 86 -2057 87 -2055
rect 93 -2051 94 -2049
rect 93 -2057 94 -2055
rect 100 -2051 101 -2049
rect 100 -2057 101 -2055
rect 107 -2051 108 -2049
rect 110 -2051 111 -2049
rect 107 -2057 108 -2055
rect 114 -2051 115 -2049
rect 117 -2051 118 -2049
rect 114 -2057 115 -2055
rect 121 -2051 122 -2049
rect 121 -2057 122 -2055
rect 128 -2051 129 -2049
rect 131 -2051 132 -2049
rect 128 -2057 129 -2055
rect 135 -2051 136 -2049
rect 138 -2051 139 -2049
rect 142 -2051 143 -2049
rect 142 -2057 143 -2055
rect 149 -2051 150 -2049
rect 149 -2057 150 -2055
rect 156 -2051 157 -2049
rect 159 -2051 160 -2049
rect 156 -2057 157 -2055
rect 163 -2051 164 -2049
rect 166 -2051 167 -2049
rect 163 -2057 164 -2055
rect 166 -2057 167 -2055
rect 170 -2051 171 -2049
rect 170 -2057 171 -2055
rect 177 -2051 178 -2049
rect 177 -2057 178 -2055
rect 184 -2051 185 -2049
rect 184 -2057 185 -2055
rect 191 -2051 192 -2049
rect 191 -2057 192 -2055
rect 198 -2051 199 -2049
rect 198 -2057 199 -2055
rect 205 -2051 206 -2049
rect 208 -2051 209 -2049
rect 205 -2057 206 -2055
rect 208 -2057 209 -2055
rect 212 -2051 213 -2049
rect 212 -2057 213 -2055
rect 219 -2051 220 -2049
rect 219 -2057 220 -2055
rect 226 -2051 227 -2049
rect 226 -2057 227 -2055
rect 233 -2051 234 -2049
rect 233 -2057 234 -2055
rect 240 -2051 241 -2049
rect 240 -2057 241 -2055
rect 247 -2051 248 -2049
rect 247 -2057 248 -2055
rect 254 -2051 255 -2049
rect 254 -2057 255 -2055
rect 261 -2051 262 -2049
rect 261 -2057 262 -2055
rect 268 -2051 269 -2049
rect 268 -2057 269 -2055
rect 275 -2051 276 -2049
rect 275 -2057 276 -2055
rect 282 -2051 283 -2049
rect 282 -2057 283 -2055
rect 289 -2051 290 -2049
rect 289 -2057 290 -2055
rect 296 -2051 297 -2049
rect 296 -2057 297 -2055
rect 303 -2051 304 -2049
rect 303 -2057 304 -2055
rect 310 -2051 311 -2049
rect 310 -2057 311 -2055
rect 317 -2051 318 -2049
rect 317 -2057 318 -2055
rect 324 -2051 325 -2049
rect 324 -2057 325 -2055
rect 331 -2051 332 -2049
rect 331 -2057 332 -2055
rect 338 -2051 339 -2049
rect 338 -2057 339 -2055
rect 345 -2051 346 -2049
rect 345 -2057 346 -2055
rect 352 -2051 353 -2049
rect 352 -2057 353 -2055
rect 359 -2051 360 -2049
rect 359 -2057 360 -2055
rect 369 -2051 370 -2049
rect 366 -2057 367 -2055
rect 369 -2057 370 -2055
rect 373 -2051 374 -2049
rect 373 -2057 374 -2055
rect 380 -2051 381 -2049
rect 380 -2057 381 -2055
rect 387 -2051 388 -2049
rect 387 -2057 388 -2055
rect 394 -2051 395 -2049
rect 394 -2057 395 -2055
rect 401 -2051 402 -2049
rect 401 -2057 402 -2055
rect 408 -2051 409 -2049
rect 408 -2057 409 -2055
rect 415 -2051 416 -2049
rect 415 -2057 416 -2055
rect 422 -2051 423 -2049
rect 422 -2057 423 -2055
rect 429 -2051 430 -2049
rect 429 -2057 430 -2055
rect 436 -2051 437 -2049
rect 436 -2057 437 -2055
rect 443 -2051 444 -2049
rect 443 -2057 444 -2055
rect 450 -2051 451 -2049
rect 450 -2057 451 -2055
rect 457 -2051 458 -2049
rect 457 -2057 458 -2055
rect 464 -2051 465 -2049
rect 464 -2057 465 -2055
rect 471 -2051 472 -2049
rect 471 -2057 472 -2055
rect 478 -2051 479 -2049
rect 478 -2057 479 -2055
rect 485 -2051 486 -2049
rect 485 -2057 486 -2055
rect 492 -2051 493 -2049
rect 492 -2057 493 -2055
rect 499 -2051 500 -2049
rect 499 -2057 500 -2055
rect 506 -2051 507 -2049
rect 506 -2057 507 -2055
rect 513 -2051 514 -2049
rect 513 -2057 514 -2055
rect 520 -2051 521 -2049
rect 520 -2057 521 -2055
rect 530 -2051 531 -2049
rect 530 -2057 531 -2055
rect 534 -2051 535 -2049
rect 534 -2057 535 -2055
rect 541 -2051 542 -2049
rect 541 -2057 542 -2055
rect 548 -2051 549 -2049
rect 548 -2057 549 -2055
rect 555 -2051 556 -2049
rect 555 -2057 556 -2055
rect 562 -2051 563 -2049
rect 562 -2057 563 -2055
rect 569 -2051 570 -2049
rect 569 -2057 570 -2055
rect 576 -2051 577 -2049
rect 576 -2057 577 -2055
rect 583 -2051 584 -2049
rect 583 -2057 584 -2055
rect 590 -2051 591 -2049
rect 593 -2051 594 -2049
rect 593 -2057 594 -2055
rect 597 -2051 598 -2049
rect 600 -2051 601 -2049
rect 600 -2057 601 -2055
rect 604 -2051 605 -2049
rect 607 -2051 608 -2049
rect 607 -2057 608 -2055
rect 611 -2051 612 -2049
rect 611 -2057 612 -2055
rect 618 -2051 619 -2049
rect 621 -2051 622 -2049
rect 618 -2057 619 -2055
rect 621 -2057 622 -2055
rect 625 -2051 626 -2049
rect 625 -2057 626 -2055
rect 632 -2051 633 -2049
rect 635 -2051 636 -2049
rect 632 -2057 633 -2055
rect 635 -2057 636 -2055
rect 639 -2051 640 -2049
rect 639 -2057 640 -2055
rect 646 -2051 647 -2049
rect 646 -2057 647 -2055
rect 653 -2051 654 -2049
rect 653 -2057 654 -2055
rect 660 -2051 661 -2049
rect 663 -2051 664 -2049
rect 660 -2057 661 -2055
rect 663 -2057 664 -2055
rect 667 -2051 668 -2049
rect 670 -2051 671 -2049
rect 667 -2057 668 -2055
rect 670 -2057 671 -2055
rect 674 -2051 675 -2049
rect 674 -2057 675 -2055
rect 681 -2051 682 -2049
rect 681 -2057 682 -2055
rect 688 -2051 689 -2049
rect 691 -2051 692 -2049
rect 688 -2057 689 -2055
rect 691 -2057 692 -2055
rect 695 -2051 696 -2049
rect 695 -2057 696 -2055
rect 702 -2051 703 -2049
rect 702 -2057 703 -2055
rect 709 -2051 710 -2049
rect 709 -2057 710 -2055
rect 716 -2051 717 -2049
rect 716 -2057 717 -2055
rect 723 -2051 724 -2049
rect 723 -2057 724 -2055
rect 730 -2051 731 -2049
rect 730 -2057 731 -2055
rect 737 -2051 738 -2049
rect 737 -2057 738 -2055
rect 744 -2051 745 -2049
rect 744 -2057 745 -2055
rect 751 -2051 752 -2049
rect 754 -2051 755 -2049
rect 751 -2057 752 -2055
rect 754 -2057 755 -2055
rect 758 -2051 759 -2049
rect 758 -2057 759 -2055
rect 765 -2051 766 -2049
rect 768 -2051 769 -2049
rect 765 -2057 766 -2055
rect 772 -2051 773 -2049
rect 772 -2057 773 -2055
rect 782 -2051 783 -2049
rect 779 -2057 780 -2055
rect 782 -2057 783 -2055
rect 786 -2051 787 -2049
rect 786 -2057 787 -2055
rect 793 -2051 794 -2049
rect 793 -2057 794 -2055
rect 800 -2051 801 -2049
rect 803 -2051 804 -2049
rect 800 -2057 801 -2055
rect 803 -2057 804 -2055
rect 807 -2051 808 -2049
rect 807 -2057 808 -2055
rect 814 -2051 815 -2049
rect 817 -2051 818 -2049
rect 814 -2057 815 -2055
rect 817 -2057 818 -2055
rect 821 -2051 822 -2049
rect 821 -2057 822 -2055
rect 828 -2051 829 -2049
rect 828 -2057 829 -2055
rect 835 -2051 836 -2049
rect 835 -2057 836 -2055
rect 842 -2051 843 -2049
rect 842 -2057 843 -2055
rect 849 -2051 850 -2049
rect 849 -2057 850 -2055
rect 856 -2051 857 -2049
rect 856 -2057 857 -2055
rect 863 -2051 864 -2049
rect 863 -2057 864 -2055
rect 870 -2051 871 -2049
rect 870 -2057 871 -2055
rect 877 -2051 878 -2049
rect 877 -2057 878 -2055
rect 884 -2051 885 -2049
rect 884 -2057 885 -2055
rect 891 -2051 892 -2049
rect 891 -2057 892 -2055
rect 898 -2051 899 -2049
rect 898 -2057 899 -2055
rect 905 -2051 906 -2049
rect 908 -2051 909 -2049
rect 905 -2057 906 -2055
rect 908 -2057 909 -2055
rect 912 -2051 913 -2049
rect 912 -2057 913 -2055
rect 919 -2051 920 -2049
rect 919 -2057 920 -2055
rect 926 -2051 927 -2049
rect 929 -2051 930 -2049
rect 926 -2057 927 -2055
rect 933 -2051 934 -2049
rect 936 -2051 937 -2049
rect 933 -2057 934 -2055
rect 936 -2057 937 -2055
rect 940 -2051 941 -2049
rect 950 -2051 951 -2049
rect 947 -2057 948 -2055
rect 950 -2057 951 -2055
rect 954 -2051 955 -2049
rect 954 -2057 955 -2055
rect 961 -2051 962 -2049
rect 961 -2057 962 -2055
rect 968 -2051 969 -2049
rect 968 -2057 969 -2055
rect 975 -2051 976 -2049
rect 975 -2057 976 -2055
rect 985 -2051 986 -2049
rect 982 -2057 983 -2055
rect 985 -2057 986 -2055
rect 989 -2051 990 -2049
rect 989 -2057 990 -2055
rect 996 -2051 997 -2049
rect 996 -2057 997 -2055
rect 1003 -2051 1004 -2049
rect 1003 -2057 1004 -2055
rect 1010 -2051 1011 -2049
rect 1010 -2057 1011 -2055
rect 1017 -2051 1018 -2049
rect 1020 -2051 1021 -2049
rect 1017 -2057 1018 -2055
rect 1020 -2057 1021 -2055
rect 1024 -2051 1025 -2049
rect 1024 -2057 1025 -2055
rect 1031 -2051 1032 -2049
rect 1031 -2057 1032 -2055
rect 1038 -2051 1039 -2049
rect 1038 -2057 1039 -2055
rect 1045 -2051 1046 -2049
rect 1045 -2057 1046 -2055
rect 1052 -2051 1053 -2049
rect 1052 -2057 1053 -2055
rect 1059 -2051 1060 -2049
rect 1059 -2057 1060 -2055
rect 1066 -2051 1067 -2049
rect 1066 -2057 1067 -2055
rect 1073 -2051 1074 -2049
rect 1073 -2057 1074 -2055
rect 1080 -2051 1081 -2049
rect 1080 -2057 1081 -2055
rect 1087 -2051 1088 -2049
rect 1087 -2057 1088 -2055
rect 1090 -2057 1091 -2055
rect 1094 -2051 1095 -2049
rect 1094 -2057 1095 -2055
rect 1101 -2051 1102 -2049
rect 1101 -2057 1102 -2055
rect 1108 -2051 1109 -2049
rect 1108 -2057 1109 -2055
rect 1115 -2051 1116 -2049
rect 1115 -2057 1116 -2055
rect 1122 -2051 1123 -2049
rect 1122 -2057 1123 -2055
rect 1129 -2051 1130 -2049
rect 1129 -2057 1130 -2055
rect 1136 -2051 1137 -2049
rect 1136 -2057 1137 -2055
rect 1143 -2051 1144 -2049
rect 1143 -2057 1144 -2055
rect 1150 -2051 1151 -2049
rect 1150 -2057 1151 -2055
rect 1157 -2051 1158 -2049
rect 1157 -2057 1158 -2055
rect 1164 -2051 1165 -2049
rect 1164 -2057 1165 -2055
rect 1171 -2051 1172 -2049
rect 1171 -2057 1172 -2055
rect 1178 -2051 1179 -2049
rect 1178 -2057 1179 -2055
rect 1185 -2051 1186 -2049
rect 1185 -2057 1186 -2055
rect 1192 -2051 1193 -2049
rect 1192 -2057 1193 -2055
rect 1199 -2051 1200 -2049
rect 1199 -2057 1200 -2055
rect 1206 -2051 1207 -2049
rect 1206 -2057 1207 -2055
rect 1213 -2051 1214 -2049
rect 1213 -2057 1214 -2055
rect 1220 -2051 1221 -2049
rect 1220 -2057 1221 -2055
rect 1227 -2051 1228 -2049
rect 1227 -2057 1228 -2055
rect 1234 -2051 1235 -2049
rect 1234 -2057 1235 -2055
rect 1241 -2051 1242 -2049
rect 1241 -2057 1242 -2055
rect 1248 -2051 1249 -2049
rect 1248 -2057 1249 -2055
rect 1255 -2051 1256 -2049
rect 1258 -2051 1259 -2049
rect 1255 -2057 1256 -2055
rect 1258 -2057 1259 -2055
rect 1262 -2051 1263 -2049
rect 1262 -2057 1263 -2055
rect 1269 -2051 1270 -2049
rect 1269 -2057 1270 -2055
rect 1276 -2051 1277 -2049
rect 1276 -2057 1277 -2055
rect 1283 -2051 1284 -2049
rect 1283 -2057 1284 -2055
rect 1290 -2051 1291 -2049
rect 1290 -2057 1291 -2055
rect 1297 -2051 1298 -2049
rect 1297 -2057 1298 -2055
rect 1304 -2051 1305 -2049
rect 1304 -2057 1305 -2055
rect 1311 -2051 1312 -2049
rect 1311 -2057 1312 -2055
rect 1318 -2051 1319 -2049
rect 1318 -2057 1319 -2055
rect 1325 -2051 1326 -2049
rect 1325 -2057 1326 -2055
rect 1332 -2051 1333 -2049
rect 1332 -2057 1333 -2055
rect 1339 -2051 1340 -2049
rect 1339 -2057 1340 -2055
rect 1346 -2051 1347 -2049
rect 1346 -2057 1347 -2055
rect 1353 -2051 1354 -2049
rect 1353 -2057 1354 -2055
rect 1360 -2051 1361 -2049
rect 1360 -2057 1361 -2055
rect 1367 -2051 1368 -2049
rect 1367 -2057 1368 -2055
rect 1374 -2051 1375 -2049
rect 1374 -2057 1375 -2055
rect 1381 -2051 1382 -2049
rect 1381 -2057 1382 -2055
rect 1388 -2051 1389 -2049
rect 1388 -2057 1389 -2055
rect 1395 -2051 1396 -2049
rect 1395 -2057 1396 -2055
rect 1402 -2051 1403 -2049
rect 1402 -2057 1403 -2055
rect 1409 -2051 1410 -2049
rect 1409 -2057 1410 -2055
rect 1416 -2051 1417 -2049
rect 1416 -2057 1417 -2055
rect 1423 -2051 1424 -2049
rect 1423 -2057 1424 -2055
rect 1430 -2051 1431 -2049
rect 1430 -2057 1431 -2055
rect 1437 -2051 1438 -2049
rect 1437 -2057 1438 -2055
rect 1444 -2051 1445 -2049
rect 1444 -2057 1445 -2055
rect 1451 -2057 1452 -2055
rect 1458 -2051 1459 -2049
rect 1458 -2057 1459 -2055
rect 1465 -2051 1466 -2049
rect 1465 -2057 1466 -2055
rect 1472 -2051 1473 -2049
rect 1472 -2057 1473 -2055
rect 1479 -2051 1480 -2049
rect 1479 -2057 1480 -2055
rect 1486 -2051 1487 -2049
rect 1486 -2057 1487 -2055
rect 1493 -2051 1494 -2049
rect 1493 -2057 1494 -2055
rect 1500 -2051 1501 -2049
rect 1500 -2057 1501 -2055
rect 1507 -2051 1508 -2049
rect 1507 -2057 1508 -2055
rect 1514 -2051 1515 -2049
rect 1514 -2057 1515 -2055
rect 1521 -2051 1522 -2049
rect 1521 -2057 1522 -2055
rect 1528 -2051 1529 -2049
rect 1528 -2057 1529 -2055
rect 1535 -2051 1536 -2049
rect 1535 -2057 1536 -2055
rect 1542 -2051 1543 -2049
rect 1542 -2057 1543 -2055
rect 1549 -2051 1550 -2049
rect 1549 -2057 1550 -2055
rect 1556 -2051 1557 -2049
rect 1556 -2057 1557 -2055
rect 1563 -2051 1564 -2049
rect 1563 -2057 1564 -2055
rect 1570 -2051 1571 -2049
rect 1570 -2057 1571 -2055
rect 1577 -2051 1578 -2049
rect 1577 -2057 1578 -2055
rect 1584 -2051 1585 -2049
rect 1584 -2057 1585 -2055
rect 1591 -2051 1592 -2049
rect 1591 -2057 1592 -2055
rect 1598 -2051 1599 -2049
rect 1598 -2057 1599 -2055
rect 1605 -2051 1606 -2049
rect 1605 -2057 1606 -2055
rect 1612 -2051 1613 -2049
rect 1612 -2057 1613 -2055
rect 1619 -2051 1620 -2049
rect 1619 -2057 1620 -2055
rect 1626 -2051 1627 -2049
rect 1626 -2057 1627 -2055
rect 1629 -2057 1630 -2055
rect 1633 -2051 1634 -2049
rect 1633 -2057 1634 -2055
rect 1640 -2051 1641 -2049
rect 1640 -2057 1641 -2055
rect 1647 -2051 1648 -2049
rect 1647 -2057 1648 -2055
rect 1654 -2051 1655 -2049
rect 1654 -2057 1655 -2055
rect 1661 -2051 1662 -2049
rect 1661 -2057 1662 -2055
rect 1668 -2051 1669 -2049
rect 1668 -2057 1669 -2055
rect 1675 -2051 1676 -2049
rect 1675 -2057 1676 -2055
rect 1682 -2051 1683 -2049
rect 1682 -2057 1683 -2055
rect 1689 -2051 1690 -2049
rect 1689 -2057 1690 -2055
rect 1696 -2051 1697 -2049
rect 1696 -2057 1697 -2055
rect 1703 -2051 1704 -2049
rect 1703 -2057 1704 -2055
rect 1710 -2051 1711 -2049
rect 1710 -2057 1711 -2055
rect 1717 -2051 1718 -2049
rect 1717 -2057 1718 -2055
rect 1724 -2051 1725 -2049
rect 1724 -2057 1725 -2055
rect 1731 -2051 1732 -2049
rect 1731 -2057 1732 -2055
rect 1738 -2051 1739 -2049
rect 1738 -2057 1739 -2055
rect 1745 -2051 1746 -2049
rect 1745 -2057 1746 -2055
rect 1748 -2057 1749 -2055
rect 1752 -2051 1753 -2049
rect 1752 -2057 1753 -2055
rect 1759 -2051 1760 -2049
rect 1762 -2051 1763 -2049
rect 1762 -2057 1763 -2055
rect 1766 -2051 1767 -2049
rect 1766 -2057 1767 -2055
rect 1773 -2051 1774 -2049
rect 1773 -2057 1774 -2055
rect 30 -2190 31 -2188
rect 30 -2196 31 -2194
rect 40 -2190 41 -2188
rect 40 -2196 41 -2194
rect 47 -2190 48 -2188
rect 44 -2196 45 -2194
rect 51 -2190 52 -2188
rect 54 -2190 55 -2188
rect 51 -2196 52 -2194
rect 58 -2190 59 -2188
rect 58 -2196 59 -2194
rect 65 -2190 66 -2188
rect 68 -2190 69 -2188
rect 68 -2196 69 -2194
rect 72 -2190 73 -2188
rect 72 -2196 73 -2194
rect 79 -2190 80 -2188
rect 79 -2196 80 -2194
rect 86 -2190 87 -2188
rect 86 -2196 87 -2194
rect 89 -2196 90 -2194
rect 93 -2190 94 -2188
rect 96 -2190 97 -2188
rect 96 -2196 97 -2194
rect 100 -2190 101 -2188
rect 100 -2196 101 -2194
rect 107 -2190 108 -2188
rect 107 -2196 108 -2194
rect 114 -2190 115 -2188
rect 114 -2196 115 -2194
rect 121 -2190 122 -2188
rect 121 -2196 122 -2194
rect 128 -2190 129 -2188
rect 131 -2190 132 -2188
rect 128 -2196 129 -2194
rect 131 -2196 132 -2194
rect 135 -2190 136 -2188
rect 135 -2196 136 -2194
rect 142 -2190 143 -2188
rect 142 -2196 143 -2194
rect 152 -2190 153 -2188
rect 149 -2196 150 -2194
rect 152 -2196 153 -2194
rect 156 -2190 157 -2188
rect 156 -2196 157 -2194
rect 163 -2190 164 -2188
rect 163 -2196 164 -2194
rect 170 -2190 171 -2188
rect 173 -2190 174 -2188
rect 170 -2196 171 -2194
rect 173 -2196 174 -2194
rect 177 -2190 178 -2188
rect 177 -2196 178 -2194
rect 184 -2190 185 -2188
rect 184 -2196 185 -2194
rect 191 -2190 192 -2188
rect 191 -2196 192 -2194
rect 198 -2190 199 -2188
rect 198 -2196 199 -2194
rect 205 -2190 206 -2188
rect 205 -2196 206 -2194
rect 212 -2190 213 -2188
rect 212 -2196 213 -2194
rect 219 -2190 220 -2188
rect 219 -2196 220 -2194
rect 226 -2190 227 -2188
rect 229 -2190 230 -2188
rect 229 -2196 230 -2194
rect 233 -2190 234 -2188
rect 233 -2196 234 -2194
rect 240 -2190 241 -2188
rect 240 -2196 241 -2194
rect 247 -2190 248 -2188
rect 247 -2196 248 -2194
rect 254 -2190 255 -2188
rect 254 -2196 255 -2194
rect 261 -2190 262 -2188
rect 261 -2196 262 -2194
rect 271 -2196 272 -2194
rect 275 -2190 276 -2188
rect 275 -2196 276 -2194
rect 282 -2190 283 -2188
rect 282 -2196 283 -2194
rect 289 -2190 290 -2188
rect 289 -2196 290 -2194
rect 296 -2190 297 -2188
rect 296 -2196 297 -2194
rect 303 -2190 304 -2188
rect 303 -2196 304 -2194
rect 310 -2190 311 -2188
rect 310 -2196 311 -2194
rect 317 -2190 318 -2188
rect 317 -2196 318 -2194
rect 324 -2190 325 -2188
rect 324 -2196 325 -2194
rect 331 -2190 332 -2188
rect 331 -2196 332 -2194
rect 338 -2190 339 -2188
rect 338 -2196 339 -2194
rect 345 -2190 346 -2188
rect 345 -2196 346 -2194
rect 352 -2190 353 -2188
rect 352 -2196 353 -2194
rect 359 -2190 360 -2188
rect 362 -2190 363 -2188
rect 359 -2196 360 -2194
rect 362 -2196 363 -2194
rect 366 -2190 367 -2188
rect 366 -2196 367 -2194
rect 373 -2190 374 -2188
rect 373 -2196 374 -2194
rect 380 -2190 381 -2188
rect 380 -2196 381 -2194
rect 387 -2190 388 -2188
rect 387 -2196 388 -2194
rect 394 -2190 395 -2188
rect 394 -2196 395 -2194
rect 401 -2190 402 -2188
rect 401 -2196 402 -2194
rect 408 -2190 409 -2188
rect 415 -2190 416 -2188
rect 415 -2196 416 -2194
rect 422 -2190 423 -2188
rect 422 -2196 423 -2194
rect 429 -2190 430 -2188
rect 429 -2196 430 -2194
rect 436 -2190 437 -2188
rect 436 -2196 437 -2194
rect 443 -2190 444 -2188
rect 443 -2196 444 -2194
rect 450 -2190 451 -2188
rect 453 -2190 454 -2188
rect 450 -2196 451 -2194
rect 453 -2196 454 -2194
rect 457 -2190 458 -2188
rect 457 -2196 458 -2194
rect 464 -2190 465 -2188
rect 464 -2196 465 -2194
rect 471 -2190 472 -2188
rect 471 -2196 472 -2194
rect 478 -2190 479 -2188
rect 478 -2196 479 -2194
rect 485 -2190 486 -2188
rect 485 -2196 486 -2194
rect 492 -2190 493 -2188
rect 492 -2196 493 -2194
rect 499 -2190 500 -2188
rect 499 -2196 500 -2194
rect 506 -2190 507 -2188
rect 506 -2196 507 -2194
rect 513 -2190 514 -2188
rect 513 -2196 514 -2194
rect 520 -2190 521 -2188
rect 520 -2196 521 -2194
rect 523 -2196 524 -2194
rect 527 -2190 528 -2188
rect 527 -2196 528 -2194
rect 534 -2190 535 -2188
rect 534 -2196 535 -2194
rect 541 -2190 542 -2188
rect 541 -2196 542 -2194
rect 548 -2190 549 -2188
rect 548 -2196 549 -2194
rect 555 -2190 556 -2188
rect 555 -2196 556 -2194
rect 562 -2190 563 -2188
rect 562 -2196 563 -2194
rect 569 -2190 570 -2188
rect 569 -2196 570 -2194
rect 576 -2190 577 -2188
rect 576 -2196 577 -2194
rect 583 -2190 584 -2188
rect 583 -2196 584 -2194
rect 590 -2190 591 -2188
rect 590 -2196 591 -2194
rect 597 -2190 598 -2188
rect 597 -2196 598 -2194
rect 604 -2196 605 -2194
rect 607 -2196 608 -2194
rect 611 -2190 612 -2188
rect 611 -2196 612 -2194
rect 618 -2190 619 -2188
rect 621 -2190 622 -2188
rect 618 -2196 619 -2194
rect 625 -2190 626 -2188
rect 625 -2196 626 -2194
rect 632 -2190 633 -2188
rect 632 -2196 633 -2194
rect 639 -2190 640 -2188
rect 639 -2196 640 -2194
rect 646 -2190 647 -2188
rect 646 -2196 647 -2194
rect 653 -2190 654 -2188
rect 653 -2196 654 -2194
rect 660 -2190 661 -2188
rect 660 -2196 661 -2194
rect 667 -2190 668 -2188
rect 667 -2196 668 -2194
rect 674 -2190 675 -2188
rect 674 -2196 675 -2194
rect 681 -2190 682 -2188
rect 681 -2196 682 -2194
rect 688 -2190 689 -2188
rect 688 -2196 689 -2194
rect 695 -2190 696 -2188
rect 695 -2196 696 -2194
rect 702 -2190 703 -2188
rect 705 -2190 706 -2188
rect 702 -2196 703 -2194
rect 705 -2196 706 -2194
rect 709 -2190 710 -2188
rect 709 -2196 710 -2194
rect 716 -2190 717 -2188
rect 716 -2196 717 -2194
rect 723 -2190 724 -2188
rect 726 -2190 727 -2188
rect 723 -2196 724 -2194
rect 730 -2190 731 -2188
rect 733 -2190 734 -2188
rect 730 -2196 731 -2194
rect 733 -2196 734 -2194
rect 737 -2190 738 -2188
rect 737 -2196 738 -2194
rect 744 -2190 745 -2188
rect 747 -2190 748 -2188
rect 744 -2196 745 -2194
rect 747 -2196 748 -2194
rect 751 -2190 752 -2188
rect 751 -2196 752 -2194
rect 758 -2190 759 -2188
rect 761 -2190 762 -2188
rect 761 -2196 762 -2194
rect 765 -2190 766 -2188
rect 765 -2196 766 -2194
rect 772 -2190 773 -2188
rect 772 -2196 773 -2194
rect 775 -2196 776 -2194
rect 779 -2190 780 -2188
rect 779 -2196 780 -2194
rect 786 -2190 787 -2188
rect 786 -2196 787 -2194
rect 793 -2196 794 -2194
rect 796 -2196 797 -2194
rect 800 -2190 801 -2188
rect 800 -2196 801 -2194
rect 807 -2190 808 -2188
rect 807 -2196 808 -2194
rect 814 -2190 815 -2188
rect 817 -2190 818 -2188
rect 814 -2196 815 -2194
rect 821 -2190 822 -2188
rect 821 -2196 822 -2194
rect 831 -2190 832 -2188
rect 828 -2196 829 -2194
rect 831 -2196 832 -2194
rect 835 -2190 836 -2188
rect 835 -2196 836 -2194
rect 842 -2190 843 -2188
rect 842 -2196 843 -2194
rect 849 -2190 850 -2188
rect 849 -2196 850 -2194
rect 856 -2190 857 -2188
rect 856 -2196 857 -2194
rect 863 -2190 864 -2188
rect 863 -2196 864 -2194
rect 873 -2190 874 -2188
rect 870 -2196 871 -2194
rect 873 -2196 874 -2194
rect 877 -2190 878 -2188
rect 877 -2196 878 -2194
rect 884 -2190 885 -2188
rect 884 -2196 885 -2194
rect 891 -2190 892 -2188
rect 891 -2196 892 -2194
rect 898 -2190 899 -2188
rect 898 -2196 899 -2194
rect 905 -2190 906 -2188
rect 905 -2196 906 -2194
rect 912 -2190 913 -2188
rect 912 -2196 913 -2194
rect 919 -2190 920 -2188
rect 919 -2196 920 -2194
rect 926 -2190 927 -2188
rect 926 -2196 927 -2194
rect 933 -2190 934 -2188
rect 936 -2190 937 -2188
rect 933 -2196 934 -2194
rect 936 -2196 937 -2194
rect 940 -2196 941 -2194
rect 947 -2190 948 -2188
rect 947 -2196 948 -2194
rect 954 -2190 955 -2188
rect 954 -2196 955 -2194
rect 961 -2190 962 -2188
rect 961 -2196 962 -2194
rect 968 -2190 969 -2188
rect 968 -2196 969 -2194
rect 978 -2190 979 -2188
rect 975 -2196 976 -2194
rect 978 -2196 979 -2194
rect 982 -2190 983 -2188
rect 982 -2196 983 -2194
rect 989 -2190 990 -2188
rect 989 -2196 990 -2194
rect 996 -2190 997 -2188
rect 996 -2196 997 -2194
rect 999 -2196 1000 -2194
rect 1003 -2190 1004 -2188
rect 1003 -2196 1004 -2194
rect 1013 -2190 1014 -2188
rect 1010 -2196 1011 -2194
rect 1013 -2196 1014 -2194
rect 1017 -2190 1018 -2188
rect 1017 -2196 1018 -2194
rect 1024 -2190 1025 -2188
rect 1024 -2196 1025 -2194
rect 1031 -2190 1032 -2188
rect 1031 -2196 1032 -2194
rect 1038 -2190 1039 -2188
rect 1038 -2196 1039 -2194
rect 1045 -2190 1046 -2188
rect 1045 -2196 1046 -2194
rect 1052 -2190 1053 -2188
rect 1052 -2196 1053 -2194
rect 1059 -2190 1060 -2188
rect 1059 -2196 1060 -2194
rect 1066 -2190 1067 -2188
rect 1066 -2196 1067 -2194
rect 1073 -2190 1074 -2188
rect 1073 -2196 1074 -2194
rect 1080 -2190 1081 -2188
rect 1080 -2196 1081 -2194
rect 1087 -2190 1088 -2188
rect 1087 -2196 1088 -2194
rect 1094 -2190 1095 -2188
rect 1094 -2196 1095 -2194
rect 1104 -2190 1105 -2188
rect 1101 -2196 1102 -2194
rect 1104 -2196 1105 -2194
rect 1108 -2190 1109 -2188
rect 1108 -2196 1109 -2194
rect 1115 -2190 1116 -2188
rect 1118 -2190 1119 -2188
rect 1115 -2196 1116 -2194
rect 1118 -2196 1119 -2194
rect 1122 -2190 1123 -2188
rect 1122 -2196 1123 -2194
rect 1129 -2190 1130 -2188
rect 1129 -2196 1130 -2194
rect 1136 -2190 1137 -2188
rect 1136 -2196 1137 -2194
rect 1143 -2190 1144 -2188
rect 1143 -2196 1144 -2194
rect 1150 -2190 1151 -2188
rect 1150 -2196 1151 -2194
rect 1157 -2190 1158 -2188
rect 1157 -2196 1158 -2194
rect 1164 -2190 1165 -2188
rect 1164 -2196 1165 -2194
rect 1171 -2190 1172 -2188
rect 1171 -2196 1172 -2194
rect 1178 -2190 1179 -2188
rect 1178 -2196 1179 -2194
rect 1185 -2190 1186 -2188
rect 1185 -2196 1186 -2194
rect 1192 -2190 1193 -2188
rect 1192 -2196 1193 -2194
rect 1199 -2190 1200 -2188
rect 1199 -2196 1200 -2194
rect 1206 -2190 1207 -2188
rect 1206 -2196 1207 -2194
rect 1213 -2190 1214 -2188
rect 1213 -2196 1214 -2194
rect 1220 -2190 1221 -2188
rect 1220 -2196 1221 -2194
rect 1227 -2190 1228 -2188
rect 1227 -2196 1228 -2194
rect 1234 -2190 1235 -2188
rect 1234 -2196 1235 -2194
rect 1241 -2190 1242 -2188
rect 1241 -2196 1242 -2194
rect 1248 -2190 1249 -2188
rect 1248 -2196 1249 -2194
rect 1255 -2190 1256 -2188
rect 1255 -2196 1256 -2194
rect 1262 -2190 1263 -2188
rect 1262 -2196 1263 -2194
rect 1269 -2190 1270 -2188
rect 1269 -2196 1270 -2194
rect 1276 -2190 1277 -2188
rect 1276 -2196 1277 -2194
rect 1283 -2190 1284 -2188
rect 1283 -2196 1284 -2194
rect 1290 -2190 1291 -2188
rect 1290 -2196 1291 -2194
rect 1297 -2190 1298 -2188
rect 1297 -2196 1298 -2194
rect 1304 -2190 1305 -2188
rect 1304 -2196 1305 -2194
rect 1311 -2190 1312 -2188
rect 1311 -2196 1312 -2194
rect 1318 -2190 1319 -2188
rect 1318 -2196 1319 -2194
rect 1325 -2190 1326 -2188
rect 1325 -2196 1326 -2194
rect 1332 -2190 1333 -2188
rect 1332 -2196 1333 -2194
rect 1339 -2190 1340 -2188
rect 1339 -2196 1340 -2194
rect 1346 -2190 1347 -2188
rect 1346 -2196 1347 -2194
rect 1353 -2190 1354 -2188
rect 1353 -2196 1354 -2194
rect 1360 -2190 1361 -2188
rect 1360 -2196 1361 -2194
rect 1367 -2190 1368 -2188
rect 1367 -2196 1368 -2194
rect 1374 -2190 1375 -2188
rect 1374 -2196 1375 -2194
rect 1381 -2190 1382 -2188
rect 1381 -2196 1382 -2194
rect 1388 -2190 1389 -2188
rect 1388 -2196 1389 -2194
rect 1395 -2190 1396 -2188
rect 1395 -2196 1396 -2194
rect 1402 -2190 1403 -2188
rect 1402 -2196 1403 -2194
rect 1409 -2190 1410 -2188
rect 1409 -2196 1410 -2194
rect 1416 -2190 1417 -2188
rect 1416 -2196 1417 -2194
rect 1423 -2190 1424 -2188
rect 1423 -2196 1424 -2194
rect 1430 -2190 1431 -2188
rect 1430 -2196 1431 -2194
rect 1437 -2190 1438 -2188
rect 1437 -2196 1438 -2194
rect 1444 -2190 1445 -2188
rect 1444 -2196 1445 -2194
rect 1451 -2190 1452 -2188
rect 1451 -2196 1452 -2194
rect 1458 -2190 1459 -2188
rect 1458 -2196 1459 -2194
rect 1465 -2190 1466 -2188
rect 1465 -2196 1466 -2194
rect 1472 -2190 1473 -2188
rect 1472 -2196 1473 -2194
rect 1479 -2190 1480 -2188
rect 1479 -2196 1480 -2194
rect 1486 -2190 1487 -2188
rect 1486 -2196 1487 -2194
rect 1493 -2190 1494 -2188
rect 1493 -2196 1494 -2194
rect 1500 -2190 1501 -2188
rect 1500 -2196 1501 -2194
rect 1507 -2190 1508 -2188
rect 1507 -2196 1508 -2194
rect 1514 -2190 1515 -2188
rect 1514 -2196 1515 -2194
rect 1521 -2190 1522 -2188
rect 1521 -2196 1522 -2194
rect 1528 -2190 1529 -2188
rect 1528 -2196 1529 -2194
rect 1535 -2190 1536 -2188
rect 1535 -2196 1536 -2194
rect 1542 -2190 1543 -2188
rect 1542 -2196 1543 -2194
rect 1549 -2190 1550 -2188
rect 1549 -2196 1550 -2194
rect 1556 -2190 1557 -2188
rect 1556 -2196 1557 -2194
rect 1563 -2190 1564 -2188
rect 1563 -2196 1564 -2194
rect 1570 -2190 1571 -2188
rect 1570 -2196 1571 -2194
rect 1577 -2190 1578 -2188
rect 1577 -2196 1578 -2194
rect 1584 -2190 1585 -2188
rect 1584 -2196 1585 -2194
rect 1591 -2190 1592 -2188
rect 1591 -2196 1592 -2194
rect 1598 -2190 1599 -2188
rect 1598 -2196 1599 -2194
rect 1605 -2190 1606 -2188
rect 1605 -2196 1606 -2194
rect 1612 -2190 1613 -2188
rect 1612 -2196 1613 -2194
rect 1619 -2190 1620 -2188
rect 1619 -2196 1620 -2194
rect 1626 -2190 1627 -2188
rect 1629 -2190 1630 -2188
rect 1626 -2196 1627 -2194
rect 1633 -2190 1634 -2188
rect 1633 -2196 1634 -2194
rect 1640 -2190 1641 -2188
rect 1640 -2196 1641 -2194
rect 1647 -2190 1648 -2188
rect 1647 -2196 1648 -2194
rect 1654 -2190 1655 -2188
rect 1654 -2196 1655 -2194
rect 1661 -2190 1662 -2188
rect 1661 -2196 1662 -2194
rect 1668 -2190 1669 -2188
rect 1668 -2196 1669 -2194
rect 1675 -2190 1676 -2188
rect 1675 -2196 1676 -2194
rect 1682 -2190 1683 -2188
rect 1682 -2196 1683 -2194
rect 1689 -2190 1690 -2188
rect 1689 -2196 1690 -2194
rect 1696 -2190 1697 -2188
rect 1696 -2196 1697 -2194
rect 1703 -2190 1704 -2188
rect 1703 -2196 1704 -2194
rect 1710 -2190 1711 -2188
rect 1710 -2196 1711 -2194
rect 1717 -2190 1718 -2188
rect 1717 -2196 1718 -2194
rect 1724 -2190 1725 -2188
rect 1724 -2196 1725 -2194
rect 1731 -2190 1732 -2188
rect 1731 -2196 1732 -2194
rect 1738 -2190 1739 -2188
rect 1738 -2196 1739 -2194
rect 1745 -2190 1746 -2188
rect 1745 -2196 1746 -2194
rect 1755 -2190 1756 -2188
rect 1752 -2196 1753 -2194
rect 1755 -2196 1756 -2194
rect 1759 -2190 1760 -2188
rect 1759 -2196 1760 -2194
rect 1766 -2190 1767 -2188
rect 1766 -2196 1767 -2194
rect 44 -2325 45 -2323
rect 44 -2331 45 -2329
rect 51 -2325 52 -2323
rect 51 -2331 52 -2329
rect 58 -2325 59 -2323
rect 58 -2331 59 -2329
rect 65 -2325 66 -2323
rect 65 -2331 66 -2329
rect 72 -2325 73 -2323
rect 72 -2331 73 -2329
rect 79 -2325 80 -2323
rect 79 -2331 80 -2329
rect 89 -2325 90 -2323
rect 86 -2331 87 -2329
rect 93 -2325 94 -2323
rect 96 -2325 97 -2323
rect 93 -2331 94 -2329
rect 96 -2331 97 -2329
rect 100 -2325 101 -2323
rect 100 -2331 101 -2329
rect 107 -2325 108 -2323
rect 107 -2331 108 -2329
rect 114 -2325 115 -2323
rect 117 -2325 118 -2323
rect 114 -2331 115 -2329
rect 117 -2331 118 -2329
rect 121 -2325 122 -2323
rect 121 -2331 122 -2329
rect 128 -2325 129 -2323
rect 128 -2331 129 -2329
rect 135 -2325 136 -2323
rect 138 -2325 139 -2323
rect 135 -2331 136 -2329
rect 138 -2331 139 -2329
rect 142 -2325 143 -2323
rect 142 -2331 143 -2329
rect 149 -2325 150 -2323
rect 149 -2331 150 -2329
rect 156 -2325 157 -2323
rect 156 -2331 157 -2329
rect 163 -2325 164 -2323
rect 163 -2331 164 -2329
rect 170 -2325 171 -2323
rect 173 -2325 174 -2323
rect 170 -2331 171 -2329
rect 173 -2331 174 -2329
rect 177 -2325 178 -2323
rect 177 -2331 178 -2329
rect 184 -2325 185 -2323
rect 184 -2331 185 -2329
rect 191 -2325 192 -2323
rect 191 -2331 192 -2329
rect 198 -2325 199 -2323
rect 198 -2331 199 -2329
rect 205 -2325 206 -2323
rect 205 -2331 206 -2329
rect 215 -2325 216 -2323
rect 212 -2331 213 -2329
rect 215 -2331 216 -2329
rect 219 -2325 220 -2323
rect 219 -2331 220 -2329
rect 226 -2325 227 -2323
rect 226 -2331 227 -2329
rect 233 -2325 234 -2323
rect 236 -2325 237 -2323
rect 236 -2331 237 -2329
rect 240 -2325 241 -2323
rect 240 -2331 241 -2329
rect 247 -2325 248 -2323
rect 247 -2331 248 -2329
rect 254 -2325 255 -2323
rect 254 -2331 255 -2329
rect 261 -2325 262 -2323
rect 261 -2331 262 -2329
rect 268 -2325 269 -2323
rect 268 -2331 269 -2329
rect 275 -2325 276 -2323
rect 275 -2331 276 -2329
rect 282 -2325 283 -2323
rect 282 -2331 283 -2329
rect 289 -2325 290 -2323
rect 289 -2331 290 -2329
rect 296 -2325 297 -2323
rect 296 -2331 297 -2329
rect 303 -2325 304 -2323
rect 303 -2331 304 -2329
rect 310 -2325 311 -2323
rect 310 -2331 311 -2329
rect 317 -2325 318 -2323
rect 317 -2331 318 -2329
rect 324 -2325 325 -2323
rect 324 -2331 325 -2329
rect 331 -2325 332 -2323
rect 331 -2331 332 -2329
rect 338 -2325 339 -2323
rect 338 -2331 339 -2329
rect 345 -2325 346 -2323
rect 345 -2331 346 -2329
rect 352 -2325 353 -2323
rect 352 -2331 353 -2329
rect 359 -2325 360 -2323
rect 359 -2331 360 -2329
rect 366 -2325 367 -2323
rect 366 -2331 367 -2329
rect 373 -2325 374 -2323
rect 373 -2331 374 -2329
rect 380 -2325 381 -2323
rect 380 -2331 381 -2329
rect 387 -2325 388 -2323
rect 387 -2331 388 -2329
rect 394 -2325 395 -2323
rect 394 -2331 395 -2329
rect 401 -2325 402 -2323
rect 401 -2331 402 -2329
rect 408 -2325 409 -2323
rect 408 -2331 409 -2329
rect 415 -2325 416 -2323
rect 415 -2331 416 -2329
rect 422 -2325 423 -2323
rect 422 -2331 423 -2329
rect 429 -2325 430 -2323
rect 429 -2331 430 -2329
rect 436 -2325 437 -2323
rect 436 -2331 437 -2329
rect 443 -2325 444 -2323
rect 443 -2331 444 -2329
rect 450 -2325 451 -2323
rect 450 -2331 451 -2329
rect 457 -2325 458 -2323
rect 457 -2331 458 -2329
rect 464 -2325 465 -2323
rect 464 -2331 465 -2329
rect 471 -2325 472 -2323
rect 471 -2331 472 -2329
rect 478 -2325 479 -2323
rect 478 -2331 479 -2329
rect 485 -2325 486 -2323
rect 485 -2331 486 -2329
rect 492 -2325 493 -2323
rect 492 -2331 493 -2329
rect 499 -2325 500 -2323
rect 499 -2331 500 -2329
rect 506 -2325 507 -2323
rect 506 -2331 507 -2329
rect 513 -2325 514 -2323
rect 513 -2331 514 -2329
rect 520 -2325 521 -2323
rect 520 -2331 521 -2329
rect 527 -2325 528 -2323
rect 527 -2331 528 -2329
rect 534 -2325 535 -2323
rect 534 -2331 535 -2329
rect 537 -2331 538 -2329
rect 541 -2325 542 -2323
rect 541 -2331 542 -2329
rect 548 -2325 549 -2323
rect 548 -2331 549 -2329
rect 555 -2325 556 -2323
rect 555 -2331 556 -2329
rect 562 -2325 563 -2323
rect 562 -2331 563 -2329
rect 569 -2325 570 -2323
rect 569 -2331 570 -2329
rect 576 -2325 577 -2323
rect 576 -2331 577 -2329
rect 583 -2325 584 -2323
rect 586 -2325 587 -2323
rect 583 -2331 584 -2329
rect 590 -2325 591 -2323
rect 590 -2331 591 -2329
rect 597 -2325 598 -2323
rect 597 -2331 598 -2329
rect 604 -2325 605 -2323
rect 604 -2331 605 -2329
rect 611 -2325 612 -2323
rect 611 -2331 612 -2329
rect 618 -2325 619 -2323
rect 618 -2331 619 -2329
rect 625 -2325 626 -2323
rect 625 -2331 626 -2329
rect 632 -2325 633 -2323
rect 632 -2331 633 -2329
rect 639 -2325 640 -2323
rect 642 -2331 643 -2329
rect 646 -2325 647 -2323
rect 646 -2331 647 -2329
rect 653 -2325 654 -2323
rect 656 -2325 657 -2323
rect 653 -2331 654 -2329
rect 656 -2331 657 -2329
rect 660 -2325 661 -2323
rect 660 -2331 661 -2329
rect 667 -2325 668 -2323
rect 667 -2331 668 -2329
rect 674 -2325 675 -2323
rect 674 -2331 675 -2329
rect 681 -2325 682 -2323
rect 681 -2331 682 -2329
rect 688 -2325 689 -2323
rect 691 -2325 692 -2323
rect 688 -2331 689 -2329
rect 691 -2331 692 -2329
rect 695 -2325 696 -2323
rect 695 -2331 696 -2329
rect 702 -2325 703 -2323
rect 705 -2325 706 -2323
rect 702 -2331 703 -2329
rect 705 -2331 706 -2329
rect 709 -2325 710 -2323
rect 709 -2331 710 -2329
rect 716 -2325 717 -2323
rect 716 -2331 717 -2329
rect 723 -2325 724 -2323
rect 723 -2331 724 -2329
rect 730 -2325 731 -2323
rect 733 -2325 734 -2323
rect 730 -2331 731 -2329
rect 733 -2331 734 -2329
rect 737 -2325 738 -2323
rect 737 -2331 738 -2329
rect 744 -2325 745 -2323
rect 747 -2325 748 -2323
rect 744 -2331 745 -2329
rect 747 -2331 748 -2329
rect 751 -2325 752 -2323
rect 751 -2331 752 -2329
rect 758 -2325 759 -2323
rect 758 -2331 759 -2329
rect 765 -2325 766 -2323
rect 765 -2331 766 -2329
rect 772 -2325 773 -2323
rect 772 -2331 773 -2329
rect 775 -2331 776 -2329
rect 779 -2325 780 -2323
rect 779 -2331 780 -2329
rect 786 -2325 787 -2323
rect 786 -2331 787 -2329
rect 793 -2325 794 -2323
rect 793 -2331 794 -2329
rect 800 -2325 801 -2323
rect 800 -2331 801 -2329
rect 807 -2325 808 -2323
rect 807 -2331 808 -2329
rect 814 -2325 815 -2323
rect 814 -2331 815 -2329
rect 821 -2325 822 -2323
rect 821 -2331 822 -2329
rect 828 -2325 829 -2323
rect 828 -2331 829 -2329
rect 835 -2325 836 -2323
rect 835 -2331 836 -2329
rect 842 -2325 843 -2323
rect 842 -2331 843 -2329
rect 849 -2325 850 -2323
rect 852 -2325 853 -2323
rect 849 -2331 850 -2329
rect 856 -2325 857 -2323
rect 856 -2331 857 -2329
rect 863 -2325 864 -2323
rect 863 -2331 864 -2329
rect 870 -2325 871 -2323
rect 873 -2325 874 -2323
rect 873 -2331 874 -2329
rect 877 -2325 878 -2323
rect 877 -2331 878 -2329
rect 884 -2325 885 -2323
rect 884 -2331 885 -2329
rect 891 -2325 892 -2323
rect 891 -2331 892 -2329
rect 898 -2325 899 -2323
rect 901 -2325 902 -2323
rect 898 -2331 899 -2329
rect 901 -2331 902 -2329
rect 905 -2325 906 -2323
rect 905 -2331 906 -2329
rect 912 -2325 913 -2323
rect 912 -2331 913 -2329
rect 919 -2325 920 -2323
rect 919 -2331 920 -2329
rect 926 -2325 927 -2323
rect 926 -2331 927 -2329
rect 933 -2325 934 -2323
rect 933 -2331 934 -2329
rect 940 -2325 941 -2323
rect 940 -2331 941 -2329
rect 947 -2325 948 -2323
rect 947 -2331 948 -2329
rect 954 -2325 955 -2323
rect 957 -2325 958 -2323
rect 954 -2331 955 -2329
rect 957 -2331 958 -2329
rect 961 -2325 962 -2323
rect 961 -2331 962 -2329
rect 968 -2325 969 -2323
rect 971 -2331 972 -2329
rect 975 -2325 976 -2323
rect 975 -2331 976 -2329
rect 982 -2325 983 -2323
rect 982 -2331 983 -2329
rect 989 -2325 990 -2323
rect 989 -2331 990 -2329
rect 996 -2325 997 -2323
rect 999 -2325 1000 -2323
rect 996 -2331 997 -2329
rect 999 -2331 1000 -2329
rect 1003 -2325 1004 -2323
rect 1003 -2331 1004 -2329
rect 1010 -2325 1011 -2323
rect 1010 -2331 1011 -2329
rect 1017 -2325 1018 -2323
rect 1017 -2331 1018 -2329
rect 1024 -2325 1025 -2323
rect 1024 -2331 1025 -2329
rect 1031 -2325 1032 -2323
rect 1031 -2331 1032 -2329
rect 1038 -2325 1039 -2323
rect 1038 -2331 1039 -2329
rect 1045 -2325 1046 -2323
rect 1045 -2331 1046 -2329
rect 1052 -2325 1053 -2323
rect 1052 -2331 1053 -2329
rect 1059 -2325 1060 -2323
rect 1059 -2331 1060 -2329
rect 1066 -2325 1067 -2323
rect 1066 -2331 1067 -2329
rect 1073 -2325 1074 -2323
rect 1073 -2331 1074 -2329
rect 1083 -2325 1084 -2323
rect 1080 -2331 1081 -2329
rect 1083 -2331 1084 -2329
rect 1087 -2325 1088 -2323
rect 1087 -2331 1088 -2329
rect 1094 -2325 1095 -2323
rect 1094 -2331 1095 -2329
rect 1097 -2331 1098 -2329
rect 1101 -2325 1102 -2323
rect 1101 -2331 1102 -2329
rect 1108 -2325 1109 -2323
rect 1108 -2331 1109 -2329
rect 1115 -2325 1116 -2323
rect 1115 -2331 1116 -2329
rect 1122 -2325 1123 -2323
rect 1122 -2331 1123 -2329
rect 1125 -2331 1126 -2329
rect 1129 -2325 1130 -2323
rect 1129 -2331 1130 -2329
rect 1136 -2325 1137 -2323
rect 1136 -2331 1137 -2329
rect 1143 -2325 1144 -2323
rect 1146 -2325 1147 -2323
rect 1143 -2331 1144 -2329
rect 1146 -2331 1147 -2329
rect 1150 -2325 1151 -2323
rect 1150 -2331 1151 -2329
rect 1157 -2325 1158 -2323
rect 1157 -2331 1158 -2329
rect 1164 -2325 1165 -2323
rect 1164 -2331 1165 -2329
rect 1171 -2331 1172 -2329
rect 1178 -2325 1179 -2323
rect 1178 -2331 1179 -2329
rect 1185 -2325 1186 -2323
rect 1185 -2331 1186 -2329
rect 1192 -2325 1193 -2323
rect 1192 -2331 1193 -2329
rect 1199 -2325 1200 -2323
rect 1199 -2331 1200 -2329
rect 1206 -2325 1207 -2323
rect 1206 -2331 1207 -2329
rect 1213 -2325 1214 -2323
rect 1213 -2331 1214 -2329
rect 1220 -2325 1221 -2323
rect 1220 -2331 1221 -2329
rect 1227 -2325 1228 -2323
rect 1227 -2331 1228 -2329
rect 1237 -2325 1238 -2323
rect 1234 -2331 1235 -2329
rect 1241 -2325 1242 -2323
rect 1241 -2331 1242 -2329
rect 1248 -2325 1249 -2323
rect 1248 -2331 1249 -2329
rect 1255 -2325 1256 -2323
rect 1255 -2331 1256 -2329
rect 1262 -2325 1263 -2323
rect 1262 -2331 1263 -2329
rect 1269 -2325 1270 -2323
rect 1269 -2331 1270 -2329
rect 1276 -2325 1277 -2323
rect 1276 -2331 1277 -2329
rect 1283 -2325 1284 -2323
rect 1283 -2331 1284 -2329
rect 1290 -2325 1291 -2323
rect 1290 -2331 1291 -2329
rect 1297 -2325 1298 -2323
rect 1297 -2331 1298 -2329
rect 1304 -2325 1305 -2323
rect 1304 -2331 1305 -2329
rect 1307 -2331 1308 -2329
rect 1311 -2325 1312 -2323
rect 1311 -2331 1312 -2329
rect 1318 -2325 1319 -2323
rect 1318 -2331 1319 -2329
rect 1325 -2325 1326 -2323
rect 1325 -2331 1326 -2329
rect 1332 -2325 1333 -2323
rect 1335 -2325 1336 -2323
rect 1332 -2331 1333 -2329
rect 1335 -2331 1336 -2329
rect 1339 -2325 1340 -2323
rect 1339 -2331 1340 -2329
rect 1346 -2325 1347 -2323
rect 1346 -2331 1347 -2329
rect 1353 -2325 1354 -2323
rect 1353 -2331 1354 -2329
rect 1360 -2325 1361 -2323
rect 1360 -2331 1361 -2329
rect 1367 -2325 1368 -2323
rect 1367 -2331 1368 -2329
rect 1374 -2325 1375 -2323
rect 1374 -2331 1375 -2329
rect 1381 -2325 1382 -2323
rect 1381 -2331 1382 -2329
rect 1388 -2325 1389 -2323
rect 1388 -2331 1389 -2329
rect 1395 -2325 1396 -2323
rect 1395 -2331 1396 -2329
rect 1402 -2325 1403 -2323
rect 1402 -2331 1403 -2329
rect 1409 -2325 1410 -2323
rect 1409 -2331 1410 -2329
rect 1416 -2325 1417 -2323
rect 1416 -2331 1417 -2329
rect 1423 -2325 1424 -2323
rect 1423 -2331 1424 -2329
rect 1430 -2325 1431 -2323
rect 1430 -2331 1431 -2329
rect 1437 -2325 1438 -2323
rect 1437 -2331 1438 -2329
rect 1444 -2325 1445 -2323
rect 1444 -2331 1445 -2329
rect 1451 -2325 1452 -2323
rect 1451 -2331 1452 -2329
rect 1458 -2325 1459 -2323
rect 1458 -2331 1459 -2329
rect 1465 -2325 1466 -2323
rect 1465 -2331 1466 -2329
rect 1472 -2325 1473 -2323
rect 1472 -2331 1473 -2329
rect 1479 -2325 1480 -2323
rect 1479 -2331 1480 -2329
rect 1486 -2325 1487 -2323
rect 1486 -2331 1487 -2329
rect 1493 -2325 1494 -2323
rect 1493 -2331 1494 -2329
rect 1500 -2325 1501 -2323
rect 1500 -2331 1501 -2329
rect 1507 -2325 1508 -2323
rect 1507 -2331 1508 -2329
rect 1514 -2325 1515 -2323
rect 1514 -2331 1515 -2329
rect 1521 -2325 1522 -2323
rect 1521 -2331 1522 -2329
rect 1528 -2325 1529 -2323
rect 1528 -2331 1529 -2329
rect 1535 -2325 1536 -2323
rect 1535 -2331 1536 -2329
rect 1542 -2325 1543 -2323
rect 1542 -2331 1543 -2329
rect 1549 -2325 1550 -2323
rect 1549 -2331 1550 -2329
rect 1556 -2325 1557 -2323
rect 1556 -2331 1557 -2329
rect 1563 -2325 1564 -2323
rect 1563 -2331 1564 -2329
rect 1570 -2325 1571 -2323
rect 1570 -2331 1571 -2329
rect 1577 -2325 1578 -2323
rect 1577 -2331 1578 -2329
rect 1584 -2325 1585 -2323
rect 1584 -2331 1585 -2329
rect 1591 -2325 1592 -2323
rect 1591 -2331 1592 -2329
rect 1598 -2325 1599 -2323
rect 1598 -2331 1599 -2329
rect 1605 -2325 1606 -2323
rect 1605 -2331 1606 -2329
rect 1612 -2325 1613 -2323
rect 1612 -2331 1613 -2329
rect 1619 -2325 1620 -2323
rect 1619 -2331 1620 -2329
rect 1626 -2325 1627 -2323
rect 1626 -2331 1627 -2329
rect 1633 -2325 1634 -2323
rect 1633 -2331 1634 -2329
rect 1640 -2325 1641 -2323
rect 1640 -2331 1641 -2329
rect 1647 -2325 1648 -2323
rect 1647 -2331 1648 -2329
rect 1654 -2325 1655 -2323
rect 1654 -2331 1655 -2329
rect 1661 -2325 1662 -2323
rect 1661 -2331 1662 -2329
rect 1668 -2325 1669 -2323
rect 1668 -2331 1669 -2329
rect 1675 -2325 1676 -2323
rect 1675 -2331 1676 -2329
rect 1682 -2325 1683 -2323
rect 1682 -2331 1683 -2329
rect 1689 -2325 1690 -2323
rect 1689 -2331 1690 -2329
rect 1696 -2325 1697 -2323
rect 1696 -2331 1697 -2329
rect 1703 -2325 1704 -2323
rect 1706 -2325 1707 -2323
rect 1703 -2331 1704 -2329
rect 1706 -2331 1707 -2329
rect 1710 -2325 1711 -2323
rect 1713 -2325 1714 -2323
rect 1710 -2331 1711 -2329
rect 1717 -2325 1718 -2323
rect 1717 -2331 1718 -2329
rect 1724 -2325 1725 -2323
rect 1724 -2331 1725 -2329
rect 1731 -2325 1732 -2323
rect 1731 -2331 1732 -2329
rect 1738 -2325 1739 -2323
rect 1738 -2331 1739 -2329
rect 51 -2440 52 -2438
rect 51 -2446 52 -2444
rect 58 -2440 59 -2438
rect 58 -2446 59 -2444
rect 65 -2440 66 -2438
rect 65 -2446 66 -2444
rect 72 -2440 73 -2438
rect 72 -2446 73 -2444
rect 79 -2440 80 -2438
rect 79 -2446 80 -2444
rect 86 -2440 87 -2438
rect 86 -2446 87 -2444
rect 93 -2440 94 -2438
rect 93 -2446 94 -2444
rect 100 -2440 101 -2438
rect 100 -2446 101 -2444
rect 107 -2440 108 -2438
rect 107 -2446 108 -2444
rect 114 -2440 115 -2438
rect 114 -2446 115 -2444
rect 121 -2440 122 -2438
rect 121 -2446 122 -2444
rect 128 -2440 129 -2438
rect 128 -2446 129 -2444
rect 135 -2440 136 -2438
rect 135 -2446 136 -2444
rect 142 -2440 143 -2438
rect 142 -2446 143 -2444
rect 149 -2440 150 -2438
rect 149 -2446 150 -2444
rect 156 -2440 157 -2438
rect 156 -2446 157 -2444
rect 163 -2440 164 -2438
rect 163 -2446 164 -2444
rect 170 -2440 171 -2438
rect 170 -2446 171 -2444
rect 177 -2440 178 -2438
rect 180 -2440 181 -2438
rect 180 -2446 181 -2444
rect 184 -2440 185 -2438
rect 184 -2446 185 -2444
rect 191 -2440 192 -2438
rect 191 -2446 192 -2444
rect 198 -2440 199 -2438
rect 198 -2446 199 -2444
rect 205 -2440 206 -2438
rect 205 -2446 206 -2444
rect 212 -2440 213 -2438
rect 215 -2440 216 -2438
rect 212 -2446 213 -2444
rect 215 -2446 216 -2444
rect 219 -2440 220 -2438
rect 219 -2446 220 -2444
rect 226 -2440 227 -2438
rect 226 -2446 227 -2444
rect 233 -2440 234 -2438
rect 233 -2446 234 -2444
rect 240 -2440 241 -2438
rect 240 -2446 241 -2444
rect 247 -2440 248 -2438
rect 247 -2446 248 -2444
rect 254 -2440 255 -2438
rect 257 -2446 258 -2444
rect 261 -2440 262 -2438
rect 261 -2446 262 -2444
rect 268 -2440 269 -2438
rect 268 -2446 269 -2444
rect 275 -2440 276 -2438
rect 275 -2446 276 -2444
rect 282 -2440 283 -2438
rect 282 -2446 283 -2444
rect 289 -2440 290 -2438
rect 289 -2446 290 -2444
rect 296 -2440 297 -2438
rect 296 -2446 297 -2444
rect 303 -2440 304 -2438
rect 303 -2446 304 -2444
rect 310 -2440 311 -2438
rect 313 -2446 314 -2444
rect 317 -2440 318 -2438
rect 317 -2446 318 -2444
rect 324 -2440 325 -2438
rect 324 -2446 325 -2444
rect 331 -2440 332 -2438
rect 331 -2446 332 -2444
rect 338 -2440 339 -2438
rect 338 -2446 339 -2444
rect 345 -2440 346 -2438
rect 345 -2446 346 -2444
rect 352 -2440 353 -2438
rect 352 -2446 353 -2444
rect 359 -2440 360 -2438
rect 359 -2446 360 -2444
rect 366 -2440 367 -2438
rect 366 -2446 367 -2444
rect 373 -2440 374 -2438
rect 373 -2446 374 -2444
rect 380 -2440 381 -2438
rect 380 -2446 381 -2444
rect 387 -2440 388 -2438
rect 387 -2446 388 -2444
rect 394 -2440 395 -2438
rect 394 -2446 395 -2444
rect 401 -2440 402 -2438
rect 401 -2446 402 -2444
rect 408 -2440 409 -2438
rect 408 -2446 409 -2444
rect 415 -2440 416 -2438
rect 415 -2446 416 -2444
rect 422 -2440 423 -2438
rect 422 -2446 423 -2444
rect 432 -2440 433 -2438
rect 429 -2446 430 -2444
rect 432 -2446 433 -2444
rect 436 -2440 437 -2438
rect 436 -2446 437 -2444
rect 443 -2440 444 -2438
rect 443 -2446 444 -2444
rect 450 -2440 451 -2438
rect 450 -2446 451 -2444
rect 457 -2440 458 -2438
rect 457 -2446 458 -2444
rect 464 -2440 465 -2438
rect 464 -2446 465 -2444
rect 471 -2440 472 -2438
rect 474 -2440 475 -2438
rect 474 -2446 475 -2444
rect 478 -2440 479 -2438
rect 478 -2446 479 -2444
rect 485 -2440 486 -2438
rect 485 -2446 486 -2444
rect 492 -2440 493 -2438
rect 492 -2446 493 -2444
rect 499 -2440 500 -2438
rect 502 -2440 503 -2438
rect 499 -2446 500 -2444
rect 502 -2446 503 -2444
rect 506 -2440 507 -2438
rect 506 -2446 507 -2444
rect 513 -2440 514 -2438
rect 513 -2446 514 -2444
rect 520 -2440 521 -2438
rect 520 -2446 521 -2444
rect 530 -2440 531 -2438
rect 527 -2446 528 -2444
rect 530 -2446 531 -2444
rect 534 -2440 535 -2438
rect 534 -2446 535 -2444
rect 541 -2440 542 -2438
rect 541 -2446 542 -2444
rect 548 -2440 549 -2438
rect 548 -2446 549 -2444
rect 555 -2440 556 -2438
rect 555 -2446 556 -2444
rect 562 -2440 563 -2438
rect 562 -2446 563 -2444
rect 569 -2440 570 -2438
rect 569 -2446 570 -2444
rect 576 -2440 577 -2438
rect 576 -2446 577 -2444
rect 583 -2440 584 -2438
rect 583 -2446 584 -2444
rect 590 -2440 591 -2438
rect 590 -2446 591 -2444
rect 597 -2440 598 -2438
rect 597 -2446 598 -2444
rect 604 -2440 605 -2438
rect 604 -2446 605 -2444
rect 611 -2440 612 -2438
rect 614 -2440 615 -2438
rect 611 -2446 612 -2444
rect 618 -2440 619 -2438
rect 618 -2446 619 -2444
rect 625 -2440 626 -2438
rect 625 -2446 626 -2444
rect 632 -2440 633 -2438
rect 632 -2446 633 -2444
rect 639 -2440 640 -2438
rect 642 -2446 643 -2444
rect 646 -2440 647 -2438
rect 646 -2446 647 -2444
rect 653 -2440 654 -2438
rect 653 -2446 654 -2444
rect 660 -2440 661 -2438
rect 660 -2446 661 -2444
rect 667 -2440 668 -2438
rect 667 -2446 668 -2444
rect 674 -2440 675 -2438
rect 677 -2440 678 -2438
rect 674 -2446 675 -2444
rect 677 -2446 678 -2444
rect 684 -2440 685 -2438
rect 681 -2446 682 -2444
rect 684 -2446 685 -2444
rect 688 -2440 689 -2438
rect 688 -2446 689 -2444
rect 695 -2440 696 -2438
rect 695 -2446 696 -2444
rect 705 -2440 706 -2438
rect 705 -2446 706 -2444
rect 709 -2440 710 -2438
rect 709 -2446 710 -2444
rect 716 -2440 717 -2438
rect 716 -2446 717 -2444
rect 723 -2440 724 -2438
rect 723 -2446 724 -2444
rect 730 -2440 731 -2438
rect 733 -2440 734 -2438
rect 730 -2446 731 -2444
rect 733 -2446 734 -2444
rect 737 -2440 738 -2438
rect 737 -2446 738 -2444
rect 744 -2440 745 -2438
rect 747 -2440 748 -2438
rect 747 -2446 748 -2444
rect 751 -2440 752 -2438
rect 751 -2446 752 -2444
rect 758 -2440 759 -2438
rect 758 -2446 759 -2444
rect 765 -2440 766 -2438
rect 765 -2446 766 -2444
rect 772 -2440 773 -2438
rect 772 -2446 773 -2444
rect 779 -2440 780 -2438
rect 779 -2446 780 -2444
rect 786 -2440 787 -2438
rect 786 -2446 787 -2444
rect 793 -2440 794 -2438
rect 793 -2446 794 -2444
rect 800 -2440 801 -2438
rect 800 -2446 801 -2444
rect 807 -2440 808 -2438
rect 810 -2440 811 -2438
rect 807 -2446 808 -2444
rect 810 -2446 811 -2444
rect 814 -2440 815 -2438
rect 814 -2446 815 -2444
rect 821 -2440 822 -2438
rect 824 -2440 825 -2438
rect 821 -2446 822 -2444
rect 824 -2446 825 -2444
rect 828 -2440 829 -2438
rect 828 -2446 829 -2444
rect 835 -2440 836 -2438
rect 835 -2446 836 -2444
rect 842 -2440 843 -2438
rect 845 -2440 846 -2438
rect 845 -2446 846 -2444
rect 849 -2440 850 -2438
rect 852 -2440 853 -2438
rect 849 -2446 850 -2444
rect 852 -2446 853 -2444
rect 856 -2440 857 -2438
rect 856 -2446 857 -2444
rect 859 -2446 860 -2444
rect 863 -2440 864 -2438
rect 863 -2446 864 -2444
rect 870 -2440 871 -2438
rect 870 -2446 871 -2444
rect 877 -2440 878 -2438
rect 877 -2446 878 -2444
rect 884 -2440 885 -2438
rect 884 -2446 885 -2444
rect 891 -2440 892 -2438
rect 891 -2446 892 -2444
rect 894 -2446 895 -2444
rect 898 -2440 899 -2438
rect 901 -2440 902 -2438
rect 898 -2446 899 -2444
rect 901 -2446 902 -2444
rect 905 -2440 906 -2438
rect 905 -2446 906 -2444
rect 912 -2440 913 -2438
rect 912 -2446 913 -2444
rect 919 -2440 920 -2438
rect 919 -2446 920 -2444
rect 926 -2440 927 -2438
rect 926 -2446 927 -2444
rect 933 -2440 934 -2438
rect 933 -2446 934 -2444
rect 940 -2440 941 -2438
rect 940 -2446 941 -2444
rect 947 -2440 948 -2438
rect 947 -2446 948 -2444
rect 954 -2440 955 -2438
rect 954 -2446 955 -2444
rect 961 -2440 962 -2438
rect 961 -2446 962 -2444
rect 968 -2440 969 -2438
rect 971 -2440 972 -2438
rect 968 -2446 969 -2444
rect 971 -2446 972 -2444
rect 975 -2440 976 -2438
rect 975 -2446 976 -2444
rect 982 -2440 983 -2438
rect 982 -2446 983 -2444
rect 989 -2440 990 -2438
rect 989 -2446 990 -2444
rect 996 -2440 997 -2438
rect 996 -2446 997 -2444
rect 1003 -2440 1004 -2438
rect 1003 -2446 1004 -2444
rect 1010 -2440 1011 -2438
rect 1010 -2446 1011 -2444
rect 1017 -2440 1018 -2438
rect 1017 -2446 1018 -2444
rect 1024 -2440 1025 -2438
rect 1024 -2446 1025 -2444
rect 1031 -2440 1032 -2438
rect 1031 -2446 1032 -2444
rect 1038 -2440 1039 -2438
rect 1038 -2446 1039 -2444
rect 1045 -2440 1046 -2438
rect 1045 -2446 1046 -2444
rect 1052 -2440 1053 -2438
rect 1052 -2446 1053 -2444
rect 1059 -2440 1060 -2438
rect 1059 -2446 1060 -2444
rect 1066 -2440 1067 -2438
rect 1066 -2446 1067 -2444
rect 1073 -2440 1074 -2438
rect 1076 -2440 1077 -2438
rect 1073 -2446 1074 -2444
rect 1076 -2446 1077 -2444
rect 1080 -2440 1081 -2438
rect 1080 -2446 1081 -2444
rect 1087 -2440 1088 -2438
rect 1087 -2446 1088 -2444
rect 1094 -2440 1095 -2438
rect 1094 -2446 1095 -2444
rect 1101 -2440 1102 -2438
rect 1101 -2446 1102 -2444
rect 1108 -2440 1109 -2438
rect 1108 -2446 1109 -2444
rect 1115 -2440 1116 -2438
rect 1115 -2446 1116 -2444
rect 1122 -2440 1123 -2438
rect 1122 -2446 1123 -2444
rect 1129 -2440 1130 -2438
rect 1129 -2446 1130 -2444
rect 1136 -2440 1137 -2438
rect 1136 -2446 1137 -2444
rect 1143 -2440 1144 -2438
rect 1143 -2446 1144 -2444
rect 1150 -2440 1151 -2438
rect 1150 -2446 1151 -2444
rect 1157 -2440 1158 -2438
rect 1157 -2446 1158 -2444
rect 1164 -2440 1165 -2438
rect 1164 -2446 1165 -2444
rect 1171 -2440 1172 -2438
rect 1171 -2446 1172 -2444
rect 1178 -2440 1179 -2438
rect 1178 -2446 1179 -2444
rect 1185 -2440 1186 -2438
rect 1185 -2446 1186 -2444
rect 1192 -2440 1193 -2438
rect 1195 -2440 1196 -2438
rect 1192 -2446 1193 -2444
rect 1195 -2446 1196 -2444
rect 1199 -2440 1200 -2438
rect 1199 -2446 1200 -2444
rect 1206 -2440 1207 -2438
rect 1206 -2446 1207 -2444
rect 1209 -2446 1210 -2444
rect 1213 -2440 1214 -2438
rect 1213 -2446 1214 -2444
rect 1220 -2440 1221 -2438
rect 1220 -2446 1221 -2444
rect 1227 -2440 1228 -2438
rect 1227 -2446 1228 -2444
rect 1234 -2440 1235 -2438
rect 1234 -2446 1235 -2444
rect 1241 -2440 1242 -2438
rect 1244 -2440 1245 -2438
rect 1244 -2446 1245 -2444
rect 1248 -2440 1249 -2438
rect 1248 -2446 1249 -2444
rect 1255 -2440 1256 -2438
rect 1255 -2446 1256 -2444
rect 1262 -2440 1263 -2438
rect 1262 -2446 1263 -2444
rect 1269 -2440 1270 -2438
rect 1269 -2446 1270 -2444
rect 1276 -2440 1277 -2438
rect 1276 -2446 1277 -2444
rect 1283 -2440 1284 -2438
rect 1283 -2446 1284 -2444
rect 1290 -2440 1291 -2438
rect 1290 -2446 1291 -2444
rect 1297 -2446 1298 -2444
rect 1300 -2446 1301 -2444
rect 1304 -2440 1305 -2438
rect 1304 -2446 1305 -2444
rect 1314 -2440 1315 -2438
rect 1311 -2446 1312 -2444
rect 1314 -2446 1315 -2444
rect 1318 -2440 1319 -2438
rect 1318 -2446 1319 -2444
rect 1325 -2440 1326 -2438
rect 1325 -2446 1326 -2444
rect 1332 -2440 1333 -2438
rect 1332 -2446 1333 -2444
rect 1339 -2440 1340 -2438
rect 1339 -2446 1340 -2444
rect 1346 -2440 1347 -2438
rect 1346 -2446 1347 -2444
rect 1353 -2440 1354 -2438
rect 1353 -2446 1354 -2444
rect 1360 -2440 1361 -2438
rect 1360 -2446 1361 -2444
rect 1367 -2440 1368 -2438
rect 1367 -2446 1368 -2444
rect 1374 -2440 1375 -2438
rect 1374 -2446 1375 -2444
rect 1381 -2440 1382 -2438
rect 1384 -2440 1385 -2438
rect 1381 -2446 1382 -2444
rect 1388 -2440 1389 -2438
rect 1388 -2446 1389 -2444
rect 1395 -2440 1396 -2438
rect 1395 -2446 1396 -2444
rect 1402 -2440 1403 -2438
rect 1402 -2446 1403 -2444
rect 1409 -2440 1410 -2438
rect 1409 -2446 1410 -2444
rect 1416 -2440 1417 -2438
rect 1416 -2446 1417 -2444
rect 1423 -2440 1424 -2438
rect 1423 -2446 1424 -2444
rect 1430 -2440 1431 -2438
rect 1430 -2446 1431 -2444
rect 1437 -2440 1438 -2438
rect 1437 -2446 1438 -2444
rect 1444 -2440 1445 -2438
rect 1444 -2446 1445 -2444
rect 1451 -2440 1452 -2438
rect 1451 -2446 1452 -2444
rect 1458 -2440 1459 -2438
rect 1458 -2446 1459 -2444
rect 1465 -2440 1466 -2438
rect 1465 -2446 1466 -2444
rect 1472 -2440 1473 -2438
rect 1472 -2446 1473 -2444
rect 1479 -2440 1480 -2438
rect 1479 -2446 1480 -2444
rect 1486 -2440 1487 -2438
rect 1486 -2446 1487 -2444
rect 1493 -2440 1494 -2438
rect 1493 -2446 1494 -2444
rect 1500 -2440 1501 -2438
rect 1500 -2446 1501 -2444
rect 1507 -2440 1508 -2438
rect 1507 -2446 1508 -2444
rect 1514 -2440 1515 -2438
rect 1514 -2446 1515 -2444
rect 1521 -2440 1522 -2438
rect 1521 -2446 1522 -2444
rect 1528 -2440 1529 -2438
rect 1528 -2446 1529 -2444
rect 1538 -2440 1539 -2438
rect 1535 -2446 1536 -2444
rect 1538 -2446 1539 -2444
rect 1542 -2440 1543 -2438
rect 1542 -2446 1543 -2444
rect 1549 -2440 1550 -2438
rect 1549 -2446 1550 -2444
rect 1556 -2440 1557 -2438
rect 1556 -2446 1557 -2444
rect 1563 -2440 1564 -2438
rect 1563 -2446 1564 -2444
rect 1570 -2440 1571 -2438
rect 1570 -2446 1571 -2444
rect 1577 -2440 1578 -2438
rect 1577 -2446 1578 -2444
rect 1580 -2446 1581 -2444
rect 1584 -2440 1585 -2438
rect 1584 -2446 1585 -2444
rect 1591 -2440 1592 -2438
rect 1591 -2446 1592 -2444
rect 1598 -2440 1599 -2438
rect 1598 -2446 1599 -2444
rect 1605 -2440 1606 -2438
rect 1605 -2446 1606 -2444
rect 1675 -2440 1676 -2438
rect 1675 -2446 1676 -2444
rect 44 -2557 45 -2555
rect 44 -2563 45 -2561
rect 51 -2557 52 -2555
rect 51 -2563 52 -2561
rect 58 -2557 59 -2555
rect 58 -2563 59 -2561
rect 65 -2557 66 -2555
rect 68 -2557 69 -2555
rect 75 -2557 76 -2555
rect 72 -2563 73 -2561
rect 75 -2563 76 -2561
rect 79 -2557 80 -2555
rect 79 -2563 80 -2561
rect 86 -2557 87 -2555
rect 86 -2563 87 -2561
rect 93 -2557 94 -2555
rect 93 -2563 94 -2561
rect 100 -2557 101 -2555
rect 103 -2557 104 -2555
rect 100 -2563 101 -2561
rect 107 -2557 108 -2555
rect 107 -2563 108 -2561
rect 114 -2557 115 -2555
rect 114 -2563 115 -2561
rect 121 -2557 122 -2555
rect 121 -2563 122 -2561
rect 128 -2557 129 -2555
rect 128 -2563 129 -2561
rect 135 -2557 136 -2555
rect 135 -2563 136 -2561
rect 142 -2557 143 -2555
rect 142 -2563 143 -2561
rect 149 -2557 150 -2555
rect 152 -2557 153 -2555
rect 149 -2563 150 -2561
rect 152 -2563 153 -2561
rect 156 -2557 157 -2555
rect 156 -2563 157 -2561
rect 163 -2557 164 -2555
rect 166 -2557 167 -2555
rect 163 -2563 164 -2561
rect 166 -2563 167 -2561
rect 173 -2557 174 -2555
rect 170 -2563 171 -2561
rect 177 -2557 178 -2555
rect 177 -2563 178 -2561
rect 184 -2557 185 -2555
rect 184 -2563 185 -2561
rect 191 -2557 192 -2555
rect 191 -2563 192 -2561
rect 198 -2557 199 -2555
rect 198 -2563 199 -2561
rect 205 -2557 206 -2555
rect 205 -2563 206 -2561
rect 212 -2557 213 -2555
rect 212 -2563 213 -2561
rect 219 -2557 220 -2555
rect 219 -2563 220 -2561
rect 226 -2557 227 -2555
rect 226 -2563 227 -2561
rect 233 -2557 234 -2555
rect 233 -2563 234 -2561
rect 240 -2557 241 -2555
rect 240 -2563 241 -2561
rect 247 -2557 248 -2555
rect 247 -2563 248 -2561
rect 254 -2563 255 -2561
rect 257 -2563 258 -2561
rect 261 -2557 262 -2555
rect 261 -2563 262 -2561
rect 268 -2557 269 -2555
rect 268 -2563 269 -2561
rect 275 -2557 276 -2555
rect 275 -2563 276 -2561
rect 282 -2557 283 -2555
rect 282 -2563 283 -2561
rect 289 -2557 290 -2555
rect 289 -2563 290 -2561
rect 296 -2557 297 -2555
rect 296 -2563 297 -2561
rect 303 -2557 304 -2555
rect 303 -2563 304 -2561
rect 310 -2557 311 -2555
rect 310 -2563 311 -2561
rect 317 -2557 318 -2555
rect 317 -2563 318 -2561
rect 324 -2557 325 -2555
rect 324 -2563 325 -2561
rect 331 -2557 332 -2555
rect 331 -2563 332 -2561
rect 338 -2557 339 -2555
rect 338 -2563 339 -2561
rect 345 -2557 346 -2555
rect 345 -2563 346 -2561
rect 352 -2557 353 -2555
rect 352 -2563 353 -2561
rect 359 -2557 360 -2555
rect 359 -2563 360 -2561
rect 366 -2557 367 -2555
rect 366 -2563 367 -2561
rect 373 -2557 374 -2555
rect 373 -2563 374 -2561
rect 380 -2557 381 -2555
rect 380 -2563 381 -2561
rect 387 -2557 388 -2555
rect 387 -2563 388 -2561
rect 394 -2557 395 -2555
rect 394 -2563 395 -2561
rect 401 -2557 402 -2555
rect 401 -2563 402 -2561
rect 408 -2557 409 -2555
rect 411 -2557 412 -2555
rect 408 -2563 409 -2561
rect 415 -2557 416 -2555
rect 415 -2563 416 -2561
rect 422 -2557 423 -2555
rect 422 -2563 423 -2561
rect 432 -2557 433 -2555
rect 429 -2563 430 -2561
rect 432 -2563 433 -2561
rect 436 -2557 437 -2555
rect 436 -2563 437 -2561
rect 443 -2557 444 -2555
rect 446 -2557 447 -2555
rect 443 -2563 444 -2561
rect 446 -2563 447 -2561
rect 450 -2557 451 -2555
rect 450 -2563 451 -2561
rect 457 -2557 458 -2555
rect 457 -2563 458 -2561
rect 464 -2557 465 -2555
rect 464 -2563 465 -2561
rect 471 -2557 472 -2555
rect 471 -2563 472 -2561
rect 478 -2557 479 -2555
rect 478 -2563 479 -2561
rect 485 -2557 486 -2555
rect 485 -2563 486 -2561
rect 492 -2557 493 -2555
rect 492 -2563 493 -2561
rect 499 -2557 500 -2555
rect 499 -2563 500 -2561
rect 506 -2557 507 -2555
rect 506 -2563 507 -2561
rect 513 -2557 514 -2555
rect 513 -2563 514 -2561
rect 520 -2557 521 -2555
rect 520 -2563 521 -2561
rect 527 -2557 528 -2555
rect 527 -2563 528 -2561
rect 534 -2557 535 -2555
rect 534 -2563 535 -2561
rect 541 -2557 542 -2555
rect 541 -2563 542 -2561
rect 548 -2557 549 -2555
rect 551 -2557 552 -2555
rect 548 -2563 549 -2561
rect 551 -2563 552 -2561
rect 555 -2557 556 -2555
rect 555 -2563 556 -2561
rect 562 -2557 563 -2555
rect 562 -2563 563 -2561
rect 569 -2557 570 -2555
rect 569 -2563 570 -2561
rect 576 -2557 577 -2555
rect 576 -2563 577 -2561
rect 583 -2557 584 -2555
rect 583 -2563 584 -2561
rect 590 -2557 591 -2555
rect 593 -2557 594 -2555
rect 590 -2563 591 -2561
rect 593 -2563 594 -2561
rect 597 -2557 598 -2555
rect 597 -2563 598 -2561
rect 604 -2557 605 -2555
rect 604 -2563 605 -2561
rect 611 -2557 612 -2555
rect 611 -2563 612 -2561
rect 618 -2557 619 -2555
rect 618 -2563 619 -2561
rect 625 -2557 626 -2555
rect 628 -2557 629 -2555
rect 625 -2563 626 -2561
rect 632 -2557 633 -2555
rect 632 -2563 633 -2561
rect 639 -2557 640 -2555
rect 639 -2563 640 -2561
rect 646 -2557 647 -2555
rect 649 -2557 650 -2555
rect 646 -2563 647 -2561
rect 649 -2563 650 -2561
rect 653 -2557 654 -2555
rect 653 -2563 654 -2561
rect 660 -2557 661 -2555
rect 663 -2557 664 -2555
rect 660 -2563 661 -2561
rect 663 -2563 664 -2561
rect 667 -2557 668 -2555
rect 667 -2563 668 -2561
rect 674 -2557 675 -2555
rect 674 -2563 675 -2561
rect 681 -2557 682 -2555
rect 681 -2563 682 -2561
rect 688 -2557 689 -2555
rect 688 -2563 689 -2561
rect 695 -2557 696 -2555
rect 695 -2563 696 -2561
rect 702 -2557 703 -2555
rect 702 -2563 703 -2561
rect 709 -2557 710 -2555
rect 709 -2563 710 -2561
rect 716 -2557 717 -2555
rect 716 -2563 717 -2561
rect 723 -2557 724 -2555
rect 723 -2563 724 -2561
rect 730 -2557 731 -2555
rect 733 -2557 734 -2555
rect 730 -2563 731 -2561
rect 733 -2563 734 -2561
rect 737 -2557 738 -2555
rect 740 -2557 741 -2555
rect 737 -2563 738 -2561
rect 740 -2563 741 -2561
rect 744 -2557 745 -2555
rect 747 -2557 748 -2555
rect 747 -2563 748 -2561
rect 751 -2557 752 -2555
rect 754 -2557 755 -2555
rect 751 -2563 752 -2561
rect 754 -2563 755 -2561
rect 758 -2557 759 -2555
rect 758 -2563 759 -2561
rect 765 -2557 766 -2555
rect 765 -2563 766 -2561
rect 772 -2557 773 -2555
rect 772 -2563 773 -2561
rect 779 -2557 780 -2555
rect 779 -2563 780 -2561
rect 786 -2557 787 -2555
rect 789 -2557 790 -2555
rect 786 -2563 787 -2561
rect 789 -2563 790 -2561
rect 793 -2557 794 -2555
rect 793 -2563 794 -2561
rect 800 -2557 801 -2555
rect 800 -2563 801 -2561
rect 807 -2557 808 -2555
rect 807 -2563 808 -2561
rect 814 -2557 815 -2555
rect 814 -2563 815 -2561
rect 821 -2557 822 -2555
rect 824 -2557 825 -2555
rect 821 -2563 822 -2561
rect 824 -2563 825 -2561
rect 828 -2557 829 -2555
rect 828 -2563 829 -2561
rect 835 -2557 836 -2555
rect 835 -2563 836 -2561
rect 842 -2557 843 -2555
rect 842 -2563 843 -2561
rect 849 -2557 850 -2555
rect 849 -2563 850 -2561
rect 856 -2557 857 -2555
rect 856 -2563 857 -2561
rect 863 -2557 864 -2555
rect 863 -2563 864 -2561
rect 870 -2557 871 -2555
rect 873 -2557 874 -2555
rect 870 -2563 871 -2561
rect 873 -2563 874 -2561
rect 877 -2557 878 -2555
rect 877 -2563 878 -2561
rect 884 -2557 885 -2555
rect 884 -2563 885 -2561
rect 891 -2557 892 -2555
rect 891 -2563 892 -2561
rect 898 -2557 899 -2555
rect 898 -2563 899 -2561
rect 905 -2557 906 -2555
rect 905 -2563 906 -2561
rect 912 -2557 913 -2555
rect 912 -2563 913 -2561
rect 919 -2557 920 -2555
rect 919 -2563 920 -2561
rect 926 -2557 927 -2555
rect 929 -2557 930 -2555
rect 926 -2563 927 -2561
rect 929 -2563 930 -2561
rect 933 -2557 934 -2555
rect 933 -2563 934 -2561
rect 940 -2557 941 -2555
rect 940 -2563 941 -2561
rect 947 -2557 948 -2555
rect 947 -2563 948 -2561
rect 954 -2557 955 -2555
rect 957 -2557 958 -2555
rect 954 -2563 955 -2561
rect 957 -2563 958 -2561
rect 961 -2557 962 -2555
rect 961 -2563 962 -2561
rect 968 -2557 969 -2555
rect 968 -2563 969 -2561
rect 975 -2557 976 -2555
rect 975 -2563 976 -2561
rect 982 -2557 983 -2555
rect 982 -2563 983 -2561
rect 989 -2557 990 -2555
rect 989 -2563 990 -2561
rect 996 -2557 997 -2555
rect 996 -2563 997 -2561
rect 1003 -2557 1004 -2555
rect 1003 -2563 1004 -2561
rect 1010 -2557 1011 -2555
rect 1010 -2563 1011 -2561
rect 1017 -2557 1018 -2555
rect 1017 -2563 1018 -2561
rect 1024 -2557 1025 -2555
rect 1024 -2563 1025 -2561
rect 1031 -2557 1032 -2555
rect 1031 -2563 1032 -2561
rect 1038 -2557 1039 -2555
rect 1038 -2563 1039 -2561
rect 1045 -2557 1046 -2555
rect 1045 -2563 1046 -2561
rect 1052 -2557 1053 -2555
rect 1052 -2563 1053 -2561
rect 1059 -2557 1060 -2555
rect 1062 -2557 1063 -2555
rect 1059 -2563 1060 -2561
rect 1062 -2563 1063 -2561
rect 1066 -2557 1067 -2555
rect 1066 -2563 1067 -2561
rect 1073 -2557 1074 -2555
rect 1073 -2563 1074 -2561
rect 1080 -2557 1081 -2555
rect 1083 -2557 1084 -2555
rect 1083 -2563 1084 -2561
rect 1087 -2557 1088 -2555
rect 1090 -2557 1091 -2555
rect 1090 -2563 1091 -2561
rect 1094 -2557 1095 -2555
rect 1094 -2563 1095 -2561
rect 1101 -2557 1102 -2555
rect 1101 -2563 1102 -2561
rect 1108 -2557 1109 -2555
rect 1108 -2563 1109 -2561
rect 1115 -2557 1116 -2555
rect 1115 -2563 1116 -2561
rect 1122 -2557 1123 -2555
rect 1122 -2563 1123 -2561
rect 1129 -2557 1130 -2555
rect 1129 -2563 1130 -2561
rect 1136 -2557 1137 -2555
rect 1136 -2563 1137 -2561
rect 1143 -2557 1144 -2555
rect 1143 -2563 1144 -2561
rect 1150 -2557 1151 -2555
rect 1150 -2563 1151 -2561
rect 1157 -2557 1158 -2555
rect 1157 -2563 1158 -2561
rect 1164 -2557 1165 -2555
rect 1167 -2557 1168 -2555
rect 1164 -2563 1165 -2561
rect 1167 -2563 1168 -2561
rect 1171 -2557 1172 -2555
rect 1171 -2563 1172 -2561
rect 1178 -2557 1179 -2555
rect 1178 -2563 1179 -2561
rect 1185 -2557 1186 -2555
rect 1188 -2557 1189 -2555
rect 1185 -2563 1186 -2561
rect 1192 -2557 1193 -2555
rect 1192 -2563 1193 -2561
rect 1199 -2557 1200 -2555
rect 1199 -2563 1200 -2561
rect 1206 -2557 1207 -2555
rect 1206 -2563 1207 -2561
rect 1213 -2557 1214 -2555
rect 1213 -2563 1214 -2561
rect 1220 -2557 1221 -2555
rect 1220 -2563 1221 -2561
rect 1227 -2557 1228 -2555
rect 1227 -2563 1228 -2561
rect 1234 -2557 1235 -2555
rect 1234 -2563 1235 -2561
rect 1241 -2557 1242 -2555
rect 1241 -2563 1242 -2561
rect 1248 -2557 1249 -2555
rect 1248 -2563 1249 -2561
rect 1255 -2557 1256 -2555
rect 1255 -2563 1256 -2561
rect 1262 -2557 1263 -2555
rect 1262 -2563 1263 -2561
rect 1269 -2557 1270 -2555
rect 1269 -2563 1270 -2561
rect 1276 -2557 1277 -2555
rect 1276 -2563 1277 -2561
rect 1283 -2557 1284 -2555
rect 1283 -2563 1284 -2561
rect 1290 -2557 1291 -2555
rect 1290 -2563 1291 -2561
rect 1297 -2557 1298 -2555
rect 1297 -2563 1298 -2561
rect 1304 -2557 1305 -2555
rect 1304 -2563 1305 -2561
rect 1311 -2557 1312 -2555
rect 1311 -2563 1312 -2561
rect 1318 -2557 1319 -2555
rect 1318 -2563 1319 -2561
rect 1325 -2557 1326 -2555
rect 1325 -2563 1326 -2561
rect 1332 -2557 1333 -2555
rect 1332 -2563 1333 -2561
rect 1339 -2557 1340 -2555
rect 1339 -2563 1340 -2561
rect 1346 -2557 1347 -2555
rect 1346 -2563 1347 -2561
rect 1353 -2557 1354 -2555
rect 1353 -2563 1354 -2561
rect 1360 -2557 1361 -2555
rect 1360 -2563 1361 -2561
rect 1367 -2557 1368 -2555
rect 1367 -2563 1368 -2561
rect 1374 -2557 1375 -2555
rect 1374 -2563 1375 -2561
rect 1381 -2557 1382 -2555
rect 1381 -2563 1382 -2561
rect 1388 -2557 1389 -2555
rect 1388 -2563 1389 -2561
rect 1395 -2557 1396 -2555
rect 1395 -2563 1396 -2561
rect 1402 -2557 1403 -2555
rect 1402 -2563 1403 -2561
rect 1409 -2557 1410 -2555
rect 1409 -2563 1410 -2561
rect 1416 -2557 1417 -2555
rect 1416 -2563 1417 -2561
rect 1423 -2557 1424 -2555
rect 1423 -2563 1424 -2561
rect 1430 -2557 1431 -2555
rect 1430 -2563 1431 -2561
rect 1437 -2557 1438 -2555
rect 1437 -2563 1438 -2561
rect 1444 -2557 1445 -2555
rect 1444 -2563 1445 -2561
rect 1451 -2557 1452 -2555
rect 1451 -2563 1452 -2561
rect 1458 -2557 1459 -2555
rect 1458 -2563 1459 -2561
rect 1465 -2557 1466 -2555
rect 1465 -2563 1466 -2561
rect 1472 -2557 1473 -2555
rect 1472 -2563 1473 -2561
rect 1479 -2557 1480 -2555
rect 1479 -2563 1480 -2561
rect 1486 -2557 1487 -2555
rect 1486 -2563 1487 -2561
rect 1493 -2557 1494 -2555
rect 1493 -2563 1494 -2561
rect 1500 -2557 1501 -2555
rect 1500 -2563 1501 -2561
rect 1507 -2557 1508 -2555
rect 1507 -2563 1508 -2561
rect 1514 -2557 1515 -2555
rect 1514 -2563 1515 -2561
rect 1521 -2557 1522 -2555
rect 1521 -2563 1522 -2561
rect 1528 -2557 1529 -2555
rect 1528 -2563 1529 -2561
rect 1535 -2557 1536 -2555
rect 1535 -2563 1536 -2561
rect 1542 -2557 1543 -2555
rect 1542 -2563 1543 -2561
rect 1549 -2557 1550 -2555
rect 1549 -2563 1550 -2561
rect 1556 -2557 1557 -2555
rect 1556 -2563 1557 -2561
rect 1563 -2557 1564 -2555
rect 1563 -2563 1564 -2561
rect 1570 -2557 1571 -2555
rect 1570 -2563 1571 -2561
rect 1577 -2557 1578 -2555
rect 1577 -2563 1578 -2561
rect 1584 -2557 1585 -2555
rect 1584 -2563 1585 -2561
rect 1591 -2557 1592 -2555
rect 1591 -2563 1592 -2561
rect 1598 -2557 1599 -2555
rect 1598 -2563 1599 -2561
rect 1605 -2557 1606 -2555
rect 1605 -2563 1606 -2561
rect 1612 -2557 1613 -2555
rect 1612 -2563 1613 -2561
rect 1619 -2557 1620 -2555
rect 1619 -2563 1620 -2561
rect 1626 -2557 1627 -2555
rect 1626 -2563 1627 -2561
rect 1633 -2557 1634 -2555
rect 1633 -2563 1634 -2561
rect 1640 -2557 1641 -2555
rect 1640 -2563 1641 -2561
rect 1647 -2557 1648 -2555
rect 1647 -2563 1648 -2561
rect 1654 -2557 1655 -2555
rect 1654 -2563 1655 -2561
rect 1661 -2557 1662 -2555
rect 1661 -2563 1662 -2561
rect 1668 -2557 1669 -2555
rect 1668 -2563 1669 -2561
rect 1678 -2557 1679 -2555
rect 1675 -2563 1676 -2561
rect 1678 -2563 1679 -2561
rect 1682 -2557 1683 -2555
rect 1682 -2563 1683 -2561
rect 1689 -2557 1690 -2555
rect 1689 -2563 1690 -2561
rect 1696 -2557 1697 -2555
rect 1696 -2563 1697 -2561
rect 1706 -2557 1707 -2555
rect 1703 -2563 1704 -2561
rect 1710 -2557 1711 -2555
rect 1710 -2563 1711 -2561
rect 1717 -2557 1718 -2555
rect 1717 -2563 1718 -2561
rect 1724 -2557 1725 -2555
rect 1724 -2563 1725 -2561
rect 1731 -2557 1732 -2555
rect 1731 -2563 1732 -2561
rect 1738 -2557 1739 -2555
rect 1738 -2563 1739 -2561
rect 44 -2686 45 -2684
rect 44 -2692 45 -2690
rect 51 -2686 52 -2684
rect 51 -2692 52 -2690
rect 58 -2686 59 -2684
rect 58 -2692 59 -2690
rect 65 -2686 66 -2684
rect 68 -2686 69 -2684
rect 65 -2692 66 -2690
rect 68 -2692 69 -2690
rect 72 -2686 73 -2684
rect 72 -2692 73 -2690
rect 82 -2686 83 -2684
rect 79 -2692 80 -2690
rect 82 -2692 83 -2690
rect 86 -2686 87 -2684
rect 89 -2686 90 -2684
rect 86 -2692 87 -2690
rect 89 -2692 90 -2690
rect 93 -2686 94 -2684
rect 93 -2692 94 -2690
rect 100 -2686 101 -2684
rect 100 -2692 101 -2690
rect 107 -2686 108 -2684
rect 107 -2692 108 -2690
rect 117 -2686 118 -2684
rect 114 -2692 115 -2690
rect 117 -2692 118 -2690
rect 121 -2686 122 -2684
rect 121 -2692 122 -2690
rect 128 -2686 129 -2684
rect 128 -2692 129 -2690
rect 135 -2686 136 -2684
rect 135 -2692 136 -2690
rect 142 -2686 143 -2684
rect 142 -2692 143 -2690
rect 149 -2686 150 -2684
rect 149 -2692 150 -2690
rect 156 -2686 157 -2684
rect 156 -2692 157 -2690
rect 163 -2686 164 -2684
rect 166 -2686 167 -2684
rect 163 -2692 164 -2690
rect 166 -2692 167 -2690
rect 170 -2686 171 -2684
rect 170 -2692 171 -2690
rect 177 -2686 178 -2684
rect 177 -2692 178 -2690
rect 184 -2686 185 -2684
rect 184 -2692 185 -2690
rect 191 -2686 192 -2684
rect 201 -2686 202 -2684
rect 198 -2692 199 -2690
rect 201 -2692 202 -2690
rect 205 -2686 206 -2684
rect 205 -2692 206 -2690
rect 212 -2686 213 -2684
rect 212 -2692 213 -2690
rect 219 -2686 220 -2684
rect 219 -2692 220 -2690
rect 226 -2686 227 -2684
rect 226 -2692 227 -2690
rect 233 -2686 234 -2684
rect 233 -2692 234 -2690
rect 240 -2686 241 -2684
rect 240 -2692 241 -2690
rect 247 -2692 248 -2690
rect 250 -2692 251 -2690
rect 254 -2686 255 -2684
rect 254 -2692 255 -2690
rect 261 -2686 262 -2684
rect 261 -2692 262 -2690
rect 268 -2686 269 -2684
rect 268 -2692 269 -2690
rect 275 -2686 276 -2684
rect 275 -2692 276 -2690
rect 278 -2692 279 -2690
rect 282 -2686 283 -2684
rect 282 -2692 283 -2690
rect 289 -2686 290 -2684
rect 289 -2692 290 -2690
rect 296 -2686 297 -2684
rect 296 -2692 297 -2690
rect 303 -2686 304 -2684
rect 303 -2692 304 -2690
rect 310 -2686 311 -2684
rect 310 -2692 311 -2690
rect 317 -2686 318 -2684
rect 317 -2692 318 -2690
rect 324 -2686 325 -2684
rect 324 -2692 325 -2690
rect 331 -2686 332 -2684
rect 331 -2692 332 -2690
rect 338 -2686 339 -2684
rect 338 -2692 339 -2690
rect 345 -2686 346 -2684
rect 345 -2692 346 -2690
rect 352 -2686 353 -2684
rect 352 -2692 353 -2690
rect 359 -2686 360 -2684
rect 359 -2692 360 -2690
rect 366 -2686 367 -2684
rect 366 -2692 367 -2690
rect 373 -2686 374 -2684
rect 373 -2692 374 -2690
rect 380 -2686 381 -2684
rect 380 -2692 381 -2690
rect 387 -2686 388 -2684
rect 387 -2692 388 -2690
rect 394 -2686 395 -2684
rect 394 -2692 395 -2690
rect 401 -2686 402 -2684
rect 401 -2692 402 -2690
rect 408 -2686 409 -2684
rect 411 -2686 412 -2684
rect 411 -2692 412 -2690
rect 418 -2686 419 -2684
rect 415 -2692 416 -2690
rect 418 -2692 419 -2690
rect 422 -2686 423 -2684
rect 422 -2692 423 -2690
rect 429 -2686 430 -2684
rect 429 -2692 430 -2690
rect 436 -2686 437 -2684
rect 436 -2692 437 -2690
rect 443 -2686 444 -2684
rect 443 -2692 444 -2690
rect 450 -2686 451 -2684
rect 450 -2692 451 -2690
rect 453 -2692 454 -2690
rect 457 -2686 458 -2684
rect 460 -2686 461 -2684
rect 457 -2692 458 -2690
rect 464 -2686 465 -2684
rect 464 -2692 465 -2690
rect 467 -2692 468 -2690
rect 471 -2686 472 -2684
rect 471 -2692 472 -2690
rect 478 -2686 479 -2684
rect 481 -2692 482 -2690
rect 485 -2686 486 -2684
rect 485 -2692 486 -2690
rect 492 -2686 493 -2684
rect 492 -2692 493 -2690
rect 499 -2686 500 -2684
rect 499 -2692 500 -2690
rect 506 -2686 507 -2684
rect 506 -2692 507 -2690
rect 513 -2686 514 -2684
rect 513 -2692 514 -2690
rect 520 -2686 521 -2684
rect 520 -2692 521 -2690
rect 527 -2686 528 -2684
rect 527 -2692 528 -2690
rect 534 -2686 535 -2684
rect 534 -2692 535 -2690
rect 541 -2686 542 -2684
rect 541 -2692 542 -2690
rect 548 -2686 549 -2684
rect 548 -2692 549 -2690
rect 555 -2686 556 -2684
rect 555 -2692 556 -2690
rect 562 -2686 563 -2684
rect 562 -2692 563 -2690
rect 569 -2686 570 -2684
rect 569 -2692 570 -2690
rect 576 -2686 577 -2684
rect 579 -2692 580 -2690
rect 583 -2686 584 -2684
rect 583 -2692 584 -2690
rect 590 -2686 591 -2684
rect 590 -2692 591 -2690
rect 597 -2686 598 -2684
rect 600 -2686 601 -2684
rect 597 -2692 598 -2690
rect 600 -2692 601 -2690
rect 604 -2686 605 -2684
rect 604 -2692 605 -2690
rect 611 -2686 612 -2684
rect 611 -2692 612 -2690
rect 618 -2686 619 -2684
rect 618 -2692 619 -2690
rect 625 -2686 626 -2684
rect 628 -2686 629 -2684
rect 625 -2692 626 -2690
rect 628 -2692 629 -2690
rect 632 -2686 633 -2684
rect 632 -2692 633 -2690
rect 639 -2686 640 -2684
rect 639 -2692 640 -2690
rect 646 -2686 647 -2684
rect 646 -2692 647 -2690
rect 653 -2686 654 -2684
rect 653 -2692 654 -2690
rect 660 -2686 661 -2684
rect 660 -2692 661 -2690
rect 667 -2686 668 -2684
rect 670 -2686 671 -2684
rect 667 -2692 668 -2690
rect 670 -2692 671 -2690
rect 674 -2686 675 -2684
rect 677 -2686 678 -2684
rect 674 -2692 675 -2690
rect 677 -2692 678 -2690
rect 681 -2686 682 -2684
rect 681 -2692 682 -2690
rect 688 -2686 689 -2684
rect 691 -2686 692 -2684
rect 688 -2692 689 -2690
rect 695 -2686 696 -2684
rect 695 -2692 696 -2690
rect 702 -2686 703 -2684
rect 702 -2692 703 -2690
rect 709 -2686 710 -2684
rect 709 -2692 710 -2690
rect 716 -2686 717 -2684
rect 716 -2692 717 -2690
rect 723 -2686 724 -2684
rect 723 -2692 724 -2690
rect 733 -2686 734 -2684
rect 730 -2692 731 -2690
rect 733 -2692 734 -2690
rect 737 -2686 738 -2684
rect 737 -2692 738 -2690
rect 744 -2686 745 -2684
rect 744 -2692 745 -2690
rect 751 -2686 752 -2684
rect 751 -2692 752 -2690
rect 754 -2692 755 -2690
rect 758 -2686 759 -2684
rect 758 -2692 759 -2690
rect 765 -2686 766 -2684
rect 768 -2686 769 -2684
rect 765 -2692 766 -2690
rect 768 -2692 769 -2690
rect 772 -2686 773 -2684
rect 772 -2692 773 -2690
rect 779 -2686 780 -2684
rect 779 -2692 780 -2690
rect 786 -2686 787 -2684
rect 786 -2692 787 -2690
rect 793 -2686 794 -2684
rect 793 -2692 794 -2690
rect 800 -2686 801 -2684
rect 803 -2686 804 -2684
rect 800 -2692 801 -2690
rect 803 -2692 804 -2690
rect 807 -2686 808 -2684
rect 807 -2692 808 -2690
rect 814 -2686 815 -2684
rect 814 -2692 815 -2690
rect 821 -2686 822 -2684
rect 821 -2692 822 -2690
rect 828 -2686 829 -2684
rect 828 -2692 829 -2690
rect 838 -2686 839 -2684
rect 835 -2692 836 -2690
rect 838 -2692 839 -2690
rect 842 -2686 843 -2684
rect 845 -2686 846 -2684
rect 842 -2692 843 -2690
rect 845 -2692 846 -2690
rect 849 -2686 850 -2684
rect 849 -2692 850 -2690
rect 856 -2686 857 -2684
rect 856 -2692 857 -2690
rect 863 -2686 864 -2684
rect 863 -2692 864 -2690
rect 870 -2686 871 -2684
rect 873 -2686 874 -2684
rect 870 -2692 871 -2690
rect 873 -2692 874 -2690
rect 877 -2686 878 -2684
rect 877 -2692 878 -2690
rect 884 -2686 885 -2684
rect 884 -2692 885 -2690
rect 891 -2686 892 -2684
rect 894 -2686 895 -2684
rect 894 -2692 895 -2690
rect 898 -2686 899 -2684
rect 898 -2692 899 -2690
rect 905 -2686 906 -2684
rect 905 -2692 906 -2690
rect 912 -2686 913 -2684
rect 912 -2692 913 -2690
rect 919 -2686 920 -2684
rect 919 -2692 920 -2690
rect 926 -2686 927 -2684
rect 926 -2692 927 -2690
rect 933 -2686 934 -2684
rect 933 -2692 934 -2690
rect 940 -2686 941 -2684
rect 940 -2692 941 -2690
rect 947 -2686 948 -2684
rect 947 -2692 948 -2690
rect 954 -2686 955 -2684
rect 957 -2686 958 -2684
rect 954 -2692 955 -2690
rect 957 -2692 958 -2690
rect 961 -2686 962 -2684
rect 961 -2692 962 -2690
rect 968 -2686 969 -2684
rect 968 -2692 969 -2690
rect 975 -2686 976 -2684
rect 975 -2692 976 -2690
rect 982 -2686 983 -2684
rect 982 -2692 983 -2690
rect 989 -2686 990 -2684
rect 989 -2692 990 -2690
rect 996 -2686 997 -2684
rect 996 -2692 997 -2690
rect 1003 -2686 1004 -2684
rect 1003 -2692 1004 -2690
rect 1010 -2686 1011 -2684
rect 1010 -2692 1011 -2690
rect 1017 -2686 1018 -2684
rect 1017 -2692 1018 -2690
rect 1024 -2686 1025 -2684
rect 1024 -2692 1025 -2690
rect 1031 -2686 1032 -2684
rect 1034 -2686 1035 -2684
rect 1031 -2692 1032 -2690
rect 1034 -2692 1035 -2690
rect 1038 -2686 1039 -2684
rect 1038 -2692 1039 -2690
rect 1045 -2686 1046 -2684
rect 1045 -2692 1046 -2690
rect 1052 -2686 1053 -2684
rect 1052 -2692 1053 -2690
rect 1059 -2686 1060 -2684
rect 1059 -2692 1060 -2690
rect 1066 -2686 1067 -2684
rect 1066 -2692 1067 -2690
rect 1073 -2686 1074 -2684
rect 1073 -2692 1074 -2690
rect 1080 -2686 1081 -2684
rect 1080 -2692 1081 -2690
rect 1087 -2686 1088 -2684
rect 1087 -2692 1088 -2690
rect 1094 -2686 1095 -2684
rect 1097 -2686 1098 -2684
rect 1094 -2692 1095 -2690
rect 1101 -2686 1102 -2684
rect 1101 -2692 1102 -2690
rect 1108 -2686 1109 -2684
rect 1108 -2692 1109 -2690
rect 1115 -2686 1116 -2684
rect 1115 -2692 1116 -2690
rect 1122 -2686 1123 -2684
rect 1122 -2692 1123 -2690
rect 1129 -2686 1130 -2684
rect 1129 -2692 1130 -2690
rect 1136 -2686 1137 -2684
rect 1136 -2692 1137 -2690
rect 1143 -2686 1144 -2684
rect 1143 -2692 1144 -2690
rect 1150 -2686 1151 -2684
rect 1150 -2692 1151 -2690
rect 1157 -2686 1158 -2684
rect 1157 -2692 1158 -2690
rect 1164 -2686 1165 -2684
rect 1164 -2692 1165 -2690
rect 1171 -2686 1172 -2684
rect 1171 -2692 1172 -2690
rect 1178 -2686 1179 -2684
rect 1178 -2692 1179 -2690
rect 1185 -2686 1186 -2684
rect 1185 -2692 1186 -2690
rect 1192 -2686 1193 -2684
rect 1192 -2692 1193 -2690
rect 1199 -2686 1200 -2684
rect 1199 -2692 1200 -2690
rect 1206 -2686 1207 -2684
rect 1206 -2692 1207 -2690
rect 1213 -2686 1214 -2684
rect 1213 -2692 1214 -2690
rect 1220 -2686 1221 -2684
rect 1220 -2692 1221 -2690
rect 1227 -2686 1228 -2684
rect 1227 -2692 1228 -2690
rect 1234 -2686 1235 -2684
rect 1234 -2692 1235 -2690
rect 1241 -2686 1242 -2684
rect 1241 -2692 1242 -2690
rect 1248 -2686 1249 -2684
rect 1248 -2692 1249 -2690
rect 1255 -2686 1256 -2684
rect 1255 -2692 1256 -2690
rect 1262 -2686 1263 -2684
rect 1262 -2692 1263 -2690
rect 1269 -2686 1270 -2684
rect 1269 -2692 1270 -2690
rect 1276 -2686 1277 -2684
rect 1276 -2692 1277 -2690
rect 1283 -2686 1284 -2684
rect 1283 -2692 1284 -2690
rect 1290 -2686 1291 -2684
rect 1290 -2692 1291 -2690
rect 1297 -2686 1298 -2684
rect 1297 -2692 1298 -2690
rect 1304 -2686 1305 -2684
rect 1304 -2692 1305 -2690
rect 1311 -2686 1312 -2684
rect 1311 -2692 1312 -2690
rect 1318 -2686 1319 -2684
rect 1318 -2692 1319 -2690
rect 1325 -2686 1326 -2684
rect 1325 -2692 1326 -2690
rect 1332 -2686 1333 -2684
rect 1332 -2692 1333 -2690
rect 1339 -2686 1340 -2684
rect 1339 -2692 1340 -2690
rect 1346 -2686 1347 -2684
rect 1346 -2692 1347 -2690
rect 1353 -2686 1354 -2684
rect 1353 -2692 1354 -2690
rect 1360 -2686 1361 -2684
rect 1360 -2692 1361 -2690
rect 1367 -2686 1368 -2684
rect 1367 -2692 1368 -2690
rect 1374 -2686 1375 -2684
rect 1374 -2692 1375 -2690
rect 1381 -2686 1382 -2684
rect 1381 -2692 1382 -2690
rect 1388 -2686 1389 -2684
rect 1388 -2692 1389 -2690
rect 1395 -2686 1396 -2684
rect 1395 -2692 1396 -2690
rect 1402 -2686 1403 -2684
rect 1402 -2692 1403 -2690
rect 1409 -2686 1410 -2684
rect 1409 -2692 1410 -2690
rect 1416 -2686 1417 -2684
rect 1416 -2692 1417 -2690
rect 1423 -2686 1424 -2684
rect 1423 -2692 1424 -2690
rect 1430 -2686 1431 -2684
rect 1430 -2692 1431 -2690
rect 1437 -2686 1438 -2684
rect 1437 -2692 1438 -2690
rect 1444 -2686 1445 -2684
rect 1444 -2692 1445 -2690
rect 1451 -2686 1452 -2684
rect 1451 -2692 1452 -2690
rect 1458 -2686 1459 -2684
rect 1458 -2692 1459 -2690
rect 1465 -2686 1466 -2684
rect 1465 -2692 1466 -2690
rect 1472 -2686 1473 -2684
rect 1472 -2692 1473 -2690
rect 1479 -2686 1480 -2684
rect 1479 -2692 1480 -2690
rect 1486 -2686 1487 -2684
rect 1486 -2692 1487 -2690
rect 1493 -2686 1494 -2684
rect 1493 -2692 1494 -2690
rect 1500 -2686 1501 -2684
rect 1500 -2692 1501 -2690
rect 1507 -2686 1508 -2684
rect 1507 -2692 1508 -2690
rect 1514 -2686 1515 -2684
rect 1514 -2692 1515 -2690
rect 1521 -2686 1522 -2684
rect 1521 -2692 1522 -2690
rect 1528 -2686 1529 -2684
rect 1528 -2692 1529 -2690
rect 1535 -2686 1536 -2684
rect 1535 -2692 1536 -2690
rect 1542 -2686 1543 -2684
rect 1542 -2692 1543 -2690
rect 1549 -2686 1550 -2684
rect 1549 -2692 1550 -2690
rect 1556 -2686 1557 -2684
rect 1556 -2692 1557 -2690
rect 1563 -2686 1564 -2684
rect 1563 -2692 1564 -2690
rect 1570 -2686 1571 -2684
rect 1570 -2692 1571 -2690
rect 1577 -2686 1578 -2684
rect 1577 -2692 1578 -2690
rect 1584 -2686 1585 -2684
rect 1584 -2692 1585 -2690
rect 1591 -2686 1592 -2684
rect 1591 -2692 1592 -2690
rect 1598 -2686 1599 -2684
rect 1598 -2692 1599 -2690
rect 1605 -2686 1606 -2684
rect 1605 -2692 1606 -2690
rect 1612 -2686 1613 -2684
rect 1612 -2692 1613 -2690
rect 1619 -2686 1620 -2684
rect 1619 -2692 1620 -2690
rect 1626 -2686 1627 -2684
rect 1626 -2692 1627 -2690
rect 1633 -2686 1634 -2684
rect 1633 -2692 1634 -2690
rect 1640 -2686 1641 -2684
rect 1640 -2692 1641 -2690
rect 1647 -2686 1648 -2684
rect 1647 -2692 1648 -2690
rect 1654 -2686 1655 -2684
rect 1654 -2692 1655 -2690
rect 1661 -2686 1662 -2684
rect 1661 -2692 1662 -2690
rect 1668 -2686 1669 -2684
rect 1668 -2692 1669 -2690
rect 1675 -2686 1676 -2684
rect 1675 -2692 1676 -2690
rect 1682 -2686 1683 -2684
rect 1682 -2692 1683 -2690
rect 1689 -2686 1690 -2684
rect 1689 -2692 1690 -2690
rect 1696 -2686 1697 -2684
rect 1696 -2692 1697 -2690
rect 1703 -2686 1704 -2684
rect 1703 -2692 1704 -2690
rect 37 -2835 38 -2833
rect 37 -2841 38 -2839
rect 44 -2835 45 -2833
rect 44 -2841 45 -2839
rect 51 -2835 52 -2833
rect 51 -2841 52 -2839
rect 58 -2835 59 -2833
rect 58 -2841 59 -2839
rect 65 -2835 66 -2833
rect 65 -2841 66 -2839
rect 72 -2835 73 -2833
rect 72 -2841 73 -2839
rect 79 -2835 80 -2833
rect 79 -2841 80 -2839
rect 86 -2835 87 -2833
rect 89 -2835 90 -2833
rect 93 -2835 94 -2833
rect 96 -2835 97 -2833
rect 93 -2841 94 -2839
rect 96 -2841 97 -2839
rect 100 -2835 101 -2833
rect 100 -2841 101 -2839
rect 107 -2835 108 -2833
rect 110 -2835 111 -2833
rect 107 -2841 108 -2839
rect 110 -2841 111 -2839
rect 114 -2835 115 -2833
rect 114 -2841 115 -2839
rect 121 -2835 122 -2833
rect 121 -2841 122 -2839
rect 128 -2835 129 -2833
rect 131 -2835 132 -2833
rect 128 -2841 129 -2839
rect 135 -2835 136 -2833
rect 135 -2841 136 -2839
rect 142 -2835 143 -2833
rect 142 -2841 143 -2839
rect 149 -2835 150 -2833
rect 149 -2841 150 -2839
rect 156 -2835 157 -2833
rect 156 -2841 157 -2839
rect 163 -2835 164 -2833
rect 166 -2835 167 -2833
rect 163 -2841 164 -2839
rect 170 -2835 171 -2833
rect 170 -2841 171 -2839
rect 180 -2835 181 -2833
rect 177 -2841 178 -2839
rect 180 -2841 181 -2839
rect 184 -2835 185 -2833
rect 184 -2841 185 -2839
rect 191 -2841 192 -2839
rect 198 -2835 199 -2833
rect 198 -2841 199 -2839
rect 205 -2835 206 -2833
rect 205 -2841 206 -2839
rect 212 -2835 213 -2833
rect 212 -2841 213 -2839
rect 219 -2835 220 -2833
rect 219 -2841 220 -2839
rect 226 -2835 227 -2833
rect 229 -2835 230 -2833
rect 226 -2841 227 -2839
rect 229 -2841 230 -2839
rect 233 -2835 234 -2833
rect 233 -2841 234 -2839
rect 240 -2835 241 -2833
rect 240 -2841 241 -2839
rect 247 -2835 248 -2833
rect 250 -2835 251 -2833
rect 250 -2841 251 -2839
rect 254 -2835 255 -2833
rect 254 -2841 255 -2839
rect 261 -2835 262 -2833
rect 261 -2841 262 -2839
rect 268 -2835 269 -2833
rect 268 -2841 269 -2839
rect 275 -2835 276 -2833
rect 278 -2835 279 -2833
rect 275 -2841 276 -2839
rect 282 -2835 283 -2833
rect 282 -2841 283 -2839
rect 289 -2835 290 -2833
rect 289 -2841 290 -2839
rect 296 -2835 297 -2833
rect 296 -2841 297 -2839
rect 303 -2835 304 -2833
rect 303 -2841 304 -2839
rect 310 -2835 311 -2833
rect 310 -2841 311 -2839
rect 317 -2835 318 -2833
rect 317 -2841 318 -2839
rect 324 -2835 325 -2833
rect 324 -2841 325 -2839
rect 331 -2835 332 -2833
rect 331 -2841 332 -2839
rect 338 -2835 339 -2833
rect 338 -2841 339 -2839
rect 345 -2835 346 -2833
rect 345 -2841 346 -2839
rect 352 -2835 353 -2833
rect 352 -2841 353 -2839
rect 359 -2835 360 -2833
rect 359 -2841 360 -2839
rect 366 -2835 367 -2833
rect 366 -2841 367 -2839
rect 373 -2835 374 -2833
rect 373 -2841 374 -2839
rect 380 -2835 381 -2833
rect 383 -2835 384 -2833
rect 380 -2841 381 -2839
rect 387 -2835 388 -2833
rect 387 -2841 388 -2839
rect 394 -2835 395 -2833
rect 394 -2841 395 -2839
rect 401 -2835 402 -2833
rect 401 -2841 402 -2839
rect 408 -2835 409 -2833
rect 408 -2841 409 -2839
rect 415 -2835 416 -2833
rect 415 -2841 416 -2839
rect 422 -2835 423 -2833
rect 422 -2841 423 -2839
rect 429 -2835 430 -2833
rect 429 -2841 430 -2839
rect 436 -2835 437 -2833
rect 436 -2841 437 -2839
rect 443 -2835 444 -2833
rect 443 -2841 444 -2839
rect 450 -2835 451 -2833
rect 450 -2841 451 -2839
rect 457 -2835 458 -2833
rect 457 -2841 458 -2839
rect 464 -2835 465 -2833
rect 464 -2841 465 -2839
rect 471 -2835 472 -2833
rect 471 -2841 472 -2839
rect 478 -2835 479 -2833
rect 478 -2841 479 -2839
rect 485 -2835 486 -2833
rect 485 -2841 486 -2839
rect 492 -2835 493 -2833
rect 492 -2841 493 -2839
rect 499 -2835 500 -2833
rect 499 -2841 500 -2839
rect 506 -2835 507 -2833
rect 506 -2841 507 -2839
rect 513 -2835 514 -2833
rect 513 -2841 514 -2839
rect 520 -2835 521 -2833
rect 523 -2835 524 -2833
rect 520 -2841 521 -2839
rect 523 -2841 524 -2839
rect 527 -2835 528 -2833
rect 527 -2841 528 -2839
rect 534 -2835 535 -2833
rect 534 -2841 535 -2839
rect 541 -2835 542 -2833
rect 541 -2841 542 -2839
rect 548 -2835 549 -2833
rect 548 -2841 549 -2839
rect 555 -2835 556 -2833
rect 555 -2841 556 -2839
rect 562 -2835 563 -2833
rect 562 -2841 563 -2839
rect 569 -2835 570 -2833
rect 569 -2841 570 -2839
rect 576 -2835 577 -2833
rect 576 -2841 577 -2839
rect 583 -2835 584 -2833
rect 583 -2841 584 -2839
rect 590 -2835 591 -2833
rect 593 -2835 594 -2833
rect 590 -2841 591 -2839
rect 593 -2841 594 -2839
rect 597 -2835 598 -2833
rect 597 -2841 598 -2839
rect 604 -2835 605 -2833
rect 604 -2841 605 -2839
rect 611 -2835 612 -2833
rect 611 -2841 612 -2839
rect 618 -2835 619 -2833
rect 618 -2841 619 -2839
rect 625 -2835 626 -2833
rect 625 -2841 626 -2839
rect 632 -2835 633 -2833
rect 632 -2841 633 -2839
rect 639 -2835 640 -2833
rect 639 -2841 640 -2839
rect 649 -2835 650 -2833
rect 646 -2841 647 -2839
rect 649 -2841 650 -2839
rect 653 -2835 654 -2833
rect 653 -2841 654 -2839
rect 656 -2841 657 -2839
rect 660 -2835 661 -2833
rect 660 -2841 661 -2839
rect 667 -2835 668 -2833
rect 667 -2841 668 -2839
rect 674 -2835 675 -2833
rect 674 -2841 675 -2839
rect 681 -2835 682 -2833
rect 684 -2835 685 -2833
rect 684 -2841 685 -2839
rect 688 -2835 689 -2833
rect 688 -2841 689 -2839
rect 695 -2835 696 -2833
rect 695 -2841 696 -2839
rect 702 -2835 703 -2833
rect 702 -2841 703 -2839
rect 709 -2835 710 -2833
rect 709 -2841 710 -2839
rect 716 -2835 717 -2833
rect 716 -2841 717 -2839
rect 723 -2835 724 -2833
rect 723 -2841 724 -2839
rect 730 -2835 731 -2833
rect 730 -2841 731 -2839
rect 737 -2835 738 -2833
rect 737 -2841 738 -2839
rect 744 -2835 745 -2833
rect 744 -2841 745 -2839
rect 751 -2835 752 -2833
rect 751 -2841 752 -2839
rect 758 -2835 759 -2833
rect 761 -2835 762 -2833
rect 758 -2841 759 -2839
rect 761 -2841 762 -2839
rect 765 -2835 766 -2833
rect 768 -2835 769 -2833
rect 765 -2841 766 -2839
rect 768 -2841 769 -2839
rect 772 -2835 773 -2833
rect 775 -2835 776 -2833
rect 775 -2841 776 -2839
rect 779 -2835 780 -2833
rect 779 -2841 780 -2839
rect 786 -2835 787 -2833
rect 786 -2841 787 -2839
rect 793 -2835 794 -2833
rect 793 -2841 794 -2839
rect 800 -2835 801 -2833
rect 803 -2835 804 -2833
rect 800 -2841 801 -2839
rect 803 -2841 804 -2839
rect 807 -2835 808 -2833
rect 807 -2841 808 -2839
rect 814 -2835 815 -2833
rect 814 -2841 815 -2839
rect 821 -2835 822 -2833
rect 821 -2841 822 -2839
rect 828 -2835 829 -2833
rect 828 -2841 829 -2839
rect 835 -2835 836 -2833
rect 835 -2841 836 -2839
rect 842 -2835 843 -2833
rect 842 -2841 843 -2839
rect 849 -2835 850 -2833
rect 849 -2841 850 -2839
rect 856 -2835 857 -2833
rect 856 -2841 857 -2839
rect 863 -2835 864 -2833
rect 863 -2841 864 -2839
rect 870 -2835 871 -2833
rect 870 -2841 871 -2839
rect 877 -2835 878 -2833
rect 877 -2841 878 -2839
rect 884 -2835 885 -2833
rect 887 -2835 888 -2833
rect 884 -2841 885 -2839
rect 887 -2841 888 -2839
rect 891 -2835 892 -2833
rect 894 -2835 895 -2833
rect 891 -2841 892 -2839
rect 898 -2835 899 -2833
rect 901 -2835 902 -2833
rect 898 -2841 899 -2839
rect 901 -2841 902 -2839
rect 905 -2835 906 -2833
rect 905 -2841 906 -2839
rect 912 -2835 913 -2833
rect 912 -2841 913 -2839
rect 919 -2835 920 -2833
rect 919 -2841 920 -2839
rect 926 -2835 927 -2833
rect 926 -2841 927 -2839
rect 933 -2835 934 -2833
rect 933 -2841 934 -2839
rect 940 -2835 941 -2833
rect 940 -2841 941 -2839
rect 947 -2835 948 -2833
rect 947 -2841 948 -2839
rect 954 -2835 955 -2833
rect 954 -2841 955 -2839
rect 961 -2835 962 -2833
rect 961 -2841 962 -2839
rect 968 -2835 969 -2833
rect 968 -2841 969 -2839
rect 975 -2835 976 -2833
rect 975 -2841 976 -2839
rect 982 -2835 983 -2833
rect 985 -2835 986 -2833
rect 982 -2841 983 -2839
rect 989 -2835 990 -2833
rect 989 -2841 990 -2839
rect 996 -2835 997 -2833
rect 999 -2835 1000 -2833
rect 996 -2841 997 -2839
rect 999 -2841 1000 -2839
rect 1003 -2835 1004 -2833
rect 1003 -2841 1004 -2839
rect 1010 -2835 1011 -2833
rect 1010 -2841 1011 -2839
rect 1017 -2835 1018 -2833
rect 1017 -2841 1018 -2839
rect 1024 -2835 1025 -2833
rect 1024 -2841 1025 -2839
rect 1031 -2835 1032 -2833
rect 1031 -2841 1032 -2839
rect 1038 -2835 1039 -2833
rect 1038 -2841 1039 -2839
rect 1045 -2835 1046 -2833
rect 1048 -2835 1049 -2833
rect 1045 -2841 1046 -2839
rect 1048 -2841 1049 -2839
rect 1052 -2835 1053 -2833
rect 1052 -2841 1053 -2839
rect 1059 -2835 1060 -2833
rect 1059 -2841 1060 -2839
rect 1066 -2835 1067 -2833
rect 1066 -2841 1067 -2839
rect 1073 -2835 1074 -2833
rect 1073 -2841 1074 -2839
rect 1080 -2835 1081 -2833
rect 1080 -2841 1081 -2839
rect 1087 -2835 1088 -2833
rect 1087 -2841 1088 -2839
rect 1094 -2835 1095 -2833
rect 1097 -2835 1098 -2833
rect 1097 -2841 1098 -2839
rect 1101 -2835 1102 -2833
rect 1101 -2841 1102 -2839
rect 1108 -2835 1109 -2833
rect 1108 -2841 1109 -2839
rect 1115 -2835 1116 -2833
rect 1115 -2841 1116 -2839
rect 1118 -2841 1119 -2839
rect 1122 -2835 1123 -2833
rect 1122 -2841 1123 -2839
rect 1129 -2835 1130 -2833
rect 1129 -2841 1130 -2839
rect 1136 -2835 1137 -2833
rect 1136 -2841 1137 -2839
rect 1143 -2835 1144 -2833
rect 1143 -2841 1144 -2839
rect 1150 -2835 1151 -2833
rect 1150 -2841 1151 -2839
rect 1157 -2835 1158 -2833
rect 1157 -2841 1158 -2839
rect 1164 -2835 1165 -2833
rect 1164 -2841 1165 -2839
rect 1171 -2835 1172 -2833
rect 1171 -2841 1172 -2839
rect 1178 -2835 1179 -2833
rect 1178 -2841 1179 -2839
rect 1185 -2835 1186 -2833
rect 1188 -2835 1189 -2833
rect 1185 -2841 1186 -2839
rect 1188 -2841 1189 -2839
rect 1192 -2835 1193 -2833
rect 1192 -2841 1193 -2839
rect 1199 -2835 1200 -2833
rect 1199 -2841 1200 -2839
rect 1206 -2835 1207 -2833
rect 1206 -2841 1207 -2839
rect 1213 -2835 1214 -2833
rect 1213 -2841 1214 -2839
rect 1220 -2835 1221 -2833
rect 1220 -2841 1221 -2839
rect 1227 -2835 1228 -2833
rect 1227 -2841 1228 -2839
rect 1234 -2835 1235 -2833
rect 1234 -2841 1235 -2839
rect 1241 -2835 1242 -2833
rect 1241 -2841 1242 -2839
rect 1248 -2835 1249 -2833
rect 1248 -2841 1249 -2839
rect 1255 -2835 1256 -2833
rect 1255 -2841 1256 -2839
rect 1262 -2835 1263 -2833
rect 1262 -2841 1263 -2839
rect 1269 -2835 1270 -2833
rect 1269 -2841 1270 -2839
rect 1276 -2835 1277 -2833
rect 1279 -2835 1280 -2833
rect 1279 -2841 1280 -2839
rect 1283 -2835 1284 -2833
rect 1283 -2841 1284 -2839
rect 1290 -2835 1291 -2833
rect 1290 -2841 1291 -2839
rect 1297 -2835 1298 -2833
rect 1297 -2841 1298 -2839
rect 1304 -2835 1305 -2833
rect 1304 -2841 1305 -2839
rect 1311 -2835 1312 -2833
rect 1311 -2841 1312 -2839
rect 1318 -2835 1319 -2833
rect 1318 -2841 1319 -2839
rect 1325 -2835 1326 -2833
rect 1325 -2841 1326 -2839
rect 1332 -2835 1333 -2833
rect 1332 -2841 1333 -2839
rect 1339 -2835 1340 -2833
rect 1339 -2841 1340 -2839
rect 1346 -2835 1347 -2833
rect 1346 -2841 1347 -2839
rect 1353 -2835 1354 -2833
rect 1353 -2841 1354 -2839
rect 1360 -2835 1361 -2833
rect 1360 -2841 1361 -2839
rect 1367 -2835 1368 -2833
rect 1367 -2841 1368 -2839
rect 1374 -2835 1375 -2833
rect 1374 -2841 1375 -2839
rect 1381 -2835 1382 -2833
rect 1381 -2841 1382 -2839
rect 1388 -2835 1389 -2833
rect 1388 -2841 1389 -2839
rect 1395 -2835 1396 -2833
rect 1395 -2841 1396 -2839
rect 1402 -2835 1403 -2833
rect 1402 -2841 1403 -2839
rect 1409 -2835 1410 -2833
rect 1409 -2841 1410 -2839
rect 1416 -2835 1417 -2833
rect 1416 -2841 1417 -2839
rect 1423 -2835 1424 -2833
rect 1423 -2841 1424 -2839
rect 1430 -2835 1431 -2833
rect 1430 -2841 1431 -2839
rect 1437 -2835 1438 -2833
rect 1437 -2841 1438 -2839
rect 1444 -2835 1445 -2833
rect 1444 -2841 1445 -2839
rect 1451 -2835 1452 -2833
rect 1451 -2841 1452 -2839
rect 1458 -2835 1459 -2833
rect 1458 -2841 1459 -2839
rect 1465 -2835 1466 -2833
rect 1465 -2841 1466 -2839
rect 1472 -2835 1473 -2833
rect 1472 -2841 1473 -2839
rect 1479 -2835 1480 -2833
rect 1479 -2841 1480 -2839
rect 1486 -2835 1487 -2833
rect 1486 -2841 1487 -2839
rect 1493 -2835 1494 -2833
rect 1493 -2841 1494 -2839
rect 1500 -2835 1501 -2833
rect 1500 -2841 1501 -2839
rect 1507 -2835 1508 -2833
rect 1510 -2835 1511 -2833
rect 1507 -2841 1508 -2839
rect 1510 -2841 1511 -2839
rect 1514 -2835 1515 -2833
rect 1514 -2841 1515 -2839
rect 1521 -2835 1522 -2833
rect 1521 -2841 1522 -2839
rect 1528 -2835 1529 -2833
rect 1528 -2841 1529 -2839
rect 1535 -2835 1536 -2833
rect 1535 -2841 1536 -2839
rect 1542 -2835 1543 -2833
rect 1542 -2841 1543 -2839
rect 1549 -2835 1550 -2833
rect 1549 -2841 1550 -2839
rect 1556 -2835 1557 -2833
rect 1556 -2841 1557 -2839
rect 30 -2946 31 -2944
rect 30 -2952 31 -2950
rect 37 -2946 38 -2944
rect 37 -2952 38 -2950
rect 44 -2946 45 -2944
rect 44 -2952 45 -2950
rect 51 -2946 52 -2944
rect 51 -2952 52 -2950
rect 58 -2946 59 -2944
rect 58 -2952 59 -2950
rect 65 -2946 66 -2944
rect 65 -2952 66 -2950
rect 72 -2946 73 -2944
rect 75 -2946 76 -2944
rect 79 -2946 80 -2944
rect 79 -2952 80 -2950
rect 86 -2946 87 -2944
rect 86 -2952 87 -2950
rect 93 -2946 94 -2944
rect 93 -2952 94 -2950
rect 100 -2946 101 -2944
rect 100 -2952 101 -2950
rect 107 -2946 108 -2944
rect 107 -2952 108 -2950
rect 114 -2946 115 -2944
rect 117 -2946 118 -2944
rect 114 -2952 115 -2950
rect 121 -2946 122 -2944
rect 121 -2952 122 -2950
rect 128 -2946 129 -2944
rect 128 -2952 129 -2950
rect 135 -2946 136 -2944
rect 135 -2952 136 -2950
rect 142 -2946 143 -2944
rect 142 -2952 143 -2950
rect 149 -2946 150 -2944
rect 149 -2952 150 -2950
rect 159 -2952 160 -2950
rect 163 -2946 164 -2944
rect 163 -2952 164 -2950
rect 170 -2946 171 -2944
rect 170 -2952 171 -2950
rect 177 -2946 178 -2944
rect 177 -2952 178 -2950
rect 180 -2952 181 -2950
rect 184 -2946 185 -2944
rect 184 -2952 185 -2950
rect 191 -2946 192 -2944
rect 191 -2952 192 -2950
rect 198 -2946 199 -2944
rect 198 -2952 199 -2950
rect 205 -2946 206 -2944
rect 205 -2952 206 -2950
rect 212 -2946 213 -2944
rect 212 -2952 213 -2950
rect 219 -2946 220 -2944
rect 219 -2952 220 -2950
rect 226 -2946 227 -2944
rect 226 -2952 227 -2950
rect 233 -2946 234 -2944
rect 233 -2952 234 -2950
rect 240 -2946 241 -2944
rect 240 -2952 241 -2950
rect 247 -2946 248 -2944
rect 250 -2946 251 -2944
rect 250 -2952 251 -2950
rect 254 -2946 255 -2944
rect 257 -2946 258 -2944
rect 254 -2952 255 -2950
rect 257 -2952 258 -2950
rect 264 -2946 265 -2944
rect 261 -2952 262 -2950
rect 264 -2952 265 -2950
rect 268 -2946 269 -2944
rect 268 -2952 269 -2950
rect 275 -2946 276 -2944
rect 275 -2952 276 -2950
rect 282 -2946 283 -2944
rect 282 -2952 283 -2950
rect 289 -2946 290 -2944
rect 289 -2952 290 -2950
rect 296 -2946 297 -2944
rect 296 -2952 297 -2950
rect 303 -2946 304 -2944
rect 303 -2952 304 -2950
rect 310 -2946 311 -2944
rect 310 -2952 311 -2950
rect 317 -2946 318 -2944
rect 317 -2952 318 -2950
rect 324 -2946 325 -2944
rect 324 -2952 325 -2950
rect 331 -2946 332 -2944
rect 331 -2952 332 -2950
rect 338 -2946 339 -2944
rect 338 -2952 339 -2950
rect 345 -2946 346 -2944
rect 345 -2952 346 -2950
rect 352 -2946 353 -2944
rect 352 -2952 353 -2950
rect 359 -2946 360 -2944
rect 359 -2952 360 -2950
rect 366 -2946 367 -2944
rect 366 -2952 367 -2950
rect 373 -2952 374 -2950
rect 376 -2952 377 -2950
rect 380 -2946 381 -2944
rect 380 -2952 381 -2950
rect 387 -2946 388 -2944
rect 387 -2952 388 -2950
rect 394 -2946 395 -2944
rect 394 -2952 395 -2950
rect 401 -2946 402 -2944
rect 404 -2946 405 -2944
rect 401 -2952 402 -2950
rect 404 -2952 405 -2950
rect 408 -2946 409 -2944
rect 411 -2946 412 -2944
rect 408 -2952 409 -2950
rect 415 -2946 416 -2944
rect 415 -2952 416 -2950
rect 422 -2946 423 -2944
rect 422 -2952 423 -2950
rect 429 -2946 430 -2944
rect 429 -2952 430 -2950
rect 436 -2946 437 -2944
rect 436 -2952 437 -2950
rect 443 -2946 444 -2944
rect 443 -2952 444 -2950
rect 450 -2946 451 -2944
rect 450 -2952 451 -2950
rect 457 -2946 458 -2944
rect 457 -2952 458 -2950
rect 464 -2946 465 -2944
rect 464 -2952 465 -2950
rect 471 -2946 472 -2944
rect 474 -2946 475 -2944
rect 471 -2952 472 -2950
rect 474 -2952 475 -2950
rect 478 -2946 479 -2944
rect 478 -2952 479 -2950
rect 481 -2952 482 -2950
rect 485 -2946 486 -2944
rect 485 -2952 486 -2950
rect 492 -2946 493 -2944
rect 492 -2952 493 -2950
rect 499 -2946 500 -2944
rect 502 -2946 503 -2944
rect 502 -2952 503 -2950
rect 506 -2946 507 -2944
rect 506 -2952 507 -2950
rect 513 -2946 514 -2944
rect 513 -2952 514 -2950
rect 520 -2946 521 -2944
rect 520 -2952 521 -2950
rect 527 -2946 528 -2944
rect 527 -2952 528 -2950
rect 534 -2946 535 -2944
rect 534 -2952 535 -2950
rect 541 -2946 542 -2944
rect 541 -2952 542 -2950
rect 548 -2946 549 -2944
rect 548 -2952 549 -2950
rect 555 -2946 556 -2944
rect 555 -2952 556 -2950
rect 562 -2946 563 -2944
rect 565 -2946 566 -2944
rect 565 -2952 566 -2950
rect 569 -2946 570 -2944
rect 569 -2952 570 -2950
rect 576 -2946 577 -2944
rect 576 -2952 577 -2950
rect 583 -2946 584 -2944
rect 583 -2952 584 -2950
rect 590 -2946 591 -2944
rect 590 -2952 591 -2950
rect 597 -2946 598 -2944
rect 597 -2952 598 -2950
rect 607 -2946 608 -2944
rect 604 -2952 605 -2950
rect 607 -2952 608 -2950
rect 611 -2946 612 -2944
rect 611 -2952 612 -2950
rect 618 -2946 619 -2944
rect 618 -2952 619 -2950
rect 625 -2946 626 -2944
rect 625 -2952 626 -2950
rect 632 -2946 633 -2944
rect 632 -2952 633 -2950
rect 635 -2952 636 -2950
rect 639 -2946 640 -2944
rect 639 -2952 640 -2950
rect 646 -2946 647 -2944
rect 646 -2952 647 -2950
rect 653 -2946 654 -2944
rect 653 -2952 654 -2950
rect 660 -2946 661 -2944
rect 660 -2952 661 -2950
rect 667 -2946 668 -2944
rect 670 -2946 671 -2944
rect 667 -2952 668 -2950
rect 670 -2952 671 -2950
rect 674 -2946 675 -2944
rect 674 -2952 675 -2950
rect 681 -2946 682 -2944
rect 681 -2952 682 -2950
rect 688 -2952 689 -2950
rect 691 -2952 692 -2950
rect 695 -2946 696 -2944
rect 695 -2952 696 -2950
rect 702 -2946 703 -2944
rect 702 -2952 703 -2950
rect 705 -2952 706 -2950
rect 709 -2946 710 -2944
rect 709 -2952 710 -2950
rect 716 -2946 717 -2944
rect 716 -2952 717 -2950
rect 723 -2946 724 -2944
rect 723 -2952 724 -2950
rect 730 -2946 731 -2944
rect 733 -2946 734 -2944
rect 730 -2952 731 -2950
rect 733 -2952 734 -2950
rect 737 -2946 738 -2944
rect 737 -2952 738 -2950
rect 744 -2946 745 -2944
rect 744 -2952 745 -2950
rect 751 -2946 752 -2944
rect 751 -2952 752 -2950
rect 761 -2946 762 -2944
rect 758 -2952 759 -2950
rect 761 -2952 762 -2950
rect 765 -2946 766 -2944
rect 765 -2952 766 -2950
rect 772 -2946 773 -2944
rect 772 -2952 773 -2950
rect 779 -2946 780 -2944
rect 779 -2952 780 -2950
rect 786 -2946 787 -2944
rect 786 -2952 787 -2950
rect 793 -2946 794 -2944
rect 793 -2952 794 -2950
rect 800 -2946 801 -2944
rect 800 -2952 801 -2950
rect 807 -2946 808 -2944
rect 807 -2952 808 -2950
rect 814 -2946 815 -2944
rect 814 -2952 815 -2950
rect 821 -2946 822 -2944
rect 821 -2952 822 -2950
rect 828 -2946 829 -2944
rect 828 -2952 829 -2950
rect 835 -2946 836 -2944
rect 835 -2952 836 -2950
rect 842 -2946 843 -2944
rect 842 -2952 843 -2950
rect 849 -2946 850 -2944
rect 849 -2952 850 -2950
rect 856 -2946 857 -2944
rect 856 -2952 857 -2950
rect 863 -2946 864 -2944
rect 866 -2946 867 -2944
rect 863 -2952 864 -2950
rect 866 -2952 867 -2950
rect 870 -2946 871 -2944
rect 870 -2952 871 -2950
rect 877 -2946 878 -2944
rect 877 -2952 878 -2950
rect 884 -2946 885 -2944
rect 884 -2952 885 -2950
rect 891 -2946 892 -2944
rect 891 -2952 892 -2950
rect 898 -2946 899 -2944
rect 898 -2952 899 -2950
rect 905 -2946 906 -2944
rect 905 -2952 906 -2950
rect 912 -2946 913 -2944
rect 915 -2946 916 -2944
rect 912 -2952 913 -2950
rect 919 -2946 920 -2944
rect 919 -2952 920 -2950
rect 926 -2946 927 -2944
rect 929 -2946 930 -2944
rect 926 -2952 927 -2950
rect 929 -2952 930 -2950
rect 936 -2946 937 -2944
rect 933 -2952 934 -2950
rect 936 -2952 937 -2950
rect 940 -2946 941 -2944
rect 940 -2952 941 -2950
rect 947 -2946 948 -2944
rect 947 -2952 948 -2950
rect 954 -2946 955 -2944
rect 954 -2952 955 -2950
rect 961 -2946 962 -2944
rect 961 -2952 962 -2950
rect 968 -2946 969 -2944
rect 968 -2952 969 -2950
rect 975 -2946 976 -2944
rect 975 -2952 976 -2950
rect 982 -2946 983 -2944
rect 982 -2952 983 -2950
rect 989 -2946 990 -2944
rect 989 -2952 990 -2950
rect 996 -2946 997 -2944
rect 996 -2952 997 -2950
rect 999 -2952 1000 -2950
rect 1003 -2946 1004 -2944
rect 1003 -2952 1004 -2950
rect 1010 -2946 1011 -2944
rect 1010 -2952 1011 -2950
rect 1017 -2946 1018 -2944
rect 1017 -2952 1018 -2950
rect 1020 -2952 1021 -2950
rect 1024 -2946 1025 -2944
rect 1027 -2946 1028 -2944
rect 1024 -2952 1025 -2950
rect 1031 -2946 1032 -2944
rect 1031 -2952 1032 -2950
rect 1038 -2946 1039 -2944
rect 1038 -2952 1039 -2950
rect 1045 -2946 1046 -2944
rect 1045 -2952 1046 -2950
rect 1052 -2946 1053 -2944
rect 1052 -2952 1053 -2950
rect 1059 -2946 1060 -2944
rect 1059 -2952 1060 -2950
rect 1066 -2946 1067 -2944
rect 1066 -2952 1067 -2950
rect 1073 -2946 1074 -2944
rect 1073 -2952 1074 -2950
rect 1080 -2946 1081 -2944
rect 1080 -2952 1081 -2950
rect 1087 -2946 1088 -2944
rect 1087 -2952 1088 -2950
rect 1094 -2946 1095 -2944
rect 1094 -2952 1095 -2950
rect 1101 -2946 1102 -2944
rect 1101 -2952 1102 -2950
rect 1108 -2946 1109 -2944
rect 1108 -2952 1109 -2950
rect 1115 -2946 1116 -2944
rect 1115 -2952 1116 -2950
rect 1122 -2946 1123 -2944
rect 1122 -2952 1123 -2950
rect 1129 -2946 1130 -2944
rect 1129 -2952 1130 -2950
rect 1136 -2946 1137 -2944
rect 1136 -2952 1137 -2950
rect 1143 -2946 1144 -2944
rect 1143 -2952 1144 -2950
rect 1150 -2946 1151 -2944
rect 1150 -2952 1151 -2950
rect 1157 -2946 1158 -2944
rect 1157 -2952 1158 -2950
rect 1164 -2946 1165 -2944
rect 1164 -2952 1165 -2950
rect 1171 -2946 1172 -2944
rect 1171 -2952 1172 -2950
rect 1178 -2946 1179 -2944
rect 1178 -2952 1179 -2950
rect 1185 -2946 1186 -2944
rect 1185 -2952 1186 -2950
rect 1192 -2946 1193 -2944
rect 1192 -2952 1193 -2950
rect 1199 -2946 1200 -2944
rect 1202 -2946 1203 -2944
rect 1206 -2946 1207 -2944
rect 1206 -2952 1207 -2950
rect 1213 -2946 1214 -2944
rect 1213 -2952 1214 -2950
rect 1220 -2946 1221 -2944
rect 1220 -2952 1221 -2950
rect 1227 -2946 1228 -2944
rect 1227 -2952 1228 -2950
rect 1234 -2946 1235 -2944
rect 1234 -2952 1235 -2950
rect 1241 -2946 1242 -2944
rect 1241 -2952 1242 -2950
rect 1248 -2946 1249 -2944
rect 1248 -2952 1249 -2950
rect 1255 -2946 1256 -2944
rect 1255 -2952 1256 -2950
rect 1262 -2946 1263 -2944
rect 1262 -2952 1263 -2950
rect 1269 -2946 1270 -2944
rect 1269 -2952 1270 -2950
rect 1276 -2946 1277 -2944
rect 1276 -2952 1277 -2950
rect 1283 -2946 1284 -2944
rect 1283 -2952 1284 -2950
rect 1290 -2946 1291 -2944
rect 1290 -2952 1291 -2950
rect 1297 -2946 1298 -2944
rect 1297 -2952 1298 -2950
rect 1304 -2946 1305 -2944
rect 1304 -2952 1305 -2950
rect 1311 -2946 1312 -2944
rect 1311 -2952 1312 -2950
rect 1318 -2946 1319 -2944
rect 1318 -2952 1319 -2950
rect 1325 -2946 1326 -2944
rect 1325 -2952 1326 -2950
rect 1332 -2946 1333 -2944
rect 1332 -2952 1333 -2950
rect 1339 -2946 1340 -2944
rect 1339 -2952 1340 -2950
rect 1346 -2946 1347 -2944
rect 1346 -2952 1347 -2950
rect 1353 -2946 1354 -2944
rect 1353 -2952 1354 -2950
rect 1360 -2946 1361 -2944
rect 1360 -2952 1361 -2950
rect 1367 -2946 1368 -2944
rect 1367 -2952 1368 -2950
rect 1374 -2946 1375 -2944
rect 1374 -2952 1375 -2950
rect 1381 -2946 1382 -2944
rect 1381 -2952 1382 -2950
rect 1388 -2946 1389 -2944
rect 1388 -2952 1389 -2950
rect 1395 -2946 1396 -2944
rect 1395 -2952 1396 -2950
rect 1402 -2946 1403 -2944
rect 1402 -2952 1403 -2950
rect 1409 -2946 1410 -2944
rect 1409 -2952 1410 -2950
rect 1416 -2946 1417 -2944
rect 1416 -2952 1417 -2950
rect 1423 -2946 1424 -2944
rect 1423 -2952 1424 -2950
rect 1430 -2946 1431 -2944
rect 1430 -2952 1431 -2950
rect 1437 -2946 1438 -2944
rect 1437 -2952 1438 -2950
rect 1447 -2946 1448 -2944
rect 1444 -2952 1445 -2950
rect 1447 -2952 1448 -2950
rect 1451 -2946 1452 -2944
rect 1451 -2952 1452 -2950
rect 1458 -2946 1459 -2944
rect 1458 -2952 1459 -2950
rect 1465 -2946 1466 -2944
rect 1465 -2952 1466 -2950
rect 1479 -2946 1480 -2944
rect 1479 -2952 1480 -2950
rect 1486 -2946 1487 -2944
rect 1486 -2952 1487 -2950
rect 1493 -2946 1494 -2944
rect 1493 -2952 1494 -2950
rect 1500 -2946 1501 -2944
rect 1500 -2952 1501 -2950
rect 37 -3065 38 -3063
rect 37 -3071 38 -3069
rect 44 -3065 45 -3063
rect 44 -3071 45 -3069
rect 51 -3065 52 -3063
rect 51 -3071 52 -3069
rect 58 -3065 59 -3063
rect 58 -3071 59 -3069
rect 65 -3065 66 -3063
rect 65 -3071 66 -3069
rect 72 -3065 73 -3063
rect 72 -3071 73 -3069
rect 79 -3065 80 -3063
rect 79 -3071 80 -3069
rect 86 -3065 87 -3063
rect 86 -3071 87 -3069
rect 96 -3065 97 -3063
rect 93 -3071 94 -3069
rect 96 -3071 97 -3069
rect 100 -3065 101 -3063
rect 100 -3071 101 -3069
rect 107 -3065 108 -3063
rect 107 -3071 108 -3069
rect 114 -3065 115 -3063
rect 114 -3071 115 -3069
rect 121 -3065 122 -3063
rect 124 -3065 125 -3063
rect 121 -3071 122 -3069
rect 128 -3065 129 -3063
rect 128 -3071 129 -3069
rect 135 -3065 136 -3063
rect 135 -3071 136 -3069
rect 142 -3065 143 -3063
rect 142 -3071 143 -3069
rect 149 -3065 150 -3063
rect 149 -3071 150 -3069
rect 156 -3065 157 -3063
rect 156 -3071 157 -3069
rect 163 -3065 164 -3063
rect 163 -3071 164 -3069
rect 170 -3065 171 -3063
rect 170 -3071 171 -3069
rect 177 -3065 178 -3063
rect 177 -3071 178 -3069
rect 180 -3071 181 -3069
rect 184 -3065 185 -3063
rect 184 -3071 185 -3069
rect 191 -3065 192 -3063
rect 191 -3071 192 -3069
rect 201 -3065 202 -3063
rect 198 -3071 199 -3069
rect 201 -3071 202 -3069
rect 205 -3065 206 -3063
rect 205 -3071 206 -3069
rect 212 -3065 213 -3063
rect 212 -3071 213 -3069
rect 222 -3071 223 -3069
rect 226 -3065 227 -3063
rect 226 -3071 227 -3069
rect 233 -3065 234 -3063
rect 233 -3071 234 -3069
rect 243 -3065 244 -3063
rect 240 -3071 241 -3069
rect 243 -3071 244 -3069
rect 247 -3065 248 -3063
rect 250 -3065 251 -3063
rect 247 -3071 248 -3069
rect 250 -3071 251 -3069
rect 254 -3065 255 -3063
rect 254 -3071 255 -3069
rect 261 -3065 262 -3063
rect 264 -3065 265 -3063
rect 261 -3071 262 -3069
rect 268 -3065 269 -3063
rect 268 -3071 269 -3069
rect 275 -3065 276 -3063
rect 275 -3071 276 -3069
rect 282 -3065 283 -3063
rect 282 -3071 283 -3069
rect 289 -3065 290 -3063
rect 289 -3071 290 -3069
rect 296 -3065 297 -3063
rect 296 -3071 297 -3069
rect 299 -3071 300 -3069
rect 303 -3065 304 -3063
rect 303 -3071 304 -3069
rect 310 -3065 311 -3063
rect 310 -3071 311 -3069
rect 317 -3065 318 -3063
rect 317 -3071 318 -3069
rect 324 -3065 325 -3063
rect 324 -3071 325 -3069
rect 331 -3065 332 -3063
rect 331 -3071 332 -3069
rect 338 -3065 339 -3063
rect 338 -3071 339 -3069
rect 345 -3065 346 -3063
rect 345 -3071 346 -3069
rect 352 -3065 353 -3063
rect 355 -3065 356 -3063
rect 352 -3071 353 -3069
rect 355 -3071 356 -3069
rect 359 -3065 360 -3063
rect 359 -3071 360 -3069
rect 366 -3065 367 -3063
rect 366 -3071 367 -3069
rect 373 -3065 374 -3063
rect 373 -3071 374 -3069
rect 380 -3065 381 -3063
rect 380 -3071 381 -3069
rect 387 -3065 388 -3063
rect 387 -3071 388 -3069
rect 394 -3065 395 -3063
rect 394 -3071 395 -3069
rect 401 -3065 402 -3063
rect 401 -3071 402 -3069
rect 408 -3065 409 -3063
rect 411 -3065 412 -3063
rect 408 -3071 409 -3069
rect 415 -3065 416 -3063
rect 415 -3071 416 -3069
rect 422 -3065 423 -3063
rect 422 -3071 423 -3069
rect 429 -3065 430 -3063
rect 429 -3071 430 -3069
rect 436 -3065 437 -3063
rect 436 -3071 437 -3069
rect 443 -3065 444 -3063
rect 443 -3071 444 -3069
rect 450 -3065 451 -3063
rect 450 -3071 451 -3069
rect 457 -3065 458 -3063
rect 457 -3071 458 -3069
rect 464 -3065 465 -3063
rect 464 -3071 465 -3069
rect 471 -3065 472 -3063
rect 471 -3071 472 -3069
rect 478 -3065 479 -3063
rect 478 -3071 479 -3069
rect 485 -3065 486 -3063
rect 485 -3071 486 -3069
rect 492 -3065 493 -3063
rect 492 -3071 493 -3069
rect 499 -3065 500 -3063
rect 499 -3071 500 -3069
rect 506 -3065 507 -3063
rect 506 -3071 507 -3069
rect 513 -3065 514 -3063
rect 513 -3071 514 -3069
rect 520 -3065 521 -3063
rect 523 -3065 524 -3063
rect 520 -3071 521 -3069
rect 523 -3071 524 -3069
rect 527 -3065 528 -3063
rect 527 -3071 528 -3069
rect 534 -3065 535 -3063
rect 534 -3071 535 -3069
rect 541 -3065 542 -3063
rect 541 -3071 542 -3069
rect 548 -3065 549 -3063
rect 548 -3071 549 -3069
rect 555 -3065 556 -3063
rect 555 -3071 556 -3069
rect 562 -3065 563 -3063
rect 562 -3071 563 -3069
rect 569 -3065 570 -3063
rect 569 -3071 570 -3069
rect 576 -3065 577 -3063
rect 576 -3071 577 -3069
rect 583 -3065 584 -3063
rect 583 -3071 584 -3069
rect 590 -3065 591 -3063
rect 590 -3071 591 -3069
rect 597 -3065 598 -3063
rect 597 -3071 598 -3069
rect 604 -3065 605 -3063
rect 607 -3065 608 -3063
rect 604 -3071 605 -3069
rect 611 -3065 612 -3063
rect 611 -3071 612 -3069
rect 618 -3065 619 -3063
rect 621 -3065 622 -3063
rect 618 -3071 619 -3069
rect 621 -3071 622 -3069
rect 625 -3065 626 -3063
rect 625 -3071 626 -3069
rect 632 -3065 633 -3063
rect 632 -3071 633 -3069
rect 639 -3065 640 -3063
rect 642 -3065 643 -3063
rect 642 -3071 643 -3069
rect 646 -3065 647 -3063
rect 646 -3071 647 -3069
rect 653 -3065 654 -3063
rect 653 -3071 654 -3069
rect 660 -3065 661 -3063
rect 660 -3071 661 -3069
rect 667 -3065 668 -3063
rect 667 -3071 668 -3069
rect 674 -3065 675 -3063
rect 674 -3071 675 -3069
rect 681 -3065 682 -3063
rect 684 -3065 685 -3063
rect 681 -3071 682 -3069
rect 684 -3071 685 -3069
rect 688 -3065 689 -3063
rect 688 -3071 689 -3069
rect 695 -3065 696 -3063
rect 695 -3071 696 -3069
rect 702 -3065 703 -3063
rect 705 -3065 706 -3063
rect 702 -3071 703 -3069
rect 705 -3071 706 -3069
rect 709 -3065 710 -3063
rect 709 -3071 710 -3069
rect 716 -3065 717 -3063
rect 716 -3071 717 -3069
rect 723 -3065 724 -3063
rect 723 -3071 724 -3069
rect 730 -3065 731 -3063
rect 730 -3071 731 -3069
rect 740 -3065 741 -3063
rect 737 -3071 738 -3069
rect 740 -3071 741 -3069
rect 744 -3065 745 -3063
rect 744 -3071 745 -3069
rect 751 -3065 752 -3063
rect 751 -3071 752 -3069
rect 758 -3065 759 -3063
rect 758 -3071 759 -3069
rect 765 -3065 766 -3063
rect 765 -3071 766 -3069
rect 772 -3065 773 -3063
rect 772 -3071 773 -3069
rect 779 -3065 780 -3063
rect 779 -3071 780 -3069
rect 786 -3065 787 -3063
rect 786 -3071 787 -3069
rect 796 -3065 797 -3063
rect 793 -3071 794 -3069
rect 796 -3071 797 -3069
rect 800 -3065 801 -3063
rect 800 -3071 801 -3069
rect 807 -3065 808 -3063
rect 807 -3071 808 -3069
rect 814 -3065 815 -3063
rect 814 -3071 815 -3069
rect 821 -3065 822 -3063
rect 821 -3071 822 -3069
rect 828 -3065 829 -3063
rect 828 -3071 829 -3069
rect 835 -3065 836 -3063
rect 835 -3071 836 -3069
rect 842 -3065 843 -3063
rect 842 -3071 843 -3069
rect 849 -3065 850 -3063
rect 852 -3065 853 -3063
rect 849 -3071 850 -3069
rect 856 -3065 857 -3063
rect 856 -3071 857 -3069
rect 863 -3065 864 -3063
rect 863 -3071 864 -3069
rect 870 -3065 871 -3063
rect 873 -3065 874 -3063
rect 870 -3071 871 -3069
rect 873 -3071 874 -3069
rect 877 -3065 878 -3063
rect 877 -3071 878 -3069
rect 884 -3065 885 -3063
rect 884 -3071 885 -3069
rect 891 -3065 892 -3063
rect 891 -3071 892 -3069
rect 898 -3065 899 -3063
rect 898 -3071 899 -3069
rect 905 -3065 906 -3063
rect 905 -3071 906 -3069
rect 912 -3065 913 -3063
rect 912 -3071 913 -3069
rect 919 -3065 920 -3063
rect 922 -3065 923 -3063
rect 919 -3071 920 -3069
rect 926 -3065 927 -3063
rect 926 -3071 927 -3069
rect 929 -3071 930 -3069
rect 933 -3065 934 -3063
rect 933 -3071 934 -3069
rect 940 -3065 941 -3063
rect 940 -3071 941 -3069
rect 947 -3065 948 -3063
rect 947 -3071 948 -3069
rect 954 -3065 955 -3063
rect 954 -3071 955 -3069
rect 961 -3065 962 -3063
rect 961 -3071 962 -3069
rect 964 -3071 965 -3069
rect 968 -3065 969 -3063
rect 968 -3071 969 -3069
rect 975 -3065 976 -3063
rect 975 -3071 976 -3069
rect 982 -3065 983 -3063
rect 982 -3071 983 -3069
rect 989 -3065 990 -3063
rect 989 -3071 990 -3069
rect 996 -3065 997 -3063
rect 999 -3065 1000 -3063
rect 996 -3071 997 -3069
rect 1003 -3065 1004 -3063
rect 1003 -3071 1004 -3069
rect 1010 -3065 1011 -3063
rect 1010 -3071 1011 -3069
rect 1017 -3065 1018 -3063
rect 1017 -3071 1018 -3069
rect 1024 -3065 1025 -3063
rect 1024 -3071 1025 -3069
rect 1031 -3065 1032 -3063
rect 1031 -3071 1032 -3069
rect 1038 -3065 1039 -3063
rect 1038 -3071 1039 -3069
rect 1045 -3065 1046 -3063
rect 1045 -3071 1046 -3069
rect 1052 -3065 1053 -3063
rect 1052 -3071 1053 -3069
rect 1062 -3065 1063 -3063
rect 1062 -3071 1063 -3069
rect 1066 -3065 1067 -3063
rect 1066 -3071 1067 -3069
rect 1073 -3065 1074 -3063
rect 1073 -3071 1074 -3069
rect 1080 -3065 1081 -3063
rect 1080 -3071 1081 -3069
rect 1087 -3065 1088 -3063
rect 1090 -3065 1091 -3063
rect 1087 -3071 1088 -3069
rect 1094 -3065 1095 -3063
rect 1094 -3071 1095 -3069
rect 1101 -3065 1102 -3063
rect 1101 -3071 1102 -3069
rect 1108 -3065 1109 -3063
rect 1108 -3071 1109 -3069
rect 1115 -3065 1116 -3063
rect 1115 -3071 1116 -3069
rect 1122 -3065 1123 -3063
rect 1122 -3071 1123 -3069
rect 1129 -3065 1130 -3063
rect 1129 -3071 1130 -3069
rect 1136 -3065 1137 -3063
rect 1136 -3071 1137 -3069
rect 1143 -3065 1144 -3063
rect 1143 -3071 1144 -3069
rect 1150 -3065 1151 -3063
rect 1150 -3071 1151 -3069
rect 1157 -3065 1158 -3063
rect 1157 -3071 1158 -3069
rect 1164 -3065 1165 -3063
rect 1164 -3071 1165 -3069
rect 1171 -3065 1172 -3063
rect 1171 -3071 1172 -3069
rect 1178 -3065 1179 -3063
rect 1178 -3071 1179 -3069
rect 1185 -3065 1186 -3063
rect 1185 -3071 1186 -3069
rect 1192 -3065 1193 -3063
rect 1192 -3071 1193 -3069
rect 1199 -3065 1200 -3063
rect 1199 -3071 1200 -3069
rect 1206 -3065 1207 -3063
rect 1206 -3071 1207 -3069
rect 1213 -3065 1214 -3063
rect 1213 -3071 1214 -3069
rect 1220 -3065 1221 -3063
rect 1223 -3065 1224 -3063
rect 1220 -3071 1221 -3069
rect 1223 -3071 1224 -3069
rect 1227 -3065 1228 -3063
rect 1227 -3071 1228 -3069
rect 1234 -3065 1235 -3063
rect 1234 -3071 1235 -3069
rect 1241 -3065 1242 -3063
rect 1241 -3071 1242 -3069
rect 1248 -3065 1249 -3063
rect 1248 -3071 1249 -3069
rect 1255 -3065 1256 -3063
rect 1255 -3071 1256 -3069
rect 1262 -3065 1263 -3063
rect 1262 -3071 1263 -3069
rect 1269 -3065 1270 -3063
rect 1269 -3071 1270 -3069
rect 1276 -3065 1277 -3063
rect 1276 -3071 1277 -3069
rect 1283 -3065 1284 -3063
rect 1283 -3071 1284 -3069
rect 1286 -3071 1287 -3069
rect 1290 -3065 1291 -3063
rect 1290 -3071 1291 -3069
rect 1297 -3065 1298 -3063
rect 1297 -3071 1298 -3069
rect 1304 -3065 1305 -3063
rect 1304 -3071 1305 -3069
rect 1311 -3065 1312 -3063
rect 1311 -3071 1312 -3069
rect 1318 -3065 1319 -3063
rect 1318 -3071 1319 -3069
rect 1325 -3065 1326 -3063
rect 1325 -3071 1326 -3069
rect 1332 -3065 1333 -3063
rect 1332 -3071 1333 -3069
rect 1339 -3065 1340 -3063
rect 1339 -3071 1340 -3069
rect 1346 -3065 1347 -3063
rect 1346 -3071 1347 -3069
rect 1374 -3065 1375 -3063
rect 1374 -3071 1375 -3069
rect 1381 -3065 1382 -3063
rect 1381 -3071 1382 -3069
rect 1416 -3065 1417 -3063
rect 1416 -3071 1417 -3069
rect 1458 -3065 1459 -3063
rect 1458 -3071 1459 -3069
rect 1465 -3065 1466 -3063
rect 1465 -3071 1466 -3069
rect 1472 -3065 1473 -3063
rect 1472 -3071 1473 -3069
rect 79 -3154 80 -3152
rect 79 -3160 80 -3158
rect 86 -3154 87 -3152
rect 86 -3160 87 -3158
rect 93 -3154 94 -3152
rect 93 -3160 94 -3158
rect 100 -3154 101 -3152
rect 100 -3160 101 -3158
rect 107 -3154 108 -3152
rect 107 -3160 108 -3158
rect 114 -3154 115 -3152
rect 114 -3160 115 -3158
rect 121 -3154 122 -3152
rect 121 -3160 122 -3158
rect 128 -3154 129 -3152
rect 128 -3160 129 -3158
rect 135 -3154 136 -3152
rect 135 -3160 136 -3158
rect 142 -3154 143 -3152
rect 142 -3160 143 -3158
rect 149 -3154 150 -3152
rect 149 -3160 150 -3158
rect 156 -3154 157 -3152
rect 156 -3160 157 -3158
rect 163 -3154 164 -3152
rect 163 -3160 164 -3158
rect 170 -3154 171 -3152
rect 170 -3160 171 -3158
rect 177 -3154 178 -3152
rect 177 -3160 178 -3158
rect 187 -3154 188 -3152
rect 187 -3160 188 -3158
rect 191 -3154 192 -3152
rect 191 -3160 192 -3158
rect 198 -3154 199 -3152
rect 198 -3160 199 -3158
rect 205 -3154 206 -3152
rect 205 -3160 206 -3158
rect 215 -3154 216 -3152
rect 212 -3160 213 -3158
rect 215 -3160 216 -3158
rect 219 -3154 220 -3152
rect 222 -3154 223 -3152
rect 222 -3160 223 -3158
rect 226 -3154 227 -3152
rect 226 -3160 227 -3158
rect 233 -3154 234 -3152
rect 233 -3160 234 -3158
rect 240 -3154 241 -3152
rect 240 -3160 241 -3158
rect 247 -3154 248 -3152
rect 247 -3160 248 -3158
rect 254 -3154 255 -3152
rect 254 -3160 255 -3158
rect 261 -3154 262 -3152
rect 261 -3160 262 -3158
rect 268 -3154 269 -3152
rect 268 -3160 269 -3158
rect 275 -3154 276 -3152
rect 275 -3160 276 -3158
rect 282 -3154 283 -3152
rect 282 -3160 283 -3158
rect 289 -3154 290 -3152
rect 289 -3160 290 -3158
rect 296 -3154 297 -3152
rect 296 -3160 297 -3158
rect 303 -3154 304 -3152
rect 306 -3160 307 -3158
rect 310 -3154 311 -3152
rect 310 -3160 311 -3158
rect 317 -3154 318 -3152
rect 317 -3160 318 -3158
rect 324 -3154 325 -3152
rect 324 -3160 325 -3158
rect 331 -3154 332 -3152
rect 331 -3160 332 -3158
rect 338 -3154 339 -3152
rect 338 -3160 339 -3158
rect 345 -3154 346 -3152
rect 345 -3160 346 -3158
rect 352 -3154 353 -3152
rect 352 -3160 353 -3158
rect 359 -3154 360 -3152
rect 362 -3154 363 -3152
rect 359 -3160 360 -3158
rect 362 -3160 363 -3158
rect 366 -3154 367 -3152
rect 366 -3160 367 -3158
rect 373 -3154 374 -3152
rect 373 -3160 374 -3158
rect 380 -3154 381 -3152
rect 380 -3160 381 -3158
rect 387 -3154 388 -3152
rect 387 -3160 388 -3158
rect 394 -3154 395 -3152
rect 394 -3160 395 -3158
rect 401 -3154 402 -3152
rect 401 -3160 402 -3158
rect 408 -3154 409 -3152
rect 408 -3160 409 -3158
rect 415 -3154 416 -3152
rect 415 -3160 416 -3158
rect 422 -3154 423 -3152
rect 422 -3160 423 -3158
rect 432 -3160 433 -3158
rect 436 -3154 437 -3152
rect 436 -3160 437 -3158
rect 443 -3154 444 -3152
rect 443 -3160 444 -3158
rect 450 -3154 451 -3152
rect 450 -3160 451 -3158
rect 457 -3154 458 -3152
rect 457 -3160 458 -3158
rect 464 -3154 465 -3152
rect 464 -3160 465 -3158
rect 471 -3154 472 -3152
rect 471 -3160 472 -3158
rect 478 -3154 479 -3152
rect 478 -3160 479 -3158
rect 485 -3154 486 -3152
rect 485 -3160 486 -3158
rect 492 -3154 493 -3152
rect 492 -3160 493 -3158
rect 499 -3154 500 -3152
rect 499 -3160 500 -3158
rect 506 -3154 507 -3152
rect 506 -3160 507 -3158
rect 513 -3154 514 -3152
rect 513 -3160 514 -3158
rect 520 -3154 521 -3152
rect 527 -3154 528 -3152
rect 527 -3160 528 -3158
rect 534 -3154 535 -3152
rect 534 -3160 535 -3158
rect 541 -3154 542 -3152
rect 541 -3160 542 -3158
rect 548 -3154 549 -3152
rect 548 -3160 549 -3158
rect 555 -3154 556 -3152
rect 555 -3160 556 -3158
rect 562 -3154 563 -3152
rect 562 -3160 563 -3158
rect 569 -3154 570 -3152
rect 569 -3160 570 -3158
rect 576 -3154 577 -3152
rect 579 -3154 580 -3152
rect 579 -3160 580 -3158
rect 583 -3154 584 -3152
rect 583 -3160 584 -3158
rect 590 -3154 591 -3152
rect 590 -3160 591 -3158
rect 597 -3154 598 -3152
rect 597 -3160 598 -3158
rect 604 -3154 605 -3152
rect 607 -3154 608 -3152
rect 604 -3160 605 -3158
rect 611 -3154 612 -3152
rect 611 -3160 612 -3158
rect 621 -3154 622 -3152
rect 618 -3160 619 -3158
rect 625 -3154 626 -3152
rect 625 -3160 626 -3158
rect 632 -3154 633 -3152
rect 635 -3154 636 -3152
rect 632 -3160 633 -3158
rect 639 -3154 640 -3152
rect 639 -3160 640 -3158
rect 646 -3154 647 -3152
rect 646 -3160 647 -3158
rect 653 -3154 654 -3152
rect 656 -3154 657 -3152
rect 656 -3160 657 -3158
rect 660 -3154 661 -3152
rect 660 -3160 661 -3158
rect 663 -3160 664 -3158
rect 667 -3154 668 -3152
rect 667 -3160 668 -3158
rect 674 -3154 675 -3152
rect 674 -3160 675 -3158
rect 681 -3154 682 -3152
rect 681 -3160 682 -3158
rect 688 -3160 689 -3158
rect 695 -3154 696 -3152
rect 695 -3160 696 -3158
rect 705 -3154 706 -3152
rect 702 -3160 703 -3158
rect 705 -3160 706 -3158
rect 709 -3154 710 -3152
rect 709 -3160 710 -3158
rect 716 -3154 717 -3152
rect 716 -3160 717 -3158
rect 723 -3154 724 -3152
rect 723 -3160 724 -3158
rect 730 -3154 731 -3152
rect 730 -3160 731 -3158
rect 733 -3160 734 -3158
rect 737 -3154 738 -3152
rect 737 -3160 738 -3158
rect 744 -3154 745 -3152
rect 744 -3160 745 -3158
rect 751 -3154 752 -3152
rect 751 -3160 752 -3158
rect 758 -3154 759 -3152
rect 758 -3160 759 -3158
rect 765 -3154 766 -3152
rect 765 -3160 766 -3158
rect 772 -3154 773 -3152
rect 775 -3154 776 -3152
rect 772 -3160 773 -3158
rect 775 -3160 776 -3158
rect 779 -3154 780 -3152
rect 782 -3154 783 -3152
rect 779 -3160 780 -3158
rect 782 -3160 783 -3158
rect 786 -3154 787 -3152
rect 786 -3160 787 -3158
rect 793 -3154 794 -3152
rect 793 -3160 794 -3158
rect 800 -3154 801 -3152
rect 800 -3160 801 -3158
rect 807 -3154 808 -3152
rect 807 -3160 808 -3158
rect 814 -3154 815 -3152
rect 814 -3160 815 -3158
rect 821 -3154 822 -3152
rect 821 -3160 822 -3158
rect 828 -3154 829 -3152
rect 828 -3160 829 -3158
rect 835 -3154 836 -3152
rect 835 -3160 836 -3158
rect 842 -3154 843 -3152
rect 845 -3154 846 -3152
rect 845 -3160 846 -3158
rect 849 -3154 850 -3152
rect 849 -3160 850 -3158
rect 856 -3154 857 -3152
rect 856 -3160 857 -3158
rect 863 -3154 864 -3152
rect 863 -3160 864 -3158
rect 870 -3154 871 -3152
rect 870 -3160 871 -3158
rect 877 -3154 878 -3152
rect 880 -3154 881 -3152
rect 880 -3160 881 -3158
rect 884 -3154 885 -3152
rect 884 -3160 885 -3158
rect 891 -3154 892 -3152
rect 891 -3160 892 -3158
rect 898 -3154 899 -3152
rect 898 -3160 899 -3158
rect 905 -3154 906 -3152
rect 905 -3160 906 -3158
rect 912 -3154 913 -3152
rect 912 -3160 913 -3158
rect 919 -3154 920 -3152
rect 919 -3160 920 -3158
rect 926 -3154 927 -3152
rect 926 -3160 927 -3158
rect 933 -3154 934 -3152
rect 933 -3160 934 -3158
rect 940 -3154 941 -3152
rect 940 -3160 941 -3158
rect 947 -3154 948 -3152
rect 947 -3160 948 -3158
rect 954 -3154 955 -3152
rect 954 -3160 955 -3158
rect 961 -3154 962 -3152
rect 964 -3154 965 -3152
rect 961 -3160 962 -3158
rect 964 -3160 965 -3158
rect 968 -3154 969 -3152
rect 968 -3160 969 -3158
rect 975 -3154 976 -3152
rect 975 -3160 976 -3158
rect 982 -3154 983 -3152
rect 982 -3160 983 -3158
rect 989 -3154 990 -3152
rect 989 -3160 990 -3158
rect 996 -3160 997 -3158
rect 999 -3160 1000 -3158
rect 1003 -3154 1004 -3152
rect 1003 -3160 1004 -3158
rect 1010 -3154 1011 -3152
rect 1010 -3160 1011 -3158
rect 1017 -3154 1018 -3152
rect 1017 -3160 1018 -3158
rect 1024 -3154 1025 -3152
rect 1024 -3160 1025 -3158
rect 1031 -3154 1032 -3152
rect 1031 -3160 1032 -3158
rect 1038 -3154 1039 -3152
rect 1038 -3160 1039 -3158
rect 1045 -3154 1046 -3152
rect 1045 -3160 1046 -3158
rect 1052 -3154 1053 -3152
rect 1052 -3160 1053 -3158
rect 1059 -3154 1060 -3152
rect 1059 -3160 1060 -3158
rect 1066 -3154 1067 -3152
rect 1066 -3160 1067 -3158
rect 1073 -3154 1074 -3152
rect 1073 -3160 1074 -3158
rect 1080 -3154 1081 -3152
rect 1080 -3160 1081 -3158
rect 1090 -3154 1091 -3152
rect 1094 -3154 1095 -3152
rect 1094 -3160 1095 -3158
rect 1097 -3160 1098 -3158
rect 1101 -3154 1102 -3152
rect 1101 -3160 1102 -3158
rect 1108 -3154 1109 -3152
rect 1108 -3160 1109 -3158
rect 1115 -3154 1116 -3152
rect 1115 -3160 1116 -3158
rect 1122 -3154 1123 -3152
rect 1122 -3160 1123 -3158
rect 1129 -3154 1130 -3152
rect 1129 -3160 1130 -3158
rect 1136 -3154 1137 -3152
rect 1136 -3160 1137 -3158
rect 1143 -3154 1144 -3152
rect 1143 -3160 1144 -3158
rect 1150 -3154 1151 -3152
rect 1150 -3160 1151 -3158
rect 1157 -3154 1158 -3152
rect 1157 -3160 1158 -3158
rect 1164 -3154 1165 -3152
rect 1164 -3160 1165 -3158
rect 1171 -3154 1172 -3152
rect 1171 -3160 1172 -3158
rect 1178 -3154 1179 -3152
rect 1178 -3160 1179 -3158
rect 1188 -3154 1189 -3152
rect 1185 -3160 1186 -3158
rect 1188 -3160 1189 -3158
rect 1192 -3154 1193 -3152
rect 1192 -3160 1193 -3158
rect 1199 -3154 1200 -3152
rect 1199 -3160 1200 -3158
rect 1206 -3154 1207 -3152
rect 1206 -3160 1207 -3158
rect 1213 -3154 1214 -3152
rect 1213 -3160 1214 -3158
rect 1220 -3154 1221 -3152
rect 1220 -3160 1221 -3158
rect 1227 -3154 1228 -3152
rect 1230 -3154 1231 -3152
rect 1227 -3160 1228 -3158
rect 1237 -3160 1238 -3158
rect 1241 -3154 1242 -3152
rect 1241 -3160 1242 -3158
rect 1244 -3160 1245 -3158
rect 1262 -3154 1263 -3152
rect 1262 -3160 1263 -3158
rect 1276 -3154 1277 -3152
rect 1276 -3160 1277 -3158
rect 1290 -3154 1291 -3152
rect 1293 -3154 1294 -3152
rect 1293 -3160 1294 -3158
rect 1346 -3154 1347 -3152
rect 1346 -3160 1347 -3158
rect 1353 -3154 1354 -3152
rect 1353 -3160 1354 -3158
rect 1367 -3154 1368 -3152
rect 1367 -3160 1368 -3158
rect 1409 -3154 1410 -3152
rect 1409 -3160 1410 -3158
rect 1451 -3154 1452 -3152
rect 1451 -3160 1452 -3158
rect 1458 -3154 1459 -3152
rect 1458 -3160 1459 -3158
rect 1465 -3154 1466 -3152
rect 1465 -3160 1466 -3158
rect 58 -3215 59 -3213
rect 58 -3221 59 -3219
rect 65 -3215 66 -3213
rect 65 -3221 66 -3219
rect 72 -3215 73 -3213
rect 72 -3221 73 -3219
rect 79 -3215 80 -3213
rect 79 -3221 80 -3219
rect 86 -3215 87 -3213
rect 86 -3221 87 -3219
rect 93 -3215 94 -3213
rect 93 -3221 94 -3219
rect 100 -3215 101 -3213
rect 100 -3221 101 -3219
rect 107 -3215 108 -3213
rect 107 -3221 108 -3219
rect 114 -3221 115 -3219
rect 117 -3221 118 -3219
rect 121 -3215 122 -3213
rect 121 -3221 122 -3219
rect 128 -3215 129 -3213
rect 131 -3215 132 -3213
rect 128 -3221 129 -3219
rect 131 -3221 132 -3219
rect 135 -3215 136 -3213
rect 135 -3221 136 -3219
rect 142 -3215 143 -3213
rect 145 -3215 146 -3213
rect 152 -3215 153 -3213
rect 149 -3221 150 -3219
rect 152 -3221 153 -3219
rect 156 -3215 157 -3213
rect 156 -3221 157 -3219
rect 163 -3215 164 -3213
rect 163 -3221 164 -3219
rect 173 -3215 174 -3213
rect 173 -3221 174 -3219
rect 180 -3215 181 -3213
rect 180 -3221 181 -3219
rect 184 -3215 185 -3213
rect 184 -3221 185 -3219
rect 191 -3215 192 -3213
rect 194 -3215 195 -3213
rect 191 -3221 192 -3219
rect 198 -3215 199 -3213
rect 201 -3215 202 -3213
rect 198 -3221 199 -3219
rect 201 -3221 202 -3219
rect 205 -3215 206 -3213
rect 208 -3215 209 -3213
rect 208 -3221 209 -3219
rect 212 -3215 213 -3213
rect 212 -3221 213 -3219
rect 219 -3215 220 -3213
rect 219 -3221 220 -3219
rect 226 -3215 227 -3213
rect 226 -3221 227 -3219
rect 233 -3215 234 -3213
rect 233 -3221 234 -3219
rect 240 -3215 241 -3213
rect 240 -3221 241 -3219
rect 247 -3215 248 -3213
rect 250 -3215 251 -3213
rect 247 -3221 248 -3219
rect 250 -3221 251 -3219
rect 254 -3215 255 -3213
rect 261 -3215 262 -3213
rect 264 -3215 265 -3213
rect 261 -3221 262 -3219
rect 264 -3221 265 -3219
rect 268 -3215 269 -3213
rect 268 -3221 269 -3219
rect 275 -3215 276 -3213
rect 275 -3221 276 -3219
rect 282 -3215 283 -3213
rect 282 -3221 283 -3219
rect 289 -3215 290 -3213
rect 289 -3221 290 -3219
rect 296 -3215 297 -3213
rect 296 -3221 297 -3219
rect 303 -3215 304 -3213
rect 303 -3221 304 -3219
rect 310 -3215 311 -3213
rect 310 -3221 311 -3219
rect 317 -3215 318 -3213
rect 317 -3221 318 -3219
rect 324 -3215 325 -3213
rect 327 -3215 328 -3213
rect 324 -3221 325 -3219
rect 331 -3215 332 -3213
rect 331 -3221 332 -3219
rect 338 -3215 339 -3213
rect 338 -3221 339 -3219
rect 345 -3215 346 -3213
rect 352 -3215 353 -3213
rect 352 -3221 353 -3219
rect 359 -3215 360 -3213
rect 359 -3221 360 -3219
rect 366 -3215 367 -3213
rect 366 -3221 367 -3219
rect 373 -3215 374 -3213
rect 373 -3221 374 -3219
rect 380 -3215 381 -3213
rect 380 -3221 381 -3219
rect 387 -3215 388 -3213
rect 387 -3221 388 -3219
rect 394 -3215 395 -3213
rect 394 -3221 395 -3219
rect 401 -3215 402 -3213
rect 401 -3221 402 -3219
rect 408 -3215 409 -3213
rect 408 -3221 409 -3219
rect 415 -3215 416 -3213
rect 415 -3221 416 -3219
rect 422 -3215 423 -3213
rect 422 -3221 423 -3219
rect 429 -3215 430 -3213
rect 429 -3221 430 -3219
rect 436 -3215 437 -3213
rect 436 -3221 437 -3219
rect 443 -3215 444 -3213
rect 443 -3221 444 -3219
rect 450 -3215 451 -3213
rect 450 -3221 451 -3219
rect 457 -3215 458 -3213
rect 457 -3221 458 -3219
rect 464 -3215 465 -3213
rect 464 -3221 465 -3219
rect 471 -3215 472 -3213
rect 471 -3221 472 -3219
rect 478 -3215 479 -3213
rect 478 -3221 479 -3219
rect 485 -3215 486 -3213
rect 485 -3221 486 -3219
rect 492 -3215 493 -3213
rect 492 -3221 493 -3219
rect 499 -3215 500 -3213
rect 499 -3221 500 -3219
rect 506 -3215 507 -3213
rect 506 -3221 507 -3219
rect 513 -3215 514 -3213
rect 513 -3221 514 -3219
rect 520 -3221 521 -3219
rect 527 -3215 528 -3213
rect 527 -3221 528 -3219
rect 534 -3215 535 -3213
rect 534 -3221 535 -3219
rect 537 -3221 538 -3219
rect 541 -3215 542 -3213
rect 541 -3221 542 -3219
rect 548 -3215 549 -3213
rect 548 -3221 549 -3219
rect 555 -3215 556 -3213
rect 555 -3221 556 -3219
rect 558 -3221 559 -3219
rect 562 -3215 563 -3213
rect 562 -3221 563 -3219
rect 569 -3215 570 -3213
rect 569 -3221 570 -3219
rect 576 -3221 577 -3219
rect 579 -3221 580 -3219
rect 583 -3215 584 -3213
rect 583 -3221 584 -3219
rect 590 -3215 591 -3213
rect 590 -3221 591 -3219
rect 597 -3215 598 -3213
rect 597 -3221 598 -3219
rect 604 -3215 605 -3213
rect 607 -3215 608 -3213
rect 604 -3221 605 -3219
rect 607 -3221 608 -3219
rect 611 -3215 612 -3213
rect 611 -3221 612 -3219
rect 618 -3215 619 -3213
rect 618 -3221 619 -3219
rect 625 -3215 626 -3213
rect 628 -3221 629 -3219
rect 632 -3215 633 -3213
rect 635 -3215 636 -3213
rect 632 -3221 633 -3219
rect 635 -3221 636 -3219
rect 639 -3215 640 -3213
rect 639 -3221 640 -3219
rect 646 -3215 647 -3213
rect 646 -3221 647 -3219
rect 653 -3215 654 -3213
rect 653 -3221 654 -3219
rect 660 -3215 661 -3213
rect 660 -3221 661 -3219
rect 663 -3221 664 -3219
rect 667 -3215 668 -3213
rect 667 -3221 668 -3219
rect 674 -3215 675 -3213
rect 674 -3221 675 -3219
rect 681 -3215 682 -3213
rect 681 -3221 682 -3219
rect 688 -3215 689 -3213
rect 688 -3221 689 -3219
rect 695 -3215 696 -3213
rect 695 -3221 696 -3219
rect 702 -3215 703 -3213
rect 702 -3221 703 -3219
rect 709 -3215 710 -3213
rect 709 -3221 710 -3219
rect 716 -3215 717 -3213
rect 716 -3221 717 -3219
rect 723 -3215 724 -3213
rect 723 -3221 724 -3219
rect 730 -3215 731 -3213
rect 730 -3221 731 -3219
rect 737 -3215 738 -3213
rect 737 -3221 738 -3219
rect 744 -3215 745 -3213
rect 744 -3221 745 -3219
rect 751 -3215 752 -3213
rect 751 -3221 752 -3219
rect 758 -3215 759 -3213
rect 761 -3215 762 -3213
rect 758 -3221 759 -3219
rect 765 -3215 766 -3213
rect 765 -3221 766 -3219
rect 772 -3215 773 -3213
rect 772 -3221 773 -3219
rect 779 -3215 780 -3213
rect 779 -3221 780 -3219
rect 786 -3215 787 -3213
rect 786 -3221 787 -3219
rect 793 -3215 794 -3213
rect 793 -3221 794 -3219
rect 800 -3215 801 -3213
rect 800 -3221 801 -3219
rect 807 -3215 808 -3213
rect 807 -3221 808 -3219
rect 814 -3215 815 -3213
rect 814 -3221 815 -3219
rect 821 -3215 822 -3213
rect 821 -3221 822 -3219
rect 828 -3215 829 -3213
rect 828 -3221 829 -3219
rect 835 -3215 836 -3213
rect 835 -3221 836 -3219
rect 842 -3215 843 -3213
rect 842 -3221 843 -3219
rect 849 -3215 850 -3213
rect 849 -3221 850 -3219
rect 856 -3215 857 -3213
rect 856 -3221 857 -3219
rect 863 -3215 864 -3213
rect 866 -3215 867 -3213
rect 863 -3221 864 -3219
rect 866 -3221 867 -3219
rect 870 -3215 871 -3213
rect 870 -3221 871 -3219
rect 877 -3215 878 -3213
rect 877 -3221 878 -3219
rect 884 -3215 885 -3213
rect 884 -3221 885 -3219
rect 891 -3215 892 -3213
rect 891 -3221 892 -3219
rect 898 -3215 899 -3213
rect 898 -3221 899 -3219
rect 905 -3215 906 -3213
rect 905 -3221 906 -3219
rect 912 -3215 913 -3213
rect 912 -3221 913 -3219
rect 919 -3215 920 -3213
rect 919 -3221 920 -3219
rect 926 -3215 927 -3213
rect 926 -3221 927 -3219
rect 933 -3215 934 -3213
rect 933 -3221 934 -3219
rect 940 -3215 941 -3213
rect 940 -3221 941 -3219
rect 947 -3215 948 -3213
rect 947 -3221 948 -3219
rect 954 -3215 955 -3213
rect 954 -3221 955 -3219
rect 961 -3215 962 -3213
rect 961 -3221 962 -3219
rect 968 -3215 969 -3213
rect 968 -3221 969 -3219
rect 975 -3215 976 -3213
rect 975 -3221 976 -3219
rect 982 -3215 983 -3213
rect 985 -3215 986 -3213
rect 982 -3221 983 -3219
rect 985 -3221 986 -3219
rect 989 -3215 990 -3213
rect 989 -3221 990 -3219
rect 996 -3215 997 -3213
rect 996 -3221 997 -3219
rect 1003 -3215 1004 -3213
rect 1006 -3215 1007 -3213
rect 1003 -3221 1004 -3219
rect 1010 -3215 1011 -3213
rect 1010 -3221 1011 -3219
rect 1017 -3215 1018 -3213
rect 1017 -3221 1018 -3219
rect 1024 -3215 1025 -3213
rect 1024 -3221 1025 -3219
rect 1031 -3215 1032 -3213
rect 1031 -3221 1032 -3219
rect 1038 -3215 1039 -3213
rect 1038 -3221 1039 -3219
rect 1045 -3215 1046 -3213
rect 1045 -3221 1046 -3219
rect 1052 -3215 1053 -3213
rect 1052 -3221 1053 -3219
rect 1059 -3215 1060 -3213
rect 1059 -3221 1060 -3219
rect 1062 -3221 1063 -3219
rect 1073 -3215 1074 -3213
rect 1073 -3221 1074 -3219
rect 1080 -3215 1081 -3213
rect 1080 -3221 1081 -3219
rect 1087 -3215 1088 -3213
rect 1087 -3221 1088 -3219
rect 1094 -3215 1095 -3213
rect 1097 -3215 1098 -3213
rect 1094 -3221 1095 -3219
rect 1101 -3215 1102 -3213
rect 1101 -3221 1102 -3219
rect 1111 -3215 1112 -3213
rect 1108 -3221 1109 -3219
rect 1111 -3221 1112 -3219
rect 1115 -3215 1116 -3213
rect 1115 -3221 1116 -3219
rect 1122 -3215 1123 -3213
rect 1122 -3221 1123 -3219
rect 1129 -3215 1130 -3213
rect 1129 -3221 1130 -3219
rect 1136 -3215 1137 -3213
rect 1136 -3221 1137 -3219
rect 1143 -3215 1144 -3213
rect 1143 -3221 1144 -3219
rect 1150 -3215 1151 -3213
rect 1150 -3221 1151 -3219
rect 1157 -3215 1158 -3213
rect 1157 -3221 1158 -3219
rect 1164 -3215 1165 -3213
rect 1167 -3215 1168 -3213
rect 1164 -3221 1165 -3219
rect 1167 -3221 1168 -3219
rect 1171 -3215 1172 -3213
rect 1171 -3221 1172 -3219
rect 1185 -3215 1186 -3213
rect 1185 -3221 1186 -3219
rect 1192 -3215 1193 -3213
rect 1192 -3221 1193 -3219
rect 1199 -3215 1200 -3213
rect 1199 -3221 1200 -3219
rect 1206 -3215 1207 -3213
rect 1206 -3221 1207 -3219
rect 1213 -3215 1214 -3213
rect 1213 -3221 1214 -3219
rect 1234 -3215 1235 -3213
rect 1234 -3221 1235 -3219
rect 1332 -3215 1333 -3213
rect 1332 -3221 1333 -3219
rect 1360 -3215 1361 -3213
rect 1360 -3221 1361 -3219
rect 1367 -3215 1368 -3213
rect 1367 -3221 1368 -3219
rect 1409 -3215 1410 -3213
rect 1409 -3221 1410 -3219
rect 1451 -3215 1452 -3213
rect 1451 -3221 1452 -3219
rect 1454 -3221 1455 -3219
rect 1458 -3215 1459 -3213
rect 1458 -3221 1459 -3219
rect 1465 -3215 1466 -3213
rect 1465 -3221 1466 -3219
rect 156 -3270 157 -3268
rect 156 -3276 157 -3274
rect 163 -3270 164 -3268
rect 163 -3276 164 -3274
rect 170 -3270 171 -3268
rect 170 -3276 171 -3274
rect 177 -3270 178 -3268
rect 177 -3276 178 -3274
rect 187 -3270 188 -3268
rect 184 -3276 185 -3274
rect 187 -3276 188 -3274
rect 191 -3270 192 -3268
rect 191 -3276 192 -3274
rect 198 -3270 199 -3268
rect 198 -3276 199 -3274
rect 208 -3270 209 -3268
rect 208 -3276 209 -3274
rect 212 -3270 213 -3268
rect 212 -3276 213 -3274
rect 219 -3270 220 -3268
rect 219 -3276 220 -3274
rect 226 -3270 227 -3268
rect 226 -3276 227 -3274
rect 233 -3270 234 -3268
rect 233 -3276 234 -3274
rect 240 -3270 241 -3268
rect 243 -3270 244 -3268
rect 243 -3276 244 -3274
rect 247 -3270 248 -3268
rect 250 -3270 251 -3268
rect 254 -3276 255 -3274
rect 261 -3270 262 -3268
rect 264 -3270 265 -3268
rect 268 -3270 269 -3268
rect 268 -3276 269 -3274
rect 275 -3270 276 -3268
rect 275 -3276 276 -3274
rect 282 -3270 283 -3268
rect 282 -3276 283 -3274
rect 289 -3270 290 -3268
rect 289 -3276 290 -3274
rect 296 -3270 297 -3268
rect 296 -3276 297 -3274
rect 303 -3270 304 -3268
rect 303 -3276 304 -3274
rect 310 -3270 311 -3268
rect 310 -3276 311 -3274
rect 317 -3270 318 -3268
rect 317 -3276 318 -3274
rect 324 -3270 325 -3268
rect 324 -3276 325 -3274
rect 331 -3270 332 -3268
rect 331 -3276 332 -3274
rect 338 -3270 339 -3268
rect 338 -3276 339 -3274
rect 345 -3276 346 -3274
rect 352 -3270 353 -3268
rect 352 -3276 353 -3274
rect 359 -3270 360 -3268
rect 359 -3276 360 -3274
rect 366 -3270 367 -3268
rect 366 -3276 367 -3274
rect 373 -3270 374 -3268
rect 373 -3276 374 -3274
rect 380 -3270 381 -3268
rect 380 -3276 381 -3274
rect 387 -3270 388 -3268
rect 387 -3276 388 -3274
rect 394 -3270 395 -3268
rect 397 -3270 398 -3268
rect 394 -3276 395 -3274
rect 401 -3270 402 -3268
rect 404 -3270 405 -3268
rect 401 -3276 402 -3274
rect 408 -3270 409 -3268
rect 408 -3276 409 -3274
rect 415 -3270 416 -3268
rect 415 -3276 416 -3274
rect 422 -3270 423 -3268
rect 422 -3276 423 -3274
rect 429 -3270 430 -3268
rect 429 -3276 430 -3274
rect 436 -3270 437 -3268
rect 436 -3276 437 -3274
rect 443 -3270 444 -3268
rect 443 -3276 444 -3274
rect 450 -3270 451 -3268
rect 450 -3276 451 -3274
rect 457 -3270 458 -3268
rect 457 -3276 458 -3274
rect 464 -3270 465 -3268
rect 464 -3276 465 -3274
rect 471 -3270 472 -3268
rect 474 -3270 475 -3268
rect 474 -3276 475 -3274
rect 478 -3270 479 -3268
rect 478 -3276 479 -3274
rect 485 -3270 486 -3268
rect 488 -3270 489 -3268
rect 485 -3276 486 -3274
rect 488 -3276 489 -3274
rect 492 -3270 493 -3268
rect 492 -3276 493 -3274
rect 499 -3270 500 -3268
rect 499 -3276 500 -3274
rect 506 -3270 507 -3268
rect 506 -3276 507 -3274
rect 513 -3270 514 -3268
rect 513 -3276 514 -3274
rect 520 -3270 521 -3268
rect 520 -3276 521 -3274
rect 527 -3270 528 -3268
rect 527 -3276 528 -3274
rect 534 -3270 535 -3268
rect 537 -3270 538 -3268
rect 534 -3276 535 -3274
rect 541 -3270 542 -3268
rect 541 -3276 542 -3274
rect 548 -3270 549 -3268
rect 548 -3276 549 -3274
rect 555 -3270 556 -3268
rect 555 -3276 556 -3274
rect 562 -3270 563 -3268
rect 562 -3276 563 -3274
rect 569 -3270 570 -3268
rect 569 -3276 570 -3274
rect 576 -3270 577 -3268
rect 576 -3276 577 -3274
rect 583 -3270 584 -3268
rect 583 -3276 584 -3274
rect 590 -3276 591 -3274
rect 593 -3276 594 -3274
rect 597 -3270 598 -3268
rect 597 -3276 598 -3274
rect 604 -3270 605 -3268
rect 604 -3276 605 -3274
rect 611 -3270 612 -3268
rect 611 -3276 612 -3274
rect 618 -3270 619 -3268
rect 618 -3276 619 -3274
rect 625 -3270 626 -3268
rect 625 -3276 626 -3274
rect 632 -3270 633 -3268
rect 635 -3270 636 -3268
rect 632 -3276 633 -3274
rect 635 -3276 636 -3274
rect 639 -3270 640 -3268
rect 639 -3276 640 -3274
rect 646 -3270 647 -3268
rect 646 -3276 647 -3274
rect 653 -3270 654 -3268
rect 653 -3276 654 -3274
rect 660 -3270 661 -3268
rect 660 -3276 661 -3274
rect 667 -3270 668 -3268
rect 667 -3276 668 -3274
rect 674 -3270 675 -3268
rect 674 -3276 675 -3274
rect 681 -3270 682 -3268
rect 681 -3276 682 -3274
rect 688 -3270 689 -3268
rect 688 -3276 689 -3274
rect 695 -3270 696 -3268
rect 695 -3276 696 -3274
rect 702 -3270 703 -3268
rect 702 -3276 703 -3274
rect 709 -3270 710 -3268
rect 709 -3276 710 -3274
rect 716 -3270 717 -3268
rect 716 -3276 717 -3274
rect 726 -3270 727 -3268
rect 723 -3276 724 -3274
rect 733 -3270 734 -3268
rect 730 -3276 731 -3274
rect 737 -3270 738 -3268
rect 737 -3276 738 -3274
rect 744 -3270 745 -3268
rect 744 -3276 745 -3274
rect 751 -3270 752 -3268
rect 751 -3276 752 -3274
rect 758 -3270 759 -3268
rect 758 -3276 759 -3274
rect 765 -3270 766 -3268
rect 765 -3276 766 -3274
rect 772 -3270 773 -3268
rect 772 -3276 773 -3274
rect 782 -3270 783 -3268
rect 779 -3276 780 -3274
rect 782 -3276 783 -3274
rect 786 -3270 787 -3268
rect 786 -3276 787 -3274
rect 793 -3270 794 -3268
rect 793 -3276 794 -3274
rect 800 -3270 801 -3268
rect 800 -3276 801 -3274
rect 807 -3270 808 -3268
rect 807 -3276 808 -3274
rect 814 -3270 815 -3268
rect 814 -3276 815 -3274
rect 821 -3270 822 -3268
rect 821 -3276 822 -3274
rect 828 -3270 829 -3268
rect 828 -3276 829 -3274
rect 842 -3270 843 -3268
rect 842 -3276 843 -3274
rect 870 -3270 871 -3268
rect 870 -3276 871 -3274
rect 877 -3270 878 -3268
rect 880 -3270 881 -3268
rect 877 -3276 878 -3274
rect 880 -3276 881 -3274
rect 884 -3270 885 -3268
rect 884 -3276 885 -3274
rect 891 -3270 892 -3268
rect 891 -3276 892 -3274
rect 898 -3270 899 -3268
rect 898 -3276 899 -3274
rect 905 -3270 906 -3268
rect 905 -3276 906 -3274
rect 912 -3270 913 -3268
rect 912 -3276 913 -3274
rect 919 -3270 920 -3268
rect 919 -3276 920 -3274
rect 926 -3270 927 -3268
rect 926 -3276 927 -3274
rect 933 -3270 934 -3268
rect 933 -3276 934 -3274
rect 940 -3270 941 -3268
rect 940 -3276 941 -3274
rect 947 -3270 948 -3268
rect 947 -3276 948 -3274
rect 954 -3270 955 -3268
rect 954 -3276 955 -3274
rect 961 -3270 962 -3268
rect 961 -3276 962 -3274
rect 982 -3270 983 -3268
rect 982 -3276 983 -3274
rect 992 -3270 993 -3268
rect 992 -3276 993 -3274
rect 996 -3270 997 -3268
rect 996 -3276 997 -3274
rect 1003 -3270 1004 -3268
rect 1003 -3276 1004 -3274
rect 1066 -3270 1067 -3268
rect 1066 -3276 1067 -3274
rect 1073 -3270 1074 -3268
rect 1073 -3276 1074 -3274
rect 1080 -3270 1081 -3268
rect 1080 -3276 1081 -3274
rect 1094 -3270 1095 -3268
rect 1094 -3276 1095 -3274
rect 1101 -3270 1102 -3268
rect 1101 -3276 1102 -3274
rect 1108 -3270 1109 -3268
rect 1108 -3276 1109 -3274
rect 1122 -3270 1123 -3268
rect 1125 -3270 1126 -3268
rect 1122 -3276 1123 -3274
rect 1125 -3276 1126 -3274
rect 1129 -3270 1130 -3268
rect 1129 -3276 1130 -3274
rect 1136 -3270 1137 -3268
rect 1136 -3276 1137 -3274
rect 1143 -3270 1144 -3268
rect 1143 -3276 1144 -3274
rect 1150 -3270 1151 -3268
rect 1150 -3276 1151 -3274
rect 1160 -3270 1161 -3268
rect 1157 -3276 1158 -3274
rect 1164 -3270 1165 -3268
rect 1164 -3276 1165 -3274
rect 1171 -3270 1172 -3268
rect 1171 -3276 1172 -3274
rect 1185 -3270 1186 -3268
rect 1188 -3270 1189 -3268
rect 1185 -3276 1186 -3274
rect 1206 -3270 1207 -3268
rect 1206 -3276 1207 -3274
rect 1216 -3270 1217 -3268
rect 1216 -3276 1217 -3274
rect 1220 -3270 1221 -3268
rect 1220 -3276 1221 -3274
rect 1234 -3270 1235 -3268
rect 1251 -3270 1252 -3268
rect 1251 -3276 1252 -3274
rect 1290 -3270 1291 -3268
rect 1290 -3276 1291 -3274
rect 1325 -3270 1326 -3268
rect 1328 -3270 1329 -3268
rect 1360 -3270 1361 -3268
rect 1360 -3276 1361 -3274
rect 1367 -3270 1368 -3268
rect 1367 -3276 1368 -3274
rect 1409 -3270 1410 -3268
rect 1409 -3276 1410 -3274
rect 1451 -3270 1452 -3268
rect 1454 -3270 1455 -3268
rect 1451 -3276 1452 -3274
rect 1458 -3270 1459 -3268
rect 1458 -3276 1459 -3274
rect 1461 -3276 1462 -3274
rect 1465 -3270 1466 -3268
rect 1465 -3276 1466 -3274
rect 177 -3333 178 -3331
rect 177 -3339 178 -3337
rect 184 -3333 185 -3331
rect 184 -3339 185 -3337
rect 191 -3333 192 -3331
rect 191 -3339 192 -3337
rect 198 -3333 199 -3331
rect 198 -3339 199 -3337
rect 205 -3333 206 -3331
rect 205 -3339 206 -3337
rect 212 -3333 213 -3331
rect 212 -3339 213 -3337
rect 219 -3333 220 -3331
rect 219 -3339 220 -3337
rect 226 -3333 227 -3331
rect 229 -3333 230 -3331
rect 233 -3333 234 -3331
rect 240 -3333 241 -3331
rect 240 -3339 241 -3337
rect 247 -3333 248 -3331
rect 247 -3339 248 -3337
rect 254 -3333 255 -3331
rect 254 -3339 255 -3337
rect 261 -3339 262 -3337
rect 264 -3339 265 -3337
rect 268 -3333 269 -3331
rect 268 -3339 269 -3337
rect 275 -3333 276 -3331
rect 275 -3339 276 -3337
rect 282 -3333 283 -3331
rect 282 -3339 283 -3337
rect 289 -3333 290 -3331
rect 289 -3339 290 -3337
rect 296 -3333 297 -3331
rect 296 -3339 297 -3337
rect 303 -3333 304 -3331
rect 303 -3339 304 -3337
rect 306 -3339 307 -3337
rect 310 -3333 311 -3331
rect 310 -3339 311 -3337
rect 317 -3333 318 -3331
rect 317 -3339 318 -3337
rect 324 -3333 325 -3331
rect 324 -3339 325 -3337
rect 331 -3333 332 -3331
rect 331 -3339 332 -3337
rect 338 -3333 339 -3331
rect 338 -3339 339 -3337
rect 345 -3333 346 -3331
rect 345 -3339 346 -3337
rect 352 -3333 353 -3331
rect 352 -3339 353 -3337
rect 359 -3333 360 -3331
rect 359 -3339 360 -3337
rect 366 -3333 367 -3331
rect 366 -3339 367 -3337
rect 373 -3333 374 -3331
rect 373 -3339 374 -3337
rect 380 -3333 381 -3331
rect 383 -3333 384 -3331
rect 383 -3339 384 -3337
rect 387 -3333 388 -3331
rect 387 -3339 388 -3337
rect 394 -3333 395 -3331
rect 394 -3339 395 -3337
rect 401 -3333 402 -3331
rect 401 -3339 402 -3337
rect 408 -3333 409 -3331
rect 411 -3333 412 -3331
rect 408 -3339 409 -3337
rect 411 -3339 412 -3337
rect 415 -3333 416 -3331
rect 415 -3339 416 -3337
rect 422 -3333 423 -3331
rect 422 -3339 423 -3337
rect 429 -3333 430 -3331
rect 429 -3339 430 -3337
rect 436 -3333 437 -3331
rect 436 -3339 437 -3337
rect 443 -3333 444 -3331
rect 446 -3333 447 -3331
rect 443 -3339 444 -3337
rect 446 -3339 447 -3337
rect 450 -3333 451 -3331
rect 450 -3339 451 -3337
rect 457 -3333 458 -3331
rect 457 -3339 458 -3337
rect 464 -3333 465 -3331
rect 467 -3333 468 -3331
rect 467 -3339 468 -3337
rect 471 -3333 472 -3331
rect 471 -3339 472 -3337
rect 478 -3333 479 -3331
rect 478 -3339 479 -3337
rect 485 -3333 486 -3331
rect 485 -3339 486 -3337
rect 492 -3333 493 -3331
rect 492 -3339 493 -3337
rect 499 -3333 500 -3331
rect 499 -3339 500 -3337
rect 506 -3333 507 -3331
rect 506 -3339 507 -3337
rect 513 -3333 514 -3331
rect 513 -3339 514 -3337
rect 520 -3333 521 -3331
rect 520 -3339 521 -3337
rect 527 -3333 528 -3331
rect 527 -3339 528 -3337
rect 534 -3333 535 -3331
rect 534 -3339 535 -3337
rect 541 -3333 542 -3331
rect 544 -3339 545 -3337
rect 548 -3333 549 -3331
rect 548 -3339 549 -3337
rect 555 -3333 556 -3331
rect 555 -3339 556 -3337
rect 562 -3333 563 -3331
rect 562 -3339 563 -3337
rect 572 -3333 573 -3331
rect 569 -3339 570 -3337
rect 572 -3339 573 -3337
rect 576 -3333 577 -3331
rect 576 -3339 577 -3337
rect 583 -3333 584 -3331
rect 583 -3339 584 -3337
rect 590 -3333 591 -3331
rect 593 -3333 594 -3331
rect 593 -3339 594 -3337
rect 597 -3333 598 -3331
rect 597 -3339 598 -3337
rect 604 -3333 605 -3331
rect 604 -3339 605 -3337
rect 611 -3333 612 -3331
rect 611 -3339 612 -3337
rect 618 -3333 619 -3331
rect 618 -3339 619 -3337
rect 621 -3339 622 -3337
rect 625 -3333 626 -3331
rect 625 -3339 626 -3337
rect 632 -3333 633 -3331
rect 632 -3339 633 -3337
rect 639 -3333 640 -3331
rect 639 -3339 640 -3337
rect 646 -3333 647 -3331
rect 646 -3339 647 -3337
rect 653 -3333 654 -3331
rect 653 -3339 654 -3337
rect 660 -3333 661 -3331
rect 660 -3339 661 -3337
rect 667 -3333 668 -3331
rect 670 -3333 671 -3331
rect 667 -3339 668 -3337
rect 674 -3333 675 -3331
rect 674 -3339 675 -3337
rect 681 -3333 682 -3331
rect 684 -3333 685 -3331
rect 681 -3339 682 -3337
rect 688 -3333 689 -3331
rect 688 -3339 689 -3337
rect 695 -3333 696 -3331
rect 695 -3339 696 -3337
rect 702 -3333 703 -3331
rect 702 -3339 703 -3337
rect 709 -3333 710 -3331
rect 712 -3333 713 -3331
rect 709 -3339 710 -3337
rect 712 -3339 713 -3337
rect 716 -3333 717 -3331
rect 716 -3339 717 -3337
rect 723 -3333 724 -3331
rect 723 -3339 724 -3337
rect 730 -3333 731 -3331
rect 730 -3339 731 -3337
rect 737 -3333 738 -3331
rect 737 -3339 738 -3337
rect 740 -3339 741 -3337
rect 744 -3333 745 -3331
rect 744 -3339 745 -3337
rect 751 -3333 752 -3331
rect 751 -3339 752 -3337
rect 758 -3333 759 -3331
rect 758 -3339 759 -3337
rect 765 -3333 766 -3331
rect 765 -3339 766 -3337
rect 772 -3333 773 -3331
rect 772 -3339 773 -3337
rect 779 -3333 780 -3331
rect 779 -3339 780 -3337
rect 786 -3333 787 -3331
rect 786 -3339 787 -3337
rect 793 -3333 794 -3331
rect 793 -3339 794 -3337
rect 800 -3333 801 -3331
rect 800 -3339 801 -3337
rect 807 -3333 808 -3331
rect 807 -3339 808 -3337
rect 814 -3333 815 -3331
rect 814 -3339 815 -3337
rect 821 -3333 822 -3331
rect 821 -3339 822 -3337
rect 828 -3333 829 -3331
rect 828 -3339 829 -3337
rect 835 -3333 836 -3331
rect 838 -3333 839 -3331
rect 842 -3333 843 -3331
rect 845 -3333 846 -3331
rect 842 -3339 843 -3337
rect 845 -3339 846 -3337
rect 849 -3333 850 -3331
rect 849 -3339 850 -3337
rect 856 -3333 857 -3331
rect 856 -3339 857 -3337
rect 863 -3333 864 -3331
rect 863 -3339 864 -3337
rect 870 -3333 871 -3331
rect 870 -3339 871 -3337
rect 877 -3333 878 -3331
rect 877 -3339 878 -3337
rect 884 -3333 885 -3331
rect 884 -3339 885 -3337
rect 891 -3333 892 -3331
rect 891 -3339 892 -3337
rect 898 -3333 899 -3331
rect 898 -3339 899 -3337
rect 905 -3333 906 -3331
rect 905 -3339 906 -3337
rect 912 -3333 913 -3331
rect 912 -3339 913 -3337
rect 919 -3333 920 -3331
rect 919 -3339 920 -3337
rect 926 -3333 927 -3331
rect 926 -3339 927 -3337
rect 933 -3333 934 -3331
rect 936 -3333 937 -3331
rect 933 -3339 934 -3337
rect 936 -3339 937 -3337
rect 940 -3333 941 -3331
rect 940 -3339 941 -3337
rect 947 -3339 948 -3337
rect 954 -3333 955 -3331
rect 954 -3339 955 -3337
rect 961 -3333 962 -3331
rect 961 -3339 962 -3337
rect 975 -3333 976 -3331
rect 975 -3339 976 -3337
rect 989 -3333 990 -3331
rect 989 -3339 990 -3337
rect 1059 -3333 1060 -3331
rect 1059 -3339 1060 -3337
rect 1062 -3339 1063 -3337
rect 1066 -3333 1067 -3331
rect 1066 -3339 1067 -3337
rect 1073 -3333 1074 -3331
rect 1073 -3339 1074 -3337
rect 1080 -3333 1081 -3331
rect 1080 -3339 1081 -3337
rect 1094 -3333 1095 -3331
rect 1097 -3333 1098 -3331
rect 1097 -3339 1098 -3337
rect 1108 -3333 1109 -3331
rect 1108 -3339 1109 -3337
rect 1115 -3333 1116 -3331
rect 1115 -3339 1116 -3337
rect 1136 -3333 1137 -3331
rect 1139 -3339 1140 -3337
rect 1143 -3333 1144 -3331
rect 1143 -3339 1144 -3337
rect 1213 -3333 1214 -3331
rect 1213 -3339 1214 -3337
rect 1290 -3333 1291 -3331
rect 1290 -3339 1291 -3337
rect 1360 -3333 1361 -3331
rect 1360 -3339 1361 -3337
rect 1367 -3333 1368 -3331
rect 1367 -3339 1368 -3337
rect 1409 -3333 1410 -3331
rect 1409 -3339 1410 -3337
rect 177 -3398 178 -3396
rect 177 -3404 178 -3402
rect 184 -3398 185 -3396
rect 184 -3404 185 -3402
rect 191 -3398 192 -3396
rect 191 -3404 192 -3402
rect 198 -3398 199 -3396
rect 198 -3404 199 -3402
rect 205 -3398 206 -3396
rect 205 -3404 206 -3402
rect 212 -3398 213 -3396
rect 212 -3404 213 -3402
rect 219 -3398 220 -3396
rect 219 -3404 220 -3402
rect 226 -3398 227 -3396
rect 229 -3398 230 -3396
rect 226 -3404 227 -3402
rect 229 -3404 230 -3402
rect 233 -3404 234 -3402
rect 240 -3398 241 -3396
rect 240 -3404 241 -3402
rect 247 -3398 248 -3396
rect 247 -3404 248 -3402
rect 254 -3398 255 -3396
rect 254 -3404 255 -3402
rect 261 -3398 262 -3396
rect 261 -3404 262 -3402
rect 268 -3398 269 -3396
rect 268 -3404 269 -3402
rect 275 -3398 276 -3396
rect 275 -3404 276 -3402
rect 282 -3398 283 -3396
rect 282 -3404 283 -3402
rect 289 -3398 290 -3396
rect 289 -3404 290 -3402
rect 296 -3398 297 -3396
rect 296 -3404 297 -3402
rect 303 -3398 304 -3396
rect 306 -3398 307 -3396
rect 303 -3404 304 -3402
rect 310 -3398 311 -3396
rect 310 -3404 311 -3402
rect 317 -3398 318 -3396
rect 317 -3404 318 -3402
rect 324 -3398 325 -3396
rect 324 -3404 325 -3402
rect 331 -3398 332 -3396
rect 331 -3404 332 -3402
rect 341 -3404 342 -3402
rect 345 -3398 346 -3396
rect 345 -3404 346 -3402
rect 352 -3398 353 -3396
rect 355 -3398 356 -3396
rect 355 -3404 356 -3402
rect 359 -3398 360 -3396
rect 359 -3404 360 -3402
rect 366 -3398 367 -3396
rect 366 -3404 367 -3402
rect 373 -3398 374 -3396
rect 373 -3404 374 -3402
rect 380 -3398 381 -3396
rect 383 -3404 384 -3402
rect 387 -3398 388 -3396
rect 387 -3404 388 -3402
rect 394 -3398 395 -3396
rect 397 -3398 398 -3396
rect 394 -3404 395 -3402
rect 401 -3398 402 -3396
rect 401 -3404 402 -3402
rect 408 -3398 409 -3396
rect 408 -3404 409 -3402
rect 415 -3398 416 -3396
rect 415 -3404 416 -3402
rect 422 -3398 423 -3396
rect 422 -3404 423 -3402
rect 429 -3398 430 -3396
rect 429 -3404 430 -3402
rect 436 -3398 437 -3396
rect 436 -3404 437 -3402
rect 443 -3398 444 -3396
rect 443 -3404 444 -3402
rect 450 -3398 451 -3396
rect 450 -3404 451 -3402
rect 457 -3398 458 -3396
rect 457 -3404 458 -3402
rect 464 -3398 465 -3396
rect 467 -3404 468 -3402
rect 471 -3398 472 -3396
rect 471 -3404 472 -3402
rect 478 -3398 479 -3396
rect 478 -3404 479 -3402
rect 485 -3398 486 -3396
rect 488 -3398 489 -3396
rect 488 -3404 489 -3402
rect 495 -3398 496 -3396
rect 495 -3404 496 -3402
rect 499 -3398 500 -3396
rect 499 -3404 500 -3402
rect 506 -3404 507 -3402
rect 513 -3398 514 -3396
rect 513 -3404 514 -3402
rect 520 -3398 521 -3396
rect 520 -3404 521 -3402
rect 527 -3398 528 -3396
rect 527 -3404 528 -3402
rect 534 -3398 535 -3396
rect 537 -3398 538 -3396
rect 534 -3404 535 -3402
rect 541 -3398 542 -3396
rect 541 -3404 542 -3402
rect 548 -3398 549 -3396
rect 548 -3404 549 -3402
rect 558 -3398 559 -3396
rect 558 -3404 559 -3402
rect 562 -3398 563 -3396
rect 562 -3404 563 -3402
rect 569 -3398 570 -3396
rect 569 -3404 570 -3402
rect 576 -3398 577 -3396
rect 576 -3404 577 -3402
rect 583 -3398 584 -3396
rect 583 -3404 584 -3402
rect 590 -3398 591 -3396
rect 590 -3404 591 -3402
rect 597 -3398 598 -3396
rect 597 -3404 598 -3402
rect 604 -3398 605 -3396
rect 604 -3404 605 -3402
rect 611 -3398 612 -3396
rect 611 -3404 612 -3402
rect 618 -3398 619 -3396
rect 618 -3404 619 -3402
rect 625 -3398 626 -3396
rect 625 -3404 626 -3402
rect 632 -3398 633 -3396
rect 632 -3404 633 -3402
rect 639 -3398 640 -3396
rect 639 -3404 640 -3402
rect 646 -3398 647 -3396
rect 646 -3404 647 -3402
rect 653 -3398 654 -3396
rect 653 -3404 654 -3402
rect 660 -3398 661 -3396
rect 660 -3404 661 -3402
rect 667 -3398 668 -3396
rect 674 -3398 675 -3396
rect 674 -3404 675 -3402
rect 681 -3398 682 -3396
rect 681 -3404 682 -3402
rect 688 -3398 689 -3396
rect 688 -3404 689 -3402
rect 695 -3398 696 -3396
rect 695 -3404 696 -3402
rect 702 -3398 703 -3396
rect 709 -3398 710 -3396
rect 709 -3404 710 -3402
rect 716 -3398 717 -3396
rect 716 -3404 717 -3402
rect 723 -3398 724 -3396
rect 723 -3404 724 -3402
rect 730 -3398 731 -3396
rect 730 -3404 731 -3402
rect 733 -3404 734 -3402
rect 737 -3398 738 -3396
rect 737 -3404 738 -3402
rect 744 -3398 745 -3396
rect 744 -3404 745 -3402
rect 751 -3398 752 -3396
rect 751 -3404 752 -3402
rect 758 -3398 759 -3396
rect 758 -3404 759 -3402
rect 765 -3398 766 -3396
rect 765 -3404 766 -3402
rect 775 -3398 776 -3396
rect 772 -3404 773 -3402
rect 775 -3404 776 -3402
rect 779 -3398 780 -3396
rect 779 -3404 780 -3402
rect 814 -3398 815 -3396
rect 814 -3404 815 -3402
rect 821 -3398 822 -3396
rect 821 -3404 822 -3402
rect 828 -3398 829 -3396
rect 831 -3398 832 -3396
rect 835 -3398 836 -3396
rect 835 -3404 836 -3402
rect 845 -3398 846 -3396
rect 842 -3404 843 -3402
rect 845 -3404 846 -3402
rect 849 -3398 850 -3396
rect 849 -3404 850 -3402
rect 856 -3398 857 -3396
rect 856 -3404 857 -3402
rect 863 -3398 864 -3396
rect 866 -3398 867 -3396
rect 863 -3404 864 -3402
rect 870 -3398 871 -3396
rect 870 -3404 871 -3402
rect 877 -3398 878 -3396
rect 877 -3404 878 -3402
rect 884 -3398 885 -3396
rect 884 -3404 885 -3402
rect 894 -3398 895 -3396
rect 891 -3404 892 -3402
rect 905 -3398 906 -3396
rect 905 -3404 906 -3402
rect 912 -3398 913 -3396
rect 912 -3404 913 -3402
rect 919 -3398 920 -3396
rect 919 -3404 920 -3402
rect 926 -3398 927 -3396
rect 926 -3404 927 -3402
rect 940 -3398 941 -3396
rect 940 -3404 941 -3402
rect 989 -3398 990 -3396
rect 989 -3404 990 -3402
rect 996 -3398 997 -3396
rect 996 -3404 997 -3402
rect 1073 -3398 1074 -3396
rect 1073 -3404 1074 -3402
rect 1115 -3398 1116 -3396
rect 1115 -3404 1116 -3402
rect 1122 -3398 1123 -3396
rect 1122 -3404 1123 -3402
rect 1213 -3398 1214 -3396
rect 1213 -3404 1214 -3402
rect 1353 -3398 1354 -3396
rect 1353 -3404 1354 -3402
rect 1360 -3398 1361 -3396
rect 1360 -3404 1361 -3402
rect 1367 -3398 1368 -3396
rect 1367 -3404 1368 -3402
rect 1409 -3398 1410 -3396
rect 1409 -3404 1410 -3402
rect 222 -3441 223 -3439
rect 222 -3447 223 -3445
rect 240 -3441 241 -3439
rect 240 -3447 241 -3445
rect 254 -3441 255 -3439
rect 254 -3447 255 -3445
rect 264 -3441 265 -3439
rect 264 -3447 265 -3445
rect 268 -3441 269 -3439
rect 268 -3447 269 -3445
rect 275 -3441 276 -3439
rect 275 -3447 276 -3445
rect 282 -3441 283 -3439
rect 282 -3447 283 -3445
rect 289 -3447 290 -3445
rect 292 -3447 293 -3445
rect 296 -3441 297 -3439
rect 296 -3447 297 -3445
rect 303 -3441 304 -3439
rect 306 -3447 307 -3445
rect 310 -3441 311 -3439
rect 310 -3447 311 -3445
rect 317 -3441 318 -3439
rect 317 -3447 318 -3445
rect 324 -3441 325 -3439
rect 327 -3441 328 -3439
rect 327 -3447 328 -3445
rect 338 -3441 339 -3439
rect 341 -3441 342 -3439
rect 345 -3441 346 -3439
rect 345 -3447 346 -3445
rect 352 -3441 353 -3439
rect 352 -3447 353 -3445
rect 359 -3441 360 -3439
rect 359 -3447 360 -3445
rect 373 -3441 374 -3439
rect 373 -3447 374 -3445
rect 387 -3441 388 -3439
rect 387 -3447 388 -3445
rect 394 -3441 395 -3439
rect 394 -3447 395 -3445
rect 401 -3441 402 -3439
rect 401 -3447 402 -3445
rect 408 -3441 409 -3439
rect 408 -3447 409 -3445
rect 422 -3441 423 -3439
rect 422 -3447 423 -3445
rect 429 -3441 430 -3439
rect 429 -3447 430 -3445
rect 436 -3441 437 -3439
rect 436 -3447 437 -3445
rect 443 -3441 444 -3439
rect 443 -3447 444 -3445
rect 450 -3441 451 -3439
rect 450 -3447 451 -3445
rect 471 -3441 472 -3439
rect 471 -3447 472 -3445
rect 485 -3441 486 -3439
rect 485 -3447 486 -3445
rect 492 -3441 493 -3439
rect 492 -3447 493 -3445
rect 499 -3441 500 -3439
rect 502 -3447 503 -3445
rect 534 -3441 535 -3439
rect 534 -3447 535 -3445
rect 541 -3441 542 -3439
rect 541 -3447 542 -3445
rect 548 -3441 549 -3439
rect 548 -3447 549 -3445
rect 555 -3441 556 -3439
rect 555 -3447 556 -3445
rect 562 -3441 563 -3439
rect 562 -3447 563 -3445
rect 569 -3441 570 -3439
rect 569 -3447 570 -3445
rect 572 -3447 573 -3445
rect 576 -3441 577 -3439
rect 576 -3447 577 -3445
rect 583 -3441 584 -3439
rect 583 -3447 584 -3445
rect 597 -3441 598 -3439
rect 597 -3447 598 -3445
rect 625 -3441 626 -3439
rect 625 -3447 626 -3445
rect 632 -3441 633 -3439
rect 632 -3447 633 -3445
rect 639 -3441 640 -3439
rect 642 -3441 643 -3439
rect 639 -3447 640 -3445
rect 642 -3447 643 -3445
rect 646 -3441 647 -3439
rect 646 -3447 647 -3445
rect 653 -3441 654 -3439
rect 653 -3447 654 -3445
rect 660 -3441 661 -3439
rect 660 -3447 661 -3445
rect 667 -3447 668 -3445
rect 674 -3441 675 -3439
rect 674 -3447 675 -3445
rect 681 -3441 682 -3439
rect 681 -3447 682 -3445
rect 688 -3441 689 -3439
rect 688 -3447 689 -3445
rect 695 -3441 696 -3439
rect 695 -3447 696 -3445
rect 702 -3441 703 -3439
rect 702 -3447 703 -3445
rect 709 -3441 710 -3439
rect 709 -3447 710 -3445
rect 719 -3441 720 -3439
rect 716 -3447 717 -3445
rect 719 -3447 720 -3445
rect 723 -3441 724 -3439
rect 723 -3447 724 -3445
rect 726 -3447 727 -3445
rect 730 -3441 731 -3439
rect 733 -3441 734 -3439
rect 730 -3447 731 -3445
rect 737 -3447 738 -3445
rect 740 -3447 741 -3445
rect 744 -3441 745 -3439
rect 744 -3447 745 -3445
rect 751 -3441 752 -3439
rect 751 -3447 752 -3445
rect 758 -3441 759 -3439
rect 758 -3447 759 -3445
rect 765 -3441 766 -3439
rect 765 -3447 766 -3445
rect 772 -3441 773 -3439
rect 779 -3441 780 -3439
rect 782 -3441 783 -3439
rect 779 -3447 780 -3445
rect 782 -3447 783 -3445
rect 821 -3441 822 -3439
rect 821 -3447 822 -3445
rect 831 -3441 832 -3439
rect 828 -3447 829 -3445
rect 831 -3447 832 -3445
rect 835 -3441 836 -3439
rect 835 -3447 836 -3445
rect 842 -3441 843 -3439
rect 842 -3447 843 -3445
rect 849 -3441 850 -3439
rect 849 -3447 850 -3445
rect 856 -3441 857 -3439
rect 856 -3447 857 -3445
rect 863 -3441 864 -3439
rect 863 -3447 864 -3445
rect 870 -3441 871 -3439
rect 870 -3447 871 -3445
rect 884 -3441 885 -3439
rect 884 -3447 885 -3445
rect 912 -3441 913 -3439
rect 912 -3447 913 -3445
rect 919 -3441 920 -3439
rect 919 -3447 920 -3445
rect 926 -3441 927 -3439
rect 926 -3447 927 -3445
rect 940 -3441 941 -3439
rect 940 -3447 941 -3445
rect 947 -3441 948 -3439
rect 947 -3447 948 -3445
rect 954 -3441 955 -3439
rect 954 -3447 955 -3445
rect 957 -3447 958 -3445
rect 961 -3441 962 -3439
rect 964 -3441 965 -3439
rect 961 -3447 962 -3445
rect 964 -3447 965 -3445
rect 968 -3441 969 -3439
rect 968 -3447 969 -3445
rect 975 -3441 976 -3439
rect 975 -3447 976 -3445
rect 982 -3441 983 -3439
rect 982 -3447 983 -3445
rect 989 -3441 990 -3439
rect 989 -3447 990 -3445
rect 996 -3441 997 -3439
rect 996 -3447 997 -3445
rect 1010 -3441 1011 -3439
rect 1010 -3447 1011 -3445
rect 1073 -3441 1074 -3439
rect 1073 -3447 1074 -3445
rect 1094 -3441 1095 -3439
rect 1094 -3447 1095 -3445
rect 1115 -3441 1116 -3439
rect 1115 -3447 1116 -3445
rect 1122 -3441 1123 -3439
rect 1122 -3447 1123 -3445
rect 1213 -3441 1214 -3439
rect 1213 -3447 1214 -3445
rect 1353 -3441 1354 -3439
rect 1353 -3447 1354 -3445
rect 1360 -3441 1361 -3439
rect 1360 -3447 1361 -3445
rect 1395 -3441 1396 -3439
rect 1395 -3447 1396 -3445
rect 1409 -3441 1410 -3439
rect 1409 -3447 1410 -3445
rect 254 -3468 255 -3466
rect 254 -3474 255 -3472
rect 261 -3468 262 -3466
rect 261 -3474 262 -3472
rect 303 -3468 304 -3466
rect 303 -3474 304 -3472
rect 317 -3468 318 -3466
rect 317 -3474 318 -3472
rect 327 -3468 328 -3466
rect 327 -3474 328 -3472
rect 331 -3468 332 -3466
rect 331 -3474 332 -3472
rect 338 -3468 339 -3466
rect 338 -3474 339 -3472
rect 352 -3468 353 -3466
rect 352 -3474 353 -3472
rect 359 -3468 360 -3466
rect 359 -3474 360 -3472
rect 380 -3468 381 -3466
rect 380 -3474 381 -3472
rect 394 -3468 395 -3466
rect 394 -3474 395 -3472
rect 401 -3468 402 -3466
rect 401 -3474 402 -3472
rect 408 -3474 409 -3472
rect 411 -3474 412 -3472
rect 415 -3468 416 -3466
rect 415 -3474 416 -3472
rect 422 -3468 423 -3466
rect 425 -3468 426 -3466
rect 429 -3468 430 -3466
rect 429 -3474 430 -3472
rect 436 -3474 437 -3472
rect 439 -3474 440 -3472
rect 443 -3468 444 -3466
rect 443 -3474 444 -3472
rect 457 -3468 458 -3466
rect 460 -3468 461 -3466
rect 464 -3468 465 -3466
rect 467 -3474 468 -3472
rect 471 -3468 472 -3466
rect 471 -3474 472 -3472
rect 478 -3468 479 -3466
rect 478 -3474 479 -3472
rect 485 -3468 486 -3466
rect 485 -3474 486 -3472
rect 492 -3468 493 -3466
rect 492 -3474 493 -3472
rect 499 -3474 500 -3472
rect 502 -3474 503 -3472
rect 506 -3468 507 -3466
rect 506 -3474 507 -3472
rect 513 -3474 514 -3472
rect 516 -3474 517 -3472
rect 520 -3468 521 -3466
rect 520 -3474 521 -3472
rect 541 -3468 542 -3466
rect 541 -3474 542 -3472
rect 548 -3468 549 -3466
rect 548 -3474 549 -3472
rect 555 -3468 556 -3466
rect 562 -3468 563 -3466
rect 562 -3474 563 -3472
rect 569 -3468 570 -3466
rect 569 -3474 570 -3472
rect 576 -3468 577 -3466
rect 576 -3474 577 -3472
rect 583 -3468 584 -3466
rect 583 -3474 584 -3472
rect 604 -3468 605 -3466
rect 604 -3474 605 -3472
rect 614 -3468 615 -3466
rect 611 -3474 612 -3472
rect 614 -3474 615 -3472
rect 621 -3468 622 -3466
rect 621 -3474 622 -3472
rect 625 -3468 626 -3466
rect 625 -3474 626 -3472
rect 646 -3468 647 -3466
rect 646 -3474 647 -3472
rect 653 -3468 654 -3466
rect 653 -3474 654 -3472
rect 660 -3468 661 -3466
rect 660 -3474 661 -3472
rect 674 -3468 675 -3466
rect 674 -3474 675 -3472
rect 681 -3468 682 -3466
rect 681 -3474 682 -3472
rect 688 -3468 689 -3466
rect 691 -3468 692 -3466
rect 695 -3468 696 -3466
rect 698 -3468 699 -3466
rect 695 -3474 696 -3472
rect 698 -3474 699 -3472
rect 709 -3468 710 -3466
rect 709 -3474 710 -3472
rect 737 -3468 738 -3466
rect 737 -3474 738 -3472
rect 758 -3468 759 -3466
rect 758 -3474 759 -3472
rect 821 -3468 822 -3466
rect 824 -3468 825 -3466
rect 821 -3474 822 -3472
rect 835 -3468 836 -3466
rect 835 -3474 836 -3472
rect 842 -3468 843 -3466
rect 842 -3474 843 -3472
rect 849 -3468 850 -3466
rect 852 -3474 853 -3472
rect 856 -3468 857 -3466
rect 856 -3474 857 -3472
rect 870 -3468 871 -3466
rect 870 -3474 871 -3472
rect 884 -3468 885 -3466
rect 884 -3474 885 -3472
rect 891 -3468 892 -3466
rect 891 -3474 892 -3472
rect 912 -3468 913 -3466
rect 912 -3474 913 -3472
rect 919 -3468 920 -3466
rect 919 -3474 920 -3472
rect 926 -3468 927 -3466
rect 926 -3474 927 -3472
rect 933 -3468 934 -3466
rect 933 -3474 934 -3472
rect 940 -3468 941 -3466
rect 940 -3474 941 -3472
rect 989 -3468 990 -3466
rect 989 -3474 990 -3472
rect 996 -3468 997 -3466
rect 996 -3474 997 -3472
rect 1066 -3468 1067 -3466
rect 1066 -3474 1067 -3472
rect 1073 -3468 1074 -3466
rect 1076 -3468 1077 -3466
rect 1115 -3468 1116 -3466
rect 1115 -3474 1116 -3472
rect 1122 -3468 1123 -3466
rect 1122 -3474 1123 -3472
rect 1213 -3468 1214 -3466
rect 1213 -3474 1214 -3472
rect 1220 -3468 1221 -3466
rect 1223 -3468 1224 -3466
rect 1220 -3474 1221 -3472
rect 1227 -3468 1228 -3466
rect 1227 -3474 1228 -3472
rect 1353 -3468 1354 -3466
rect 1353 -3474 1354 -3472
rect 1360 -3468 1361 -3466
rect 1360 -3474 1361 -3472
rect 1409 -3468 1410 -3466
rect 1409 -3474 1410 -3472
rect 1412 -3474 1413 -3472
rect 1416 -3468 1417 -3466
rect 1416 -3474 1417 -3472
rect 261 -3491 262 -3489
rect 261 -3497 262 -3495
rect 268 -3491 269 -3489
rect 268 -3497 269 -3495
rect 310 -3491 311 -3489
rect 310 -3497 311 -3495
rect 331 -3491 332 -3489
rect 331 -3497 332 -3495
rect 338 -3491 339 -3489
rect 338 -3497 339 -3495
rect 345 -3497 346 -3495
rect 352 -3491 353 -3489
rect 352 -3497 353 -3495
rect 408 -3491 409 -3489
rect 408 -3497 409 -3495
rect 418 -3491 419 -3489
rect 418 -3497 419 -3495
rect 429 -3491 430 -3489
rect 429 -3497 430 -3495
rect 436 -3491 437 -3489
rect 436 -3497 437 -3495
rect 478 -3491 479 -3489
rect 478 -3497 479 -3495
rect 541 -3491 542 -3489
rect 541 -3497 542 -3495
rect 548 -3491 549 -3489
rect 548 -3497 549 -3495
rect 555 -3497 556 -3495
rect 569 -3491 570 -3489
rect 569 -3497 570 -3495
rect 576 -3491 577 -3489
rect 576 -3497 577 -3495
rect 583 -3491 584 -3489
rect 583 -3497 584 -3495
rect 590 -3491 591 -3489
rect 590 -3497 591 -3495
rect 597 -3491 598 -3489
rect 597 -3497 598 -3495
rect 646 -3491 647 -3489
rect 646 -3497 647 -3495
rect 653 -3491 654 -3489
rect 653 -3497 654 -3495
rect 660 -3491 661 -3489
rect 660 -3497 661 -3495
rect 681 -3491 682 -3489
rect 681 -3497 682 -3495
rect 688 -3491 689 -3489
rect 688 -3497 689 -3495
rect 716 -3491 717 -3489
rect 716 -3497 717 -3495
rect 726 -3491 727 -3489
rect 723 -3497 724 -3495
rect 828 -3491 829 -3489
rect 828 -3497 829 -3495
rect 835 -3491 836 -3489
rect 835 -3497 836 -3495
rect 842 -3497 843 -3495
rect 849 -3491 850 -3489
rect 849 -3497 850 -3495
rect 877 -3491 878 -3489
rect 877 -3497 878 -3495
rect 884 -3491 885 -3489
rect 887 -3491 888 -3489
rect 898 -3491 899 -3489
rect 898 -3497 899 -3495
rect 905 -3491 906 -3489
rect 905 -3497 906 -3495
rect 912 -3491 913 -3489
rect 912 -3497 913 -3495
rect 919 -3491 920 -3489
rect 919 -3497 920 -3495
rect 926 -3491 927 -3489
rect 926 -3497 927 -3495
rect 940 -3491 941 -3489
rect 940 -3497 941 -3495
rect 950 -3491 951 -3489
rect 950 -3497 951 -3495
rect 992 -3491 993 -3489
rect 989 -3497 990 -3495
rect 996 -3491 997 -3489
rect 996 -3497 997 -3495
rect 1094 -3491 1095 -3489
rect 1094 -3497 1095 -3495
rect 1115 -3491 1116 -3489
rect 1115 -3497 1116 -3495
rect 1118 -3497 1119 -3495
rect 1122 -3491 1123 -3489
rect 1122 -3497 1123 -3495
rect 1220 -3491 1221 -3489
rect 1353 -3491 1354 -3489
rect 1353 -3497 1354 -3495
rect 1360 -3491 1361 -3489
rect 1360 -3497 1361 -3495
rect 1409 -3491 1410 -3489
rect 1412 -3491 1413 -3489
rect 1412 -3497 1413 -3495
rect 1416 -3491 1417 -3489
rect 1416 -3497 1417 -3495
rect 271 -3506 272 -3504
rect 271 -3512 272 -3510
rect 275 -3506 276 -3504
rect 275 -3512 276 -3510
rect 324 -3506 325 -3504
rect 327 -3512 328 -3510
rect 331 -3506 332 -3504
rect 331 -3512 332 -3510
rect 355 -3506 356 -3504
rect 355 -3512 356 -3510
rect 359 -3506 360 -3504
rect 359 -3512 360 -3510
rect 541 -3506 542 -3504
rect 541 -3512 542 -3510
rect 551 -3506 552 -3504
rect 555 -3512 556 -3510
rect 565 -3506 566 -3504
rect 565 -3512 566 -3510
rect 569 -3506 570 -3504
rect 569 -3512 570 -3510
rect 576 -3506 577 -3504
rect 579 -3512 580 -3510
rect 583 -3506 584 -3504
rect 583 -3512 584 -3510
rect 660 -3512 661 -3510
rect 667 -3506 668 -3504
rect 667 -3512 668 -3510
rect 688 -3506 689 -3504
rect 691 -3506 692 -3504
rect 859 -3506 860 -3504
rect 856 -3512 857 -3510
rect 870 -3506 871 -3504
rect 870 -3512 871 -3510
rect 877 -3506 878 -3504
rect 877 -3512 878 -3510
rect 912 -3506 913 -3504
rect 915 -3512 916 -3510
rect 919 -3506 920 -3504
rect 922 -3506 923 -3504
rect 1353 -3506 1354 -3504
rect 1353 -3512 1354 -3510
rect 1360 -3512 1361 -3510
rect 1363 -3512 1364 -3510
rect 1367 -3506 1368 -3504
rect 1367 -3512 1368 -3510
<< metal1 >>
rect 282 0 346 1
rect 425 0 451 1
rect 464 0 479 1
rect 905 0 951 1
rect 317 -2 353 -1
rect 436 -2 514 -1
rect 947 -2 990 -1
rect 443 -4 458 -3
rect 226 -15 286 -14
rect 303 -15 318 -14
rect 338 -15 360 -14
rect 366 -15 437 -14
rect 450 -15 458 -14
rect 478 -15 500 -14
rect 506 -15 612 -14
rect 618 -15 626 -14
rect 891 -15 906 -14
rect 989 -15 1004 -14
rect 345 -17 374 -16
rect 380 -17 426 -16
rect 436 -17 444 -16
rect 450 -17 465 -16
rect 513 -17 549 -16
rect 579 -17 591 -16
rect 597 -17 640 -16
rect 289 -19 346 -18
rect 348 -19 409 -18
rect 422 -19 510 -18
rect 527 -19 542 -18
rect 583 -19 605 -18
rect 352 -21 388 -20
rect 394 -21 419 -20
rect 460 -21 465 -20
rect 509 -21 514 -20
rect 537 -21 675 -20
rect 352 -23 363 -22
rect 219 -34 227 -33
rect 275 -34 290 -33
rect 324 -34 367 -33
rect 387 -34 402 -33
rect 415 -34 437 -33
rect 443 -34 458 -33
rect 464 -34 472 -33
rect 492 -34 566 -33
rect 576 -34 598 -33
rect 611 -34 654 -33
rect 674 -34 724 -33
rect 758 -34 829 -33
rect 884 -34 892 -33
rect 1003 -34 1011 -33
rect 282 -36 297 -35
rect 331 -36 342 -35
rect 359 -36 433 -35
rect 436 -36 458 -35
rect 499 -36 503 -35
rect 513 -36 521 -35
rect 541 -36 556 -35
rect 583 -36 622 -35
rect 625 -36 633 -35
rect 639 -36 675 -35
rect 338 -38 346 -37
rect 366 -38 381 -37
rect 387 -38 486 -37
rect 499 -38 507 -37
rect 520 -38 528 -37
rect 551 -38 731 -37
rect 338 -40 423 -39
rect 450 -40 465 -39
rect 502 -40 507 -39
rect 523 -40 542 -39
rect 590 -40 598 -39
rect 625 -40 682 -39
rect 380 -42 395 -41
rect 408 -42 451 -41
rect 548 -42 591 -41
rect 635 -42 640 -41
rect 394 -44 538 -43
rect 408 -46 419 -45
rect 422 -46 430 -45
rect 191 -57 255 -56
rect 278 -57 283 -56
rect 289 -57 465 -56
rect 506 -57 517 -56
rect 523 -57 738 -56
rect 789 -57 864 -56
rect 884 -57 892 -56
rect 1010 -57 1018 -56
rect 205 -59 241 -58
rect 243 -59 262 -58
rect 275 -59 283 -58
rect 296 -59 304 -58
rect 317 -59 391 -58
rect 464 -59 500 -58
rect 513 -59 521 -58
rect 527 -59 587 -58
rect 597 -59 661 -58
rect 709 -59 759 -58
rect 793 -59 801 -58
rect 828 -59 899 -58
rect 219 -61 248 -60
rect 275 -61 311 -60
rect 341 -61 346 -60
rect 390 -61 479 -60
rect 562 -61 780 -60
rect 233 -63 321 -62
rect 345 -63 381 -62
rect 471 -63 500 -62
rect 569 -63 626 -62
rect 632 -63 647 -62
rect 653 -63 703 -62
rect 730 -63 808 -62
rect 299 -65 339 -64
rect 373 -65 381 -64
rect 471 -65 510 -64
rect 569 -65 584 -64
rect 590 -65 598 -64
rect 604 -65 633 -64
rect 639 -65 654 -64
rect 723 -65 731 -64
rect 219 -67 300 -66
rect 303 -67 325 -66
rect 338 -67 549 -66
rect 576 -67 591 -66
rect 604 -67 629 -66
rect 681 -67 724 -66
rect 324 -69 535 -68
rect 555 -69 577 -68
rect 611 -69 619 -68
rect 621 -69 689 -68
rect 373 -71 444 -70
rect 485 -71 549 -70
rect 572 -71 612 -70
rect 614 -71 668 -70
rect 674 -71 682 -70
rect 436 -73 444 -72
rect 457 -73 486 -72
rect 520 -73 640 -72
rect 383 -75 458 -74
rect 541 -75 556 -74
rect 422 -77 437 -76
rect 422 -79 493 -78
rect 429 -81 493 -80
rect 415 -83 430 -82
rect 415 -85 451 -84
rect 331 -87 451 -86
rect 331 -89 360 -88
rect 352 -91 360 -90
rect 352 -93 367 -92
rect 366 -95 395 -94
rect 394 -97 783 -96
rect 114 -108 192 -107
rect 198 -108 297 -107
rect 299 -108 391 -107
rect 471 -108 563 -107
rect 565 -108 696 -107
rect 723 -108 787 -107
rect 793 -108 857 -107
rect 891 -108 920 -107
rect 1010 -108 1137 -107
rect 121 -110 384 -109
rect 387 -110 451 -109
rect 509 -110 563 -109
rect 572 -110 745 -109
rect 782 -110 1172 -109
rect 135 -112 300 -111
rect 334 -112 724 -111
rect 737 -112 843 -111
rect 898 -112 941 -111
rect 1017 -112 1025 -111
rect 142 -114 521 -113
rect 537 -114 822 -113
rect 863 -114 899 -113
rect 149 -116 374 -115
rect 380 -116 542 -115
rect 558 -116 605 -115
rect 611 -116 773 -115
rect 800 -116 878 -115
rect 156 -118 311 -117
rect 369 -118 535 -117
rect 583 -118 591 -117
rect 593 -118 759 -117
rect 807 -118 871 -117
rect 163 -120 206 -119
rect 212 -120 454 -119
rect 516 -120 801 -119
rect 863 -120 1014 -119
rect 170 -122 290 -121
rect 310 -122 409 -121
rect 443 -122 472 -121
rect 614 -122 738 -121
rect 177 -124 230 -123
rect 240 -124 304 -123
rect 408 -124 605 -123
rect 618 -124 794 -123
rect 184 -126 220 -125
rect 226 -126 514 -125
rect 586 -126 619 -125
rect 625 -126 850 -125
rect 191 -128 395 -127
rect 415 -128 444 -127
rect 450 -128 500 -127
rect 513 -128 542 -127
rect 576 -128 626 -127
rect 628 -128 717 -127
rect 205 -130 234 -129
rect 247 -130 374 -129
rect 394 -130 549 -129
rect 639 -130 780 -129
rect 219 -132 325 -131
rect 415 -132 507 -131
rect 639 -132 647 -131
rect 660 -132 766 -131
rect 233 -134 612 -133
rect 667 -134 752 -133
rect 247 -136 258 -135
rect 268 -136 423 -135
rect 464 -136 517 -135
rect 597 -136 647 -135
rect 688 -136 815 -135
rect 271 -138 276 -137
rect 289 -138 531 -137
rect 555 -138 598 -137
rect 632 -138 668 -137
rect 702 -138 808 -137
rect 275 -140 339 -139
rect 390 -140 423 -139
rect 464 -140 528 -139
rect 555 -140 675 -139
rect 702 -140 731 -139
rect 303 -142 524 -141
rect 527 -142 829 -141
rect 324 -144 353 -143
rect 478 -144 661 -143
rect 730 -144 836 -143
rect 338 -146 367 -145
rect 478 -146 486 -145
rect 492 -146 549 -145
rect 632 -146 710 -145
rect 128 -148 367 -147
rect 457 -148 486 -147
rect 492 -148 503 -147
rect 653 -148 689 -147
rect 345 -150 353 -149
rect 436 -150 458 -149
rect 499 -150 577 -149
rect 583 -150 654 -149
rect 656 -150 710 -149
rect 345 -152 402 -151
rect 359 -154 437 -153
rect 359 -156 430 -155
rect 317 -158 430 -157
rect 254 -160 318 -159
rect 401 -160 787 -159
rect 254 -162 332 -161
rect 331 -164 507 -163
rect 72 -175 570 -174
rect 597 -175 601 -174
rect 709 -175 885 -174
rect 898 -175 934 -174
rect 940 -175 990 -174
rect 1024 -175 1039 -174
rect 1136 -175 1186 -174
rect 86 -177 657 -176
rect 751 -177 1018 -176
rect 1171 -177 1326 -176
rect 93 -179 269 -178
rect 275 -179 297 -178
rect 310 -179 454 -178
rect 478 -179 531 -178
rect 548 -179 591 -178
rect 597 -179 633 -178
rect 772 -179 913 -178
rect 919 -179 983 -178
rect 100 -181 199 -180
rect 205 -181 402 -180
rect 446 -181 941 -180
rect 107 -183 416 -182
rect 513 -183 773 -182
rect 793 -183 1004 -182
rect 114 -185 209 -184
rect 222 -185 892 -184
rect 121 -187 237 -186
rect 240 -187 335 -186
rect 401 -187 479 -186
rect 520 -187 731 -186
rect 800 -187 899 -186
rect 121 -189 143 -188
rect 149 -189 570 -188
rect 576 -189 710 -188
rect 716 -189 794 -188
rect 807 -189 927 -188
rect 142 -191 507 -190
rect 523 -191 594 -190
rect 600 -191 633 -190
rect 674 -191 920 -190
rect 149 -193 185 -192
rect 191 -193 528 -192
rect 534 -193 577 -192
rect 625 -193 675 -192
rect 681 -193 717 -192
rect 737 -193 801 -192
rect 814 -193 1011 -192
rect 79 -195 626 -194
rect 681 -195 689 -194
rect 702 -195 738 -194
rect 744 -195 815 -194
rect 821 -195 962 -194
rect 163 -197 276 -196
rect 289 -197 297 -196
rect 310 -197 391 -196
rect 422 -197 514 -196
rect 555 -197 615 -196
rect 667 -197 745 -196
rect 828 -197 948 -196
rect 163 -199 178 -198
rect 184 -199 220 -198
rect 233 -199 416 -198
rect 432 -199 808 -198
rect 835 -199 906 -198
rect 114 -201 220 -200
rect 233 -201 370 -200
rect 436 -201 521 -200
rect 558 -201 654 -200
rect 688 -201 752 -200
rect 765 -201 836 -200
rect 856 -201 969 -200
rect 170 -203 199 -202
rect 243 -203 423 -202
rect 464 -203 535 -202
rect 562 -203 605 -202
rect 618 -203 766 -202
rect 870 -203 976 -202
rect 156 -205 171 -204
rect 177 -205 405 -204
rect 443 -205 465 -204
rect 471 -205 668 -204
rect 702 -205 759 -204
rect 786 -205 871 -204
rect 877 -205 1025 -204
rect 128 -207 444 -206
rect 471 -207 493 -206
rect 607 -207 759 -206
rect 842 -207 878 -206
rect 128 -209 227 -208
rect 229 -209 843 -208
rect 191 -211 206 -210
rect 261 -211 269 -210
rect 289 -211 353 -210
rect 387 -211 787 -210
rect 247 -213 262 -212
rect 331 -213 339 -212
rect 352 -213 367 -212
rect 380 -213 388 -212
rect 394 -213 437 -212
rect 485 -213 507 -212
rect 618 -213 647 -212
rect 660 -213 857 -212
rect 212 -215 339 -214
rect 373 -215 381 -214
rect 394 -215 552 -214
rect 611 -215 661 -214
rect 723 -215 822 -214
rect 212 -217 500 -216
rect 611 -217 955 -216
rect 247 -219 325 -218
rect 359 -219 374 -218
rect 429 -219 647 -218
rect 723 -219 864 -218
rect 135 -221 430 -220
rect 492 -221 542 -220
rect 779 -221 864 -220
rect 135 -223 255 -222
rect 317 -223 332 -222
rect 345 -223 360 -222
rect 499 -223 563 -222
rect 695 -223 780 -222
rect 254 -225 304 -224
rect 317 -225 409 -224
rect 541 -225 640 -224
rect 695 -225 832 -224
rect 303 -227 451 -226
rect 583 -227 640 -226
rect 324 -229 486 -228
rect 583 -229 850 -228
rect 345 -231 409 -230
rect 450 -231 629 -230
rect 849 -231 997 -230
rect 93 -242 486 -241
rect 488 -242 857 -241
rect 884 -242 1116 -241
rect 1185 -242 1207 -241
rect 1307 -242 1459 -241
rect 93 -244 143 -243
rect 145 -244 402 -243
rect 446 -244 493 -243
rect 502 -244 913 -243
rect 919 -244 1053 -243
rect 1325 -244 1382 -243
rect 100 -246 174 -245
rect 177 -246 479 -245
rect 485 -246 748 -245
rect 754 -246 1081 -245
rect 100 -248 237 -247
rect 247 -248 402 -247
rect 453 -248 1004 -247
rect 1038 -248 1067 -247
rect 107 -250 444 -249
rect 492 -250 507 -249
rect 537 -250 1102 -249
rect 107 -252 143 -251
rect 159 -252 258 -251
rect 303 -252 552 -251
rect 600 -252 913 -251
rect 954 -252 1109 -251
rect 128 -254 241 -253
rect 247 -254 367 -253
rect 369 -254 458 -253
rect 506 -254 528 -253
rect 551 -254 619 -253
rect 628 -254 920 -253
rect 968 -254 1032 -253
rect 79 -256 129 -255
rect 138 -256 689 -255
rect 737 -256 752 -255
rect 765 -256 1095 -255
rect 79 -258 150 -257
rect 163 -258 178 -257
rect 191 -258 195 -257
rect 205 -258 227 -257
rect 233 -258 290 -257
rect 303 -258 577 -257
rect 618 -258 629 -257
rect 632 -258 689 -257
rect 716 -258 738 -257
rect 786 -258 857 -257
rect 877 -258 955 -257
rect 975 -258 1074 -257
rect 114 -260 150 -259
rect 163 -260 185 -259
rect 191 -260 220 -259
rect 226 -260 563 -259
rect 632 -260 1018 -259
rect 114 -262 122 -261
rect 170 -262 500 -261
rect 541 -262 563 -261
rect 670 -262 808 -261
rect 821 -262 885 -261
rect 891 -262 1046 -261
rect 121 -264 353 -263
rect 366 -264 374 -263
rect 376 -264 521 -263
rect 541 -264 556 -263
rect 674 -264 969 -263
rect 982 -264 1039 -263
rect 194 -266 220 -265
rect 289 -266 395 -265
rect 450 -266 528 -265
rect 646 -266 675 -265
rect 695 -266 717 -265
rect 779 -266 822 -265
rect 835 -266 892 -265
rect 905 -266 1004 -265
rect 198 -268 577 -267
rect 625 -268 780 -267
rect 793 -268 878 -267
rect 905 -268 1025 -267
rect 198 -270 262 -269
rect 331 -270 353 -269
rect 380 -270 556 -269
rect 646 -270 983 -269
rect 989 -270 1060 -269
rect 208 -272 262 -271
rect 380 -272 1123 -271
rect 86 -274 209 -273
rect 212 -274 332 -273
rect 383 -274 605 -273
rect 709 -274 787 -273
rect 898 -274 990 -273
rect 996 -274 1088 -273
rect 86 -276 430 -275
rect 450 -276 549 -275
rect 604 -276 1011 -275
rect 184 -278 213 -277
rect 387 -278 409 -277
rect 415 -278 430 -277
rect 457 -278 465 -277
rect 478 -278 766 -277
rect 926 -278 1011 -277
rect 187 -280 465 -279
rect 499 -280 598 -279
rect 607 -280 927 -279
rect 933 -280 976 -279
rect 317 -282 416 -281
rect 513 -282 521 -281
rect 534 -282 598 -281
rect 611 -282 710 -281
rect 723 -282 794 -281
rect 842 -282 934 -281
rect 940 -282 1018 -281
rect 65 -284 535 -283
rect 590 -284 612 -283
rect 660 -284 724 -283
rect 744 -284 899 -283
rect 947 -284 997 -283
rect 317 -286 325 -285
rect 387 -286 850 -285
rect 863 -286 941 -285
rect 961 -286 1025 -285
rect 324 -288 346 -287
rect 390 -288 668 -287
rect 744 -288 836 -287
rect 870 -288 948 -287
rect 72 -290 346 -289
rect 394 -290 472 -289
rect 590 -290 871 -289
rect 72 -292 157 -291
rect 275 -292 472 -291
rect 653 -292 661 -291
rect 667 -292 773 -291
rect 800 -292 843 -291
rect 156 -294 255 -293
rect 275 -294 297 -293
rect 411 -294 850 -293
rect 170 -296 801 -295
rect 814 -296 864 -295
rect 254 -298 374 -297
rect 422 -298 514 -297
rect 639 -298 654 -297
rect 730 -298 815 -297
rect 828 -298 962 -297
rect 282 -300 297 -299
rect 422 -300 437 -299
rect 481 -300 773 -299
rect 135 -302 283 -301
rect 583 -302 640 -301
rect 681 -302 731 -301
rect 758 -302 829 -301
rect 243 -304 437 -303
rect 446 -304 759 -303
rect 569 -306 584 -305
rect 681 -306 703 -305
rect 338 -308 570 -307
rect 695 -308 703 -307
rect 338 -310 360 -309
rect 310 -312 360 -311
rect 310 -314 808 -313
rect 65 -325 381 -324
rect 446 -325 577 -324
rect 590 -325 1095 -324
rect 1101 -325 1214 -324
rect 1381 -325 1410 -324
rect 1458 -325 1522 -324
rect 72 -327 363 -326
rect 369 -327 570 -326
rect 597 -327 899 -326
rect 912 -327 1151 -326
rect 1171 -327 1224 -326
rect 72 -329 122 -328
rect 135 -329 290 -328
rect 345 -329 535 -328
rect 548 -329 1053 -328
rect 1059 -329 1165 -328
rect 1199 -329 1308 -328
rect 79 -331 188 -330
rect 205 -331 1109 -330
rect 1122 -331 1389 -330
rect 58 -333 206 -332
rect 250 -333 535 -332
rect 541 -333 549 -332
rect 551 -333 969 -332
rect 989 -333 1123 -332
rect 79 -335 150 -334
rect 166 -335 577 -334
rect 597 -335 790 -334
rect 807 -335 899 -334
rect 926 -335 990 -334
rect 1003 -335 1130 -334
rect 86 -337 384 -336
rect 478 -337 542 -336
rect 565 -337 1179 -336
rect 86 -339 594 -338
rect 604 -339 619 -338
rect 625 -339 1046 -338
rect 1066 -339 1109 -338
rect 93 -341 538 -340
rect 618 -341 661 -340
rect 667 -341 689 -340
rect 702 -341 745 -340
rect 821 -341 969 -340
rect 975 -341 1046 -340
rect 1073 -341 1186 -340
rect 93 -343 419 -342
rect 464 -343 605 -342
rect 625 -343 808 -342
rect 835 -343 913 -342
rect 961 -343 1004 -342
rect 1017 -343 1144 -342
rect 100 -345 188 -344
rect 191 -345 384 -344
rect 464 -345 556 -344
rect 583 -345 661 -344
rect 702 -345 787 -344
rect 856 -345 927 -344
rect 947 -345 1018 -344
rect 1024 -345 1095 -344
rect 100 -347 157 -346
rect 170 -347 850 -346
rect 856 -347 906 -346
rect 947 -347 1011 -346
rect 1031 -347 1137 -346
rect 121 -349 129 -348
rect 149 -349 311 -348
rect 345 -349 451 -348
rect 495 -349 514 -348
rect 555 -349 654 -348
rect 758 -349 850 -348
rect 870 -349 1053 -348
rect 1080 -349 1193 -348
rect 128 -351 304 -350
rect 310 -351 360 -350
rect 373 -351 486 -350
rect 506 -351 591 -350
rect 628 -351 731 -350
rect 765 -351 822 -350
rect 884 -351 962 -350
rect 982 -351 1067 -350
rect 1080 -351 1116 -350
rect 173 -353 570 -352
rect 583 -353 766 -352
rect 772 -353 1032 -352
rect 1038 -353 1060 -352
rect 1087 -353 1158 -352
rect 107 -355 1088 -354
rect 107 -357 115 -356
rect 173 -357 507 -356
rect 513 -357 528 -356
rect 632 -357 650 -356
rect 709 -357 773 -356
rect 786 -357 1102 -356
rect 114 -359 472 -358
rect 481 -359 654 -358
rect 730 -359 801 -358
rect 814 -359 906 -358
rect 919 -359 983 -358
rect 996 -359 1025 -358
rect 184 -361 1074 -360
rect 138 -363 185 -362
rect 194 -363 486 -362
rect 520 -363 528 -362
rect 572 -363 815 -362
rect 828 -363 885 -362
rect 891 -363 976 -362
rect 247 -365 759 -364
rect 793 -365 829 -364
rect 842 -365 892 -364
rect 940 -365 1011 -364
rect 156 -367 248 -366
rect 282 -367 391 -366
rect 415 -367 521 -366
rect 646 -367 836 -366
rect 842 -367 934 -366
rect 954 -367 1039 -366
rect 142 -369 416 -368
rect 436 -369 451 -368
rect 586 -369 934 -368
rect 142 -371 164 -370
rect 233 -371 283 -370
rect 289 -371 692 -370
rect 723 -371 794 -370
rect 863 -371 941 -370
rect 233 -373 636 -372
rect 670 -373 997 -372
rect 303 -375 339 -374
rect 376 -375 472 -374
rect 737 -375 920 -374
rect 261 -377 339 -376
rect 387 -377 801 -376
rect 877 -377 955 -376
rect 212 -379 262 -378
rect 313 -379 388 -378
rect 408 -379 724 -378
rect 747 -379 1116 -378
rect 212 -381 220 -380
rect 366 -381 409 -380
rect 436 -381 612 -380
rect 716 -381 738 -380
rect 779 -381 864 -380
rect 177 -383 220 -382
rect 443 -383 710 -382
rect 716 -383 871 -382
rect 177 -385 255 -384
rect 422 -385 444 -384
rect 562 -385 612 -384
rect 751 -385 780 -384
rect 240 -387 423 -386
rect 600 -387 878 -386
rect 240 -389 395 -388
rect 632 -389 752 -388
rect 254 -391 269 -390
rect 394 -391 402 -390
rect 198 -393 269 -392
rect 401 -393 696 -392
rect 198 -395 493 -394
rect 681 -395 696 -394
rect 275 -397 493 -396
rect 639 -397 682 -396
rect 275 -399 325 -398
rect 639 -399 675 -398
rect 324 -401 332 -400
rect 499 -401 675 -400
rect 226 -403 500 -402
rect 226 -405 318 -404
rect 331 -405 353 -404
rect 296 -407 318 -406
rect 352 -407 458 -406
rect 208 -409 458 -408
rect 296 -411 430 -410
rect 429 -413 689 -412
rect 51 -424 188 -423
rect 194 -424 759 -423
rect 838 -424 1214 -423
rect 1388 -424 1487 -423
rect 1521 -424 1543 -423
rect 58 -426 146 -425
rect 149 -426 213 -425
rect 250 -426 318 -425
rect 359 -426 591 -425
rect 611 -426 622 -425
rect 656 -426 731 -425
rect 754 -426 1123 -425
rect 1157 -426 1228 -425
rect 1409 -426 1431 -425
rect 65 -428 122 -427
rect 124 -428 1144 -427
rect 1185 -428 1214 -427
rect 72 -430 426 -429
rect 450 -430 542 -429
rect 544 -430 794 -429
rect 919 -430 1235 -429
rect 72 -432 563 -431
rect 572 -432 703 -431
rect 737 -432 794 -431
rect 870 -432 920 -431
rect 1073 -432 1158 -431
rect 1192 -432 1242 -431
rect 86 -434 174 -433
rect 177 -434 391 -433
rect 415 -434 521 -433
rect 541 -434 675 -433
rect 688 -434 843 -433
rect 1031 -434 1074 -433
rect 1080 -434 1256 -433
rect 86 -436 108 -435
rect 114 -436 150 -435
rect 163 -436 423 -435
rect 450 -436 552 -435
rect 558 -436 619 -435
rect 628 -436 703 -435
rect 821 -436 871 -435
rect 1108 -436 1186 -435
rect 1206 -436 1224 -435
rect 93 -438 685 -437
rect 691 -438 1130 -437
rect 1136 -438 1144 -437
rect 1164 -438 1193 -437
rect 93 -440 101 -439
rect 114 -440 437 -439
rect 464 -440 521 -439
rect 548 -440 563 -439
rect 583 -440 969 -439
rect 1101 -440 1130 -439
rect 1164 -440 1200 -439
rect 100 -442 199 -441
rect 212 -442 276 -441
rect 296 -442 587 -441
rect 590 -442 647 -441
rect 663 -442 787 -441
rect 824 -442 1081 -441
rect 1115 -442 1123 -441
rect 1171 -442 1207 -441
rect 121 -444 1088 -443
rect 1094 -444 1116 -443
rect 1150 -444 1172 -443
rect 135 -446 493 -445
rect 495 -446 1109 -445
rect 107 -448 136 -447
rect 138 -448 846 -447
rect 852 -448 1032 -447
rect 1045 -448 1088 -447
rect 142 -450 164 -449
rect 166 -450 248 -449
rect 257 -450 339 -449
rect 359 -450 514 -449
rect 548 -450 605 -449
rect 632 -450 1151 -449
rect 152 -452 339 -451
rect 366 -452 731 -451
rect 947 -452 1095 -451
rect 166 -454 1221 -453
rect 170 -456 300 -455
rect 317 -456 325 -455
rect 366 -456 570 -455
rect 632 -456 1252 -455
rect 177 -458 626 -457
rect 667 -458 759 -457
rect 905 -458 948 -457
rect 968 -458 983 -457
rect 1024 -458 1102 -457
rect 184 -460 220 -459
rect 247 -460 594 -459
rect 667 -460 752 -459
rect 835 -460 906 -459
rect 961 -460 983 -459
rect 989 -460 1025 -459
rect 1038 -460 1046 -459
rect 191 -462 195 -461
rect 219 -462 353 -461
rect 380 -462 605 -461
rect 695 -462 738 -461
rect 779 -462 836 -461
rect 898 -462 990 -461
rect 1017 -462 1039 -461
rect 142 -464 780 -463
rect 814 -464 899 -463
rect 954 -464 962 -463
rect 1010 -464 1018 -463
rect 191 -466 675 -465
rect 698 -466 1053 -465
rect 261 -468 325 -467
rect 331 -468 353 -467
rect 383 -468 395 -467
rect 401 -468 437 -467
rect 464 -468 661 -467
rect 723 -468 1200 -467
rect 261 -470 311 -469
rect 345 -470 381 -469
rect 394 -470 409 -469
rect 415 -470 619 -469
rect 726 -470 1137 -469
rect 275 -472 283 -471
rect 296 -472 388 -471
rect 408 -472 822 -471
rect 877 -472 1011 -471
rect 156 -474 283 -473
rect 303 -474 332 -473
rect 345 -474 468 -473
rect 471 -474 514 -473
rect 569 -474 752 -473
rect 765 -474 815 -473
rect 940 -474 955 -473
rect 1003 -474 1053 -473
rect 198 -476 388 -475
rect 418 -476 717 -475
rect 744 -476 766 -475
rect 800 -476 878 -475
rect 912 -476 1004 -475
rect 303 -478 650 -477
rect 653 -478 745 -477
rect 772 -478 801 -477
rect 863 -478 941 -477
rect 310 -480 405 -479
rect 422 -480 682 -479
rect 807 -480 864 -479
rect 884 -480 913 -479
rect 429 -482 472 -481
rect 478 -482 612 -481
rect 653 -482 689 -481
rect 709 -482 808 -481
rect 828 -482 885 -481
rect 226 -484 430 -483
rect 478 -484 500 -483
rect 506 -484 584 -483
rect 597 -484 829 -483
rect 226 -486 241 -485
rect 373 -486 507 -485
rect 534 -486 710 -485
rect 205 -488 241 -487
rect 373 -488 444 -487
rect 485 -488 598 -487
rect 681 -488 1179 -487
rect 128 -490 486 -489
rect 499 -490 720 -489
rect 1059 -490 1179 -489
rect 128 -492 363 -491
rect 443 -492 458 -491
rect 527 -492 535 -491
rect 555 -492 773 -491
rect 1059 -492 1067 -491
rect 205 -494 234 -493
rect 289 -494 528 -493
rect 555 -494 626 -493
rect 975 -494 1067 -493
rect 268 -496 290 -495
rect 457 -496 790 -495
rect 933 -496 976 -495
rect 254 -498 269 -497
rect 576 -498 724 -497
rect 926 -498 934 -497
rect 156 -500 255 -499
rect 576 -500 640 -499
rect 849 -500 927 -499
rect 369 -502 640 -501
rect 44 -513 87 -512
rect 93 -513 1389 -512
rect 1419 -513 1620 -512
rect 58 -515 647 -514
rect 649 -515 1263 -514
rect 1430 -515 1459 -514
rect 1486 -515 1529 -514
rect 1542 -515 1550 -514
rect 58 -517 748 -516
rect 751 -517 1074 -516
rect 1087 -517 1221 -516
rect 1227 -517 1438 -516
rect 65 -519 192 -518
rect 254 -519 381 -518
rect 387 -519 1158 -518
rect 1178 -519 1361 -518
rect 65 -521 237 -520
rect 264 -521 1319 -520
rect 72 -523 328 -522
rect 401 -523 570 -522
rect 590 -523 850 -522
rect 863 -523 1452 -522
rect 72 -525 661 -524
rect 663 -525 899 -524
rect 905 -525 1333 -524
rect 86 -527 150 -526
rect 156 -527 381 -526
rect 425 -527 570 -526
rect 593 -527 1067 -526
rect 1115 -527 1305 -526
rect 93 -529 234 -528
rect 268 -529 293 -528
rect 296 -529 426 -528
rect 450 -529 591 -528
rect 618 -529 1445 -528
rect 121 -531 391 -530
rect 429 -531 451 -530
rect 527 -531 619 -530
rect 621 -531 1375 -530
rect 128 -533 699 -532
rect 730 -533 804 -532
rect 821 -533 1466 -532
rect 128 -535 206 -534
rect 296 -535 643 -534
rect 646 -535 1018 -534
rect 1024 -535 1431 -534
rect 124 -537 206 -536
rect 299 -537 507 -536
rect 534 -537 549 -536
rect 555 -537 766 -536
rect 789 -537 1284 -536
rect 135 -539 657 -538
rect 660 -539 1224 -538
rect 1241 -539 1252 -538
rect 142 -541 185 -540
rect 191 -541 227 -540
rect 359 -541 528 -540
rect 555 -541 710 -540
rect 716 -541 822 -540
rect 856 -541 899 -540
rect 933 -541 1291 -540
rect 142 -543 458 -542
rect 471 -543 535 -542
rect 625 -543 717 -542
rect 744 -543 864 -542
rect 873 -543 990 -542
rect 1010 -543 1088 -542
rect 1122 -543 1354 -542
rect 114 -545 626 -544
rect 653 -545 1095 -544
rect 1129 -545 1242 -544
rect 100 -547 115 -546
rect 145 -547 1424 -546
rect 100 -549 108 -548
rect 149 -549 290 -548
rect 359 -549 395 -548
rect 471 -549 584 -548
rect 632 -549 654 -548
rect 667 -549 906 -548
rect 919 -549 990 -548
rect 1017 -549 1165 -548
rect 1185 -549 1312 -548
rect 156 -551 650 -550
rect 674 -551 752 -550
rect 754 -551 1270 -550
rect 110 -553 675 -552
rect 684 -553 1249 -552
rect 163 -555 1340 -554
rect 163 -557 234 -556
rect 268 -557 458 -556
rect 478 -557 633 -556
rect 684 -557 1004 -556
rect 1024 -557 1256 -556
rect 166 -559 248 -558
rect 355 -559 584 -558
rect 611 -559 668 -558
rect 688 -559 766 -558
rect 800 -559 1116 -558
rect 1143 -559 1368 -558
rect 184 -561 304 -560
rect 373 -561 430 -560
rect 443 -561 612 -560
rect 698 -561 1235 -560
rect 194 -563 1235 -562
rect 219 -565 374 -564
rect 394 -565 598 -564
rect 702 -565 710 -564
rect 744 -565 1277 -564
rect 219 -567 346 -566
rect 366 -567 444 -566
rect 478 -567 1228 -566
rect 198 -569 346 -568
rect 366 -569 416 -568
rect 485 -569 703 -568
rect 758 -569 857 -568
rect 884 -569 934 -568
rect 954 -569 1004 -568
rect 1034 -569 1095 -568
rect 1108 -569 1165 -568
rect 1171 -569 1186 -568
rect 1192 -569 1382 -568
rect 226 -571 325 -570
rect 495 -571 689 -570
rect 761 -571 1193 -570
rect 1199 -571 1396 -570
rect 247 -573 332 -572
rect 506 -573 514 -572
rect 562 -573 598 -572
rect 828 -573 885 -572
rect 891 -573 1011 -572
rect 1031 -573 1200 -572
rect 1206 -573 1326 -572
rect 303 -575 759 -574
rect 786 -575 829 -574
rect 835 -575 892 -574
rect 926 -575 955 -574
rect 961 -575 1074 -574
rect 1080 -575 1256 -574
rect 310 -577 416 -576
rect 481 -577 927 -576
rect 968 -577 1158 -576
rect 1213 -577 1410 -576
rect 240 -579 311 -578
rect 324 -579 1123 -578
rect 1136 -579 1207 -578
rect 240 -581 283 -580
rect 331 -581 461 -580
rect 492 -581 514 -580
rect 723 -581 836 -580
rect 842 -581 920 -580
rect 940 -581 969 -580
rect 975 -581 1144 -580
rect 1150 -581 1347 -580
rect 261 -583 283 -582
rect 317 -583 493 -582
rect 499 -583 1214 -582
rect 79 -585 262 -584
rect 275 -585 318 -584
rect 576 -585 976 -584
rect 982 -585 1403 -584
rect 79 -587 486 -586
rect 639 -587 724 -586
rect 824 -587 1081 -586
rect 1101 -587 1151 -586
rect 275 -589 423 -588
rect 436 -589 577 -588
rect 639 -589 773 -588
rect 870 -589 962 -588
rect 996 -589 1109 -588
rect 51 -591 423 -590
rect 467 -591 1102 -590
rect 51 -593 171 -592
rect 289 -593 500 -592
rect 562 -593 871 -592
rect 912 -593 997 -592
rect 1038 -593 1130 -592
rect 107 -595 437 -594
rect 681 -595 941 -594
rect 1045 -595 1172 -594
rect 170 -597 199 -596
rect 390 -597 983 -596
rect 1052 -597 1179 -596
rect 772 -599 808 -598
rect 814 -599 913 -598
rect 947 -599 1046 -598
rect 1059 -599 1137 -598
rect 607 -601 808 -600
rect 845 -601 1053 -600
rect 695 -603 1060 -602
rect 695 -605 1067 -604
rect 737 -607 815 -606
rect 845 -607 1298 -606
rect 604 -609 738 -608
rect 779 -609 1039 -608
rect 464 -611 605 -610
rect 779 -611 853 -610
rect 877 -611 948 -610
rect 408 -613 465 -612
rect 793 -613 878 -612
rect 338 -615 409 -614
rect 338 -617 353 -616
rect 404 -617 794 -616
rect 212 -619 353 -618
rect 212 -621 542 -620
rect 387 -623 542 -622
rect 65 -634 265 -633
rect 310 -634 325 -633
rect 334 -634 423 -633
rect 523 -634 612 -633
rect 618 -634 682 -633
rect 691 -634 780 -633
rect 786 -634 1340 -633
rect 1419 -634 1459 -633
rect 1549 -634 1557 -633
rect 1619 -634 1697 -633
rect 72 -636 640 -635
rect 646 -636 1480 -635
rect 1528 -636 1550 -635
rect 68 -638 73 -637
rect 121 -638 636 -637
rect 649 -638 773 -637
rect 831 -638 1410 -637
rect 1444 -638 1459 -637
rect 1465 -638 1529 -637
rect 121 -640 213 -639
rect 222 -640 1228 -639
rect 1276 -640 1487 -639
rect 128 -642 234 -641
rect 240 -642 482 -641
rect 485 -642 773 -641
rect 838 -642 1144 -641
rect 1360 -642 1410 -641
rect 1437 -642 1445 -641
rect 128 -644 283 -643
rect 296 -644 423 -643
rect 429 -644 486 -643
rect 555 -644 608 -643
rect 674 -644 1228 -643
rect 1423 -644 1438 -643
rect 159 -646 976 -645
rect 982 -646 1144 -645
rect 1164 -646 1361 -645
rect 117 -648 983 -647
rect 1017 -648 1375 -647
rect 79 -650 1018 -649
rect 1052 -650 1277 -649
rect 1318 -650 1424 -649
rect 58 -652 80 -651
rect 191 -652 619 -651
rect 674 -652 1298 -651
rect 93 -654 192 -653
rect 198 -654 1270 -653
rect 93 -656 157 -655
rect 198 -656 360 -655
rect 394 -656 458 -655
rect 492 -656 976 -655
rect 1066 -656 1165 -655
rect 1192 -656 1270 -655
rect 114 -658 493 -657
rect 555 -658 857 -657
rect 870 -658 1431 -657
rect 44 -660 115 -659
rect 201 -660 1235 -659
rect 1255 -660 1298 -659
rect 44 -662 374 -661
rect 457 -662 843 -661
rect 845 -662 1326 -661
rect 205 -664 241 -663
rect 247 -664 325 -663
rect 345 -664 573 -663
rect 590 -664 696 -663
rect 709 -664 780 -663
rect 800 -664 1319 -663
rect 149 -666 248 -665
rect 282 -666 290 -665
rect 296 -666 332 -665
rect 345 -666 608 -665
rect 677 -666 1291 -665
rect 149 -668 752 -667
rect 758 -668 1452 -667
rect 212 -670 220 -669
rect 226 -670 479 -669
rect 495 -670 843 -669
rect 926 -670 1067 -669
rect 1108 -670 1466 -669
rect 219 -672 801 -671
rect 803 -672 1375 -671
rect 1395 -672 1452 -671
rect 226 -674 262 -673
rect 275 -674 290 -673
rect 310 -674 367 -673
rect 478 -674 535 -673
rect 569 -674 612 -673
rect 653 -674 759 -673
rect 828 -674 857 -673
rect 933 -674 1032 -673
rect 1038 -674 1193 -673
rect 1206 -674 1256 -673
rect 1283 -674 1291 -673
rect 1304 -674 1396 -673
rect 170 -676 367 -675
rect 471 -676 654 -675
rect 681 -676 738 -675
rect 744 -676 1158 -675
rect 1220 -676 1326 -675
rect 142 -678 472 -677
rect 527 -678 535 -677
rect 590 -678 626 -677
rect 632 -678 745 -677
rect 751 -678 906 -677
rect 912 -678 934 -677
rect 961 -678 1109 -677
rect 1122 -678 1431 -677
rect 142 -680 437 -679
rect 527 -680 941 -679
rect 1059 -680 1158 -679
rect 1248 -680 1284 -679
rect 156 -682 1060 -681
rect 1080 -682 1207 -681
rect 1262 -682 1305 -681
rect 170 -684 451 -683
rect 597 -684 626 -683
rect 632 -684 1116 -683
rect 1129 -684 1221 -683
rect 184 -686 570 -685
rect 604 -686 1214 -685
rect 184 -688 304 -687
rect 317 -688 388 -687
rect 425 -688 738 -687
rect 761 -688 1081 -687
rect 1087 -688 1123 -687
rect 1136 -688 1340 -687
rect 86 -690 388 -689
rect 558 -690 598 -689
rect 604 -690 1333 -689
rect 86 -692 108 -691
rect 233 -692 353 -691
rect 355 -692 395 -691
rect 530 -692 1333 -691
rect 107 -694 790 -693
rect 821 -694 1039 -693
rect 1094 -694 1214 -693
rect 254 -696 353 -695
rect 359 -696 465 -695
rect 688 -696 787 -695
rect 814 -696 822 -695
rect 828 -696 1473 -695
rect 177 -698 815 -697
rect 849 -698 941 -697
rect 954 -698 1088 -697
rect 1150 -698 1235 -697
rect 177 -700 328 -699
rect 380 -700 451 -699
rect 464 -700 1417 -699
rect 254 -702 374 -701
rect 429 -702 955 -701
rect 968 -702 1116 -701
rect 1178 -702 1263 -701
rect 1388 -702 1417 -701
rect 261 -704 339 -703
rect 467 -704 969 -703
rect 989 -704 1130 -703
rect 1178 -704 1382 -703
rect 268 -706 339 -705
rect 702 -706 710 -705
rect 719 -706 1368 -705
rect 268 -708 402 -707
rect 460 -708 703 -707
rect 730 -708 1053 -707
rect 1185 -708 1389 -707
rect 135 -710 402 -709
rect 684 -710 1186 -709
rect 1311 -710 1368 -709
rect 135 -712 206 -711
rect 303 -712 416 -711
rect 733 -712 1102 -711
rect 1346 -712 1382 -711
rect 317 -714 409 -713
rect 415 -714 500 -713
rect 733 -714 1403 -713
rect 163 -716 409 -715
rect 499 -716 577 -715
rect 793 -716 850 -715
rect 873 -716 1312 -715
rect 58 -718 164 -717
rect 331 -718 381 -717
rect 576 -718 717 -717
rect 884 -718 913 -717
rect 919 -718 962 -717
rect 989 -718 1025 -717
rect 1045 -718 1151 -717
rect 1171 -718 1403 -717
rect 275 -720 717 -719
rect 877 -720 1046 -719
rect 432 -722 885 -721
rect 891 -722 920 -721
rect 929 -722 1095 -721
rect 51 -724 892 -723
rect 905 -724 1200 -723
rect 51 -726 244 -725
rect 436 -726 1025 -725
rect 1073 -726 1200 -725
rect 642 -728 1074 -727
rect 807 -730 878 -729
rect 908 -730 1347 -729
rect 723 -732 808 -731
rect 996 -732 1137 -731
rect 506 -734 724 -733
rect 947 -734 997 -733
rect 1003 -734 1172 -733
rect 257 -736 507 -735
rect 520 -736 1004 -735
rect 1010 -736 1102 -735
rect 863 -738 948 -737
rect 1020 -738 1249 -737
rect 765 -740 864 -739
rect 898 -740 1011 -739
rect 443 -742 766 -741
rect 835 -742 899 -741
rect 443 -744 661 -743
rect 835 -744 1354 -743
rect 660 -746 668 -745
rect 1241 -746 1354 -745
rect 583 -748 668 -747
rect 698 -748 1242 -747
rect 541 -750 584 -749
rect 513 -752 542 -751
rect 513 -754 563 -753
rect 562 -756 797 -755
rect 37 -767 52 -766
rect 58 -767 563 -766
rect 572 -767 1424 -766
rect 1430 -767 1585 -766
rect 1696 -767 1725 -766
rect 44 -769 433 -768
rect 485 -769 531 -768
rect 551 -769 738 -768
rect 793 -769 1193 -768
rect 1255 -769 1536 -768
rect 1549 -769 1578 -768
rect 44 -771 62 -770
rect 65 -771 346 -770
rect 366 -771 647 -770
rect 667 -771 717 -770
rect 737 -771 948 -770
rect 961 -771 1193 -770
rect 1353 -771 1431 -770
rect 1437 -771 1508 -770
rect 1528 -771 1571 -770
rect 65 -773 73 -772
rect 114 -773 360 -772
rect 366 -773 514 -772
rect 530 -773 549 -772
rect 558 -773 1039 -772
rect 1115 -773 1256 -772
rect 1262 -773 1354 -772
rect 1409 -773 1529 -772
rect 72 -775 94 -774
rect 124 -775 290 -774
rect 296 -775 556 -774
rect 607 -775 773 -774
rect 793 -775 878 -774
rect 905 -775 1438 -774
rect 1444 -775 1550 -774
rect 93 -777 185 -776
rect 187 -777 311 -776
rect 324 -777 360 -776
rect 380 -777 556 -776
rect 604 -777 906 -776
rect 908 -777 1326 -776
rect 1367 -777 1445 -776
rect 1458 -777 1515 -776
rect 135 -779 332 -778
rect 345 -779 353 -778
rect 380 -779 458 -778
rect 478 -779 514 -778
rect 534 -779 605 -778
rect 611 -779 678 -778
rect 684 -779 923 -778
rect 926 -779 1179 -778
rect 1220 -779 1263 -778
rect 1290 -779 1410 -778
rect 1416 -779 1501 -778
rect 135 -781 157 -780
rect 163 -781 332 -780
rect 394 -781 479 -780
rect 506 -781 829 -780
rect 835 -781 857 -780
rect 926 -781 990 -780
rect 1017 -781 1039 -780
rect 1115 -781 1242 -780
rect 1346 -781 1368 -780
rect 1374 -781 1417 -780
rect 1472 -781 1522 -780
rect 163 -783 783 -782
rect 796 -783 1102 -782
rect 1178 -783 1207 -782
rect 1213 -783 1221 -782
rect 1227 -783 1326 -782
rect 1479 -783 1560 -782
rect 117 -785 1214 -784
rect 1241 -785 1277 -784
rect 1311 -785 1480 -784
rect 1486 -785 1543 -784
rect 166 -787 675 -786
rect 688 -787 1046 -786
rect 1059 -787 1347 -786
rect 184 -789 1004 -788
rect 1024 -789 1375 -788
rect 191 -791 465 -790
rect 485 -791 836 -790
rect 849 -791 857 -790
rect 929 -791 1067 -790
rect 1094 -791 1207 -790
rect 1248 -791 1312 -790
rect 191 -793 549 -792
rect 569 -793 1067 -792
rect 1080 -793 1095 -792
rect 1199 -793 1277 -792
rect 205 -795 766 -794
rect 772 -795 808 -794
rect 828 -795 1494 -794
rect 208 -797 1228 -796
rect 1248 -797 1305 -796
rect 208 -799 724 -798
rect 751 -799 1004 -798
rect 1027 -799 1473 -798
rect 226 -801 311 -800
rect 352 -801 507 -800
rect 527 -801 1200 -800
rect 212 -803 227 -802
rect 240 -803 290 -802
rect 296 -803 493 -802
rect 534 -803 759 -802
rect 800 -803 1102 -802
rect 212 -805 437 -804
rect 457 -805 528 -804
rect 541 -805 1018 -804
rect 1045 -805 1088 -804
rect 233 -807 437 -806
rect 464 -807 472 -806
rect 576 -807 766 -806
rect 786 -807 801 -806
rect 807 -807 864 -806
rect 940 -807 948 -806
rect 961 -807 1340 -806
rect 121 -809 787 -808
rect 821 -809 941 -808
rect 975 -809 1025 -808
rect 1059 -809 1130 -808
rect 233 -811 412 -810
rect 415 -811 524 -810
rect 583 -811 612 -810
rect 632 -811 668 -810
rect 702 -811 724 -810
rect 814 -811 822 -810
rect 838 -811 1305 -810
rect 142 -813 524 -812
rect 583 -813 682 -812
rect 709 -813 759 -812
rect 814 -813 1459 -812
rect 142 -815 892 -814
rect 968 -815 976 -814
rect 982 -815 990 -814
rect 996 -815 1088 -814
rect 1122 -815 1130 -814
rect 79 -817 892 -816
rect 919 -817 997 -816
rect 1073 -817 1081 -816
rect 1122 -817 1137 -816
rect 79 -819 87 -818
rect 156 -819 682 -818
rect 716 -819 965 -818
rect 982 -819 1011 -818
rect 1052 -819 1074 -818
rect 1136 -819 1144 -818
rect 86 -821 101 -820
rect 240 -821 388 -820
rect 401 -821 577 -820
rect 590 -821 850 -820
rect 863 -821 885 -820
rect 933 -821 1011 -820
rect 1031 -821 1053 -820
rect 100 -823 444 -822
rect 509 -823 1340 -822
rect 152 -825 444 -824
rect 590 -825 640 -824
rect 646 -825 1466 -824
rect 149 -827 640 -826
rect 649 -827 1487 -826
rect 51 -829 150 -828
rect 261 -829 325 -828
rect 338 -829 388 -828
rect 401 -829 423 -828
rect 429 -829 720 -828
rect 744 -829 885 -828
rect 912 -829 934 -828
rect 1381 -829 1466 -828
rect 170 -831 339 -830
rect 373 -831 493 -830
rect 499 -831 745 -830
rect 838 -831 1403 -830
rect 170 -833 199 -832
rect 247 -833 262 -832
rect 282 -833 395 -832
rect 408 -833 563 -832
rect 625 -833 969 -832
rect 1283 -833 1382 -832
rect 121 -835 283 -834
rect 303 -835 416 -834
rect 422 -835 874 -834
rect 877 -835 1144 -834
rect 1269 -835 1284 -834
rect 1360 -835 1403 -834
rect 128 -837 248 -836
rect 268 -837 304 -836
rect 317 -837 430 -836
rect 499 -837 1291 -836
rect 128 -839 178 -838
rect 198 -839 206 -838
rect 268 -839 832 -838
rect 873 -839 1452 -838
rect 177 -841 276 -840
rect 317 -841 451 -840
rect 635 -841 710 -840
rect 831 -841 1396 -840
rect 107 -843 451 -842
rect 649 -843 703 -842
rect 880 -843 1396 -842
rect 107 -845 1424 -844
rect 254 -847 276 -846
rect 373 -847 731 -846
rect 898 -847 913 -846
rect 919 -847 1032 -846
rect 1164 -847 1361 -846
rect 1388 -847 1452 -846
rect 159 -849 899 -848
rect 1185 -849 1389 -848
rect 520 -851 1186 -850
rect 1234 -851 1270 -850
rect 520 -853 542 -852
rect 653 -853 731 -852
rect 870 -853 1165 -852
rect 1234 -853 1319 -852
rect 653 -855 675 -854
rect 691 -855 1319 -854
rect 660 -857 689 -856
rect 751 -857 871 -856
rect 660 -859 696 -858
rect 618 -861 696 -860
rect 597 -863 619 -862
rect 597 -865 843 -864
rect 779 -867 843 -866
rect 471 -869 780 -868
rect 30 -880 143 -879
rect 149 -880 892 -879
rect 919 -880 1452 -879
rect 1542 -880 1567 -879
rect 1570 -880 1627 -879
rect 1724 -880 1739 -879
rect 44 -882 629 -881
rect 656 -882 1571 -881
rect 1577 -882 1613 -881
rect 44 -884 52 -883
rect 79 -884 650 -883
rect 660 -884 832 -883
rect 838 -884 871 -883
rect 873 -884 1256 -883
rect 1318 -884 1634 -883
rect 51 -886 66 -885
rect 79 -886 129 -885
rect 135 -886 143 -885
rect 166 -886 1361 -885
rect 1521 -886 1543 -885
rect 1573 -886 1578 -885
rect 1584 -886 1620 -885
rect 65 -888 73 -887
rect 82 -888 234 -887
rect 257 -888 1438 -887
rect 1479 -888 1585 -887
rect 72 -890 87 -889
rect 93 -890 153 -889
rect 208 -890 353 -889
rect 408 -890 552 -889
rect 660 -890 857 -889
rect 880 -890 1529 -889
rect 58 -892 87 -891
rect 93 -892 570 -891
rect 667 -892 941 -891
rect 964 -892 1417 -891
rect 1437 -892 1445 -891
rect 1479 -892 1487 -891
rect 1493 -892 1522 -891
rect 58 -894 423 -893
rect 436 -894 643 -893
rect 667 -894 689 -893
rect 775 -894 1207 -893
rect 1346 -894 1557 -893
rect 100 -896 965 -895
rect 985 -896 1382 -895
rect 1388 -896 1445 -895
rect 1465 -896 1494 -895
rect 1514 -896 1529 -895
rect 100 -898 878 -897
rect 891 -898 955 -897
rect 961 -898 1557 -897
rect 107 -900 297 -899
rect 317 -900 321 -899
rect 338 -900 500 -899
rect 502 -900 969 -899
rect 992 -900 1452 -899
rect 1465 -900 1508 -899
rect 107 -902 213 -901
rect 219 -902 535 -901
rect 548 -902 591 -901
rect 674 -902 885 -901
rect 905 -902 920 -901
rect 926 -902 930 -901
rect 940 -902 1011 -901
rect 1069 -902 1550 -901
rect 110 -904 311 -903
rect 317 -904 325 -903
rect 352 -904 451 -903
rect 502 -904 1424 -903
rect 1472 -904 1515 -903
rect 1549 -904 1564 -903
rect 121 -906 367 -905
rect 408 -906 724 -905
rect 779 -906 843 -905
rect 856 -906 976 -905
rect 1111 -906 1487 -905
rect 1563 -906 1606 -905
rect 121 -908 125 -907
rect 128 -908 276 -907
rect 289 -908 297 -907
rect 310 -908 395 -907
rect 411 -908 923 -907
rect 926 -908 934 -907
rect 968 -908 990 -907
rect 1171 -908 1207 -907
rect 1248 -908 1382 -907
rect 1409 -908 1417 -907
rect 138 -910 381 -909
rect 394 -910 703 -909
rect 723 -910 759 -909
rect 782 -910 1396 -909
rect 163 -912 213 -911
rect 222 -912 255 -911
rect 268 -912 437 -911
rect 446 -912 871 -911
rect 877 -912 1193 -911
rect 1248 -912 1263 -911
rect 1290 -912 1347 -911
rect 1367 -912 1410 -911
rect 163 -914 178 -913
rect 191 -914 290 -913
rect 380 -914 773 -913
rect 828 -914 1361 -913
rect 1374 -914 1508 -913
rect 177 -916 388 -915
rect 450 -916 493 -915
rect 506 -916 1018 -915
rect 1164 -916 1193 -915
rect 1241 -916 1263 -915
rect 1269 -916 1291 -915
rect 1297 -916 1368 -915
rect 1395 -916 1431 -915
rect 191 -918 514 -917
rect 520 -918 1319 -917
rect 135 -920 514 -919
rect 523 -920 696 -919
rect 698 -920 955 -919
rect 975 -920 1256 -919
rect 1304 -920 1389 -919
rect 198 -922 423 -921
rect 425 -922 521 -921
rect 530 -922 1025 -921
rect 1115 -922 1298 -921
rect 198 -924 262 -923
rect 268 -924 304 -923
rect 387 -924 633 -923
rect 670 -924 829 -923
rect 845 -924 1375 -923
rect 205 -926 339 -925
rect 492 -926 685 -925
rect 688 -926 1312 -925
rect 205 -928 374 -927
rect 509 -928 517 -927
rect 534 -928 556 -927
rect 569 -928 619 -927
rect 625 -928 1424 -927
rect 184 -930 556 -929
rect 586 -930 1116 -929
rect 1157 -930 1165 -929
rect 1171 -930 1179 -929
rect 1227 -930 1270 -929
rect 1283 -930 1305 -929
rect 149 -932 185 -931
rect 226 -932 367 -931
rect 373 -932 402 -931
rect 506 -932 1284 -931
rect 233 -934 479 -933
rect 509 -934 528 -933
rect 590 -934 822 -933
rect 898 -934 906 -933
rect 933 -934 948 -933
rect 999 -934 1158 -933
rect 1234 -934 1242 -933
rect 250 -936 549 -935
rect 611 -936 633 -935
rect 674 -936 731 -935
rect 758 -936 787 -935
rect 898 -936 1354 -935
rect 254 -938 283 -937
rect 303 -938 416 -937
rect 478 -938 486 -937
rect 527 -938 815 -937
rect 835 -938 1354 -937
rect 170 -940 283 -939
rect 401 -940 430 -939
rect 485 -940 654 -939
rect 677 -940 1326 -939
rect 156 -942 171 -941
rect 261 -942 346 -941
rect 415 -942 542 -941
rect 604 -942 612 -941
rect 625 -942 650 -941
rect 684 -942 787 -941
rect 800 -942 815 -941
rect 901 -942 1312 -941
rect 1325 -942 1340 -941
rect 156 -944 248 -943
rect 275 -944 472 -943
rect 541 -944 563 -943
rect 695 -944 745 -943
rect 768 -944 1340 -943
rect 345 -946 360 -945
rect 429 -946 577 -945
rect 597 -946 745 -945
rect 772 -946 1592 -945
rect 114 -948 360 -947
rect 457 -948 605 -947
rect 702 -948 752 -947
rect 793 -948 801 -947
rect 1017 -948 1039 -947
rect 1150 -948 1179 -947
rect 1220 -948 1235 -947
rect 114 -950 241 -949
rect 443 -950 458 -949
rect 464 -950 472 -949
rect 562 -950 766 -949
rect 793 -950 808 -949
rect 1024 -950 1053 -949
rect 1108 -950 1221 -949
rect 37 -952 241 -951
rect 443 -952 1473 -951
rect 37 -954 864 -953
rect 929 -954 948 -953
rect 1038 -954 1095 -953
rect 1150 -954 1333 -953
rect 464 -956 1011 -955
rect 1052 -956 1102 -955
rect 1332 -956 1403 -955
rect 576 -958 738 -957
rect 765 -958 1599 -957
rect 583 -960 752 -959
rect 842 -960 1403 -959
rect 583 -962 850 -961
rect 1059 -962 1102 -961
rect 597 -964 1004 -963
rect 1031 -964 1060 -963
rect 1094 -964 1186 -963
rect 639 -966 1186 -965
rect 639 -968 1431 -967
rect 646 -970 864 -969
rect 982 -970 1004 -969
rect 1031 -970 1074 -969
rect 646 -972 1277 -971
rect 716 -974 822 -973
rect 849 -974 913 -973
rect 978 -974 1277 -973
rect 681 -976 913 -975
rect 982 -976 1214 -975
rect 226 -978 682 -977
rect 709 -978 717 -977
rect 730 -978 1228 -977
rect 499 -980 710 -979
rect 733 -980 836 -979
rect 1073 -980 1081 -979
rect 1199 -980 1214 -979
rect 737 -982 997 -981
rect 1045 -982 1200 -981
rect 996 -984 1536 -983
rect 653 -986 1536 -985
rect 1045 -988 1144 -987
rect 1080 -990 1088 -989
rect 1136 -990 1144 -989
rect 884 -992 1088 -991
rect 1122 -992 1137 -991
rect 1066 -994 1123 -993
rect 537 -996 1067 -995
rect 23 -1007 619 -1006
rect 628 -1007 724 -1006
rect 768 -1007 941 -1006
rect 961 -1007 1333 -1006
rect 1374 -1007 1567 -1006
rect 1570 -1007 1676 -1006
rect 1738 -1007 1746 -1006
rect 30 -1009 136 -1008
rect 149 -1009 206 -1008
rect 250 -1009 297 -1008
rect 310 -1009 517 -1008
rect 555 -1009 724 -1008
rect 786 -1009 902 -1008
rect 919 -1009 1385 -1008
rect 1528 -1009 1571 -1008
rect 1591 -1009 1683 -1008
rect 30 -1011 598 -1010
rect 611 -1011 657 -1010
rect 667 -1011 731 -1010
rect 786 -1011 801 -1010
rect 845 -1011 1200 -1010
rect 1241 -1011 1375 -1010
rect 1486 -1011 1529 -1010
rect 1535 -1011 1641 -1010
rect 37 -1013 696 -1012
rect 698 -1013 1592 -1012
rect 1626 -1013 1655 -1012
rect 44 -1015 76 -1014
rect 82 -1015 108 -1014
rect 114 -1015 216 -1014
rect 275 -1015 1000 -1014
rect 1010 -1015 1522 -1014
rect 1552 -1015 1613 -1014
rect 44 -1017 87 -1016
rect 89 -1017 409 -1016
rect 422 -1017 1606 -1016
rect 58 -1019 62 -1018
rect 72 -1019 87 -1018
rect 100 -1019 426 -1018
rect 485 -1019 612 -1018
rect 618 -1019 633 -1018
rect 684 -1019 1221 -1018
rect 1241 -1019 1298 -1018
rect 1360 -1019 1487 -1018
rect 1500 -1019 1536 -1018
rect 1556 -1019 1613 -1018
rect 51 -1021 73 -1020
rect 100 -1021 437 -1020
rect 492 -1021 776 -1020
rect 800 -1021 1249 -1020
rect 1297 -1021 1312 -1020
rect 1395 -1021 1501 -1020
rect 1563 -1021 1648 -1020
rect 51 -1023 122 -1022
rect 128 -1023 237 -1022
rect 268 -1023 409 -1022
rect 492 -1023 993 -1022
rect 996 -1023 1326 -1022
rect 1381 -1023 1396 -1022
rect 1423 -1023 1522 -1022
rect 1577 -1023 1627 -1022
rect 58 -1025 66 -1024
rect 107 -1025 482 -1024
rect 499 -1025 605 -1024
rect 632 -1025 703 -1024
rect 730 -1025 759 -1024
rect 835 -1025 997 -1024
rect 1003 -1025 1011 -1024
rect 1013 -1025 1032 -1024
rect 1108 -1025 1557 -1024
rect 1584 -1025 1606 -1024
rect 114 -1027 213 -1026
rect 275 -1027 843 -1026
rect 856 -1027 920 -1026
rect 933 -1027 962 -1026
rect 975 -1027 1067 -1026
rect 1111 -1027 1494 -1026
rect 1507 -1027 1585 -1026
rect 121 -1029 318 -1028
rect 324 -1029 510 -1028
rect 520 -1029 703 -1028
rect 733 -1029 1361 -1028
rect 1409 -1029 1424 -1028
rect 1430 -1029 1508 -1028
rect 1542 -1029 1578 -1028
rect 128 -1031 234 -1030
rect 282 -1031 444 -1030
rect 541 -1031 668 -1030
rect 688 -1031 1186 -1030
rect 1220 -1031 1256 -1030
rect 1318 -1031 1326 -1030
rect 1409 -1031 1438 -1030
rect 1444 -1031 1564 -1030
rect 138 -1033 486 -1032
rect 506 -1033 1319 -1032
rect 1416 -1033 1438 -1032
rect 1444 -1033 1452 -1032
rect 138 -1035 1473 -1034
rect 156 -1037 318 -1036
rect 331 -1037 503 -1036
rect 541 -1037 570 -1036
rect 576 -1037 696 -1036
rect 737 -1037 843 -1036
rect 863 -1037 888 -1036
rect 891 -1037 941 -1036
rect 954 -1037 1032 -1036
rect 1066 -1037 1102 -1036
rect 1115 -1037 1333 -1036
rect 1402 -1037 1417 -1036
rect 1472 -1037 1620 -1036
rect 156 -1039 388 -1038
rect 394 -1039 521 -1038
rect 548 -1039 556 -1038
rect 562 -1039 605 -1038
rect 660 -1039 759 -1038
rect 793 -1039 836 -1038
rect 866 -1039 1151 -1038
rect 1157 -1039 1312 -1038
rect 1388 -1039 1403 -1038
rect 1598 -1039 1620 -1038
rect 170 -1041 174 -1040
rect 177 -1041 269 -1040
rect 296 -1041 881 -1040
rect 891 -1041 1116 -1040
rect 1129 -1041 1133 -1040
rect 1157 -1041 1382 -1040
rect 1388 -1041 1476 -1040
rect 170 -1043 241 -1042
rect 310 -1043 398 -1042
rect 401 -1043 437 -1042
rect 457 -1043 507 -1042
rect 548 -1043 678 -1042
rect 691 -1043 773 -1042
rect 894 -1043 1081 -1042
rect 1090 -1043 1431 -1042
rect 177 -1045 213 -1044
rect 219 -1045 283 -1044
rect 331 -1045 451 -1044
rect 457 -1045 472 -1044
rect 562 -1045 1494 -1044
rect 184 -1047 206 -1046
rect 219 -1047 535 -1046
rect 569 -1047 675 -1046
rect 716 -1047 738 -1046
rect 870 -1047 1081 -1046
rect 1129 -1047 1165 -1046
rect 1185 -1047 1207 -1046
rect 1234 -1047 1249 -1046
rect 1255 -1047 1305 -1046
rect 142 -1049 185 -1048
rect 191 -1049 647 -1048
rect 660 -1049 804 -1048
rect 821 -1049 871 -1048
rect 877 -1049 1305 -1048
rect 142 -1051 647 -1050
rect 733 -1051 1599 -1050
rect 191 -1053 255 -1052
rect 338 -1053 388 -1052
rect 394 -1053 1354 -1052
rect 198 -1055 325 -1054
rect 352 -1055 622 -1054
rect 625 -1055 717 -1054
rect 744 -1055 822 -1054
rect 877 -1055 1200 -1054
rect 1206 -1055 1550 -1054
rect 163 -1057 199 -1056
rect 254 -1057 416 -1056
rect 446 -1057 626 -1056
rect 744 -1057 780 -1056
rect 912 -1057 1543 -1056
rect 163 -1059 381 -1058
rect 401 -1059 591 -1058
rect 597 -1059 1056 -1058
rect 1073 -1059 1102 -1058
rect 1227 -1059 1235 -1058
rect 1353 -1059 1368 -1058
rect 1465 -1059 1550 -1058
rect 261 -1061 353 -1060
rect 359 -1061 416 -1060
rect 450 -1061 650 -1060
rect 653 -1061 780 -1060
rect 926 -1061 955 -1060
rect 982 -1061 1109 -1060
rect 1213 -1061 1228 -1060
rect 1346 -1061 1368 -1060
rect 1465 -1061 1480 -1060
rect 359 -1063 888 -1062
rect 905 -1063 983 -1062
rect 985 -1063 1515 -1062
rect 373 -1065 444 -1064
rect 464 -1065 591 -1064
rect 649 -1065 927 -1064
rect 933 -1065 1018 -1064
rect 1024 -1065 1028 -1064
rect 1073 -1065 1137 -1064
rect 1171 -1065 1214 -1064
rect 1458 -1065 1515 -1064
rect 226 -1067 374 -1066
rect 380 -1067 430 -1066
rect 471 -1067 913 -1066
rect 968 -1067 1018 -1066
rect 1024 -1067 1039 -1066
rect 1136 -1067 1179 -1066
rect 226 -1069 304 -1068
rect 429 -1069 479 -1068
rect 534 -1069 699 -1068
rect 863 -1069 1480 -1068
rect 289 -1071 465 -1070
rect 576 -1071 1452 -1070
rect 289 -1073 528 -1072
rect 583 -1073 857 -1072
rect 905 -1073 1004 -1072
rect 1122 -1073 1179 -1072
rect 250 -1075 528 -1074
rect 586 -1075 794 -1074
rect 947 -1075 969 -1074
rect 989 -1075 1263 -1074
rect 303 -1077 766 -1076
rect 947 -1077 1053 -1076
rect 1132 -1077 1165 -1076
rect 1171 -1077 1193 -1076
rect 1262 -1077 1291 -1076
rect 131 -1079 766 -1078
rect 1045 -1079 1123 -1078
rect 1143 -1079 1193 -1078
rect 1283 -1079 1291 -1078
rect 338 -1081 990 -1080
rect 1045 -1081 1060 -1080
rect 1094 -1081 1144 -1080
rect 1276 -1081 1284 -1080
rect 513 -1083 584 -1082
rect 642 -1083 1459 -1082
rect 513 -1085 682 -1084
rect 828 -1085 1095 -1084
rect 79 -1087 682 -1086
rect 814 -1087 829 -1086
rect 978 -1087 1060 -1086
rect 79 -1089 94 -1088
rect 653 -1089 710 -1088
rect 807 -1089 815 -1088
rect 1006 -1089 1277 -1088
rect 93 -1091 640 -1090
rect 674 -1091 1347 -1090
rect 499 -1093 640 -1092
rect 709 -1093 899 -1092
rect 807 -1095 885 -1094
rect 898 -1095 1088 -1094
rect 1087 -1097 1151 -1096
rect 23 -1108 440 -1107
rect 471 -1108 703 -1107
rect 730 -1108 1242 -1107
rect 1255 -1108 1382 -1107
rect 1384 -1108 1627 -1107
rect 1640 -1108 1725 -1107
rect 1745 -1108 1760 -1107
rect 23 -1110 244 -1109
rect 275 -1110 479 -1109
rect 499 -1110 626 -1109
rect 649 -1110 745 -1109
rect 765 -1110 867 -1109
rect 887 -1110 1375 -1109
rect 1444 -1110 1662 -1109
rect 1675 -1110 1704 -1109
rect 37 -1112 213 -1111
rect 219 -1112 251 -1111
rect 275 -1112 304 -1111
rect 324 -1112 342 -1111
rect 401 -1112 678 -1111
rect 681 -1112 801 -1111
rect 817 -1112 1186 -1111
rect 1213 -1112 1382 -1111
rect 1444 -1112 1767 -1111
rect 72 -1114 542 -1113
rect 656 -1114 1347 -1113
rect 1451 -1114 1564 -1113
rect 1570 -1114 1718 -1113
rect 75 -1116 1676 -1115
rect 1682 -1116 1770 -1115
rect 89 -1118 514 -1117
rect 516 -1118 598 -1117
rect 681 -1118 773 -1117
rect 835 -1118 878 -1117
rect 929 -1118 1298 -1117
rect 1318 -1118 1452 -1117
rect 1465 -1118 1683 -1117
rect 93 -1120 545 -1119
rect 548 -1120 878 -1119
rect 933 -1120 1375 -1119
rect 1437 -1120 1564 -1119
rect 1570 -1120 1606 -1119
rect 1612 -1120 1753 -1119
rect 93 -1122 139 -1121
rect 173 -1122 668 -1121
rect 688 -1122 825 -1121
rect 859 -1122 899 -1121
rect 912 -1122 934 -1121
rect 950 -1122 1305 -1121
rect 1311 -1122 1438 -1121
rect 1479 -1122 1606 -1121
rect 1654 -1122 1781 -1121
rect 100 -1124 423 -1123
rect 506 -1124 731 -1123
rect 737 -1124 745 -1123
rect 758 -1124 913 -1123
rect 1045 -1124 1235 -1123
rect 1248 -1124 1613 -1123
rect 58 -1126 101 -1125
rect 107 -1126 234 -1125
rect 236 -1126 1473 -1125
rect 1493 -1126 1620 -1125
rect 58 -1128 171 -1127
rect 177 -1128 626 -1127
rect 653 -1128 773 -1127
rect 891 -1128 1312 -1127
rect 1332 -1128 1455 -1127
rect 1496 -1128 1648 -1127
rect 68 -1130 1249 -1129
rect 1290 -1130 1620 -1129
rect 89 -1132 1494 -1131
rect 1500 -1132 1641 -1131
rect 110 -1134 325 -1133
rect 380 -1134 549 -1133
rect 698 -1134 787 -1133
rect 891 -1134 1291 -1133
rect 1325 -1134 1501 -1133
rect 1507 -1134 1648 -1133
rect 121 -1136 398 -1135
rect 401 -1136 409 -1135
rect 415 -1136 636 -1135
rect 716 -1136 1214 -1135
rect 1220 -1136 1711 -1135
rect 121 -1138 1627 -1137
rect 128 -1140 136 -1139
rect 180 -1140 311 -1139
rect 380 -1140 570 -1139
rect 649 -1140 1221 -1139
rect 1325 -1140 1431 -1139
rect 1514 -1140 1669 -1139
rect 128 -1142 230 -1141
rect 233 -1142 430 -1141
rect 485 -1142 787 -1141
rect 919 -1142 1046 -1141
rect 1048 -1142 1200 -1141
rect 1339 -1142 1508 -1141
rect 1528 -1142 1690 -1141
rect 184 -1144 304 -1143
rect 387 -1144 409 -1143
rect 415 -1144 451 -1143
rect 492 -1144 717 -1143
rect 723 -1144 836 -1143
rect 968 -1144 1333 -1143
rect 1367 -1144 1515 -1143
rect 1549 -1144 1697 -1143
rect 79 -1146 388 -1145
rect 443 -1146 451 -1145
rect 499 -1146 738 -1145
rect 758 -1146 832 -1145
rect 1055 -1146 1354 -1145
rect 1402 -1146 1529 -1145
rect 1556 -1146 1739 -1145
rect 51 -1148 1354 -1147
rect 1409 -1148 1655 -1147
rect 51 -1150 598 -1149
rect 611 -1150 724 -1149
rect 765 -1150 885 -1149
rect 1055 -1150 1186 -1149
rect 1269 -1150 1368 -1149
rect 1416 -1150 1550 -1149
rect 1577 -1150 1732 -1149
rect 65 -1152 80 -1151
rect 124 -1152 969 -1151
rect 1066 -1152 1256 -1151
rect 1276 -1152 1403 -1151
rect 1416 -1152 1746 -1151
rect 65 -1154 1480 -1153
rect 1535 -1154 1557 -1153
rect 1577 -1154 1634 -1153
rect 142 -1156 493 -1155
rect 520 -1156 668 -1155
rect 768 -1156 843 -1155
rect 905 -1156 1270 -1155
rect 1283 -1156 1410 -1155
rect 1486 -1156 1634 -1155
rect 184 -1158 584 -1157
rect 779 -1158 1431 -1157
rect 1598 -1158 1788 -1157
rect 198 -1160 311 -1159
rect 338 -1160 843 -1159
rect 880 -1160 1284 -1159
rect 1388 -1160 1536 -1159
rect 198 -1162 255 -1161
rect 282 -1162 647 -1161
rect 793 -1162 920 -1161
rect 1003 -1162 1277 -1161
rect 1458 -1162 1599 -1161
rect 177 -1164 255 -1163
rect 261 -1164 1004 -1163
rect 1052 -1164 1487 -1163
rect 212 -1166 804 -1165
rect 821 -1166 906 -1165
rect 1066 -1166 1543 -1165
rect 219 -1168 265 -1167
rect 282 -1168 426 -1167
rect 443 -1168 696 -1167
rect 793 -1168 1074 -1167
rect 1087 -1168 1130 -1167
rect 1143 -1168 1389 -1167
rect 1458 -1168 1592 -1167
rect 226 -1170 640 -1169
rect 688 -1170 822 -1169
rect 961 -1170 1074 -1169
rect 1094 -1170 1347 -1169
rect 1521 -1170 1543 -1169
rect 1584 -1170 1592 -1169
rect 30 -1172 227 -1171
rect 247 -1172 486 -1171
rect 520 -1172 895 -1171
rect 996 -1172 1095 -1171
rect 1101 -1172 1200 -1171
rect 1395 -1172 1522 -1171
rect 30 -1174 87 -1173
rect 205 -1174 248 -1173
rect 296 -1174 430 -1173
rect 471 -1174 895 -1173
rect 1010 -1174 1130 -1173
rect 1150 -1174 1242 -1173
rect 86 -1176 164 -1175
rect 205 -1176 458 -1175
rect 527 -1176 612 -1175
rect 618 -1176 640 -1175
rect 695 -1176 1361 -1175
rect 149 -1178 164 -1177
rect 289 -1178 297 -1177
rect 338 -1178 437 -1177
rect 457 -1178 535 -1177
rect 569 -1178 710 -1177
rect 828 -1178 962 -1177
rect 982 -1178 1011 -1177
rect 1017 -1178 1088 -1177
rect 1101 -1178 1137 -1177
rect 1157 -1178 1235 -1177
rect 1360 -1178 1749 -1177
rect 145 -1180 150 -1179
rect 170 -1180 1137 -1179
rect 1164 -1180 1466 -1179
rect 268 -1182 437 -1181
rect 464 -1182 535 -1181
rect 562 -1182 710 -1181
rect 740 -1182 1165 -1181
rect 1171 -1182 1319 -1181
rect 142 -1184 269 -1183
rect 331 -1184 465 -1183
rect 562 -1184 675 -1183
rect 849 -1184 1018 -1183
rect 1038 -1184 1172 -1183
rect 1178 -1184 1340 -1183
rect 331 -1186 360 -1185
rect 576 -1186 780 -1185
rect 856 -1186 983 -1185
rect 1059 -1186 1144 -1185
rect 1178 -1186 1207 -1185
rect 1227 -1186 1396 -1185
rect 345 -1188 360 -1187
rect 555 -1188 577 -1187
rect 583 -1188 734 -1187
rect 751 -1188 850 -1187
rect 856 -1188 997 -1187
rect 1080 -1188 1207 -1187
rect 1227 -1188 1263 -1187
rect 345 -1190 482 -1189
rect 555 -1190 633 -1189
rect 674 -1190 808 -1189
rect 926 -1190 1060 -1189
rect 1108 -1190 1151 -1189
rect 1192 -1190 1585 -1189
rect 394 -1192 1081 -1191
rect 1115 -1192 1298 -1191
rect 352 -1194 395 -1193
rect 618 -1194 829 -1193
rect 898 -1194 927 -1193
rect 940 -1194 1039 -1193
rect 1122 -1194 1305 -1193
rect 352 -1196 374 -1195
rect 691 -1196 1109 -1195
rect 1262 -1196 1476 -1195
rect 317 -1198 374 -1197
rect 702 -1198 1116 -1197
rect 44 -1200 318 -1199
rect 751 -1200 864 -1199
rect 947 -1200 1158 -1199
rect 44 -1202 157 -1201
rect 541 -1202 864 -1201
rect 947 -1202 1025 -1201
rect 1031 -1202 1123 -1201
rect 156 -1204 591 -1203
rect 796 -1204 808 -1203
rect 954 -1204 1032 -1203
rect 590 -1206 661 -1205
rect 698 -1206 955 -1205
rect 975 -1206 1025 -1205
rect 604 -1208 661 -1207
rect 814 -1208 976 -1207
rect 989 -1208 1193 -1207
rect 527 -1210 605 -1209
rect 814 -1210 941 -1209
rect 870 -1212 990 -1211
rect 240 -1214 871 -1213
rect 240 -1216 290 -1215
rect 16 -1227 447 -1226
rect 506 -1227 864 -1226
rect 891 -1227 1088 -1226
rect 1094 -1227 1203 -1226
rect 1290 -1227 1294 -1226
rect 1311 -1227 1315 -1226
rect 1703 -1227 1749 -1226
rect 1766 -1227 1788 -1226
rect 44 -1229 265 -1228
rect 289 -1229 510 -1228
rect 548 -1229 566 -1228
rect 590 -1229 598 -1228
rect 607 -1229 1270 -1228
rect 1290 -1229 1305 -1228
rect 1311 -1229 1319 -1228
rect 1696 -1229 1704 -1228
rect 1745 -1229 1760 -1228
rect 44 -1231 90 -1230
rect 103 -1231 304 -1230
rect 345 -1231 797 -1230
rect 800 -1231 864 -1230
rect 894 -1231 1613 -1230
rect 1745 -1231 1777 -1230
rect 65 -1233 1354 -1232
rect 1612 -1233 1718 -1232
rect 54 -1235 66 -1234
rect 68 -1235 80 -1234
rect 107 -1235 115 -1234
rect 121 -1235 1375 -1234
rect 1717 -1235 1732 -1234
rect 72 -1237 654 -1236
rect 709 -1237 794 -1236
rect 817 -1237 962 -1236
rect 1010 -1237 1095 -1236
rect 1146 -1237 1466 -1236
rect 51 -1239 73 -1238
rect 110 -1239 661 -1238
rect 667 -1239 794 -1238
rect 821 -1239 1620 -1238
rect 114 -1241 941 -1240
rect 947 -1241 1536 -1240
rect 121 -1243 454 -1242
rect 551 -1243 1137 -1242
rect 1248 -1243 1270 -1242
rect 1314 -1243 1319 -1242
rect 1353 -1243 1480 -1242
rect 1486 -1243 1536 -1242
rect 124 -1245 479 -1244
rect 565 -1245 717 -1244
rect 737 -1245 745 -1244
rect 751 -1245 766 -1244
rect 779 -1245 801 -1244
rect 821 -1245 1543 -1244
rect 61 -1247 738 -1246
rect 740 -1247 1333 -1246
rect 1360 -1247 1375 -1246
rect 1458 -1247 1732 -1246
rect 145 -1249 1557 -1248
rect 170 -1251 178 -1250
rect 180 -1251 1739 -1250
rect 142 -1253 171 -1252
rect 177 -1253 199 -1252
rect 208 -1253 241 -1252
rect 243 -1253 1158 -1252
rect 1220 -1253 1249 -1252
rect 1325 -1253 1557 -1252
rect 142 -1255 213 -1254
rect 226 -1255 1004 -1254
rect 1010 -1255 1046 -1254
rect 1052 -1255 1585 -1254
rect 128 -1257 213 -1256
rect 226 -1257 255 -1256
rect 261 -1257 437 -1256
rect 443 -1257 1021 -1256
rect 1059 -1257 1158 -1256
rect 1171 -1257 1221 -1256
rect 1325 -1257 1770 -1256
rect 163 -1259 255 -1258
rect 292 -1259 871 -1258
rect 933 -1259 1060 -1258
rect 1087 -1259 1501 -1258
rect 1542 -1259 1550 -1258
rect 1584 -1259 1592 -1258
rect 163 -1261 706 -1260
rect 723 -1261 745 -1260
rect 751 -1261 769 -1260
rect 824 -1261 1056 -1260
rect 1101 -1261 1333 -1260
rect 1402 -1261 1459 -1260
rect 1465 -1261 1508 -1260
rect 1549 -1261 1599 -1260
rect 184 -1263 710 -1262
rect 740 -1263 1431 -1262
rect 1479 -1263 1641 -1262
rect 184 -1265 619 -1264
rect 632 -1265 1347 -1264
rect 1402 -1265 1445 -1264
rect 1486 -1265 1529 -1264
rect 1570 -1265 1592 -1264
rect 1598 -1265 1634 -1264
rect 1640 -1265 1655 -1264
rect 198 -1267 780 -1266
rect 828 -1267 1361 -1266
rect 1423 -1267 1508 -1266
rect 1528 -1267 1578 -1266
rect 1633 -1267 1648 -1266
rect 1654 -1267 1676 -1266
rect 296 -1269 605 -1268
rect 611 -1269 633 -1268
rect 639 -1269 661 -1268
rect 831 -1269 1256 -1268
rect 1339 -1269 1347 -1268
rect 1423 -1269 1515 -1268
rect 1577 -1269 1627 -1268
rect 1647 -1269 1669 -1268
rect 1675 -1269 1690 -1268
rect 58 -1271 605 -1270
rect 611 -1271 913 -1270
rect 922 -1271 1571 -1270
rect 1682 -1271 1690 -1270
rect 58 -1273 101 -1272
rect 296 -1273 353 -1272
rect 380 -1273 696 -1272
rect 702 -1273 1340 -1272
rect 1500 -1273 1522 -1272
rect 1682 -1273 1711 -1272
rect 205 -1275 353 -1274
rect 380 -1275 598 -1274
rect 600 -1275 640 -1274
rect 688 -1275 703 -1274
rect 831 -1275 1263 -1274
rect 1710 -1275 1725 -1274
rect 23 -1277 206 -1276
rect 303 -1277 332 -1276
rect 345 -1277 374 -1276
rect 387 -1277 591 -1276
rect 681 -1277 689 -1276
rect 835 -1277 892 -1276
rect 912 -1277 983 -1276
rect 996 -1277 1046 -1276
rect 1101 -1277 1473 -1276
rect 1724 -1277 1753 -1276
rect 23 -1279 542 -1278
rect 548 -1279 1256 -1278
rect 1752 -1279 1781 -1278
rect 310 -1281 717 -1280
rect 852 -1281 920 -1280
rect 929 -1281 1669 -1280
rect 156 -1283 311 -1282
rect 317 -1283 388 -1282
rect 415 -1283 507 -1282
rect 513 -1283 871 -1282
rect 933 -1283 1697 -1282
rect 149 -1285 157 -1284
rect 317 -1285 790 -1284
rect 856 -1285 1494 -1284
rect 100 -1287 1494 -1286
rect 149 -1289 878 -1288
rect 936 -1289 1298 -1288
rect 331 -1291 360 -1290
rect 366 -1291 542 -1290
rect 625 -1291 682 -1290
rect 807 -1291 878 -1290
rect 940 -1291 1007 -1290
rect 1017 -1291 1053 -1290
rect 1104 -1291 1620 -1290
rect 275 -1293 626 -1292
rect 667 -1293 983 -1292
rect 1038 -1293 1627 -1292
rect 135 -1295 276 -1294
rect 282 -1295 367 -1294
rect 373 -1295 465 -1294
rect 499 -1295 724 -1294
rect 772 -1295 808 -1294
rect 842 -1295 857 -1294
rect 859 -1295 1074 -1294
rect 1115 -1295 1739 -1294
rect 82 -1297 136 -1296
rect 187 -1297 500 -1296
rect 635 -1297 1039 -1296
rect 1108 -1297 1116 -1296
rect 1129 -1297 1137 -1296
rect 1150 -1297 1298 -1296
rect 191 -1299 465 -1298
rect 558 -1299 1130 -1298
rect 1143 -1299 1151 -1298
rect 1164 -1299 1172 -1298
rect 1192 -1299 1522 -1298
rect 191 -1301 976 -1300
rect 1031 -1301 1074 -1300
rect 1080 -1301 1109 -1300
rect 1164 -1301 1207 -1300
rect 1227 -1301 1473 -1300
rect 247 -1303 283 -1302
rect 338 -1303 416 -1302
rect 422 -1303 836 -1302
rect 950 -1303 1515 -1302
rect 173 -1305 339 -1304
rect 359 -1305 657 -1304
rect 674 -1305 773 -1304
rect 950 -1305 962 -1304
rect 989 -1305 1032 -1304
rect 1080 -1305 1186 -1304
rect 1206 -1305 1214 -1304
rect 1234 -1305 1431 -1304
rect 86 -1307 675 -1306
rect 695 -1307 1214 -1306
rect 1241 -1307 1263 -1306
rect 86 -1309 528 -1308
rect 562 -1309 1193 -1308
rect 247 -1311 269 -1310
rect 408 -1311 843 -1310
rect 926 -1311 1235 -1310
rect 222 -1313 269 -1312
rect 324 -1313 409 -1312
rect 422 -1313 755 -1312
rect 898 -1313 927 -1312
rect 954 -1313 990 -1312
rect 1003 -1313 1186 -1312
rect 324 -1315 969 -1314
rect 1024 -1315 1242 -1314
rect 436 -1317 759 -1316
rect 849 -1317 1025 -1316
rect 450 -1319 479 -1318
rect 485 -1319 563 -1318
rect 572 -1319 1228 -1318
rect 450 -1321 997 -1320
rect 457 -1323 514 -1322
rect 555 -1323 759 -1322
rect 884 -1323 969 -1322
rect 401 -1325 556 -1324
rect 583 -1325 899 -1324
rect 905 -1325 955 -1324
rect 394 -1327 402 -1326
rect 429 -1327 885 -1326
rect 219 -1329 430 -1328
rect 457 -1329 535 -1328
rect 618 -1329 850 -1328
rect 394 -1331 577 -1330
rect 698 -1331 976 -1330
rect 37 -1333 577 -1332
rect 786 -1333 906 -1332
rect 492 -1335 528 -1334
rect 534 -1335 815 -1334
rect 233 -1337 493 -1336
rect 520 -1337 584 -1336
rect 646 -1337 815 -1336
rect 30 -1339 234 -1338
rect 520 -1339 731 -1338
rect 786 -1339 1368 -1338
rect 30 -1341 570 -1340
rect 730 -1341 1067 -1340
rect 1367 -1341 1382 -1340
rect 485 -1343 570 -1342
rect 1066 -1343 1123 -1342
rect 1381 -1343 1389 -1342
rect 1122 -1345 1200 -1344
rect 1388 -1345 1396 -1344
rect 1199 -1347 1445 -1346
rect 1395 -1349 1410 -1348
rect 1409 -1351 1417 -1350
rect 1416 -1353 1438 -1352
rect 1437 -1355 1564 -1354
rect 1563 -1357 1606 -1356
rect 817 -1359 1606 -1358
rect 16 -1370 111 -1369
rect 121 -1370 209 -1369
rect 219 -1370 1039 -1369
rect 1048 -1370 1095 -1369
rect 1104 -1370 1690 -1369
rect 1738 -1370 1802 -1369
rect 51 -1372 94 -1371
rect 107 -1372 647 -1371
rect 719 -1372 1025 -1371
rect 1038 -1372 1109 -1371
rect 1146 -1372 1662 -1371
rect 1689 -1372 1697 -1371
rect 51 -1374 150 -1373
rect 159 -1374 178 -1373
rect 187 -1374 766 -1373
rect 814 -1374 1137 -1373
rect 1199 -1374 1347 -1373
rect 1591 -1374 1697 -1373
rect 58 -1376 619 -1375
rect 646 -1376 661 -1375
rect 751 -1376 1291 -1375
rect 1346 -1376 1396 -1375
rect 1591 -1376 1634 -1375
rect 65 -1378 80 -1377
rect 82 -1378 1375 -1377
rect 1395 -1378 1403 -1377
rect 1528 -1378 1634 -1377
rect 79 -1380 941 -1379
rect 978 -1380 1501 -1379
rect 1612 -1380 1662 -1379
rect 93 -1382 521 -1381
rect 551 -1382 836 -1381
rect 849 -1382 1326 -1381
rect 1374 -1382 1410 -1381
rect 1437 -1382 1529 -1381
rect 1612 -1382 1648 -1381
rect 124 -1384 717 -1383
rect 751 -1384 759 -1383
rect 761 -1384 1627 -1383
rect 1647 -1384 1683 -1383
rect 149 -1386 825 -1385
rect 831 -1386 1221 -1385
rect 1227 -1386 1410 -1385
rect 1500 -1386 1557 -1385
rect 1626 -1386 1676 -1385
rect 156 -1388 178 -1387
rect 194 -1388 283 -1387
rect 289 -1388 472 -1387
rect 478 -1388 517 -1387
rect 520 -1388 1032 -1387
rect 1034 -1388 1683 -1387
rect 103 -1390 1032 -1389
rect 1066 -1390 1095 -1389
rect 1108 -1390 1249 -1389
rect 1402 -1390 1588 -1389
rect 156 -1392 293 -1391
rect 317 -1392 619 -1391
rect 625 -1392 661 -1391
rect 758 -1392 1326 -1391
rect 1556 -1392 1564 -1391
rect 170 -1394 206 -1393
rect 219 -1394 311 -1393
rect 324 -1394 671 -1393
rect 786 -1394 1137 -1393
rect 1202 -1394 1704 -1393
rect 114 -1396 206 -1395
rect 222 -1396 1340 -1395
rect 1563 -1396 1669 -1395
rect 114 -1398 717 -1397
rect 789 -1398 941 -1397
rect 982 -1398 1732 -1397
rect 170 -1400 640 -1399
rect 817 -1400 1221 -1399
rect 1227 -1400 1256 -1399
rect 1339 -1400 1382 -1399
rect 1584 -1400 1669 -1399
rect 1731 -1400 1746 -1399
rect 163 -1402 640 -1401
rect 821 -1402 1333 -1401
rect 1381 -1402 1431 -1401
rect 1584 -1402 1704 -1401
rect 163 -1404 255 -1403
rect 257 -1404 612 -1403
rect 849 -1404 892 -1403
rect 919 -1404 1609 -1403
rect 198 -1406 542 -1405
rect 555 -1406 906 -1405
rect 919 -1406 927 -1405
rect 982 -1406 997 -1405
rect 1003 -1406 1214 -1405
rect 1216 -1406 1508 -1405
rect 54 -1408 997 -1407
rect 1006 -1408 1473 -1407
rect 1507 -1408 1599 -1407
rect 135 -1410 199 -1409
rect 201 -1410 1438 -1409
rect 1472 -1410 1606 -1409
rect 135 -1412 143 -1411
rect 226 -1412 283 -1411
rect 310 -1412 458 -1411
rect 471 -1412 486 -1411
rect 506 -1412 556 -1411
rect 558 -1412 1571 -1411
rect 1598 -1412 1725 -1411
rect 142 -1414 213 -1413
rect 229 -1414 304 -1413
rect 366 -1414 486 -1413
rect 541 -1414 934 -1413
rect 1010 -1414 1025 -1413
rect 1066 -1414 1116 -1413
rect 1157 -1414 1606 -1413
rect 191 -1416 213 -1415
rect 215 -1416 367 -1415
rect 380 -1416 507 -1415
rect 562 -1416 836 -1415
rect 891 -1416 955 -1415
rect 1010 -1416 1060 -1415
rect 1115 -1416 1151 -1415
rect 1157 -1416 1193 -1415
rect 1213 -1416 1263 -1415
rect 1332 -1416 1536 -1415
rect 37 -1418 192 -1417
rect 240 -1418 325 -1417
rect 380 -1418 514 -1417
rect 562 -1418 682 -1417
rect 730 -1418 927 -1417
rect 933 -1418 1291 -1417
rect 1318 -1418 1536 -1417
rect 86 -1420 731 -1419
rect 922 -1420 1235 -1419
rect 1248 -1420 1277 -1419
rect 1318 -1420 1417 -1419
rect 1430 -1420 1452 -1419
rect 1479 -1420 1571 -1419
rect 86 -1422 794 -1421
rect 950 -1422 1452 -1421
rect 1479 -1422 1655 -1421
rect 254 -1424 304 -1423
rect 387 -1424 815 -1423
rect 954 -1424 969 -1423
rect 1017 -1424 1676 -1423
rect 61 -1426 388 -1425
rect 408 -1426 766 -1425
rect 793 -1426 801 -1425
rect 968 -1426 1046 -1425
rect 1059 -1426 1130 -1425
rect 1192 -1426 1270 -1425
rect 1276 -1426 1578 -1425
rect 268 -1428 1102 -1427
rect 1129 -1428 1172 -1427
rect 1255 -1428 1298 -1427
rect 1416 -1428 1515 -1427
rect 1538 -1428 1655 -1427
rect 268 -1430 297 -1429
rect 408 -1430 605 -1429
rect 611 -1430 741 -1429
rect 1017 -1430 1074 -1429
rect 1080 -1430 1151 -1429
rect 1171 -1430 1207 -1429
rect 1262 -1430 1305 -1429
rect 1577 -1430 1620 -1429
rect 184 -1432 1620 -1431
rect 275 -1434 482 -1433
rect 499 -1434 801 -1433
rect 975 -1434 1074 -1433
rect 1143 -1434 1515 -1433
rect 275 -1436 829 -1435
rect 1020 -1436 1123 -1435
rect 1143 -1436 1179 -1435
rect 1297 -1436 1494 -1435
rect 296 -1438 465 -1437
rect 478 -1438 1207 -1437
rect 1304 -1438 1354 -1437
rect 1360 -1438 1494 -1437
rect 44 -1440 465 -1439
rect 499 -1440 535 -1439
rect 569 -1440 1053 -1439
rect 1178 -1440 1186 -1439
rect 1353 -1440 1445 -1439
rect 44 -1442 73 -1441
rect 415 -1442 573 -1441
rect 597 -1442 738 -1441
rect 779 -1442 1081 -1441
rect 1185 -1442 1312 -1441
rect 1360 -1442 1466 -1441
rect 72 -1444 227 -1443
rect 240 -1444 738 -1443
rect 1045 -1444 1459 -1443
rect 1465 -1444 1641 -1443
rect 247 -1446 416 -1445
rect 436 -1446 948 -1445
rect 1052 -1446 1242 -1445
rect 1444 -1446 1487 -1445
rect 247 -1448 339 -1447
rect 436 -1448 937 -1447
rect 947 -1448 1718 -1447
rect 261 -1450 339 -1449
rect 450 -1450 668 -1449
rect 674 -1450 1725 -1449
rect 261 -1452 332 -1451
rect 453 -1452 843 -1451
rect 1241 -1452 1284 -1451
rect 1458 -1452 1543 -1451
rect 1710 -1452 1718 -1451
rect 233 -1454 843 -1453
rect 1283 -1454 1368 -1453
rect 1486 -1454 1522 -1453
rect 1542 -1454 1550 -1453
rect 1643 -1454 1711 -1453
rect 233 -1456 423 -1455
rect 457 -1456 906 -1455
rect 1367 -1456 1424 -1455
rect 1549 -1456 1753 -1455
rect 331 -1458 549 -1457
rect 569 -1458 591 -1457
rect 604 -1458 871 -1457
rect 1388 -1458 1424 -1457
rect 422 -1460 937 -1459
rect 460 -1462 1235 -1461
rect 513 -1464 1270 -1463
rect 527 -1466 598 -1465
rect 653 -1466 675 -1465
rect 681 -1466 808 -1465
rect 852 -1466 1522 -1465
rect 373 -1468 528 -1467
rect 534 -1468 825 -1467
rect 870 -1468 878 -1467
rect 373 -1470 493 -1469
rect 548 -1470 951 -1469
rect 30 -1472 493 -1471
rect 576 -1472 780 -1471
rect 877 -1472 885 -1471
rect 30 -1474 132 -1473
rect 576 -1474 633 -1473
rect 653 -1474 1088 -1473
rect 131 -1476 584 -1475
rect 590 -1476 986 -1475
rect 394 -1478 584 -1477
rect 632 -1478 990 -1477
rect 394 -1480 430 -1479
rect 443 -1480 1088 -1479
rect 359 -1482 430 -1481
rect 443 -1482 703 -1481
rect 726 -1482 1123 -1481
rect 352 -1484 360 -1483
rect 695 -1484 1102 -1483
rect 352 -1486 402 -1485
rect 695 -1486 724 -1485
rect 740 -1486 1389 -1485
rect 345 -1488 402 -1487
rect 702 -1488 829 -1487
rect 884 -1488 899 -1487
rect 912 -1488 990 -1487
rect 23 -1490 346 -1489
rect 754 -1490 808 -1489
rect 856 -1490 899 -1489
rect 912 -1490 962 -1489
rect 23 -1492 129 -1491
rect 856 -1492 864 -1491
rect 961 -1492 1553 -1491
rect 128 -1494 1312 -1493
rect 772 -1496 864 -1495
rect 709 -1498 773 -1497
rect 709 -1500 867 -1499
rect 23 -1511 230 -1510
rect 240 -1511 321 -1510
rect 373 -1511 377 -1510
rect 401 -1511 458 -1510
rect 460 -1511 1228 -1510
rect 1451 -1511 1455 -1510
rect 1521 -1511 1550 -1510
rect 1584 -1511 1669 -1510
rect 1706 -1511 1711 -1510
rect 1801 -1511 1823 -1510
rect 23 -1513 419 -1512
rect 436 -1513 762 -1512
rect 779 -1513 829 -1512
rect 866 -1513 1424 -1512
rect 1451 -1513 1473 -1512
rect 1521 -1513 1606 -1512
rect 1640 -1513 1732 -1512
rect 37 -1515 727 -1514
rect 737 -1515 1221 -1514
rect 1227 -1515 1256 -1514
rect 1304 -1515 1424 -1514
rect 1535 -1515 1697 -1514
rect 37 -1517 66 -1516
rect 93 -1517 318 -1516
rect 373 -1517 486 -1516
rect 492 -1517 671 -1516
rect 681 -1517 979 -1516
rect 1020 -1517 1466 -1516
rect 1535 -1517 1543 -1516
rect 1577 -1517 1585 -1516
rect 1598 -1517 1697 -1516
rect 51 -1519 626 -1518
rect 688 -1519 951 -1518
rect 1031 -1519 1200 -1518
rect 1255 -1519 1263 -1518
rect 1454 -1519 1473 -1518
rect 1507 -1519 1543 -1518
rect 1577 -1519 1613 -1518
rect 1640 -1519 1648 -1518
rect 1650 -1519 1725 -1518
rect 51 -1521 262 -1520
rect 264 -1521 521 -1520
rect 527 -1521 657 -1520
rect 716 -1521 1263 -1520
rect 1311 -1521 1508 -1520
rect 1591 -1521 1599 -1520
rect 1612 -1521 1627 -1520
rect 1643 -1521 1711 -1520
rect 1717 -1521 1725 -1520
rect 58 -1523 958 -1522
rect 989 -1523 1032 -1522
rect 1034 -1523 1109 -1522
rect 1157 -1523 1200 -1522
rect 1311 -1523 1319 -1522
rect 1479 -1523 1592 -1522
rect 1668 -1523 1683 -1522
rect 1703 -1523 1718 -1522
rect 65 -1525 871 -1524
rect 880 -1525 1018 -1524
rect 1045 -1525 1067 -1524
rect 1188 -1525 1459 -1524
rect 1514 -1525 1627 -1524
rect 1633 -1525 1683 -1524
rect 93 -1527 542 -1526
rect 607 -1527 920 -1526
rect 936 -1527 1186 -1526
rect 1192 -1527 1221 -1526
rect 1318 -1527 1648 -1526
rect 124 -1529 314 -1528
rect 380 -1529 458 -1528
rect 481 -1529 1609 -1528
rect 44 -1531 125 -1530
rect 128 -1531 199 -1530
rect 212 -1531 241 -1530
rect 310 -1531 727 -1530
rect 737 -1531 745 -1530
rect 747 -1531 934 -1530
rect 947 -1531 1235 -1530
rect 1332 -1531 1515 -1530
rect 1563 -1531 1634 -1530
rect 44 -1533 62 -1532
rect 79 -1533 129 -1532
rect 131 -1533 297 -1532
rect 415 -1533 570 -1532
rect 611 -1533 682 -1532
rect 702 -1533 717 -1532
rect 723 -1533 1361 -1532
rect 1416 -1533 1480 -1532
rect 1556 -1533 1564 -1532
rect 79 -1535 1007 -1534
rect 1048 -1535 1284 -1534
rect 1325 -1535 1333 -1534
rect 1395 -1535 1417 -1534
rect 1430 -1535 1459 -1534
rect 1556 -1535 1571 -1534
rect 149 -1537 612 -1536
rect 625 -1537 822 -1536
rect 831 -1537 1606 -1536
rect 135 -1539 150 -1538
rect 156 -1539 1550 -1538
rect 159 -1541 381 -1540
rect 415 -1541 472 -1540
rect 506 -1541 528 -1540
rect 569 -1541 1655 -1540
rect 184 -1543 444 -1542
rect 506 -1543 556 -1542
rect 604 -1543 703 -1542
rect 709 -1543 1067 -1542
rect 1073 -1543 1193 -1542
rect 1206 -1543 1284 -1542
rect 1290 -1543 1326 -1542
rect 1381 -1543 1396 -1542
rect 1493 -1543 1571 -1542
rect 1654 -1543 1662 -1542
rect 184 -1545 1431 -1544
rect 1661 -1545 1676 -1544
rect 191 -1547 402 -1546
rect 422 -1547 521 -1546
rect 544 -1547 1382 -1546
rect 1675 -1547 1690 -1546
rect 86 -1549 423 -1548
rect 436 -1549 997 -1548
rect 1059 -1549 1074 -1548
rect 1164 -1549 1235 -1548
rect 1269 -1549 1291 -1548
rect 1685 -1549 1690 -1548
rect 68 -1551 87 -1550
rect 191 -1551 248 -1550
rect 387 -1551 472 -1550
rect 478 -1551 1494 -1550
rect 194 -1553 1466 -1552
rect 198 -1555 451 -1554
rect 653 -1555 920 -1554
rect 947 -1555 1539 -1554
rect 205 -1557 934 -1556
rect 968 -1557 990 -1556
rect 996 -1557 1123 -1556
rect 1178 -1557 1270 -1556
rect 121 -1559 206 -1558
rect 212 -1559 325 -1558
rect 387 -1559 465 -1558
rect 541 -1559 1123 -1558
rect 1136 -1559 1179 -1558
rect 1185 -1559 1305 -1558
rect 121 -1561 157 -1560
rect 215 -1561 409 -1560
rect 443 -1561 563 -1560
rect 632 -1561 969 -1560
rect 1062 -1561 1445 -1560
rect 219 -1563 689 -1562
rect 709 -1563 836 -1562
rect 863 -1563 1361 -1562
rect 1367 -1563 1445 -1562
rect 30 -1565 220 -1564
rect 222 -1565 734 -1564
rect 740 -1565 1102 -1564
rect 1136 -1565 1144 -1564
rect 1346 -1565 1368 -1564
rect 30 -1567 629 -1566
rect 653 -1567 675 -1566
rect 754 -1567 1053 -1566
rect 1101 -1567 1151 -1566
rect 1346 -1567 1403 -1566
rect 233 -1569 297 -1568
rect 324 -1569 818 -1568
rect 863 -1569 1158 -1568
rect 1388 -1569 1403 -1568
rect 233 -1571 430 -1570
rect 446 -1571 479 -1570
rect 499 -1571 633 -1570
rect 667 -1571 1165 -1570
rect 1388 -1571 1501 -1570
rect 247 -1573 311 -1572
rect 429 -1573 822 -1572
rect 870 -1573 1004 -1572
rect 1094 -1573 1151 -1572
rect 1409 -1573 1501 -1572
rect 275 -1575 409 -1574
rect 464 -1575 605 -1574
rect 758 -1575 857 -1574
rect 894 -1575 1242 -1574
rect 1353 -1575 1410 -1574
rect 142 -1577 276 -1576
rect 499 -1577 640 -1576
rect 730 -1577 759 -1576
rect 779 -1577 1018 -1576
rect 1094 -1577 1130 -1576
rect 1297 -1577 1354 -1576
rect 142 -1579 164 -1578
rect 548 -1579 668 -1578
rect 730 -1579 1340 -1578
rect 163 -1581 1242 -1580
rect 1297 -1581 1340 -1580
rect 548 -1583 584 -1582
rect 590 -1583 675 -1582
rect 786 -1583 927 -1582
rect 940 -1583 1004 -1582
rect 1115 -1583 1130 -1582
rect 187 -1585 591 -1584
rect 639 -1585 892 -1584
rect 912 -1585 927 -1584
rect 940 -1585 1081 -1584
rect 1087 -1585 1116 -1584
rect 1125 -1585 1144 -1584
rect 492 -1587 892 -1586
rect 898 -1587 913 -1586
rect 975 -1587 1053 -1586
rect 1080 -1587 1207 -1586
rect 562 -1589 577 -1588
rect 583 -1589 661 -1588
rect 786 -1589 825 -1588
rect 884 -1589 899 -1588
rect 954 -1589 976 -1588
rect 1024 -1589 1088 -1588
rect 135 -1591 825 -1590
rect 849 -1591 885 -1590
rect 954 -1591 1277 -1590
rect 450 -1593 850 -1592
rect 1010 -1593 1025 -1592
rect 1213 -1593 1277 -1592
rect 551 -1595 1214 -1594
rect 576 -1597 766 -1596
rect 789 -1597 843 -1596
rect 982 -1597 1011 -1596
rect 597 -1599 661 -1598
rect 800 -1599 836 -1598
rect 982 -1599 1039 -1598
rect 72 -1601 1039 -1600
rect 72 -1603 255 -1602
rect 618 -1603 766 -1602
rect 793 -1603 801 -1602
rect 807 -1603 867 -1602
rect 100 -1605 619 -1604
rect 772 -1605 794 -1604
rect 814 -1605 843 -1604
rect 100 -1607 227 -1606
rect 513 -1607 808 -1606
rect 114 -1609 227 -1608
rect 359 -1609 514 -1608
rect 555 -1609 815 -1608
rect 114 -1611 332 -1610
rect 359 -1611 367 -1610
rect 751 -1611 773 -1610
rect 166 -1613 255 -1612
rect 366 -1613 752 -1612
rect 170 -1615 598 -1614
rect 170 -1617 290 -1616
rect 107 -1619 290 -1618
rect 107 -1621 395 -1620
rect 268 -1623 395 -1622
rect 268 -1625 283 -1624
rect 282 -1627 339 -1626
rect 338 -1629 346 -1628
rect 345 -1631 535 -1630
rect 534 -1633 878 -1632
rect 331 -1635 878 -1634
rect 30 -1646 311 -1645
rect 324 -1646 384 -1645
rect 387 -1646 608 -1645
rect 660 -1646 734 -1645
rect 789 -1646 1298 -1645
rect 1300 -1646 1459 -1645
rect 1549 -1646 1704 -1645
rect 1822 -1646 1840 -1645
rect 30 -1648 199 -1647
rect 219 -1648 503 -1647
rect 548 -1648 1711 -1647
rect 23 -1650 199 -1649
rect 236 -1650 1795 -1649
rect 23 -1652 234 -1651
rect 275 -1652 311 -1651
rect 352 -1652 451 -1651
rect 551 -1652 1116 -1651
rect 1122 -1652 1459 -1651
rect 1598 -1652 1732 -1651
rect 58 -1654 731 -1653
rect 800 -1654 818 -1653
rect 856 -1654 885 -1653
rect 891 -1654 1788 -1653
rect 107 -1656 892 -1655
rect 954 -1656 1112 -1655
rect 1125 -1656 1256 -1655
rect 1423 -1656 1550 -1655
rect 1605 -1656 1746 -1655
rect 93 -1658 108 -1657
rect 121 -1658 1172 -1657
rect 1185 -1658 1837 -1657
rect 93 -1660 538 -1659
rect 576 -1660 801 -1659
rect 814 -1660 1641 -1659
rect 1647 -1660 1781 -1659
rect 121 -1662 720 -1661
rect 782 -1662 1606 -1661
rect 1619 -1662 1753 -1661
rect 124 -1664 888 -1663
rect 957 -1664 1739 -1663
rect 135 -1666 678 -1665
rect 681 -1666 752 -1665
rect 835 -1666 1172 -1665
rect 1185 -1666 1235 -1665
rect 1304 -1666 1424 -1665
rect 1451 -1666 1711 -1665
rect 135 -1668 1063 -1667
rect 1066 -1668 1084 -1667
rect 1101 -1668 1256 -1667
rect 1332 -1668 1452 -1667
rect 1479 -1668 1620 -1667
rect 1626 -1668 1760 -1667
rect 159 -1670 580 -1669
rect 590 -1670 752 -1669
rect 835 -1670 850 -1669
rect 859 -1670 997 -1669
rect 1003 -1670 1564 -1669
rect 1633 -1670 1767 -1669
rect 184 -1672 213 -1671
rect 275 -1672 521 -1671
rect 604 -1672 727 -1671
rect 863 -1672 1088 -1671
rect 1101 -1672 1690 -1671
rect 1696 -1672 1830 -1671
rect 145 -1674 185 -1673
rect 187 -1674 535 -1673
rect 611 -1674 661 -1673
rect 674 -1674 815 -1673
rect 828 -1674 864 -1673
rect 877 -1674 1361 -1673
rect 1374 -1674 1480 -1673
rect 1521 -1674 1641 -1673
rect 1650 -1674 1725 -1673
rect 44 -1676 675 -1675
rect 681 -1676 780 -1675
rect 786 -1676 829 -1675
rect 877 -1676 906 -1675
rect 950 -1676 1634 -1675
rect 1654 -1676 1809 -1675
rect 44 -1678 640 -1677
rect 716 -1678 731 -1677
rect 779 -1678 825 -1677
rect 880 -1678 1326 -1677
rect 1395 -1678 1522 -1677
rect 1528 -1678 1690 -1677
rect 212 -1680 556 -1679
rect 611 -1680 843 -1679
rect 901 -1680 997 -1679
rect 1017 -1680 1130 -1679
rect 1146 -1680 1578 -1679
rect 1584 -1680 1725 -1679
rect 303 -1682 325 -1681
rect 352 -1682 545 -1681
rect 618 -1682 906 -1681
rect 947 -1682 1018 -1681
rect 1020 -1682 1235 -1681
rect 1262 -1682 1326 -1681
rect 1402 -1682 1529 -1681
rect 1542 -1682 1697 -1681
rect 205 -1684 1403 -1683
rect 1416 -1684 1543 -1683
rect 1661 -1684 1802 -1683
rect 37 -1686 1662 -1685
rect 1668 -1686 1816 -1685
rect 37 -1688 507 -1687
rect 534 -1688 1088 -1687
rect 1108 -1688 1592 -1687
rect 1675 -1688 1823 -1687
rect 79 -1690 206 -1689
rect 254 -1690 304 -1689
rect 331 -1690 619 -1689
rect 639 -1690 647 -1689
rect 716 -1690 1032 -1689
rect 1038 -1690 1599 -1689
rect 1682 -1690 1718 -1689
rect 79 -1692 367 -1691
rect 387 -1692 493 -1691
rect 499 -1692 521 -1691
rect 646 -1692 654 -1691
rect 723 -1692 1067 -1691
rect 1080 -1692 1417 -1691
rect 1437 -1692 1564 -1691
rect 1570 -1692 1592 -1691
rect 254 -1694 465 -1693
rect 485 -1694 545 -1693
rect 632 -1694 654 -1693
rect 747 -1694 1396 -1693
rect 1444 -1694 1585 -1693
rect 331 -1696 360 -1695
rect 362 -1696 1004 -1695
rect 1010 -1696 1081 -1695
rect 1129 -1696 1249 -1695
rect 1269 -1696 1333 -1695
rect 1388 -1696 1676 -1695
rect 366 -1698 381 -1697
rect 394 -1698 594 -1697
rect 807 -1698 843 -1697
rect 975 -1698 1032 -1697
rect 1038 -1698 1060 -1697
rect 1136 -1698 1270 -1697
rect 1290 -1698 1389 -1697
rect 1472 -1698 1627 -1697
rect 394 -1700 598 -1699
rect 754 -1700 1137 -1699
rect 1157 -1700 1445 -1699
rect 1493 -1700 1655 -1699
rect 401 -1702 598 -1701
rect 726 -1702 1494 -1701
rect 1500 -1702 1578 -1701
rect 240 -1704 402 -1703
rect 408 -1704 552 -1703
rect 765 -1704 808 -1703
rect 824 -1704 969 -1703
rect 978 -1704 1648 -1703
rect 114 -1706 241 -1705
rect 408 -1706 885 -1705
rect 898 -1706 969 -1705
rect 989 -1706 1109 -1705
rect 1157 -1706 1319 -1705
rect 1339 -1706 1473 -1705
rect 1507 -1706 1571 -1705
rect 415 -1708 451 -1707
rect 457 -1708 493 -1707
rect 506 -1708 542 -1707
rect 758 -1708 766 -1707
rect 919 -1708 990 -1707
rect 1010 -1708 1144 -1707
rect 1164 -1708 1249 -1707
rect 1276 -1708 1340 -1707
rect 1381 -1708 1501 -1707
rect 1514 -1708 1669 -1707
rect 219 -1710 1515 -1709
rect 1535 -1710 1683 -1709
rect 415 -1712 577 -1711
rect 635 -1712 1382 -1711
rect 1409 -1712 1536 -1711
rect 1556 -1712 1718 -1711
rect 429 -1714 1305 -1713
rect 1311 -1714 1508 -1713
rect 436 -1716 745 -1715
rect 758 -1716 773 -1715
rect 786 -1716 1277 -1715
rect 1430 -1716 1557 -1715
rect 114 -1718 773 -1717
rect 849 -1718 1144 -1717
rect 1178 -1718 1312 -1717
rect 1367 -1718 1431 -1717
rect 436 -1720 570 -1719
rect 695 -1720 745 -1719
rect 870 -1720 920 -1719
rect 933 -1720 1060 -1719
rect 1206 -1720 1613 -1719
rect 89 -1722 1207 -1721
rect 1220 -1722 1319 -1721
rect 1353 -1722 1613 -1721
rect 446 -1724 514 -1723
rect 541 -1724 556 -1723
rect 562 -1724 570 -1723
rect 695 -1724 794 -1723
rect 870 -1724 948 -1723
rect 1006 -1724 1410 -1723
rect 317 -1726 794 -1725
rect 933 -1726 962 -1725
rect 1024 -1726 1375 -1725
rect 268 -1728 1025 -1727
rect 1027 -1728 1123 -1727
rect 1227 -1728 1368 -1727
rect 268 -1730 549 -1729
rect 562 -1730 899 -1729
rect 940 -1730 1179 -1729
rect 1241 -1730 1263 -1729
rect 1283 -1730 1354 -1729
rect 100 -1732 1242 -1731
rect 100 -1734 171 -1733
rect 261 -1734 941 -1733
rect 1045 -1734 1165 -1733
rect 1213 -1734 1284 -1733
rect 317 -1736 1210 -1735
rect 453 -1738 1221 -1737
rect 457 -1740 479 -1739
rect 485 -1740 528 -1739
rect 1045 -1740 1200 -1739
rect 163 -1742 1200 -1741
rect 163 -1744 192 -1743
rect 289 -1744 528 -1743
rect 1052 -1744 1116 -1743
rect 1150 -1744 1214 -1743
rect 156 -1746 192 -1745
rect 222 -1746 290 -1745
rect 464 -1746 472 -1745
rect 478 -1746 584 -1745
rect 982 -1746 1151 -1745
rect 156 -1748 430 -1747
rect 471 -1748 626 -1747
rect 912 -1748 983 -1747
rect 1052 -1748 1487 -1747
rect 170 -1750 223 -1749
rect 499 -1750 962 -1749
rect 1055 -1750 1361 -1749
rect 1465 -1750 1487 -1749
rect 513 -1752 668 -1751
rect 702 -1752 913 -1751
rect 1094 -1752 1228 -1751
rect 1346 -1752 1466 -1751
rect 296 -1754 1095 -1753
rect 1192 -1754 1347 -1753
rect 226 -1756 297 -1755
rect 422 -1756 703 -1755
rect 1073 -1756 1193 -1755
rect 51 -1758 227 -1757
rect 422 -1758 738 -1757
rect 51 -1760 927 -1759
rect 65 -1762 927 -1761
rect 65 -1764 374 -1763
rect 583 -1764 1438 -1763
rect 247 -1766 374 -1765
rect 625 -1766 1686 -1765
rect 72 -1768 248 -1767
rect 667 -1768 706 -1767
rect 709 -1768 1074 -1767
rect 72 -1770 1774 -1769
rect 688 -1772 738 -1771
rect 128 -1774 689 -1773
rect 709 -1774 867 -1773
rect 86 -1776 129 -1775
rect 86 -1778 150 -1777
rect 149 -1780 178 -1779
rect 142 -1782 178 -1781
rect 37 -1793 538 -1792
rect 541 -1793 685 -1792
rect 695 -1793 916 -1792
rect 947 -1793 1207 -1792
rect 1230 -1793 1641 -1792
rect 37 -1795 612 -1794
rect 621 -1795 1088 -1794
rect 1143 -1795 1193 -1794
rect 1395 -1795 1756 -1794
rect 30 -1797 612 -1796
rect 635 -1797 647 -1796
rect 656 -1797 892 -1796
rect 898 -1797 1214 -1796
rect 1423 -1797 1427 -1796
rect 1640 -1797 1830 -1796
rect 30 -1799 94 -1798
rect 100 -1799 118 -1798
rect 142 -1799 1053 -1798
rect 1192 -1799 1326 -1798
rect 1423 -1799 1536 -1798
rect 65 -1801 265 -1800
rect 268 -1801 647 -1800
rect 674 -1801 696 -1800
rect 716 -1801 1445 -1800
rect 68 -1803 374 -1802
rect 394 -1803 503 -1802
rect 548 -1803 1179 -1802
rect 1213 -1803 1284 -1802
rect 1325 -1803 1494 -1802
rect 72 -1805 129 -1804
rect 145 -1805 360 -1804
rect 373 -1805 710 -1804
rect 723 -1805 993 -1804
rect 1024 -1805 1690 -1804
rect 72 -1807 458 -1806
rect 499 -1807 1102 -1806
rect 1178 -1807 1228 -1806
rect 1234 -1807 1494 -1806
rect 1689 -1807 1788 -1806
rect 75 -1809 815 -1808
rect 821 -1809 836 -1808
rect 884 -1809 1669 -1808
rect 79 -1811 83 -1810
rect 89 -1811 178 -1810
rect 184 -1811 237 -1810
rect 250 -1811 458 -1810
rect 548 -1811 598 -1810
rect 674 -1811 773 -1810
rect 782 -1811 1795 -1810
rect 58 -1813 178 -1812
rect 184 -1813 318 -1812
rect 338 -1813 433 -1812
rect 576 -1813 668 -1812
rect 677 -1813 1067 -1812
rect 1101 -1813 1165 -1812
rect 1283 -1813 1333 -1812
rect 1444 -1813 1725 -1812
rect 1794 -1813 1837 -1812
rect 58 -1815 1662 -1814
rect 1668 -1815 1746 -1814
rect 79 -1817 444 -1816
rect 583 -1817 626 -1816
rect 726 -1817 1228 -1816
rect 1332 -1817 1382 -1816
rect 1661 -1817 1739 -1816
rect 1745 -1817 1816 -1816
rect 93 -1819 479 -1818
rect 534 -1819 584 -1818
rect 597 -1819 773 -1818
rect 786 -1819 1375 -1818
rect 1381 -1819 1809 -1818
rect 100 -1821 416 -1820
rect 422 -1821 671 -1820
rect 726 -1821 1028 -1820
rect 1052 -1821 1151 -1820
rect 1374 -1821 1417 -1820
rect 1577 -1821 1739 -1820
rect 110 -1823 1235 -1822
rect 1416 -1823 1585 -1822
rect 128 -1825 150 -1824
rect 159 -1825 1840 -1824
rect 149 -1827 521 -1826
rect 527 -1827 535 -1826
rect 730 -1827 759 -1826
rect 765 -1827 888 -1826
rect 891 -1827 955 -1826
rect 975 -1827 1270 -1826
rect 1293 -1827 1585 -1826
rect 170 -1829 1126 -1828
rect 1150 -1829 1165 -1828
rect 1269 -1829 1459 -1828
rect 1577 -1829 1620 -1828
rect 212 -1831 444 -1830
rect 471 -1831 626 -1830
rect 733 -1831 829 -1830
rect 831 -1831 1781 -1830
rect 114 -1833 829 -1832
rect 856 -1833 885 -1832
rect 898 -1833 920 -1832
rect 947 -1833 1385 -1832
rect 1426 -1833 1536 -1832
rect 219 -1835 325 -1834
rect 341 -1835 1095 -1834
rect 1290 -1835 1620 -1834
rect 135 -1837 325 -1836
rect 359 -1837 563 -1836
rect 758 -1837 794 -1836
rect 810 -1837 1312 -1836
rect 1458 -1837 1466 -1836
rect 135 -1839 164 -1838
rect 222 -1839 717 -1838
rect 765 -1839 1060 -1838
rect 1066 -1839 1158 -1838
rect 1311 -1839 1354 -1838
rect 1465 -1839 1473 -1838
rect 163 -1841 192 -1840
rect 222 -1841 1599 -1840
rect 191 -1843 255 -1842
rect 261 -1843 500 -1842
rect 527 -1843 1207 -1842
rect 1353 -1843 1403 -1842
rect 1430 -1843 1473 -1842
rect 1570 -1843 1599 -1842
rect 61 -1845 262 -1844
rect 268 -1845 486 -1844
rect 544 -1845 1291 -1844
rect 1297 -1845 1431 -1844
rect 1570 -1845 1823 -1844
rect 173 -1847 1403 -1846
rect 226 -1849 405 -1848
rect 415 -1849 594 -1848
rect 786 -1849 1648 -1848
rect 23 -1851 594 -1850
rect 793 -1851 843 -1850
rect 856 -1851 1098 -1850
rect 1157 -1851 1718 -1850
rect 226 -1853 633 -1852
rect 814 -1853 871 -1852
rect 901 -1853 1655 -1852
rect 233 -1855 290 -1854
rect 303 -1855 381 -1854
rect 394 -1855 790 -1854
rect 821 -1855 1137 -1854
rect 1297 -1855 1340 -1854
rect 1605 -1855 1718 -1854
rect 44 -1857 790 -1856
rect 824 -1857 1060 -1856
rect 1080 -1857 1137 -1856
rect 1605 -1857 1767 -1856
rect 44 -1859 745 -1858
rect 842 -1859 906 -1858
rect 919 -1859 969 -1858
rect 975 -1859 1018 -1858
rect 1024 -1859 1410 -1858
rect 1647 -1859 1711 -1858
rect 219 -1861 304 -1860
rect 317 -1861 507 -1860
rect 562 -1861 801 -1860
rect 870 -1861 1088 -1860
rect 1094 -1861 1627 -1860
rect 1654 -1861 1704 -1860
rect 1710 -1861 1774 -1860
rect 198 -1863 507 -1862
rect 632 -1863 640 -1862
rect 702 -1863 745 -1862
rect 800 -1863 850 -1862
rect 877 -1863 969 -1862
rect 1017 -1863 1074 -1862
rect 1080 -1863 1116 -1862
rect 1346 -1863 1767 -1862
rect 86 -1865 1074 -1864
rect 1409 -1865 1438 -1864
rect 1626 -1865 1683 -1864
rect 1703 -1865 1760 -1864
rect 86 -1867 409 -1866
rect 422 -1867 451 -1866
rect 471 -1867 986 -1866
rect 1045 -1867 1116 -1866
rect 1437 -1867 1522 -1866
rect 1591 -1867 1683 -1866
rect 156 -1869 1347 -1868
rect 1521 -1869 1543 -1868
rect 1591 -1869 1613 -1868
rect 1633 -1869 1760 -1868
rect 156 -1871 248 -1870
rect 254 -1871 720 -1870
rect 849 -1871 1305 -1870
rect 1542 -1871 1550 -1870
rect 1612 -1871 1676 -1870
rect 198 -1873 346 -1872
rect 366 -1873 836 -1872
rect 877 -1873 1011 -1872
rect 1045 -1873 1172 -1872
rect 1304 -1873 1319 -1872
rect 1549 -1873 1557 -1872
rect 1633 -1873 1697 -1872
rect 240 -1875 290 -1874
rect 296 -1875 409 -1874
rect 429 -1875 710 -1874
rect 905 -1875 1147 -1874
rect 1171 -1875 1221 -1874
rect 1318 -1875 1368 -1874
rect 1675 -1875 1732 -1874
rect 275 -1877 521 -1876
rect 618 -1877 640 -1876
rect 702 -1877 962 -1876
rect 1010 -1877 1032 -1876
rect 1360 -1877 1557 -1876
rect 1696 -1877 1753 -1876
rect 275 -1879 661 -1878
rect 688 -1879 962 -1878
rect 1360 -1879 1389 -1878
rect 1731 -1879 1802 -1878
rect 282 -1881 363 -1880
rect 366 -1881 605 -1880
rect 618 -1881 1340 -1880
rect 1367 -1881 1480 -1880
rect 282 -1883 311 -1882
rect 331 -1883 451 -1882
rect 478 -1883 493 -1882
rect 579 -1883 1389 -1882
rect 1479 -1883 1501 -1882
rect 205 -1885 311 -1884
rect 331 -1885 339 -1884
rect 345 -1885 1161 -1884
rect 1500 -1885 1508 -1884
rect 205 -1887 941 -1886
rect 954 -1887 1004 -1886
rect 1507 -1887 1515 -1886
rect 296 -1889 465 -1888
rect 485 -1889 654 -1888
rect 660 -1889 682 -1888
rect 688 -1889 979 -1888
rect 1514 -1889 1529 -1888
rect 121 -1891 654 -1890
rect 681 -1891 1039 -1890
rect 1486 -1891 1529 -1890
rect 121 -1893 738 -1892
rect 779 -1893 1221 -1892
rect 380 -1895 384 -1894
rect 401 -1895 465 -1894
rect 492 -1895 913 -1894
rect 933 -1895 1032 -1894
rect 1038 -1895 1109 -1894
rect 1129 -1895 1487 -1894
rect 401 -1897 1725 -1896
rect 436 -1899 605 -1898
rect 737 -1899 808 -1898
rect 912 -1899 1396 -1898
rect 51 -1901 808 -1900
rect 933 -1901 983 -1900
rect 1108 -1901 1277 -1900
rect 51 -1903 244 -1902
rect 436 -1903 556 -1902
rect 751 -1903 780 -1902
rect 940 -1903 997 -1902
rect 1122 -1903 1277 -1902
rect 551 -1905 1004 -1904
rect 1129 -1905 1200 -1904
rect 555 -1907 570 -1906
rect 751 -1907 927 -1906
rect 1199 -1907 1256 -1906
rect 513 -1909 570 -1908
rect 926 -1909 990 -1908
rect 1241 -1909 1256 -1908
rect 107 -1911 514 -1910
rect 1185 -1911 1242 -1910
rect 107 -1913 864 -1912
rect 1185 -1913 1249 -1912
rect 233 -1915 990 -1914
rect 1248 -1915 1263 -1914
rect 590 -1917 1263 -1916
rect 590 -1919 997 -1918
rect 863 -1921 1168 -1920
rect 23 -1932 937 -1931
rect 950 -1932 1137 -1931
rect 1157 -1932 1767 -1931
rect 30 -1934 62 -1933
rect 65 -1934 507 -1933
rect 534 -1934 608 -1933
rect 618 -1934 1291 -1933
rect 1381 -1934 1676 -1933
rect 1738 -1934 1774 -1933
rect 37 -1936 171 -1935
rect 219 -1936 395 -1935
rect 408 -1936 601 -1935
rect 656 -1936 1718 -1935
rect 37 -1938 87 -1937
rect 93 -1938 769 -1937
rect 772 -1938 934 -1937
rect 985 -1938 1361 -1937
rect 1381 -1938 1396 -1937
rect 1640 -1938 1739 -1937
rect 58 -1940 605 -1939
rect 716 -1940 804 -1939
rect 849 -1940 899 -1939
rect 912 -1940 1592 -1939
rect 1640 -1940 1655 -1939
rect 1675 -1940 1711 -1939
rect 1717 -1940 1746 -1939
rect 68 -1942 1690 -1941
rect 1710 -1942 1725 -1941
rect 79 -1944 94 -1943
rect 100 -1944 535 -1943
rect 604 -1944 682 -1943
rect 716 -1944 731 -1943
rect 754 -1944 822 -1943
rect 873 -1944 1109 -1943
rect 1122 -1944 1494 -1943
rect 1500 -1944 1690 -1943
rect 79 -1946 136 -1945
rect 138 -1946 640 -1945
rect 646 -1946 682 -1945
rect 723 -1946 934 -1945
rect 989 -1946 1368 -1945
rect 1384 -1946 1529 -1945
rect 1549 -1946 1592 -1945
rect 1654 -1946 1662 -1945
rect 1682 -1946 1746 -1945
rect 100 -1948 143 -1947
rect 149 -1948 909 -1947
rect 912 -1948 955 -1947
rect 1059 -1948 1767 -1947
rect 107 -1950 318 -1949
rect 359 -1950 871 -1949
rect 898 -1950 941 -1949
rect 947 -1950 990 -1949
rect 1080 -1950 1109 -1949
rect 1157 -1950 1172 -1949
rect 1185 -1950 1189 -1949
rect 1227 -1950 1417 -1949
rect 1423 -1950 1501 -1949
rect 1528 -1950 1763 -1949
rect 135 -1952 1221 -1951
rect 1290 -1952 1473 -1951
rect 1570 -1952 1725 -1951
rect 142 -1954 542 -1953
rect 597 -1954 955 -1953
rect 1066 -1954 1081 -1953
rect 1087 -1954 1123 -1953
rect 1160 -1954 1760 -1953
rect 149 -1956 164 -1955
rect 166 -1956 710 -1955
rect 730 -1956 1021 -1955
rect 1097 -1956 1438 -1955
rect 1661 -1956 1669 -1955
rect 1682 -1956 1753 -1955
rect 1759 -1956 1795 -1955
rect 65 -1958 164 -1957
rect 170 -1958 416 -1957
rect 432 -1958 1137 -1957
rect 1167 -1958 1648 -1957
rect 1668 -1958 1704 -1957
rect 159 -1960 353 -1959
rect 359 -1960 528 -1959
rect 639 -1960 920 -1959
rect 929 -1960 1571 -1959
rect 1696 -1960 1704 -1959
rect 72 -1962 353 -1961
rect 380 -1962 622 -1961
rect 646 -1962 661 -1961
rect 670 -1962 1697 -1961
rect 72 -1964 132 -1963
rect 219 -1964 374 -1963
rect 394 -1964 437 -1963
rect 471 -1964 542 -1963
rect 621 -1964 1536 -1963
rect 51 -1966 472 -1965
rect 492 -1966 594 -1965
rect 660 -1966 1151 -1965
rect 1171 -1966 1179 -1965
rect 1185 -1966 1242 -1965
rect 1325 -1966 1473 -1965
rect 51 -1968 346 -1967
rect 373 -1968 818 -1967
rect 821 -1968 857 -1967
rect 877 -1968 1151 -1967
rect 1178 -1968 1564 -1967
rect 117 -1970 437 -1969
rect 450 -1970 493 -1969
rect 506 -1970 570 -1969
rect 593 -1970 1396 -1969
rect 1444 -1970 1648 -1969
rect 226 -1972 311 -1971
rect 324 -1972 381 -1971
rect 401 -1972 1067 -1971
rect 1101 -1972 1417 -1971
rect 1444 -1972 1466 -1971
rect 1514 -1972 1564 -1971
rect 177 -1974 227 -1973
rect 240 -1974 339 -1973
rect 345 -1974 514 -1973
rect 555 -1974 570 -1973
rect 670 -1974 906 -1973
rect 915 -1974 1249 -1973
rect 1353 -1974 1550 -1973
rect 156 -1976 514 -1975
rect 691 -1976 1515 -1975
rect 156 -1978 727 -1977
rect 765 -1978 1494 -1977
rect 177 -1980 986 -1979
rect 1024 -1980 1354 -1979
rect 1360 -1980 1375 -1979
rect 1388 -1980 1424 -1979
rect 184 -1982 339 -1981
rect 401 -1982 685 -1981
rect 695 -1982 710 -1981
rect 765 -1982 1060 -1981
rect 1073 -1982 1102 -1981
rect 1115 -1982 1221 -1981
rect 1230 -1982 1249 -1981
rect 1367 -1982 1452 -1981
rect 184 -1984 836 -1983
rect 856 -1984 1207 -1983
rect 1213 -1984 1228 -1983
rect 1374 -1984 1480 -1983
rect 205 -1986 836 -1985
rect 905 -1986 1613 -1985
rect 205 -1988 209 -1987
rect 233 -1988 696 -1987
rect 702 -1988 871 -1987
rect 940 -1988 976 -1987
rect 1038 -1988 1074 -1987
rect 1087 -1988 1116 -1987
rect 1192 -1988 1242 -1987
rect 1388 -1988 1403 -1987
rect 1409 -1988 1466 -1987
rect 1584 -1988 1613 -1987
rect 233 -1990 598 -1989
rect 702 -1990 997 -1989
rect 1017 -1990 1039 -1989
rect 1188 -1990 1193 -1989
rect 1213 -1990 1340 -1989
rect 1402 -1990 1543 -1989
rect 240 -1992 388 -1991
rect 408 -1992 654 -1991
rect 688 -1992 997 -1991
rect 1017 -1992 1284 -1991
rect 1409 -1992 1459 -1991
rect 1542 -1992 1606 -1991
rect 247 -1994 311 -1993
rect 324 -1994 675 -1993
rect 772 -1994 843 -1993
rect 975 -1994 1004 -1993
rect 1129 -1994 1340 -1993
rect 1430 -1994 1480 -1993
rect 1598 -1994 1606 -1993
rect 107 -1996 675 -1995
rect 789 -1996 1025 -1995
rect 1052 -1996 1130 -1995
rect 1276 -1996 1284 -1995
rect 1332 -1996 1431 -1995
rect 1556 -1996 1599 -1995
rect 243 -1998 248 -1997
rect 250 -1998 1256 -1997
rect 1332 -1998 1347 -1997
rect 1556 -1998 1578 -1997
rect 254 -2000 416 -1999
rect 450 -2000 636 -1999
rect 667 -2000 1053 -1999
rect 1255 -2000 1438 -1999
rect 1577 -2000 1732 -1999
rect 254 -2002 290 -2001
rect 303 -2002 318 -2001
rect 387 -2002 549 -2001
rect 576 -2002 654 -2001
rect 667 -2002 1326 -2001
rect 1346 -2002 1508 -2001
rect 1521 -2002 1732 -2001
rect 268 -2004 619 -2003
rect 800 -2004 983 -2003
rect 1003 -2004 1011 -2003
rect 1262 -2004 1508 -2003
rect 198 -2006 269 -2005
rect 275 -2006 531 -2005
rect 548 -2006 689 -2005
rect 800 -2006 878 -2005
rect 1010 -2006 1165 -2005
rect 1311 -2006 1522 -2005
rect 110 -2008 276 -2007
rect 282 -2008 370 -2007
rect 457 -2008 577 -2007
rect 590 -2008 1585 -2007
rect 114 -2010 199 -2009
rect 229 -2010 1312 -2009
rect 114 -2012 1277 -2011
rect 282 -2014 783 -2013
rect 807 -2014 920 -2013
rect 1045 -2014 1263 -2013
rect 289 -2016 430 -2015
rect 457 -2016 626 -2015
rect 793 -2016 808 -2015
rect 810 -2016 1536 -2015
rect 303 -2018 332 -2017
rect 404 -2018 1046 -2017
rect 1164 -2018 1259 -2017
rect 331 -2020 367 -2019
rect 429 -2020 612 -2019
rect 625 -2020 864 -2019
rect 485 -2022 612 -2021
rect 814 -2022 843 -2021
rect 863 -2022 892 -2021
rect 443 -2024 486 -2023
rect 499 -2024 1207 -2023
rect 422 -2026 444 -2025
rect 478 -2026 500 -2025
rect 530 -2026 556 -2025
rect 562 -2026 794 -2025
rect 814 -2026 1487 -2025
rect 44 -2028 423 -2027
rect 562 -2028 962 -2027
rect 1125 -2028 1487 -2027
rect 44 -2030 129 -2029
rect 212 -2030 479 -2029
rect 590 -2030 759 -2029
rect 891 -2030 927 -2029
rect 961 -2030 1032 -2029
rect 128 -2032 192 -2031
rect 212 -2032 262 -2031
rect 737 -2032 927 -2031
rect 121 -2034 738 -2033
rect 758 -2034 780 -2033
rect 828 -2034 1032 -2033
rect 121 -2036 1095 -2035
rect 173 -2038 1095 -2037
rect 191 -2040 297 -2039
rect 786 -2040 829 -2039
rect 261 -2042 521 -2041
rect 751 -2042 787 -2041
rect 296 -2044 465 -2043
rect 520 -2044 664 -2043
rect 751 -2044 1459 -2043
rect 464 -2046 633 -2045
rect 86 -2048 633 -2047
rect 40 -2059 1550 -2058
rect 1626 -2059 1630 -2058
rect 1759 -2059 1767 -2058
rect 44 -2061 153 -2060
rect 163 -2061 563 -2060
rect 632 -2061 1522 -2060
rect 1626 -2061 1655 -2060
rect 1766 -2061 1774 -2060
rect 23 -2063 563 -2062
rect 663 -2063 717 -2062
rect 726 -2063 1018 -2062
rect 1090 -2063 1291 -2062
rect 1346 -2063 1522 -2062
rect 47 -2065 682 -2064
rect 688 -2065 738 -2064
rect 782 -2065 1179 -2064
rect 1206 -2065 1753 -2064
rect 68 -2067 136 -2066
rect 142 -2067 801 -2066
rect 803 -2067 1564 -2066
rect 100 -2069 780 -2068
rect 786 -2069 801 -2068
rect 873 -2069 1763 -2068
rect 100 -2071 857 -2070
rect 919 -2071 923 -2070
rect 926 -2071 1417 -2070
rect 1451 -2071 1599 -2070
rect 107 -2073 706 -2072
rect 716 -2073 745 -2072
rect 758 -2073 787 -2072
rect 856 -2073 878 -2072
rect 912 -2073 927 -2072
rect 936 -2073 1704 -2072
rect 107 -2075 370 -2074
rect 436 -2075 762 -2074
rect 779 -2075 871 -2074
rect 877 -2075 955 -2074
rect 985 -2075 1550 -2074
rect 1703 -2075 1711 -2074
rect 114 -2077 297 -2076
rect 352 -2077 437 -2076
rect 453 -2077 500 -2076
rect 506 -2077 682 -2076
rect 744 -2077 1592 -2076
rect 1696 -2077 1711 -2076
rect 54 -2079 115 -2078
rect 128 -2079 1466 -2078
rect 1570 -2079 1592 -2078
rect 1682 -2079 1697 -2078
rect 128 -2081 276 -2080
rect 289 -2081 353 -2080
rect 359 -2081 622 -2080
rect 667 -2081 808 -2080
rect 898 -2081 913 -2080
rect 919 -2081 941 -2080
rect 947 -2081 1340 -2080
rect 1395 -2081 1417 -2080
rect 1451 -2081 1557 -2080
rect 1605 -2081 1683 -2080
rect 121 -2083 668 -2082
rect 674 -2083 755 -2082
rect 758 -2083 1263 -2082
rect 1269 -2083 1466 -2082
rect 1528 -2083 1557 -2082
rect 1605 -2083 1613 -2082
rect 1629 -2083 1655 -2082
rect 121 -2085 150 -2084
rect 163 -2085 822 -2084
rect 884 -2085 948 -2084
rect 989 -2085 1021 -2084
rect 1104 -2085 1690 -2084
rect 173 -2087 1424 -2086
rect 1500 -2087 1529 -2086
rect 1535 -2087 1571 -2086
rect 1612 -2087 1634 -2086
rect 177 -2089 818 -2088
rect 821 -2089 843 -2088
rect 936 -2089 1263 -2088
rect 1311 -2089 1347 -2088
rect 1353 -2089 1396 -2088
rect 1402 -2089 1564 -2088
rect 1619 -2089 1634 -2088
rect 177 -2091 325 -2090
rect 331 -2091 507 -2090
rect 534 -2091 748 -2090
rect 989 -2091 1039 -2090
rect 1157 -2091 1179 -2090
rect 1199 -2091 1207 -2090
rect 1227 -2091 1291 -2090
rect 1325 -2091 1354 -2090
rect 1402 -2091 1445 -2090
rect 1584 -2091 1620 -2090
rect 51 -2093 535 -2092
rect 555 -2093 955 -2092
rect 1010 -2093 1039 -2092
rect 1073 -2093 1228 -2092
rect 1255 -2093 1599 -2092
rect 184 -2095 738 -2094
rect 950 -2095 1200 -2094
rect 1258 -2095 1732 -2094
rect 184 -2097 374 -2096
rect 408 -2097 843 -2096
rect 1017 -2097 1032 -2096
rect 1073 -2097 1221 -2096
rect 1339 -2097 1368 -2096
rect 1423 -2097 1648 -2096
rect 1717 -2097 1732 -2096
rect 191 -2099 636 -2098
rect 674 -2099 724 -2098
rect 817 -2099 1718 -2098
rect 142 -2101 724 -2100
rect 1031 -2101 1046 -2100
rect 1118 -2101 1326 -2100
rect 1444 -2101 1749 -2100
rect 191 -2103 262 -2102
rect 289 -2103 815 -2102
rect 1045 -2103 1053 -2102
rect 1129 -2103 1368 -2102
rect 1542 -2103 1648 -2102
rect 205 -2105 1515 -2104
rect 1584 -2105 1669 -2104
rect 96 -2107 1669 -2106
rect 205 -2109 269 -2108
rect 296 -2109 304 -2108
rect 310 -2109 332 -2108
rect 345 -2109 360 -2108
rect 366 -2109 1256 -2108
rect 1374 -2109 1515 -2108
rect 208 -2111 633 -2110
rect 691 -2111 899 -2110
rect 1052 -2111 1109 -2110
rect 1115 -2111 1130 -2110
rect 1157 -2111 1214 -2110
rect 1220 -2111 1235 -2110
rect 1332 -2111 1375 -2110
rect 1507 -2111 1543 -2110
rect 212 -2113 304 -2112
rect 310 -2113 318 -2112
rect 324 -2113 1014 -2112
rect 1101 -2113 1109 -2112
rect 1115 -2113 1501 -2112
rect 79 -2115 318 -2114
rect 338 -2115 367 -2114
rect 373 -2115 395 -2114
rect 408 -2115 549 -2114
rect 555 -2115 570 -2114
rect 576 -2115 689 -2114
rect 1171 -2115 1312 -2114
rect 1472 -2115 1508 -2114
rect 79 -2117 1746 -2116
rect 156 -2119 395 -2118
rect 422 -2119 808 -2118
rect 1192 -2119 1214 -2118
rect 1234 -2119 1249 -2118
rect 1437 -2119 1473 -2118
rect 1724 -2119 1746 -2118
rect 131 -2121 157 -2120
rect 166 -2121 577 -2120
rect 593 -2121 1333 -2120
rect 1409 -2121 1438 -2120
rect 1577 -2121 1725 -2120
rect 212 -2123 832 -2122
rect 905 -2123 1578 -2122
rect 233 -2125 528 -2124
rect 541 -2125 549 -2124
rect 569 -2125 773 -2124
rect 1192 -2125 1277 -2124
rect 1388 -2125 1410 -2124
rect 233 -2127 255 -2126
rect 338 -2127 416 -2126
rect 429 -2127 500 -2126
rect 530 -2127 542 -2126
rect 607 -2127 1536 -2126
rect 86 -2129 255 -2128
rect 345 -2129 734 -2128
rect 765 -2129 1172 -2128
rect 1276 -2129 1641 -2128
rect 37 -2131 766 -2130
rect 772 -2131 1494 -2130
rect 86 -2133 479 -2132
rect 485 -2133 598 -2132
rect 618 -2133 906 -2132
rect 1381 -2133 1389 -2132
rect 1479 -2133 1494 -2132
rect 30 -2135 619 -2134
rect 621 -2135 647 -2134
rect 660 -2135 1249 -2134
rect 1360 -2135 1382 -2134
rect 1458 -2135 1480 -2134
rect 1486 -2135 1641 -2134
rect 51 -2137 479 -2136
rect 485 -2137 731 -2136
rect 1059 -2137 1487 -2136
rect 240 -2139 276 -2138
rect 387 -2139 423 -2138
rect 429 -2139 969 -2138
rect 1059 -2139 1088 -2138
rect 1318 -2139 1361 -2138
rect 170 -2141 241 -2140
rect 247 -2141 262 -2140
rect 387 -2141 444 -2140
rect 457 -2141 885 -2140
rect 968 -2141 1004 -2140
rect 1087 -2141 1095 -2140
rect 1304 -2141 1319 -2140
rect 93 -2143 458 -2142
rect 464 -2143 591 -2142
rect 653 -2143 731 -2142
rect 814 -2143 1004 -2142
rect 1094 -2143 1144 -2142
rect 1297 -2143 1305 -2142
rect 93 -2145 997 -2144
rect 1122 -2145 1144 -2144
rect 1283 -2145 1298 -2144
rect 58 -2147 997 -2146
rect 1241 -2147 1284 -2146
rect 58 -2149 626 -2148
rect 670 -2149 1459 -2148
rect 170 -2151 1690 -2150
rect 219 -2153 444 -2152
rect 471 -2153 909 -2152
rect 1185 -2153 1242 -2152
rect 198 -2155 220 -2154
rect 226 -2155 248 -2154
rect 362 -2155 465 -2154
rect 520 -2155 647 -2154
rect 751 -2155 1123 -2154
rect 1164 -2155 1186 -2154
rect 198 -2157 1756 -2156
rect 226 -2159 1431 -2158
rect 229 -2161 472 -2160
rect 513 -2161 521 -2160
rect 583 -2161 654 -2160
rect 751 -2161 829 -2160
rect 1150 -2161 1165 -2160
rect 65 -2163 514 -2162
rect 583 -2163 696 -2162
rect 1136 -2163 1151 -2162
rect 65 -2165 1025 -2164
rect 415 -2167 979 -2166
rect 982 -2167 1137 -2166
rect 600 -2169 1431 -2168
rect 625 -2171 892 -2170
rect 961 -2171 1025 -2170
rect 695 -2173 710 -2172
rect 849 -2173 892 -2172
rect 975 -2173 983 -2172
rect 282 -2175 710 -2174
rect 849 -2175 864 -2174
rect 282 -2177 402 -2176
rect 639 -2177 864 -2176
rect 72 -2179 640 -2178
rect 702 -2179 962 -2178
rect 72 -2181 934 -2180
rect 380 -2183 402 -2182
rect 702 -2183 794 -2182
rect 933 -2183 1270 -2182
rect 380 -2185 451 -2184
rect 450 -2187 661 -2186
rect 30 -2198 451 -2197
rect 453 -2198 654 -2197
rect 688 -2198 794 -2197
rect 796 -2198 1396 -2197
rect 1640 -2198 1707 -2197
rect 1752 -2198 1767 -2197
rect 44 -2200 871 -2199
rect 873 -2200 1466 -2199
rect 1640 -2200 1697 -2199
rect 51 -2202 73 -2201
rect 89 -2202 104 -2201
rect 117 -2202 1445 -2201
rect 1465 -2202 1515 -2201
rect 1682 -2202 1714 -2201
rect 51 -2204 395 -2203
rect 408 -2204 780 -2203
rect 786 -2204 815 -2203
rect 828 -2204 1368 -2203
rect 1514 -2204 1550 -2203
rect 1682 -2204 1718 -2203
rect 58 -2206 958 -2205
rect 978 -2206 1424 -2205
rect 1549 -2206 1592 -2205
rect 1696 -2206 1739 -2205
rect 58 -2208 640 -2207
rect 691 -2208 717 -2207
rect 723 -2208 1347 -2207
rect 1423 -2208 1473 -2207
rect 1738 -2208 1760 -2207
rect 65 -2210 605 -2209
rect 607 -2210 808 -2209
rect 814 -2210 822 -2209
rect 828 -2210 843 -2209
rect 852 -2210 1032 -2209
rect 1118 -2210 1662 -2209
rect 68 -2212 563 -2211
rect 611 -2212 748 -2211
rect 758 -2212 1130 -2211
rect 1146 -2212 1732 -2211
rect 72 -2214 122 -2213
rect 131 -2214 1018 -2213
rect 1031 -2214 1102 -2213
rect 1129 -2214 1207 -2213
rect 1227 -2214 1732 -2213
rect 89 -2216 178 -2215
rect 184 -2216 605 -2215
rect 618 -2216 1368 -2215
rect 1507 -2216 1662 -2215
rect 93 -2218 885 -2217
rect 891 -2218 937 -2217
rect 999 -2218 1277 -2217
rect 1335 -2218 1655 -2217
rect 96 -2220 1123 -2219
rect 1192 -2220 1396 -2219
rect 96 -2222 185 -2221
rect 226 -2222 416 -2221
rect 450 -2222 647 -2221
rect 695 -2222 731 -2221
rect 733 -2222 1704 -2221
rect 121 -2224 234 -2223
rect 236 -2224 794 -2223
rect 807 -2224 836 -2223
rect 842 -2224 878 -2223
rect 884 -2224 1067 -2223
rect 1122 -2224 1746 -2223
rect 142 -2226 146 -2225
rect 152 -2226 1445 -2225
rect 142 -2228 626 -2227
rect 639 -2228 1039 -2227
rect 1066 -2228 1756 -2227
rect 170 -2230 318 -2229
rect 362 -2230 874 -2229
rect 877 -2230 906 -2229
rect 933 -2230 1284 -2229
rect 1346 -2230 1403 -2229
rect 170 -2232 524 -2231
rect 569 -2232 696 -2231
rect 702 -2232 1634 -2231
rect 177 -2234 206 -2233
rect 229 -2234 955 -2233
rect 999 -2234 1718 -2233
rect 205 -2236 346 -2235
rect 464 -2236 612 -2235
rect 618 -2236 675 -2235
rect 702 -2236 1214 -2235
rect 1227 -2236 1298 -2235
rect 1339 -2236 1403 -2235
rect 1626 -2236 1634 -2235
rect 100 -2238 675 -2237
rect 716 -2238 752 -2237
rect 772 -2238 1508 -2237
rect 1612 -2238 1627 -2237
rect 44 -2240 773 -2239
rect 786 -2240 801 -2239
rect 821 -2240 850 -2239
rect 891 -2240 1046 -2239
rect 1206 -2240 1319 -2239
rect 1339 -2240 1389 -2239
rect 1542 -2240 1613 -2239
rect 100 -2242 136 -2241
rect 191 -2242 346 -2241
rect 422 -2242 465 -2241
rect 471 -2242 563 -2241
rect 569 -2242 1060 -2241
rect 1213 -2242 1256 -2241
rect 1276 -2242 1487 -2241
rect 1542 -2242 1578 -2241
rect 135 -2244 1620 -2243
rect 191 -2246 241 -2245
rect 268 -2246 556 -2245
rect 586 -2246 1193 -2245
rect 1237 -2246 1676 -2245
rect 107 -2248 241 -2247
rect 271 -2248 542 -2247
rect 548 -2248 556 -2247
rect 646 -2248 661 -2247
rect 730 -2248 1473 -2247
rect 1486 -2248 1522 -2247
rect 1577 -2248 1704 -2247
rect 107 -2250 164 -2249
rect 233 -2250 262 -2249
rect 282 -2250 776 -2249
rect 800 -2250 927 -2249
rect 933 -2250 969 -2249
rect 1003 -2250 1102 -2249
rect 1255 -2250 1431 -2249
rect 1521 -2250 1725 -2249
rect 114 -2252 262 -2251
rect 282 -2252 437 -2251
rect 506 -2252 734 -2251
rect 737 -2252 780 -2251
rect 835 -2252 962 -2251
rect 1003 -2252 1151 -2251
rect 1283 -2252 1417 -2251
rect 163 -2254 633 -2253
rect 656 -2254 661 -2253
rect 747 -2254 1676 -2253
rect 215 -2256 738 -2255
rect 751 -2256 857 -2255
rect 898 -2256 962 -2255
rect 1010 -2256 1361 -2255
rect 1388 -2256 1599 -2255
rect 156 -2258 899 -2257
rect 905 -2258 920 -2257
rect 926 -2258 1025 -2257
rect 1038 -2258 1200 -2257
rect 1290 -2258 1725 -2257
rect 156 -2260 535 -2259
rect 541 -2260 983 -2259
rect 1010 -2260 1109 -2259
rect 1199 -2260 1235 -2259
rect 1290 -2260 1375 -2259
rect 1584 -2260 1599 -2259
rect 128 -2262 1585 -2261
rect 40 -2264 129 -2263
rect 289 -2264 626 -2263
rect 761 -2264 920 -2263
rect 982 -2264 1137 -2263
rect 1297 -2264 1382 -2263
rect 173 -2266 1382 -2265
rect 173 -2268 902 -2267
rect 1013 -2268 1025 -2267
rect 1045 -2268 1095 -2267
rect 1108 -2268 1669 -2267
rect 289 -2270 381 -2269
rect 436 -2270 514 -2269
rect 520 -2270 1620 -2269
rect 1668 -2270 1711 -2269
rect 114 -2272 514 -2271
rect 548 -2272 682 -2271
rect 849 -2272 1655 -2271
rect 149 -2274 521 -2273
rect 681 -2274 832 -2273
rect 1017 -2274 1053 -2273
rect 1059 -2274 1186 -2273
rect 1318 -2274 1459 -2273
rect 1591 -2274 1711 -2273
rect 149 -2276 255 -2275
rect 296 -2276 360 -2275
rect 478 -2276 633 -2275
rect 1052 -2276 1081 -2275
rect 1094 -2276 1564 -2275
rect 219 -2278 381 -2277
rect 478 -2278 598 -2277
rect 1073 -2278 1151 -2277
rect 1185 -2278 1249 -2277
rect 1332 -2278 1417 -2277
rect 1458 -2278 1480 -2277
rect 1556 -2278 1564 -2277
rect 145 -2280 220 -2279
rect 247 -2280 255 -2279
rect 296 -2280 710 -2279
rect 1073 -2280 1165 -2279
rect 1353 -2280 1431 -2279
rect 1479 -2280 1529 -2279
rect 1556 -2280 1606 -2279
rect 79 -2282 248 -2281
rect 303 -2282 395 -2281
rect 457 -2282 710 -2281
rect 968 -2282 1354 -2281
rect 1360 -2282 1410 -2281
rect 1493 -2282 1606 -2281
rect 79 -2284 199 -2283
rect 310 -2284 976 -2283
rect 1136 -2284 1263 -2283
rect 1304 -2284 1529 -2283
rect 86 -2286 458 -2285
rect 492 -2286 535 -2285
rect 723 -2286 1305 -2285
rect 1374 -2286 1452 -2285
rect 1493 -2286 1690 -2285
rect 138 -2288 304 -2287
rect 310 -2288 486 -2287
rect 499 -2288 507 -2287
rect 653 -2288 1690 -2287
rect 198 -2290 1105 -2289
rect 1157 -2290 1249 -2289
rect 1269 -2290 1452 -2289
rect 317 -2292 689 -2291
rect 744 -2292 1410 -2291
rect 324 -2294 857 -2293
rect 975 -2294 990 -2293
rect 1083 -2294 1263 -2293
rect 324 -2296 367 -2295
rect 373 -2296 486 -2295
rect 499 -2296 864 -2295
rect 989 -2296 1312 -2295
rect 275 -2298 367 -2297
rect 429 -2298 493 -2297
rect 744 -2298 948 -2297
rect 954 -2298 1312 -2297
rect 212 -2300 276 -2299
rect 331 -2300 423 -2299
rect 429 -2300 706 -2299
rect 863 -2300 1144 -2299
rect 1157 -2300 1221 -2299
rect 331 -2302 1116 -2301
rect 1164 -2302 1242 -2301
rect 338 -2304 374 -2303
rect 415 -2304 706 -2303
rect 912 -2304 1116 -2303
rect 1171 -2304 1221 -2303
rect 1241 -2304 1326 -2303
rect 338 -2306 402 -2305
rect 912 -2306 941 -2305
rect 947 -2306 1333 -2305
rect 352 -2308 402 -2307
rect 940 -2308 1088 -2307
rect 1143 -2308 1326 -2307
rect 352 -2310 577 -2309
rect 1087 -2310 1179 -2309
rect 359 -2312 388 -2311
rect 576 -2312 668 -2311
rect 996 -2312 1179 -2311
rect 387 -2314 528 -2313
rect 667 -2314 766 -2313
rect 996 -2314 1270 -2313
rect 443 -2316 766 -2315
rect 443 -2318 584 -2317
rect 471 -2320 584 -2319
rect 527 -2322 871 -2321
rect 51 -2333 181 -2332
rect 215 -2333 976 -2332
rect 982 -2333 997 -2332
rect 999 -2333 1487 -2332
rect 1514 -2333 1539 -2332
rect 1605 -2333 1707 -2332
rect 51 -2335 227 -2334
rect 443 -2335 825 -2334
rect 856 -2335 972 -2334
rect 982 -2335 1046 -2334
rect 1076 -2335 1438 -2334
rect 1493 -2335 1515 -2334
rect 1605 -2335 1676 -2334
rect 79 -2337 703 -2336
rect 733 -2337 1123 -2336
rect 1171 -2337 1452 -2336
rect 1612 -2337 1676 -2336
rect 79 -2339 94 -2338
rect 100 -2339 1126 -2338
rect 1171 -2339 1179 -2338
rect 1244 -2339 1669 -2338
rect 86 -2341 1690 -2340
rect 86 -2343 129 -2342
rect 135 -2343 381 -2342
rect 415 -2343 444 -2342
rect 450 -2343 584 -2342
rect 597 -2343 657 -2342
rect 660 -2343 678 -2342
rect 684 -2343 1585 -2342
rect 93 -2345 423 -2344
rect 464 -2345 468 -2344
rect 492 -2345 731 -2344
rect 775 -2345 1396 -2344
rect 1437 -2345 1473 -2344
rect 100 -2347 262 -2346
rect 345 -2347 451 -2346
rect 457 -2347 493 -2346
rect 502 -2347 535 -2346
rect 548 -2347 584 -2346
rect 597 -2347 643 -2346
rect 691 -2347 1564 -2346
rect 65 -2349 458 -2348
rect 464 -2349 486 -2348
rect 527 -2349 1046 -2348
rect 1080 -2349 1529 -2348
rect 1556 -2349 1564 -2348
rect 65 -2351 150 -2350
rect 163 -2351 237 -2350
rect 240 -2351 381 -2350
rect 422 -2351 731 -2350
rect 733 -2351 1473 -2350
rect 1521 -2351 1557 -2350
rect 96 -2353 1529 -2352
rect 107 -2355 535 -2354
rect 548 -2355 563 -2354
rect 569 -2355 654 -2354
rect 800 -2355 1196 -2354
rect 1304 -2355 1627 -2354
rect 107 -2357 139 -2356
rect 149 -2357 206 -2356
rect 212 -2357 416 -2356
rect 467 -2357 486 -2356
rect 530 -2357 976 -2356
rect 989 -2357 1585 -2356
rect 58 -2359 206 -2358
rect 212 -2359 1193 -2358
rect 1304 -2359 1354 -2358
rect 1384 -2359 1571 -2358
rect 114 -2361 500 -2360
rect 576 -2361 661 -2360
rect 779 -2361 801 -2360
rect 856 -2361 1634 -2360
rect 44 -2363 577 -2362
rect 618 -2363 689 -2362
rect 695 -2363 780 -2362
rect 863 -2363 1147 -2362
rect 1178 -2363 1308 -2362
rect 1314 -2363 1697 -2362
rect 114 -2365 360 -2364
rect 432 -2365 619 -2364
rect 625 -2365 1487 -2364
rect 1521 -2365 1655 -2364
rect 117 -2367 234 -2366
rect 240 -2367 388 -2366
rect 471 -2367 563 -2366
rect 590 -2367 626 -2366
rect 632 -2367 748 -2366
rect 863 -2367 1144 -2366
rect 1283 -2367 1354 -2366
rect 1388 -2367 1494 -2366
rect 1570 -2367 1599 -2366
rect 128 -2369 157 -2368
rect 163 -2369 836 -2368
rect 870 -2369 878 -2368
rect 898 -2369 1683 -2368
rect 135 -2371 605 -2370
rect 632 -2371 948 -2370
rect 954 -2371 1662 -2370
rect 142 -2373 878 -2372
rect 898 -2373 1312 -2372
rect 1332 -2373 1648 -2372
rect 142 -2375 479 -2374
rect 499 -2375 1084 -2374
rect 1097 -2375 1256 -2374
rect 1388 -2375 1410 -2374
rect 1451 -2375 1550 -2374
rect 1598 -2375 1704 -2374
rect 170 -2377 521 -2376
rect 541 -2377 748 -2376
rect 828 -2377 836 -2376
rect 873 -2377 1501 -2376
rect 170 -2379 199 -2378
rect 215 -2379 675 -2378
rect 688 -2379 724 -2378
rect 828 -2379 1067 -2378
rect 1080 -2379 1102 -2378
rect 1108 -2379 1501 -2378
rect 156 -2381 675 -2380
rect 695 -2381 710 -2380
rect 723 -2381 815 -2380
rect 919 -2381 990 -2380
rect 996 -2381 1032 -2380
rect 1066 -2381 1151 -2380
rect 1192 -2381 1284 -2380
rect 1395 -2381 1424 -2380
rect 198 -2383 297 -2382
rect 345 -2383 374 -2382
rect 387 -2383 475 -2382
rect 478 -2383 682 -2382
rect 709 -2383 717 -2382
rect 793 -2383 1102 -2382
rect 1122 -2383 1130 -2382
rect 1143 -2383 1200 -2382
rect 1255 -2383 1340 -2382
rect 1374 -2383 1424 -2382
rect 226 -2385 248 -2384
rect 254 -2385 262 -2384
rect 268 -2385 570 -2384
rect 590 -2385 612 -2384
rect 639 -2385 1620 -2384
rect 184 -2387 248 -2386
rect 254 -2387 402 -2386
rect 471 -2387 766 -2386
rect 786 -2387 794 -2386
rect 919 -2387 1214 -2386
rect 1339 -2387 1361 -2386
rect 1374 -2387 1445 -2386
rect 184 -2389 850 -2388
rect 901 -2389 1445 -2388
rect 268 -2391 430 -2390
rect 513 -2391 1151 -2390
rect 1185 -2391 1214 -2390
rect 1360 -2391 1403 -2390
rect 1409 -2391 1480 -2390
rect 282 -2393 514 -2392
rect 520 -2393 745 -2392
rect 786 -2393 822 -2392
rect 901 -2393 1431 -2392
rect 1479 -2393 1578 -2392
rect 282 -2395 290 -2394
rect 296 -2395 773 -2394
rect 814 -2395 850 -2394
rect 926 -2395 955 -2394
rect 957 -2395 1333 -2394
rect 1346 -2395 1403 -2394
rect 1430 -2395 1592 -2394
rect 173 -2397 290 -2396
rect 303 -2397 402 -2396
rect 555 -2397 612 -2396
rect 646 -2397 766 -2396
rect 772 -2397 853 -2396
rect 884 -2397 927 -2396
rect 933 -2397 948 -2396
rect 971 -2397 1459 -2396
rect 1577 -2397 1739 -2396
rect 177 -2399 304 -2398
rect 310 -2399 556 -2398
rect 604 -2399 752 -2398
rect 821 -2399 1732 -2398
rect 58 -2401 311 -2400
rect 338 -2401 374 -2400
rect 653 -2401 668 -2400
rect 716 -2401 738 -2400
rect 744 -2401 913 -2400
rect 1024 -2401 1109 -2400
rect 1115 -2401 1592 -2400
rect 177 -2403 437 -2402
rect 667 -2403 808 -2402
rect 842 -2403 885 -2402
rect 891 -2403 913 -2402
rect 1017 -2403 1025 -2402
rect 1031 -2403 1228 -2402
rect 1318 -2403 1347 -2402
rect 1458 -2403 1543 -2402
rect 191 -2405 339 -2404
rect 352 -2405 647 -2404
rect 737 -2405 811 -2404
rect 842 -2405 1004 -2404
rect 1038 -2405 1130 -2404
rect 1136 -2405 1228 -2404
rect 1535 -2405 1543 -2404
rect 191 -2407 332 -2406
rect 359 -2407 367 -2406
rect 436 -2407 507 -2406
rect 751 -2407 969 -2406
rect 1003 -2407 1291 -2406
rect 219 -2409 353 -2408
rect 506 -2409 542 -2408
rect 758 -2409 1018 -2408
rect 1038 -2409 1060 -2408
rect 1115 -2409 1158 -2408
rect 1185 -2409 1326 -2408
rect 219 -2411 318 -2410
rect 324 -2411 367 -2410
rect 758 -2411 1235 -2410
rect 1290 -2411 1382 -2410
rect 121 -2413 318 -2412
rect 324 -2413 808 -2412
rect 891 -2413 1011 -2412
rect 1059 -2413 1088 -2412
rect 1136 -2413 1718 -2412
rect 72 -2415 122 -2414
rect 331 -2415 615 -2414
rect 961 -2415 1011 -2414
rect 1073 -2415 1088 -2414
rect 1157 -2415 1165 -2414
rect 1199 -2415 1207 -2414
rect 1220 -2415 1319 -2414
rect 1325 -2415 1336 -2414
rect 1381 -2415 1417 -2414
rect 72 -2417 1095 -2416
rect 1164 -2417 1725 -2416
rect 537 -2419 1221 -2418
rect 1234 -2419 1242 -2418
rect 1276 -2419 1417 -2418
rect 933 -2421 1074 -2420
rect 1206 -2421 1298 -2420
rect 940 -2423 1095 -2422
rect 1241 -2423 1550 -2422
rect 940 -2425 1711 -2424
rect 961 -2427 1053 -2426
rect 1262 -2427 1277 -2426
rect 705 -2429 1053 -2428
rect 1262 -2429 1270 -2428
rect 408 -2431 706 -2430
rect 1269 -2431 1368 -2430
rect 275 -2433 409 -2432
rect 1367 -2433 1466 -2432
rect 275 -2435 395 -2434
rect 1465 -2435 1508 -2434
rect 394 -2437 846 -2436
rect 1507 -2437 1641 -2436
rect 44 -2448 164 -2447
rect 184 -2448 650 -2447
rect 681 -2448 745 -2447
rect 754 -2448 780 -2447
rect 786 -2448 874 -2447
rect 912 -2448 1697 -2447
rect 86 -2450 178 -2449
rect 240 -2450 860 -2449
rect 870 -2450 913 -2449
rect 957 -2450 997 -2449
rect 1062 -2450 1613 -2449
rect 1675 -2450 1732 -2449
rect 86 -2452 598 -2451
rect 611 -2452 1522 -2451
rect 1528 -2452 1679 -2451
rect 100 -2454 241 -2453
rect 257 -2454 682 -2453
rect 688 -2454 741 -2453
rect 779 -2454 801 -2453
rect 807 -2454 955 -2453
rect 971 -2454 1585 -2453
rect 1605 -2454 1725 -2453
rect 107 -2456 871 -2455
rect 891 -2456 997 -2455
rect 1076 -2456 1347 -2455
rect 1367 -2456 1522 -2455
rect 1538 -2456 1564 -2455
rect 1577 -2456 1739 -2455
rect 72 -2458 108 -2457
rect 142 -2458 167 -2457
rect 180 -2458 801 -2457
rect 821 -2458 1606 -2457
rect 142 -2460 629 -2459
rect 642 -2460 1193 -2459
rect 1227 -2460 1368 -2459
rect 1381 -2460 1480 -2459
rect 1500 -2460 1578 -2459
rect 152 -2462 1291 -2461
rect 1300 -2462 1431 -2461
rect 1458 -2462 1620 -2461
rect 282 -2464 552 -2463
rect 562 -2464 612 -2463
rect 702 -2464 829 -2463
rect 842 -2464 1074 -2463
rect 1115 -2464 1228 -2463
rect 1244 -2464 1305 -2463
rect 1311 -2464 1529 -2463
rect 1556 -2464 1711 -2463
rect 261 -2466 283 -2465
rect 296 -2466 472 -2465
rect 492 -2466 563 -2465
rect 593 -2466 1137 -2465
rect 1157 -2466 1641 -2465
rect 226 -2468 262 -2467
rect 296 -2468 353 -2467
rect 411 -2468 465 -2467
rect 502 -2468 1662 -2467
rect 93 -2470 353 -2469
rect 422 -2470 465 -2469
rect 506 -2470 689 -2469
rect 716 -2470 829 -2469
rect 845 -2470 1270 -2469
rect 1276 -2470 1347 -2469
rect 1395 -2470 1683 -2469
rect 65 -2472 94 -2471
rect 226 -2472 318 -2471
rect 324 -2472 500 -2471
rect 506 -2472 685 -2471
rect 730 -2472 1095 -2471
rect 1129 -2472 1193 -2471
rect 1199 -2472 1312 -2471
rect 1314 -2472 1487 -2471
rect 1507 -2472 1690 -2471
rect 65 -2474 80 -2473
rect 100 -2474 318 -2473
rect 324 -2474 409 -2473
rect 422 -2474 486 -2473
rect 513 -2474 542 -2473
rect 583 -2474 717 -2473
rect 751 -2474 1459 -2473
rect 1465 -2474 1585 -2473
rect 58 -2476 486 -2475
rect 513 -2476 591 -2475
rect 597 -2476 654 -2475
rect 751 -2476 1564 -2475
rect 58 -2478 633 -2477
rect 765 -2478 892 -2477
rect 919 -2478 1270 -2477
rect 1276 -2478 1452 -2477
rect 1507 -2478 1571 -2477
rect 79 -2480 346 -2479
rect 401 -2480 766 -2479
rect 793 -2480 808 -2479
rect 852 -2480 1123 -2479
rect 1129 -2480 1599 -2479
rect 121 -2482 402 -2481
rect 408 -2482 899 -2481
rect 929 -2482 1501 -2481
rect 1514 -2482 1669 -2481
rect 121 -2484 129 -2483
rect 215 -2484 1487 -2483
rect 128 -2486 150 -2485
rect 303 -2486 433 -2485
rect 436 -2486 493 -2485
rect 520 -2486 675 -2485
rect 677 -2486 1571 -2485
rect 75 -2488 437 -2487
rect 450 -2488 654 -2487
rect 674 -2488 787 -2487
rect 877 -2488 899 -2487
rect 1024 -2488 1095 -2487
rect 1167 -2488 1410 -2487
rect 1416 -2488 1515 -2487
rect 149 -2490 185 -2489
rect 303 -2490 388 -2489
rect 429 -2490 1627 -2489
rect 310 -2492 374 -2491
rect 387 -2492 458 -2491
rect 474 -2492 500 -2491
rect 520 -2492 962 -2491
rect 982 -2492 1025 -2491
rect 1031 -2492 1305 -2491
rect 1332 -2492 1410 -2491
rect 1472 -2492 1599 -2491
rect 103 -2494 374 -2493
rect 432 -2494 1718 -2493
rect 313 -2496 360 -2495
rect 443 -2496 451 -2495
rect 527 -2496 570 -2495
rect 576 -2496 1417 -2495
rect 247 -2498 360 -2497
rect 366 -2498 528 -2497
rect 541 -2498 724 -2497
rect 877 -2498 895 -2497
rect 933 -2498 962 -2497
rect 1031 -2498 1189 -2497
rect 1199 -2498 1256 -2497
rect 1290 -2498 1389 -2497
rect 1395 -2498 1550 -2497
rect 219 -2500 248 -2499
rect 275 -2500 367 -2499
rect 415 -2500 444 -2499
rect 534 -2500 724 -2499
rect 810 -2500 1389 -2499
rect 1542 -2500 1550 -2499
rect 198 -2502 220 -2501
rect 275 -2502 734 -2501
rect 884 -2502 920 -2501
rect 933 -2502 1298 -2501
rect 1325 -2502 1333 -2501
rect 1339 -2502 1655 -2501
rect 173 -2504 199 -2503
rect 331 -2504 458 -2503
rect 534 -2504 850 -2503
rect 1038 -2504 1158 -2503
rect 1178 -2504 1298 -2503
rect 1339 -2504 1581 -2503
rect 51 -2506 850 -2505
rect 1003 -2506 1039 -2505
rect 1052 -2506 1137 -2505
rect 1185 -2506 1382 -2505
rect 1444 -2506 1543 -2505
rect 51 -2508 171 -2507
rect 268 -2508 332 -2507
rect 338 -2508 342 -2507
rect 415 -2508 531 -2507
rect 548 -2508 584 -2507
rect 590 -2508 640 -2507
rect 663 -2508 1179 -2507
rect 1185 -2508 1424 -2507
rect 268 -2510 290 -2509
rect 338 -2510 381 -2509
rect 548 -2510 1116 -2509
rect 1206 -2510 1445 -2509
rect 163 -2512 1207 -2511
rect 1209 -2512 1452 -2511
rect 289 -2514 447 -2513
rect 569 -2514 605 -2513
rect 625 -2514 633 -2513
rect 695 -2514 794 -2513
rect 821 -2514 1424 -2513
rect 156 -2516 626 -2515
rect 733 -2516 1707 -2515
rect 156 -2518 748 -2517
rect 835 -2518 885 -2517
rect 926 -2518 1004 -2517
rect 1010 -2518 1053 -2517
rect 1059 -2518 1074 -2517
rect 1083 -2518 1123 -2517
rect 1213 -2518 1473 -2517
rect 341 -2520 381 -2519
rect 555 -2520 696 -2519
rect 709 -2520 836 -2519
rect 926 -2520 983 -2519
rect 1059 -2520 1151 -2519
rect 1213 -2520 1319 -2519
rect 1360 -2520 1466 -2519
rect 576 -2522 738 -2521
rect 863 -2522 1319 -2521
rect 135 -2524 738 -2523
rect 863 -2524 906 -2523
rect 975 -2524 1011 -2523
rect 1066 -2524 1431 -2523
rect 135 -2526 192 -2525
rect 394 -2526 1067 -2525
rect 1087 -2526 1151 -2525
rect 1220 -2526 1326 -2525
rect 114 -2528 192 -2527
rect 394 -2528 668 -2527
rect 705 -2528 906 -2527
rect 1087 -2528 1634 -2527
rect 114 -2530 619 -2529
rect 660 -2530 748 -2529
rect 814 -2530 976 -2529
rect 1090 -2530 1557 -2529
rect 68 -2532 619 -2531
rect 660 -2532 1375 -2531
rect 604 -2534 941 -2533
rect 1220 -2534 1592 -2533
rect 478 -2536 941 -2535
rect 1248 -2536 1648 -2535
rect 205 -2538 479 -2537
rect 667 -2538 902 -2537
rect 1143 -2538 1249 -2537
rect 1255 -2538 1354 -2537
rect 1374 -2538 1494 -2537
rect 1535 -2538 1592 -2537
rect 205 -2540 969 -2539
rect 1045 -2540 1144 -2539
rect 1234 -2540 1354 -2539
rect 1402 -2540 1494 -2539
rect 709 -2542 790 -2541
rect 814 -2542 825 -2541
rect 856 -2542 969 -2541
rect 989 -2542 1046 -2541
rect 1171 -2542 1235 -2541
rect 1262 -2542 1361 -2541
rect 1437 -2542 1536 -2541
rect 555 -2544 825 -2543
rect 856 -2544 955 -2543
rect 989 -2544 1109 -2543
rect 1164 -2544 1263 -2543
rect 1283 -2544 1403 -2543
rect 758 -2546 1284 -2545
rect 730 -2548 759 -2547
rect 1017 -2548 1109 -2547
rect 1164 -2548 1480 -2547
rect 772 -2550 1018 -2549
rect 1101 -2550 1172 -2549
rect 1195 -2550 1438 -2549
rect 646 -2552 773 -2551
rect 1080 -2552 1102 -2551
rect 345 -2554 647 -2553
rect 1080 -2554 1242 -2553
rect 72 -2565 479 -2564
rect 513 -2565 787 -2564
rect 789 -2565 1431 -2564
rect 1678 -2565 1732 -2564
rect 75 -2567 1564 -2566
rect 1703 -2567 1739 -2566
rect 79 -2569 447 -2568
rect 460 -2569 605 -2568
rect 618 -2569 1186 -2568
rect 1430 -2569 1501 -2568
rect 1563 -2569 1627 -2568
rect 1703 -2569 1718 -2568
rect 100 -2571 850 -2570
rect 873 -2571 1242 -2570
rect 1500 -2571 1585 -2570
rect 1626 -2571 1662 -2570
rect 100 -2573 136 -2572
rect 149 -2573 1067 -2572
rect 1080 -2573 1130 -2572
rect 1178 -2573 1186 -2572
rect 1374 -2573 1585 -2572
rect 128 -2575 150 -2574
rect 170 -2575 402 -2574
rect 429 -2575 857 -2574
rect 873 -2575 1263 -2574
rect 1374 -2575 1424 -2574
rect 58 -2577 430 -2576
rect 432 -2577 528 -2576
rect 548 -2577 1459 -2576
rect 58 -2579 325 -2578
rect 373 -2579 377 -2578
rect 436 -2579 549 -2578
rect 555 -2579 787 -2578
rect 800 -2579 1424 -2578
rect 1458 -2579 1690 -2578
rect 44 -2581 556 -2580
rect 576 -2581 825 -2580
rect 845 -2581 1655 -2580
rect 44 -2583 90 -2582
rect 121 -2583 171 -2582
rect 201 -2583 1417 -2582
rect 1542 -2583 1655 -2582
rect 128 -2585 395 -2584
rect 436 -2585 479 -2584
rect 506 -2585 850 -2584
rect 856 -2585 892 -2584
rect 926 -2585 1648 -2584
rect 135 -2587 664 -2586
rect 670 -2587 1683 -2586
rect 152 -2589 1690 -2588
rect 240 -2591 577 -2590
rect 593 -2591 612 -2590
rect 625 -2591 1697 -2590
rect 240 -2593 262 -2592
rect 268 -2593 528 -2592
rect 600 -2593 1144 -2592
rect 1178 -2593 1228 -2592
rect 1262 -2593 1305 -2592
rect 1395 -2593 1662 -2592
rect 1696 -2593 1725 -2592
rect 226 -2595 269 -2594
rect 303 -2595 395 -2594
rect 401 -2595 892 -2594
rect 905 -2595 927 -2594
rect 954 -2595 1452 -2594
rect 212 -2597 227 -2596
rect 233 -2597 304 -2596
rect 324 -2597 381 -2596
rect 506 -2597 591 -2596
rect 604 -2597 675 -2596
rect 730 -2597 941 -2596
rect 1034 -2597 1130 -2596
rect 1213 -2597 1305 -2596
rect 1395 -2597 1438 -2596
rect 1451 -2597 1522 -2596
rect 117 -2599 941 -2598
rect 1038 -2599 1084 -2598
rect 1087 -2599 1284 -2598
rect 1416 -2599 1494 -2598
rect 163 -2601 591 -2600
rect 611 -2601 696 -2600
rect 733 -2601 1683 -2600
rect 163 -2603 552 -2602
rect 632 -2603 647 -2602
rect 649 -2603 1354 -2602
rect 1437 -2603 1515 -2602
rect 68 -2605 1354 -2604
rect 1493 -2605 1550 -2604
rect 166 -2607 675 -2606
rect 695 -2607 839 -2606
rect 884 -2607 930 -2606
rect 1010 -2607 1039 -2606
rect 1059 -2607 1641 -2606
rect 166 -2609 1571 -2608
rect 198 -2611 234 -2610
rect 254 -2611 283 -2610
rect 296 -2611 906 -2610
rect 1003 -2611 1011 -2610
rect 1059 -2611 1102 -2610
rect 1122 -2611 1168 -2610
rect 1227 -2611 1249 -2610
rect 1276 -2611 1571 -2610
rect 65 -2613 1004 -2612
rect 1066 -2613 1340 -2612
rect 1507 -2613 1641 -2612
rect 156 -2615 297 -2614
rect 373 -2615 423 -2614
rect 520 -2615 1091 -2614
rect 1094 -2615 1242 -2614
rect 1276 -2615 1326 -2614
rect 1507 -2615 1711 -2614
rect 156 -2617 346 -2616
rect 376 -2617 423 -2616
rect 520 -2617 563 -2616
rect 632 -2617 717 -2616
rect 733 -2617 759 -2616
rect 772 -2617 955 -2616
rect 957 -2617 1249 -2616
rect 1283 -2617 1319 -2616
rect 1325 -2617 1382 -2616
rect 1514 -2617 1592 -2616
rect 212 -2619 360 -2618
rect 380 -2619 388 -2618
rect 464 -2619 759 -2618
rect 772 -2619 808 -2618
rect 821 -2619 1221 -2618
rect 1255 -2619 1382 -2618
rect 1549 -2619 1613 -2618
rect 191 -2621 360 -2620
rect 492 -2621 563 -2620
rect 639 -2621 692 -2620
rect 716 -2621 1109 -2620
rect 1122 -2621 1151 -2620
rect 1157 -2621 1221 -2620
rect 1255 -2621 1298 -2620
rect 1318 -2621 1361 -2620
rect 1612 -2621 1634 -2620
rect 184 -2623 192 -2622
rect 254 -2623 258 -2622
rect 261 -2623 276 -2622
rect 282 -2623 500 -2622
rect 646 -2623 1165 -2622
rect 1199 -2623 1340 -2622
rect 142 -2625 185 -2624
rect 275 -2625 409 -2624
rect 418 -2625 500 -2624
rect 660 -2625 815 -2624
rect 821 -2625 829 -2624
rect 884 -2625 934 -2624
rect 957 -2625 1543 -2624
rect 107 -2627 409 -2626
rect 457 -2627 493 -2626
rect 569 -2627 829 -2626
rect 894 -2627 1522 -2626
rect 107 -2629 206 -2628
rect 310 -2629 458 -2628
rect 471 -2629 570 -2628
rect 744 -2629 766 -2628
rect 779 -2629 815 -2628
rect 933 -2629 962 -2628
rect 989 -2629 1165 -2628
rect 1199 -2629 1207 -2628
rect 1269 -2629 1634 -2628
rect 72 -2631 766 -2630
rect 803 -2631 990 -2630
rect 1024 -2631 1109 -2630
rect 1150 -2631 1676 -2630
rect 142 -2633 668 -2632
rect 747 -2633 1648 -2632
rect 177 -2635 472 -2634
rect 485 -2635 640 -2634
rect 653 -2635 668 -2634
rect 751 -2635 1487 -2634
rect 1556 -2635 1676 -2634
rect 51 -2637 178 -2636
rect 205 -2637 290 -2636
rect 317 -2637 661 -2636
rect 751 -2637 1144 -2636
rect 1157 -2637 1172 -2636
rect 1206 -2637 1235 -2636
rect 1269 -2637 1312 -2636
rect 1486 -2637 1669 -2636
rect 51 -2639 542 -2638
rect 597 -2639 780 -2638
rect 807 -2639 836 -2638
rect 947 -2639 962 -2638
rect 982 -2639 1172 -2638
rect 1297 -2639 1403 -2638
rect 1556 -2639 1620 -2638
rect 121 -2641 598 -2640
rect 625 -2641 1620 -2640
rect 247 -2643 311 -2642
rect 317 -2643 451 -2642
rect 534 -2643 654 -2642
rect 702 -2643 983 -2642
rect 1017 -2643 1025 -2642
rect 1062 -2643 1592 -2642
rect 86 -2645 703 -2644
rect 737 -2645 1669 -2644
rect 86 -2647 1578 -2646
rect 289 -2649 465 -2648
rect 534 -2649 801 -2648
rect 1017 -2649 1032 -2648
rect 1094 -2649 1235 -2648
rect 1290 -2649 1403 -2648
rect 338 -2651 388 -2650
rect 411 -2651 486 -2650
rect 541 -2651 864 -2650
rect 1031 -2651 1361 -2650
rect 219 -2653 339 -2652
rect 345 -2653 710 -2652
rect 737 -2653 878 -2652
rect 1097 -2653 1473 -2652
rect 82 -2655 220 -2654
rect 450 -2655 1214 -2654
rect 1290 -2655 1333 -2654
rect 1472 -2655 1536 -2654
rect 628 -2657 948 -2656
rect 1101 -2657 1116 -2656
rect 1311 -2657 1368 -2656
rect 1535 -2657 1606 -2656
rect 443 -2659 1606 -2658
rect 331 -2661 444 -2660
rect 709 -2661 724 -2660
rect 754 -2661 1578 -2660
rect 331 -2663 353 -2662
rect 723 -2663 843 -2662
rect 863 -2663 1046 -2662
rect 1115 -2663 1137 -2662
rect 1332 -2663 1389 -2662
rect 114 -2665 353 -2664
rect 366 -2665 1046 -2664
rect 1073 -2665 1137 -2664
rect 1367 -2665 1410 -2664
rect 366 -2667 584 -2666
rect 768 -2667 1074 -2666
rect 1388 -2667 1466 -2666
rect 415 -2669 584 -2668
rect 877 -2669 913 -2668
rect 1409 -2669 1480 -2668
rect 513 -2671 843 -2670
rect 912 -2671 920 -2670
rect 1465 -2671 1529 -2670
rect 740 -2673 1480 -2672
rect 1528 -2673 1599 -2672
rect 919 -2675 969 -2674
rect 1444 -2675 1599 -2674
rect 870 -2677 1445 -2676
rect 688 -2679 871 -2678
rect 968 -2679 997 -2678
rect 618 -2681 689 -2680
rect 677 -2683 997 -2682
rect 37 -2694 570 -2693
rect 579 -2694 794 -2693
rect 803 -2694 1396 -2693
rect 51 -2696 902 -2695
rect 926 -2696 1098 -2695
rect 1395 -2696 1487 -2695
rect 51 -2698 213 -2697
rect 250 -2698 703 -2697
rect 733 -2698 1067 -2697
rect 1094 -2698 1704 -2697
rect 58 -2700 629 -2699
rect 649 -2700 850 -2699
rect 954 -2700 1242 -2699
rect 1486 -2700 1697 -2699
rect 58 -2702 241 -2701
rect 250 -2702 633 -2701
rect 660 -2702 703 -2701
rect 758 -2702 1049 -2701
rect 1066 -2702 1123 -2701
rect 1241 -2702 1291 -2701
rect 65 -2704 654 -2703
rect 660 -2704 671 -2703
rect 674 -2704 1298 -2703
rect 65 -2706 888 -2705
rect 954 -2706 1102 -2705
rect 1290 -2706 1431 -2705
rect 68 -2708 1046 -2707
rect 1094 -2708 1669 -2707
rect 72 -2710 419 -2709
rect 453 -2710 521 -2709
rect 523 -2710 1186 -2709
rect 1297 -2710 1417 -2709
rect 1430 -2710 1557 -2709
rect 82 -2712 787 -2711
rect 793 -2712 948 -2711
rect 957 -2712 1550 -2711
rect 1556 -2712 1578 -2711
rect 110 -2714 1284 -2713
rect 1416 -2714 1620 -2713
rect 114 -2716 556 -2715
rect 583 -2716 1511 -2715
rect 1549 -2716 1599 -2715
rect 114 -2718 640 -2717
rect 653 -2718 1123 -2717
rect 1283 -2718 1424 -2717
rect 117 -2720 619 -2719
rect 625 -2720 885 -2719
rect 947 -2720 1151 -2719
rect 1423 -2720 1627 -2719
rect 121 -2722 801 -2721
rect 814 -2722 846 -2721
rect 849 -2722 1004 -2721
rect 1034 -2722 1382 -2721
rect 121 -2724 248 -2723
rect 275 -2724 279 -2723
rect 289 -2724 479 -2723
rect 481 -2724 563 -2723
rect 583 -2724 983 -2723
rect 989 -2724 1655 -2723
rect 107 -2726 290 -2725
rect 331 -2726 776 -2725
rect 786 -2726 941 -2725
rect 989 -2726 1228 -2725
rect 1381 -2726 1613 -2725
rect 86 -2728 108 -2727
rect 128 -2728 755 -2727
rect 758 -2728 934 -2727
rect 940 -2728 1130 -2727
rect 1150 -2728 1277 -2727
rect 86 -2730 1676 -2729
rect 93 -2732 129 -2731
rect 142 -2732 678 -2731
rect 688 -2732 1200 -2731
rect 1227 -2732 1410 -2731
rect 72 -2734 94 -2733
rect 149 -2734 153 -2733
rect 166 -2734 332 -2733
rect 352 -2734 640 -2733
rect 667 -2734 682 -2733
rect 765 -2734 1193 -2733
rect 1199 -2734 1326 -2733
rect 89 -2736 143 -2735
rect 149 -2736 199 -2735
rect 201 -2736 731 -2735
rect 814 -2736 864 -2735
rect 873 -2736 1130 -2735
rect 1192 -2736 1340 -2735
rect 89 -2738 339 -2737
rect 373 -2738 416 -2737
rect 429 -2738 801 -2737
rect 835 -2738 899 -2737
rect 933 -2738 1074 -2737
rect 1101 -2738 1312 -2737
rect 1325 -2738 1501 -2737
rect 166 -2740 577 -2739
rect 593 -2740 1186 -2739
rect 1311 -2740 1606 -2739
rect 180 -2742 1634 -2741
rect 184 -2744 199 -2743
rect 205 -2744 339 -2743
rect 359 -2744 374 -2743
rect 401 -2744 570 -2743
rect 597 -2744 1690 -2743
rect 156 -2746 206 -2745
rect 212 -2746 227 -2745
rect 240 -2746 262 -2745
rect 268 -2746 353 -2745
rect 359 -2746 486 -2745
rect 506 -2746 633 -2745
rect 667 -2746 1018 -2745
rect 1045 -2746 1585 -2745
rect 44 -2748 227 -2747
rect 254 -2748 262 -2747
rect 268 -2748 468 -2747
rect 485 -2748 724 -2747
rect 730 -2748 857 -2747
rect 863 -2748 1189 -2747
rect 1339 -2748 1543 -2747
rect 44 -2750 101 -2749
rect 131 -2750 724 -2749
rect 835 -2750 997 -2749
rect 1003 -2750 1137 -2749
rect 1374 -2750 1543 -2749
rect 96 -2752 157 -2751
rect 184 -2752 192 -2751
rect 254 -2752 384 -2751
rect 401 -2752 437 -2751
rect 450 -2752 983 -2751
rect 1017 -2752 1172 -2751
rect 1374 -2752 1438 -2751
rect 1458 -2752 1501 -2751
rect 100 -2754 283 -2753
rect 345 -2754 997 -2753
rect 1073 -2754 1256 -2753
rect 1437 -2754 1564 -2753
rect 275 -2756 325 -2755
rect 345 -2756 493 -2755
rect 520 -2756 689 -2755
rect 716 -2756 857 -2755
rect 884 -2756 1256 -2755
rect 1458 -2756 1662 -2755
rect 233 -2758 493 -2757
rect 534 -2758 1032 -2757
rect 1136 -2758 1270 -2757
rect 177 -2760 234 -2759
rect 282 -2760 451 -2759
rect 457 -2760 1410 -2759
rect 229 -2762 458 -2761
rect 534 -2762 976 -2761
rect 1031 -2762 1088 -2761
rect 1171 -2762 1361 -2761
rect 317 -2764 325 -2763
rect 366 -2764 507 -2763
rect 541 -2764 895 -2763
rect 898 -2764 927 -2763
rect 975 -2764 1053 -2763
rect 1269 -2764 1452 -2763
rect 296 -2766 367 -2765
rect 408 -2766 1280 -2765
rect 1360 -2766 1592 -2765
rect 296 -2768 423 -2767
rect 429 -2768 612 -2767
rect 618 -2768 1109 -2767
rect 1451 -2768 1641 -2767
rect 317 -2770 444 -2769
rect 499 -2770 612 -2769
rect 625 -2770 710 -2769
rect 716 -2770 752 -2769
rect 870 -2770 1088 -2769
rect 1108 -2770 1263 -2769
rect 278 -2772 444 -2771
rect 499 -2772 745 -2771
rect 751 -2772 773 -2771
rect 870 -2772 1165 -2771
rect 1262 -2772 1473 -2771
rect 411 -2774 528 -2773
rect 541 -2774 591 -2773
rect 597 -2774 920 -2773
rect 1052 -2774 1333 -2773
rect 1472 -2774 1508 -2773
rect 415 -2776 685 -2775
rect 709 -2776 878 -2775
rect 894 -2776 1683 -2775
rect 247 -2778 878 -2777
rect 919 -2778 1214 -2777
rect 1332 -2778 1536 -2777
rect 422 -2780 804 -2779
rect 1164 -2780 1368 -2779
rect 1493 -2780 1508 -2779
rect 436 -2782 549 -2781
rect 555 -2782 808 -2781
rect 1213 -2782 1445 -2781
rect 1493 -2782 1648 -2781
rect 219 -2784 549 -2783
rect 562 -2784 780 -2783
rect 807 -2784 962 -2783
rect 1248 -2784 1445 -2783
rect 170 -2786 220 -2785
rect 527 -2786 986 -2785
rect 1206 -2786 1249 -2785
rect 1346 -2786 1536 -2785
rect 170 -2788 769 -2787
rect 842 -2788 1207 -2787
rect 1346 -2788 1515 -2787
rect 79 -2790 1515 -2789
rect 79 -2792 395 -2791
rect 590 -2792 822 -2791
rect 842 -2792 913 -2791
rect 961 -2792 1116 -2791
rect 1367 -2792 1389 -2791
rect 394 -2794 472 -2793
rect 600 -2794 738 -2793
rect 744 -2794 829 -2793
rect 912 -2794 969 -2793
rect 1115 -2794 1389 -2793
rect 135 -2796 472 -2795
rect 674 -2796 1081 -2795
rect 135 -2798 647 -2797
rect 681 -2798 1319 -2797
rect 464 -2800 738 -2799
rect 761 -2800 780 -2799
rect 821 -2800 1011 -2799
rect 1318 -2800 1480 -2799
rect 163 -2802 1480 -2801
rect 163 -2804 906 -2803
rect 999 -2804 1081 -2803
rect 310 -2806 465 -2805
rect 765 -2806 969 -2805
rect 303 -2808 311 -2807
rect 768 -2808 1025 -2807
rect 303 -2810 514 -2809
rect 772 -2810 829 -2809
rect 838 -2810 906 -2809
rect 1024 -2810 1158 -2809
rect 513 -2812 605 -2811
rect 891 -2812 1011 -2811
rect 1157 -2812 1179 -2811
rect 604 -2814 696 -2813
rect 1178 -2814 1221 -2813
rect 695 -2816 1039 -2815
rect 1220 -2816 1466 -2815
rect 1038 -2818 1060 -2817
rect 1465 -2818 1522 -2817
rect 1059 -2820 1354 -2819
rect 1304 -2822 1522 -2821
rect 1234 -2824 1305 -2823
rect 1353 -2824 1571 -2823
rect 1234 -2826 1403 -2825
rect 1402 -2828 1529 -2827
rect 1143 -2830 1529 -2829
rect 1143 -2832 1277 -2831
rect 30 -2843 458 -2842
rect 506 -2843 657 -2842
rect 765 -2843 843 -2842
rect 887 -2843 930 -2842
rect 982 -2843 1403 -2842
rect 1514 -2843 1557 -2842
rect 37 -2845 503 -2844
rect 583 -2845 654 -2844
rect 702 -2845 843 -2844
rect 898 -2845 1375 -2844
rect 1395 -2845 1403 -2844
rect 37 -2847 500 -2846
rect 569 -2847 584 -2846
rect 593 -2847 794 -2846
rect 803 -2847 962 -2846
rect 996 -2847 1193 -2846
rect 1202 -2847 1368 -2846
rect 44 -2849 118 -2848
rect 121 -2849 566 -2848
rect 607 -2849 682 -2848
rect 751 -2849 766 -2848
rect 775 -2849 1200 -2848
rect 1276 -2849 1333 -2848
rect 1367 -2849 1389 -2848
rect 51 -2851 227 -2850
rect 250 -2851 1375 -2850
rect 1388 -2851 1445 -2850
rect 51 -2853 626 -2852
rect 653 -2853 829 -2852
rect 877 -2853 1396 -2852
rect 72 -2855 1116 -2854
rect 1118 -2855 1501 -2854
rect 75 -2857 528 -2856
rect 618 -2857 885 -2856
rect 898 -2857 1508 -2856
rect 86 -2859 304 -2858
rect 345 -2859 685 -2858
rect 751 -2859 787 -2858
rect 807 -2859 916 -2858
rect 947 -2859 983 -2858
rect 996 -2859 1067 -2858
rect 1097 -2859 1438 -2858
rect 1500 -2859 1550 -2858
rect 93 -2861 108 -2860
rect 121 -2861 265 -2860
rect 268 -2861 759 -2860
rect 828 -2861 1032 -2860
rect 1038 -2861 1095 -2860
rect 1164 -2861 1186 -2860
rect 1188 -2861 1431 -2860
rect 93 -2863 605 -2862
rect 618 -2863 717 -2862
rect 779 -2863 1039 -2862
rect 1048 -2863 1137 -2862
rect 1185 -2863 1207 -2862
rect 1279 -2863 1452 -2862
rect 96 -2865 535 -2864
rect 625 -2865 689 -2864
rect 695 -2865 808 -2864
rect 856 -2865 878 -2864
rect 905 -2865 1067 -2864
rect 1192 -2865 1214 -2864
rect 1248 -2865 1452 -2864
rect 100 -2867 178 -2866
rect 226 -2867 262 -2866
rect 268 -2867 395 -2866
rect 411 -2867 1207 -2866
rect 1213 -2867 1284 -2866
rect 1318 -2867 1333 -2866
rect 1430 -2867 1459 -2866
rect 100 -2869 230 -2868
rect 275 -2869 304 -2868
rect 345 -2869 388 -2868
rect 429 -2869 570 -2868
rect 576 -2869 696 -2868
rect 709 -2869 787 -2868
rect 800 -2869 1165 -2868
rect 1283 -2869 1511 -2868
rect 107 -2871 542 -2870
rect 646 -2871 1438 -2870
rect 1458 -2871 1536 -2870
rect 128 -2873 794 -2872
rect 800 -2873 850 -2872
rect 866 -2873 885 -2872
rect 905 -2873 934 -2872
rect 940 -2873 1032 -2872
rect 1129 -2873 1249 -2872
rect 1311 -2873 1319 -2872
rect 128 -2875 241 -2874
rect 275 -2875 311 -2874
rect 359 -2875 388 -2874
rect 450 -2875 1410 -2874
rect 135 -2877 535 -2876
rect 541 -2877 640 -2876
rect 646 -2877 990 -2876
rect 1003 -2877 1137 -2876
rect 1311 -2877 1361 -2876
rect 1409 -2877 1424 -2876
rect 135 -2879 181 -2878
rect 191 -2879 311 -2878
rect 331 -2879 451 -2878
rect 457 -2879 591 -2878
rect 660 -2879 710 -2878
rect 716 -2879 769 -2878
rect 779 -2879 864 -2878
rect 912 -2879 1046 -2878
rect 1080 -2879 1130 -2878
rect 1360 -2879 1382 -2878
rect 1423 -2879 1487 -2878
rect 142 -2881 773 -2880
rect 863 -2881 1151 -2880
rect 1381 -2881 1417 -2880
rect 1486 -2881 1522 -2880
rect 142 -2883 213 -2882
rect 219 -2883 395 -2882
rect 474 -2883 1116 -2882
rect 1150 -2883 1228 -2882
rect 1416 -2883 1448 -2882
rect 72 -2885 213 -2884
rect 219 -2885 1000 -2884
rect 1003 -2885 1074 -2884
rect 1080 -2885 1242 -2884
rect 170 -2887 500 -2886
rect 523 -2887 941 -2886
rect 961 -2887 976 -2886
rect 1010 -2887 1046 -2886
rect 1122 -2887 1228 -2886
rect 1241 -2887 1263 -2886
rect 170 -2889 1200 -2888
rect 177 -2891 241 -2890
rect 282 -2891 577 -2890
rect 660 -2891 745 -2890
rect 870 -2891 1074 -2890
rect 1087 -2891 1263 -2890
rect 163 -2893 283 -2892
rect 331 -2893 367 -2892
rect 373 -2893 521 -2892
rect 527 -2893 549 -2892
rect 555 -2893 640 -2892
rect 667 -2893 850 -2892
rect 912 -2893 1494 -2892
rect 114 -2895 521 -2894
rect 548 -2895 612 -2894
rect 667 -2895 745 -2894
rect 926 -2895 990 -2894
rect 1010 -2895 1179 -2894
rect 1493 -2895 1529 -2894
rect 163 -2897 248 -2896
rect 250 -2897 871 -2896
rect 926 -2897 1305 -2896
rect 191 -2899 206 -2898
rect 359 -2899 937 -2898
rect 975 -2899 1158 -2898
rect 1178 -2899 1291 -2898
rect 1304 -2899 1354 -2898
rect 205 -2901 255 -2900
rect 366 -2901 650 -2900
rect 674 -2901 703 -2900
rect 737 -2901 857 -2900
rect 968 -2901 1354 -2900
rect 254 -2903 339 -2902
rect 380 -2903 430 -2902
rect 485 -2903 591 -2902
rect 597 -2903 675 -2902
rect 761 -2903 969 -2902
rect 1027 -2903 1480 -2902
rect 289 -2905 339 -2904
rect 380 -2905 479 -2904
rect 485 -2905 563 -2904
rect 611 -2905 815 -2904
rect 1052 -2905 1123 -2904
rect 1157 -2905 1340 -2904
rect 1479 -2905 1543 -2904
rect 44 -2907 563 -2906
rect 761 -2907 948 -2906
rect 1052 -2907 1102 -2906
rect 1255 -2907 1340 -2906
rect 65 -2909 290 -2908
rect 408 -2909 738 -2908
rect 814 -2909 836 -2908
rect 1059 -2909 1088 -2908
rect 1101 -2909 1144 -2908
rect 1255 -2909 1298 -2908
rect 65 -2911 416 -2910
rect 436 -2911 598 -2910
rect 733 -2911 1298 -2910
rect 110 -2913 836 -2912
rect 1059 -2913 1109 -2912
rect 1143 -2913 1172 -2912
rect 1290 -2913 1347 -2912
rect 401 -2915 416 -2914
rect 436 -2915 493 -2914
rect 555 -2915 920 -2914
rect 1171 -2915 1235 -2914
rect 58 -2917 402 -2916
rect 408 -2917 465 -2916
rect 478 -2917 902 -2916
rect 919 -2917 955 -2916
rect 1220 -2917 1235 -2916
rect 58 -2919 633 -2918
rect 723 -2919 1109 -2918
rect 1220 -2919 1270 -2918
rect 114 -2921 633 -2920
rect 723 -2921 731 -2920
rect 891 -2921 1347 -2920
rect 149 -2923 892 -2922
rect 954 -2923 1018 -2922
rect 1269 -2923 1326 -2922
rect 149 -2925 185 -2924
rect 317 -2925 465 -2924
rect 471 -2925 731 -2924
rect 1017 -2925 1025 -2924
rect 184 -2927 199 -2926
rect 257 -2927 318 -2926
rect 404 -2927 1326 -2926
rect 198 -2929 297 -2928
rect 422 -2929 493 -2928
rect 1024 -2929 1466 -2928
rect 79 -2931 297 -2930
rect 422 -2931 671 -2930
rect 1465 -2931 1473 -2930
rect 79 -2933 325 -2932
rect 471 -2933 507 -2932
rect 233 -2935 325 -2934
rect 233 -2937 353 -2936
rect 352 -2939 514 -2938
rect 443 -2941 514 -2940
rect 156 -2943 444 -2942
rect 30 -2954 73 -2953
rect 79 -2954 475 -2953
rect 523 -2954 633 -2953
rect 635 -2954 969 -2953
rect 982 -2954 1025 -2953
rect 1038 -2954 1042 -2953
rect 1062 -2954 1431 -2953
rect 1444 -2954 1487 -2953
rect 37 -2956 97 -2955
rect 100 -2956 703 -2955
rect 758 -2956 766 -2955
rect 828 -2956 864 -2955
rect 870 -2956 1000 -2955
rect 1020 -2956 1151 -2955
rect 1199 -2956 1277 -2955
rect 1447 -2956 1501 -2955
rect 37 -2958 122 -2957
rect 124 -2958 311 -2957
rect 366 -2958 853 -2957
rect 870 -2958 1438 -2957
rect 1472 -2958 1494 -2957
rect 44 -2960 251 -2959
rect 254 -2960 325 -2959
rect 373 -2960 451 -2959
rect 464 -2960 671 -2959
rect 684 -2960 1284 -2959
rect 44 -2962 150 -2961
rect 156 -2962 381 -2961
rect 429 -2962 479 -2961
rect 534 -2962 643 -2961
rect 646 -2962 934 -2961
rect 936 -2962 983 -2961
rect 996 -2962 1186 -2961
rect 1255 -2962 1284 -2961
rect 51 -2964 608 -2963
rect 611 -2964 731 -2963
rect 758 -2964 836 -2963
rect 877 -2964 1025 -2963
rect 1038 -2964 1123 -2963
rect 1143 -2964 1186 -2963
rect 1255 -2964 1396 -2963
rect 51 -2966 409 -2965
rect 429 -2966 797 -2965
rect 828 -2966 1375 -2965
rect 65 -2968 80 -2967
rect 93 -2968 622 -2967
rect 625 -2968 766 -2967
rect 793 -2968 878 -2967
rect 922 -2968 1053 -2967
rect 1073 -2968 1123 -2967
rect 1143 -2968 1242 -2967
rect 1276 -2968 1319 -2967
rect 1374 -2968 1459 -2967
rect 65 -2970 251 -2969
rect 254 -2970 276 -2969
rect 289 -2970 367 -2969
rect 373 -2970 598 -2969
rect 632 -2970 724 -2969
rect 933 -2970 990 -2969
rect 996 -2970 1333 -2969
rect 1458 -2970 1466 -2969
rect 100 -2972 542 -2971
rect 555 -2972 864 -2971
rect 954 -2972 969 -2971
rect 1041 -2972 1074 -2971
rect 1090 -2972 1410 -2971
rect 1465 -2972 1480 -2971
rect 114 -2974 150 -2973
rect 159 -2974 521 -2973
rect 527 -2974 542 -2973
rect 555 -2974 874 -2973
rect 954 -2974 1004 -2973
rect 1052 -2974 1130 -2973
rect 1136 -2974 1319 -2973
rect 1332 -2974 1452 -2973
rect 114 -2976 136 -2975
rect 177 -2976 290 -2975
rect 352 -2976 608 -2975
rect 646 -2976 696 -2975
rect 723 -2976 913 -2975
rect 1003 -2976 1060 -2975
rect 1129 -2976 1172 -2975
rect 121 -2978 136 -2977
rect 177 -2978 1326 -2977
rect 180 -2980 395 -2979
rect 408 -2980 465 -2979
rect 534 -2980 745 -2979
rect 912 -2980 976 -2979
rect 1080 -2980 1172 -2979
rect 198 -2982 605 -2981
rect 653 -2982 990 -2981
rect 1080 -2982 1109 -2981
rect 1136 -2982 1228 -2981
rect 201 -2984 514 -2983
rect 562 -2984 801 -2983
rect 1108 -2984 1270 -2983
rect 219 -2986 381 -2985
rect 394 -2986 867 -2985
rect 1150 -2986 1263 -2985
rect 226 -2988 325 -2987
rect 352 -2988 416 -2987
rect 422 -2988 528 -2987
rect 565 -2988 738 -2987
rect 800 -2988 815 -2987
rect 1094 -2988 1263 -2987
rect 170 -2990 227 -2989
rect 233 -2990 311 -2989
rect 355 -2990 479 -2989
rect 506 -2990 815 -2989
rect 1094 -2990 1193 -2989
rect 1213 -2990 1270 -2989
rect 128 -2992 234 -2991
rect 243 -2992 762 -2991
rect 1157 -2992 1214 -2991
rect 1227 -2992 1305 -2991
rect 58 -2994 129 -2993
rect 170 -2994 206 -2993
rect 257 -2994 423 -2993
rect 443 -2994 500 -2993
rect 506 -2994 717 -2993
rect 1031 -2994 1305 -2993
rect 58 -2996 164 -2995
rect 205 -2996 521 -2995
rect 569 -2996 689 -2995
rect 691 -2996 1088 -2995
rect 1157 -2996 1179 -2995
rect 1192 -2996 1235 -2995
rect 86 -2998 444 -2997
rect 450 -2998 549 -2997
rect 569 -2998 584 -2997
rect 590 -2998 741 -2997
rect 1031 -2998 1067 -2997
rect 1087 -2998 1326 -2997
rect 86 -3000 377 -2999
rect 401 -3000 745 -2999
rect 1066 -3000 1102 -2999
rect 1178 -3000 1382 -2999
rect 163 -3002 619 -3001
rect 639 -3002 654 -3001
rect 667 -3002 1354 -3001
rect 1381 -3002 1417 -3001
rect 261 -3004 549 -3003
rect 590 -3004 899 -3003
rect 926 -3004 1102 -3003
rect 1234 -3004 1340 -3003
rect 1416 -3004 1424 -3003
rect 142 -3006 262 -3005
rect 264 -3006 269 -3005
rect 275 -3006 458 -3005
rect 502 -3006 584 -3005
rect 597 -3006 850 -3005
rect 898 -3006 1224 -3005
rect 1311 -3006 1340 -3005
rect 107 -3008 458 -3007
rect 604 -3008 892 -3007
rect 1311 -3008 1389 -3007
rect 107 -3010 493 -3009
rect 611 -3010 927 -3009
rect 142 -3012 185 -3011
rect 264 -3012 773 -3011
rect 891 -3012 920 -3011
rect 184 -3014 192 -3013
rect 268 -3014 339 -3013
rect 359 -3014 626 -3013
rect 639 -3014 1347 -3013
rect 191 -3016 486 -3015
rect 492 -3016 661 -3015
rect 667 -3016 941 -3015
rect 1346 -3016 1403 -3015
rect 282 -3018 773 -3017
rect 940 -3018 962 -3017
rect 282 -3020 332 -3019
rect 338 -3020 346 -3019
rect 401 -3020 472 -3019
rect 485 -3020 734 -3019
rect 807 -3020 962 -3019
rect 296 -3022 360 -3021
rect 404 -3022 514 -3021
rect 576 -3022 920 -3021
rect 296 -3024 836 -3023
rect 317 -3026 577 -3025
rect 618 -3026 976 -3025
rect 303 -3028 318 -3027
rect 331 -3028 482 -3027
rect 660 -3028 710 -3027
rect 716 -3028 780 -3027
rect 303 -3030 1000 -3029
rect 345 -3032 437 -3031
rect 471 -3032 706 -3031
rect 779 -3032 787 -3031
rect 212 -3034 437 -3033
rect 674 -3034 731 -3033
rect 786 -3034 850 -3033
rect 212 -3036 241 -3035
rect 247 -3036 675 -3035
rect 681 -3036 710 -3035
rect 411 -3038 416 -3037
rect 681 -3038 885 -3037
rect 688 -3040 843 -3039
rect 856 -3040 885 -3039
rect 695 -3042 752 -3041
rect 842 -3042 948 -3041
rect 702 -3044 808 -3043
rect 856 -3044 1018 -3043
rect 705 -3046 1242 -3045
rect 751 -3048 930 -3047
rect 947 -3048 1011 -3047
rect 1017 -3048 1116 -3047
rect 1010 -3050 1046 -3049
rect 1115 -3050 1207 -3049
rect 1045 -3052 1165 -3051
rect 1206 -3052 1368 -3051
rect 1164 -3054 1221 -3053
rect 1220 -3056 1249 -3055
rect 1248 -3058 1298 -3057
rect 1290 -3060 1298 -3059
rect 1290 -3062 1361 -3061
rect 37 -3073 97 -3072
rect 100 -3073 580 -3072
rect 621 -3073 745 -3072
rect 775 -3073 1249 -3072
rect 1262 -3073 1287 -3072
rect 1293 -3073 1298 -3072
rect 1339 -3073 1354 -3072
rect 1367 -3073 1382 -3072
rect 1409 -3073 1417 -3072
rect 1451 -3073 1459 -3072
rect 44 -3075 220 -3074
rect 240 -3075 983 -3074
rect 1010 -3075 1088 -3074
rect 1090 -3075 1270 -3074
rect 1283 -3075 1347 -3074
rect 1458 -3075 1466 -3074
rect 51 -3077 216 -3076
rect 226 -3077 241 -3076
rect 243 -3077 339 -3076
rect 373 -3077 622 -3076
rect 639 -3077 808 -3076
rect 849 -3077 969 -3076
rect 982 -3077 1116 -3076
rect 1220 -3077 1291 -3076
rect 1346 -3077 1375 -3076
rect 1465 -3077 1473 -3076
rect 58 -3079 181 -3078
rect 191 -3079 251 -3078
rect 289 -3079 608 -3078
rect 653 -3079 706 -3078
rect 740 -3079 969 -3078
rect 1010 -3079 1053 -3078
rect 1059 -3079 1242 -3078
rect 1262 -3079 1333 -3078
rect 72 -3081 188 -3080
rect 191 -3081 269 -3080
rect 299 -3081 325 -3080
rect 338 -3081 465 -3080
rect 513 -3081 738 -3080
rect 744 -3081 801 -3080
rect 807 -3081 857 -3080
rect 870 -3081 948 -3080
rect 961 -3081 1137 -3080
rect 1164 -3081 1221 -3080
rect 1230 -3081 1312 -3080
rect 79 -3083 409 -3082
rect 436 -3083 1063 -3082
rect 1066 -3083 1116 -3082
rect 1136 -3083 1235 -3082
rect 79 -3085 94 -3084
rect 100 -3085 115 -3084
rect 121 -3085 738 -3084
rect 782 -3085 1039 -3084
rect 1052 -3085 1256 -3084
rect 86 -3087 356 -3086
rect 373 -3087 472 -3086
rect 478 -3087 801 -3086
rect 873 -3087 906 -3086
rect 929 -3087 1277 -3086
rect 65 -3089 87 -3088
rect 93 -3089 164 -3088
rect 177 -3089 416 -3088
rect 436 -3089 521 -3088
rect 523 -3089 878 -3088
rect 884 -3089 920 -3088
rect 933 -3089 948 -3088
rect 964 -3089 1186 -3088
rect 1276 -3089 1326 -3088
rect 114 -3091 129 -3090
rect 142 -3091 223 -3090
rect 226 -3091 636 -3090
rect 656 -3091 829 -3090
rect 884 -3091 892 -3090
rect 905 -3091 965 -3090
rect 996 -3091 1039 -3090
rect 1066 -3091 1095 -3090
rect 1101 -3091 1291 -3090
rect 121 -3093 157 -3092
rect 163 -3093 206 -3092
rect 247 -3093 363 -3092
rect 366 -3093 479 -3092
rect 520 -3093 612 -3092
rect 618 -3093 878 -3092
rect 912 -3093 934 -3092
rect 940 -3093 962 -3092
rect 975 -3093 1095 -3092
rect 1101 -3093 1200 -3092
rect 142 -3095 171 -3094
rect 177 -3095 185 -3094
rect 198 -3095 689 -3094
rect 702 -3095 1074 -3094
rect 1129 -3095 1200 -3094
rect 156 -3097 297 -3096
rect 303 -3097 514 -3096
rect 527 -3097 920 -3096
rect 940 -3097 955 -3096
rect 1073 -3097 1207 -3096
rect 128 -3099 304 -3098
rect 366 -3099 857 -3098
rect 898 -3099 955 -3098
rect 1164 -3099 1224 -3098
rect 170 -3101 276 -3100
rect 296 -3101 388 -3100
rect 394 -3101 416 -3100
rect 464 -3101 643 -3100
rect 674 -3101 871 -3100
rect 898 -3101 1032 -3100
rect 1206 -3101 1305 -3100
rect 198 -3103 283 -3102
rect 352 -3103 675 -3102
rect 684 -3103 773 -3102
rect 786 -3103 850 -3102
rect 912 -3103 1081 -3102
rect 201 -3105 325 -3104
rect 352 -3105 430 -3104
rect 471 -3105 598 -3104
rect 765 -3105 787 -3104
rect 793 -3105 1025 -3104
rect 1031 -3105 1109 -3104
rect 233 -3107 248 -3106
rect 261 -3107 395 -3106
rect 401 -3107 846 -3106
rect 1024 -3107 1123 -3106
rect 212 -3109 262 -3108
rect 268 -3109 311 -3108
rect 380 -3109 384 -3108
rect 387 -3109 682 -3108
rect 723 -3109 766 -3108
rect 796 -3109 881 -3108
rect 1080 -3109 1228 -3108
rect 222 -3111 402 -3110
rect 408 -3111 486 -3110
rect 506 -3111 598 -3110
rect 681 -3111 696 -3110
rect 723 -3111 759 -3110
rect 835 -3111 892 -3110
rect 1108 -3111 1151 -3110
rect 233 -3113 332 -3112
rect 380 -3113 605 -3112
rect 695 -3113 710 -3112
rect 758 -3113 843 -3112
rect 1122 -3113 1179 -3112
rect 275 -3115 346 -3114
rect 485 -3115 654 -3114
rect 709 -3115 731 -3114
rect 828 -3115 843 -3114
rect 1129 -3115 1228 -3114
rect 282 -3117 556 -3116
rect 576 -3117 612 -3116
rect 835 -3117 927 -3116
rect 1150 -3117 1189 -3116
rect 289 -3119 731 -3118
rect 814 -3119 927 -3118
rect 1178 -3119 1193 -3118
rect 310 -3121 458 -3120
rect 506 -3121 633 -3120
rect 814 -3121 822 -3120
rect 1192 -3121 1319 -3120
rect 317 -3123 332 -3122
rect 345 -3123 360 -3122
rect 457 -3123 773 -3122
rect 821 -3123 1046 -3122
rect 135 -3125 318 -3124
rect 527 -3125 626 -3124
rect 1045 -3125 1214 -3124
rect 205 -3127 360 -3126
rect 534 -3127 633 -3126
rect 1157 -3127 1214 -3126
rect 450 -3129 535 -3128
rect 541 -3129 556 -3128
rect 583 -3129 794 -3128
rect 1157 -3129 1242 -3128
rect 450 -3131 549 -3130
rect 604 -3131 864 -3130
rect 422 -3133 549 -3132
rect 625 -3133 717 -3132
rect 863 -3133 990 -3132
rect 422 -3135 577 -3134
rect 716 -3135 780 -3134
rect 989 -3135 1004 -3134
rect 492 -3137 1004 -3136
rect 443 -3139 493 -3138
rect 499 -3139 584 -3138
rect 779 -3139 976 -3138
rect 383 -3141 444 -3140
rect 499 -3141 570 -3140
rect 541 -3143 647 -3142
rect 562 -3145 647 -3144
rect 562 -3147 752 -3146
rect 569 -3149 661 -3148
rect 667 -3149 752 -3148
rect 135 -3151 661 -3150
rect 667 -3151 706 -3150
rect 58 -3162 199 -3161
rect 219 -3162 353 -3161
rect 373 -3162 430 -3161
rect 432 -3162 556 -3161
rect 569 -3162 580 -3161
rect 611 -3162 664 -3161
rect 667 -3162 780 -3161
rect 793 -3162 843 -3161
rect 845 -3162 1018 -3161
rect 1080 -3162 1088 -3161
rect 1094 -3162 1098 -3161
rect 1188 -3162 1263 -3161
rect 1332 -3162 1347 -3161
rect 1353 -3162 1361 -3161
rect 65 -3164 136 -3163
rect 145 -3164 188 -3163
rect 306 -3164 339 -3163
rect 352 -3164 388 -3163
rect 415 -3164 419 -3163
rect 471 -3164 636 -3163
rect 653 -3164 738 -3163
rect 751 -3164 794 -3163
rect 856 -3164 1053 -3163
rect 1080 -3164 1109 -3163
rect 1220 -3164 1242 -3163
rect 72 -3166 206 -3165
rect 296 -3166 339 -3165
rect 373 -3166 500 -3165
rect 513 -3166 612 -3165
rect 618 -3166 710 -3165
rect 716 -3166 738 -3165
rect 761 -3166 773 -3165
rect 775 -3166 836 -3165
rect 856 -3166 871 -3165
rect 877 -3166 969 -3165
rect 985 -3166 1123 -3165
rect 1227 -3166 1235 -3165
rect 1237 -3166 1277 -3165
rect 79 -3168 216 -3167
rect 250 -3168 717 -3167
rect 733 -3168 913 -3167
rect 919 -3168 1053 -3167
rect 1094 -3168 1130 -3167
rect 79 -3170 157 -3169
rect 180 -3170 668 -3169
rect 688 -3170 892 -3169
rect 912 -3170 948 -3169
rect 964 -3170 990 -3169
rect 999 -3170 1039 -3169
rect 1122 -3170 1193 -3169
rect 93 -3172 206 -3171
rect 327 -3172 363 -3171
rect 387 -3172 657 -3171
rect 660 -3172 822 -3171
rect 835 -3172 955 -3171
rect 968 -3172 1060 -3171
rect 1129 -3172 1137 -3171
rect 1192 -3172 1294 -3171
rect 93 -3174 171 -3173
rect 201 -3174 297 -3173
rect 401 -3174 472 -3173
rect 492 -3174 500 -3173
rect 534 -3174 538 -3173
rect 541 -3174 867 -3173
rect 870 -3174 899 -3173
rect 933 -3174 948 -3173
rect 989 -3174 1046 -3173
rect 100 -3176 153 -3175
rect 156 -3176 192 -3175
rect 324 -3176 402 -3175
rect 415 -3176 465 -3175
rect 534 -3176 549 -3175
rect 569 -3176 808 -3175
rect 863 -3176 920 -3175
rect 933 -3176 1032 -3175
rect 1045 -3176 1074 -3175
rect 100 -3178 265 -3177
rect 268 -3178 325 -3177
rect 422 -3178 514 -3177
rect 541 -3178 647 -3177
rect 660 -3178 1025 -3177
rect 1031 -3178 1245 -3177
rect 114 -3180 209 -3179
rect 247 -3180 269 -3179
rect 422 -3180 444 -3179
rect 464 -3180 486 -3179
rect 492 -3180 864 -3179
rect 880 -3180 899 -3179
rect 940 -3180 955 -3179
rect 1006 -3180 1067 -3179
rect 1073 -3180 1151 -3179
rect 121 -3182 199 -3181
rect 436 -3182 773 -3181
rect 779 -3182 927 -3181
rect 1010 -3182 1039 -3181
rect 1115 -3182 1151 -3181
rect 121 -3184 227 -3183
rect 282 -3184 437 -3183
rect 443 -3184 703 -3183
rect 705 -3184 1018 -3183
rect 1024 -3184 1158 -3183
rect 131 -3186 185 -3185
rect 282 -3186 346 -3185
rect 485 -3186 521 -3185
rect 548 -3186 675 -3185
rect 681 -3186 689 -3185
rect 695 -3186 710 -3185
rect 765 -3186 822 -3185
rect 884 -3186 997 -3185
rect 1115 -3186 1186 -3185
rect 135 -3188 458 -3187
rect 506 -3188 682 -3187
rect 800 -3188 892 -3187
rect 905 -3188 941 -3187
rect 1097 -3188 1137 -3187
rect 1143 -3188 1186 -3187
rect 142 -3190 192 -3189
rect 331 -3190 346 -3189
rect 359 -3190 997 -3189
rect 1143 -3190 1165 -3189
rect 86 -3192 143 -3191
rect 149 -3192 195 -3191
rect 359 -3192 395 -3191
rect 408 -3192 458 -3191
rect 506 -3192 584 -3191
rect 597 -3192 619 -3191
rect 625 -3192 696 -3191
rect 786 -3192 801 -3191
rect 807 -3192 815 -3191
rect 884 -3192 962 -3191
rect 1157 -3192 1172 -3191
rect 86 -3194 108 -3193
rect 163 -3194 332 -3193
rect 380 -3194 395 -3193
rect 478 -3194 598 -3193
rect 607 -3194 1011 -3193
rect 1164 -3194 1179 -3193
rect 107 -3196 234 -3195
rect 303 -3196 626 -3195
rect 632 -3196 1004 -3195
rect 1171 -3196 1207 -3195
rect 163 -3198 255 -3197
rect 317 -3198 409 -3197
rect 562 -3198 703 -3197
rect 730 -3198 787 -3197
rect 814 -3198 850 -3197
rect 905 -3198 1112 -3197
rect 1167 -3198 1207 -3197
rect 173 -3200 227 -3199
rect 254 -3200 262 -3199
rect 366 -3200 381 -3199
rect 527 -3200 563 -3199
rect 583 -3200 591 -3199
rect 639 -3200 752 -3199
rect 828 -3200 850 -3199
rect 926 -3200 983 -3199
rect 212 -3202 318 -3201
rect 366 -3202 605 -3201
rect 632 -3202 640 -3201
rect 646 -3202 783 -3201
rect 828 -3202 1004 -3201
rect 177 -3204 213 -3203
rect 222 -3204 234 -3203
rect 310 -3204 605 -3203
rect 730 -3204 745 -3203
rect 961 -3204 1060 -3203
rect 240 -3206 311 -3205
rect 450 -3206 528 -3205
rect 555 -3206 591 -3205
rect 744 -3206 759 -3205
rect 240 -3208 276 -3207
rect 289 -3208 451 -3207
rect 478 -3208 983 -3207
rect 247 -3210 290 -3209
rect 758 -3210 766 -3209
rect 261 -3212 276 -3211
rect 58 -3223 248 -3222
rect 338 -3223 342 -3222
rect 359 -3223 363 -3222
rect 380 -3223 398 -3222
rect 408 -3223 664 -3222
rect 702 -3223 759 -3222
rect 782 -3223 1032 -3222
rect 1038 -3223 1063 -3222
rect 1066 -3223 1081 -3222
rect 1101 -3223 1112 -3222
rect 1136 -3223 1158 -3222
rect 1206 -3223 1252 -3222
rect 1290 -3223 1326 -3222
rect 1328 -3223 1333 -3222
rect 1451 -3223 1455 -3222
rect 65 -3225 262 -3224
rect 338 -3225 346 -3224
rect 359 -3225 444 -3224
rect 464 -3225 580 -3224
rect 604 -3225 920 -3224
rect 982 -3225 1217 -3224
rect 1451 -3225 1459 -3224
rect 72 -3227 118 -3226
rect 121 -3227 325 -3226
rect 380 -3227 416 -3226
rect 429 -3227 489 -3226
rect 534 -3227 538 -3226
rect 548 -3227 727 -3226
rect 737 -3227 864 -3226
rect 866 -3227 934 -3226
rect 982 -3227 990 -3226
rect 992 -3227 1046 -3226
rect 1052 -3227 1102 -3226
rect 1125 -3227 1137 -3226
rect 1150 -3227 1189 -3226
rect 1213 -3227 1221 -3226
rect 79 -3229 174 -3228
rect 177 -3229 192 -3228
rect 201 -3229 388 -3228
rect 422 -3229 430 -3228
rect 443 -3229 458 -3228
rect 534 -3229 647 -3228
rect 730 -3229 738 -3228
rect 758 -3229 766 -3228
rect 786 -3229 1004 -3228
rect 1017 -3229 1168 -3228
rect 1185 -3229 1207 -3228
rect 86 -3231 129 -3230
rect 131 -3231 325 -3230
rect 352 -3231 416 -3230
rect 450 -3231 458 -3230
rect 541 -3231 647 -3230
rect 733 -3231 787 -3230
rect 849 -3231 986 -3230
rect 996 -3231 1109 -3230
rect 1150 -3231 1172 -3230
rect 1185 -3231 1200 -3230
rect 93 -3233 181 -3232
rect 187 -3233 367 -3232
rect 387 -3233 402 -3232
rect 450 -3233 472 -3232
rect 548 -3233 598 -3232
rect 604 -3233 633 -3232
rect 639 -3233 703 -3232
rect 765 -3233 829 -3232
rect 880 -3233 927 -3232
rect 933 -3233 969 -3232
rect 996 -3233 1165 -3232
rect 100 -3235 244 -3234
rect 247 -3235 276 -3234
rect 282 -3235 353 -3234
rect 366 -3235 405 -3234
rect 474 -3235 598 -3234
rect 611 -3235 640 -3234
rect 807 -3235 829 -3234
rect 898 -3235 927 -3234
rect 940 -3235 1004 -3234
rect 1059 -3235 1123 -3234
rect 1160 -3235 1172 -3234
rect 114 -3237 493 -3236
rect 555 -3237 892 -3236
rect 898 -3237 913 -3236
rect 919 -3237 1123 -3236
rect 1164 -3237 1193 -3236
rect 135 -3239 171 -3238
rect 191 -3239 402 -3238
rect 555 -3239 563 -3238
rect 569 -3239 577 -3238
rect 611 -3239 654 -3238
rect 800 -3239 808 -3238
rect 856 -3239 892 -3238
rect 940 -3239 955 -3238
rect 1080 -3239 1116 -3238
rect 149 -3241 465 -3240
rect 527 -3241 570 -3240
rect 618 -3241 626 -3240
rect 628 -3241 745 -3240
rect 793 -3241 801 -3240
rect 884 -3241 913 -3240
rect 947 -3241 955 -3240
rect 1087 -3241 1109 -3240
rect 152 -3243 577 -3242
rect 618 -3243 636 -3242
rect 653 -3243 689 -3242
rect 744 -3243 752 -3242
rect 793 -3243 822 -3242
rect 842 -3243 948 -3242
rect 226 -3245 230 -3244
rect 264 -3245 276 -3244
rect 296 -3245 423 -3244
rect 513 -3245 528 -3244
rect 558 -3245 675 -3244
rect 751 -3245 780 -3244
rect 821 -3245 962 -3244
rect 107 -3247 265 -3246
rect 268 -3247 283 -3246
rect 296 -3247 304 -3246
rect 394 -3247 633 -3246
rect 635 -3247 773 -3246
rect 842 -3247 871 -3246
rect 884 -3247 906 -3246
rect 961 -3247 1025 -3246
rect 156 -3249 395 -3248
rect 506 -3249 514 -3248
rect 562 -3249 584 -3248
rect 660 -3249 689 -3248
rect 772 -3249 815 -3248
rect 870 -3249 878 -3248
rect 905 -3249 976 -3248
rect 156 -3251 262 -3250
rect 268 -3251 290 -3250
rect 436 -3251 584 -3250
rect 660 -3251 696 -3250
rect 877 -3251 1011 -3250
rect 198 -3253 290 -3252
rect 373 -3253 437 -3252
rect 506 -3253 608 -3252
rect 667 -3253 815 -3252
rect 184 -3255 199 -3254
rect 219 -3255 304 -3254
rect 331 -3255 374 -3254
rect 590 -3255 696 -3254
rect 212 -3257 220 -3256
rect 226 -3257 255 -3256
rect 310 -3257 332 -3256
rect 667 -3257 717 -3256
rect 212 -3259 234 -3258
rect 310 -3259 479 -3258
rect 674 -3259 682 -3258
rect 709 -3259 717 -3258
rect 1454 -3259 1459 -3258
rect 163 -3261 234 -3260
rect 478 -3261 486 -3260
rect 681 -3261 724 -3260
rect 163 -3263 209 -3262
rect 408 -3263 486 -3262
rect 709 -3263 836 -3262
rect 208 -3265 241 -3264
rect 240 -3267 493 -3266
rect 163 -3278 230 -3277
rect 243 -3278 535 -3277
rect 593 -3278 647 -3277
rect 670 -3278 675 -3277
rect 684 -3278 703 -3277
rect 723 -3278 920 -3277
rect 936 -3278 941 -3277
rect 947 -3278 976 -3277
rect 982 -3278 990 -3277
rect 1003 -3278 1060 -3277
rect 1073 -3278 1077 -3277
rect 1108 -3278 1116 -3277
rect 1122 -3278 1130 -3277
rect 1136 -3278 1158 -3277
rect 1171 -3278 1186 -3277
rect 1206 -3278 1214 -3277
rect 1216 -3278 1221 -3277
rect 1251 -3278 1291 -3277
rect 1451 -3278 1462 -3277
rect 177 -3280 206 -3279
rect 208 -3280 241 -3279
rect 289 -3280 412 -3279
rect 415 -3280 647 -3279
rect 688 -3280 703 -3279
rect 730 -3280 752 -3279
rect 779 -3280 801 -3279
rect 807 -3280 836 -3279
rect 838 -3280 997 -3279
rect 1073 -3280 1081 -3279
rect 1097 -3280 1291 -3279
rect 1458 -3280 1466 -3279
rect 177 -3282 269 -3281
rect 282 -3282 290 -3281
rect 331 -3282 384 -3281
rect 394 -3282 619 -3281
rect 639 -3282 675 -3281
rect 681 -3282 689 -3281
rect 751 -3282 759 -3281
rect 779 -3282 787 -3281
rect 793 -3282 801 -3281
rect 814 -3282 850 -3281
rect 856 -3282 878 -3281
rect 912 -3282 920 -3281
rect 940 -3282 955 -3281
rect 1076 -3282 1081 -3281
rect 1101 -3282 1109 -3281
rect 1125 -3282 1165 -3281
rect 184 -3284 192 -3283
rect 226 -3284 248 -3283
rect 282 -3284 297 -3283
rect 324 -3284 395 -3283
rect 415 -3284 430 -3283
rect 457 -3284 591 -3283
rect 593 -3284 710 -3283
rect 712 -3284 815 -3283
rect 863 -3284 885 -3283
rect 912 -3284 934 -3283
rect 954 -3284 962 -3283
rect 1136 -3284 1151 -3283
rect 156 -3286 192 -3285
rect 226 -3286 619 -3285
rect 639 -3286 661 -3285
rect 681 -3286 808 -3285
rect 870 -3286 885 -3285
rect 926 -3286 962 -3285
rect 184 -3288 199 -3287
rect 296 -3288 573 -3287
rect 576 -3288 934 -3287
rect 187 -3290 269 -3289
rect 331 -3290 346 -3289
rect 366 -3290 591 -3289
rect 597 -3290 724 -3289
rect 744 -3290 787 -3289
rect 793 -3290 822 -3289
rect 877 -3290 899 -3289
rect 198 -3292 220 -3291
rect 338 -3292 346 -3291
rect 366 -3292 388 -3291
rect 422 -3292 458 -3291
rect 471 -3292 479 -3291
rect 488 -3292 584 -3291
rect 635 -3292 871 -3291
rect 891 -3292 927 -3291
rect 170 -3294 339 -3293
rect 373 -3294 430 -3293
rect 446 -3294 745 -3293
rect 758 -3294 766 -3293
rect 821 -3294 843 -3293
rect 898 -3294 906 -3293
rect 219 -3296 234 -3295
rect 275 -3296 388 -3295
rect 422 -3296 507 -3295
rect 534 -3296 542 -3295
rect 555 -3296 598 -3295
rect 660 -3296 717 -3295
rect 765 -3296 773 -3295
rect 842 -3296 846 -3295
rect 880 -3296 906 -3295
rect 233 -3298 409 -3297
rect 464 -3298 556 -3297
rect 576 -3298 710 -3297
rect 716 -3298 738 -3297
rect 254 -3300 276 -3299
rect 317 -3300 374 -3299
rect 464 -3300 605 -3299
rect 695 -3300 773 -3299
rect 254 -3302 353 -3301
rect 401 -3302 696 -3301
rect 737 -3302 892 -3301
rect 310 -3304 318 -3303
rect 352 -3304 486 -3303
rect 492 -3304 542 -3303
rect 583 -3304 633 -3303
rect 303 -3306 311 -3305
rect 380 -3306 486 -3305
rect 604 -3306 783 -3305
rect 303 -3308 993 -3307
rect 380 -3310 731 -3309
rect 401 -3312 451 -3311
rect 467 -3312 633 -3311
rect 436 -3314 493 -3313
rect 436 -3316 444 -3315
rect 450 -3316 626 -3315
rect 324 -3318 444 -3317
rect 474 -3318 514 -3317
rect 625 -3318 654 -3317
rect 478 -3320 500 -3319
rect 513 -3320 668 -3319
rect 499 -3322 521 -3321
rect 548 -3322 654 -3321
rect 506 -3324 668 -3323
rect 520 -3326 528 -3325
rect 548 -3326 563 -3325
rect 408 -3328 563 -3327
rect 527 -3330 570 -3329
rect 191 -3341 195 -3340
rect 261 -3341 619 -3340
rect 621 -3341 787 -3340
rect 807 -3341 867 -3340
rect 870 -3341 1098 -3340
rect 1115 -3341 1123 -3340
rect 1139 -3341 1144 -3340
rect 1353 -3341 1368 -3340
rect 191 -3343 234 -3342
rect 240 -3343 262 -3342
rect 264 -3343 276 -3342
rect 282 -3343 412 -3342
rect 471 -3343 570 -3342
rect 576 -3343 591 -3342
rect 604 -3343 619 -3342
rect 709 -3343 741 -3342
rect 821 -3343 836 -3342
rect 842 -3343 885 -3342
rect 894 -3343 927 -3342
rect 947 -3343 962 -3342
rect 975 -3343 997 -3342
rect 1059 -3343 1074 -3342
rect 1108 -3343 1116 -3342
rect 1290 -3343 1368 -3342
rect 198 -3345 241 -3344
rect 254 -3345 276 -3344
rect 282 -3345 290 -3344
rect 303 -3345 307 -3344
rect 338 -3345 465 -3344
rect 471 -3345 521 -3344
rect 541 -3345 934 -3344
rect 1062 -3345 1067 -3344
rect 1073 -3345 1081 -3344
rect 198 -3347 353 -3346
rect 355 -3347 507 -3346
rect 520 -3347 528 -3346
rect 558 -3347 570 -3346
rect 604 -3347 647 -3346
rect 660 -3347 710 -3346
rect 712 -3347 794 -3346
rect 828 -3347 832 -3346
rect 870 -3347 906 -3346
rect 926 -3347 955 -3346
rect 226 -3349 647 -3348
rect 737 -3349 801 -3348
rect 884 -3349 892 -3348
rect 905 -3349 913 -3348
rect 247 -3351 255 -3350
rect 268 -3351 444 -3350
rect 492 -3351 545 -3350
rect 555 -3351 661 -3350
rect 737 -3351 759 -3350
rect 775 -3351 822 -3350
rect 877 -3351 913 -3350
rect 212 -3353 269 -3352
rect 289 -3353 318 -3352
rect 366 -3353 381 -3352
rect 383 -3353 388 -3352
rect 394 -3353 468 -3352
rect 495 -3353 528 -3352
rect 744 -3353 829 -3352
rect 863 -3353 878 -3352
rect 177 -3355 395 -3354
rect 397 -3355 682 -3354
rect 744 -3355 773 -3354
rect 863 -3355 899 -3354
rect 177 -3357 230 -3356
rect 296 -3357 367 -3356
rect 373 -3357 388 -3356
rect 443 -3357 573 -3356
rect 576 -3357 682 -3356
rect 758 -3357 766 -3356
rect 205 -3359 213 -3358
rect 219 -3359 248 -3358
rect 296 -3359 360 -3358
rect 373 -3359 458 -3358
rect 499 -3359 594 -3358
rect 751 -3359 766 -3358
rect 205 -3361 325 -3360
rect 359 -3361 489 -3360
rect 499 -3361 563 -3360
rect 730 -3361 752 -3360
rect 219 -3363 332 -3362
rect 415 -3363 458 -3362
rect 716 -3363 731 -3362
rect 303 -3365 311 -3364
rect 317 -3365 409 -3364
rect 450 -3365 563 -3364
rect 639 -3365 717 -3364
rect 310 -3367 423 -3366
rect 450 -3367 479 -3366
rect 639 -3367 675 -3366
rect 306 -3369 423 -3368
rect 478 -3369 535 -3368
rect 667 -3369 675 -3368
rect 324 -3371 346 -3370
rect 352 -3371 416 -3370
rect 625 -3371 668 -3370
rect 331 -3373 437 -3372
rect 611 -3373 626 -3372
rect 345 -3375 538 -3374
rect 611 -3375 724 -3374
rect 401 -3377 437 -3376
rect 723 -3377 846 -3376
rect 401 -3379 535 -3378
rect 814 -3379 846 -3378
rect 408 -3381 486 -3380
rect 814 -3381 937 -3380
rect 485 -3383 654 -3382
rect 653 -3385 689 -3384
rect 583 -3387 689 -3386
rect 583 -3389 633 -3388
rect 548 -3391 633 -3390
rect 548 -3393 598 -3392
rect 446 -3395 598 -3394
rect 177 -3406 227 -3405
rect 247 -3406 356 -3405
rect 366 -3406 384 -3405
rect 457 -3406 496 -3405
rect 499 -3406 507 -3405
rect 513 -3406 577 -3405
rect 632 -3406 636 -3405
rect 695 -3406 703 -3405
rect 719 -3406 738 -3405
rect 765 -3406 773 -3405
rect 782 -3406 983 -3405
rect 1367 -3406 1396 -3405
rect 184 -3408 230 -3407
rect 264 -3408 269 -3407
rect 275 -3408 395 -3407
rect 467 -3408 605 -3407
rect 632 -3408 654 -3407
rect 681 -3408 766 -3407
rect 772 -3408 780 -3407
rect 831 -3408 857 -3407
rect 891 -3408 927 -3407
rect 947 -3408 965 -3407
rect 968 -3408 976 -3407
rect 212 -3410 223 -3409
rect 233 -3410 276 -3409
rect 310 -3410 395 -3409
rect 471 -3410 486 -3409
rect 499 -3410 556 -3409
rect 558 -3410 626 -3409
rect 653 -3410 668 -3409
rect 688 -3410 780 -3409
rect 842 -3410 871 -3409
rect 912 -3410 927 -3409
rect 954 -3410 1011 -3409
rect 254 -3412 311 -3411
rect 317 -3412 339 -3411
rect 341 -3412 388 -3411
rect 408 -3412 472 -3411
rect 478 -3412 493 -3411
rect 520 -3412 542 -3411
rect 569 -3412 577 -3411
rect 625 -3412 640 -3411
rect 660 -3412 682 -3411
rect 688 -3412 724 -3411
rect 730 -3412 734 -3411
rect 842 -3412 846 -3411
rect 856 -3412 885 -3411
rect 905 -3412 913 -3411
rect 961 -3412 1095 -3411
rect 191 -3414 342 -3413
rect 352 -3414 402 -3413
rect 534 -3414 549 -3413
rect 569 -3414 591 -3413
rect 597 -3414 661 -3413
rect 695 -3414 717 -3413
rect 723 -3414 815 -3413
rect 863 -3414 871 -3413
rect 877 -3414 885 -3413
rect 240 -3416 255 -3415
rect 261 -3416 269 -3415
rect 289 -3416 318 -3415
rect 327 -3416 416 -3415
rect 488 -3416 535 -3415
rect 541 -3416 643 -3415
rect 730 -3416 759 -3415
rect 821 -3416 864 -3415
rect 198 -3418 241 -3417
rect 331 -3418 402 -3417
rect 527 -3418 549 -3417
rect 562 -3418 598 -3417
rect 639 -3418 776 -3417
rect 821 -3418 836 -3417
rect 359 -3420 388 -3419
rect 562 -3420 584 -3419
rect 646 -3420 836 -3419
rect 296 -3422 360 -3421
rect 373 -3422 409 -3421
rect 583 -3422 612 -3421
rect 618 -3422 647 -3421
rect 733 -3422 759 -3421
rect 219 -3424 297 -3423
rect 303 -3424 374 -3423
rect 303 -3426 430 -3425
rect 429 -3428 437 -3427
rect 436 -3430 451 -3429
rect 422 -3432 451 -3431
rect 345 -3434 423 -3433
rect 324 -3436 346 -3435
rect 205 -3438 325 -3437
rect 222 -3449 328 -3448
rect 338 -3449 353 -3448
rect 359 -3449 381 -3448
rect 401 -3449 465 -3448
rect 478 -3449 486 -3448
rect 506 -3449 542 -3448
rect 597 -3449 605 -3448
rect 614 -3449 626 -3448
rect 642 -3449 689 -3448
rect 698 -3449 703 -3448
rect 709 -3449 738 -3448
rect 740 -3449 759 -3448
rect 765 -3449 780 -3448
rect 782 -3449 965 -3448
rect 982 -3449 1067 -3448
rect 1073 -3449 1077 -3448
rect 1094 -3449 1221 -3448
rect 1223 -3449 1228 -3448
rect 1409 -3449 1417 -3448
rect 254 -3451 262 -3450
rect 264 -3451 461 -3450
rect 471 -3451 486 -3450
rect 520 -3451 573 -3450
rect 621 -3451 724 -3450
rect 737 -3451 752 -3450
rect 821 -3451 829 -3450
rect 831 -3451 850 -3450
rect 933 -3451 955 -3450
rect 957 -3451 969 -3450
rect 1010 -3451 1074 -3450
rect 1395 -3451 1410 -3450
rect 240 -3453 255 -3452
rect 268 -3453 290 -3452
rect 292 -3453 360 -3452
rect 373 -3453 402 -3452
rect 408 -3453 416 -3452
rect 422 -3453 503 -3452
rect 541 -3453 570 -3452
rect 625 -3453 633 -3452
rect 674 -3453 692 -3452
rect 695 -3453 710 -3452
rect 719 -3453 731 -3452
rect 824 -3453 962 -3452
rect 275 -3455 307 -3454
rect 317 -3455 328 -3454
rect 345 -3455 353 -3454
rect 394 -3455 472 -3454
rect 569 -3455 584 -3454
rect 667 -3455 675 -3454
rect 681 -3455 717 -3454
rect 835 -3455 892 -3454
rect 947 -3455 976 -3454
rect 282 -3457 304 -3456
rect 310 -3457 318 -3456
rect 387 -3457 395 -3456
rect 422 -3457 430 -3456
rect 450 -3457 458 -3456
rect 576 -3457 584 -3456
rect 660 -3457 682 -3456
rect 688 -3457 745 -3456
rect 821 -3457 836 -3456
rect 849 -3457 871 -3456
rect 296 -3459 332 -3458
rect 425 -3459 640 -3458
rect 660 -3459 727 -3458
rect 863 -3459 871 -3458
rect 429 -3461 437 -3460
rect 555 -3461 577 -3460
rect 695 -3461 759 -3460
rect 555 -3463 563 -3462
rect 534 -3465 563 -3464
rect 261 -3476 269 -3475
rect 303 -3476 311 -3475
rect 317 -3476 328 -3475
rect 380 -3476 412 -3475
rect 415 -3476 437 -3475
rect 467 -3476 521 -3475
rect 548 -3476 552 -3475
rect 583 -3476 591 -3475
rect 597 -3476 661 -3475
rect 681 -3476 689 -3475
rect 695 -3476 829 -3475
rect 842 -3476 850 -3475
rect 852 -3476 857 -3475
rect 870 -3476 888 -3475
rect 891 -3476 951 -3475
rect 989 -3476 993 -3475
rect 1066 -3476 1095 -3475
rect 1115 -3476 1119 -3475
rect 1213 -3476 1221 -3475
rect 1409 -3476 1413 -3475
rect 254 -3478 262 -3477
rect 394 -3478 409 -3477
rect 418 -3478 699 -3477
rect 709 -3478 717 -3477
rect 726 -3478 738 -3477
rect 758 -3478 822 -3477
rect 877 -3478 899 -3477
rect 905 -3478 934 -3477
rect 1115 -3478 1123 -3477
rect 1220 -3478 1228 -3477
rect 1409 -3478 1417 -3477
rect 401 -3480 409 -3479
rect 429 -3480 440 -3479
rect 471 -3480 507 -3479
rect 548 -3480 556 -3479
rect 576 -3480 584 -3479
rect 604 -3480 622 -3479
rect 646 -3480 661 -3479
rect 674 -3480 682 -3479
rect 359 -3482 430 -3481
rect 436 -3482 444 -3481
rect 478 -3482 503 -3481
rect 513 -3482 647 -3481
rect 1412 -3482 1417 -3481
rect 478 -3484 615 -3483
rect 485 -3486 517 -3485
rect 562 -3486 577 -3485
rect 611 -3486 626 -3485
rect 492 -3488 500 -3487
rect 261 -3499 272 -3498
rect 310 -3499 325 -3498
rect 331 -3499 346 -3498
rect 352 -3499 360 -3498
rect 408 -3499 419 -3498
rect 429 -3499 437 -3498
rect 541 -3499 552 -3498
rect 555 -3499 566 -3498
rect 583 -3499 598 -3498
rect 646 -3499 654 -3498
rect 660 -3499 668 -3498
rect 681 -3499 692 -3498
rect 716 -3499 724 -3498
rect 828 -3499 871 -3498
rect 898 -3499 906 -3498
rect 922 -3499 927 -3498
rect 940 -3499 951 -3498
rect 989 -3499 997 -3498
rect 1094 -3499 1116 -3498
rect 1118 -3499 1123 -3498
rect 1360 -3499 1368 -3498
rect 1412 -3499 1417 -3498
rect 268 -3501 276 -3500
rect 331 -3501 339 -3500
rect 355 -3501 479 -3500
rect 541 -3501 549 -3500
rect 576 -3501 584 -3500
rect 835 -3501 860 -3500
rect 576 -3503 591 -3502
rect 842 -3503 850 -3502
rect 271 -3514 276 -3513
rect 327 -3514 332 -3513
rect 355 -3514 360 -3513
rect 541 -3514 556 -3513
rect 565 -3514 570 -3513
rect 579 -3514 584 -3513
rect 660 -3514 668 -3513
rect 856 -3514 878 -3513
rect 1353 -3514 1361 -3513
rect 1363 -3514 1368 -3513
rect 870 -3516 916 -3515
<< m2contact >>
rect 282 0 283 1
rect 345 0 346 1
rect 425 0 426 1
rect 450 0 451 1
rect 464 0 465 1
rect 478 0 479 1
rect 905 0 906 1
rect 950 0 951 1
rect 317 -2 318 -1
rect 352 -2 353 -1
rect 436 -2 437 -1
rect 513 -2 514 -1
rect 947 -2 948 -1
rect 989 -2 990 -1
rect 443 -4 444 -3
rect 457 -4 458 -3
rect 226 -15 227 -14
rect 285 -15 286 -14
rect 303 -15 304 -14
rect 317 -15 318 -14
rect 338 -15 339 -14
rect 359 -15 360 -14
rect 366 -15 367 -14
rect 436 -15 437 -14
rect 450 -15 451 -14
rect 457 -15 458 -14
rect 478 -15 479 -14
rect 499 -15 500 -14
rect 506 -15 507 -14
rect 611 -15 612 -14
rect 618 -15 619 -14
rect 625 -15 626 -14
rect 891 -15 892 -14
rect 905 -15 906 -14
rect 989 -15 990 -14
rect 1003 -15 1004 -14
rect 345 -17 346 -16
rect 373 -17 374 -16
rect 380 -17 381 -16
rect 425 -17 426 -16
rect 436 -17 437 -16
rect 443 -17 444 -16
rect 450 -17 451 -16
rect 464 -17 465 -16
rect 513 -17 514 -16
rect 548 -17 549 -16
rect 579 -17 580 -16
rect 590 -17 591 -16
rect 597 -17 598 -16
rect 639 -17 640 -16
rect 289 -19 290 -18
rect 345 -19 346 -18
rect 348 -19 349 -18
rect 408 -19 409 -18
rect 422 -19 423 -18
rect 509 -19 510 -18
rect 527 -19 528 -18
rect 541 -19 542 -18
rect 583 -19 584 -18
rect 604 -19 605 -18
rect 352 -21 353 -20
rect 387 -21 388 -20
rect 394 -21 395 -20
rect 418 -21 419 -20
rect 460 -21 461 -20
rect 464 -21 465 -20
rect 509 -21 510 -20
rect 513 -21 514 -20
rect 537 -21 538 -20
rect 674 -21 675 -20
rect 352 -23 353 -22
rect 362 -23 363 -22
rect 219 -34 220 -33
rect 226 -34 227 -33
rect 275 -34 276 -33
rect 289 -34 290 -33
rect 324 -34 325 -33
rect 366 -34 367 -33
rect 387 -34 388 -33
rect 401 -34 402 -33
rect 415 -34 416 -33
rect 436 -34 437 -33
rect 443 -34 444 -33
rect 457 -34 458 -33
rect 464 -34 465 -33
rect 471 -34 472 -33
rect 492 -34 493 -33
rect 565 -34 566 -33
rect 576 -34 577 -33
rect 597 -34 598 -33
rect 611 -34 612 -33
rect 653 -34 654 -33
rect 674 -34 675 -33
rect 723 -34 724 -33
rect 758 -34 759 -33
rect 828 -34 829 -33
rect 884 -34 885 -33
rect 891 -34 892 -33
rect 1003 -34 1004 -33
rect 1010 -34 1011 -33
rect 282 -36 283 -35
rect 296 -36 297 -35
rect 331 -36 332 -35
rect 341 -36 342 -35
rect 359 -36 360 -35
rect 432 -36 433 -35
rect 436 -36 437 -35
rect 457 -36 458 -35
rect 499 -36 500 -35
rect 502 -36 503 -35
rect 513 -36 514 -35
rect 520 -36 521 -35
rect 541 -36 542 -35
rect 555 -36 556 -35
rect 583 -36 584 -35
rect 621 -36 622 -35
rect 625 -36 626 -35
rect 632 -36 633 -35
rect 639 -36 640 -35
rect 674 -36 675 -35
rect 338 -38 339 -37
rect 345 -38 346 -37
rect 366 -38 367 -37
rect 380 -38 381 -37
rect 387 -38 388 -37
rect 485 -38 486 -37
rect 499 -38 500 -37
rect 506 -38 507 -37
rect 520 -38 521 -37
rect 527 -38 528 -37
rect 551 -38 552 -37
rect 730 -38 731 -37
rect 338 -40 339 -39
rect 422 -40 423 -39
rect 450 -40 451 -39
rect 464 -40 465 -39
rect 502 -40 503 -39
rect 506 -40 507 -39
rect 523 -40 524 -39
rect 541 -40 542 -39
rect 590 -40 591 -39
rect 597 -40 598 -39
rect 625 -40 626 -39
rect 681 -40 682 -39
rect 380 -42 381 -41
rect 394 -42 395 -41
rect 408 -42 409 -41
rect 450 -42 451 -41
rect 548 -42 549 -41
rect 590 -42 591 -41
rect 635 -42 636 -41
rect 639 -42 640 -41
rect 394 -44 395 -43
rect 537 -44 538 -43
rect 408 -46 409 -45
rect 418 -46 419 -45
rect 422 -46 423 -45
rect 429 -46 430 -45
rect 191 -57 192 -56
rect 254 -57 255 -56
rect 278 -57 279 -56
rect 282 -57 283 -56
rect 289 -57 290 -56
rect 464 -57 465 -56
rect 506 -57 507 -56
rect 516 -57 517 -56
rect 523 -57 524 -56
rect 737 -57 738 -56
rect 789 -57 790 -56
rect 863 -57 864 -56
rect 884 -57 885 -56
rect 891 -57 892 -56
rect 1010 -57 1011 -56
rect 1017 -57 1018 -56
rect 205 -59 206 -58
rect 240 -59 241 -58
rect 243 -59 244 -58
rect 261 -59 262 -58
rect 275 -59 276 -58
rect 282 -59 283 -58
rect 296 -59 297 -58
rect 303 -59 304 -58
rect 317 -59 318 -58
rect 390 -59 391 -58
rect 464 -59 465 -58
rect 499 -59 500 -58
rect 513 -59 514 -58
rect 520 -59 521 -58
rect 527 -59 528 -58
rect 586 -59 587 -58
rect 597 -59 598 -58
rect 660 -59 661 -58
rect 709 -59 710 -58
rect 758 -59 759 -58
rect 793 -59 794 -58
rect 800 -59 801 -58
rect 828 -59 829 -58
rect 898 -59 899 -58
rect 219 -61 220 -60
rect 247 -61 248 -60
rect 275 -61 276 -60
rect 310 -61 311 -60
rect 341 -61 342 -60
rect 345 -61 346 -60
rect 390 -61 391 -60
rect 478 -61 479 -60
rect 562 -61 563 -60
rect 779 -61 780 -60
rect 233 -63 234 -62
rect 320 -63 321 -62
rect 345 -63 346 -62
rect 380 -63 381 -62
rect 471 -63 472 -62
rect 499 -63 500 -62
rect 569 -63 570 -62
rect 625 -63 626 -62
rect 632 -63 633 -62
rect 646 -63 647 -62
rect 653 -63 654 -62
rect 702 -63 703 -62
rect 730 -63 731 -62
rect 807 -63 808 -62
rect 299 -65 300 -64
rect 338 -65 339 -64
rect 373 -65 374 -64
rect 380 -65 381 -64
rect 471 -65 472 -64
rect 509 -65 510 -64
rect 569 -65 570 -64
rect 583 -65 584 -64
rect 590 -65 591 -64
rect 597 -65 598 -64
rect 604 -65 605 -64
rect 632 -65 633 -64
rect 639 -65 640 -64
rect 653 -65 654 -64
rect 723 -65 724 -64
rect 730 -65 731 -64
rect 219 -67 220 -66
rect 299 -67 300 -66
rect 303 -67 304 -66
rect 324 -67 325 -66
rect 338 -67 339 -66
rect 548 -67 549 -66
rect 576 -67 577 -66
rect 590 -67 591 -66
rect 604 -67 605 -66
rect 628 -67 629 -66
rect 681 -67 682 -66
rect 723 -67 724 -66
rect 324 -69 325 -68
rect 534 -69 535 -68
rect 555 -69 556 -68
rect 576 -69 577 -68
rect 611 -69 612 -68
rect 618 -69 619 -68
rect 621 -69 622 -68
rect 688 -69 689 -68
rect 373 -71 374 -70
rect 443 -71 444 -70
rect 485 -71 486 -70
rect 548 -71 549 -70
rect 572 -71 573 -70
rect 611 -71 612 -70
rect 614 -71 615 -70
rect 667 -71 668 -70
rect 674 -71 675 -70
rect 681 -71 682 -70
rect 436 -73 437 -72
rect 443 -73 444 -72
rect 457 -73 458 -72
rect 485 -73 486 -72
rect 520 -73 521 -72
rect 639 -73 640 -72
rect 383 -75 384 -74
rect 457 -75 458 -74
rect 541 -75 542 -74
rect 555 -75 556 -74
rect 422 -77 423 -76
rect 436 -77 437 -76
rect 422 -79 423 -78
rect 492 -79 493 -78
rect 429 -81 430 -80
rect 492 -81 493 -80
rect 415 -83 416 -82
rect 429 -83 430 -82
rect 415 -85 416 -84
rect 450 -85 451 -84
rect 331 -87 332 -86
rect 450 -87 451 -86
rect 331 -89 332 -88
rect 359 -89 360 -88
rect 352 -91 353 -90
rect 359 -91 360 -90
rect 352 -93 353 -92
rect 366 -93 367 -92
rect 366 -95 367 -94
rect 394 -95 395 -94
rect 394 -97 395 -96
rect 782 -97 783 -96
rect 114 -108 115 -107
rect 191 -108 192 -107
rect 198 -108 199 -107
rect 296 -108 297 -107
rect 299 -108 300 -107
rect 390 -108 391 -107
rect 471 -108 472 -107
rect 562 -108 563 -107
rect 565 -108 566 -107
rect 695 -108 696 -107
rect 723 -108 724 -107
rect 786 -108 787 -107
rect 793 -108 794 -107
rect 856 -108 857 -107
rect 891 -108 892 -107
rect 919 -108 920 -107
rect 1010 -108 1011 -107
rect 1136 -108 1137 -107
rect 121 -110 122 -109
rect 383 -110 384 -109
rect 387 -110 388 -109
rect 450 -110 451 -109
rect 509 -110 510 -109
rect 562 -110 563 -109
rect 572 -110 573 -109
rect 744 -110 745 -109
rect 782 -110 783 -109
rect 1171 -110 1172 -109
rect 135 -112 136 -111
rect 299 -112 300 -111
rect 334 -112 335 -111
rect 723 -112 724 -111
rect 737 -112 738 -111
rect 842 -112 843 -111
rect 898 -112 899 -111
rect 940 -112 941 -111
rect 1017 -112 1018 -111
rect 1024 -112 1025 -111
rect 142 -114 143 -113
rect 520 -114 521 -113
rect 537 -114 538 -113
rect 821 -114 822 -113
rect 863 -114 864 -113
rect 898 -114 899 -113
rect 149 -116 150 -115
rect 373 -116 374 -115
rect 380 -116 381 -115
rect 541 -116 542 -115
rect 558 -116 559 -115
rect 604 -116 605 -115
rect 611 -116 612 -115
rect 772 -116 773 -115
rect 800 -116 801 -115
rect 877 -116 878 -115
rect 156 -118 157 -117
rect 310 -118 311 -117
rect 369 -118 370 -117
rect 534 -118 535 -117
rect 583 -118 584 -117
rect 590 -118 591 -117
rect 593 -118 594 -117
rect 758 -118 759 -117
rect 807 -118 808 -117
rect 870 -118 871 -117
rect 163 -120 164 -119
rect 205 -120 206 -119
rect 212 -120 213 -119
rect 453 -120 454 -119
rect 516 -120 517 -119
rect 800 -120 801 -119
rect 863 -120 864 -119
rect 1013 -120 1014 -119
rect 170 -122 171 -121
rect 289 -122 290 -121
rect 310 -122 311 -121
rect 408 -122 409 -121
rect 443 -122 444 -121
rect 471 -122 472 -121
rect 614 -122 615 -121
rect 737 -122 738 -121
rect 177 -124 178 -123
rect 229 -124 230 -123
rect 240 -124 241 -123
rect 303 -124 304 -123
rect 408 -124 409 -123
rect 604 -124 605 -123
rect 618 -124 619 -123
rect 793 -124 794 -123
rect 184 -126 185 -125
rect 219 -126 220 -125
rect 226 -126 227 -125
rect 513 -126 514 -125
rect 586 -126 587 -125
rect 618 -126 619 -125
rect 625 -126 626 -125
rect 849 -126 850 -125
rect 191 -128 192 -127
rect 394 -128 395 -127
rect 415 -128 416 -127
rect 443 -128 444 -127
rect 450 -128 451 -127
rect 499 -128 500 -127
rect 513 -128 514 -127
rect 541 -128 542 -127
rect 576 -128 577 -127
rect 625 -128 626 -127
rect 628 -128 629 -127
rect 716 -128 717 -127
rect 205 -130 206 -129
rect 233 -130 234 -129
rect 247 -130 248 -129
rect 373 -130 374 -129
rect 394 -130 395 -129
rect 548 -130 549 -129
rect 639 -130 640 -129
rect 779 -130 780 -129
rect 219 -132 220 -131
rect 324 -132 325 -131
rect 415 -132 416 -131
rect 506 -132 507 -131
rect 639 -132 640 -131
rect 646 -132 647 -131
rect 660 -132 661 -131
rect 765 -132 766 -131
rect 233 -134 234 -133
rect 611 -134 612 -133
rect 667 -134 668 -133
rect 751 -134 752 -133
rect 247 -136 248 -135
rect 257 -136 258 -135
rect 268 -136 269 -135
rect 422 -136 423 -135
rect 464 -136 465 -135
rect 516 -136 517 -135
rect 597 -136 598 -135
rect 646 -136 647 -135
rect 688 -136 689 -135
rect 814 -136 815 -135
rect 271 -138 272 -137
rect 275 -138 276 -137
rect 289 -138 290 -137
rect 530 -138 531 -137
rect 555 -138 556 -137
rect 597 -138 598 -137
rect 632 -138 633 -137
rect 667 -138 668 -137
rect 702 -138 703 -137
rect 807 -138 808 -137
rect 275 -140 276 -139
rect 338 -140 339 -139
rect 390 -140 391 -139
rect 422 -140 423 -139
rect 464 -140 465 -139
rect 527 -140 528 -139
rect 555 -140 556 -139
rect 674 -140 675 -139
rect 702 -140 703 -139
rect 730 -140 731 -139
rect 303 -142 304 -141
rect 523 -142 524 -141
rect 527 -142 528 -141
rect 828 -142 829 -141
rect 324 -144 325 -143
rect 352 -144 353 -143
rect 478 -144 479 -143
rect 660 -144 661 -143
rect 730 -144 731 -143
rect 835 -144 836 -143
rect 338 -146 339 -145
rect 366 -146 367 -145
rect 478 -146 479 -145
rect 485 -146 486 -145
rect 492 -146 493 -145
rect 548 -146 549 -145
rect 632 -146 633 -145
rect 709 -146 710 -145
rect 128 -148 129 -147
rect 366 -148 367 -147
rect 457 -148 458 -147
rect 485 -148 486 -147
rect 492 -148 493 -147
rect 502 -148 503 -147
rect 653 -148 654 -147
rect 688 -148 689 -147
rect 345 -150 346 -149
rect 352 -150 353 -149
rect 436 -150 437 -149
rect 457 -150 458 -149
rect 499 -150 500 -149
rect 576 -150 577 -149
rect 583 -150 584 -149
rect 653 -150 654 -149
rect 656 -150 657 -149
rect 709 -150 710 -149
rect 345 -152 346 -151
rect 401 -152 402 -151
rect 359 -154 360 -153
rect 436 -154 437 -153
rect 359 -156 360 -155
rect 429 -156 430 -155
rect 317 -158 318 -157
rect 429 -158 430 -157
rect 254 -160 255 -159
rect 317 -160 318 -159
rect 401 -160 402 -159
rect 786 -160 787 -159
rect 254 -162 255 -161
rect 331 -162 332 -161
rect 331 -164 332 -163
rect 506 -164 507 -163
rect 72 -175 73 -174
rect 569 -175 570 -174
rect 597 -175 598 -174
rect 600 -175 601 -174
rect 709 -175 710 -174
rect 884 -175 885 -174
rect 898 -175 899 -174
rect 933 -175 934 -174
rect 940 -175 941 -174
rect 989 -175 990 -174
rect 1024 -175 1025 -174
rect 1038 -175 1039 -174
rect 1136 -175 1137 -174
rect 1185 -175 1186 -174
rect 86 -177 87 -176
rect 656 -177 657 -176
rect 751 -177 752 -176
rect 1017 -177 1018 -176
rect 1171 -177 1172 -176
rect 1325 -177 1326 -176
rect 93 -179 94 -178
rect 268 -179 269 -178
rect 275 -179 276 -178
rect 296 -179 297 -178
rect 310 -179 311 -178
rect 453 -179 454 -178
rect 478 -179 479 -178
rect 530 -179 531 -178
rect 548 -179 549 -178
rect 590 -179 591 -178
rect 597 -179 598 -178
rect 632 -179 633 -178
rect 772 -179 773 -178
rect 912 -179 913 -178
rect 919 -179 920 -178
rect 982 -179 983 -178
rect 100 -181 101 -180
rect 198 -181 199 -180
rect 205 -181 206 -180
rect 401 -181 402 -180
rect 446 -181 447 -180
rect 940 -181 941 -180
rect 107 -183 108 -182
rect 415 -183 416 -182
rect 513 -183 514 -182
rect 772 -183 773 -182
rect 793 -183 794 -182
rect 1003 -183 1004 -182
rect 114 -185 115 -184
rect 208 -185 209 -184
rect 222 -185 223 -184
rect 891 -185 892 -184
rect 121 -187 122 -186
rect 236 -187 237 -186
rect 240 -187 241 -186
rect 334 -187 335 -186
rect 401 -187 402 -186
rect 478 -187 479 -186
rect 520 -187 521 -186
rect 730 -187 731 -186
rect 800 -187 801 -186
rect 898 -187 899 -186
rect 121 -189 122 -188
rect 142 -189 143 -188
rect 149 -189 150 -188
rect 569 -189 570 -188
rect 576 -189 577 -188
rect 709 -189 710 -188
rect 716 -189 717 -188
rect 793 -189 794 -188
rect 807 -189 808 -188
rect 926 -189 927 -188
rect 142 -191 143 -190
rect 506 -191 507 -190
rect 523 -191 524 -190
rect 593 -191 594 -190
rect 600 -191 601 -190
rect 632 -191 633 -190
rect 674 -191 675 -190
rect 919 -191 920 -190
rect 149 -193 150 -192
rect 184 -193 185 -192
rect 191 -193 192 -192
rect 527 -193 528 -192
rect 534 -193 535 -192
rect 576 -193 577 -192
rect 625 -193 626 -192
rect 674 -193 675 -192
rect 681 -193 682 -192
rect 716 -193 717 -192
rect 737 -193 738 -192
rect 800 -193 801 -192
rect 814 -193 815 -192
rect 1010 -193 1011 -192
rect 79 -195 80 -194
rect 625 -195 626 -194
rect 681 -195 682 -194
rect 688 -195 689 -194
rect 702 -195 703 -194
rect 737 -195 738 -194
rect 744 -195 745 -194
rect 814 -195 815 -194
rect 821 -195 822 -194
rect 961 -195 962 -194
rect 163 -197 164 -196
rect 275 -197 276 -196
rect 289 -197 290 -196
rect 296 -197 297 -196
rect 310 -197 311 -196
rect 390 -197 391 -196
rect 422 -197 423 -196
rect 513 -197 514 -196
rect 555 -197 556 -196
rect 614 -197 615 -196
rect 667 -197 668 -196
rect 744 -197 745 -196
rect 828 -197 829 -196
rect 947 -197 948 -196
rect 163 -199 164 -198
rect 177 -199 178 -198
rect 184 -199 185 -198
rect 219 -199 220 -198
rect 233 -199 234 -198
rect 415 -199 416 -198
rect 432 -199 433 -198
rect 807 -199 808 -198
rect 835 -199 836 -198
rect 905 -199 906 -198
rect 114 -201 115 -200
rect 219 -201 220 -200
rect 233 -201 234 -200
rect 369 -201 370 -200
rect 436 -201 437 -200
rect 520 -201 521 -200
rect 558 -201 559 -200
rect 653 -201 654 -200
rect 688 -201 689 -200
rect 751 -201 752 -200
rect 765 -201 766 -200
rect 835 -201 836 -200
rect 856 -201 857 -200
rect 968 -201 969 -200
rect 170 -203 171 -202
rect 198 -203 199 -202
rect 243 -203 244 -202
rect 422 -203 423 -202
rect 464 -203 465 -202
rect 534 -203 535 -202
rect 562 -203 563 -202
rect 604 -203 605 -202
rect 618 -203 619 -202
rect 765 -203 766 -202
rect 870 -203 871 -202
rect 975 -203 976 -202
rect 156 -205 157 -204
rect 170 -205 171 -204
rect 177 -205 178 -204
rect 404 -205 405 -204
rect 443 -205 444 -204
rect 464 -205 465 -204
rect 471 -205 472 -204
rect 667 -205 668 -204
rect 702 -205 703 -204
rect 758 -205 759 -204
rect 786 -205 787 -204
rect 870 -205 871 -204
rect 877 -205 878 -204
rect 1024 -205 1025 -204
rect 128 -207 129 -206
rect 443 -207 444 -206
rect 471 -207 472 -206
rect 492 -207 493 -206
rect 607 -207 608 -206
rect 758 -207 759 -206
rect 842 -207 843 -206
rect 877 -207 878 -206
rect 128 -209 129 -208
rect 226 -209 227 -208
rect 229 -209 230 -208
rect 842 -209 843 -208
rect 191 -211 192 -210
rect 205 -211 206 -210
rect 261 -211 262 -210
rect 268 -211 269 -210
rect 289 -211 290 -210
rect 352 -211 353 -210
rect 387 -211 388 -210
rect 786 -211 787 -210
rect 247 -213 248 -212
rect 261 -213 262 -212
rect 331 -213 332 -212
rect 338 -213 339 -212
rect 352 -213 353 -212
rect 366 -213 367 -212
rect 380 -213 381 -212
rect 387 -213 388 -212
rect 394 -213 395 -212
rect 436 -213 437 -212
rect 485 -213 486 -212
rect 506 -213 507 -212
rect 618 -213 619 -212
rect 646 -213 647 -212
rect 660 -213 661 -212
rect 856 -213 857 -212
rect 212 -215 213 -214
rect 338 -215 339 -214
rect 373 -215 374 -214
rect 380 -215 381 -214
rect 394 -215 395 -214
rect 551 -215 552 -214
rect 611 -215 612 -214
rect 660 -215 661 -214
rect 723 -215 724 -214
rect 821 -215 822 -214
rect 212 -217 213 -216
rect 499 -217 500 -216
rect 611 -217 612 -216
rect 954 -217 955 -216
rect 247 -219 248 -218
rect 324 -219 325 -218
rect 359 -219 360 -218
rect 373 -219 374 -218
rect 429 -219 430 -218
rect 646 -219 647 -218
rect 723 -219 724 -218
rect 863 -219 864 -218
rect 135 -221 136 -220
rect 429 -221 430 -220
rect 492 -221 493 -220
rect 541 -221 542 -220
rect 779 -221 780 -220
rect 863 -221 864 -220
rect 135 -223 136 -222
rect 254 -223 255 -222
rect 317 -223 318 -222
rect 331 -223 332 -222
rect 345 -223 346 -222
rect 359 -223 360 -222
rect 499 -223 500 -222
rect 562 -223 563 -222
rect 695 -223 696 -222
rect 779 -223 780 -222
rect 254 -225 255 -224
rect 303 -225 304 -224
rect 317 -225 318 -224
rect 408 -225 409 -224
rect 541 -225 542 -224
rect 639 -225 640 -224
rect 695 -225 696 -224
rect 831 -225 832 -224
rect 303 -227 304 -226
rect 450 -227 451 -226
rect 583 -227 584 -226
rect 639 -227 640 -226
rect 324 -229 325 -228
rect 485 -229 486 -228
rect 583 -229 584 -228
rect 849 -229 850 -228
rect 345 -231 346 -230
rect 408 -231 409 -230
rect 450 -231 451 -230
rect 628 -231 629 -230
rect 849 -231 850 -230
rect 996 -231 997 -230
rect 93 -242 94 -241
rect 485 -242 486 -241
rect 488 -242 489 -241
rect 856 -242 857 -241
rect 884 -242 885 -241
rect 1115 -242 1116 -241
rect 1185 -242 1186 -241
rect 1206 -242 1207 -241
rect 1307 -242 1308 -241
rect 1458 -242 1459 -241
rect 93 -244 94 -243
rect 142 -244 143 -243
rect 145 -244 146 -243
rect 401 -244 402 -243
rect 446 -244 447 -243
rect 492 -244 493 -243
rect 502 -244 503 -243
rect 912 -244 913 -243
rect 919 -244 920 -243
rect 1052 -244 1053 -243
rect 1325 -244 1326 -243
rect 1381 -244 1382 -243
rect 100 -246 101 -245
rect 173 -246 174 -245
rect 177 -246 178 -245
rect 478 -246 479 -245
rect 485 -246 486 -245
rect 747 -246 748 -245
rect 754 -246 755 -245
rect 1080 -246 1081 -245
rect 100 -248 101 -247
rect 236 -248 237 -247
rect 247 -248 248 -247
rect 401 -248 402 -247
rect 453 -248 454 -247
rect 1003 -248 1004 -247
rect 1038 -248 1039 -247
rect 1066 -248 1067 -247
rect 107 -250 108 -249
rect 443 -250 444 -249
rect 492 -250 493 -249
rect 506 -250 507 -249
rect 537 -250 538 -249
rect 1101 -250 1102 -249
rect 107 -252 108 -251
rect 142 -252 143 -251
rect 159 -252 160 -251
rect 257 -252 258 -251
rect 303 -252 304 -251
rect 551 -252 552 -251
rect 600 -252 601 -251
rect 912 -252 913 -251
rect 954 -252 955 -251
rect 1108 -252 1109 -251
rect 128 -254 129 -253
rect 240 -254 241 -253
rect 247 -254 248 -253
rect 366 -254 367 -253
rect 369 -254 370 -253
rect 457 -254 458 -253
rect 506 -254 507 -253
rect 527 -254 528 -253
rect 551 -254 552 -253
rect 618 -254 619 -253
rect 628 -254 629 -253
rect 919 -254 920 -253
rect 968 -254 969 -253
rect 1031 -254 1032 -253
rect 79 -256 80 -255
rect 128 -256 129 -255
rect 138 -256 139 -255
rect 688 -256 689 -255
rect 737 -256 738 -255
rect 751 -256 752 -255
rect 765 -256 766 -255
rect 1094 -256 1095 -255
rect 79 -258 80 -257
rect 149 -258 150 -257
rect 163 -258 164 -257
rect 177 -258 178 -257
rect 191 -258 192 -257
rect 194 -258 195 -257
rect 205 -258 206 -257
rect 226 -258 227 -257
rect 233 -258 234 -257
rect 289 -258 290 -257
rect 303 -258 304 -257
rect 576 -258 577 -257
rect 618 -258 619 -257
rect 628 -258 629 -257
rect 632 -258 633 -257
rect 688 -258 689 -257
rect 716 -258 717 -257
rect 737 -258 738 -257
rect 786 -258 787 -257
rect 856 -258 857 -257
rect 877 -258 878 -257
rect 954 -258 955 -257
rect 975 -258 976 -257
rect 1073 -258 1074 -257
rect 114 -260 115 -259
rect 149 -260 150 -259
rect 163 -260 164 -259
rect 184 -260 185 -259
rect 191 -260 192 -259
rect 219 -260 220 -259
rect 226 -260 227 -259
rect 562 -260 563 -259
rect 632 -260 633 -259
rect 1017 -260 1018 -259
rect 114 -262 115 -261
rect 121 -262 122 -261
rect 170 -262 171 -261
rect 499 -262 500 -261
rect 541 -262 542 -261
rect 562 -262 563 -261
rect 670 -262 671 -261
rect 807 -262 808 -261
rect 821 -262 822 -261
rect 884 -262 885 -261
rect 891 -262 892 -261
rect 1045 -262 1046 -261
rect 121 -264 122 -263
rect 352 -264 353 -263
rect 366 -264 367 -263
rect 373 -264 374 -263
rect 376 -264 377 -263
rect 520 -264 521 -263
rect 541 -264 542 -263
rect 555 -264 556 -263
rect 674 -264 675 -263
rect 968 -264 969 -263
rect 982 -264 983 -263
rect 1038 -264 1039 -263
rect 194 -266 195 -265
rect 219 -266 220 -265
rect 289 -266 290 -265
rect 394 -266 395 -265
rect 450 -266 451 -265
rect 527 -266 528 -265
rect 646 -266 647 -265
rect 674 -266 675 -265
rect 695 -266 696 -265
rect 716 -266 717 -265
rect 779 -266 780 -265
rect 821 -266 822 -265
rect 835 -266 836 -265
rect 891 -266 892 -265
rect 905 -266 906 -265
rect 1003 -266 1004 -265
rect 198 -268 199 -267
rect 576 -268 577 -267
rect 625 -268 626 -267
rect 779 -268 780 -267
rect 793 -268 794 -267
rect 877 -268 878 -267
rect 905 -268 906 -267
rect 1024 -268 1025 -267
rect 198 -270 199 -269
rect 261 -270 262 -269
rect 331 -270 332 -269
rect 352 -270 353 -269
rect 380 -270 381 -269
rect 555 -270 556 -269
rect 646 -270 647 -269
rect 982 -270 983 -269
rect 989 -270 990 -269
rect 1059 -270 1060 -269
rect 208 -272 209 -271
rect 261 -272 262 -271
rect 380 -272 381 -271
rect 1122 -272 1123 -271
rect 86 -274 87 -273
rect 208 -274 209 -273
rect 212 -274 213 -273
rect 331 -274 332 -273
rect 383 -274 384 -273
rect 604 -274 605 -273
rect 709 -274 710 -273
rect 786 -274 787 -273
rect 898 -274 899 -273
rect 989 -274 990 -273
rect 996 -274 997 -273
rect 1087 -274 1088 -273
rect 86 -276 87 -275
rect 429 -276 430 -275
rect 450 -276 451 -275
rect 548 -276 549 -275
rect 604 -276 605 -275
rect 1010 -276 1011 -275
rect 184 -278 185 -277
rect 212 -278 213 -277
rect 387 -278 388 -277
rect 408 -278 409 -277
rect 415 -278 416 -277
rect 429 -278 430 -277
rect 457 -278 458 -277
rect 464 -278 465 -277
rect 478 -278 479 -277
rect 765 -278 766 -277
rect 926 -278 927 -277
rect 1010 -278 1011 -277
rect 187 -280 188 -279
rect 464 -280 465 -279
rect 499 -280 500 -279
rect 597 -280 598 -279
rect 607 -280 608 -279
rect 926 -280 927 -279
rect 933 -280 934 -279
rect 975 -280 976 -279
rect 317 -282 318 -281
rect 415 -282 416 -281
rect 513 -282 514 -281
rect 520 -282 521 -281
rect 534 -282 535 -281
rect 597 -282 598 -281
rect 611 -282 612 -281
rect 709 -282 710 -281
rect 723 -282 724 -281
rect 793 -282 794 -281
rect 842 -282 843 -281
rect 933 -282 934 -281
rect 940 -282 941 -281
rect 1017 -282 1018 -281
rect 65 -284 66 -283
rect 534 -284 535 -283
rect 590 -284 591 -283
rect 611 -284 612 -283
rect 660 -284 661 -283
rect 723 -284 724 -283
rect 744 -284 745 -283
rect 898 -284 899 -283
rect 947 -284 948 -283
rect 996 -284 997 -283
rect 317 -286 318 -285
rect 324 -286 325 -285
rect 387 -286 388 -285
rect 849 -286 850 -285
rect 863 -286 864 -285
rect 940 -286 941 -285
rect 961 -286 962 -285
rect 1024 -286 1025 -285
rect 324 -288 325 -287
rect 345 -288 346 -287
rect 390 -288 391 -287
rect 667 -288 668 -287
rect 744 -288 745 -287
rect 835 -288 836 -287
rect 870 -288 871 -287
rect 947 -288 948 -287
rect 72 -290 73 -289
rect 345 -290 346 -289
rect 394 -290 395 -289
rect 471 -290 472 -289
rect 590 -290 591 -289
rect 870 -290 871 -289
rect 72 -292 73 -291
rect 156 -292 157 -291
rect 275 -292 276 -291
rect 471 -292 472 -291
rect 653 -292 654 -291
rect 660 -292 661 -291
rect 667 -292 668 -291
rect 772 -292 773 -291
rect 800 -292 801 -291
rect 842 -292 843 -291
rect 156 -294 157 -293
rect 254 -294 255 -293
rect 275 -294 276 -293
rect 296 -294 297 -293
rect 411 -294 412 -293
rect 849 -294 850 -293
rect 170 -296 171 -295
rect 800 -296 801 -295
rect 814 -296 815 -295
rect 863 -296 864 -295
rect 254 -298 255 -297
rect 373 -298 374 -297
rect 422 -298 423 -297
rect 513 -298 514 -297
rect 639 -298 640 -297
rect 653 -298 654 -297
rect 730 -298 731 -297
rect 814 -298 815 -297
rect 828 -298 829 -297
rect 961 -298 962 -297
rect 282 -300 283 -299
rect 296 -300 297 -299
rect 422 -300 423 -299
rect 436 -300 437 -299
rect 481 -300 482 -299
rect 772 -300 773 -299
rect 135 -302 136 -301
rect 282 -302 283 -301
rect 583 -302 584 -301
rect 639 -302 640 -301
rect 681 -302 682 -301
rect 730 -302 731 -301
rect 758 -302 759 -301
rect 828 -302 829 -301
rect 243 -304 244 -303
rect 436 -304 437 -303
rect 446 -304 447 -303
rect 758 -304 759 -303
rect 569 -306 570 -305
rect 583 -306 584 -305
rect 681 -306 682 -305
rect 702 -306 703 -305
rect 338 -308 339 -307
rect 569 -308 570 -307
rect 695 -308 696 -307
rect 702 -308 703 -307
rect 338 -310 339 -309
rect 359 -310 360 -309
rect 310 -312 311 -311
rect 359 -312 360 -311
rect 310 -314 311 -313
rect 807 -314 808 -313
rect 65 -325 66 -324
rect 380 -325 381 -324
rect 446 -325 447 -324
rect 576 -325 577 -324
rect 590 -325 591 -324
rect 1094 -325 1095 -324
rect 1101 -325 1102 -324
rect 1213 -325 1214 -324
rect 1381 -325 1382 -324
rect 1409 -325 1410 -324
rect 1458 -325 1459 -324
rect 1521 -325 1522 -324
rect 72 -327 73 -326
rect 362 -327 363 -326
rect 369 -327 370 -326
rect 569 -327 570 -326
rect 597 -327 598 -326
rect 898 -327 899 -326
rect 912 -327 913 -326
rect 1150 -327 1151 -326
rect 1171 -327 1172 -326
rect 1223 -327 1224 -326
rect 72 -329 73 -328
rect 121 -329 122 -328
rect 135 -329 136 -328
rect 289 -329 290 -328
rect 345 -329 346 -328
rect 534 -329 535 -328
rect 548 -329 549 -328
rect 1052 -329 1053 -328
rect 1059 -329 1060 -328
rect 1164 -329 1165 -328
rect 1199 -329 1200 -328
rect 1307 -329 1308 -328
rect 79 -331 80 -330
rect 187 -331 188 -330
rect 205 -331 206 -330
rect 1108 -331 1109 -330
rect 1122 -331 1123 -330
rect 1388 -331 1389 -330
rect 58 -333 59 -332
rect 205 -333 206 -332
rect 250 -333 251 -332
rect 534 -333 535 -332
rect 541 -333 542 -332
rect 548 -333 549 -332
rect 551 -333 552 -332
rect 968 -333 969 -332
rect 989 -333 990 -332
rect 1122 -333 1123 -332
rect 79 -335 80 -334
rect 149 -335 150 -334
rect 166 -335 167 -334
rect 576 -335 577 -334
rect 597 -335 598 -334
rect 789 -335 790 -334
rect 807 -335 808 -334
rect 898 -335 899 -334
rect 926 -335 927 -334
rect 989 -335 990 -334
rect 1003 -335 1004 -334
rect 1129 -335 1130 -334
rect 86 -337 87 -336
rect 383 -337 384 -336
rect 478 -337 479 -336
rect 541 -337 542 -336
rect 565 -337 566 -336
rect 1178 -337 1179 -336
rect 86 -339 87 -338
rect 593 -339 594 -338
rect 604 -339 605 -338
rect 618 -339 619 -338
rect 625 -339 626 -338
rect 1045 -339 1046 -338
rect 1066 -339 1067 -338
rect 1108 -339 1109 -338
rect 93 -341 94 -340
rect 537 -341 538 -340
rect 618 -341 619 -340
rect 660 -341 661 -340
rect 667 -341 668 -340
rect 688 -341 689 -340
rect 702 -341 703 -340
rect 744 -341 745 -340
rect 821 -341 822 -340
rect 968 -341 969 -340
rect 975 -341 976 -340
rect 1045 -341 1046 -340
rect 1073 -341 1074 -340
rect 1185 -341 1186 -340
rect 93 -343 94 -342
rect 418 -343 419 -342
rect 464 -343 465 -342
rect 604 -343 605 -342
rect 625 -343 626 -342
rect 807 -343 808 -342
rect 835 -343 836 -342
rect 912 -343 913 -342
rect 961 -343 962 -342
rect 1003 -343 1004 -342
rect 1017 -343 1018 -342
rect 1143 -343 1144 -342
rect 100 -345 101 -344
rect 187 -345 188 -344
rect 191 -345 192 -344
rect 383 -345 384 -344
rect 464 -345 465 -344
rect 555 -345 556 -344
rect 583 -345 584 -344
rect 660 -345 661 -344
rect 702 -345 703 -344
rect 786 -345 787 -344
rect 856 -345 857 -344
rect 926 -345 927 -344
rect 947 -345 948 -344
rect 1017 -345 1018 -344
rect 1024 -345 1025 -344
rect 1094 -345 1095 -344
rect 100 -347 101 -346
rect 156 -347 157 -346
rect 170 -347 171 -346
rect 849 -347 850 -346
rect 856 -347 857 -346
rect 905 -347 906 -346
rect 947 -347 948 -346
rect 1010 -347 1011 -346
rect 1031 -347 1032 -346
rect 1136 -347 1137 -346
rect 121 -349 122 -348
rect 128 -349 129 -348
rect 149 -349 150 -348
rect 310 -349 311 -348
rect 345 -349 346 -348
rect 450 -349 451 -348
rect 495 -349 496 -348
rect 513 -349 514 -348
rect 555 -349 556 -348
rect 653 -349 654 -348
rect 758 -349 759 -348
rect 849 -349 850 -348
rect 870 -349 871 -348
rect 1052 -349 1053 -348
rect 1080 -349 1081 -348
rect 1192 -349 1193 -348
rect 128 -351 129 -350
rect 303 -351 304 -350
rect 310 -351 311 -350
rect 359 -351 360 -350
rect 373 -351 374 -350
rect 485 -351 486 -350
rect 506 -351 507 -350
rect 590 -351 591 -350
rect 628 -351 629 -350
rect 730 -351 731 -350
rect 765 -351 766 -350
rect 821 -351 822 -350
rect 884 -351 885 -350
rect 961 -351 962 -350
rect 982 -351 983 -350
rect 1066 -351 1067 -350
rect 1080 -351 1081 -350
rect 1115 -351 1116 -350
rect 173 -353 174 -352
rect 569 -353 570 -352
rect 583 -353 584 -352
rect 765 -353 766 -352
rect 772 -353 773 -352
rect 1031 -353 1032 -352
rect 1038 -353 1039 -352
rect 1059 -353 1060 -352
rect 1087 -353 1088 -352
rect 1157 -353 1158 -352
rect 107 -355 108 -354
rect 1087 -355 1088 -354
rect 107 -357 108 -356
rect 114 -357 115 -356
rect 173 -357 174 -356
rect 506 -357 507 -356
rect 513 -357 514 -356
rect 527 -357 528 -356
rect 632 -357 633 -356
rect 649 -357 650 -356
rect 709 -357 710 -356
rect 772 -357 773 -356
rect 786 -357 787 -356
rect 1101 -357 1102 -356
rect 114 -359 115 -358
rect 471 -359 472 -358
rect 481 -359 482 -358
rect 653 -359 654 -358
rect 730 -359 731 -358
rect 800 -359 801 -358
rect 814 -359 815 -358
rect 905 -359 906 -358
rect 919 -359 920 -358
rect 982 -359 983 -358
rect 996 -359 997 -358
rect 1024 -359 1025 -358
rect 184 -361 185 -360
rect 1073 -361 1074 -360
rect 138 -363 139 -362
rect 184 -363 185 -362
rect 194 -363 195 -362
rect 485 -363 486 -362
rect 520 -363 521 -362
rect 527 -363 528 -362
rect 572 -363 573 -362
rect 814 -363 815 -362
rect 828 -363 829 -362
rect 884 -363 885 -362
rect 891 -363 892 -362
rect 975 -363 976 -362
rect 247 -365 248 -364
rect 758 -365 759 -364
rect 793 -365 794 -364
rect 828 -365 829 -364
rect 842 -365 843 -364
rect 891 -365 892 -364
rect 940 -365 941 -364
rect 1010 -365 1011 -364
rect 156 -367 157 -366
rect 247 -367 248 -366
rect 282 -367 283 -366
rect 390 -367 391 -366
rect 415 -367 416 -366
rect 520 -367 521 -366
rect 646 -367 647 -366
rect 835 -367 836 -366
rect 842 -367 843 -366
rect 933 -367 934 -366
rect 954 -367 955 -366
rect 1038 -367 1039 -366
rect 142 -369 143 -368
rect 415 -369 416 -368
rect 436 -369 437 -368
rect 450 -369 451 -368
rect 586 -369 587 -368
rect 933 -369 934 -368
rect 142 -371 143 -370
rect 163 -371 164 -370
rect 233 -371 234 -370
rect 282 -371 283 -370
rect 289 -371 290 -370
rect 691 -371 692 -370
rect 723 -371 724 -370
rect 793 -371 794 -370
rect 863 -371 864 -370
rect 940 -371 941 -370
rect 233 -373 234 -372
rect 635 -373 636 -372
rect 670 -373 671 -372
rect 996 -373 997 -372
rect 303 -375 304 -374
rect 338 -375 339 -374
rect 376 -375 377 -374
rect 471 -375 472 -374
rect 737 -375 738 -374
rect 919 -375 920 -374
rect 261 -377 262 -376
rect 338 -377 339 -376
rect 387 -377 388 -376
rect 800 -377 801 -376
rect 877 -377 878 -376
rect 954 -377 955 -376
rect 212 -379 213 -378
rect 261 -379 262 -378
rect 313 -379 314 -378
rect 387 -379 388 -378
rect 408 -379 409 -378
rect 723 -379 724 -378
rect 747 -379 748 -378
rect 1115 -379 1116 -378
rect 212 -381 213 -380
rect 219 -381 220 -380
rect 366 -381 367 -380
rect 408 -381 409 -380
rect 436 -381 437 -380
rect 611 -381 612 -380
rect 716 -381 717 -380
rect 737 -381 738 -380
rect 779 -381 780 -380
rect 863 -381 864 -380
rect 177 -383 178 -382
rect 219 -383 220 -382
rect 443 -383 444 -382
rect 709 -383 710 -382
rect 716 -383 717 -382
rect 870 -383 871 -382
rect 177 -385 178 -384
rect 254 -385 255 -384
rect 422 -385 423 -384
rect 443 -385 444 -384
rect 562 -385 563 -384
rect 611 -385 612 -384
rect 751 -385 752 -384
rect 779 -385 780 -384
rect 240 -387 241 -386
rect 422 -387 423 -386
rect 600 -387 601 -386
rect 877 -387 878 -386
rect 240 -389 241 -388
rect 394 -389 395 -388
rect 632 -389 633 -388
rect 751 -389 752 -388
rect 254 -391 255 -390
rect 268 -391 269 -390
rect 394 -391 395 -390
rect 401 -391 402 -390
rect 198 -393 199 -392
rect 268 -393 269 -392
rect 401 -393 402 -392
rect 695 -393 696 -392
rect 198 -395 199 -394
rect 492 -395 493 -394
rect 681 -395 682 -394
rect 695 -395 696 -394
rect 275 -397 276 -396
rect 492 -397 493 -396
rect 639 -397 640 -396
rect 681 -397 682 -396
rect 275 -399 276 -398
rect 324 -399 325 -398
rect 639 -399 640 -398
rect 674 -399 675 -398
rect 324 -401 325 -400
rect 331 -401 332 -400
rect 499 -401 500 -400
rect 674 -401 675 -400
rect 226 -403 227 -402
rect 499 -403 500 -402
rect 226 -405 227 -404
rect 317 -405 318 -404
rect 331 -405 332 -404
rect 352 -405 353 -404
rect 296 -407 297 -406
rect 317 -407 318 -406
rect 352 -407 353 -406
rect 457 -407 458 -406
rect 208 -409 209 -408
rect 457 -409 458 -408
rect 296 -411 297 -410
rect 429 -411 430 -410
rect 429 -413 430 -412
rect 688 -413 689 -412
rect 51 -424 52 -423
rect 187 -424 188 -423
rect 194 -424 195 -423
rect 758 -424 759 -423
rect 838 -424 839 -423
rect 1213 -424 1214 -423
rect 1388 -424 1389 -423
rect 1486 -424 1487 -423
rect 1521 -424 1522 -423
rect 1542 -424 1543 -423
rect 58 -426 59 -425
rect 145 -426 146 -425
rect 149 -426 150 -425
rect 212 -426 213 -425
rect 250 -426 251 -425
rect 317 -426 318 -425
rect 359 -426 360 -425
rect 590 -426 591 -425
rect 611 -426 612 -425
rect 621 -426 622 -425
rect 656 -426 657 -425
rect 730 -426 731 -425
rect 754 -426 755 -425
rect 1122 -426 1123 -425
rect 1157 -426 1158 -425
rect 1227 -426 1228 -425
rect 1409 -426 1410 -425
rect 1430 -426 1431 -425
rect 65 -428 66 -427
rect 121 -428 122 -427
rect 124 -428 125 -427
rect 1143 -428 1144 -427
rect 1185 -428 1186 -427
rect 1213 -428 1214 -427
rect 72 -430 73 -429
rect 425 -430 426 -429
rect 450 -430 451 -429
rect 541 -430 542 -429
rect 544 -430 545 -429
rect 793 -430 794 -429
rect 919 -430 920 -429
rect 1234 -430 1235 -429
rect 72 -432 73 -431
rect 562 -432 563 -431
rect 572 -432 573 -431
rect 702 -432 703 -431
rect 737 -432 738 -431
rect 793 -432 794 -431
rect 870 -432 871 -431
rect 919 -432 920 -431
rect 1073 -432 1074 -431
rect 1157 -432 1158 -431
rect 1192 -432 1193 -431
rect 1241 -432 1242 -431
rect 86 -434 87 -433
rect 173 -434 174 -433
rect 177 -434 178 -433
rect 390 -434 391 -433
rect 415 -434 416 -433
rect 520 -434 521 -433
rect 541 -434 542 -433
rect 674 -434 675 -433
rect 688 -434 689 -433
rect 842 -434 843 -433
rect 1031 -434 1032 -433
rect 1073 -434 1074 -433
rect 1080 -434 1081 -433
rect 1255 -434 1256 -433
rect 86 -436 87 -435
rect 107 -436 108 -435
rect 114 -436 115 -435
rect 149 -436 150 -435
rect 163 -436 164 -435
rect 422 -436 423 -435
rect 450 -436 451 -435
rect 551 -436 552 -435
rect 558 -436 559 -435
rect 618 -436 619 -435
rect 628 -436 629 -435
rect 702 -436 703 -435
rect 821 -436 822 -435
rect 870 -436 871 -435
rect 1108 -436 1109 -435
rect 1185 -436 1186 -435
rect 1206 -436 1207 -435
rect 1223 -436 1224 -435
rect 93 -438 94 -437
rect 684 -438 685 -437
rect 691 -438 692 -437
rect 1129 -438 1130 -437
rect 1136 -438 1137 -437
rect 1143 -438 1144 -437
rect 1164 -438 1165 -437
rect 1192 -438 1193 -437
rect 93 -440 94 -439
rect 100 -440 101 -439
rect 114 -440 115 -439
rect 436 -440 437 -439
rect 464 -440 465 -439
rect 520 -440 521 -439
rect 548 -440 549 -439
rect 562 -440 563 -439
rect 583 -440 584 -439
rect 968 -440 969 -439
rect 1101 -440 1102 -439
rect 1129 -440 1130 -439
rect 1164 -440 1165 -439
rect 1199 -440 1200 -439
rect 100 -442 101 -441
rect 198 -442 199 -441
rect 212 -442 213 -441
rect 275 -442 276 -441
rect 296 -442 297 -441
rect 586 -442 587 -441
rect 590 -442 591 -441
rect 646 -442 647 -441
rect 663 -442 664 -441
rect 786 -442 787 -441
rect 824 -442 825 -441
rect 1080 -442 1081 -441
rect 1115 -442 1116 -441
rect 1122 -442 1123 -441
rect 1171 -442 1172 -441
rect 1206 -442 1207 -441
rect 121 -444 122 -443
rect 1087 -444 1088 -443
rect 1094 -444 1095 -443
rect 1115 -444 1116 -443
rect 1150 -444 1151 -443
rect 1171 -444 1172 -443
rect 135 -446 136 -445
rect 492 -446 493 -445
rect 495 -446 496 -445
rect 1108 -446 1109 -445
rect 107 -448 108 -447
rect 135 -448 136 -447
rect 138 -448 139 -447
rect 845 -448 846 -447
rect 852 -448 853 -447
rect 1031 -448 1032 -447
rect 1045 -448 1046 -447
rect 1087 -448 1088 -447
rect 142 -450 143 -449
rect 163 -450 164 -449
rect 166 -450 167 -449
rect 247 -450 248 -449
rect 257 -450 258 -449
rect 338 -450 339 -449
rect 359 -450 360 -449
rect 513 -450 514 -449
rect 548 -450 549 -449
rect 604 -450 605 -449
rect 632 -450 633 -449
rect 1150 -450 1151 -449
rect 152 -452 153 -451
rect 338 -452 339 -451
rect 366 -452 367 -451
rect 730 -452 731 -451
rect 947 -452 948 -451
rect 1094 -452 1095 -451
rect 166 -454 167 -453
rect 1220 -454 1221 -453
rect 170 -456 171 -455
rect 299 -456 300 -455
rect 317 -456 318 -455
rect 324 -456 325 -455
rect 366 -456 367 -455
rect 569 -456 570 -455
rect 632 -456 633 -455
rect 1251 -456 1252 -455
rect 177 -458 178 -457
rect 625 -458 626 -457
rect 667 -458 668 -457
rect 758 -458 759 -457
rect 905 -458 906 -457
rect 947 -458 948 -457
rect 968 -458 969 -457
rect 982 -458 983 -457
rect 1024 -458 1025 -457
rect 1101 -458 1102 -457
rect 184 -460 185 -459
rect 219 -460 220 -459
rect 247 -460 248 -459
rect 593 -460 594 -459
rect 667 -460 668 -459
rect 751 -460 752 -459
rect 835 -460 836 -459
rect 905 -460 906 -459
rect 961 -460 962 -459
rect 982 -460 983 -459
rect 989 -460 990 -459
rect 1024 -460 1025 -459
rect 1038 -460 1039 -459
rect 1045 -460 1046 -459
rect 191 -462 192 -461
rect 194 -462 195 -461
rect 219 -462 220 -461
rect 352 -462 353 -461
rect 380 -462 381 -461
rect 604 -462 605 -461
rect 695 -462 696 -461
rect 737 -462 738 -461
rect 779 -462 780 -461
rect 835 -462 836 -461
rect 898 -462 899 -461
rect 989 -462 990 -461
rect 1017 -462 1018 -461
rect 1038 -462 1039 -461
rect 142 -464 143 -463
rect 779 -464 780 -463
rect 814 -464 815 -463
rect 898 -464 899 -463
rect 954 -464 955 -463
rect 961 -464 962 -463
rect 1010 -464 1011 -463
rect 1017 -464 1018 -463
rect 191 -466 192 -465
rect 674 -466 675 -465
rect 698 -466 699 -465
rect 1052 -466 1053 -465
rect 261 -468 262 -467
rect 324 -468 325 -467
rect 331 -468 332 -467
rect 352 -468 353 -467
rect 383 -468 384 -467
rect 394 -468 395 -467
rect 401 -468 402 -467
rect 436 -468 437 -467
rect 464 -468 465 -467
rect 660 -468 661 -467
rect 723 -468 724 -467
rect 1199 -468 1200 -467
rect 261 -470 262 -469
rect 310 -470 311 -469
rect 345 -470 346 -469
rect 380 -470 381 -469
rect 394 -470 395 -469
rect 408 -470 409 -469
rect 415 -470 416 -469
rect 618 -470 619 -469
rect 726 -470 727 -469
rect 1136 -470 1137 -469
rect 275 -472 276 -471
rect 282 -472 283 -471
rect 296 -472 297 -471
rect 387 -472 388 -471
rect 408 -472 409 -471
rect 821 -472 822 -471
rect 877 -472 878 -471
rect 1010 -472 1011 -471
rect 156 -474 157 -473
rect 282 -474 283 -473
rect 303 -474 304 -473
rect 331 -474 332 -473
rect 345 -474 346 -473
rect 467 -474 468 -473
rect 471 -474 472 -473
rect 513 -474 514 -473
rect 569 -474 570 -473
rect 751 -474 752 -473
rect 765 -474 766 -473
rect 814 -474 815 -473
rect 940 -474 941 -473
rect 954 -474 955 -473
rect 1003 -474 1004 -473
rect 1052 -474 1053 -473
rect 198 -476 199 -475
rect 387 -476 388 -475
rect 418 -476 419 -475
rect 716 -476 717 -475
rect 744 -476 745 -475
rect 765 -476 766 -475
rect 800 -476 801 -475
rect 877 -476 878 -475
rect 912 -476 913 -475
rect 1003 -476 1004 -475
rect 303 -478 304 -477
rect 649 -478 650 -477
rect 653 -478 654 -477
rect 744 -478 745 -477
rect 772 -478 773 -477
rect 800 -478 801 -477
rect 863 -478 864 -477
rect 940 -478 941 -477
rect 310 -480 311 -479
rect 404 -480 405 -479
rect 422 -480 423 -479
rect 681 -480 682 -479
rect 807 -480 808 -479
rect 863 -480 864 -479
rect 884 -480 885 -479
rect 912 -480 913 -479
rect 429 -482 430 -481
rect 471 -482 472 -481
rect 478 -482 479 -481
rect 611 -482 612 -481
rect 653 -482 654 -481
rect 688 -482 689 -481
rect 709 -482 710 -481
rect 807 -482 808 -481
rect 828 -482 829 -481
rect 884 -482 885 -481
rect 226 -484 227 -483
rect 429 -484 430 -483
rect 478 -484 479 -483
rect 499 -484 500 -483
rect 506 -484 507 -483
rect 583 -484 584 -483
rect 597 -484 598 -483
rect 828 -484 829 -483
rect 226 -486 227 -485
rect 240 -486 241 -485
rect 373 -486 374 -485
rect 506 -486 507 -485
rect 534 -486 535 -485
rect 709 -486 710 -485
rect 205 -488 206 -487
rect 240 -488 241 -487
rect 373 -488 374 -487
rect 443 -488 444 -487
rect 485 -488 486 -487
rect 597 -488 598 -487
rect 681 -488 682 -487
rect 1178 -488 1179 -487
rect 128 -490 129 -489
rect 485 -490 486 -489
rect 499 -490 500 -489
rect 719 -490 720 -489
rect 1059 -490 1060 -489
rect 1178 -490 1179 -489
rect 128 -492 129 -491
rect 362 -492 363 -491
rect 443 -492 444 -491
rect 457 -492 458 -491
rect 527 -492 528 -491
rect 534 -492 535 -491
rect 555 -492 556 -491
rect 772 -492 773 -491
rect 1059 -492 1060 -491
rect 1066 -492 1067 -491
rect 205 -494 206 -493
rect 233 -494 234 -493
rect 289 -494 290 -493
rect 527 -494 528 -493
rect 555 -494 556 -493
rect 625 -494 626 -493
rect 975 -494 976 -493
rect 1066 -494 1067 -493
rect 268 -496 269 -495
rect 289 -496 290 -495
rect 457 -496 458 -495
rect 789 -496 790 -495
rect 933 -496 934 -495
rect 975 -496 976 -495
rect 254 -498 255 -497
rect 268 -498 269 -497
rect 576 -498 577 -497
rect 723 -498 724 -497
rect 926 -498 927 -497
rect 933 -498 934 -497
rect 156 -500 157 -499
rect 254 -500 255 -499
rect 576 -500 577 -499
rect 639 -500 640 -499
rect 849 -500 850 -499
rect 926 -500 927 -499
rect 369 -502 370 -501
rect 639 -502 640 -501
rect 44 -513 45 -512
rect 86 -513 87 -512
rect 93 -513 94 -512
rect 1388 -513 1389 -512
rect 1419 -513 1420 -512
rect 1619 -513 1620 -512
rect 58 -515 59 -514
rect 646 -515 647 -514
rect 649 -515 650 -514
rect 1262 -515 1263 -514
rect 1430 -515 1431 -514
rect 1458 -515 1459 -514
rect 1486 -515 1487 -514
rect 1528 -515 1529 -514
rect 1542 -515 1543 -514
rect 1549 -515 1550 -514
rect 58 -517 59 -516
rect 747 -517 748 -516
rect 751 -517 752 -516
rect 1073 -517 1074 -516
rect 1087 -517 1088 -516
rect 1220 -517 1221 -516
rect 1227 -517 1228 -516
rect 1437 -517 1438 -516
rect 65 -519 66 -518
rect 191 -519 192 -518
rect 254 -519 255 -518
rect 380 -519 381 -518
rect 387 -519 388 -518
rect 1157 -519 1158 -518
rect 1178 -519 1179 -518
rect 1360 -519 1361 -518
rect 65 -521 66 -520
rect 236 -521 237 -520
rect 264 -521 265 -520
rect 1318 -521 1319 -520
rect 72 -523 73 -522
rect 327 -523 328 -522
rect 401 -523 402 -522
rect 569 -523 570 -522
rect 590 -523 591 -522
rect 849 -523 850 -522
rect 863 -523 864 -522
rect 1451 -523 1452 -522
rect 72 -525 73 -524
rect 660 -525 661 -524
rect 663 -525 664 -524
rect 898 -525 899 -524
rect 905 -525 906 -524
rect 1332 -525 1333 -524
rect 86 -527 87 -526
rect 149 -527 150 -526
rect 156 -527 157 -526
rect 380 -527 381 -526
rect 425 -527 426 -526
rect 569 -527 570 -526
rect 593 -527 594 -526
rect 1066 -527 1067 -526
rect 1115 -527 1116 -526
rect 1304 -527 1305 -526
rect 93 -529 94 -528
rect 233 -529 234 -528
rect 268 -529 269 -528
rect 292 -529 293 -528
rect 296 -529 297 -528
rect 425 -529 426 -528
rect 450 -529 451 -528
rect 590 -529 591 -528
rect 618 -529 619 -528
rect 1444 -529 1445 -528
rect 121 -531 122 -530
rect 390 -531 391 -530
rect 429 -531 430 -530
rect 450 -531 451 -530
rect 527 -531 528 -530
rect 618 -531 619 -530
rect 621 -531 622 -530
rect 1374 -531 1375 -530
rect 128 -533 129 -532
rect 698 -533 699 -532
rect 730 -533 731 -532
rect 803 -533 804 -532
rect 821 -533 822 -532
rect 1465 -533 1466 -532
rect 128 -535 129 -534
rect 205 -535 206 -534
rect 296 -535 297 -534
rect 642 -535 643 -534
rect 646 -535 647 -534
rect 1017 -535 1018 -534
rect 1024 -535 1025 -534
rect 1430 -535 1431 -534
rect 124 -537 125 -536
rect 205 -537 206 -536
rect 299 -537 300 -536
rect 506 -537 507 -536
rect 534 -537 535 -536
rect 548 -537 549 -536
rect 555 -537 556 -536
rect 765 -537 766 -536
rect 789 -537 790 -536
rect 1283 -537 1284 -536
rect 135 -539 136 -538
rect 656 -539 657 -538
rect 660 -539 661 -538
rect 1223 -539 1224 -538
rect 1241 -539 1242 -538
rect 1251 -539 1252 -538
rect 142 -541 143 -540
rect 184 -541 185 -540
rect 191 -541 192 -540
rect 226 -541 227 -540
rect 359 -541 360 -540
rect 527 -541 528 -540
rect 555 -541 556 -540
rect 709 -541 710 -540
rect 716 -541 717 -540
rect 821 -541 822 -540
rect 856 -541 857 -540
rect 898 -541 899 -540
rect 933 -541 934 -540
rect 1290 -541 1291 -540
rect 142 -543 143 -542
rect 457 -543 458 -542
rect 471 -543 472 -542
rect 534 -543 535 -542
rect 625 -543 626 -542
rect 716 -543 717 -542
rect 744 -543 745 -542
rect 863 -543 864 -542
rect 873 -543 874 -542
rect 989 -543 990 -542
rect 1010 -543 1011 -542
rect 1087 -543 1088 -542
rect 1122 -543 1123 -542
rect 1353 -543 1354 -542
rect 114 -545 115 -544
rect 625 -545 626 -544
rect 653 -545 654 -544
rect 1094 -545 1095 -544
rect 1129 -545 1130 -544
rect 1241 -545 1242 -544
rect 100 -547 101 -546
rect 114 -547 115 -546
rect 145 -547 146 -546
rect 1423 -547 1424 -546
rect 100 -549 101 -548
rect 107 -549 108 -548
rect 149 -549 150 -548
rect 289 -549 290 -548
rect 359 -549 360 -548
rect 394 -549 395 -548
rect 471 -549 472 -548
rect 583 -549 584 -548
rect 632 -549 633 -548
rect 653 -549 654 -548
rect 667 -549 668 -548
rect 905 -549 906 -548
rect 919 -549 920 -548
rect 989 -549 990 -548
rect 1017 -549 1018 -548
rect 1164 -549 1165 -548
rect 1185 -549 1186 -548
rect 1311 -549 1312 -548
rect 156 -551 157 -550
rect 649 -551 650 -550
rect 674 -551 675 -550
rect 751 -551 752 -550
rect 754 -551 755 -550
rect 1269 -551 1270 -550
rect 110 -553 111 -552
rect 674 -553 675 -552
rect 684 -553 685 -552
rect 1248 -553 1249 -552
rect 163 -555 164 -554
rect 1339 -555 1340 -554
rect 163 -557 164 -556
rect 233 -557 234 -556
rect 268 -557 269 -556
rect 457 -557 458 -556
rect 478 -557 479 -556
rect 632 -557 633 -556
rect 684 -557 685 -556
rect 1003 -557 1004 -556
rect 1024 -557 1025 -556
rect 1255 -557 1256 -556
rect 166 -559 167 -558
rect 247 -559 248 -558
rect 355 -559 356 -558
rect 583 -559 584 -558
rect 611 -559 612 -558
rect 667 -559 668 -558
rect 688 -559 689 -558
rect 765 -559 766 -558
rect 800 -559 801 -558
rect 1115 -559 1116 -558
rect 1143 -559 1144 -558
rect 1367 -559 1368 -558
rect 184 -561 185 -560
rect 303 -561 304 -560
rect 373 -561 374 -560
rect 429 -561 430 -560
rect 443 -561 444 -560
rect 611 -561 612 -560
rect 698 -561 699 -560
rect 1234 -561 1235 -560
rect 194 -563 195 -562
rect 1234 -563 1235 -562
rect 219 -565 220 -564
rect 373 -565 374 -564
rect 394 -565 395 -564
rect 597 -565 598 -564
rect 702 -565 703 -564
rect 709 -565 710 -564
rect 744 -565 745 -564
rect 1276 -565 1277 -564
rect 219 -567 220 -566
rect 345 -567 346 -566
rect 366 -567 367 -566
rect 443 -567 444 -566
rect 478 -567 479 -566
rect 1227 -567 1228 -566
rect 198 -569 199 -568
rect 345 -569 346 -568
rect 366 -569 367 -568
rect 415 -569 416 -568
rect 485 -569 486 -568
rect 702 -569 703 -568
rect 758 -569 759 -568
rect 856 -569 857 -568
rect 884 -569 885 -568
rect 933 -569 934 -568
rect 954 -569 955 -568
rect 1003 -569 1004 -568
rect 1034 -569 1035 -568
rect 1094 -569 1095 -568
rect 1108 -569 1109 -568
rect 1164 -569 1165 -568
rect 1171 -569 1172 -568
rect 1185 -569 1186 -568
rect 1192 -569 1193 -568
rect 1381 -569 1382 -568
rect 226 -571 227 -570
rect 324 -571 325 -570
rect 495 -571 496 -570
rect 688 -571 689 -570
rect 761 -571 762 -570
rect 1192 -571 1193 -570
rect 1199 -571 1200 -570
rect 1395 -571 1396 -570
rect 247 -573 248 -572
rect 331 -573 332 -572
rect 506 -573 507 -572
rect 513 -573 514 -572
rect 562 -573 563 -572
rect 597 -573 598 -572
rect 828 -573 829 -572
rect 884 -573 885 -572
rect 891 -573 892 -572
rect 1010 -573 1011 -572
rect 1031 -573 1032 -572
rect 1199 -573 1200 -572
rect 1206 -573 1207 -572
rect 1325 -573 1326 -572
rect 303 -575 304 -574
rect 758 -575 759 -574
rect 786 -575 787 -574
rect 828 -575 829 -574
rect 835 -575 836 -574
rect 891 -575 892 -574
rect 926 -575 927 -574
rect 954 -575 955 -574
rect 961 -575 962 -574
rect 1073 -575 1074 -574
rect 1080 -575 1081 -574
rect 1255 -575 1256 -574
rect 310 -577 311 -576
rect 415 -577 416 -576
rect 481 -577 482 -576
rect 926 -577 927 -576
rect 968 -577 969 -576
rect 1157 -577 1158 -576
rect 1213 -577 1214 -576
rect 1409 -577 1410 -576
rect 240 -579 241 -578
rect 310 -579 311 -578
rect 324 -579 325 -578
rect 1122 -579 1123 -578
rect 1136 -579 1137 -578
rect 1206 -579 1207 -578
rect 240 -581 241 -580
rect 282 -581 283 -580
rect 331 -581 332 -580
rect 460 -581 461 -580
rect 492 -581 493 -580
rect 513 -581 514 -580
rect 723 -581 724 -580
rect 835 -581 836 -580
rect 842 -581 843 -580
rect 919 -581 920 -580
rect 940 -581 941 -580
rect 968 -581 969 -580
rect 975 -581 976 -580
rect 1143 -581 1144 -580
rect 1150 -581 1151 -580
rect 1346 -581 1347 -580
rect 261 -583 262 -582
rect 282 -583 283 -582
rect 317 -583 318 -582
rect 492 -583 493 -582
rect 499 -583 500 -582
rect 1213 -583 1214 -582
rect 79 -585 80 -584
rect 261 -585 262 -584
rect 275 -585 276 -584
rect 317 -585 318 -584
rect 576 -585 577 -584
rect 975 -585 976 -584
rect 982 -585 983 -584
rect 1402 -585 1403 -584
rect 79 -587 80 -586
rect 485 -587 486 -586
rect 639 -587 640 -586
rect 723 -587 724 -586
rect 824 -587 825 -586
rect 1080 -587 1081 -586
rect 1101 -587 1102 -586
rect 1150 -587 1151 -586
rect 275 -589 276 -588
rect 422 -589 423 -588
rect 436 -589 437 -588
rect 576 -589 577 -588
rect 639 -589 640 -588
rect 772 -589 773 -588
rect 870 -589 871 -588
rect 961 -589 962 -588
rect 996 -589 997 -588
rect 1108 -589 1109 -588
rect 51 -591 52 -590
rect 422 -591 423 -590
rect 467 -591 468 -590
rect 1101 -591 1102 -590
rect 51 -593 52 -592
rect 170 -593 171 -592
rect 289 -593 290 -592
rect 499 -593 500 -592
rect 562 -593 563 -592
rect 870 -593 871 -592
rect 912 -593 913 -592
rect 996 -593 997 -592
rect 1038 -593 1039 -592
rect 1129 -593 1130 -592
rect 107 -595 108 -594
rect 436 -595 437 -594
rect 681 -595 682 -594
rect 940 -595 941 -594
rect 1045 -595 1046 -594
rect 1171 -595 1172 -594
rect 170 -597 171 -596
rect 198 -597 199 -596
rect 390 -597 391 -596
rect 982 -597 983 -596
rect 1052 -597 1053 -596
rect 1178 -597 1179 -596
rect 772 -599 773 -598
rect 807 -599 808 -598
rect 814 -599 815 -598
rect 912 -599 913 -598
rect 947 -599 948 -598
rect 1045 -599 1046 -598
rect 1059 -599 1060 -598
rect 1136 -599 1137 -598
rect 607 -601 608 -600
rect 807 -601 808 -600
rect 845 -601 846 -600
rect 1052 -601 1053 -600
rect 695 -603 696 -602
rect 1059 -603 1060 -602
rect 695 -605 696 -604
rect 1066 -605 1067 -604
rect 737 -607 738 -606
rect 814 -607 815 -606
rect 845 -607 846 -606
rect 1297 -607 1298 -606
rect 604 -609 605 -608
rect 737 -609 738 -608
rect 779 -609 780 -608
rect 1038 -609 1039 -608
rect 464 -611 465 -610
rect 604 -611 605 -610
rect 779 -611 780 -610
rect 852 -611 853 -610
rect 877 -611 878 -610
rect 947 -611 948 -610
rect 408 -613 409 -612
rect 464 -613 465 -612
rect 793 -613 794 -612
rect 877 -613 878 -612
rect 338 -615 339 -614
rect 408 -615 409 -614
rect 338 -617 339 -616
rect 352 -617 353 -616
rect 404 -617 405 -616
rect 793 -617 794 -616
rect 212 -619 213 -618
rect 352 -619 353 -618
rect 212 -621 213 -620
rect 541 -621 542 -620
rect 387 -623 388 -622
rect 541 -623 542 -622
rect 65 -634 66 -633
rect 264 -634 265 -633
rect 310 -634 311 -633
rect 324 -634 325 -633
rect 334 -634 335 -633
rect 422 -634 423 -633
rect 523 -634 524 -633
rect 611 -634 612 -633
rect 618 -634 619 -633
rect 681 -634 682 -633
rect 691 -634 692 -633
rect 779 -634 780 -633
rect 786 -634 787 -633
rect 1339 -634 1340 -633
rect 1419 -634 1420 -633
rect 1458 -634 1459 -633
rect 1549 -634 1550 -633
rect 1556 -634 1557 -633
rect 1619 -634 1620 -633
rect 1696 -634 1697 -633
rect 72 -636 73 -635
rect 639 -636 640 -635
rect 646 -636 647 -635
rect 1479 -636 1480 -635
rect 1528 -636 1529 -635
rect 1549 -636 1550 -635
rect 68 -638 69 -637
rect 72 -638 73 -637
rect 121 -638 122 -637
rect 635 -638 636 -637
rect 649 -638 650 -637
rect 772 -638 773 -637
rect 831 -638 832 -637
rect 1409 -638 1410 -637
rect 1444 -638 1445 -637
rect 1458 -638 1459 -637
rect 1465 -638 1466 -637
rect 1528 -638 1529 -637
rect 121 -640 122 -639
rect 212 -640 213 -639
rect 222 -640 223 -639
rect 1227 -640 1228 -639
rect 1276 -640 1277 -639
rect 1486 -640 1487 -639
rect 128 -642 129 -641
rect 233 -642 234 -641
rect 240 -642 241 -641
rect 481 -642 482 -641
rect 485 -642 486 -641
rect 772 -642 773 -641
rect 838 -642 839 -641
rect 1143 -642 1144 -641
rect 1360 -642 1361 -641
rect 1409 -642 1410 -641
rect 1437 -642 1438 -641
rect 1444 -642 1445 -641
rect 128 -644 129 -643
rect 282 -644 283 -643
rect 296 -644 297 -643
rect 422 -644 423 -643
rect 429 -644 430 -643
rect 485 -644 486 -643
rect 555 -644 556 -643
rect 607 -644 608 -643
rect 674 -644 675 -643
rect 1227 -644 1228 -643
rect 1423 -644 1424 -643
rect 1437 -644 1438 -643
rect 159 -646 160 -645
rect 975 -646 976 -645
rect 982 -646 983 -645
rect 1143 -646 1144 -645
rect 1164 -646 1165 -645
rect 1360 -646 1361 -645
rect 117 -648 118 -647
rect 982 -648 983 -647
rect 1017 -648 1018 -647
rect 1374 -648 1375 -647
rect 79 -650 80 -649
rect 1017 -650 1018 -649
rect 1052 -650 1053 -649
rect 1276 -650 1277 -649
rect 1318 -650 1319 -649
rect 1423 -650 1424 -649
rect 58 -652 59 -651
rect 79 -652 80 -651
rect 191 -652 192 -651
rect 618 -652 619 -651
rect 674 -652 675 -651
rect 1297 -652 1298 -651
rect 93 -654 94 -653
rect 191 -654 192 -653
rect 198 -654 199 -653
rect 1269 -654 1270 -653
rect 93 -656 94 -655
rect 156 -656 157 -655
rect 198 -656 199 -655
rect 359 -656 360 -655
rect 394 -656 395 -655
rect 457 -656 458 -655
rect 492 -656 493 -655
rect 975 -656 976 -655
rect 1066 -656 1067 -655
rect 1164 -656 1165 -655
rect 1192 -656 1193 -655
rect 1269 -656 1270 -655
rect 114 -658 115 -657
rect 492 -658 493 -657
rect 555 -658 556 -657
rect 856 -658 857 -657
rect 870 -658 871 -657
rect 1430 -658 1431 -657
rect 44 -660 45 -659
rect 114 -660 115 -659
rect 201 -660 202 -659
rect 1234 -660 1235 -659
rect 1255 -660 1256 -659
rect 1297 -660 1298 -659
rect 44 -662 45 -661
rect 373 -662 374 -661
rect 457 -662 458 -661
rect 842 -662 843 -661
rect 845 -662 846 -661
rect 1325 -662 1326 -661
rect 205 -664 206 -663
rect 240 -664 241 -663
rect 247 -664 248 -663
rect 324 -664 325 -663
rect 345 -664 346 -663
rect 572 -664 573 -663
rect 590 -664 591 -663
rect 695 -664 696 -663
rect 709 -664 710 -663
rect 779 -664 780 -663
rect 800 -664 801 -663
rect 1318 -664 1319 -663
rect 149 -666 150 -665
rect 247 -666 248 -665
rect 282 -666 283 -665
rect 289 -666 290 -665
rect 296 -666 297 -665
rect 331 -666 332 -665
rect 345 -666 346 -665
rect 607 -666 608 -665
rect 677 -666 678 -665
rect 1290 -666 1291 -665
rect 149 -668 150 -667
rect 751 -668 752 -667
rect 758 -668 759 -667
rect 1451 -668 1452 -667
rect 212 -670 213 -669
rect 219 -670 220 -669
rect 226 -670 227 -669
rect 478 -670 479 -669
rect 495 -670 496 -669
rect 842 -670 843 -669
rect 926 -670 927 -669
rect 1066 -670 1067 -669
rect 1108 -670 1109 -669
rect 1465 -670 1466 -669
rect 219 -672 220 -671
rect 800 -672 801 -671
rect 803 -672 804 -671
rect 1374 -672 1375 -671
rect 1395 -672 1396 -671
rect 1451 -672 1452 -671
rect 226 -674 227 -673
rect 261 -674 262 -673
rect 275 -674 276 -673
rect 289 -674 290 -673
rect 310 -674 311 -673
rect 366 -674 367 -673
rect 478 -674 479 -673
rect 534 -674 535 -673
rect 569 -674 570 -673
rect 611 -674 612 -673
rect 653 -674 654 -673
rect 758 -674 759 -673
rect 828 -674 829 -673
rect 856 -674 857 -673
rect 933 -674 934 -673
rect 1031 -674 1032 -673
rect 1038 -674 1039 -673
rect 1192 -674 1193 -673
rect 1206 -674 1207 -673
rect 1255 -674 1256 -673
rect 1283 -674 1284 -673
rect 1290 -674 1291 -673
rect 1304 -674 1305 -673
rect 1395 -674 1396 -673
rect 170 -676 171 -675
rect 366 -676 367 -675
rect 471 -676 472 -675
rect 653 -676 654 -675
rect 681 -676 682 -675
rect 737 -676 738 -675
rect 744 -676 745 -675
rect 1157 -676 1158 -675
rect 1220 -676 1221 -675
rect 1325 -676 1326 -675
rect 142 -678 143 -677
rect 471 -678 472 -677
rect 527 -678 528 -677
rect 534 -678 535 -677
rect 590 -678 591 -677
rect 625 -678 626 -677
rect 632 -678 633 -677
rect 744 -678 745 -677
rect 751 -678 752 -677
rect 905 -678 906 -677
rect 912 -678 913 -677
rect 933 -678 934 -677
rect 961 -678 962 -677
rect 1108 -678 1109 -677
rect 1122 -678 1123 -677
rect 1430 -678 1431 -677
rect 142 -680 143 -679
rect 436 -680 437 -679
rect 527 -680 528 -679
rect 940 -680 941 -679
rect 1059 -680 1060 -679
rect 1157 -680 1158 -679
rect 1248 -680 1249 -679
rect 1283 -680 1284 -679
rect 156 -682 157 -681
rect 1059 -682 1060 -681
rect 1080 -682 1081 -681
rect 1206 -682 1207 -681
rect 1262 -682 1263 -681
rect 1304 -682 1305 -681
rect 170 -684 171 -683
rect 450 -684 451 -683
rect 597 -684 598 -683
rect 625 -684 626 -683
rect 632 -684 633 -683
rect 1115 -684 1116 -683
rect 1129 -684 1130 -683
rect 1220 -684 1221 -683
rect 184 -686 185 -685
rect 569 -686 570 -685
rect 604 -686 605 -685
rect 1213 -686 1214 -685
rect 184 -688 185 -687
rect 303 -688 304 -687
rect 317 -688 318 -687
rect 387 -688 388 -687
rect 425 -688 426 -687
rect 737 -688 738 -687
rect 761 -688 762 -687
rect 1080 -688 1081 -687
rect 1087 -688 1088 -687
rect 1122 -688 1123 -687
rect 1136 -688 1137 -687
rect 1339 -688 1340 -687
rect 86 -690 87 -689
rect 387 -690 388 -689
rect 558 -690 559 -689
rect 597 -690 598 -689
rect 604 -690 605 -689
rect 1332 -690 1333 -689
rect 86 -692 87 -691
rect 107 -692 108 -691
rect 233 -692 234 -691
rect 352 -692 353 -691
rect 355 -692 356 -691
rect 394 -692 395 -691
rect 530 -692 531 -691
rect 1332 -692 1333 -691
rect 107 -694 108 -693
rect 789 -694 790 -693
rect 821 -694 822 -693
rect 1038 -694 1039 -693
rect 1094 -694 1095 -693
rect 1213 -694 1214 -693
rect 254 -696 255 -695
rect 352 -696 353 -695
rect 359 -696 360 -695
rect 464 -696 465 -695
rect 688 -696 689 -695
rect 786 -696 787 -695
rect 814 -696 815 -695
rect 821 -696 822 -695
rect 828 -696 829 -695
rect 1472 -696 1473 -695
rect 177 -698 178 -697
rect 814 -698 815 -697
rect 849 -698 850 -697
rect 940 -698 941 -697
rect 954 -698 955 -697
rect 1087 -698 1088 -697
rect 1150 -698 1151 -697
rect 1234 -698 1235 -697
rect 177 -700 178 -699
rect 327 -700 328 -699
rect 380 -700 381 -699
rect 450 -700 451 -699
rect 464 -700 465 -699
rect 1416 -700 1417 -699
rect 254 -702 255 -701
rect 373 -702 374 -701
rect 429 -702 430 -701
rect 954 -702 955 -701
rect 968 -702 969 -701
rect 1115 -702 1116 -701
rect 1178 -702 1179 -701
rect 1262 -702 1263 -701
rect 1388 -702 1389 -701
rect 1416 -702 1417 -701
rect 261 -704 262 -703
rect 338 -704 339 -703
rect 467 -704 468 -703
rect 968 -704 969 -703
rect 989 -704 990 -703
rect 1129 -704 1130 -703
rect 1178 -704 1179 -703
rect 1381 -704 1382 -703
rect 268 -706 269 -705
rect 338 -706 339 -705
rect 702 -706 703 -705
rect 709 -706 710 -705
rect 719 -706 720 -705
rect 1367 -706 1368 -705
rect 268 -708 269 -707
rect 401 -708 402 -707
rect 460 -708 461 -707
rect 702 -708 703 -707
rect 730 -708 731 -707
rect 1052 -708 1053 -707
rect 1185 -708 1186 -707
rect 1388 -708 1389 -707
rect 135 -710 136 -709
rect 401 -710 402 -709
rect 684 -710 685 -709
rect 1185 -710 1186 -709
rect 1311 -710 1312 -709
rect 1367 -710 1368 -709
rect 135 -712 136 -711
rect 205 -712 206 -711
rect 303 -712 304 -711
rect 415 -712 416 -711
rect 733 -712 734 -711
rect 1101 -712 1102 -711
rect 1346 -712 1347 -711
rect 1381 -712 1382 -711
rect 317 -714 318 -713
rect 408 -714 409 -713
rect 415 -714 416 -713
rect 499 -714 500 -713
rect 733 -714 734 -713
rect 1402 -714 1403 -713
rect 163 -716 164 -715
rect 408 -716 409 -715
rect 499 -716 500 -715
rect 576 -716 577 -715
rect 793 -716 794 -715
rect 849 -716 850 -715
rect 873 -716 874 -715
rect 1311 -716 1312 -715
rect 58 -718 59 -717
rect 163 -718 164 -717
rect 331 -718 332 -717
rect 380 -718 381 -717
rect 576 -718 577 -717
rect 716 -718 717 -717
rect 884 -718 885 -717
rect 912 -718 913 -717
rect 919 -718 920 -717
rect 961 -718 962 -717
rect 989 -718 990 -717
rect 1024 -718 1025 -717
rect 1045 -718 1046 -717
rect 1150 -718 1151 -717
rect 1171 -718 1172 -717
rect 1402 -718 1403 -717
rect 275 -720 276 -719
rect 716 -720 717 -719
rect 877 -720 878 -719
rect 1045 -720 1046 -719
rect 432 -722 433 -721
rect 884 -722 885 -721
rect 891 -722 892 -721
rect 919 -722 920 -721
rect 929 -722 930 -721
rect 1094 -722 1095 -721
rect 51 -724 52 -723
rect 891 -724 892 -723
rect 905 -724 906 -723
rect 1199 -724 1200 -723
rect 51 -726 52 -725
rect 243 -726 244 -725
rect 436 -726 437 -725
rect 1024 -726 1025 -725
rect 1073 -726 1074 -725
rect 1199 -726 1200 -725
rect 642 -728 643 -727
rect 1073 -728 1074 -727
rect 807 -730 808 -729
rect 877 -730 878 -729
rect 908 -730 909 -729
rect 1346 -730 1347 -729
rect 723 -732 724 -731
rect 807 -732 808 -731
rect 996 -732 997 -731
rect 1136 -732 1137 -731
rect 506 -734 507 -733
rect 723 -734 724 -733
rect 947 -734 948 -733
rect 996 -734 997 -733
rect 1003 -734 1004 -733
rect 1171 -734 1172 -733
rect 257 -736 258 -735
rect 506 -736 507 -735
rect 520 -736 521 -735
rect 1003 -736 1004 -735
rect 1010 -736 1011 -735
rect 1101 -736 1102 -735
rect 863 -738 864 -737
rect 947 -738 948 -737
rect 1020 -738 1021 -737
rect 1248 -738 1249 -737
rect 765 -740 766 -739
rect 863 -740 864 -739
rect 898 -740 899 -739
rect 1010 -740 1011 -739
rect 443 -742 444 -741
rect 765 -742 766 -741
rect 835 -742 836 -741
rect 898 -742 899 -741
rect 443 -744 444 -743
rect 660 -744 661 -743
rect 835 -744 836 -743
rect 1353 -744 1354 -743
rect 660 -746 661 -745
rect 667 -746 668 -745
rect 1241 -746 1242 -745
rect 1353 -746 1354 -745
rect 583 -748 584 -747
rect 667 -748 668 -747
rect 698 -748 699 -747
rect 1241 -748 1242 -747
rect 541 -750 542 -749
rect 583 -750 584 -749
rect 513 -752 514 -751
rect 541 -752 542 -751
rect 513 -754 514 -753
rect 562 -754 563 -753
rect 562 -756 563 -755
rect 796 -756 797 -755
rect 37 -767 38 -766
rect 51 -767 52 -766
rect 58 -767 59 -766
rect 562 -767 563 -766
rect 572 -767 573 -766
rect 1423 -767 1424 -766
rect 1430 -767 1431 -766
rect 1584 -767 1585 -766
rect 1696 -767 1697 -766
rect 1724 -767 1725 -766
rect 44 -769 45 -768
rect 432 -769 433 -768
rect 485 -769 486 -768
rect 530 -769 531 -768
rect 551 -769 552 -768
rect 737 -769 738 -768
rect 793 -769 794 -768
rect 1192 -769 1193 -768
rect 1255 -769 1256 -768
rect 1535 -769 1536 -768
rect 1549 -769 1550 -768
rect 1577 -769 1578 -768
rect 44 -771 45 -770
rect 61 -771 62 -770
rect 65 -771 66 -770
rect 345 -771 346 -770
rect 366 -771 367 -770
rect 646 -771 647 -770
rect 667 -771 668 -770
rect 716 -771 717 -770
rect 737 -771 738 -770
rect 947 -771 948 -770
rect 961 -771 962 -770
rect 1192 -771 1193 -770
rect 1353 -771 1354 -770
rect 1430 -771 1431 -770
rect 1437 -771 1438 -770
rect 1507 -771 1508 -770
rect 1528 -771 1529 -770
rect 1570 -771 1571 -770
rect 65 -773 66 -772
rect 72 -773 73 -772
rect 114 -773 115 -772
rect 359 -773 360 -772
rect 366 -773 367 -772
rect 513 -773 514 -772
rect 530 -773 531 -772
rect 548 -773 549 -772
rect 558 -773 559 -772
rect 1038 -773 1039 -772
rect 1115 -773 1116 -772
rect 1255 -773 1256 -772
rect 1262 -773 1263 -772
rect 1353 -773 1354 -772
rect 1409 -773 1410 -772
rect 1528 -773 1529 -772
rect 72 -775 73 -774
rect 93 -775 94 -774
rect 124 -775 125 -774
rect 289 -775 290 -774
rect 296 -775 297 -774
rect 555 -775 556 -774
rect 607 -775 608 -774
rect 772 -775 773 -774
rect 793 -775 794 -774
rect 877 -775 878 -774
rect 905 -775 906 -774
rect 1437 -775 1438 -774
rect 1444 -775 1445 -774
rect 1549 -775 1550 -774
rect 93 -777 94 -776
rect 184 -777 185 -776
rect 187 -777 188 -776
rect 310 -777 311 -776
rect 324 -777 325 -776
rect 359 -777 360 -776
rect 380 -777 381 -776
rect 555 -777 556 -776
rect 604 -777 605 -776
rect 905 -777 906 -776
rect 908 -777 909 -776
rect 1325 -777 1326 -776
rect 1367 -777 1368 -776
rect 1444 -777 1445 -776
rect 1458 -777 1459 -776
rect 1514 -777 1515 -776
rect 135 -779 136 -778
rect 331 -779 332 -778
rect 345 -779 346 -778
rect 352 -779 353 -778
rect 380 -779 381 -778
rect 457 -779 458 -778
rect 478 -779 479 -778
rect 513 -779 514 -778
rect 534 -779 535 -778
rect 604 -779 605 -778
rect 611 -779 612 -778
rect 677 -779 678 -778
rect 684 -779 685 -778
rect 922 -779 923 -778
rect 926 -779 927 -778
rect 1178 -779 1179 -778
rect 1220 -779 1221 -778
rect 1262 -779 1263 -778
rect 1290 -779 1291 -778
rect 1409 -779 1410 -778
rect 1416 -779 1417 -778
rect 1500 -779 1501 -778
rect 135 -781 136 -780
rect 156 -781 157 -780
rect 163 -781 164 -780
rect 331 -781 332 -780
rect 394 -781 395 -780
rect 478 -781 479 -780
rect 506 -781 507 -780
rect 828 -781 829 -780
rect 835 -781 836 -780
rect 856 -781 857 -780
rect 926 -781 927 -780
rect 989 -781 990 -780
rect 1017 -781 1018 -780
rect 1038 -781 1039 -780
rect 1115 -781 1116 -780
rect 1241 -781 1242 -780
rect 1346 -781 1347 -780
rect 1367 -781 1368 -780
rect 1374 -781 1375 -780
rect 1416 -781 1417 -780
rect 1472 -781 1473 -780
rect 1521 -781 1522 -780
rect 163 -783 164 -782
rect 782 -783 783 -782
rect 796 -783 797 -782
rect 1101 -783 1102 -782
rect 1178 -783 1179 -782
rect 1206 -783 1207 -782
rect 1213 -783 1214 -782
rect 1220 -783 1221 -782
rect 1227 -783 1228 -782
rect 1325 -783 1326 -782
rect 1479 -783 1480 -782
rect 1559 -783 1560 -782
rect 117 -785 118 -784
rect 1213 -785 1214 -784
rect 1241 -785 1242 -784
rect 1276 -785 1277 -784
rect 1311 -785 1312 -784
rect 1479 -785 1480 -784
rect 1486 -785 1487 -784
rect 1542 -785 1543 -784
rect 166 -787 167 -786
rect 674 -787 675 -786
rect 688 -787 689 -786
rect 1045 -787 1046 -786
rect 1059 -787 1060 -786
rect 1346 -787 1347 -786
rect 184 -789 185 -788
rect 1003 -789 1004 -788
rect 1024 -789 1025 -788
rect 1374 -789 1375 -788
rect 191 -791 192 -790
rect 464 -791 465 -790
rect 485 -791 486 -790
rect 835 -791 836 -790
rect 849 -791 850 -790
rect 856 -791 857 -790
rect 929 -791 930 -790
rect 1066 -791 1067 -790
rect 1094 -791 1095 -790
rect 1206 -791 1207 -790
rect 1248 -791 1249 -790
rect 1311 -791 1312 -790
rect 191 -793 192 -792
rect 548 -793 549 -792
rect 569 -793 570 -792
rect 1066 -793 1067 -792
rect 1080 -793 1081 -792
rect 1094 -793 1095 -792
rect 1199 -793 1200 -792
rect 1276 -793 1277 -792
rect 205 -795 206 -794
rect 765 -795 766 -794
rect 772 -795 773 -794
rect 807 -795 808 -794
rect 828 -795 829 -794
rect 1493 -795 1494 -794
rect 208 -797 209 -796
rect 1227 -797 1228 -796
rect 1248 -797 1249 -796
rect 1304 -797 1305 -796
rect 208 -799 209 -798
rect 723 -799 724 -798
rect 751 -799 752 -798
rect 1003 -799 1004 -798
rect 1027 -799 1028 -798
rect 1472 -799 1473 -798
rect 226 -801 227 -800
rect 310 -801 311 -800
rect 352 -801 353 -800
rect 506 -801 507 -800
rect 527 -801 528 -800
rect 1199 -801 1200 -800
rect 212 -803 213 -802
rect 226 -803 227 -802
rect 240 -803 241 -802
rect 289 -803 290 -802
rect 296 -803 297 -802
rect 492 -803 493 -802
rect 534 -803 535 -802
rect 758 -803 759 -802
rect 800 -803 801 -802
rect 1101 -803 1102 -802
rect 212 -805 213 -804
rect 436 -805 437 -804
rect 457 -805 458 -804
rect 527 -805 528 -804
rect 541 -805 542 -804
rect 1017 -805 1018 -804
rect 1045 -805 1046 -804
rect 1087 -805 1088 -804
rect 233 -807 234 -806
rect 436 -807 437 -806
rect 464 -807 465 -806
rect 471 -807 472 -806
rect 576 -807 577 -806
rect 765 -807 766 -806
rect 786 -807 787 -806
rect 800 -807 801 -806
rect 807 -807 808 -806
rect 863 -807 864 -806
rect 940 -807 941 -806
rect 947 -807 948 -806
rect 961 -807 962 -806
rect 1339 -807 1340 -806
rect 121 -809 122 -808
rect 786 -809 787 -808
rect 821 -809 822 -808
rect 940 -809 941 -808
rect 975 -809 976 -808
rect 1024 -809 1025 -808
rect 1059 -809 1060 -808
rect 1129 -809 1130 -808
rect 233 -811 234 -810
rect 411 -811 412 -810
rect 415 -811 416 -810
rect 523 -811 524 -810
rect 583 -811 584 -810
rect 611 -811 612 -810
rect 632 -811 633 -810
rect 667 -811 668 -810
rect 702 -811 703 -810
rect 723 -811 724 -810
rect 814 -811 815 -810
rect 821 -811 822 -810
rect 838 -811 839 -810
rect 1304 -811 1305 -810
rect 142 -813 143 -812
rect 523 -813 524 -812
rect 583 -813 584 -812
rect 681 -813 682 -812
rect 709 -813 710 -812
rect 758 -813 759 -812
rect 814 -813 815 -812
rect 1458 -813 1459 -812
rect 142 -815 143 -814
rect 891 -815 892 -814
rect 968 -815 969 -814
rect 975 -815 976 -814
rect 982 -815 983 -814
rect 989 -815 990 -814
rect 996 -815 997 -814
rect 1087 -815 1088 -814
rect 1122 -815 1123 -814
rect 1129 -815 1130 -814
rect 79 -817 80 -816
rect 891 -817 892 -816
rect 919 -817 920 -816
rect 996 -817 997 -816
rect 1073 -817 1074 -816
rect 1080 -817 1081 -816
rect 1122 -817 1123 -816
rect 1136 -817 1137 -816
rect 79 -819 80 -818
rect 86 -819 87 -818
rect 156 -819 157 -818
rect 681 -819 682 -818
rect 716 -819 717 -818
rect 964 -819 965 -818
rect 982 -819 983 -818
rect 1010 -819 1011 -818
rect 1052 -819 1053 -818
rect 1073 -819 1074 -818
rect 1136 -819 1137 -818
rect 1143 -819 1144 -818
rect 86 -821 87 -820
rect 100 -821 101 -820
rect 240 -821 241 -820
rect 387 -821 388 -820
rect 401 -821 402 -820
rect 576 -821 577 -820
rect 590 -821 591 -820
rect 849 -821 850 -820
rect 863 -821 864 -820
rect 884 -821 885 -820
rect 933 -821 934 -820
rect 1010 -821 1011 -820
rect 1031 -821 1032 -820
rect 1052 -821 1053 -820
rect 100 -823 101 -822
rect 443 -823 444 -822
rect 509 -823 510 -822
rect 1339 -823 1340 -822
rect 152 -825 153 -824
rect 443 -825 444 -824
rect 590 -825 591 -824
rect 639 -825 640 -824
rect 646 -825 647 -824
rect 1465 -825 1466 -824
rect 149 -827 150 -826
rect 639 -827 640 -826
rect 649 -827 650 -826
rect 1486 -827 1487 -826
rect 51 -829 52 -828
rect 149 -829 150 -828
rect 261 -829 262 -828
rect 324 -829 325 -828
rect 338 -829 339 -828
rect 387 -829 388 -828
rect 401 -829 402 -828
rect 422 -829 423 -828
rect 429 -829 430 -828
rect 719 -829 720 -828
rect 744 -829 745 -828
rect 884 -829 885 -828
rect 912 -829 913 -828
rect 933 -829 934 -828
rect 1381 -829 1382 -828
rect 1465 -829 1466 -828
rect 170 -831 171 -830
rect 338 -831 339 -830
rect 373 -831 374 -830
rect 492 -831 493 -830
rect 499 -831 500 -830
rect 744 -831 745 -830
rect 838 -831 839 -830
rect 1402 -831 1403 -830
rect 170 -833 171 -832
rect 198 -833 199 -832
rect 247 -833 248 -832
rect 261 -833 262 -832
rect 282 -833 283 -832
rect 394 -833 395 -832
rect 408 -833 409 -832
rect 562 -833 563 -832
rect 625 -833 626 -832
rect 968 -833 969 -832
rect 1283 -833 1284 -832
rect 1381 -833 1382 -832
rect 121 -835 122 -834
rect 282 -835 283 -834
rect 303 -835 304 -834
rect 415 -835 416 -834
rect 422 -835 423 -834
rect 873 -835 874 -834
rect 877 -835 878 -834
rect 1143 -835 1144 -834
rect 1269 -835 1270 -834
rect 1283 -835 1284 -834
rect 1360 -835 1361 -834
rect 1402 -835 1403 -834
rect 128 -837 129 -836
rect 247 -837 248 -836
rect 268 -837 269 -836
rect 303 -837 304 -836
rect 317 -837 318 -836
rect 429 -837 430 -836
rect 499 -837 500 -836
rect 1290 -837 1291 -836
rect 128 -839 129 -838
rect 177 -839 178 -838
rect 198 -839 199 -838
rect 205 -839 206 -838
rect 268 -839 269 -838
rect 831 -839 832 -838
rect 873 -839 874 -838
rect 1451 -839 1452 -838
rect 177 -841 178 -840
rect 275 -841 276 -840
rect 317 -841 318 -840
rect 450 -841 451 -840
rect 635 -841 636 -840
rect 709 -841 710 -840
rect 831 -841 832 -840
rect 1395 -841 1396 -840
rect 107 -843 108 -842
rect 450 -843 451 -842
rect 649 -843 650 -842
rect 702 -843 703 -842
rect 880 -843 881 -842
rect 1395 -843 1396 -842
rect 107 -845 108 -844
rect 1423 -845 1424 -844
rect 254 -847 255 -846
rect 275 -847 276 -846
rect 373 -847 374 -846
rect 730 -847 731 -846
rect 898 -847 899 -846
rect 912 -847 913 -846
rect 919 -847 920 -846
rect 1031 -847 1032 -846
rect 1164 -847 1165 -846
rect 1360 -847 1361 -846
rect 1388 -847 1389 -846
rect 1451 -847 1452 -846
rect 159 -849 160 -848
rect 898 -849 899 -848
rect 1185 -849 1186 -848
rect 1388 -849 1389 -848
rect 520 -851 521 -850
rect 1185 -851 1186 -850
rect 1234 -851 1235 -850
rect 1269 -851 1270 -850
rect 520 -853 521 -852
rect 541 -853 542 -852
rect 653 -853 654 -852
rect 730 -853 731 -852
rect 870 -853 871 -852
rect 1164 -853 1165 -852
rect 1234 -853 1235 -852
rect 1318 -853 1319 -852
rect 653 -855 654 -854
rect 674 -855 675 -854
rect 691 -855 692 -854
rect 1318 -855 1319 -854
rect 660 -857 661 -856
rect 688 -857 689 -856
rect 751 -857 752 -856
rect 870 -857 871 -856
rect 660 -859 661 -858
rect 695 -859 696 -858
rect 618 -861 619 -860
rect 695 -861 696 -860
rect 597 -863 598 -862
rect 618 -863 619 -862
rect 597 -865 598 -864
rect 842 -865 843 -864
rect 779 -867 780 -866
rect 842 -867 843 -866
rect 471 -869 472 -868
rect 779 -869 780 -868
rect 30 -880 31 -879
rect 142 -880 143 -879
rect 149 -880 150 -879
rect 891 -880 892 -879
rect 919 -880 920 -879
rect 1451 -880 1452 -879
rect 1542 -880 1543 -879
rect 1566 -880 1567 -879
rect 1570 -880 1571 -879
rect 1626 -880 1627 -879
rect 1724 -880 1725 -879
rect 1738 -880 1739 -879
rect 44 -882 45 -881
rect 628 -882 629 -881
rect 656 -882 657 -881
rect 1570 -882 1571 -881
rect 1577 -882 1578 -881
rect 1612 -882 1613 -881
rect 44 -884 45 -883
rect 51 -884 52 -883
rect 79 -884 80 -883
rect 649 -884 650 -883
rect 660 -884 661 -883
rect 831 -884 832 -883
rect 838 -884 839 -883
rect 870 -884 871 -883
rect 873 -884 874 -883
rect 1255 -884 1256 -883
rect 1318 -884 1319 -883
rect 1633 -884 1634 -883
rect 51 -886 52 -885
rect 65 -886 66 -885
rect 79 -886 80 -885
rect 128 -886 129 -885
rect 135 -886 136 -885
rect 142 -886 143 -885
rect 166 -886 167 -885
rect 1360 -886 1361 -885
rect 1521 -886 1522 -885
rect 1542 -886 1543 -885
rect 1573 -886 1574 -885
rect 1577 -886 1578 -885
rect 1584 -886 1585 -885
rect 1619 -886 1620 -885
rect 65 -888 66 -887
rect 72 -888 73 -887
rect 82 -888 83 -887
rect 233 -888 234 -887
rect 257 -888 258 -887
rect 1437 -888 1438 -887
rect 1479 -888 1480 -887
rect 1584 -888 1585 -887
rect 72 -890 73 -889
rect 86 -890 87 -889
rect 93 -890 94 -889
rect 152 -890 153 -889
rect 208 -890 209 -889
rect 352 -890 353 -889
rect 408 -890 409 -889
rect 551 -890 552 -889
rect 660 -890 661 -889
rect 856 -890 857 -889
rect 880 -890 881 -889
rect 1528 -890 1529 -889
rect 58 -892 59 -891
rect 86 -892 87 -891
rect 93 -892 94 -891
rect 569 -892 570 -891
rect 667 -892 668 -891
rect 940 -892 941 -891
rect 964 -892 965 -891
rect 1416 -892 1417 -891
rect 1437 -892 1438 -891
rect 1444 -892 1445 -891
rect 1479 -892 1480 -891
rect 1486 -892 1487 -891
rect 1493 -892 1494 -891
rect 1521 -892 1522 -891
rect 58 -894 59 -893
rect 422 -894 423 -893
rect 436 -894 437 -893
rect 642 -894 643 -893
rect 667 -894 668 -893
rect 688 -894 689 -893
rect 775 -894 776 -893
rect 1206 -894 1207 -893
rect 1346 -894 1347 -893
rect 1556 -894 1557 -893
rect 100 -896 101 -895
rect 964 -896 965 -895
rect 985 -896 986 -895
rect 1381 -896 1382 -895
rect 1388 -896 1389 -895
rect 1444 -896 1445 -895
rect 1465 -896 1466 -895
rect 1493 -896 1494 -895
rect 1514 -896 1515 -895
rect 1528 -896 1529 -895
rect 100 -898 101 -897
rect 877 -898 878 -897
rect 891 -898 892 -897
rect 954 -898 955 -897
rect 961 -898 962 -897
rect 1556 -898 1557 -897
rect 107 -900 108 -899
rect 296 -900 297 -899
rect 317 -900 318 -899
rect 320 -900 321 -899
rect 338 -900 339 -899
rect 499 -900 500 -899
rect 502 -900 503 -899
rect 968 -900 969 -899
rect 992 -900 993 -899
rect 1451 -900 1452 -899
rect 1465 -900 1466 -899
rect 1507 -900 1508 -899
rect 107 -902 108 -901
rect 212 -902 213 -901
rect 219 -902 220 -901
rect 534 -902 535 -901
rect 548 -902 549 -901
rect 590 -902 591 -901
rect 674 -902 675 -901
rect 884 -902 885 -901
rect 905 -902 906 -901
rect 919 -902 920 -901
rect 926 -902 927 -901
rect 929 -902 930 -901
rect 940 -902 941 -901
rect 1010 -902 1011 -901
rect 1069 -902 1070 -901
rect 1549 -902 1550 -901
rect 110 -904 111 -903
rect 310 -904 311 -903
rect 317 -904 318 -903
rect 324 -904 325 -903
rect 352 -904 353 -903
rect 450 -904 451 -903
rect 502 -904 503 -903
rect 1423 -904 1424 -903
rect 1472 -904 1473 -903
rect 1514 -904 1515 -903
rect 1549 -904 1550 -903
rect 1563 -904 1564 -903
rect 121 -906 122 -905
rect 366 -906 367 -905
rect 408 -906 409 -905
rect 723 -906 724 -905
rect 779 -906 780 -905
rect 842 -906 843 -905
rect 856 -906 857 -905
rect 975 -906 976 -905
rect 1111 -906 1112 -905
rect 1486 -906 1487 -905
rect 1563 -906 1564 -905
rect 1605 -906 1606 -905
rect 121 -908 122 -907
rect 124 -908 125 -907
rect 128 -908 129 -907
rect 275 -908 276 -907
rect 289 -908 290 -907
rect 296 -908 297 -907
rect 310 -908 311 -907
rect 394 -908 395 -907
rect 411 -908 412 -907
rect 922 -908 923 -907
rect 926 -908 927 -907
rect 933 -908 934 -907
rect 968 -908 969 -907
rect 989 -908 990 -907
rect 1171 -908 1172 -907
rect 1206 -908 1207 -907
rect 1248 -908 1249 -907
rect 1381 -908 1382 -907
rect 1409 -908 1410 -907
rect 1416 -908 1417 -907
rect 138 -910 139 -909
rect 380 -910 381 -909
rect 394 -910 395 -909
rect 702 -910 703 -909
rect 723 -910 724 -909
rect 758 -910 759 -909
rect 782 -910 783 -909
rect 1395 -910 1396 -909
rect 163 -912 164 -911
rect 212 -912 213 -911
rect 222 -912 223 -911
rect 254 -912 255 -911
rect 268 -912 269 -911
rect 436 -912 437 -911
rect 446 -912 447 -911
rect 870 -912 871 -911
rect 877 -912 878 -911
rect 1192 -912 1193 -911
rect 1248 -912 1249 -911
rect 1262 -912 1263 -911
rect 1290 -912 1291 -911
rect 1346 -912 1347 -911
rect 1367 -912 1368 -911
rect 1409 -912 1410 -911
rect 163 -914 164 -913
rect 177 -914 178 -913
rect 191 -914 192 -913
rect 289 -914 290 -913
rect 380 -914 381 -913
rect 772 -914 773 -913
rect 828 -914 829 -913
rect 1360 -914 1361 -913
rect 1374 -914 1375 -913
rect 1507 -914 1508 -913
rect 177 -916 178 -915
rect 387 -916 388 -915
rect 450 -916 451 -915
rect 492 -916 493 -915
rect 506 -916 507 -915
rect 1017 -916 1018 -915
rect 1164 -916 1165 -915
rect 1192 -916 1193 -915
rect 1241 -916 1242 -915
rect 1262 -916 1263 -915
rect 1269 -916 1270 -915
rect 1290 -916 1291 -915
rect 1297 -916 1298 -915
rect 1367 -916 1368 -915
rect 1395 -916 1396 -915
rect 1430 -916 1431 -915
rect 191 -918 192 -917
rect 513 -918 514 -917
rect 520 -918 521 -917
rect 1318 -918 1319 -917
rect 135 -920 136 -919
rect 513 -920 514 -919
rect 523 -920 524 -919
rect 695 -920 696 -919
rect 698 -920 699 -919
rect 954 -920 955 -919
rect 975 -920 976 -919
rect 1255 -920 1256 -919
rect 1304 -920 1305 -919
rect 1388 -920 1389 -919
rect 198 -922 199 -921
rect 422 -922 423 -921
rect 425 -922 426 -921
rect 520 -922 521 -921
rect 530 -922 531 -921
rect 1024 -922 1025 -921
rect 1115 -922 1116 -921
rect 1297 -922 1298 -921
rect 198 -924 199 -923
rect 261 -924 262 -923
rect 268 -924 269 -923
rect 303 -924 304 -923
rect 387 -924 388 -923
rect 632 -924 633 -923
rect 670 -924 671 -923
rect 828 -924 829 -923
rect 845 -924 846 -923
rect 1374 -924 1375 -923
rect 205 -926 206 -925
rect 338 -926 339 -925
rect 492 -926 493 -925
rect 684 -926 685 -925
rect 688 -926 689 -925
rect 1311 -926 1312 -925
rect 205 -928 206 -927
rect 373 -928 374 -927
rect 509 -928 510 -927
rect 516 -928 517 -927
rect 534 -928 535 -927
rect 555 -928 556 -927
rect 569 -928 570 -927
rect 618 -928 619 -927
rect 625 -928 626 -927
rect 1423 -928 1424 -927
rect 184 -930 185 -929
rect 555 -930 556 -929
rect 586 -930 587 -929
rect 1115 -930 1116 -929
rect 1157 -930 1158 -929
rect 1164 -930 1165 -929
rect 1171 -930 1172 -929
rect 1178 -930 1179 -929
rect 1227 -930 1228 -929
rect 1269 -930 1270 -929
rect 1283 -930 1284 -929
rect 1304 -930 1305 -929
rect 149 -932 150 -931
rect 184 -932 185 -931
rect 226 -932 227 -931
rect 366 -932 367 -931
rect 373 -932 374 -931
rect 401 -932 402 -931
rect 506 -932 507 -931
rect 1283 -932 1284 -931
rect 233 -934 234 -933
rect 478 -934 479 -933
rect 509 -934 510 -933
rect 527 -934 528 -933
rect 590 -934 591 -933
rect 821 -934 822 -933
rect 898 -934 899 -933
rect 905 -934 906 -933
rect 933 -934 934 -933
rect 947 -934 948 -933
rect 999 -934 1000 -933
rect 1157 -934 1158 -933
rect 1234 -934 1235 -933
rect 1241 -934 1242 -933
rect 250 -936 251 -935
rect 548 -936 549 -935
rect 611 -936 612 -935
rect 632 -936 633 -935
rect 674 -936 675 -935
rect 730 -936 731 -935
rect 758 -936 759 -935
rect 786 -936 787 -935
rect 898 -936 899 -935
rect 1353 -936 1354 -935
rect 254 -938 255 -937
rect 282 -938 283 -937
rect 303 -938 304 -937
rect 415 -938 416 -937
rect 478 -938 479 -937
rect 485 -938 486 -937
rect 527 -938 528 -937
rect 814 -938 815 -937
rect 835 -938 836 -937
rect 1353 -938 1354 -937
rect 170 -940 171 -939
rect 282 -940 283 -939
rect 401 -940 402 -939
rect 429 -940 430 -939
rect 485 -940 486 -939
rect 653 -940 654 -939
rect 677 -940 678 -939
rect 1325 -940 1326 -939
rect 156 -942 157 -941
rect 170 -942 171 -941
rect 261 -942 262 -941
rect 345 -942 346 -941
rect 415 -942 416 -941
rect 541 -942 542 -941
rect 604 -942 605 -941
rect 611 -942 612 -941
rect 625 -942 626 -941
rect 649 -942 650 -941
rect 684 -942 685 -941
rect 786 -942 787 -941
rect 800 -942 801 -941
rect 814 -942 815 -941
rect 901 -942 902 -941
rect 1311 -942 1312 -941
rect 1325 -942 1326 -941
rect 1339 -942 1340 -941
rect 156 -944 157 -943
rect 247 -944 248 -943
rect 275 -944 276 -943
rect 471 -944 472 -943
rect 541 -944 542 -943
rect 562 -944 563 -943
rect 695 -944 696 -943
rect 744 -944 745 -943
rect 768 -944 769 -943
rect 1339 -944 1340 -943
rect 345 -946 346 -945
rect 359 -946 360 -945
rect 429 -946 430 -945
rect 576 -946 577 -945
rect 597 -946 598 -945
rect 744 -946 745 -945
rect 772 -946 773 -945
rect 1591 -946 1592 -945
rect 114 -948 115 -947
rect 359 -948 360 -947
rect 457 -948 458 -947
rect 604 -948 605 -947
rect 702 -948 703 -947
rect 751 -948 752 -947
rect 793 -948 794 -947
rect 800 -948 801 -947
rect 1017 -948 1018 -947
rect 1038 -948 1039 -947
rect 1150 -948 1151 -947
rect 1178 -948 1179 -947
rect 1220 -948 1221 -947
rect 1234 -948 1235 -947
rect 114 -950 115 -949
rect 240 -950 241 -949
rect 443 -950 444 -949
rect 457 -950 458 -949
rect 464 -950 465 -949
rect 471 -950 472 -949
rect 562 -950 563 -949
rect 765 -950 766 -949
rect 793 -950 794 -949
rect 807 -950 808 -949
rect 1024 -950 1025 -949
rect 1052 -950 1053 -949
rect 1108 -950 1109 -949
rect 1220 -950 1221 -949
rect 37 -952 38 -951
rect 240 -952 241 -951
rect 443 -952 444 -951
rect 1472 -952 1473 -951
rect 37 -954 38 -953
rect 863 -954 864 -953
rect 929 -954 930 -953
rect 947 -954 948 -953
rect 1038 -954 1039 -953
rect 1094 -954 1095 -953
rect 1150 -954 1151 -953
rect 1332 -954 1333 -953
rect 464 -956 465 -955
rect 1010 -956 1011 -955
rect 1052 -956 1053 -955
rect 1101 -956 1102 -955
rect 1332 -956 1333 -955
rect 1402 -956 1403 -955
rect 576 -958 577 -957
rect 737 -958 738 -957
rect 765 -958 766 -957
rect 1598 -958 1599 -957
rect 583 -960 584 -959
rect 751 -960 752 -959
rect 842 -960 843 -959
rect 1402 -960 1403 -959
rect 583 -962 584 -961
rect 849 -962 850 -961
rect 1059 -962 1060 -961
rect 1101 -962 1102 -961
rect 597 -964 598 -963
rect 1003 -964 1004 -963
rect 1031 -964 1032 -963
rect 1059 -964 1060 -963
rect 1094 -964 1095 -963
rect 1185 -964 1186 -963
rect 639 -966 640 -965
rect 1185 -966 1186 -965
rect 639 -968 640 -967
rect 1430 -968 1431 -967
rect 646 -970 647 -969
rect 863 -970 864 -969
rect 982 -970 983 -969
rect 1003 -970 1004 -969
rect 1031 -970 1032 -969
rect 1073 -970 1074 -969
rect 646 -972 647 -971
rect 1276 -972 1277 -971
rect 716 -974 717 -973
rect 821 -974 822 -973
rect 849 -974 850 -973
rect 912 -974 913 -973
rect 978 -974 979 -973
rect 1276 -974 1277 -973
rect 681 -976 682 -975
rect 912 -976 913 -975
rect 982 -976 983 -975
rect 1213 -976 1214 -975
rect 226 -978 227 -977
rect 681 -978 682 -977
rect 709 -978 710 -977
rect 716 -978 717 -977
rect 730 -978 731 -977
rect 1227 -978 1228 -977
rect 499 -980 500 -979
rect 709 -980 710 -979
rect 733 -980 734 -979
rect 835 -980 836 -979
rect 1073 -980 1074 -979
rect 1080 -980 1081 -979
rect 1199 -980 1200 -979
rect 1213 -980 1214 -979
rect 737 -982 738 -981
rect 996 -982 997 -981
rect 1045 -982 1046 -981
rect 1199 -982 1200 -981
rect 996 -984 997 -983
rect 1535 -984 1536 -983
rect 653 -986 654 -985
rect 1535 -986 1536 -985
rect 1045 -988 1046 -987
rect 1143 -988 1144 -987
rect 1080 -990 1081 -989
rect 1087 -990 1088 -989
rect 1136 -990 1137 -989
rect 1143 -990 1144 -989
rect 884 -992 885 -991
rect 1087 -992 1088 -991
rect 1122 -992 1123 -991
rect 1136 -992 1137 -991
rect 1066 -994 1067 -993
rect 1122 -994 1123 -993
rect 537 -996 538 -995
rect 1066 -996 1067 -995
rect 23 -1007 24 -1006
rect 618 -1007 619 -1006
rect 628 -1007 629 -1006
rect 723 -1007 724 -1006
rect 768 -1007 769 -1006
rect 940 -1007 941 -1006
rect 961 -1007 962 -1006
rect 1332 -1007 1333 -1006
rect 1374 -1007 1375 -1006
rect 1566 -1007 1567 -1006
rect 1570 -1007 1571 -1006
rect 1675 -1007 1676 -1006
rect 1738 -1007 1739 -1006
rect 1745 -1007 1746 -1006
rect 30 -1009 31 -1008
rect 135 -1009 136 -1008
rect 149 -1009 150 -1008
rect 205 -1009 206 -1008
rect 250 -1009 251 -1008
rect 296 -1009 297 -1008
rect 310 -1009 311 -1008
rect 516 -1009 517 -1008
rect 555 -1009 556 -1008
rect 723 -1009 724 -1008
rect 786 -1009 787 -1008
rect 901 -1009 902 -1008
rect 919 -1009 920 -1008
rect 1384 -1009 1385 -1008
rect 1528 -1009 1529 -1008
rect 1570 -1009 1571 -1008
rect 1591 -1009 1592 -1008
rect 1682 -1009 1683 -1008
rect 30 -1011 31 -1010
rect 597 -1011 598 -1010
rect 611 -1011 612 -1010
rect 656 -1011 657 -1010
rect 667 -1011 668 -1010
rect 730 -1011 731 -1010
rect 786 -1011 787 -1010
rect 800 -1011 801 -1010
rect 845 -1011 846 -1010
rect 1199 -1011 1200 -1010
rect 1241 -1011 1242 -1010
rect 1374 -1011 1375 -1010
rect 1486 -1011 1487 -1010
rect 1528 -1011 1529 -1010
rect 1535 -1011 1536 -1010
rect 1640 -1011 1641 -1010
rect 37 -1013 38 -1012
rect 695 -1013 696 -1012
rect 698 -1013 699 -1012
rect 1591 -1013 1592 -1012
rect 1626 -1013 1627 -1012
rect 1654 -1013 1655 -1012
rect 44 -1015 45 -1014
rect 75 -1015 76 -1014
rect 82 -1015 83 -1014
rect 107 -1015 108 -1014
rect 114 -1015 115 -1014
rect 215 -1015 216 -1014
rect 275 -1015 276 -1014
rect 999 -1015 1000 -1014
rect 1010 -1015 1011 -1014
rect 1521 -1015 1522 -1014
rect 1552 -1015 1553 -1014
rect 1612 -1015 1613 -1014
rect 44 -1017 45 -1016
rect 86 -1017 87 -1016
rect 89 -1017 90 -1016
rect 408 -1017 409 -1016
rect 422 -1017 423 -1016
rect 1605 -1017 1606 -1016
rect 58 -1019 59 -1018
rect 61 -1019 62 -1018
rect 72 -1019 73 -1018
rect 86 -1019 87 -1018
rect 100 -1019 101 -1018
rect 425 -1019 426 -1018
rect 485 -1019 486 -1018
rect 611 -1019 612 -1018
rect 618 -1019 619 -1018
rect 632 -1019 633 -1018
rect 684 -1019 685 -1018
rect 1220 -1019 1221 -1018
rect 1241 -1019 1242 -1018
rect 1297 -1019 1298 -1018
rect 1360 -1019 1361 -1018
rect 1486 -1019 1487 -1018
rect 1500 -1019 1501 -1018
rect 1535 -1019 1536 -1018
rect 1556 -1019 1557 -1018
rect 1612 -1019 1613 -1018
rect 51 -1021 52 -1020
rect 72 -1021 73 -1020
rect 100 -1021 101 -1020
rect 436 -1021 437 -1020
rect 492 -1021 493 -1020
rect 775 -1021 776 -1020
rect 800 -1021 801 -1020
rect 1248 -1021 1249 -1020
rect 1297 -1021 1298 -1020
rect 1311 -1021 1312 -1020
rect 1395 -1021 1396 -1020
rect 1500 -1021 1501 -1020
rect 1563 -1021 1564 -1020
rect 1647 -1021 1648 -1020
rect 51 -1023 52 -1022
rect 121 -1023 122 -1022
rect 128 -1023 129 -1022
rect 236 -1023 237 -1022
rect 268 -1023 269 -1022
rect 408 -1023 409 -1022
rect 492 -1023 493 -1022
rect 992 -1023 993 -1022
rect 996 -1023 997 -1022
rect 1325 -1023 1326 -1022
rect 1381 -1023 1382 -1022
rect 1395 -1023 1396 -1022
rect 1423 -1023 1424 -1022
rect 1521 -1023 1522 -1022
rect 1577 -1023 1578 -1022
rect 1626 -1023 1627 -1022
rect 58 -1025 59 -1024
rect 65 -1025 66 -1024
rect 107 -1025 108 -1024
rect 481 -1025 482 -1024
rect 499 -1025 500 -1024
rect 604 -1025 605 -1024
rect 632 -1025 633 -1024
rect 702 -1025 703 -1024
rect 730 -1025 731 -1024
rect 758 -1025 759 -1024
rect 835 -1025 836 -1024
rect 996 -1025 997 -1024
rect 1003 -1025 1004 -1024
rect 1010 -1025 1011 -1024
rect 1013 -1025 1014 -1024
rect 1031 -1025 1032 -1024
rect 1108 -1025 1109 -1024
rect 1556 -1025 1557 -1024
rect 1584 -1025 1585 -1024
rect 1605 -1025 1606 -1024
rect 114 -1027 115 -1026
rect 212 -1027 213 -1026
rect 275 -1027 276 -1026
rect 842 -1027 843 -1026
rect 856 -1027 857 -1026
rect 919 -1027 920 -1026
rect 933 -1027 934 -1026
rect 961 -1027 962 -1026
rect 975 -1027 976 -1026
rect 1066 -1027 1067 -1026
rect 1111 -1027 1112 -1026
rect 1493 -1027 1494 -1026
rect 1507 -1027 1508 -1026
rect 1584 -1027 1585 -1026
rect 121 -1029 122 -1028
rect 317 -1029 318 -1028
rect 324 -1029 325 -1028
rect 509 -1029 510 -1028
rect 520 -1029 521 -1028
rect 702 -1029 703 -1028
rect 733 -1029 734 -1028
rect 1360 -1029 1361 -1028
rect 1409 -1029 1410 -1028
rect 1423 -1029 1424 -1028
rect 1430 -1029 1431 -1028
rect 1507 -1029 1508 -1028
rect 1542 -1029 1543 -1028
rect 1577 -1029 1578 -1028
rect 128 -1031 129 -1030
rect 233 -1031 234 -1030
rect 282 -1031 283 -1030
rect 443 -1031 444 -1030
rect 541 -1031 542 -1030
rect 667 -1031 668 -1030
rect 688 -1031 689 -1030
rect 1185 -1031 1186 -1030
rect 1220 -1031 1221 -1030
rect 1255 -1031 1256 -1030
rect 1318 -1031 1319 -1030
rect 1325 -1031 1326 -1030
rect 1409 -1031 1410 -1030
rect 1437 -1031 1438 -1030
rect 1444 -1031 1445 -1030
rect 1563 -1031 1564 -1030
rect 138 -1033 139 -1032
rect 485 -1033 486 -1032
rect 506 -1033 507 -1032
rect 1318 -1033 1319 -1032
rect 1416 -1033 1417 -1032
rect 1437 -1033 1438 -1032
rect 1444 -1033 1445 -1032
rect 1451 -1033 1452 -1032
rect 138 -1035 139 -1034
rect 1472 -1035 1473 -1034
rect 156 -1037 157 -1036
rect 317 -1037 318 -1036
rect 331 -1037 332 -1036
rect 502 -1037 503 -1036
rect 541 -1037 542 -1036
rect 569 -1037 570 -1036
rect 576 -1037 577 -1036
rect 695 -1037 696 -1036
rect 737 -1037 738 -1036
rect 842 -1037 843 -1036
rect 863 -1037 864 -1036
rect 887 -1037 888 -1036
rect 891 -1037 892 -1036
rect 940 -1037 941 -1036
rect 954 -1037 955 -1036
rect 1031 -1037 1032 -1036
rect 1066 -1037 1067 -1036
rect 1101 -1037 1102 -1036
rect 1115 -1037 1116 -1036
rect 1332 -1037 1333 -1036
rect 1402 -1037 1403 -1036
rect 1416 -1037 1417 -1036
rect 1472 -1037 1473 -1036
rect 1619 -1037 1620 -1036
rect 156 -1039 157 -1038
rect 387 -1039 388 -1038
rect 394 -1039 395 -1038
rect 520 -1039 521 -1038
rect 548 -1039 549 -1038
rect 555 -1039 556 -1038
rect 562 -1039 563 -1038
rect 604 -1039 605 -1038
rect 660 -1039 661 -1038
rect 758 -1039 759 -1038
rect 793 -1039 794 -1038
rect 835 -1039 836 -1038
rect 866 -1039 867 -1038
rect 1150 -1039 1151 -1038
rect 1157 -1039 1158 -1038
rect 1311 -1039 1312 -1038
rect 1388 -1039 1389 -1038
rect 1402 -1039 1403 -1038
rect 1598 -1039 1599 -1038
rect 1619 -1039 1620 -1038
rect 170 -1041 171 -1040
rect 173 -1041 174 -1040
rect 177 -1041 178 -1040
rect 268 -1041 269 -1040
rect 296 -1041 297 -1040
rect 880 -1041 881 -1040
rect 891 -1041 892 -1040
rect 1115 -1041 1116 -1040
rect 1129 -1041 1130 -1040
rect 1132 -1041 1133 -1040
rect 1157 -1041 1158 -1040
rect 1381 -1041 1382 -1040
rect 1388 -1041 1389 -1040
rect 1475 -1041 1476 -1040
rect 170 -1043 171 -1042
rect 240 -1043 241 -1042
rect 310 -1043 311 -1042
rect 397 -1043 398 -1042
rect 401 -1043 402 -1042
rect 436 -1043 437 -1042
rect 457 -1043 458 -1042
rect 506 -1043 507 -1042
rect 548 -1043 549 -1042
rect 677 -1043 678 -1042
rect 691 -1043 692 -1042
rect 772 -1043 773 -1042
rect 894 -1043 895 -1042
rect 1080 -1043 1081 -1042
rect 1090 -1043 1091 -1042
rect 1430 -1043 1431 -1042
rect 177 -1045 178 -1044
rect 212 -1045 213 -1044
rect 219 -1045 220 -1044
rect 282 -1045 283 -1044
rect 331 -1045 332 -1044
rect 450 -1045 451 -1044
rect 457 -1045 458 -1044
rect 471 -1045 472 -1044
rect 562 -1045 563 -1044
rect 1493 -1045 1494 -1044
rect 184 -1047 185 -1046
rect 205 -1047 206 -1046
rect 219 -1047 220 -1046
rect 534 -1047 535 -1046
rect 569 -1047 570 -1046
rect 674 -1047 675 -1046
rect 716 -1047 717 -1046
rect 737 -1047 738 -1046
rect 870 -1047 871 -1046
rect 1080 -1047 1081 -1046
rect 1129 -1047 1130 -1046
rect 1164 -1047 1165 -1046
rect 1185 -1047 1186 -1046
rect 1206 -1047 1207 -1046
rect 1234 -1047 1235 -1046
rect 1248 -1047 1249 -1046
rect 1255 -1047 1256 -1046
rect 1304 -1047 1305 -1046
rect 142 -1049 143 -1048
rect 184 -1049 185 -1048
rect 191 -1049 192 -1048
rect 646 -1049 647 -1048
rect 660 -1049 661 -1048
rect 803 -1049 804 -1048
rect 821 -1049 822 -1048
rect 870 -1049 871 -1048
rect 877 -1049 878 -1048
rect 1304 -1049 1305 -1048
rect 142 -1051 143 -1050
rect 646 -1051 647 -1050
rect 733 -1051 734 -1050
rect 1598 -1051 1599 -1050
rect 191 -1053 192 -1052
rect 254 -1053 255 -1052
rect 338 -1053 339 -1052
rect 387 -1053 388 -1052
rect 394 -1053 395 -1052
rect 1353 -1053 1354 -1052
rect 198 -1055 199 -1054
rect 324 -1055 325 -1054
rect 352 -1055 353 -1054
rect 621 -1055 622 -1054
rect 625 -1055 626 -1054
rect 716 -1055 717 -1054
rect 744 -1055 745 -1054
rect 821 -1055 822 -1054
rect 877 -1055 878 -1054
rect 1199 -1055 1200 -1054
rect 1206 -1055 1207 -1054
rect 1549 -1055 1550 -1054
rect 163 -1057 164 -1056
rect 198 -1057 199 -1056
rect 254 -1057 255 -1056
rect 415 -1057 416 -1056
rect 446 -1057 447 -1056
rect 625 -1057 626 -1056
rect 744 -1057 745 -1056
rect 779 -1057 780 -1056
rect 912 -1057 913 -1056
rect 1542 -1057 1543 -1056
rect 163 -1059 164 -1058
rect 380 -1059 381 -1058
rect 401 -1059 402 -1058
rect 590 -1059 591 -1058
rect 597 -1059 598 -1058
rect 1055 -1059 1056 -1058
rect 1073 -1059 1074 -1058
rect 1101 -1059 1102 -1058
rect 1227 -1059 1228 -1058
rect 1234 -1059 1235 -1058
rect 1353 -1059 1354 -1058
rect 1367 -1059 1368 -1058
rect 1465 -1059 1466 -1058
rect 1549 -1059 1550 -1058
rect 261 -1061 262 -1060
rect 352 -1061 353 -1060
rect 359 -1061 360 -1060
rect 415 -1061 416 -1060
rect 450 -1061 451 -1060
rect 649 -1061 650 -1060
rect 653 -1061 654 -1060
rect 779 -1061 780 -1060
rect 926 -1061 927 -1060
rect 954 -1061 955 -1060
rect 982 -1061 983 -1060
rect 1108 -1061 1109 -1060
rect 1213 -1061 1214 -1060
rect 1227 -1061 1228 -1060
rect 1346 -1061 1347 -1060
rect 1367 -1061 1368 -1060
rect 1465 -1061 1466 -1060
rect 1479 -1061 1480 -1060
rect 359 -1063 360 -1062
rect 887 -1063 888 -1062
rect 905 -1063 906 -1062
rect 982 -1063 983 -1062
rect 985 -1063 986 -1062
rect 1514 -1063 1515 -1062
rect 373 -1065 374 -1064
rect 443 -1065 444 -1064
rect 464 -1065 465 -1064
rect 590 -1065 591 -1064
rect 649 -1065 650 -1064
rect 926 -1065 927 -1064
rect 933 -1065 934 -1064
rect 1017 -1065 1018 -1064
rect 1024 -1065 1025 -1064
rect 1027 -1065 1028 -1064
rect 1073 -1065 1074 -1064
rect 1136 -1065 1137 -1064
rect 1171 -1065 1172 -1064
rect 1213 -1065 1214 -1064
rect 1458 -1065 1459 -1064
rect 1514 -1065 1515 -1064
rect 226 -1067 227 -1066
rect 373 -1067 374 -1066
rect 380 -1067 381 -1066
rect 429 -1067 430 -1066
rect 471 -1067 472 -1066
rect 912 -1067 913 -1066
rect 968 -1067 969 -1066
rect 1017 -1067 1018 -1066
rect 1024 -1067 1025 -1066
rect 1038 -1067 1039 -1066
rect 1136 -1067 1137 -1066
rect 1178 -1067 1179 -1066
rect 226 -1069 227 -1068
rect 303 -1069 304 -1068
rect 429 -1069 430 -1068
rect 478 -1069 479 -1068
rect 534 -1069 535 -1068
rect 698 -1069 699 -1068
rect 863 -1069 864 -1068
rect 1479 -1069 1480 -1068
rect 289 -1071 290 -1070
rect 464 -1071 465 -1070
rect 576 -1071 577 -1070
rect 1451 -1071 1452 -1070
rect 289 -1073 290 -1072
rect 527 -1073 528 -1072
rect 583 -1073 584 -1072
rect 856 -1073 857 -1072
rect 905 -1073 906 -1072
rect 1003 -1073 1004 -1072
rect 1122 -1073 1123 -1072
rect 1178 -1073 1179 -1072
rect 250 -1075 251 -1074
rect 527 -1075 528 -1074
rect 586 -1075 587 -1074
rect 793 -1075 794 -1074
rect 947 -1075 948 -1074
rect 968 -1075 969 -1074
rect 989 -1075 990 -1074
rect 1262 -1075 1263 -1074
rect 303 -1077 304 -1076
rect 765 -1077 766 -1076
rect 947 -1077 948 -1076
rect 1052 -1077 1053 -1076
rect 1132 -1077 1133 -1076
rect 1164 -1077 1165 -1076
rect 1171 -1077 1172 -1076
rect 1192 -1077 1193 -1076
rect 1262 -1077 1263 -1076
rect 1290 -1077 1291 -1076
rect 131 -1079 132 -1078
rect 765 -1079 766 -1078
rect 1045 -1079 1046 -1078
rect 1122 -1079 1123 -1078
rect 1143 -1079 1144 -1078
rect 1192 -1079 1193 -1078
rect 1283 -1079 1284 -1078
rect 1290 -1079 1291 -1078
rect 338 -1081 339 -1080
rect 989 -1081 990 -1080
rect 1045 -1081 1046 -1080
rect 1059 -1081 1060 -1080
rect 1094 -1081 1095 -1080
rect 1143 -1081 1144 -1080
rect 1276 -1081 1277 -1080
rect 1283 -1081 1284 -1080
rect 513 -1083 514 -1082
rect 583 -1083 584 -1082
rect 642 -1083 643 -1082
rect 1458 -1083 1459 -1082
rect 513 -1085 514 -1084
rect 681 -1085 682 -1084
rect 828 -1085 829 -1084
rect 1094 -1085 1095 -1084
rect 79 -1087 80 -1086
rect 681 -1087 682 -1086
rect 814 -1087 815 -1086
rect 828 -1087 829 -1086
rect 978 -1087 979 -1086
rect 1059 -1087 1060 -1086
rect 79 -1089 80 -1088
rect 93 -1089 94 -1088
rect 653 -1089 654 -1088
rect 709 -1089 710 -1088
rect 807 -1089 808 -1088
rect 814 -1089 815 -1088
rect 1006 -1089 1007 -1088
rect 1276 -1089 1277 -1088
rect 93 -1091 94 -1090
rect 639 -1091 640 -1090
rect 674 -1091 675 -1090
rect 1346 -1091 1347 -1090
rect 499 -1093 500 -1092
rect 639 -1093 640 -1092
rect 709 -1093 710 -1092
rect 898 -1093 899 -1092
rect 807 -1095 808 -1094
rect 884 -1095 885 -1094
rect 898 -1095 899 -1094
rect 1087 -1095 1088 -1094
rect 1087 -1097 1088 -1096
rect 1150 -1097 1151 -1096
rect 23 -1108 24 -1107
rect 439 -1108 440 -1107
rect 471 -1108 472 -1107
rect 702 -1108 703 -1107
rect 730 -1108 731 -1107
rect 1241 -1108 1242 -1107
rect 1255 -1108 1256 -1107
rect 1381 -1108 1382 -1107
rect 1384 -1108 1385 -1107
rect 1626 -1108 1627 -1107
rect 1640 -1108 1641 -1107
rect 1724 -1108 1725 -1107
rect 1745 -1108 1746 -1107
rect 1759 -1108 1760 -1107
rect 23 -1110 24 -1109
rect 243 -1110 244 -1109
rect 275 -1110 276 -1109
rect 478 -1110 479 -1109
rect 499 -1110 500 -1109
rect 625 -1110 626 -1109
rect 649 -1110 650 -1109
rect 744 -1110 745 -1109
rect 765 -1110 766 -1109
rect 866 -1110 867 -1109
rect 887 -1110 888 -1109
rect 1374 -1110 1375 -1109
rect 1444 -1110 1445 -1109
rect 1661 -1110 1662 -1109
rect 1675 -1110 1676 -1109
rect 1703 -1110 1704 -1109
rect 37 -1112 38 -1111
rect 212 -1112 213 -1111
rect 219 -1112 220 -1111
rect 250 -1112 251 -1111
rect 275 -1112 276 -1111
rect 303 -1112 304 -1111
rect 324 -1112 325 -1111
rect 341 -1112 342 -1111
rect 401 -1112 402 -1111
rect 677 -1112 678 -1111
rect 681 -1112 682 -1111
rect 800 -1112 801 -1111
rect 817 -1112 818 -1111
rect 1185 -1112 1186 -1111
rect 1213 -1112 1214 -1111
rect 1381 -1112 1382 -1111
rect 1444 -1112 1445 -1111
rect 1766 -1112 1767 -1111
rect 72 -1114 73 -1113
rect 541 -1114 542 -1113
rect 656 -1114 657 -1113
rect 1346 -1114 1347 -1113
rect 1451 -1114 1452 -1113
rect 1563 -1114 1564 -1113
rect 1570 -1114 1571 -1113
rect 1717 -1114 1718 -1113
rect 75 -1116 76 -1115
rect 1675 -1116 1676 -1115
rect 1682 -1116 1683 -1115
rect 1769 -1116 1770 -1115
rect 89 -1118 90 -1117
rect 513 -1118 514 -1117
rect 516 -1118 517 -1117
rect 597 -1118 598 -1117
rect 681 -1118 682 -1117
rect 772 -1118 773 -1117
rect 835 -1118 836 -1117
rect 877 -1118 878 -1117
rect 929 -1118 930 -1117
rect 1297 -1118 1298 -1117
rect 1318 -1118 1319 -1117
rect 1451 -1118 1452 -1117
rect 1465 -1118 1466 -1117
rect 1682 -1118 1683 -1117
rect 93 -1120 94 -1119
rect 544 -1120 545 -1119
rect 548 -1120 549 -1119
rect 877 -1120 878 -1119
rect 933 -1120 934 -1119
rect 1374 -1120 1375 -1119
rect 1437 -1120 1438 -1119
rect 1563 -1120 1564 -1119
rect 1570 -1120 1571 -1119
rect 1605 -1120 1606 -1119
rect 1612 -1120 1613 -1119
rect 1752 -1120 1753 -1119
rect 93 -1122 94 -1121
rect 138 -1122 139 -1121
rect 173 -1122 174 -1121
rect 667 -1122 668 -1121
rect 688 -1122 689 -1121
rect 824 -1122 825 -1121
rect 859 -1122 860 -1121
rect 898 -1122 899 -1121
rect 912 -1122 913 -1121
rect 933 -1122 934 -1121
rect 950 -1122 951 -1121
rect 1304 -1122 1305 -1121
rect 1311 -1122 1312 -1121
rect 1437 -1122 1438 -1121
rect 1479 -1122 1480 -1121
rect 1605 -1122 1606 -1121
rect 1654 -1122 1655 -1121
rect 1780 -1122 1781 -1121
rect 100 -1124 101 -1123
rect 422 -1124 423 -1123
rect 506 -1124 507 -1123
rect 730 -1124 731 -1123
rect 737 -1124 738 -1123
rect 744 -1124 745 -1123
rect 758 -1124 759 -1123
rect 912 -1124 913 -1123
rect 1045 -1124 1046 -1123
rect 1234 -1124 1235 -1123
rect 1248 -1124 1249 -1123
rect 1612 -1124 1613 -1123
rect 58 -1126 59 -1125
rect 100 -1126 101 -1125
rect 107 -1126 108 -1125
rect 233 -1126 234 -1125
rect 236 -1126 237 -1125
rect 1472 -1126 1473 -1125
rect 1493 -1126 1494 -1125
rect 1619 -1126 1620 -1125
rect 58 -1128 59 -1127
rect 170 -1128 171 -1127
rect 177 -1128 178 -1127
rect 625 -1128 626 -1127
rect 653 -1128 654 -1127
rect 772 -1128 773 -1127
rect 891 -1128 892 -1127
rect 1311 -1128 1312 -1127
rect 1332 -1128 1333 -1127
rect 1454 -1128 1455 -1127
rect 1496 -1128 1497 -1127
rect 1647 -1128 1648 -1127
rect 68 -1130 69 -1129
rect 1248 -1130 1249 -1129
rect 1290 -1130 1291 -1129
rect 1619 -1130 1620 -1129
rect 89 -1132 90 -1131
rect 1493 -1132 1494 -1131
rect 1500 -1132 1501 -1131
rect 1640 -1132 1641 -1131
rect 110 -1134 111 -1133
rect 324 -1134 325 -1133
rect 380 -1134 381 -1133
rect 548 -1134 549 -1133
rect 698 -1134 699 -1133
rect 786 -1134 787 -1133
rect 891 -1134 892 -1133
rect 1290 -1134 1291 -1133
rect 1325 -1134 1326 -1133
rect 1500 -1134 1501 -1133
rect 1507 -1134 1508 -1133
rect 1647 -1134 1648 -1133
rect 121 -1136 122 -1135
rect 397 -1136 398 -1135
rect 401 -1136 402 -1135
rect 408 -1136 409 -1135
rect 415 -1136 416 -1135
rect 635 -1136 636 -1135
rect 716 -1136 717 -1135
rect 1213 -1136 1214 -1135
rect 1220 -1136 1221 -1135
rect 1710 -1136 1711 -1135
rect 121 -1138 122 -1137
rect 1626 -1138 1627 -1137
rect 128 -1140 129 -1139
rect 135 -1140 136 -1139
rect 180 -1140 181 -1139
rect 310 -1140 311 -1139
rect 380 -1140 381 -1139
rect 569 -1140 570 -1139
rect 649 -1140 650 -1139
rect 1220 -1140 1221 -1139
rect 1325 -1140 1326 -1139
rect 1430 -1140 1431 -1139
rect 1514 -1140 1515 -1139
rect 1668 -1140 1669 -1139
rect 128 -1142 129 -1141
rect 229 -1142 230 -1141
rect 233 -1142 234 -1141
rect 429 -1142 430 -1141
rect 485 -1142 486 -1141
rect 786 -1142 787 -1141
rect 919 -1142 920 -1141
rect 1045 -1142 1046 -1141
rect 1048 -1142 1049 -1141
rect 1199 -1142 1200 -1141
rect 1339 -1142 1340 -1141
rect 1507 -1142 1508 -1141
rect 1528 -1142 1529 -1141
rect 1689 -1142 1690 -1141
rect 184 -1144 185 -1143
rect 303 -1144 304 -1143
rect 387 -1144 388 -1143
rect 408 -1144 409 -1143
rect 415 -1144 416 -1143
rect 450 -1144 451 -1143
rect 492 -1144 493 -1143
rect 716 -1144 717 -1143
rect 723 -1144 724 -1143
rect 835 -1144 836 -1143
rect 968 -1144 969 -1143
rect 1332 -1144 1333 -1143
rect 1367 -1144 1368 -1143
rect 1514 -1144 1515 -1143
rect 1549 -1144 1550 -1143
rect 1696 -1144 1697 -1143
rect 79 -1146 80 -1145
rect 387 -1146 388 -1145
rect 443 -1146 444 -1145
rect 450 -1146 451 -1145
rect 499 -1146 500 -1145
rect 737 -1146 738 -1145
rect 758 -1146 759 -1145
rect 831 -1146 832 -1145
rect 1055 -1146 1056 -1145
rect 1353 -1146 1354 -1145
rect 1402 -1146 1403 -1145
rect 1528 -1146 1529 -1145
rect 1556 -1146 1557 -1145
rect 1738 -1146 1739 -1145
rect 51 -1148 52 -1147
rect 1353 -1148 1354 -1147
rect 1409 -1148 1410 -1147
rect 1654 -1148 1655 -1147
rect 51 -1150 52 -1149
rect 597 -1150 598 -1149
rect 611 -1150 612 -1149
rect 723 -1150 724 -1149
rect 765 -1150 766 -1149
rect 884 -1150 885 -1149
rect 1055 -1150 1056 -1149
rect 1185 -1150 1186 -1149
rect 1269 -1150 1270 -1149
rect 1367 -1150 1368 -1149
rect 1416 -1150 1417 -1149
rect 1549 -1150 1550 -1149
rect 1577 -1150 1578 -1149
rect 1731 -1150 1732 -1149
rect 65 -1152 66 -1151
rect 79 -1152 80 -1151
rect 124 -1152 125 -1151
rect 968 -1152 969 -1151
rect 1066 -1152 1067 -1151
rect 1255 -1152 1256 -1151
rect 1276 -1152 1277 -1151
rect 1402 -1152 1403 -1151
rect 1416 -1152 1417 -1151
rect 1745 -1152 1746 -1151
rect 65 -1154 66 -1153
rect 1479 -1154 1480 -1153
rect 1535 -1154 1536 -1153
rect 1556 -1154 1557 -1153
rect 1577 -1154 1578 -1153
rect 1633 -1154 1634 -1153
rect 142 -1156 143 -1155
rect 492 -1156 493 -1155
rect 520 -1156 521 -1155
rect 667 -1156 668 -1155
rect 768 -1156 769 -1155
rect 842 -1156 843 -1155
rect 905 -1156 906 -1155
rect 1269 -1156 1270 -1155
rect 1283 -1156 1284 -1155
rect 1409 -1156 1410 -1155
rect 1486 -1156 1487 -1155
rect 1633 -1156 1634 -1155
rect 184 -1158 185 -1157
rect 583 -1158 584 -1157
rect 779 -1158 780 -1157
rect 1430 -1158 1431 -1157
rect 1598 -1158 1599 -1157
rect 1787 -1158 1788 -1157
rect 198 -1160 199 -1159
rect 310 -1160 311 -1159
rect 338 -1160 339 -1159
rect 842 -1160 843 -1159
rect 880 -1160 881 -1159
rect 1283 -1160 1284 -1159
rect 1388 -1160 1389 -1159
rect 1535 -1160 1536 -1159
rect 198 -1162 199 -1161
rect 254 -1162 255 -1161
rect 282 -1162 283 -1161
rect 646 -1162 647 -1161
rect 793 -1162 794 -1161
rect 919 -1162 920 -1161
rect 1003 -1162 1004 -1161
rect 1276 -1162 1277 -1161
rect 1458 -1162 1459 -1161
rect 1598 -1162 1599 -1161
rect 177 -1164 178 -1163
rect 254 -1164 255 -1163
rect 261 -1164 262 -1163
rect 1003 -1164 1004 -1163
rect 1052 -1164 1053 -1163
rect 1486 -1164 1487 -1163
rect 212 -1166 213 -1165
rect 803 -1166 804 -1165
rect 821 -1166 822 -1165
rect 905 -1166 906 -1165
rect 1066 -1166 1067 -1165
rect 1542 -1166 1543 -1165
rect 219 -1168 220 -1167
rect 264 -1168 265 -1167
rect 282 -1168 283 -1167
rect 425 -1168 426 -1167
rect 443 -1168 444 -1167
rect 695 -1168 696 -1167
rect 793 -1168 794 -1167
rect 1073 -1168 1074 -1167
rect 1087 -1168 1088 -1167
rect 1129 -1168 1130 -1167
rect 1143 -1168 1144 -1167
rect 1388 -1168 1389 -1167
rect 1458 -1168 1459 -1167
rect 1591 -1168 1592 -1167
rect 226 -1170 227 -1169
rect 639 -1170 640 -1169
rect 688 -1170 689 -1169
rect 821 -1170 822 -1169
rect 961 -1170 962 -1169
rect 1073 -1170 1074 -1169
rect 1094 -1170 1095 -1169
rect 1346 -1170 1347 -1169
rect 1521 -1170 1522 -1169
rect 1542 -1170 1543 -1169
rect 1584 -1170 1585 -1169
rect 1591 -1170 1592 -1169
rect 30 -1172 31 -1171
rect 226 -1172 227 -1171
rect 247 -1172 248 -1171
rect 485 -1172 486 -1171
rect 520 -1172 521 -1171
rect 894 -1172 895 -1171
rect 996 -1172 997 -1171
rect 1094 -1172 1095 -1171
rect 1101 -1172 1102 -1171
rect 1199 -1172 1200 -1171
rect 1395 -1172 1396 -1171
rect 1521 -1172 1522 -1171
rect 30 -1174 31 -1173
rect 86 -1174 87 -1173
rect 205 -1174 206 -1173
rect 247 -1174 248 -1173
rect 296 -1174 297 -1173
rect 429 -1174 430 -1173
rect 471 -1174 472 -1173
rect 894 -1174 895 -1173
rect 1010 -1174 1011 -1173
rect 1129 -1174 1130 -1173
rect 1150 -1174 1151 -1173
rect 1241 -1174 1242 -1173
rect 86 -1176 87 -1175
rect 163 -1176 164 -1175
rect 205 -1176 206 -1175
rect 457 -1176 458 -1175
rect 527 -1176 528 -1175
rect 611 -1176 612 -1175
rect 618 -1176 619 -1175
rect 639 -1176 640 -1175
rect 695 -1176 696 -1175
rect 1360 -1176 1361 -1175
rect 149 -1178 150 -1177
rect 163 -1178 164 -1177
rect 289 -1178 290 -1177
rect 296 -1178 297 -1177
rect 338 -1178 339 -1177
rect 436 -1178 437 -1177
rect 457 -1178 458 -1177
rect 534 -1178 535 -1177
rect 569 -1178 570 -1177
rect 709 -1178 710 -1177
rect 828 -1178 829 -1177
rect 961 -1178 962 -1177
rect 982 -1178 983 -1177
rect 1010 -1178 1011 -1177
rect 1017 -1178 1018 -1177
rect 1087 -1178 1088 -1177
rect 1101 -1178 1102 -1177
rect 1136 -1178 1137 -1177
rect 1157 -1178 1158 -1177
rect 1234 -1178 1235 -1177
rect 1360 -1178 1361 -1177
rect 1748 -1178 1749 -1177
rect 145 -1180 146 -1179
rect 149 -1180 150 -1179
rect 170 -1180 171 -1179
rect 1136 -1180 1137 -1179
rect 1164 -1180 1165 -1179
rect 1465 -1180 1466 -1179
rect 268 -1182 269 -1181
rect 436 -1182 437 -1181
rect 464 -1182 465 -1181
rect 534 -1182 535 -1181
rect 562 -1182 563 -1181
rect 709 -1182 710 -1181
rect 740 -1182 741 -1181
rect 1164 -1182 1165 -1181
rect 1171 -1182 1172 -1181
rect 1318 -1182 1319 -1181
rect 142 -1184 143 -1183
rect 268 -1184 269 -1183
rect 331 -1184 332 -1183
rect 464 -1184 465 -1183
rect 562 -1184 563 -1183
rect 674 -1184 675 -1183
rect 849 -1184 850 -1183
rect 1017 -1184 1018 -1183
rect 1038 -1184 1039 -1183
rect 1171 -1184 1172 -1183
rect 1178 -1184 1179 -1183
rect 1339 -1184 1340 -1183
rect 331 -1186 332 -1185
rect 359 -1186 360 -1185
rect 576 -1186 577 -1185
rect 779 -1186 780 -1185
rect 856 -1186 857 -1185
rect 982 -1186 983 -1185
rect 1059 -1186 1060 -1185
rect 1143 -1186 1144 -1185
rect 1178 -1186 1179 -1185
rect 1206 -1186 1207 -1185
rect 1227 -1186 1228 -1185
rect 1395 -1186 1396 -1185
rect 345 -1188 346 -1187
rect 359 -1188 360 -1187
rect 555 -1188 556 -1187
rect 576 -1188 577 -1187
rect 583 -1188 584 -1187
rect 733 -1188 734 -1187
rect 751 -1188 752 -1187
rect 849 -1188 850 -1187
rect 856 -1188 857 -1187
rect 996 -1188 997 -1187
rect 1080 -1188 1081 -1187
rect 1206 -1188 1207 -1187
rect 1227 -1188 1228 -1187
rect 1262 -1188 1263 -1187
rect 345 -1190 346 -1189
rect 481 -1190 482 -1189
rect 555 -1190 556 -1189
rect 632 -1190 633 -1189
rect 674 -1190 675 -1189
rect 807 -1190 808 -1189
rect 926 -1190 927 -1189
rect 1059 -1190 1060 -1189
rect 1108 -1190 1109 -1189
rect 1150 -1190 1151 -1189
rect 1192 -1190 1193 -1189
rect 1584 -1190 1585 -1189
rect 394 -1192 395 -1191
rect 1080 -1192 1081 -1191
rect 1115 -1192 1116 -1191
rect 1297 -1192 1298 -1191
rect 352 -1194 353 -1193
rect 394 -1194 395 -1193
rect 618 -1194 619 -1193
rect 828 -1194 829 -1193
rect 898 -1194 899 -1193
rect 926 -1194 927 -1193
rect 940 -1194 941 -1193
rect 1038 -1194 1039 -1193
rect 1122 -1194 1123 -1193
rect 1304 -1194 1305 -1193
rect 352 -1196 353 -1195
rect 373 -1196 374 -1195
rect 691 -1196 692 -1195
rect 1108 -1196 1109 -1195
rect 1262 -1196 1263 -1195
rect 1475 -1196 1476 -1195
rect 317 -1198 318 -1197
rect 373 -1198 374 -1197
rect 702 -1198 703 -1197
rect 1115 -1198 1116 -1197
rect 44 -1200 45 -1199
rect 317 -1200 318 -1199
rect 751 -1200 752 -1199
rect 863 -1200 864 -1199
rect 947 -1200 948 -1199
rect 1157 -1200 1158 -1199
rect 44 -1202 45 -1201
rect 156 -1202 157 -1201
rect 541 -1202 542 -1201
rect 863 -1202 864 -1201
rect 947 -1202 948 -1201
rect 1024 -1202 1025 -1201
rect 1031 -1202 1032 -1201
rect 1122 -1202 1123 -1201
rect 156 -1204 157 -1203
rect 590 -1204 591 -1203
rect 796 -1204 797 -1203
rect 807 -1204 808 -1203
rect 954 -1204 955 -1203
rect 1031 -1204 1032 -1203
rect 590 -1206 591 -1205
rect 660 -1206 661 -1205
rect 698 -1206 699 -1205
rect 954 -1206 955 -1205
rect 975 -1206 976 -1205
rect 1024 -1206 1025 -1205
rect 604 -1208 605 -1207
rect 660 -1208 661 -1207
rect 814 -1208 815 -1207
rect 975 -1208 976 -1207
rect 989 -1208 990 -1207
rect 1192 -1208 1193 -1207
rect 527 -1210 528 -1209
rect 604 -1210 605 -1209
rect 814 -1210 815 -1209
rect 940 -1210 941 -1209
rect 870 -1212 871 -1211
rect 989 -1212 990 -1211
rect 240 -1214 241 -1213
rect 870 -1214 871 -1213
rect 240 -1216 241 -1215
rect 289 -1216 290 -1215
rect 16 -1227 17 -1226
rect 446 -1227 447 -1226
rect 506 -1227 507 -1226
rect 863 -1227 864 -1226
rect 891 -1227 892 -1226
rect 1087 -1227 1088 -1226
rect 1094 -1227 1095 -1226
rect 1202 -1227 1203 -1226
rect 1290 -1227 1291 -1226
rect 1293 -1227 1294 -1226
rect 1311 -1227 1312 -1226
rect 1314 -1227 1315 -1226
rect 1703 -1227 1704 -1226
rect 1748 -1227 1749 -1226
rect 1766 -1227 1767 -1226
rect 1787 -1227 1788 -1226
rect 44 -1229 45 -1228
rect 264 -1229 265 -1228
rect 289 -1229 290 -1228
rect 509 -1229 510 -1228
rect 548 -1229 549 -1228
rect 565 -1229 566 -1228
rect 590 -1229 591 -1228
rect 597 -1229 598 -1228
rect 607 -1229 608 -1228
rect 1269 -1229 1270 -1228
rect 1290 -1229 1291 -1228
rect 1304 -1229 1305 -1228
rect 1311 -1229 1312 -1228
rect 1318 -1229 1319 -1228
rect 1696 -1229 1697 -1228
rect 1703 -1229 1704 -1228
rect 1745 -1229 1746 -1228
rect 1759 -1229 1760 -1228
rect 44 -1231 45 -1230
rect 89 -1231 90 -1230
rect 103 -1231 104 -1230
rect 303 -1231 304 -1230
rect 345 -1231 346 -1230
rect 796 -1231 797 -1230
rect 800 -1231 801 -1230
rect 863 -1231 864 -1230
rect 894 -1231 895 -1230
rect 1612 -1231 1613 -1230
rect 1745 -1231 1746 -1230
rect 1776 -1231 1777 -1230
rect 65 -1233 66 -1232
rect 1353 -1233 1354 -1232
rect 1612 -1233 1613 -1232
rect 1717 -1233 1718 -1232
rect 54 -1235 55 -1234
rect 65 -1235 66 -1234
rect 68 -1235 69 -1234
rect 79 -1235 80 -1234
rect 107 -1235 108 -1234
rect 114 -1235 115 -1234
rect 121 -1235 122 -1234
rect 1374 -1235 1375 -1234
rect 1717 -1235 1718 -1234
rect 1731 -1235 1732 -1234
rect 72 -1237 73 -1236
rect 653 -1237 654 -1236
rect 709 -1237 710 -1236
rect 793 -1237 794 -1236
rect 817 -1237 818 -1236
rect 961 -1237 962 -1236
rect 1010 -1237 1011 -1236
rect 1094 -1237 1095 -1236
rect 1146 -1237 1147 -1236
rect 1465 -1237 1466 -1236
rect 51 -1239 52 -1238
rect 72 -1239 73 -1238
rect 110 -1239 111 -1238
rect 660 -1239 661 -1238
rect 667 -1239 668 -1238
rect 793 -1239 794 -1238
rect 821 -1239 822 -1238
rect 1619 -1239 1620 -1238
rect 114 -1241 115 -1240
rect 940 -1241 941 -1240
rect 947 -1241 948 -1240
rect 1535 -1241 1536 -1240
rect 121 -1243 122 -1242
rect 453 -1243 454 -1242
rect 551 -1243 552 -1242
rect 1136 -1243 1137 -1242
rect 1248 -1243 1249 -1242
rect 1269 -1243 1270 -1242
rect 1314 -1243 1315 -1242
rect 1318 -1243 1319 -1242
rect 1353 -1243 1354 -1242
rect 1479 -1243 1480 -1242
rect 1486 -1243 1487 -1242
rect 1535 -1243 1536 -1242
rect 124 -1245 125 -1244
rect 478 -1245 479 -1244
rect 565 -1245 566 -1244
rect 716 -1245 717 -1244
rect 737 -1245 738 -1244
rect 744 -1245 745 -1244
rect 751 -1245 752 -1244
rect 765 -1245 766 -1244
rect 779 -1245 780 -1244
rect 800 -1245 801 -1244
rect 821 -1245 822 -1244
rect 1542 -1245 1543 -1244
rect 61 -1247 62 -1246
rect 737 -1247 738 -1246
rect 740 -1247 741 -1246
rect 1332 -1247 1333 -1246
rect 1360 -1247 1361 -1246
rect 1374 -1247 1375 -1246
rect 1458 -1247 1459 -1246
rect 1731 -1247 1732 -1246
rect 145 -1249 146 -1248
rect 1556 -1249 1557 -1248
rect 170 -1251 171 -1250
rect 177 -1251 178 -1250
rect 180 -1251 181 -1250
rect 1738 -1251 1739 -1250
rect 142 -1253 143 -1252
rect 170 -1253 171 -1252
rect 177 -1253 178 -1252
rect 198 -1253 199 -1252
rect 208 -1253 209 -1252
rect 240 -1253 241 -1252
rect 243 -1253 244 -1252
rect 1157 -1253 1158 -1252
rect 1220 -1253 1221 -1252
rect 1248 -1253 1249 -1252
rect 1325 -1253 1326 -1252
rect 1556 -1253 1557 -1252
rect 142 -1255 143 -1254
rect 212 -1255 213 -1254
rect 226 -1255 227 -1254
rect 1003 -1255 1004 -1254
rect 1010 -1255 1011 -1254
rect 1045 -1255 1046 -1254
rect 1052 -1255 1053 -1254
rect 1584 -1255 1585 -1254
rect 128 -1257 129 -1256
rect 212 -1257 213 -1256
rect 226 -1257 227 -1256
rect 254 -1257 255 -1256
rect 261 -1257 262 -1256
rect 436 -1257 437 -1256
rect 443 -1257 444 -1256
rect 1020 -1257 1021 -1256
rect 1059 -1257 1060 -1256
rect 1157 -1257 1158 -1256
rect 1171 -1257 1172 -1256
rect 1220 -1257 1221 -1256
rect 1325 -1257 1326 -1256
rect 1769 -1257 1770 -1256
rect 163 -1259 164 -1258
rect 254 -1259 255 -1258
rect 292 -1259 293 -1258
rect 870 -1259 871 -1258
rect 933 -1259 934 -1258
rect 1059 -1259 1060 -1258
rect 1087 -1259 1088 -1258
rect 1500 -1259 1501 -1258
rect 1542 -1259 1543 -1258
rect 1549 -1259 1550 -1258
rect 1584 -1259 1585 -1258
rect 1591 -1259 1592 -1258
rect 163 -1261 164 -1260
rect 705 -1261 706 -1260
rect 723 -1261 724 -1260
rect 744 -1261 745 -1260
rect 751 -1261 752 -1260
rect 768 -1261 769 -1260
rect 824 -1261 825 -1260
rect 1055 -1261 1056 -1260
rect 1101 -1261 1102 -1260
rect 1332 -1261 1333 -1260
rect 1402 -1261 1403 -1260
rect 1458 -1261 1459 -1260
rect 1465 -1261 1466 -1260
rect 1507 -1261 1508 -1260
rect 1549 -1261 1550 -1260
rect 1598 -1261 1599 -1260
rect 184 -1263 185 -1262
rect 709 -1263 710 -1262
rect 740 -1263 741 -1262
rect 1430 -1263 1431 -1262
rect 1479 -1263 1480 -1262
rect 1640 -1263 1641 -1262
rect 184 -1265 185 -1264
rect 618 -1265 619 -1264
rect 632 -1265 633 -1264
rect 1346 -1265 1347 -1264
rect 1402 -1265 1403 -1264
rect 1444 -1265 1445 -1264
rect 1486 -1265 1487 -1264
rect 1528 -1265 1529 -1264
rect 1570 -1265 1571 -1264
rect 1591 -1265 1592 -1264
rect 1598 -1265 1599 -1264
rect 1633 -1265 1634 -1264
rect 1640 -1265 1641 -1264
rect 1654 -1265 1655 -1264
rect 198 -1267 199 -1266
rect 779 -1267 780 -1266
rect 828 -1267 829 -1266
rect 1360 -1267 1361 -1266
rect 1423 -1267 1424 -1266
rect 1507 -1267 1508 -1266
rect 1528 -1267 1529 -1266
rect 1577 -1267 1578 -1266
rect 1633 -1267 1634 -1266
rect 1647 -1267 1648 -1266
rect 1654 -1267 1655 -1266
rect 1675 -1267 1676 -1266
rect 296 -1269 297 -1268
rect 604 -1269 605 -1268
rect 611 -1269 612 -1268
rect 632 -1269 633 -1268
rect 639 -1269 640 -1268
rect 660 -1269 661 -1268
rect 831 -1269 832 -1268
rect 1255 -1269 1256 -1268
rect 1339 -1269 1340 -1268
rect 1346 -1269 1347 -1268
rect 1423 -1269 1424 -1268
rect 1514 -1269 1515 -1268
rect 1577 -1269 1578 -1268
rect 1626 -1269 1627 -1268
rect 1647 -1269 1648 -1268
rect 1668 -1269 1669 -1268
rect 1675 -1269 1676 -1268
rect 1689 -1269 1690 -1268
rect 58 -1271 59 -1270
rect 604 -1271 605 -1270
rect 611 -1271 612 -1270
rect 912 -1271 913 -1270
rect 922 -1271 923 -1270
rect 1570 -1271 1571 -1270
rect 1682 -1271 1683 -1270
rect 1689 -1271 1690 -1270
rect 58 -1273 59 -1272
rect 100 -1273 101 -1272
rect 296 -1273 297 -1272
rect 352 -1273 353 -1272
rect 380 -1273 381 -1272
rect 695 -1273 696 -1272
rect 702 -1273 703 -1272
rect 1339 -1273 1340 -1272
rect 1500 -1273 1501 -1272
rect 1521 -1273 1522 -1272
rect 1682 -1273 1683 -1272
rect 1710 -1273 1711 -1272
rect 205 -1275 206 -1274
rect 352 -1275 353 -1274
rect 380 -1275 381 -1274
rect 597 -1275 598 -1274
rect 600 -1275 601 -1274
rect 639 -1275 640 -1274
rect 688 -1275 689 -1274
rect 702 -1275 703 -1274
rect 831 -1275 832 -1274
rect 1262 -1275 1263 -1274
rect 1710 -1275 1711 -1274
rect 1724 -1275 1725 -1274
rect 23 -1277 24 -1276
rect 205 -1277 206 -1276
rect 303 -1277 304 -1276
rect 331 -1277 332 -1276
rect 345 -1277 346 -1276
rect 373 -1277 374 -1276
rect 387 -1277 388 -1276
rect 590 -1277 591 -1276
rect 681 -1277 682 -1276
rect 688 -1277 689 -1276
rect 835 -1277 836 -1276
rect 891 -1277 892 -1276
rect 912 -1277 913 -1276
rect 982 -1277 983 -1276
rect 996 -1277 997 -1276
rect 1045 -1277 1046 -1276
rect 1101 -1277 1102 -1276
rect 1472 -1277 1473 -1276
rect 1724 -1277 1725 -1276
rect 1752 -1277 1753 -1276
rect 23 -1279 24 -1278
rect 541 -1279 542 -1278
rect 548 -1279 549 -1278
rect 1255 -1279 1256 -1278
rect 1752 -1279 1753 -1278
rect 1780 -1279 1781 -1278
rect 310 -1281 311 -1280
rect 716 -1281 717 -1280
rect 852 -1281 853 -1280
rect 919 -1281 920 -1280
rect 929 -1281 930 -1280
rect 1668 -1281 1669 -1280
rect 156 -1283 157 -1282
rect 310 -1283 311 -1282
rect 317 -1283 318 -1282
rect 387 -1283 388 -1282
rect 415 -1283 416 -1282
rect 506 -1283 507 -1282
rect 513 -1283 514 -1282
rect 870 -1283 871 -1282
rect 933 -1283 934 -1282
rect 1696 -1283 1697 -1282
rect 149 -1285 150 -1284
rect 156 -1285 157 -1284
rect 317 -1285 318 -1284
rect 789 -1285 790 -1284
rect 856 -1285 857 -1284
rect 1493 -1285 1494 -1284
rect 100 -1287 101 -1286
rect 1493 -1287 1494 -1286
rect 149 -1289 150 -1288
rect 877 -1289 878 -1288
rect 936 -1289 937 -1288
rect 1297 -1289 1298 -1288
rect 331 -1291 332 -1290
rect 359 -1291 360 -1290
rect 366 -1291 367 -1290
rect 541 -1291 542 -1290
rect 625 -1291 626 -1290
rect 681 -1291 682 -1290
rect 807 -1291 808 -1290
rect 877 -1291 878 -1290
rect 940 -1291 941 -1290
rect 1006 -1291 1007 -1290
rect 1017 -1291 1018 -1290
rect 1052 -1291 1053 -1290
rect 1104 -1291 1105 -1290
rect 1619 -1291 1620 -1290
rect 275 -1293 276 -1292
rect 625 -1293 626 -1292
rect 667 -1293 668 -1292
rect 982 -1293 983 -1292
rect 1038 -1293 1039 -1292
rect 1626 -1293 1627 -1292
rect 135 -1295 136 -1294
rect 275 -1295 276 -1294
rect 282 -1295 283 -1294
rect 366 -1295 367 -1294
rect 373 -1295 374 -1294
rect 464 -1295 465 -1294
rect 499 -1295 500 -1294
rect 723 -1295 724 -1294
rect 772 -1295 773 -1294
rect 807 -1295 808 -1294
rect 842 -1295 843 -1294
rect 856 -1295 857 -1294
rect 859 -1295 860 -1294
rect 1073 -1295 1074 -1294
rect 1115 -1295 1116 -1294
rect 1738 -1295 1739 -1294
rect 82 -1297 83 -1296
rect 135 -1297 136 -1296
rect 187 -1297 188 -1296
rect 499 -1297 500 -1296
rect 635 -1297 636 -1296
rect 1038 -1297 1039 -1296
rect 1108 -1297 1109 -1296
rect 1115 -1297 1116 -1296
rect 1129 -1297 1130 -1296
rect 1136 -1297 1137 -1296
rect 1150 -1297 1151 -1296
rect 1297 -1297 1298 -1296
rect 191 -1299 192 -1298
rect 464 -1299 465 -1298
rect 558 -1299 559 -1298
rect 1129 -1299 1130 -1298
rect 1143 -1299 1144 -1298
rect 1150 -1299 1151 -1298
rect 1164 -1299 1165 -1298
rect 1171 -1299 1172 -1298
rect 1192 -1299 1193 -1298
rect 1521 -1299 1522 -1298
rect 191 -1301 192 -1300
rect 975 -1301 976 -1300
rect 1031 -1301 1032 -1300
rect 1073 -1301 1074 -1300
rect 1080 -1301 1081 -1300
rect 1108 -1301 1109 -1300
rect 1164 -1301 1165 -1300
rect 1206 -1301 1207 -1300
rect 1227 -1301 1228 -1300
rect 1472 -1301 1473 -1300
rect 247 -1303 248 -1302
rect 282 -1303 283 -1302
rect 338 -1303 339 -1302
rect 415 -1303 416 -1302
rect 422 -1303 423 -1302
rect 835 -1303 836 -1302
rect 950 -1303 951 -1302
rect 1514 -1303 1515 -1302
rect 173 -1305 174 -1304
rect 338 -1305 339 -1304
rect 359 -1305 360 -1304
rect 656 -1305 657 -1304
rect 674 -1305 675 -1304
rect 772 -1305 773 -1304
rect 950 -1305 951 -1304
rect 961 -1305 962 -1304
rect 989 -1305 990 -1304
rect 1031 -1305 1032 -1304
rect 1080 -1305 1081 -1304
rect 1185 -1305 1186 -1304
rect 1206 -1305 1207 -1304
rect 1213 -1305 1214 -1304
rect 1234 -1305 1235 -1304
rect 1430 -1305 1431 -1304
rect 86 -1307 87 -1306
rect 674 -1307 675 -1306
rect 695 -1307 696 -1306
rect 1213 -1307 1214 -1306
rect 1241 -1307 1242 -1306
rect 1262 -1307 1263 -1306
rect 86 -1309 87 -1308
rect 527 -1309 528 -1308
rect 562 -1309 563 -1308
rect 1192 -1309 1193 -1308
rect 247 -1311 248 -1310
rect 268 -1311 269 -1310
rect 408 -1311 409 -1310
rect 842 -1311 843 -1310
rect 926 -1311 927 -1310
rect 1234 -1311 1235 -1310
rect 222 -1313 223 -1312
rect 268 -1313 269 -1312
rect 324 -1313 325 -1312
rect 408 -1313 409 -1312
rect 422 -1313 423 -1312
rect 754 -1313 755 -1312
rect 898 -1313 899 -1312
rect 926 -1313 927 -1312
rect 954 -1313 955 -1312
rect 989 -1313 990 -1312
rect 1003 -1313 1004 -1312
rect 1185 -1313 1186 -1312
rect 324 -1315 325 -1314
rect 968 -1315 969 -1314
rect 1024 -1315 1025 -1314
rect 1241 -1315 1242 -1314
rect 436 -1317 437 -1316
rect 758 -1317 759 -1316
rect 849 -1317 850 -1316
rect 1024 -1317 1025 -1316
rect 450 -1319 451 -1318
rect 478 -1319 479 -1318
rect 485 -1319 486 -1318
rect 562 -1319 563 -1318
rect 572 -1319 573 -1318
rect 1227 -1319 1228 -1318
rect 450 -1321 451 -1320
rect 996 -1321 997 -1320
rect 457 -1323 458 -1322
rect 513 -1323 514 -1322
rect 555 -1323 556 -1322
rect 758 -1323 759 -1322
rect 884 -1323 885 -1322
rect 968 -1323 969 -1322
rect 401 -1325 402 -1324
rect 555 -1325 556 -1324
rect 583 -1325 584 -1324
rect 898 -1325 899 -1324
rect 905 -1325 906 -1324
rect 954 -1325 955 -1324
rect 394 -1327 395 -1326
rect 401 -1327 402 -1326
rect 429 -1327 430 -1326
rect 884 -1327 885 -1326
rect 219 -1329 220 -1328
rect 429 -1329 430 -1328
rect 457 -1329 458 -1328
rect 534 -1329 535 -1328
rect 618 -1329 619 -1328
rect 849 -1329 850 -1328
rect 394 -1331 395 -1330
rect 576 -1331 577 -1330
rect 698 -1331 699 -1330
rect 975 -1331 976 -1330
rect 37 -1333 38 -1332
rect 576 -1333 577 -1332
rect 786 -1333 787 -1332
rect 905 -1333 906 -1332
rect 492 -1335 493 -1334
rect 527 -1335 528 -1334
rect 534 -1335 535 -1334
rect 814 -1335 815 -1334
rect 233 -1337 234 -1336
rect 492 -1337 493 -1336
rect 520 -1337 521 -1336
rect 583 -1337 584 -1336
rect 646 -1337 647 -1336
rect 814 -1337 815 -1336
rect 30 -1339 31 -1338
rect 233 -1339 234 -1338
rect 520 -1339 521 -1338
rect 730 -1339 731 -1338
rect 786 -1339 787 -1338
rect 1367 -1339 1368 -1338
rect 30 -1341 31 -1340
rect 569 -1341 570 -1340
rect 730 -1341 731 -1340
rect 1066 -1341 1067 -1340
rect 1367 -1341 1368 -1340
rect 1381 -1341 1382 -1340
rect 485 -1343 486 -1342
rect 569 -1343 570 -1342
rect 1066 -1343 1067 -1342
rect 1122 -1343 1123 -1342
rect 1381 -1343 1382 -1342
rect 1388 -1343 1389 -1342
rect 1122 -1345 1123 -1344
rect 1199 -1345 1200 -1344
rect 1388 -1345 1389 -1344
rect 1395 -1345 1396 -1344
rect 1199 -1347 1200 -1346
rect 1444 -1347 1445 -1346
rect 1395 -1349 1396 -1348
rect 1409 -1349 1410 -1348
rect 1409 -1351 1410 -1350
rect 1416 -1351 1417 -1350
rect 1416 -1353 1417 -1352
rect 1437 -1353 1438 -1352
rect 1437 -1355 1438 -1354
rect 1563 -1355 1564 -1354
rect 1563 -1357 1564 -1356
rect 1605 -1357 1606 -1356
rect 817 -1359 818 -1358
rect 1605 -1359 1606 -1358
rect 16 -1370 17 -1369
rect 110 -1370 111 -1369
rect 121 -1370 122 -1369
rect 208 -1370 209 -1369
rect 219 -1370 220 -1369
rect 1038 -1370 1039 -1369
rect 1048 -1370 1049 -1369
rect 1094 -1370 1095 -1369
rect 1104 -1370 1105 -1369
rect 1689 -1370 1690 -1369
rect 1738 -1370 1739 -1369
rect 1801 -1370 1802 -1369
rect 51 -1372 52 -1371
rect 93 -1372 94 -1371
rect 107 -1372 108 -1371
rect 646 -1372 647 -1371
rect 719 -1372 720 -1371
rect 1024 -1372 1025 -1371
rect 1038 -1372 1039 -1371
rect 1108 -1372 1109 -1371
rect 1146 -1372 1147 -1371
rect 1661 -1372 1662 -1371
rect 1689 -1372 1690 -1371
rect 1696 -1372 1697 -1371
rect 51 -1374 52 -1373
rect 149 -1374 150 -1373
rect 159 -1374 160 -1373
rect 177 -1374 178 -1373
rect 187 -1374 188 -1373
rect 765 -1374 766 -1373
rect 814 -1374 815 -1373
rect 1136 -1374 1137 -1373
rect 1199 -1374 1200 -1373
rect 1346 -1374 1347 -1373
rect 1591 -1374 1592 -1373
rect 1696 -1374 1697 -1373
rect 58 -1376 59 -1375
rect 618 -1376 619 -1375
rect 646 -1376 647 -1375
rect 660 -1376 661 -1375
rect 751 -1376 752 -1375
rect 1290 -1376 1291 -1375
rect 1346 -1376 1347 -1375
rect 1395 -1376 1396 -1375
rect 1591 -1376 1592 -1375
rect 1633 -1376 1634 -1375
rect 65 -1378 66 -1377
rect 79 -1378 80 -1377
rect 82 -1378 83 -1377
rect 1374 -1378 1375 -1377
rect 1395 -1378 1396 -1377
rect 1402 -1378 1403 -1377
rect 1528 -1378 1529 -1377
rect 1633 -1378 1634 -1377
rect 79 -1380 80 -1379
rect 940 -1380 941 -1379
rect 978 -1380 979 -1379
rect 1500 -1380 1501 -1379
rect 1612 -1380 1613 -1379
rect 1661 -1380 1662 -1379
rect 93 -1382 94 -1381
rect 520 -1382 521 -1381
rect 551 -1382 552 -1381
rect 835 -1382 836 -1381
rect 849 -1382 850 -1381
rect 1325 -1382 1326 -1381
rect 1374 -1382 1375 -1381
rect 1409 -1382 1410 -1381
rect 1437 -1382 1438 -1381
rect 1528 -1382 1529 -1381
rect 1612 -1382 1613 -1381
rect 1647 -1382 1648 -1381
rect 124 -1384 125 -1383
rect 716 -1384 717 -1383
rect 751 -1384 752 -1383
rect 758 -1384 759 -1383
rect 761 -1384 762 -1383
rect 1626 -1384 1627 -1383
rect 1647 -1384 1648 -1383
rect 1682 -1384 1683 -1383
rect 149 -1386 150 -1385
rect 824 -1386 825 -1385
rect 831 -1386 832 -1385
rect 1220 -1386 1221 -1385
rect 1227 -1386 1228 -1385
rect 1409 -1386 1410 -1385
rect 1500 -1386 1501 -1385
rect 1556 -1386 1557 -1385
rect 1626 -1386 1627 -1385
rect 1675 -1386 1676 -1385
rect 156 -1388 157 -1387
rect 177 -1388 178 -1387
rect 194 -1388 195 -1387
rect 282 -1388 283 -1387
rect 289 -1388 290 -1387
rect 471 -1388 472 -1387
rect 478 -1388 479 -1387
rect 516 -1388 517 -1387
rect 520 -1388 521 -1387
rect 1031 -1388 1032 -1387
rect 1034 -1388 1035 -1387
rect 1682 -1388 1683 -1387
rect 103 -1390 104 -1389
rect 1031 -1390 1032 -1389
rect 1066 -1390 1067 -1389
rect 1094 -1390 1095 -1389
rect 1108 -1390 1109 -1389
rect 1248 -1390 1249 -1389
rect 1402 -1390 1403 -1389
rect 1587 -1390 1588 -1389
rect 156 -1392 157 -1391
rect 292 -1392 293 -1391
rect 317 -1392 318 -1391
rect 618 -1392 619 -1391
rect 625 -1392 626 -1391
rect 660 -1392 661 -1391
rect 758 -1392 759 -1391
rect 1325 -1392 1326 -1391
rect 1556 -1392 1557 -1391
rect 1563 -1392 1564 -1391
rect 170 -1394 171 -1393
rect 205 -1394 206 -1393
rect 219 -1394 220 -1393
rect 310 -1394 311 -1393
rect 324 -1394 325 -1393
rect 670 -1394 671 -1393
rect 786 -1394 787 -1393
rect 1136 -1394 1137 -1393
rect 1202 -1394 1203 -1393
rect 1703 -1394 1704 -1393
rect 114 -1396 115 -1395
rect 205 -1396 206 -1395
rect 222 -1396 223 -1395
rect 1339 -1396 1340 -1395
rect 1563 -1396 1564 -1395
rect 1668 -1396 1669 -1395
rect 114 -1398 115 -1397
rect 716 -1398 717 -1397
rect 789 -1398 790 -1397
rect 940 -1398 941 -1397
rect 982 -1398 983 -1397
rect 1731 -1398 1732 -1397
rect 170 -1400 171 -1399
rect 639 -1400 640 -1399
rect 817 -1400 818 -1399
rect 1220 -1400 1221 -1399
rect 1227 -1400 1228 -1399
rect 1255 -1400 1256 -1399
rect 1339 -1400 1340 -1399
rect 1381 -1400 1382 -1399
rect 1584 -1400 1585 -1399
rect 1668 -1400 1669 -1399
rect 1731 -1400 1732 -1399
rect 1745 -1400 1746 -1399
rect 163 -1402 164 -1401
rect 639 -1402 640 -1401
rect 821 -1402 822 -1401
rect 1332 -1402 1333 -1401
rect 1381 -1402 1382 -1401
rect 1430 -1402 1431 -1401
rect 1584 -1402 1585 -1401
rect 1703 -1402 1704 -1401
rect 163 -1404 164 -1403
rect 254 -1404 255 -1403
rect 257 -1404 258 -1403
rect 611 -1404 612 -1403
rect 849 -1404 850 -1403
rect 891 -1404 892 -1403
rect 919 -1404 920 -1403
rect 1608 -1404 1609 -1403
rect 198 -1406 199 -1405
rect 541 -1406 542 -1405
rect 555 -1406 556 -1405
rect 905 -1406 906 -1405
rect 919 -1406 920 -1405
rect 926 -1406 927 -1405
rect 982 -1406 983 -1405
rect 996 -1406 997 -1405
rect 1003 -1406 1004 -1405
rect 1213 -1406 1214 -1405
rect 1216 -1406 1217 -1405
rect 1507 -1406 1508 -1405
rect 54 -1408 55 -1407
rect 996 -1408 997 -1407
rect 1006 -1408 1007 -1407
rect 1472 -1408 1473 -1407
rect 1507 -1408 1508 -1407
rect 1598 -1408 1599 -1407
rect 135 -1410 136 -1409
rect 198 -1410 199 -1409
rect 201 -1410 202 -1409
rect 1437 -1410 1438 -1409
rect 1472 -1410 1473 -1409
rect 1605 -1410 1606 -1409
rect 135 -1412 136 -1411
rect 142 -1412 143 -1411
rect 226 -1412 227 -1411
rect 282 -1412 283 -1411
rect 310 -1412 311 -1411
rect 457 -1412 458 -1411
rect 471 -1412 472 -1411
rect 485 -1412 486 -1411
rect 506 -1412 507 -1411
rect 555 -1412 556 -1411
rect 558 -1412 559 -1411
rect 1570 -1412 1571 -1411
rect 1598 -1412 1599 -1411
rect 1724 -1412 1725 -1411
rect 142 -1414 143 -1413
rect 212 -1414 213 -1413
rect 229 -1414 230 -1413
rect 303 -1414 304 -1413
rect 366 -1414 367 -1413
rect 485 -1414 486 -1413
rect 541 -1414 542 -1413
rect 933 -1414 934 -1413
rect 1010 -1414 1011 -1413
rect 1024 -1414 1025 -1413
rect 1066 -1414 1067 -1413
rect 1115 -1414 1116 -1413
rect 1157 -1414 1158 -1413
rect 1605 -1414 1606 -1413
rect 191 -1416 192 -1415
rect 212 -1416 213 -1415
rect 215 -1416 216 -1415
rect 366 -1416 367 -1415
rect 380 -1416 381 -1415
rect 506 -1416 507 -1415
rect 562 -1416 563 -1415
rect 835 -1416 836 -1415
rect 891 -1416 892 -1415
rect 954 -1416 955 -1415
rect 1010 -1416 1011 -1415
rect 1059 -1416 1060 -1415
rect 1115 -1416 1116 -1415
rect 1150 -1416 1151 -1415
rect 1157 -1416 1158 -1415
rect 1192 -1416 1193 -1415
rect 1213 -1416 1214 -1415
rect 1262 -1416 1263 -1415
rect 1332 -1416 1333 -1415
rect 1535 -1416 1536 -1415
rect 37 -1418 38 -1417
rect 191 -1418 192 -1417
rect 240 -1418 241 -1417
rect 324 -1418 325 -1417
rect 380 -1418 381 -1417
rect 513 -1418 514 -1417
rect 562 -1418 563 -1417
rect 681 -1418 682 -1417
rect 730 -1418 731 -1417
rect 926 -1418 927 -1417
rect 933 -1418 934 -1417
rect 1290 -1418 1291 -1417
rect 1318 -1418 1319 -1417
rect 1535 -1418 1536 -1417
rect 86 -1420 87 -1419
rect 730 -1420 731 -1419
rect 922 -1420 923 -1419
rect 1234 -1420 1235 -1419
rect 1248 -1420 1249 -1419
rect 1276 -1420 1277 -1419
rect 1318 -1420 1319 -1419
rect 1416 -1420 1417 -1419
rect 1430 -1420 1431 -1419
rect 1451 -1420 1452 -1419
rect 1479 -1420 1480 -1419
rect 1570 -1420 1571 -1419
rect 86 -1422 87 -1421
rect 793 -1422 794 -1421
rect 950 -1422 951 -1421
rect 1451 -1422 1452 -1421
rect 1479 -1422 1480 -1421
rect 1654 -1422 1655 -1421
rect 254 -1424 255 -1423
rect 303 -1424 304 -1423
rect 387 -1424 388 -1423
rect 814 -1424 815 -1423
rect 954 -1424 955 -1423
rect 968 -1424 969 -1423
rect 1017 -1424 1018 -1423
rect 1675 -1424 1676 -1423
rect 61 -1426 62 -1425
rect 387 -1426 388 -1425
rect 408 -1426 409 -1425
rect 765 -1426 766 -1425
rect 793 -1426 794 -1425
rect 800 -1426 801 -1425
rect 968 -1426 969 -1425
rect 1045 -1426 1046 -1425
rect 1059 -1426 1060 -1425
rect 1129 -1426 1130 -1425
rect 1192 -1426 1193 -1425
rect 1269 -1426 1270 -1425
rect 1276 -1426 1277 -1425
rect 1577 -1426 1578 -1425
rect 268 -1428 269 -1427
rect 1101 -1428 1102 -1427
rect 1129 -1428 1130 -1427
rect 1171 -1428 1172 -1427
rect 1255 -1428 1256 -1427
rect 1297 -1428 1298 -1427
rect 1416 -1428 1417 -1427
rect 1514 -1428 1515 -1427
rect 1538 -1428 1539 -1427
rect 1654 -1428 1655 -1427
rect 268 -1430 269 -1429
rect 296 -1430 297 -1429
rect 408 -1430 409 -1429
rect 604 -1430 605 -1429
rect 611 -1430 612 -1429
rect 740 -1430 741 -1429
rect 1017 -1430 1018 -1429
rect 1073 -1430 1074 -1429
rect 1080 -1430 1081 -1429
rect 1150 -1430 1151 -1429
rect 1171 -1430 1172 -1429
rect 1206 -1430 1207 -1429
rect 1262 -1430 1263 -1429
rect 1304 -1430 1305 -1429
rect 1577 -1430 1578 -1429
rect 1619 -1430 1620 -1429
rect 184 -1432 185 -1431
rect 1619 -1432 1620 -1431
rect 275 -1434 276 -1433
rect 481 -1434 482 -1433
rect 499 -1434 500 -1433
rect 800 -1434 801 -1433
rect 975 -1434 976 -1433
rect 1073 -1434 1074 -1433
rect 1143 -1434 1144 -1433
rect 1514 -1434 1515 -1433
rect 275 -1436 276 -1435
rect 828 -1436 829 -1435
rect 1020 -1436 1021 -1435
rect 1122 -1436 1123 -1435
rect 1143 -1436 1144 -1435
rect 1178 -1436 1179 -1435
rect 1297 -1436 1298 -1435
rect 1493 -1436 1494 -1435
rect 296 -1438 297 -1437
rect 464 -1438 465 -1437
rect 478 -1438 479 -1437
rect 1206 -1438 1207 -1437
rect 1304 -1438 1305 -1437
rect 1353 -1438 1354 -1437
rect 1360 -1438 1361 -1437
rect 1493 -1438 1494 -1437
rect 44 -1440 45 -1439
rect 464 -1440 465 -1439
rect 499 -1440 500 -1439
rect 534 -1440 535 -1439
rect 569 -1440 570 -1439
rect 1052 -1440 1053 -1439
rect 1178 -1440 1179 -1439
rect 1185 -1440 1186 -1439
rect 1353 -1440 1354 -1439
rect 1444 -1440 1445 -1439
rect 44 -1442 45 -1441
rect 72 -1442 73 -1441
rect 415 -1442 416 -1441
rect 572 -1442 573 -1441
rect 597 -1442 598 -1441
rect 737 -1442 738 -1441
rect 779 -1442 780 -1441
rect 1080 -1442 1081 -1441
rect 1185 -1442 1186 -1441
rect 1311 -1442 1312 -1441
rect 1360 -1442 1361 -1441
rect 1465 -1442 1466 -1441
rect 72 -1444 73 -1443
rect 226 -1444 227 -1443
rect 240 -1444 241 -1443
rect 737 -1444 738 -1443
rect 1045 -1444 1046 -1443
rect 1458 -1444 1459 -1443
rect 1465 -1444 1466 -1443
rect 1640 -1444 1641 -1443
rect 247 -1446 248 -1445
rect 415 -1446 416 -1445
rect 436 -1446 437 -1445
rect 947 -1446 948 -1445
rect 1052 -1446 1053 -1445
rect 1241 -1446 1242 -1445
rect 1444 -1446 1445 -1445
rect 1486 -1446 1487 -1445
rect 247 -1448 248 -1447
rect 338 -1448 339 -1447
rect 436 -1448 437 -1447
rect 936 -1448 937 -1447
rect 947 -1448 948 -1447
rect 1717 -1448 1718 -1447
rect 261 -1450 262 -1449
rect 338 -1450 339 -1449
rect 450 -1450 451 -1449
rect 667 -1450 668 -1449
rect 674 -1450 675 -1449
rect 1724 -1450 1725 -1449
rect 261 -1452 262 -1451
rect 331 -1452 332 -1451
rect 453 -1452 454 -1451
rect 842 -1452 843 -1451
rect 1241 -1452 1242 -1451
rect 1283 -1452 1284 -1451
rect 1458 -1452 1459 -1451
rect 1542 -1452 1543 -1451
rect 1710 -1452 1711 -1451
rect 1717 -1452 1718 -1451
rect 233 -1454 234 -1453
rect 842 -1454 843 -1453
rect 1283 -1454 1284 -1453
rect 1367 -1454 1368 -1453
rect 1486 -1454 1487 -1453
rect 1521 -1454 1522 -1453
rect 1542 -1454 1543 -1453
rect 1549 -1454 1550 -1453
rect 1643 -1454 1644 -1453
rect 1710 -1454 1711 -1453
rect 233 -1456 234 -1455
rect 422 -1456 423 -1455
rect 457 -1456 458 -1455
rect 905 -1456 906 -1455
rect 1367 -1456 1368 -1455
rect 1423 -1456 1424 -1455
rect 1549 -1456 1550 -1455
rect 1752 -1456 1753 -1455
rect 331 -1458 332 -1457
rect 548 -1458 549 -1457
rect 569 -1458 570 -1457
rect 590 -1458 591 -1457
rect 604 -1458 605 -1457
rect 870 -1458 871 -1457
rect 1388 -1458 1389 -1457
rect 1423 -1458 1424 -1457
rect 422 -1460 423 -1459
rect 936 -1460 937 -1459
rect 460 -1462 461 -1461
rect 1234 -1462 1235 -1461
rect 513 -1464 514 -1463
rect 1269 -1464 1270 -1463
rect 527 -1466 528 -1465
rect 597 -1466 598 -1465
rect 653 -1466 654 -1465
rect 674 -1466 675 -1465
rect 681 -1466 682 -1465
rect 807 -1466 808 -1465
rect 852 -1466 853 -1465
rect 1521 -1466 1522 -1465
rect 373 -1468 374 -1467
rect 527 -1468 528 -1467
rect 534 -1468 535 -1467
rect 824 -1468 825 -1467
rect 870 -1468 871 -1467
rect 877 -1468 878 -1467
rect 373 -1470 374 -1469
rect 492 -1470 493 -1469
rect 548 -1470 549 -1469
rect 950 -1470 951 -1469
rect 30 -1472 31 -1471
rect 492 -1472 493 -1471
rect 576 -1472 577 -1471
rect 779 -1472 780 -1471
rect 877 -1472 878 -1471
rect 884 -1472 885 -1471
rect 30 -1474 31 -1473
rect 131 -1474 132 -1473
rect 576 -1474 577 -1473
rect 632 -1474 633 -1473
rect 653 -1474 654 -1473
rect 1087 -1474 1088 -1473
rect 131 -1476 132 -1475
rect 583 -1476 584 -1475
rect 590 -1476 591 -1475
rect 985 -1476 986 -1475
rect 394 -1478 395 -1477
rect 583 -1478 584 -1477
rect 632 -1478 633 -1477
rect 989 -1478 990 -1477
rect 394 -1480 395 -1479
rect 429 -1480 430 -1479
rect 443 -1480 444 -1479
rect 1087 -1480 1088 -1479
rect 359 -1482 360 -1481
rect 429 -1482 430 -1481
rect 443 -1482 444 -1481
rect 702 -1482 703 -1481
rect 726 -1482 727 -1481
rect 1122 -1482 1123 -1481
rect 352 -1484 353 -1483
rect 359 -1484 360 -1483
rect 695 -1484 696 -1483
rect 1101 -1484 1102 -1483
rect 352 -1486 353 -1485
rect 401 -1486 402 -1485
rect 695 -1486 696 -1485
rect 723 -1486 724 -1485
rect 740 -1486 741 -1485
rect 1388 -1486 1389 -1485
rect 345 -1488 346 -1487
rect 401 -1488 402 -1487
rect 702 -1488 703 -1487
rect 828 -1488 829 -1487
rect 884 -1488 885 -1487
rect 898 -1488 899 -1487
rect 912 -1488 913 -1487
rect 989 -1488 990 -1487
rect 23 -1490 24 -1489
rect 345 -1490 346 -1489
rect 754 -1490 755 -1489
rect 807 -1490 808 -1489
rect 856 -1490 857 -1489
rect 898 -1490 899 -1489
rect 912 -1490 913 -1489
rect 961 -1490 962 -1489
rect 23 -1492 24 -1491
rect 128 -1492 129 -1491
rect 856 -1492 857 -1491
rect 863 -1492 864 -1491
rect 961 -1492 962 -1491
rect 1552 -1492 1553 -1491
rect 128 -1494 129 -1493
rect 1311 -1494 1312 -1493
rect 772 -1496 773 -1495
rect 863 -1496 864 -1495
rect 709 -1498 710 -1497
rect 772 -1498 773 -1497
rect 709 -1500 710 -1499
rect 866 -1500 867 -1499
rect 23 -1511 24 -1510
rect 229 -1511 230 -1510
rect 240 -1511 241 -1510
rect 320 -1511 321 -1510
rect 373 -1511 374 -1510
rect 376 -1511 377 -1510
rect 401 -1511 402 -1510
rect 457 -1511 458 -1510
rect 460 -1511 461 -1510
rect 1227 -1511 1228 -1510
rect 1451 -1511 1452 -1510
rect 1454 -1511 1455 -1510
rect 1521 -1511 1522 -1510
rect 1549 -1511 1550 -1510
rect 1584 -1511 1585 -1510
rect 1668 -1511 1669 -1510
rect 1706 -1511 1707 -1510
rect 1710 -1511 1711 -1510
rect 1801 -1511 1802 -1510
rect 1822 -1511 1823 -1510
rect 23 -1513 24 -1512
rect 418 -1513 419 -1512
rect 436 -1513 437 -1512
rect 761 -1513 762 -1512
rect 779 -1513 780 -1512
rect 828 -1513 829 -1512
rect 866 -1513 867 -1512
rect 1423 -1513 1424 -1512
rect 1451 -1513 1452 -1512
rect 1472 -1513 1473 -1512
rect 1521 -1513 1522 -1512
rect 1605 -1513 1606 -1512
rect 1640 -1513 1641 -1512
rect 1731 -1513 1732 -1512
rect 37 -1515 38 -1514
rect 726 -1515 727 -1514
rect 737 -1515 738 -1514
rect 1220 -1515 1221 -1514
rect 1227 -1515 1228 -1514
rect 1255 -1515 1256 -1514
rect 1304 -1515 1305 -1514
rect 1423 -1515 1424 -1514
rect 1535 -1515 1536 -1514
rect 1696 -1515 1697 -1514
rect 37 -1517 38 -1516
rect 65 -1517 66 -1516
rect 93 -1517 94 -1516
rect 317 -1517 318 -1516
rect 373 -1517 374 -1516
rect 485 -1517 486 -1516
rect 492 -1517 493 -1516
rect 670 -1517 671 -1516
rect 681 -1517 682 -1516
rect 978 -1517 979 -1516
rect 1020 -1517 1021 -1516
rect 1465 -1517 1466 -1516
rect 1535 -1517 1536 -1516
rect 1542 -1517 1543 -1516
rect 1577 -1517 1578 -1516
rect 1584 -1517 1585 -1516
rect 1598 -1517 1599 -1516
rect 1696 -1517 1697 -1516
rect 51 -1519 52 -1518
rect 625 -1519 626 -1518
rect 688 -1519 689 -1518
rect 950 -1519 951 -1518
rect 1031 -1519 1032 -1518
rect 1199 -1519 1200 -1518
rect 1255 -1519 1256 -1518
rect 1262 -1519 1263 -1518
rect 1454 -1519 1455 -1518
rect 1472 -1519 1473 -1518
rect 1507 -1519 1508 -1518
rect 1542 -1519 1543 -1518
rect 1577 -1519 1578 -1518
rect 1612 -1519 1613 -1518
rect 1640 -1519 1641 -1518
rect 1647 -1519 1648 -1518
rect 1650 -1519 1651 -1518
rect 1724 -1519 1725 -1518
rect 51 -1521 52 -1520
rect 261 -1521 262 -1520
rect 264 -1521 265 -1520
rect 520 -1521 521 -1520
rect 527 -1521 528 -1520
rect 656 -1521 657 -1520
rect 716 -1521 717 -1520
rect 1262 -1521 1263 -1520
rect 1311 -1521 1312 -1520
rect 1507 -1521 1508 -1520
rect 1591 -1521 1592 -1520
rect 1598 -1521 1599 -1520
rect 1612 -1521 1613 -1520
rect 1626 -1521 1627 -1520
rect 1643 -1521 1644 -1520
rect 1710 -1521 1711 -1520
rect 1717 -1521 1718 -1520
rect 1724 -1521 1725 -1520
rect 58 -1523 59 -1522
rect 957 -1523 958 -1522
rect 989 -1523 990 -1522
rect 1031 -1523 1032 -1522
rect 1034 -1523 1035 -1522
rect 1108 -1523 1109 -1522
rect 1157 -1523 1158 -1522
rect 1199 -1523 1200 -1522
rect 1311 -1523 1312 -1522
rect 1318 -1523 1319 -1522
rect 1479 -1523 1480 -1522
rect 1591 -1523 1592 -1522
rect 1668 -1523 1669 -1522
rect 1682 -1523 1683 -1522
rect 1703 -1523 1704 -1522
rect 1717 -1523 1718 -1522
rect 65 -1525 66 -1524
rect 870 -1525 871 -1524
rect 880 -1525 881 -1524
rect 1017 -1525 1018 -1524
rect 1045 -1525 1046 -1524
rect 1066 -1525 1067 -1524
rect 1188 -1525 1189 -1524
rect 1458 -1525 1459 -1524
rect 1514 -1525 1515 -1524
rect 1626 -1525 1627 -1524
rect 1633 -1525 1634 -1524
rect 1682 -1525 1683 -1524
rect 93 -1527 94 -1526
rect 541 -1527 542 -1526
rect 607 -1527 608 -1526
rect 919 -1527 920 -1526
rect 936 -1527 937 -1526
rect 1185 -1527 1186 -1526
rect 1192 -1527 1193 -1526
rect 1220 -1527 1221 -1526
rect 1318 -1527 1319 -1526
rect 1647 -1527 1648 -1526
rect 124 -1529 125 -1528
rect 313 -1529 314 -1528
rect 380 -1529 381 -1528
rect 457 -1529 458 -1528
rect 481 -1529 482 -1528
rect 1608 -1529 1609 -1528
rect 44 -1531 45 -1530
rect 124 -1531 125 -1530
rect 128 -1531 129 -1530
rect 198 -1531 199 -1530
rect 212 -1531 213 -1530
rect 240 -1531 241 -1530
rect 310 -1531 311 -1530
rect 726 -1531 727 -1530
rect 737 -1531 738 -1530
rect 744 -1531 745 -1530
rect 747 -1531 748 -1530
rect 933 -1531 934 -1530
rect 947 -1531 948 -1530
rect 1234 -1531 1235 -1530
rect 1332 -1531 1333 -1530
rect 1514 -1531 1515 -1530
rect 1563 -1531 1564 -1530
rect 1633 -1531 1634 -1530
rect 44 -1533 45 -1532
rect 61 -1533 62 -1532
rect 79 -1533 80 -1532
rect 128 -1533 129 -1532
rect 131 -1533 132 -1532
rect 296 -1533 297 -1532
rect 415 -1533 416 -1532
rect 569 -1533 570 -1532
rect 611 -1533 612 -1532
rect 681 -1533 682 -1532
rect 702 -1533 703 -1532
rect 716 -1533 717 -1532
rect 723 -1533 724 -1532
rect 1360 -1533 1361 -1532
rect 1416 -1533 1417 -1532
rect 1479 -1533 1480 -1532
rect 1556 -1533 1557 -1532
rect 1563 -1533 1564 -1532
rect 79 -1535 80 -1534
rect 1006 -1535 1007 -1534
rect 1048 -1535 1049 -1534
rect 1283 -1535 1284 -1534
rect 1325 -1535 1326 -1534
rect 1332 -1535 1333 -1534
rect 1395 -1535 1396 -1534
rect 1416 -1535 1417 -1534
rect 1430 -1535 1431 -1534
rect 1458 -1535 1459 -1534
rect 1556 -1535 1557 -1534
rect 1570 -1535 1571 -1534
rect 149 -1537 150 -1536
rect 611 -1537 612 -1536
rect 625 -1537 626 -1536
rect 821 -1537 822 -1536
rect 831 -1537 832 -1536
rect 1605 -1537 1606 -1536
rect 135 -1539 136 -1538
rect 149 -1539 150 -1538
rect 156 -1539 157 -1538
rect 1549 -1539 1550 -1538
rect 159 -1541 160 -1540
rect 380 -1541 381 -1540
rect 415 -1541 416 -1540
rect 471 -1541 472 -1540
rect 506 -1541 507 -1540
rect 527 -1541 528 -1540
rect 569 -1541 570 -1540
rect 1654 -1541 1655 -1540
rect 184 -1543 185 -1542
rect 443 -1543 444 -1542
rect 506 -1543 507 -1542
rect 555 -1543 556 -1542
rect 604 -1543 605 -1542
rect 702 -1543 703 -1542
rect 709 -1543 710 -1542
rect 1066 -1543 1067 -1542
rect 1073 -1543 1074 -1542
rect 1192 -1543 1193 -1542
rect 1206 -1543 1207 -1542
rect 1283 -1543 1284 -1542
rect 1290 -1543 1291 -1542
rect 1325 -1543 1326 -1542
rect 1381 -1543 1382 -1542
rect 1395 -1543 1396 -1542
rect 1493 -1543 1494 -1542
rect 1570 -1543 1571 -1542
rect 1654 -1543 1655 -1542
rect 1661 -1543 1662 -1542
rect 184 -1545 185 -1544
rect 1430 -1545 1431 -1544
rect 1661 -1545 1662 -1544
rect 1675 -1545 1676 -1544
rect 191 -1547 192 -1546
rect 401 -1547 402 -1546
rect 422 -1547 423 -1546
rect 520 -1547 521 -1546
rect 544 -1547 545 -1546
rect 1381 -1547 1382 -1546
rect 1675 -1547 1676 -1546
rect 1689 -1547 1690 -1546
rect 86 -1549 87 -1548
rect 422 -1549 423 -1548
rect 436 -1549 437 -1548
rect 996 -1549 997 -1548
rect 1059 -1549 1060 -1548
rect 1073 -1549 1074 -1548
rect 1164 -1549 1165 -1548
rect 1234 -1549 1235 -1548
rect 1269 -1549 1270 -1548
rect 1290 -1549 1291 -1548
rect 1685 -1549 1686 -1548
rect 1689 -1549 1690 -1548
rect 68 -1551 69 -1550
rect 86 -1551 87 -1550
rect 191 -1551 192 -1550
rect 247 -1551 248 -1550
rect 387 -1551 388 -1550
rect 471 -1551 472 -1550
rect 478 -1551 479 -1550
rect 1493 -1551 1494 -1550
rect 194 -1553 195 -1552
rect 1465 -1553 1466 -1552
rect 198 -1555 199 -1554
rect 450 -1555 451 -1554
rect 653 -1555 654 -1554
rect 919 -1555 920 -1554
rect 947 -1555 948 -1554
rect 1538 -1555 1539 -1554
rect 205 -1557 206 -1556
rect 933 -1557 934 -1556
rect 968 -1557 969 -1556
rect 989 -1557 990 -1556
rect 996 -1557 997 -1556
rect 1122 -1557 1123 -1556
rect 1178 -1557 1179 -1556
rect 1269 -1557 1270 -1556
rect 121 -1559 122 -1558
rect 205 -1559 206 -1558
rect 212 -1559 213 -1558
rect 324 -1559 325 -1558
rect 387 -1559 388 -1558
rect 464 -1559 465 -1558
rect 541 -1559 542 -1558
rect 1122 -1559 1123 -1558
rect 1136 -1559 1137 -1558
rect 1178 -1559 1179 -1558
rect 1185 -1559 1186 -1558
rect 1304 -1559 1305 -1558
rect 121 -1561 122 -1560
rect 156 -1561 157 -1560
rect 215 -1561 216 -1560
rect 408 -1561 409 -1560
rect 443 -1561 444 -1560
rect 562 -1561 563 -1560
rect 632 -1561 633 -1560
rect 968 -1561 969 -1560
rect 1062 -1561 1063 -1560
rect 1444 -1561 1445 -1560
rect 219 -1563 220 -1562
rect 688 -1563 689 -1562
rect 709 -1563 710 -1562
rect 835 -1563 836 -1562
rect 863 -1563 864 -1562
rect 1360 -1563 1361 -1562
rect 1367 -1563 1368 -1562
rect 1444 -1563 1445 -1562
rect 30 -1565 31 -1564
rect 219 -1565 220 -1564
rect 222 -1565 223 -1564
rect 733 -1565 734 -1564
rect 740 -1565 741 -1564
rect 1101 -1565 1102 -1564
rect 1136 -1565 1137 -1564
rect 1143 -1565 1144 -1564
rect 1346 -1565 1347 -1564
rect 1367 -1565 1368 -1564
rect 30 -1567 31 -1566
rect 628 -1567 629 -1566
rect 653 -1567 654 -1566
rect 674 -1567 675 -1566
rect 754 -1567 755 -1566
rect 1052 -1567 1053 -1566
rect 1101 -1567 1102 -1566
rect 1150 -1567 1151 -1566
rect 1346 -1567 1347 -1566
rect 1402 -1567 1403 -1566
rect 233 -1569 234 -1568
rect 296 -1569 297 -1568
rect 324 -1569 325 -1568
rect 817 -1569 818 -1568
rect 863 -1569 864 -1568
rect 1157 -1569 1158 -1568
rect 1388 -1569 1389 -1568
rect 1402 -1569 1403 -1568
rect 233 -1571 234 -1570
rect 429 -1571 430 -1570
rect 446 -1571 447 -1570
rect 478 -1571 479 -1570
rect 499 -1571 500 -1570
rect 632 -1571 633 -1570
rect 667 -1571 668 -1570
rect 1164 -1571 1165 -1570
rect 1388 -1571 1389 -1570
rect 1500 -1571 1501 -1570
rect 247 -1573 248 -1572
rect 310 -1573 311 -1572
rect 429 -1573 430 -1572
rect 821 -1573 822 -1572
rect 870 -1573 871 -1572
rect 1003 -1573 1004 -1572
rect 1094 -1573 1095 -1572
rect 1150 -1573 1151 -1572
rect 1409 -1573 1410 -1572
rect 1500 -1573 1501 -1572
rect 275 -1575 276 -1574
rect 408 -1575 409 -1574
rect 464 -1575 465 -1574
rect 604 -1575 605 -1574
rect 758 -1575 759 -1574
rect 856 -1575 857 -1574
rect 894 -1575 895 -1574
rect 1241 -1575 1242 -1574
rect 1353 -1575 1354 -1574
rect 1409 -1575 1410 -1574
rect 142 -1577 143 -1576
rect 275 -1577 276 -1576
rect 499 -1577 500 -1576
rect 639 -1577 640 -1576
rect 730 -1577 731 -1576
rect 758 -1577 759 -1576
rect 779 -1577 780 -1576
rect 1017 -1577 1018 -1576
rect 1094 -1577 1095 -1576
rect 1129 -1577 1130 -1576
rect 1297 -1577 1298 -1576
rect 1353 -1577 1354 -1576
rect 142 -1579 143 -1578
rect 163 -1579 164 -1578
rect 548 -1579 549 -1578
rect 667 -1579 668 -1578
rect 730 -1579 731 -1578
rect 1339 -1579 1340 -1578
rect 163 -1581 164 -1580
rect 1241 -1581 1242 -1580
rect 1297 -1581 1298 -1580
rect 1339 -1581 1340 -1580
rect 548 -1583 549 -1582
rect 583 -1583 584 -1582
rect 590 -1583 591 -1582
rect 674 -1583 675 -1582
rect 786 -1583 787 -1582
rect 926 -1583 927 -1582
rect 940 -1583 941 -1582
rect 1003 -1583 1004 -1582
rect 1115 -1583 1116 -1582
rect 1129 -1583 1130 -1582
rect 187 -1585 188 -1584
rect 590 -1585 591 -1584
rect 639 -1585 640 -1584
rect 891 -1585 892 -1584
rect 912 -1585 913 -1584
rect 926 -1585 927 -1584
rect 940 -1585 941 -1584
rect 1080 -1585 1081 -1584
rect 1087 -1585 1088 -1584
rect 1115 -1585 1116 -1584
rect 1125 -1585 1126 -1584
rect 1143 -1585 1144 -1584
rect 492 -1587 493 -1586
rect 891 -1587 892 -1586
rect 898 -1587 899 -1586
rect 912 -1587 913 -1586
rect 975 -1587 976 -1586
rect 1052 -1587 1053 -1586
rect 1080 -1587 1081 -1586
rect 1206 -1587 1207 -1586
rect 562 -1589 563 -1588
rect 576 -1589 577 -1588
rect 583 -1589 584 -1588
rect 660 -1589 661 -1588
rect 786 -1589 787 -1588
rect 824 -1589 825 -1588
rect 884 -1589 885 -1588
rect 898 -1589 899 -1588
rect 954 -1589 955 -1588
rect 975 -1589 976 -1588
rect 1024 -1589 1025 -1588
rect 1087 -1589 1088 -1588
rect 135 -1591 136 -1590
rect 824 -1591 825 -1590
rect 849 -1591 850 -1590
rect 884 -1591 885 -1590
rect 954 -1591 955 -1590
rect 1276 -1591 1277 -1590
rect 450 -1593 451 -1592
rect 849 -1593 850 -1592
rect 1010 -1593 1011 -1592
rect 1024 -1593 1025 -1592
rect 1213 -1593 1214 -1592
rect 1276 -1593 1277 -1592
rect 551 -1595 552 -1594
rect 1213 -1595 1214 -1594
rect 576 -1597 577 -1596
rect 765 -1597 766 -1596
rect 789 -1597 790 -1596
rect 842 -1597 843 -1596
rect 982 -1597 983 -1596
rect 1010 -1597 1011 -1596
rect 597 -1599 598 -1598
rect 660 -1599 661 -1598
rect 800 -1599 801 -1598
rect 835 -1599 836 -1598
rect 982 -1599 983 -1598
rect 1038 -1599 1039 -1598
rect 72 -1601 73 -1600
rect 1038 -1601 1039 -1600
rect 72 -1603 73 -1602
rect 254 -1603 255 -1602
rect 618 -1603 619 -1602
rect 765 -1603 766 -1602
rect 793 -1603 794 -1602
rect 800 -1603 801 -1602
rect 807 -1603 808 -1602
rect 866 -1603 867 -1602
rect 100 -1605 101 -1604
rect 618 -1605 619 -1604
rect 772 -1605 773 -1604
rect 793 -1605 794 -1604
rect 814 -1605 815 -1604
rect 842 -1605 843 -1604
rect 100 -1607 101 -1606
rect 226 -1607 227 -1606
rect 513 -1607 514 -1606
rect 807 -1607 808 -1606
rect 114 -1609 115 -1608
rect 226 -1609 227 -1608
rect 359 -1609 360 -1608
rect 513 -1609 514 -1608
rect 555 -1609 556 -1608
rect 814 -1609 815 -1608
rect 114 -1611 115 -1610
rect 331 -1611 332 -1610
rect 359 -1611 360 -1610
rect 366 -1611 367 -1610
rect 751 -1611 752 -1610
rect 772 -1611 773 -1610
rect 166 -1613 167 -1612
rect 254 -1613 255 -1612
rect 366 -1613 367 -1612
rect 751 -1613 752 -1612
rect 170 -1615 171 -1614
rect 597 -1615 598 -1614
rect 170 -1617 171 -1616
rect 289 -1617 290 -1616
rect 107 -1619 108 -1618
rect 289 -1619 290 -1618
rect 107 -1621 108 -1620
rect 394 -1621 395 -1620
rect 268 -1623 269 -1622
rect 394 -1623 395 -1622
rect 268 -1625 269 -1624
rect 282 -1625 283 -1624
rect 282 -1627 283 -1626
rect 338 -1627 339 -1626
rect 338 -1629 339 -1628
rect 345 -1629 346 -1628
rect 345 -1631 346 -1630
rect 534 -1631 535 -1630
rect 534 -1633 535 -1632
rect 877 -1633 878 -1632
rect 331 -1635 332 -1634
rect 877 -1635 878 -1634
rect 30 -1646 31 -1645
rect 310 -1646 311 -1645
rect 324 -1646 325 -1645
rect 383 -1646 384 -1645
rect 387 -1646 388 -1645
rect 607 -1646 608 -1645
rect 660 -1646 661 -1645
rect 733 -1646 734 -1645
rect 789 -1646 790 -1645
rect 1297 -1646 1298 -1645
rect 1300 -1646 1301 -1645
rect 1458 -1646 1459 -1645
rect 1549 -1646 1550 -1645
rect 1703 -1646 1704 -1645
rect 1822 -1646 1823 -1645
rect 1839 -1646 1840 -1645
rect 30 -1648 31 -1647
rect 198 -1648 199 -1647
rect 219 -1648 220 -1647
rect 502 -1648 503 -1647
rect 548 -1648 549 -1647
rect 1710 -1648 1711 -1647
rect 23 -1650 24 -1649
rect 198 -1650 199 -1649
rect 236 -1650 237 -1649
rect 1794 -1650 1795 -1649
rect 23 -1652 24 -1651
rect 233 -1652 234 -1651
rect 275 -1652 276 -1651
rect 310 -1652 311 -1651
rect 352 -1652 353 -1651
rect 450 -1652 451 -1651
rect 551 -1652 552 -1651
rect 1115 -1652 1116 -1651
rect 1122 -1652 1123 -1651
rect 1458 -1652 1459 -1651
rect 1598 -1652 1599 -1651
rect 1731 -1652 1732 -1651
rect 58 -1654 59 -1653
rect 730 -1654 731 -1653
rect 800 -1654 801 -1653
rect 817 -1654 818 -1653
rect 856 -1654 857 -1653
rect 884 -1654 885 -1653
rect 891 -1654 892 -1653
rect 1787 -1654 1788 -1653
rect 107 -1656 108 -1655
rect 891 -1656 892 -1655
rect 954 -1656 955 -1655
rect 1111 -1656 1112 -1655
rect 1125 -1656 1126 -1655
rect 1255 -1656 1256 -1655
rect 1423 -1656 1424 -1655
rect 1549 -1656 1550 -1655
rect 1605 -1656 1606 -1655
rect 1745 -1656 1746 -1655
rect 93 -1658 94 -1657
rect 107 -1658 108 -1657
rect 121 -1658 122 -1657
rect 1171 -1658 1172 -1657
rect 1185 -1658 1186 -1657
rect 1836 -1658 1837 -1657
rect 93 -1660 94 -1659
rect 537 -1660 538 -1659
rect 576 -1660 577 -1659
rect 800 -1660 801 -1659
rect 814 -1660 815 -1659
rect 1640 -1660 1641 -1659
rect 1647 -1660 1648 -1659
rect 1780 -1660 1781 -1659
rect 121 -1662 122 -1661
rect 719 -1662 720 -1661
rect 782 -1662 783 -1661
rect 1605 -1662 1606 -1661
rect 1619 -1662 1620 -1661
rect 1752 -1662 1753 -1661
rect 124 -1664 125 -1663
rect 887 -1664 888 -1663
rect 957 -1664 958 -1663
rect 1738 -1664 1739 -1663
rect 135 -1666 136 -1665
rect 677 -1666 678 -1665
rect 681 -1666 682 -1665
rect 751 -1666 752 -1665
rect 835 -1666 836 -1665
rect 1171 -1666 1172 -1665
rect 1185 -1666 1186 -1665
rect 1234 -1666 1235 -1665
rect 1304 -1666 1305 -1665
rect 1423 -1666 1424 -1665
rect 1451 -1666 1452 -1665
rect 1710 -1666 1711 -1665
rect 135 -1668 136 -1667
rect 1062 -1668 1063 -1667
rect 1066 -1668 1067 -1667
rect 1083 -1668 1084 -1667
rect 1101 -1668 1102 -1667
rect 1255 -1668 1256 -1667
rect 1332 -1668 1333 -1667
rect 1451 -1668 1452 -1667
rect 1479 -1668 1480 -1667
rect 1619 -1668 1620 -1667
rect 1626 -1668 1627 -1667
rect 1759 -1668 1760 -1667
rect 159 -1670 160 -1669
rect 579 -1670 580 -1669
rect 590 -1670 591 -1669
rect 751 -1670 752 -1669
rect 835 -1670 836 -1669
rect 849 -1670 850 -1669
rect 859 -1670 860 -1669
rect 996 -1670 997 -1669
rect 1003 -1670 1004 -1669
rect 1563 -1670 1564 -1669
rect 1633 -1670 1634 -1669
rect 1766 -1670 1767 -1669
rect 184 -1672 185 -1671
rect 212 -1672 213 -1671
rect 275 -1672 276 -1671
rect 520 -1672 521 -1671
rect 604 -1672 605 -1671
rect 726 -1672 727 -1671
rect 863 -1672 864 -1671
rect 1087 -1672 1088 -1671
rect 1101 -1672 1102 -1671
rect 1689 -1672 1690 -1671
rect 1696 -1672 1697 -1671
rect 1829 -1672 1830 -1671
rect 145 -1674 146 -1673
rect 184 -1674 185 -1673
rect 187 -1674 188 -1673
rect 534 -1674 535 -1673
rect 611 -1674 612 -1673
rect 660 -1674 661 -1673
rect 674 -1674 675 -1673
rect 814 -1674 815 -1673
rect 828 -1674 829 -1673
rect 863 -1674 864 -1673
rect 877 -1674 878 -1673
rect 1360 -1674 1361 -1673
rect 1374 -1674 1375 -1673
rect 1479 -1674 1480 -1673
rect 1521 -1674 1522 -1673
rect 1640 -1674 1641 -1673
rect 1650 -1674 1651 -1673
rect 1724 -1674 1725 -1673
rect 44 -1676 45 -1675
rect 674 -1676 675 -1675
rect 681 -1676 682 -1675
rect 779 -1676 780 -1675
rect 786 -1676 787 -1675
rect 828 -1676 829 -1675
rect 877 -1676 878 -1675
rect 905 -1676 906 -1675
rect 950 -1676 951 -1675
rect 1633 -1676 1634 -1675
rect 1654 -1676 1655 -1675
rect 1808 -1676 1809 -1675
rect 44 -1678 45 -1677
rect 639 -1678 640 -1677
rect 716 -1678 717 -1677
rect 730 -1678 731 -1677
rect 779 -1678 780 -1677
rect 824 -1678 825 -1677
rect 880 -1678 881 -1677
rect 1325 -1678 1326 -1677
rect 1395 -1678 1396 -1677
rect 1521 -1678 1522 -1677
rect 1528 -1678 1529 -1677
rect 1689 -1678 1690 -1677
rect 212 -1680 213 -1679
rect 555 -1680 556 -1679
rect 611 -1680 612 -1679
rect 842 -1680 843 -1679
rect 901 -1680 902 -1679
rect 996 -1680 997 -1679
rect 1017 -1680 1018 -1679
rect 1129 -1680 1130 -1679
rect 1146 -1680 1147 -1679
rect 1577 -1680 1578 -1679
rect 1584 -1680 1585 -1679
rect 1724 -1680 1725 -1679
rect 303 -1682 304 -1681
rect 324 -1682 325 -1681
rect 352 -1682 353 -1681
rect 544 -1682 545 -1681
rect 618 -1682 619 -1681
rect 905 -1682 906 -1681
rect 947 -1682 948 -1681
rect 1017 -1682 1018 -1681
rect 1020 -1682 1021 -1681
rect 1234 -1682 1235 -1681
rect 1262 -1682 1263 -1681
rect 1325 -1682 1326 -1681
rect 1402 -1682 1403 -1681
rect 1528 -1682 1529 -1681
rect 1542 -1682 1543 -1681
rect 1696 -1682 1697 -1681
rect 205 -1684 206 -1683
rect 1402 -1684 1403 -1683
rect 1416 -1684 1417 -1683
rect 1542 -1684 1543 -1683
rect 1661 -1684 1662 -1683
rect 1801 -1684 1802 -1683
rect 37 -1686 38 -1685
rect 1661 -1686 1662 -1685
rect 1668 -1686 1669 -1685
rect 1815 -1686 1816 -1685
rect 37 -1688 38 -1687
rect 506 -1688 507 -1687
rect 534 -1688 535 -1687
rect 1087 -1688 1088 -1687
rect 1108 -1688 1109 -1687
rect 1591 -1688 1592 -1687
rect 1675 -1688 1676 -1687
rect 1822 -1688 1823 -1687
rect 79 -1690 80 -1689
rect 205 -1690 206 -1689
rect 254 -1690 255 -1689
rect 303 -1690 304 -1689
rect 331 -1690 332 -1689
rect 618 -1690 619 -1689
rect 639 -1690 640 -1689
rect 646 -1690 647 -1689
rect 716 -1690 717 -1689
rect 1031 -1690 1032 -1689
rect 1038 -1690 1039 -1689
rect 1598 -1690 1599 -1689
rect 1682 -1690 1683 -1689
rect 1717 -1690 1718 -1689
rect 79 -1692 80 -1691
rect 366 -1692 367 -1691
rect 387 -1692 388 -1691
rect 492 -1692 493 -1691
rect 499 -1692 500 -1691
rect 520 -1692 521 -1691
rect 646 -1692 647 -1691
rect 653 -1692 654 -1691
rect 723 -1692 724 -1691
rect 1066 -1692 1067 -1691
rect 1080 -1692 1081 -1691
rect 1416 -1692 1417 -1691
rect 1437 -1692 1438 -1691
rect 1563 -1692 1564 -1691
rect 1570 -1692 1571 -1691
rect 1591 -1692 1592 -1691
rect 254 -1694 255 -1693
rect 464 -1694 465 -1693
rect 485 -1694 486 -1693
rect 544 -1694 545 -1693
rect 632 -1694 633 -1693
rect 653 -1694 654 -1693
rect 747 -1694 748 -1693
rect 1395 -1694 1396 -1693
rect 1444 -1694 1445 -1693
rect 1584 -1694 1585 -1693
rect 331 -1696 332 -1695
rect 359 -1696 360 -1695
rect 362 -1696 363 -1695
rect 1003 -1696 1004 -1695
rect 1010 -1696 1011 -1695
rect 1080 -1696 1081 -1695
rect 1129 -1696 1130 -1695
rect 1248 -1696 1249 -1695
rect 1269 -1696 1270 -1695
rect 1332 -1696 1333 -1695
rect 1388 -1696 1389 -1695
rect 1675 -1696 1676 -1695
rect 366 -1698 367 -1697
rect 380 -1698 381 -1697
rect 394 -1698 395 -1697
rect 593 -1698 594 -1697
rect 807 -1698 808 -1697
rect 842 -1698 843 -1697
rect 975 -1698 976 -1697
rect 1031 -1698 1032 -1697
rect 1038 -1698 1039 -1697
rect 1059 -1698 1060 -1697
rect 1136 -1698 1137 -1697
rect 1269 -1698 1270 -1697
rect 1290 -1698 1291 -1697
rect 1388 -1698 1389 -1697
rect 1472 -1698 1473 -1697
rect 1626 -1698 1627 -1697
rect 394 -1700 395 -1699
rect 597 -1700 598 -1699
rect 754 -1700 755 -1699
rect 1136 -1700 1137 -1699
rect 1157 -1700 1158 -1699
rect 1444 -1700 1445 -1699
rect 1493 -1700 1494 -1699
rect 1654 -1700 1655 -1699
rect 401 -1702 402 -1701
rect 597 -1702 598 -1701
rect 726 -1702 727 -1701
rect 1493 -1702 1494 -1701
rect 1500 -1702 1501 -1701
rect 1577 -1702 1578 -1701
rect 240 -1704 241 -1703
rect 401 -1704 402 -1703
rect 408 -1704 409 -1703
rect 551 -1704 552 -1703
rect 765 -1704 766 -1703
rect 807 -1704 808 -1703
rect 824 -1704 825 -1703
rect 968 -1704 969 -1703
rect 978 -1704 979 -1703
rect 1647 -1704 1648 -1703
rect 114 -1706 115 -1705
rect 240 -1706 241 -1705
rect 408 -1706 409 -1705
rect 884 -1706 885 -1705
rect 898 -1706 899 -1705
rect 968 -1706 969 -1705
rect 989 -1706 990 -1705
rect 1108 -1706 1109 -1705
rect 1157 -1706 1158 -1705
rect 1318 -1706 1319 -1705
rect 1339 -1706 1340 -1705
rect 1472 -1706 1473 -1705
rect 1507 -1706 1508 -1705
rect 1570 -1706 1571 -1705
rect 415 -1708 416 -1707
rect 450 -1708 451 -1707
rect 457 -1708 458 -1707
rect 492 -1708 493 -1707
rect 506 -1708 507 -1707
rect 541 -1708 542 -1707
rect 758 -1708 759 -1707
rect 765 -1708 766 -1707
rect 919 -1708 920 -1707
rect 989 -1708 990 -1707
rect 1010 -1708 1011 -1707
rect 1143 -1708 1144 -1707
rect 1164 -1708 1165 -1707
rect 1248 -1708 1249 -1707
rect 1276 -1708 1277 -1707
rect 1339 -1708 1340 -1707
rect 1381 -1708 1382 -1707
rect 1500 -1708 1501 -1707
rect 1514 -1708 1515 -1707
rect 1668 -1708 1669 -1707
rect 219 -1710 220 -1709
rect 1514 -1710 1515 -1709
rect 1535 -1710 1536 -1709
rect 1682 -1710 1683 -1709
rect 415 -1712 416 -1711
rect 576 -1712 577 -1711
rect 635 -1712 636 -1711
rect 1381 -1712 1382 -1711
rect 1409 -1712 1410 -1711
rect 1535 -1712 1536 -1711
rect 1556 -1712 1557 -1711
rect 1717 -1712 1718 -1711
rect 429 -1714 430 -1713
rect 1304 -1714 1305 -1713
rect 1311 -1714 1312 -1713
rect 1507 -1714 1508 -1713
rect 436 -1716 437 -1715
rect 744 -1716 745 -1715
rect 758 -1716 759 -1715
rect 772 -1716 773 -1715
rect 786 -1716 787 -1715
rect 1276 -1716 1277 -1715
rect 1430 -1716 1431 -1715
rect 1556 -1716 1557 -1715
rect 114 -1718 115 -1717
rect 772 -1718 773 -1717
rect 849 -1718 850 -1717
rect 1143 -1718 1144 -1717
rect 1178 -1718 1179 -1717
rect 1311 -1718 1312 -1717
rect 1367 -1718 1368 -1717
rect 1430 -1718 1431 -1717
rect 436 -1720 437 -1719
rect 569 -1720 570 -1719
rect 695 -1720 696 -1719
rect 744 -1720 745 -1719
rect 870 -1720 871 -1719
rect 919 -1720 920 -1719
rect 933 -1720 934 -1719
rect 1059 -1720 1060 -1719
rect 1206 -1720 1207 -1719
rect 1612 -1720 1613 -1719
rect 89 -1722 90 -1721
rect 1206 -1722 1207 -1721
rect 1220 -1722 1221 -1721
rect 1318 -1722 1319 -1721
rect 1353 -1722 1354 -1721
rect 1612 -1722 1613 -1721
rect 446 -1724 447 -1723
rect 513 -1724 514 -1723
rect 541 -1724 542 -1723
rect 555 -1724 556 -1723
rect 562 -1724 563 -1723
rect 569 -1724 570 -1723
rect 695 -1724 696 -1723
rect 793 -1724 794 -1723
rect 870 -1724 871 -1723
rect 947 -1724 948 -1723
rect 1006 -1724 1007 -1723
rect 1409 -1724 1410 -1723
rect 317 -1726 318 -1725
rect 793 -1726 794 -1725
rect 933 -1726 934 -1725
rect 961 -1726 962 -1725
rect 1024 -1726 1025 -1725
rect 1374 -1726 1375 -1725
rect 268 -1728 269 -1727
rect 1024 -1728 1025 -1727
rect 1027 -1728 1028 -1727
rect 1122 -1728 1123 -1727
rect 1227 -1728 1228 -1727
rect 1367 -1728 1368 -1727
rect 268 -1730 269 -1729
rect 548 -1730 549 -1729
rect 562 -1730 563 -1729
rect 898 -1730 899 -1729
rect 940 -1730 941 -1729
rect 1178 -1730 1179 -1729
rect 1241 -1730 1242 -1729
rect 1262 -1730 1263 -1729
rect 1283 -1730 1284 -1729
rect 1353 -1730 1354 -1729
rect 100 -1732 101 -1731
rect 1241 -1732 1242 -1731
rect 100 -1734 101 -1733
rect 170 -1734 171 -1733
rect 261 -1734 262 -1733
rect 940 -1734 941 -1733
rect 1045 -1734 1046 -1733
rect 1164 -1734 1165 -1733
rect 1213 -1734 1214 -1733
rect 1283 -1734 1284 -1733
rect 317 -1736 318 -1735
rect 1209 -1736 1210 -1735
rect 453 -1738 454 -1737
rect 1220 -1738 1221 -1737
rect 457 -1740 458 -1739
rect 478 -1740 479 -1739
rect 485 -1740 486 -1739
rect 527 -1740 528 -1739
rect 1045 -1740 1046 -1739
rect 1199 -1740 1200 -1739
rect 163 -1742 164 -1741
rect 1199 -1742 1200 -1741
rect 163 -1744 164 -1743
rect 191 -1744 192 -1743
rect 289 -1744 290 -1743
rect 527 -1744 528 -1743
rect 1052 -1744 1053 -1743
rect 1115 -1744 1116 -1743
rect 1150 -1744 1151 -1743
rect 1213 -1744 1214 -1743
rect 156 -1746 157 -1745
rect 191 -1746 192 -1745
rect 222 -1746 223 -1745
rect 289 -1746 290 -1745
rect 464 -1746 465 -1745
rect 471 -1746 472 -1745
rect 478 -1746 479 -1745
rect 583 -1746 584 -1745
rect 982 -1746 983 -1745
rect 1150 -1746 1151 -1745
rect 156 -1748 157 -1747
rect 429 -1748 430 -1747
rect 471 -1748 472 -1747
rect 625 -1748 626 -1747
rect 912 -1748 913 -1747
rect 982 -1748 983 -1747
rect 1052 -1748 1053 -1747
rect 1486 -1748 1487 -1747
rect 170 -1750 171 -1749
rect 222 -1750 223 -1749
rect 499 -1750 500 -1749
rect 961 -1750 962 -1749
rect 1055 -1750 1056 -1749
rect 1360 -1750 1361 -1749
rect 1465 -1750 1466 -1749
rect 1486 -1750 1487 -1749
rect 513 -1752 514 -1751
rect 667 -1752 668 -1751
rect 702 -1752 703 -1751
rect 912 -1752 913 -1751
rect 1094 -1752 1095 -1751
rect 1227 -1752 1228 -1751
rect 1346 -1752 1347 -1751
rect 1465 -1752 1466 -1751
rect 296 -1754 297 -1753
rect 1094 -1754 1095 -1753
rect 1192 -1754 1193 -1753
rect 1346 -1754 1347 -1753
rect 226 -1756 227 -1755
rect 296 -1756 297 -1755
rect 422 -1756 423 -1755
rect 702 -1756 703 -1755
rect 1073 -1756 1074 -1755
rect 1192 -1756 1193 -1755
rect 51 -1758 52 -1757
rect 226 -1758 227 -1757
rect 422 -1758 423 -1757
rect 737 -1758 738 -1757
rect 51 -1760 52 -1759
rect 926 -1760 927 -1759
rect 65 -1762 66 -1761
rect 926 -1762 927 -1761
rect 65 -1764 66 -1763
rect 373 -1764 374 -1763
rect 583 -1764 584 -1763
rect 1437 -1764 1438 -1763
rect 247 -1766 248 -1765
rect 373 -1766 374 -1765
rect 625 -1766 626 -1765
rect 1685 -1766 1686 -1765
rect 72 -1768 73 -1767
rect 247 -1768 248 -1767
rect 667 -1768 668 -1767
rect 705 -1768 706 -1767
rect 709 -1768 710 -1767
rect 1073 -1768 1074 -1767
rect 72 -1770 73 -1769
rect 1773 -1770 1774 -1769
rect 688 -1772 689 -1771
rect 737 -1772 738 -1771
rect 128 -1774 129 -1773
rect 688 -1774 689 -1773
rect 709 -1774 710 -1773
rect 866 -1774 867 -1773
rect 86 -1776 87 -1775
rect 128 -1776 129 -1775
rect 86 -1778 87 -1777
rect 149 -1778 150 -1777
rect 149 -1780 150 -1779
rect 177 -1780 178 -1779
rect 142 -1782 143 -1781
rect 177 -1782 178 -1781
rect 37 -1793 38 -1792
rect 537 -1793 538 -1792
rect 541 -1793 542 -1792
rect 684 -1793 685 -1792
rect 695 -1793 696 -1792
rect 915 -1793 916 -1792
rect 947 -1793 948 -1792
rect 1206 -1793 1207 -1792
rect 1230 -1793 1231 -1792
rect 1640 -1793 1641 -1792
rect 37 -1795 38 -1794
rect 611 -1795 612 -1794
rect 621 -1795 622 -1794
rect 1087 -1795 1088 -1794
rect 1143 -1795 1144 -1794
rect 1192 -1795 1193 -1794
rect 1395 -1795 1396 -1794
rect 1755 -1795 1756 -1794
rect 30 -1797 31 -1796
rect 611 -1797 612 -1796
rect 635 -1797 636 -1796
rect 646 -1797 647 -1796
rect 656 -1797 657 -1796
rect 891 -1797 892 -1796
rect 898 -1797 899 -1796
rect 1213 -1797 1214 -1796
rect 1423 -1797 1424 -1796
rect 1426 -1797 1427 -1796
rect 1640 -1797 1641 -1796
rect 1829 -1797 1830 -1796
rect 30 -1799 31 -1798
rect 93 -1799 94 -1798
rect 100 -1799 101 -1798
rect 117 -1799 118 -1798
rect 142 -1799 143 -1798
rect 1052 -1799 1053 -1798
rect 1192 -1799 1193 -1798
rect 1325 -1799 1326 -1798
rect 1423 -1799 1424 -1798
rect 1535 -1799 1536 -1798
rect 65 -1801 66 -1800
rect 264 -1801 265 -1800
rect 268 -1801 269 -1800
rect 646 -1801 647 -1800
rect 674 -1801 675 -1800
rect 695 -1801 696 -1800
rect 716 -1801 717 -1800
rect 1444 -1801 1445 -1800
rect 68 -1803 69 -1802
rect 373 -1803 374 -1802
rect 394 -1803 395 -1802
rect 502 -1803 503 -1802
rect 548 -1803 549 -1802
rect 1178 -1803 1179 -1802
rect 1213 -1803 1214 -1802
rect 1283 -1803 1284 -1802
rect 1325 -1803 1326 -1802
rect 1493 -1803 1494 -1802
rect 72 -1805 73 -1804
rect 128 -1805 129 -1804
rect 145 -1805 146 -1804
rect 359 -1805 360 -1804
rect 373 -1805 374 -1804
rect 709 -1805 710 -1804
rect 723 -1805 724 -1804
rect 992 -1805 993 -1804
rect 1024 -1805 1025 -1804
rect 1689 -1805 1690 -1804
rect 72 -1807 73 -1806
rect 457 -1807 458 -1806
rect 499 -1807 500 -1806
rect 1101 -1807 1102 -1806
rect 1178 -1807 1179 -1806
rect 1227 -1807 1228 -1806
rect 1234 -1807 1235 -1806
rect 1493 -1807 1494 -1806
rect 1689 -1807 1690 -1806
rect 1787 -1807 1788 -1806
rect 75 -1809 76 -1808
rect 814 -1809 815 -1808
rect 821 -1809 822 -1808
rect 835 -1809 836 -1808
rect 884 -1809 885 -1808
rect 1668 -1809 1669 -1808
rect 79 -1811 80 -1810
rect 82 -1811 83 -1810
rect 89 -1811 90 -1810
rect 177 -1811 178 -1810
rect 184 -1811 185 -1810
rect 236 -1811 237 -1810
rect 250 -1811 251 -1810
rect 457 -1811 458 -1810
rect 548 -1811 549 -1810
rect 597 -1811 598 -1810
rect 674 -1811 675 -1810
rect 772 -1811 773 -1810
rect 782 -1811 783 -1810
rect 1794 -1811 1795 -1810
rect 58 -1813 59 -1812
rect 177 -1813 178 -1812
rect 184 -1813 185 -1812
rect 317 -1813 318 -1812
rect 338 -1813 339 -1812
rect 432 -1813 433 -1812
rect 576 -1813 577 -1812
rect 667 -1813 668 -1812
rect 677 -1813 678 -1812
rect 1066 -1813 1067 -1812
rect 1101 -1813 1102 -1812
rect 1164 -1813 1165 -1812
rect 1283 -1813 1284 -1812
rect 1332 -1813 1333 -1812
rect 1444 -1813 1445 -1812
rect 1724 -1813 1725 -1812
rect 1794 -1813 1795 -1812
rect 1836 -1813 1837 -1812
rect 58 -1815 59 -1814
rect 1661 -1815 1662 -1814
rect 1668 -1815 1669 -1814
rect 1745 -1815 1746 -1814
rect 79 -1817 80 -1816
rect 443 -1817 444 -1816
rect 583 -1817 584 -1816
rect 625 -1817 626 -1816
rect 726 -1817 727 -1816
rect 1227 -1817 1228 -1816
rect 1332 -1817 1333 -1816
rect 1381 -1817 1382 -1816
rect 1661 -1817 1662 -1816
rect 1738 -1817 1739 -1816
rect 1745 -1817 1746 -1816
rect 1815 -1817 1816 -1816
rect 93 -1819 94 -1818
rect 478 -1819 479 -1818
rect 534 -1819 535 -1818
rect 583 -1819 584 -1818
rect 597 -1819 598 -1818
rect 772 -1819 773 -1818
rect 786 -1819 787 -1818
rect 1374 -1819 1375 -1818
rect 1381 -1819 1382 -1818
rect 1808 -1819 1809 -1818
rect 100 -1821 101 -1820
rect 415 -1821 416 -1820
rect 422 -1821 423 -1820
rect 670 -1821 671 -1820
rect 726 -1821 727 -1820
rect 1027 -1821 1028 -1820
rect 1052 -1821 1053 -1820
rect 1150 -1821 1151 -1820
rect 1374 -1821 1375 -1820
rect 1416 -1821 1417 -1820
rect 1577 -1821 1578 -1820
rect 1738 -1821 1739 -1820
rect 110 -1823 111 -1822
rect 1234 -1823 1235 -1822
rect 1416 -1823 1417 -1822
rect 1584 -1823 1585 -1822
rect 128 -1825 129 -1824
rect 149 -1825 150 -1824
rect 159 -1825 160 -1824
rect 1839 -1825 1840 -1824
rect 149 -1827 150 -1826
rect 520 -1827 521 -1826
rect 527 -1827 528 -1826
rect 534 -1827 535 -1826
rect 730 -1827 731 -1826
rect 758 -1827 759 -1826
rect 765 -1827 766 -1826
rect 887 -1827 888 -1826
rect 891 -1827 892 -1826
rect 954 -1827 955 -1826
rect 975 -1827 976 -1826
rect 1269 -1827 1270 -1826
rect 1293 -1827 1294 -1826
rect 1584 -1827 1585 -1826
rect 170 -1829 171 -1828
rect 1125 -1829 1126 -1828
rect 1150 -1829 1151 -1828
rect 1164 -1829 1165 -1828
rect 1269 -1829 1270 -1828
rect 1458 -1829 1459 -1828
rect 1577 -1829 1578 -1828
rect 1619 -1829 1620 -1828
rect 212 -1831 213 -1830
rect 443 -1831 444 -1830
rect 471 -1831 472 -1830
rect 625 -1831 626 -1830
rect 733 -1831 734 -1830
rect 828 -1831 829 -1830
rect 831 -1831 832 -1830
rect 1780 -1831 1781 -1830
rect 114 -1833 115 -1832
rect 828 -1833 829 -1832
rect 856 -1833 857 -1832
rect 884 -1833 885 -1832
rect 898 -1833 899 -1832
rect 919 -1833 920 -1832
rect 947 -1833 948 -1832
rect 1384 -1833 1385 -1832
rect 1426 -1833 1427 -1832
rect 1535 -1833 1536 -1832
rect 219 -1835 220 -1834
rect 324 -1835 325 -1834
rect 341 -1835 342 -1834
rect 1094 -1835 1095 -1834
rect 1290 -1835 1291 -1834
rect 1619 -1835 1620 -1834
rect 135 -1837 136 -1836
rect 324 -1837 325 -1836
rect 359 -1837 360 -1836
rect 562 -1837 563 -1836
rect 758 -1837 759 -1836
rect 793 -1837 794 -1836
rect 810 -1837 811 -1836
rect 1311 -1837 1312 -1836
rect 1458 -1837 1459 -1836
rect 1465 -1837 1466 -1836
rect 135 -1839 136 -1838
rect 163 -1839 164 -1838
rect 222 -1839 223 -1838
rect 716 -1839 717 -1838
rect 765 -1839 766 -1838
rect 1059 -1839 1060 -1838
rect 1066 -1839 1067 -1838
rect 1157 -1839 1158 -1838
rect 1311 -1839 1312 -1838
rect 1353 -1839 1354 -1838
rect 1465 -1839 1466 -1838
rect 1472 -1839 1473 -1838
rect 163 -1841 164 -1840
rect 191 -1841 192 -1840
rect 222 -1841 223 -1840
rect 1598 -1841 1599 -1840
rect 191 -1843 192 -1842
rect 254 -1843 255 -1842
rect 261 -1843 262 -1842
rect 499 -1843 500 -1842
rect 527 -1843 528 -1842
rect 1206 -1843 1207 -1842
rect 1353 -1843 1354 -1842
rect 1402 -1843 1403 -1842
rect 1430 -1843 1431 -1842
rect 1472 -1843 1473 -1842
rect 1570 -1843 1571 -1842
rect 1598 -1843 1599 -1842
rect 61 -1845 62 -1844
rect 261 -1845 262 -1844
rect 268 -1845 269 -1844
rect 485 -1845 486 -1844
rect 544 -1845 545 -1844
rect 1290 -1845 1291 -1844
rect 1297 -1845 1298 -1844
rect 1430 -1845 1431 -1844
rect 1570 -1845 1571 -1844
rect 1822 -1845 1823 -1844
rect 173 -1847 174 -1846
rect 1402 -1847 1403 -1846
rect 226 -1849 227 -1848
rect 404 -1849 405 -1848
rect 415 -1849 416 -1848
rect 593 -1849 594 -1848
rect 786 -1849 787 -1848
rect 1647 -1849 1648 -1848
rect 23 -1851 24 -1850
rect 593 -1851 594 -1850
rect 793 -1851 794 -1850
rect 842 -1851 843 -1850
rect 856 -1851 857 -1850
rect 1097 -1851 1098 -1850
rect 1157 -1851 1158 -1850
rect 1717 -1851 1718 -1850
rect 226 -1853 227 -1852
rect 632 -1853 633 -1852
rect 814 -1853 815 -1852
rect 870 -1853 871 -1852
rect 901 -1853 902 -1852
rect 1654 -1853 1655 -1852
rect 233 -1855 234 -1854
rect 289 -1855 290 -1854
rect 303 -1855 304 -1854
rect 380 -1855 381 -1854
rect 394 -1855 395 -1854
rect 789 -1855 790 -1854
rect 821 -1855 822 -1854
rect 1136 -1855 1137 -1854
rect 1297 -1855 1298 -1854
rect 1339 -1855 1340 -1854
rect 1605 -1855 1606 -1854
rect 1717 -1855 1718 -1854
rect 44 -1857 45 -1856
rect 789 -1857 790 -1856
rect 824 -1857 825 -1856
rect 1059 -1857 1060 -1856
rect 1080 -1857 1081 -1856
rect 1136 -1857 1137 -1856
rect 1605 -1857 1606 -1856
rect 1766 -1857 1767 -1856
rect 44 -1859 45 -1858
rect 744 -1859 745 -1858
rect 842 -1859 843 -1858
rect 905 -1859 906 -1858
rect 919 -1859 920 -1858
rect 968 -1859 969 -1858
rect 975 -1859 976 -1858
rect 1017 -1859 1018 -1858
rect 1024 -1859 1025 -1858
rect 1409 -1859 1410 -1858
rect 1647 -1859 1648 -1858
rect 1710 -1859 1711 -1858
rect 219 -1861 220 -1860
rect 303 -1861 304 -1860
rect 317 -1861 318 -1860
rect 506 -1861 507 -1860
rect 562 -1861 563 -1860
rect 800 -1861 801 -1860
rect 870 -1861 871 -1860
rect 1087 -1861 1088 -1860
rect 1094 -1861 1095 -1860
rect 1626 -1861 1627 -1860
rect 1654 -1861 1655 -1860
rect 1703 -1861 1704 -1860
rect 1710 -1861 1711 -1860
rect 1773 -1861 1774 -1860
rect 198 -1863 199 -1862
rect 506 -1863 507 -1862
rect 632 -1863 633 -1862
rect 639 -1863 640 -1862
rect 702 -1863 703 -1862
rect 744 -1863 745 -1862
rect 800 -1863 801 -1862
rect 849 -1863 850 -1862
rect 877 -1863 878 -1862
rect 968 -1863 969 -1862
rect 1017 -1863 1018 -1862
rect 1073 -1863 1074 -1862
rect 1080 -1863 1081 -1862
rect 1115 -1863 1116 -1862
rect 1346 -1863 1347 -1862
rect 1766 -1863 1767 -1862
rect 86 -1865 87 -1864
rect 1073 -1865 1074 -1864
rect 1409 -1865 1410 -1864
rect 1437 -1865 1438 -1864
rect 1626 -1865 1627 -1864
rect 1682 -1865 1683 -1864
rect 1703 -1865 1704 -1864
rect 1759 -1865 1760 -1864
rect 86 -1867 87 -1866
rect 408 -1867 409 -1866
rect 422 -1867 423 -1866
rect 450 -1867 451 -1866
rect 471 -1867 472 -1866
rect 985 -1867 986 -1866
rect 1045 -1867 1046 -1866
rect 1115 -1867 1116 -1866
rect 1437 -1867 1438 -1866
rect 1521 -1867 1522 -1866
rect 1591 -1867 1592 -1866
rect 1682 -1867 1683 -1866
rect 156 -1869 157 -1868
rect 1346 -1869 1347 -1868
rect 1521 -1869 1522 -1868
rect 1542 -1869 1543 -1868
rect 1591 -1869 1592 -1868
rect 1612 -1869 1613 -1868
rect 1633 -1869 1634 -1868
rect 1759 -1869 1760 -1868
rect 156 -1871 157 -1870
rect 247 -1871 248 -1870
rect 254 -1871 255 -1870
rect 719 -1871 720 -1870
rect 849 -1871 850 -1870
rect 1304 -1871 1305 -1870
rect 1542 -1871 1543 -1870
rect 1549 -1871 1550 -1870
rect 1612 -1871 1613 -1870
rect 1675 -1871 1676 -1870
rect 198 -1873 199 -1872
rect 345 -1873 346 -1872
rect 366 -1873 367 -1872
rect 835 -1873 836 -1872
rect 877 -1873 878 -1872
rect 1010 -1873 1011 -1872
rect 1045 -1873 1046 -1872
rect 1171 -1873 1172 -1872
rect 1304 -1873 1305 -1872
rect 1318 -1873 1319 -1872
rect 1549 -1873 1550 -1872
rect 1556 -1873 1557 -1872
rect 1633 -1873 1634 -1872
rect 1696 -1873 1697 -1872
rect 240 -1875 241 -1874
rect 289 -1875 290 -1874
rect 296 -1875 297 -1874
rect 408 -1875 409 -1874
rect 429 -1875 430 -1874
rect 709 -1875 710 -1874
rect 905 -1875 906 -1874
rect 1146 -1875 1147 -1874
rect 1171 -1875 1172 -1874
rect 1220 -1875 1221 -1874
rect 1318 -1875 1319 -1874
rect 1367 -1875 1368 -1874
rect 1675 -1875 1676 -1874
rect 1731 -1875 1732 -1874
rect 275 -1877 276 -1876
rect 520 -1877 521 -1876
rect 618 -1877 619 -1876
rect 639 -1877 640 -1876
rect 702 -1877 703 -1876
rect 961 -1877 962 -1876
rect 1010 -1877 1011 -1876
rect 1031 -1877 1032 -1876
rect 1360 -1877 1361 -1876
rect 1556 -1877 1557 -1876
rect 1696 -1877 1697 -1876
rect 1752 -1877 1753 -1876
rect 275 -1879 276 -1878
rect 660 -1879 661 -1878
rect 688 -1879 689 -1878
rect 961 -1879 962 -1878
rect 1360 -1879 1361 -1878
rect 1388 -1879 1389 -1878
rect 1731 -1879 1732 -1878
rect 1801 -1879 1802 -1878
rect 282 -1881 283 -1880
rect 362 -1881 363 -1880
rect 366 -1881 367 -1880
rect 604 -1881 605 -1880
rect 618 -1881 619 -1880
rect 1339 -1881 1340 -1880
rect 1367 -1881 1368 -1880
rect 1479 -1881 1480 -1880
rect 282 -1883 283 -1882
rect 310 -1883 311 -1882
rect 331 -1883 332 -1882
rect 450 -1883 451 -1882
rect 478 -1883 479 -1882
rect 492 -1883 493 -1882
rect 579 -1883 580 -1882
rect 1388 -1883 1389 -1882
rect 1479 -1883 1480 -1882
rect 1500 -1883 1501 -1882
rect 205 -1885 206 -1884
rect 310 -1885 311 -1884
rect 331 -1885 332 -1884
rect 338 -1885 339 -1884
rect 345 -1885 346 -1884
rect 1160 -1885 1161 -1884
rect 1500 -1885 1501 -1884
rect 1507 -1885 1508 -1884
rect 205 -1887 206 -1886
rect 940 -1887 941 -1886
rect 954 -1887 955 -1886
rect 1003 -1887 1004 -1886
rect 1507 -1887 1508 -1886
rect 1514 -1887 1515 -1886
rect 296 -1889 297 -1888
rect 464 -1889 465 -1888
rect 485 -1889 486 -1888
rect 653 -1889 654 -1888
rect 660 -1889 661 -1888
rect 681 -1889 682 -1888
rect 688 -1889 689 -1888
rect 978 -1889 979 -1888
rect 1514 -1889 1515 -1888
rect 1528 -1889 1529 -1888
rect 121 -1891 122 -1890
rect 653 -1891 654 -1890
rect 681 -1891 682 -1890
rect 1038 -1891 1039 -1890
rect 1486 -1891 1487 -1890
rect 1528 -1891 1529 -1890
rect 121 -1893 122 -1892
rect 737 -1893 738 -1892
rect 779 -1893 780 -1892
rect 1220 -1893 1221 -1892
rect 380 -1895 381 -1894
rect 383 -1895 384 -1894
rect 401 -1895 402 -1894
rect 464 -1895 465 -1894
rect 492 -1895 493 -1894
rect 912 -1895 913 -1894
rect 933 -1895 934 -1894
rect 1031 -1895 1032 -1894
rect 1038 -1895 1039 -1894
rect 1108 -1895 1109 -1894
rect 1129 -1895 1130 -1894
rect 1486 -1895 1487 -1894
rect 401 -1897 402 -1896
rect 1724 -1897 1725 -1896
rect 436 -1899 437 -1898
rect 604 -1899 605 -1898
rect 737 -1899 738 -1898
rect 807 -1899 808 -1898
rect 912 -1899 913 -1898
rect 1395 -1899 1396 -1898
rect 51 -1901 52 -1900
rect 807 -1901 808 -1900
rect 933 -1901 934 -1900
rect 982 -1901 983 -1900
rect 1108 -1901 1109 -1900
rect 1276 -1901 1277 -1900
rect 51 -1903 52 -1902
rect 243 -1903 244 -1902
rect 436 -1903 437 -1902
rect 555 -1903 556 -1902
rect 751 -1903 752 -1902
rect 779 -1903 780 -1902
rect 940 -1903 941 -1902
rect 996 -1903 997 -1902
rect 1122 -1903 1123 -1902
rect 1276 -1903 1277 -1902
rect 551 -1905 552 -1904
rect 1003 -1905 1004 -1904
rect 1129 -1905 1130 -1904
rect 1199 -1905 1200 -1904
rect 555 -1907 556 -1906
rect 569 -1907 570 -1906
rect 751 -1907 752 -1906
rect 926 -1907 927 -1906
rect 1199 -1907 1200 -1906
rect 1255 -1907 1256 -1906
rect 513 -1909 514 -1908
rect 569 -1909 570 -1908
rect 926 -1909 927 -1908
rect 989 -1909 990 -1908
rect 1241 -1909 1242 -1908
rect 1255 -1909 1256 -1908
rect 107 -1911 108 -1910
rect 513 -1911 514 -1910
rect 1185 -1911 1186 -1910
rect 1241 -1911 1242 -1910
rect 107 -1913 108 -1912
rect 863 -1913 864 -1912
rect 1185 -1913 1186 -1912
rect 1248 -1913 1249 -1912
rect 233 -1915 234 -1914
rect 989 -1915 990 -1914
rect 1248 -1915 1249 -1914
rect 1262 -1915 1263 -1914
rect 590 -1917 591 -1916
rect 1262 -1917 1263 -1916
rect 590 -1919 591 -1918
rect 996 -1919 997 -1918
rect 863 -1921 864 -1920
rect 1167 -1921 1168 -1920
rect 23 -1932 24 -1931
rect 936 -1932 937 -1931
rect 950 -1932 951 -1931
rect 1136 -1932 1137 -1931
rect 1157 -1932 1158 -1931
rect 1766 -1932 1767 -1931
rect 30 -1934 31 -1933
rect 61 -1934 62 -1933
rect 65 -1934 66 -1933
rect 506 -1934 507 -1933
rect 534 -1934 535 -1933
rect 607 -1934 608 -1933
rect 618 -1934 619 -1933
rect 1290 -1934 1291 -1933
rect 1381 -1934 1382 -1933
rect 1675 -1934 1676 -1933
rect 1738 -1934 1739 -1933
rect 1773 -1934 1774 -1933
rect 37 -1936 38 -1935
rect 170 -1936 171 -1935
rect 219 -1936 220 -1935
rect 394 -1936 395 -1935
rect 408 -1936 409 -1935
rect 600 -1936 601 -1935
rect 656 -1936 657 -1935
rect 1717 -1936 1718 -1935
rect 37 -1938 38 -1937
rect 86 -1938 87 -1937
rect 93 -1938 94 -1937
rect 768 -1938 769 -1937
rect 772 -1938 773 -1937
rect 933 -1938 934 -1937
rect 985 -1938 986 -1937
rect 1360 -1938 1361 -1937
rect 1381 -1938 1382 -1937
rect 1395 -1938 1396 -1937
rect 1640 -1938 1641 -1937
rect 1738 -1938 1739 -1937
rect 58 -1940 59 -1939
rect 604 -1940 605 -1939
rect 716 -1940 717 -1939
rect 803 -1940 804 -1939
rect 849 -1940 850 -1939
rect 898 -1940 899 -1939
rect 912 -1940 913 -1939
rect 1591 -1940 1592 -1939
rect 1640 -1940 1641 -1939
rect 1654 -1940 1655 -1939
rect 1675 -1940 1676 -1939
rect 1710 -1940 1711 -1939
rect 1717 -1940 1718 -1939
rect 1745 -1940 1746 -1939
rect 68 -1942 69 -1941
rect 1689 -1942 1690 -1941
rect 1710 -1942 1711 -1941
rect 1724 -1942 1725 -1941
rect 79 -1944 80 -1943
rect 93 -1944 94 -1943
rect 100 -1944 101 -1943
rect 534 -1944 535 -1943
rect 604 -1944 605 -1943
rect 681 -1944 682 -1943
rect 716 -1944 717 -1943
rect 730 -1944 731 -1943
rect 754 -1944 755 -1943
rect 821 -1944 822 -1943
rect 873 -1944 874 -1943
rect 1108 -1944 1109 -1943
rect 1122 -1944 1123 -1943
rect 1493 -1944 1494 -1943
rect 1500 -1944 1501 -1943
rect 1689 -1944 1690 -1943
rect 79 -1946 80 -1945
rect 135 -1946 136 -1945
rect 138 -1946 139 -1945
rect 639 -1946 640 -1945
rect 646 -1946 647 -1945
rect 681 -1946 682 -1945
rect 723 -1946 724 -1945
rect 933 -1946 934 -1945
rect 989 -1946 990 -1945
rect 1367 -1946 1368 -1945
rect 1384 -1946 1385 -1945
rect 1528 -1946 1529 -1945
rect 1549 -1946 1550 -1945
rect 1591 -1946 1592 -1945
rect 1654 -1946 1655 -1945
rect 1661 -1946 1662 -1945
rect 1682 -1946 1683 -1945
rect 1745 -1946 1746 -1945
rect 100 -1948 101 -1947
rect 142 -1948 143 -1947
rect 149 -1948 150 -1947
rect 908 -1948 909 -1947
rect 912 -1948 913 -1947
rect 954 -1948 955 -1947
rect 1059 -1948 1060 -1947
rect 1766 -1948 1767 -1947
rect 107 -1950 108 -1949
rect 317 -1950 318 -1949
rect 359 -1950 360 -1949
rect 870 -1950 871 -1949
rect 898 -1950 899 -1949
rect 940 -1950 941 -1949
rect 947 -1950 948 -1949
rect 989 -1950 990 -1949
rect 1080 -1950 1081 -1949
rect 1108 -1950 1109 -1949
rect 1157 -1950 1158 -1949
rect 1171 -1950 1172 -1949
rect 1185 -1950 1186 -1949
rect 1188 -1950 1189 -1949
rect 1227 -1950 1228 -1949
rect 1416 -1950 1417 -1949
rect 1423 -1950 1424 -1949
rect 1500 -1950 1501 -1949
rect 1528 -1950 1529 -1949
rect 1762 -1950 1763 -1949
rect 135 -1952 136 -1951
rect 1220 -1952 1221 -1951
rect 1290 -1952 1291 -1951
rect 1472 -1952 1473 -1951
rect 1570 -1952 1571 -1951
rect 1724 -1952 1725 -1951
rect 142 -1954 143 -1953
rect 541 -1954 542 -1953
rect 597 -1954 598 -1953
rect 954 -1954 955 -1953
rect 1066 -1954 1067 -1953
rect 1080 -1954 1081 -1953
rect 1087 -1954 1088 -1953
rect 1122 -1954 1123 -1953
rect 1160 -1954 1161 -1953
rect 1759 -1954 1760 -1953
rect 149 -1956 150 -1955
rect 163 -1956 164 -1955
rect 166 -1956 167 -1955
rect 709 -1956 710 -1955
rect 730 -1956 731 -1955
rect 1020 -1956 1021 -1955
rect 1097 -1956 1098 -1955
rect 1437 -1956 1438 -1955
rect 1661 -1956 1662 -1955
rect 1668 -1956 1669 -1955
rect 1682 -1956 1683 -1955
rect 1752 -1956 1753 -1955
rect 1759 -1956 1760 -1955
rect 1794 -1956 1795 -1955
rect 65 -1958 66 -1957
rect 163 -1958 164 -1957
rect 170 -1958 171 -1957
rect 415 -1958 416 -1957
rect 432 -1958 433 -1957
rect 1136 -1958 1137 -1957
rect 1167 -1958 1168 -1957
rect 1647 -1958 1648 -1957
rect 1668 -1958 1669 -1957
rect 1703 -1958 1704 -1957
rect 159 -1960 160 -1959
rect 352 -1960 353 -1959
rect 359 -1960 360 -1959
rect 527 -1960 528 -1959
rect 639 -1960 640 -1959
rect 919 -1960 920 -1959
rect 929 -1960 930 -1959
rect 1570 -1960 1571 -1959
rect 1696 -1960 1697 -1959
rect 1703 -1960 1704 -1959
rect 72 -1962 73 -1961
rect 352 -1962 353 -1961
rect 380 -1962 381 -1961
rect 621 -1962 622 -1961
rect 646 -1962 647 -1961
rect 660 -1962 661 -1961
rect 670 -1962 671 -1961
rect 1696 -1962 1697 -1961
rect 72 -1964 73 -1963
rect 131 -1964 132 -1963
rect 219 -1964 220 -1963
rect 373 -1964 374 -1963
rect 394 -1964 395 -1963
rect 436 -1964 437 -1963
rect 471 -1964 472 -1963
rect 541 -1964 542 -1963
rect 621 -1964 622 -1963
rect 1535 -1964 1536 -1963
rect 51 -1966 52 -1965
rect 471 -1966 472 -1965
rect 492 -1966 493 -1965
rect 593 -1966 594 -1965
rect 660 -1966 661 -1965
rect 1150 -1966 1151 -1965
rect 1171 -1966 1172 -1965
rect 1178 -1966 1179 -1965
rect 1185 -1966 1186 -1965
rect 1241 -1966 1242 -1965
rect 1325 -1966 1326 -1965
rect 1472 -1966 1473 -1965
rect 51 -1968 52 -1967
rect 345 -1968 346 -1967
rect 373 -1968 374 -1967
rect 817 -1968 818 -1967
rect 821 -1968 822 -1967
rect 856 -1968 857 -1967
rect 877 -1968 878 -1967
rect 1150 -1968 1151 -1967
rect 1178 -1968 1179 -1967
rect 1563 -1968 1564 -1967
rect 117 -1970 118 -1969
rect 436 -1970 437 -1969
rect 450 -1970 451 -1969
rect 492 -1970 493 -1969
rect 506 -1970 507 -1969
rect 569 -1970 570 -1969
rect 593 -1970 594 -1969
rect 1395 -1970 1396 -1969
rect 1444 -1970 1445 -1969
rect 1647 -1970 1648 -1969
rect 226 -1972 227 -1971
rect 310 -1972 311 -1971
rect 324 -1972 325 -1971
rect 380 -1972 381 -1971
rect 401 -1972 402 -1971
rect 1066 -1972 1067 -1971
rect 1101 -1972 1102 -1971
rect 1416 -1972 1417 -1971
rect 1444 -1972 1445 -1971
rect 1465 -1972 1466 -1971
rect 1514 -1972 1515 -1971
rect 1563 -1972 1564 -1971
rect 177 -1974 178 -1973
rect 226 -1974 227 -1973
rect 240 -1974 241 -1973
rect 338 -1974 339 -1973
rect 345 -1974 346 -1973
rect 513 -1974 514 -1973
rect 555 -1974 556 -1973
rect 569 -1974 570 -1973
rect 670 -1974 671 -1973
rect 905 -1974 906 -1973
rect 915 -1974 916 -1973
rect 1248 -1974 1249 -1973
rect 1353 -1974 1354 -1973
rect 1549 -1974 1550 -1973
rect 156 -1976 157 -1975
rect 513 -1976 514 -1975
rect 691 -1976 692 -1975
rect 1514 -1976 1515 -1975
rect 156 -1978 157 -1977
rect 726 -1978 727 -1977
rect 765 -1978 766 -1977
rect 1493 -1978 1494 -1977
rect 177 -1980 178 -1979
rect 985 -1980 986 -1979
rect 1024 -1980 1025 -1979
rect 1353 -1980 1354 -1979
rect 1360 -1980 1361 -1979
rect 1374 -1980 1375 -1979
rect 1388 -1980 1389 -1979
rect 1423 -1980 1424 -1979
rect 184 -1982 185 -1981
rect 338 -1982 339 -1981
rect 401 -1982 402 -1981
rect 684 -1982 685 -1981
rect 695 -1982 696 -1981
rect 709 -1982 710 -1981
rect 765 -1982 766 -1981
rect 1059 -1982 1060 -1981
rect 1073 -1982 1074 -1981
rect 1101 -1982 1102 -1981
rect 1115 -1982 1116 -1981
rect 1220 -1982 1221 -1981
rect 1230 -1982 1231 -1981
rect 1248 -1982 1249 -1981
rect 1367 -1982 1368 -1981
rect 1451 -1982 1452 -1981
rect 184 -1984 185 -1983
rect 835 -1984 836 -1983
rect 856 -1984 857 -1983
rect 1206 -1984 1207 -1983
rect 1213 -1984 1214 -1983
rect 1227 -1984 1228 -1983
rect 1374 -1984 1375 -1983
rect 1479 -1984 1480 -1983
rect 205 -1986 206 -1985
rect 835 -1986 836 -1985
rect 905 -1986 906 -1985
rect 1612 -1986 1613 -1985
rect 205 -1988 206 -1987
rect 208 -1988 209 -1987
rect 233 -1988 234 -1987
rect 695 -1988 696 -1987
rect 702 -1988 703 -1987
rect 870 -1988 871 -1987
rect 940 -1988 941 -1987
rect 975 -1988 976 -1987
rect 1038 -1988 1039 -1987
rect 1073 -1988 1074 -1987
rect 1087 -1988 1088 -1987
rect 1115 -1988 1116 -1987
rect 1192 -1988 1193 -1987
rect 1241 -1988 1242 -1987
rect 1388 -1988 1389 -1987
rect 1402 -1988 1403 -1987
rect 1409 -1988 1410 -1987
rect 1465 -1988 1466 -1987
rect 1584 -1988 1585 -1987
rect 1612 -1988 1613 -1987
rect 233 -1990 234 -1989
rect 597 -1990 598 -1989
rect 702 -1990 703 -1989
rect 996 -1990 997 -1989
rect 1017 -1990 1018 -1989
rect 1038 -1990 1039 -1989
rect 1188 -1990 1189 -1989
rect 1192 -1990 1193 -1989
rect 1213 -1990 1214 -1989
rect 1339 -1990 1340 -1989
rect 1402 -1990 1403 -1989
rect 1542 -1990 1543 -1989
rect 240 -1992 241 -1991
rect 387 -1992 388 -1991
rect 408 -1992 409 -1991
rect 653 -1992 654 -1991
rect 688 -1992 689 -1991
rect 996 -1992 997 -1991
rect 1017 -1992 1018 -1991
rect 1283 -1992 1284 -1991
rect 1409 -1992 1410 -1991
rect 1458 -1992 1459 -1991
rect 1542 -1992 1543 -1991
rect 1605 -1992 1606 -1991
rect 247 -1994 248 -1993
rect 310 -1994 311 -1993
rect 324 -1994 325 -1993
rect 674 -1994 675 -1993
rect 772 -1994 773 -1993
rect 842 -1994 843 -1993
rect 975 -1994 976 -1993
rect 1003 -1994 1004 -1993
rect 1129 -1994 1130 -1993
rect 1339 -1994 1340 -1993
rect 1430 -1994 1431 -1993
rect 1479 -1994 1480 -1993
rect 1598 -1994 1599 -1993
rect 1605 -1994 1606 -1993
rect 107 -1996 108 -1995
rect 674 -1996 675 -1995
rect 789 -1996 790 -1995
rect 1024 -1996 1025 -1995
rect 1052 -1996 1053 -1995
rect 1129 -1996 1130 -1995
rect 1276 -1996 1277 -1995
rect 1283 -1996 1284 -1995
rect 1332 -1996 1333 -1995
rect 1430 -1996 1431 -1995
rect 1556 -1996 1557 -1995
rect 1598 -1996 1599 -1995
rect 243 -1998 244 -1997
rect 247 -1998 248 -1997
rect 250 -1998 251 -1997
rect 1255 -1998 1256 -1997
rect 1332 -1998 1333 -1997
rect 1346 -1998 1347 -1997
rect 1556 -1998 1557 -1997
rect 1577 -1998 1578 -1997
rect 254 -2000 255 -1999
rect 415 -2000 416 -1999
rect 450 -2000 451 -1999
rect 635 -2000 636 -1999
rect 667 -2000 668 -1999
rect 1052 -2000 1053 -1999
rect 1255 -2000 1256 -1999
rect 1437 -2000 1438 -1999
rect 1577 -2000 1578 -1999
rect 1731 -2000 1732 -1999
rect 254 -2002 255 -2001
rect 289 -2002 290 -2001
rect 303 -2002 304 -2001
rect 317 -2002 318 -2001
rect 387 -2002 388 -2001
rect 548 -2002 549 -2001
rect 576 -2002 577 -2001
rect 653 -2002 654 -2001
rect 667 -2002 668 -2001
rect 1325 -2002 1326 -2001
rect 1346 -2002 1347 -2001
rect 1507 -2002 1508 -2001
rect 1521 -2002 1522 -2001
rect 1731 -2002 1732 -2001
rect 268 -2004 269 -2003
rect 618 -2004 619 -2003
rect 800 -2004 801 -2003
rect 982 -2004 983 -2003
rect 1003 -2004 1004 -2003
rect 1010 -2004 1011 -2003
rect 1262 -2004 1263 -2003
rect 1507 -2004 1508 -2003
rect 198 -2006 199 -2005
rect 268 -2006 269 -2005
rect 275 -2006 276 -2005
rect 530 -2006 531 -2005
rect 548 -2006 549 -2005
rect 688 -2006 689 -2005
rect 800 -2006 801 -2005
rect 877 -2006 878 -2005
rect 1010 -2006 1011 -2005
rect 1164 -2006 1165 -2005
rect 1311 -2006 1312 -2005
rect 1521 -2006 1522 -2005
rect 110 -2008 111 -2007
rect 275 -2008 276 -2007
rect 282 -2008 283 -2007
rect 369 -2008 370 -2007
rect 457 -2008 458 -2007
rect 576 -2008 577 -2007
rect 590 -2008 591 -2007
rect 1584 -2008 1585 -2007
rect 114 -2010 115 -2009
rect 198 -2010 199 -2009
rect 229 -2010 230 -2009
rect 1311 -2010 1312 -2009
rect 114 -2012 115 -2011
rect 1276 -2012 1277 -2011
rect 282 -2014 283 -2013
rect 782 -2014 783 -2013
rect 807 -2014 808 -2013
rect 919 -2014 920 -2013
rect 1045 -2014 1046 -2013
rect 1262 -2014 1263 -2013
rect 289 -2016 290 -2015
rect 429 -2016 430 -2015
rect 457 -2016 458 -2015
rect 625 -2016 626 -2015
rect 793 -2016 794 -2015
rect 807 -2016 808 -2015
rect 810 -2016 811 -2015
rect 1535 -2016 1536 -2015
rect 303 -2018 304 -2017
rect 331 -2018 332 -2017
rect 404 -2018 405 -2017
rect 1045 -2018 1046 -2017
rect 1164 -2018 1165 -2017
rect 1258 -2018 1259 -2017
rect 331 -2020 332 -2019
rect 366 -2020 367 -2019
rect 429 -2020 430 -2019
rect 611 -2020 612 -2019
rect 625 -2020 626 -2019
rect 863 -2020 864 -2019
rect 485 -2022 486 -2021
rect 611 -2022 612 -2021
rect 814 -2022 815 -2021
rect 842 -2022 843 -2021
rect 863 -2022 864 -2021
rect 891 -2022 892 -2021
rect 443 -2024 444 -2023
rect 485 -2024 486 -2023
rect 499 -2024 500 -2023
rect 1206 -2024 1207 -2023
rect 422 -2026 423 -2025
rect 443 -2026 444 -2025
rect 478 -2026 479 -2025
rect 499 -2026 500 -2025
rect 530 -2026 531 -2025
rect 555 -2026 556 -2025
rect 562 -2026 563 -2025
rect 793 -2026 794 -2025
rect 814 -2026 815 -2025
rect 1486 -2026 1487 -2025
rect 44 -2028 45 -2027
rect 422 -2028 423 -2027
rect 562 -2028 563 -2027
rect 961 -2028 962 -2027
rect 1125 -2028 1126 -2027
rect 1486 -2028 1487 -2027
rect 44 -2030 45 -2029
rect 128 -2030 129 -2029
rect 212 -2030 213 -2029
rect 478 -2030 479 -2029
rect 590 -2030 591 -2029
rect 758 -2030 759 -2029
rect 891 -2030 892 -2029
rect 926 -2030 927 -2029
rect 961 -2030 962 -2029
rect 1031 -2030 1032 -2029
rect 128 -2032 129 -2031
rect 191 -2032 192 -2031
rect 212 -2032 213 -2031
rect 261 -2032 262 -2031
rect 737 -2032 738 -2031
rect 926 -2032 927 -2031
rect 121 -2034 122 -2033
rect 737 -2034 738 -2033
rect 758 -2034 759 -2033
rect 779 -2034 780 -2033
rect 828 -2034 829 -2033
rect 1031 -2034 1032 -2033
rect 121 -2036 122 -2035
rect 1094 -2036 1095 -2035
rect 173 -2038 174 -2037
rect 1094 -2038 1095 -2037
rect 191 -2040 192 -2039
rect 296 -2040 297 -2039
rect 786 -2040 787 -2039
rect 828 -2040 829 -2039
rect 261 -2042 262 -2041
rect 520 -2042 521 -2041
rect 751 -2042 752 -2041
rect 786 -2042 787 -2041
rect 296 -2044 297 -2043
rect 464 -2044 465 -2043
rect 520 -2044 521 -2043
rect 663 -2044 664 -2043
rect 751 -2044 752 -2043
rect 1458 -2044 1459 -2043
rect 464 -2046 465 -2045
rect 632 -2046 633 -2045
rect 86 -2048 87 -2047
rect 632 -2048 633 -2047
rect 40 -2059 41 -2058
rect 1549 -2059 1550 -2058
rect 1626 -2059 1627 -2058
rect 1629 -2059 1630 -2058
rect 1759 -2059 1760 -2058
rect 1766 -2059 1767 -2058
rect 44 -2061 45 -2060
rect 152 -2061 153 -2060
rect 163 -2061 164 -2060
rect 562 -2061 563 -2060
rect 632 -2061 633 -2060
rect 1521 -2061 1522 -2060
rect 1626 -2061 1627 -2060
rect 1654 -2061 1655 -2060
rect 1766 -2061 1767 -2060
rect 1773 -2061 1774 -2060
rect 23 -2063 24 -2062
rect 562 -2063 563 -2062
rect 663 -2063 664 -2062
rect 716 -2063 717 -2062
rect 726 -2063 727 -2062
rect 1017 -2063 1018 -2062
rect 1090 -2063 1091 -2062
rect 1290 -2063 1291 -2062
rect 1346 -2063 1347 -2062
rect 1521 -2063 1522 -2062
rect 47 -2065 48 -2064
rect 681 -2065 682 -2064
rect 688 -2065 689 -2064
rect 737 -2065 738 -2064
rect 782 -2065 783 -2064
rect 1178 -2065 1179 -2064
rect 1206 -2065 1207 -2064
rect 1752 -2065 1753 -2064
rect 68 -2067 69 -2066
rect 135 -2067 136 -2066
rect 142 -2067 143 -2066
rect 800 -2067 801 -2066
rect 803 -2067 804 -2066
rect 1563 -2067 1564 -2066
rect 100 -2069 101 -2068
rect 779 -2069 780 -2068
rect 786 -2069 787 -2068
rect 800 -2069 801 -2068
rect 873 -2069 874 -2068
rect 1762 -2069 1763 -2068
rect 100 -2071 101 -2070
rect 856 -2071 857 -2070
rect 919 -2071 920 -2070
rect 922 -2071 923 -2070
rect 926 -2071 927 -2070
rect 1416 -2071 1417 -2070
rect 1451 -2071 1452 -2070
rect 1598 -2071 1599 -2070
rect 107 -2073 108 -2072
rect 705 -2073 706 -2072
rect 716 -2073 717 -2072
rect 744 -2073 745 -2072
rect 758 -2073 759 -2072
rect 786 -2073 787 -2072
rect 856 -2073 857 -2072
rect 877 -2073 878 -2072
rect 912 -2073 913 -2072
rect 926 -2073 927 -2072
rect 936 -2073 937 -2072
rect 1703 -2073 1704 -2072
rect 107 -2075 108 -2074
rect 369 -2075 370 -2074
rect 436 -2075 437 -2074
rect 761 -2075 762 -2074
rect 779 -2075 780 -2074
rect 870 -2075 871 -2074
rect 877 -2075 878 -2074
rect 954 -2075 955 -2074
rect 985 -2075 986 -2074
rect 1549 -2075 1550 -2074
rect 1703 -2075 1704 -2074
rect 1710 -2075 1711 -2074
rect 114 -2077 115 -2076
rect 296 -2077 297 -2076
rect 352 -2077 353 -2076
rect 436 -2077 437 -2076
rect 453 -2077 454 -2076
rect 499 -2077 500 -2076
rect 506 -2077 507 -2076
rect 681 -2077 682 -2076
rect 744 -2077 745 -2076
rect 1591 -2077 1592 -2076
rect 1696 -2077 1697 -2076
rect 1710 -2077 1711 -2076
rect 54 -2079 55 -2078
rect 114 -2079 115 -2078
rect 128 -2079 129 -2078
rect 1465 -2079 1466 -2078
rect 1570 -2079 1571 -2078
rect 1591 -2079 1592 -2078
rect 1682 -2079 1683 -2078
rect 1696 -2079 1697 -2078
rect 128 -2081 129 -2080
rect 275 -2081 276 -2080
rect 289 -2081 290 -2080
rect 352 -2081 353 -2080
rect 359 -2081 360 -2080
rect 621 -2081 622 -2080
rect 667 -2081 668 -2080
rect 807 -2081 808 -2080
rect 898 -2081 899 -2080
rect 912 -2081 913 -2080
rect 919 -2081 920 -2080
rect 940 -2081 941 -2080
rect 947 -2081 948 -2080
rect 1339 -2081 1340 -2080
rect 1395 -2081 1396 -2080
rect 1416 -2081 1417 -2080
rect 1451 -2081 1452 -2080
rect 1556 -2081 1557 -2080
rect 1605 -2081 1606 -2080
rect 1682 -2081 1683 -2080
rect 121 -2083 122 -2082
rect 667 -2083 668 -2082
rect 674 -2083 675 -2082
rect 754 -2083 755 -2082
rect 758 -2083 759 -2082
rect 1262 -2083 1263 -2082
rect 1269 -2083 1270 -2082
rect 1465 -2083 1466 -2082
rect 1528 -2083 1529 -2082
rect 1556 -2083 1557 -2082
rect 1605 -2083 1606 -2082
rect 1612 -2083 1613 -2082
rect 1629 -2083 1630 -2082
rect 1654 -2083 1655 -2082
rect 121 -2085 122 -2084
rect 149 -2085 150 -2084
rect 163 -2085 164 -2084
rect 821 -2085 822 -2084
rect 884 -2085 885 -2084
rect 947 -2085 948 -2084
rect 989 -2085 990 -2084
rect 1020 -2085 1021 -2084
rect 1104 -2085 1105 -2084
rect 1689 -2085 1690 -2084
rect 173 -2087 174 -2086
rect 1423 -2087 1424 -2086
rect 1500 -2087 1501 -2086
rect 1528 -2087 1529 -2086
rect 1535 -2087 1536 -2086
rect 1570 -2087 1571 -2086
rect 1612 -2087 1613 -2086
rect 1633 -2087 1634 -2086
rect 177 -2089 178 -2088
rect 817 -2089 818 -2088
rect 821 -2089 822 -2088
rect 842 -2089 843 -2088
rect 936 -2089 937 -2088
rect 1262 -2089 1263 -2088
rect 1311 -2089 1312 -2088
rect 1346 -2089 1347 -2088
rect 1353 -2089 1354 -2088
rect 1395 -2089 1396 -2088
rect 1402 -2089 1403 -2088
rect 1563 -2089 1564 -2088
rect 1619 -2089 1620 -2088
rect 1633 -2089 1634 -2088
rect 177 -2091 178 -2090
rect 324 -2091 325 -2090
rect 331 -2091 332 -2090
rect 506 -2091 507 -2090
rect 534 -2091 535 -2090
rect 747 -2091 748 -2090
rect 989 -2091 990 -2090
rect 1038 -2091 1039 -2090
rect 1157 -2091 1158 -2090
rect 1178 -2091 1179 -2090
rect 1199 -2091 1200 -2090
rect 1206 -2091 1207 -2090
rect 1227 -2091 1228 -2090
rect 1290 -2091 1291 -2090
rect 1325 -2091 1326 -2090
rect 1353 -2091 1354 -2090
rect 1402 -2091 1403 -2090
rect 1444 -2091 1445 -2090
rect 1584 -2091 1585 -2090
rect 1619 -2091 1620 -2090
rect 51 -2093 52 -2092
rect 534 -2093 535 -2092
rect 555 -2093 556 -2092
rect 954 -2093 955 -2092
rect 1010 -2093 1011 -2092
rect 1038 -2093 1039 -2092
rect 1073 -2093 1074 -2092
rect 1227 -2093 1228 -2092
rect 1255 -2093 1256 -2092
rect 1598 -2093 1599 -2092
rect 184 -2095 185 -2094
rect 737 -2095 738 -2094
rect 950 -2095 951 -2094
rect 1199 -2095 1200 -2094
rect 1258 -2095 1259 -2094
rect 1731 -2095 1732 -2094
rect 184 -2097 185 -2096
rect 373 -2097 374 -2096
rect 408 -2097 409 -2096
rect 842 -2097 843 -2096
rect 1017 -2097 1018 -2096
rect 1031 -2097 1032 -2096
rect 1073 -2097 1074 -2096
rect 1220 -2097 1221 -2096
rect 1339 -2097 1340 -2096
rect 1367 -2097 1368 -2096
rect 1423 -2097 1424 -2096
rect 1647 -2097 1648 -2096
rect 1717 -2097 1718 -2096
rect 1731 -2097 1732 -2096
rect 191 -2099 192 -2098
rect 635 -2099 636 -2098
rect 674 -2099 675 -2098
rect 723 -2099 724 -2098
rect 817 -2099 818 -2098
rect 1717 -2099 1718 -2098
rect 142 -2101 143 -2100
rect 723 -2101 724 -2100
rect 1031 -2101 1032 -2100
rect 1045 -2101 1046 -2100
rect 1118 -2101 1119 -2100
rect 1325 -2101 1326 -2100
rect 1444 -2101 1445 -2100
rect 1748 -2101 1749 -2100
rect 191 -2103 192 -2102
rect 261 -2103 262 -2102
rect 289 -2103 290 -2102
rect 814 -2103 815 -2102
rect 1045 -2103 1046 -2102
rect 1052 -2103 1053 -2102
rect 1129 -2103 1130 -2102
rect 1367 -2103 1368 -2102
rect 1542 -2103 1543 -2102
rect 1647 -2103 1648 -2102
rect 205 -2105 206 -2104
rect 1514 -2105 1515 -2104
rect 1584 -2105 1585 -2104
rect 1668 -2105 1669 -2104
rect 96 -2107 97 -2106
rect 1668 -2107 1669 -2106
rect 205 -2109 206 -2108
rect 268 -2109 269 -2108
rect 296 -2109 297 -2108
rect 303 -2109 304 -2108
rect 310 -2109 311 -2108
rect 331 -2109 332 -2108
rect 345 -2109 346 -2108
rect 359 -2109 360 -2108
rect 366 -2109 367 -2108
rect 1255 -2109 1256 -2108
rect 1374 -2109 1375 -2108
rect 1514 -2109 1515 -2108
rect 208 -2111 209 -2110
rect 632 -2111 633 -2110
rect 691 -2111 692 -2110
rect 898 -2111 899 -2110
rect 1052 -2111 1053 -2110
rect 1108 -2111 1109 -2110
rect 1115 -2111 1116 -2110
rect 1129 -2111 1130 -2110
rect 1157 -2111 1158 -2110
rect 1213 -2111 1214 -2110
rect 1220 -2111 1221 -2110
rect 1234 -2111 1235 -2110
rect 1332 -2111 1333 -2110
rect 1374 -2111 1375 -2110
rect 1507 -2111 1508 -2110
rect 1542 -2111 1543 -2110
rect 212 -2113 213 -2112
rect 303 -2113 304 -2112
rect 310 -2113 311 -2112
rect 317 -2113 318 -2112
rect 324 -2113 325 -2112
rect 1013 -2113 1014 -2112
rect 1101 -2113 1102 -2112
rect 1108 -2113 1109 -2112
rect 1115 -2113 1116 -2112
rect 1500 -2113 1501 -2112
rect 79 -2115 80 -2114
rect 317 -2115 318 -2114
rect 338 -2115 339 -2114
rect 366 -2115 367 -2114
rect 373 -2115 374 -2114
rect 394 -2115 395 -2114
rect 408 -2115 409 -2114
rect 548 -2115 549 -2114
rect 555 -2115 556 -2114
rect 569 -2115 570 -2114
rect 576 -2115 577 -2114
rect 688 -2115 689 -2114
rect 1171 -2115 1172 -2114
rect 1311 -2115 1312 -2114
rect 1472 -2115 1473 -2114
rect 1507 -2115 1508 -2114
rect 79 -2117 80 -2116
rect 1745 -2117 1746 -2116
rect 156 -2119 157 -2118
rect 394 -2119 395 -2118
rect 422 -2119 423 -2118
rect 807 -2119 808 -2118
rect 1192 -2119 1193 -2118
rect 1213 -2119 1214 -2118
rect 1234 -2119 1235 -2118
rect 1248 -2119 1249 -2118
rect 1437 -2119 1438 -2118
rect 1472 -2119 1473 -2118
rect 1724 -2119 1725 -2118
rect 1745 -2119 1746 -2118
rect 131 -2121 132 -2120
rect 156 -2121 157 -2120
rect 166 -2121 167 -2120
rect 576 -2121 577 -2120
rect 593 -2121 594 -2120
rect 1332 -2121 1333 -2120
rect 1409 -2121 1410 -2120
rect 1437 -2121 1438 -2120
rect 1577 -2121 1578 -2120
rect 1724 -2121 1725 -2120
rect 212 -2123 213 -2122
rect 831 -2123 832 -2122
rect 905 -2123 906 -2122
rect 1577 -2123 1578 -2122
rect 233 -2125 234 -2124
rect 527 -2125 528 -2124
rect 541 -2125 542 -2124
rect 548 -2125 549 -2124
rect 569 -2125 570 -2124
rect 772 -2125 773 -2124
rect 1192 -2125 1193 -2124
rect 1276 -2125 1277 -2124
rect 1388 -2125 1389 -2124
rect 1409 -2125 1410 -2124
rect 233 -2127 234 -2126
rect 254 -2127 255 -2126
rect 338 -2127 339 -2126
rect 415 -2127 416 -2126
rect 429 -2127 430 -2126
rect 499 -2127 500 -2126
rect 530 -2127 531 -2126
rect 541 -2127 542 -2126
rect 607 -2127 608 -2126
rect 1535 -2127 1536 -2126
rect 86 -2129 87 -2128
rect 254 -2129 255 -2128
rect 345 -2129 346 -2128
rect 733 -2129 734 -2128
rect 765 -2129 766 -2128
rect 1171 -2129 1172 -2128
rect 1276 -2129 1277 -2128
rect 1640 -2129 1641 -2128
rect 37 -2131 38 -2130
rect 765 -2131 766 -2130
rect 772 -2131 773 -2130
rect 1493 -2131 1494 -2130
rect 86 -2133 87 -2132
rect 478 -2133 479 -2132
rect 485 -2133 486 -2132
rect 597 -2133 598 -2132
rect 618 -2133 619 -2132
rect 905 -2133 906 -2132
rect 1381 -2133 1382 -2132
rect 1388 -2133 1389 -2132
rect 1479 -2133 1480 -2132
rect 1493 -2133 1494 -2132
rect 30 -2135 31 -2134
rect 618 -2135 619 -2134
rect 621 -2135 622 -2134
rect 646 -2135 647 -2134
rect 660 -2135 661 -2134
rect 1248 -2135 1249 -2134
rect 1360 -2135 1361 -2134
rect 1381 -2135 1382 -2134
rect 1458 -2135 1459 -2134
rect 1479 -2135 1480 -2134
rect 1486 -2135 1487 -2134
rect 1640 -2135 1641 -2134
rect 51 -2137 52 -2136
rect 478 -2137 479 -2136
rect 485 -2137 486 -2136
rect 730 -2137 731 -2136
rect 1059 -2137 1060 -2136
rect 1486 -2137 1487 -2136
rect 240 -2139 241 -2138
rect 275 -2139 276 -2138
rect 387 -2139 388 -2138
rect 422 -2139 423 -2138
rect 429 -2139 430 -2138
rect 968 -2139 969 -2138
rect 1059 -2139 1060 -2138
rect 1087 -2139 1088 -2138
rect 1318 -2139 1319 -2138
rect 1360 -2139 1361 -2138
rect 170 -2141 171 -2140
rect 240 -2141 241 -2140
rect 247 -2141 248 -2140
rect 261 -2141 262 -2140
rect 387 -2141 388 -2140
rect 443 -2141 444 -2140
rect 457 -2141 458 -2140
rect 884 -2141 885 -2140
rect 968 -2141 969 -2140
rect 1003 -2141 1004 -2140
rect 1087 -2141 1088 -2140
rect 1094 -2141 1095 -2140
rect 1304 -2141 1305 -2140
rect 1318 -2141 1319 -2140
rect 93 -2143 94 -2142
rect 457 -2143 458 -2142
rect 464 -2143 465 -2142
rect 590 -2143 591 -2142
rect 653 -2143 654 -2142
rect 730 -2143 731 -2142
rect 814 -2143 815 -2142
rect 1003 -2143 1004 -2142
rect 1094 -2143 1095 -2142
rect 1143 -2143 1144 -2142
rect 1297 -2143 1298 -2142
rect 1304 -2143 1305 -2142
rect 93 -2145 94 -2144
rect 996 -2145 997 -2144
rect 1122 -2145 1123 -2144
rect 1143 -2145 1144 -2144
rect 1283 -2145 1284 -2144
rect 1297 -2145 1298 -2144
rect 58 -2147 59 -2146
rect 996 -2147 997 -2146
rect 1241 -2147 1242 -2146
rect 1283 -2147 1284 -2146
rect 58 -2149 59 -2148
rect 625 -2149 626 -2148
rect 670 -2149 671 -2148
rect 1458 -2149 1459 -2148
rect 170 -2151 171 -2150
rect 1689 -2151 1690 -2150
rect 219 -2153 220 -2152
rect 443 -2153 444 -2152
rect 471 -2153 472 -2152
rect 908 -2153 909 -2152
rect 1185 -2153 1186 -2152
rect 1241 -2153 1242 -2152
rect 198 -2155 199 -2154
rect 219 -2155 220 -2154
rect 226 -2155 227 -2154
rect 247 -2155 248 -2154
rect 362 -2155 363 -2154
rect 464 -2155 465 -2154
rect 520 -2155 521 -2154
rect 646 -2155 647 -2154
rect 751 -2155 752 -2154
rect 1122 -2155 1123 -2154
rect 1164 -2155 1165 -2154
rect 1185 -2155 1186 -2154
rect 198 -2157 199 -2156
rect 1755 -2157 1756 -2156
rect 226 -2159 227 -2158
rect 1430 -2159 1431 -2158
rect 229 -2161 230 -2160
rect 471 -2161 472 -2160
rect 513 -2161 514 -2160
rect 520 -2161 521 -2160
rect 583 -2161 584 -2160
rect 653 -2161 654 -2160
rect 751 -2161 752 -2160
rect 828 -2161 829 -2160
rect 1150 -2161 1151 -2160
rect 1164 -2161 1165 -2160
rect 65 -2163 66 -2162
rect 513 -2163 514 -2162
rect 583 -2163 584 -2162
rect 695 -2163 696 -2162
rect 1136 -2163 1137 -2162
rect 1150 -2163 1151 -2162
rect 65 -2165 66 -2164
rect 1024 -2165 1025 -2164
rect 415 -2167 416 -2166
rect 978 -2167 979 -2166
rect 982 -2167 983 -2166
rect 1136 -2167 1137 -2166
rect 600 -2169 601 -2168
rect 1430 -2169 1431 -2168
rect 625 -2171 626 -2170
rect 891 -2171 892 -2170
rect 961 -2171 962 -2170
rect 1024 -2171 1025 -2170
rect 695 -2173 696 -2172
rect 709 -2173 710 -2172
rect 849 -2173 850 -2172
rect 891 -2173 892 -2172
rect 975 -2173 976 -2172
rect 982 -2173 983 -2172
rect 282 -2175 283 -2174
rect 709 -2175 710 -2174
rect 849 -2175 850 -2174
rect 863 -2175 864 -2174
rect 282 -2177 283 -2176
rect 401 -2177 402 -2176
rect 639 -2177 640 -2176
rect 863 -2177 864 -2176
rect 72 -2179 73 -2178
rect 639 -2179 640 -2178
rect 702 -2179 703 -2178
rect 961 -2179 962 -2178
rect 72 -2181 73 -2180
rect 933 -2181 934 -2180
rect 380 -2183 381 -2182
rect 401 -2183 402 -2182
rect 702 -2183 703 -2182
rect 793 -2183 794 -2182
rect 933 -2183 934 -2182
rect 1269 -2183 1270 -2182
rect 380 -2185 381 -2184
rect 450 -2185 451 -2184
rect 450 -2187 451 -2186
rect 660 -2187 661 -2186
rect 30 -2198 31 -2197
rect 450 -2198 451 -2197
rect 453 -2198 454 -2197
rect 653 -2198 654 -2197
rect 688 -2198 689 -2197
rect 793 -2198 794 -2197
rect 796 -2198 797 -2197
rect 1395 -2198 1396 -2197
rect 1640 -2198 1641 -2197
rect 1706 -2198 1707 -2197
rect 1752 -2198 1753 -2197
rect 1766 -2198 1767 -2197
rect 44 -2200 45 -2199
rect 870 -2200 871 -2199
rect 873 -2200 874 -2199
rect 1465 -2200 1466 -2199
rect 1640 -2200 1641 -2199
rect 1696 -2200 1697 -2199
rect 51 -2202 52 -2201
rect 72 -2202 73 -2201
rect 89 -2202 90 -2201
rect 103 -2202 104 -2201
rect 117 -2202 118 -2201
rect 1444 -2202 1445 -2201
rect 1465 -2202 1466 -2201
rect 1514 -2202 1515 -2201
rect 1682 -2202 1683 -2201
rect 1713 -2202 1714 -2201
rect 51 -2204 52 -2203
rect 394 -2204 395 -2203
rect 408 -2204 409 -2203
rect 779 -2204 780 -2203
rect 786 -2204 787 -2203
rect 814 -2204 815 -2203
rect 828 -2204 829 -2203
rect 1367 -2204 1368 -2203
rect 1514 -2204 1515 -2203
rect 1549 -2204 1550 -2203
rect 1682 -2204 1683 -2203
rect 1717 -2204 1718 -2203
rect 58 -2206 59 -2205
rect 957 -2206 958 -2205
rect 978 -2206 979 -2205
rect 1423 -2206 1424 -2205
rect 1549 -2206 1550 -2205
rect 1591 -2206 1592 -2205
rect 1696 -2206 1697 -2205
rect 1738 -2206 1739 -2205
rect 58 -2208 59 -2207
rect 639 -2208 640 -2207
rect 691 -2208 692 -2207
rect 716 -2208 717 -2207
rect 723 -2208 724 -2207
rect 1346 -2208 1347 -2207
rect 1423 -2208 1424 -2207
rect 1472 -2208 1473 -2207
rect 1738 -2208 1739 -2207
rect 1759 -2208 1760 -2207
rect 65 -2210 66 -2209
rect 604 -2210 605 -2209
rect 607 -2210 608 -2209
rect 807 -2210 808 -2209
rect 814 -2210 815 -2209
rect 821 -2210 822 -2209
rect 828 -2210 829 -2209
rect 842 -2210 843 -2209
rect 852 -2210 853 -2209
rect 1031 -2210 1032 -2209
rect 1118 -2210 1119 -2209
rect 1661 -2210 1662 -2209
rect 68 -2212 69 -2211
rect 562 -2212 563 -2211
rect 611 -2212 612 -2211
rect 747 -2212 748 -2211
rect 758 -2212 759 -2211
rect 1129 -2212 1130 -2211
rect 1146 -2212 1147 -2211
rect 1731 -2212 1732 -2211
rect 72 -2214 73 -2213
rect 121 -2214 122 -2213
rect 131 -2214 132 -2213
rect 1017 -2214 1018 -2213
rect 1031 -2214 1032 -2213
rect 1101 -2214 1102 -2213
rect 1129 -2214 1130 -2213
rect 1206 -2214 1207 -2213
rect 1227 -2214 1228 -2213
rect 1731 -2214 1732 -2213
rect 89 -2216 90 -2215
rect 177 -2216 178 -2215
rect 184 -2216 185 -2215
rect 604 -2216 605 -2215
rect 618 -2216 619 -2215
rect 1367 -2216 1368 -2215
rect 1507 -2216 1508 -2215
rect 1661 -2216 1662 -2215
rect 93 -2218 94 -2217
rect 884 -2218 885 -2217
rect 891 -2218 892 -2217
rect 936 -2218 937 -2217
rect 999 -2218 1000 -2217
rect 1276 -2218 1277 -2217
rect 1335 -2218 1336 -2217
rect 1654 -2218 1655 -2217
rect 96 -2220 97 -2219
rect 1122 -2220 1123 -2219
rect 1192 -2220 1193 -2219
rect 1395 -2220 1396 -2219
rect 96 -2222 97 -2221
rect 184 -2222 185 -2221
rect 226 -2222 227 -2221
rect 415 -2222 416 -2221
rect 450 -2222 451 -2221
rect 646 -2222 647 -2221
rect 695 -2222 696 -2221
rect 730 -2222 731 -2221
rect 733 -2222 734 -2221
rect 1703 -2222 1704 -2221
rect 121 -2224 122 -2223
rect 233 -2224 234 -2223
rect 236 -2224 237 -2223
rect 793 -2224 794 -2223
rect 807 -2224 808 -2223
rect 835 -2224 836 -2223
rect 842 -2224 843 -2223
rect 877 -2224 878 -2223
rect 884 -2224 885 -2223
rect 1066 -2224 1067 -2223
rect 1122 -2224 1123 -2223
rect 1745 -2224 1746 -2223
rect 142 -2226 143 -2225
rect 145 -2226 146 -2225
rect 152 -2226 153 -2225
rect 1444 -2226 1445 -2225
rect 142 -2228 143 -2227
rect 625 -2228 626 -2227
rect 639 -2228 640 -2227
rect 1038 -2228 1039 -2227
rect 1066 -2228 1067 -2227
rect 1755 -2228 1756 -2227
rect 170 -2230 171 -2229
rect 317 -2230 318 -2229
rect 362 -2230 363 -2229
rect 873 -2230 874 -2229
rect 877 -2230 878 -2229
rect 905 -2230 906 -2229
rect 933 -2230 934 -2229
rect 1283 -2230 1284 -2229
rect 1346 -2230 1347 -2229
rect 1402 -2230 1403 -2229
rect 170 -2232 171 -2231
rect 523 -2232 524 -2231
rect 569 -2232 570 -2231
rect 695 -2232 696 -2231
rect 702 -2232 703 -2231
rect 1633 -2232 1634 -2231
rect 177 -2234 178 -2233
rect 205 -2234 206 -2233
rect 229 -2234 230 -2233
rect 954 -2234 955 -2233
rect 999 -2234 1000 -2233
rect 1717 -2234 1718 -2233
rect 205 -2236 206 -2235
rect 345 -2236 346 -2235
rect 464 -2236 465 -2235
rect 611 -2236 612 -2235
rect 618 -2236 619 -2235
rect 674 -2236 675 -2235
rect 702 -2236 703 -2235
rect 1213 -2236 1214 -2235
rect 1227 -2236 1228 -2235
rect 1297 -2236 1298 -2235
rect 1339 -2236 1340 -2235
rect 1402 -2236 1403 -2235
rect 1626 -2236 1627 -2235
rect 1633 -2236 1634 -2235
rect 100 -2238 101 -2237
rect 674 -2238 675 -2237
rect 716 -2238 717 -2237
rect 751 -2238 752 -2237
rect 772 -2238 773 -2237
rect 1507 -2238 1508 -2237
rect 1612 -2238 1613 -2237
rect 1626 -2238 1627 -2237
rect 44 -2240 45 -2239
rect 772 -2240 773 -2239
rect 786 -2240 787 -2239
rect 800 -2240 801 -2239
rect 821 -2240 822 -2239
rect 849 -2240 850 -2239
rect 891 -2240 892 -2239
rect 1045 -2240 1046 -2239
rect 1206 -2240 1207 -2239
rect 1318 -2240 1319 -2239
rect 1339 -2240 1340 -2239
rect 1388 -2240 1389 -2239
rect 1542 -2240 1543 -2239
rect 1612 -2240 1613 -2239
rect 100 -2242 101 -2241
rect 135 -2242 136 -2241
rect 191 -2242 192 -2241
rect 345 -2242 346 -2241
rect 422 -2242 423 -2241
rect 464 -2242 465 -2241
rect 471 -2242 472 -2241
rect 562 -2242 563 -2241
rect 569 -2242 570 -2241
rect 1059 -2242 1060 -2241
rect 1213 -2242 1214 -2241
rect 1255 -2242 1256 -2241
rect 1276 -2242 1277 -2241
rect 1486 -2242 1487 -2241
rect 1542 -2242 1543 -2241
rect 1577 -2242 1578 -2241
rect 135 -2244 136 -2243
rect 1619 -2244 1620 -2243
rect 191 -2246 192 -2245
rect 240 -2246 241 -2245
rect 268 -2246 269 -2245
rect 555 -2246 556 -2245
rect 586 -2246 587 -2245
rect 1192 -2246 1193 -2245
rect 1237 -2246 1238 -2245
rect 1675 -2246 1676 -2245
rect 107 -2248 108 -2247
rect 240 -2248 241 -2247
rect 271 -2248 272 -2247
rect 541 -2248 542 -2247
rect 548 -2248 549 -2247
rect 555 -2248 556 -2247
rect 646 -2248 647 -2247
rect 660 -2248 661 -2247
rect 730 -2248 731 -2247
rect 1472 -2248 1473 -2247
rect 1486 -2248 1487 -2247
rect 1521 -2248 1522 -2247
rect 1577 -2248 1578 -2247
rect 1703 -2248 1704 -2247
rect 107 -2250 108 -2249
rect 163 -2250 164 -2249
rect 233 -2250 234 -2249
rect 261 -2250 262 -2249
rect 282 -2250 283 -2249
rect 775 -2250 776 -2249
rect 800 -2250 801 -2249
rect 926 -2250 927 -2249
rect 933 -2250 934 -2249
rect 968 -2250 969 -2249
rect 1003 -2250 1004 -2249
rect 1101 -2250 1102 -2249
rect 1255 -2250 1256 -2249
rect 1430 -2250 1431 -2249
rect 1521 -2250 1522 -2249
rect 1724 -2250 1725 -2249
rect 114 -2252 115 -2251
rect 261 -2252 262 -2251
rect 282 -2252 283 -2251
rect 436 -2252 437 -2251
rect 506 -2252 507 -2251
rect 733 -2252 734 -2251
rect 737 -2252 738 -2251
rect 779 -2252 780 -2251
rect 835 -2252 836 -2251
rect 961 -2252 962 -2251
rect 1003 -2252 1004 -2251
rect 1150 -2252 1151 -2251
rect 1283 -2252 1284 -2251
rect 1416 -2252 1417 -2251
rect 163 -2254 164 -2253
rect 632 -2254 633 -2253
rect 656 -2254 657 -2253
rect 660 -2254 661 -2253
rect 747 -2254 748 -2253
rect 1675 -2254 1676 -2253
rect 215 -2256 216 -2255
rect 737 -2256 738 -2255
rect 751 -2256 752 -2255
rect 856 -2256 857 -2255
rect 898 -2256 899 -2255
rect 961 -2256 962 -2255
rect 1010 -2256 1011 -2255
rect 1360 -2256 1361 -2255
rect 1388 -2256 1389 -2255
rect 1598 -2256 1599 -2255
rect 156 -2258 157 -2257
rect 898 -2258 899 -2257
rect 905 -2258 906 -2257
rect 919 -2258 920 -2257
rect 926 -2258 927 -2257
rect 1024 -2258 1025 -2257
rect 1038 -2258 1039 -2257
rect 1199 -2258 1200 -2257
rect 1290 -2258 1291 -2257
rect 1724 -2258 1725 -2257
rect 156 -2260 157 -2259
rect 534 -2260 535 -2259
rect 541 -2260 542 -2259
rect 982 -2260 983 -2259
rect 1010 -2260 1011 -2259
rect 1108 -2260 1109 -2259
rect 1199 -2260 1200 -2259
rect 1234 -2260 1235 -2259
rect 1290 -2260 1291 -2259
rect 1374 -2260 1375 -2259
rect 1584 -2260 1585 -2259
rect 1598 -2260 1599 -2259
rect 128 -2262 129 -2261
rect 1584 -2262 1585 -2261
rect 40 -2264 41 -2263
rect 128 -2264 129 -2263
rect 289 -2264 290 -2263
rect 625 -2264 626 -2263
rect 761 -2264 762 -2263
rect 919 -2264 920 -2263
rect 982 -2264 983 -2263
rect 1136 -2264 1137 -2263
rect 1297 -2264 1298 -2263
rect 1381 -2264 1382 -2263
rect 173 -2266 174 -2265
rect 1381 -2266 1382 -2265
rect 173 -2268 174 -2267
rect 901 -2268 902 -2267
rect 1013 -2268 1014 -2267
rect 1024 -2268 1025 -2267
rect 1045 -2268 1046 -2267
rect 1094 -2268 1095 -2267
rect 1108 -2268 1109 -2267
rect 1668 -2268 1669 -2267
rect 289 -2270 290 -2269
rect 380 -2270 381 -2269
rect 436 -2270 437 -2269
rect 513 -2270 514 -2269
rect 520 -2270 521 -2269
rect 1619 -2270 1620 -2269
rect 1668 -2270 1669 -2269
rect 1710 -2270 1711 -2269
rect 114 -2272 115 -2271
rect 513 -2272 514 -2271
rect 548 -2272 549 -2271
rect 681 -2272 682 -2271
rect 849 -2272 850 -2271
rect 1654 -2272 1655 -2271
rect 149 -2274 150 -2273
rect 520 -2274 521 -2273
rect 681 -2274 682 -2273
rect 831 -2274 832 -2273
rect 1017 -2274 1018 -2273
rect 1052 -2274 1053 -2273
rect 1059 -2274 1060 -2273
rect 1185 -2274 1186 -2273
rect 1318 -2274 1319 -2273
rect 1458 -2274 1459 -2273
rect 1591 -2274 1592 -2273
rect 1710 -2274 1711 -2273
rect 149 -2276 150 -2275
rect 254 -2276 255 -2275
rect 296 -2276 297 -2275
rect 359 -2276 360 -2275
rect 478 -2276 479 -2275
rect 632 -2276 633 -2275
rect 1052 -2276 1053 -2275
rect 1080 -2276 1081 -2275
rect 1094 -2276 1095 -2275
rect 1563 -2276 1564 -2275
rect 219 -2278 220 -2277
rect 380 -2278 381 -2277
rect 478 -2278 479 -2277
rect 597 -2278 598 -2277
rect 1073 -2278 1074 -2277
rect 1150 -2278 1151 -2277
rect 1185 -2278 1186 -2277
rect 1248 -2278 1249 -2277
rect 1332 -2278 1333 -2277
rect 1416 -2278 1417 -2277
rect 1458 -2278 1459 -2277
rect 1479 -2278 1480 -2277
rect 1556 -2278 1557 -2277
rect 1563 -2278 1564 -2277
rect 145 -2280 146 -2279
rect 219 -2280 220 -2279
rect 247 -2280 248 -2279
rect 254 -2280 255 -2279
rect 296 -2280 297 -2279
rect 709 -2280 710 -2279
rect 1073 -2280 1074 -2279
rect 1164 -2280 1165 -2279
rect 1353 -2280 1354 -2279
rect 1430 -2280 1431 -2279
rect 1479 -2280 1480 -2279
rect 1528 -2280 1529 -2279
rect 1556 -2280 1557 -2279
rect 1605 -2280 1606 -2279
rect 79 -2282 80 -2281
rect 247 -2282 248 -2281
rect 303 -2282 304 -2281
rect 394 -2282 395 -2281
rect 457 -2282 458 -2281
rect 709 -2282 710 -2281
rect 968 -2282 969 -2281
rect 1353 -2282 1354 -2281
rect 1360 -2282 1361 -2281
rect 1409 -2282 1410 -2281
rect 1493 -2282 1494 -2281
rect 1605 -2282 1606 -2281
rect 79 -2284 80 -2283
rect 198 -2284 199 -2283
rect 310 -2284 311 -2283
rect 975 -2284 976 -2283
rect 1136 -2284 1137 -2283
rect 1262 -2284 1263 -2283
rect 1304 -2284 1305 -2283
rect 1528 -2284 1529 -2283
rect 86 -2286 87 -2285
rect 457 -2286 458 -2285
rect 492 -2286 493 -2285
rect 534 -2286 535 -2285
rect 723 -2286 724 -2285
rect 1304 -2286 1305 -2285
rect 1374 -2286 1375 -2285
rect 1451 -2286 1452 -2285
rect 1493 -2286 1494 -2285
rect 1689 -2286 1690 -2285
rect 138 -2288 139 -2287
rect 303 -2288 304 -2287
rect 310 -2288 311 -2287
rect 485 -2288 486 -2287
rect 499 -2288 500 -2287
rect 506 -2288 507 -2287
rect 653 -2288 654 -2287
rect 1689 -2288 1690 -2287
rect 198 -2290 199 -2289
rect 1104 -2290 1105 -2289
rect 1157 -2290 1158 -2289
rect 1248 -2290 1249 -2289
rect 1269 -2290 1270 -2289
rect 1451 -2290 1452 -2289
rect 317 -2292 318 -2291
rect 688 -2292 689 -2291
rect 744 -2292 745 -2291
rect 1409 -2292 1410 -2291
rect 324 -2294 325 -2293
rect 856 -2294 857 -2293
rect 975 -2294 976 -2293
rect 989 -2294 990 -2293
rect 1083 -2294 1084 -2293
rect 1262 -2294 1263 -2293
rect 324 -2296 325 -2295
rect 366 -2296 367 -2295
rect 373 -2296 374 -2295
rect 485 -2296 486 -2295
rect 499 -2296 500 -2295
rect 863 -2296 864 -2295
rect 989 -2296 990 -2295
rect 1311 -2296 1312 -2295
rect 275 -2298 276 -2297
rect 366 -2298 367 -2297
rect 429 -2298 430 -2297
rect 492 -2298 493 -2297
rect 744 -2298 745 -2297
rect 947 -2298 948 -2297
rect 954 -2298 955 -2297
rect 1311 -2298 1312 -2297
rect 212 -2300 213 -2299
rect 275 -2300 276 -2299
rect 331 -2300 332 -2299
rect 422 -2300 423 -2299
rect 429 -2300 430 -2299
rect 705 -2300 706 -2299
rect 863 -2300 864 -2299
rect 1143 -2300 1144 -2299
rect 1157 -2300 1158 -2299
rect 1220 -2300 1221 -2299
rect 331 -2302 332 -2301
rect 1115 -2302 1116 -2301
rect 1164 -2302 1165 -2301
rect 1241 -2302 1242 -2301
rect 338 -2304 339 -2303
rect 373 -2304 374 -2303
rect 415 -2304 416 -2303
rect 705 -2304 706 -2303
rect 912 -2304 913 -2303
rect 1115 -2304 1116 -2303
rect 1171 -2304 1172 -2303
rect 1220 -2304 1221 -2303
rect 1241 -2304 1242 -2303
rect 1325 -2304 1326 -2303
rect 338 -2306 339 -2305
rect 401 -2306 402 -2305
rect 912 -2306 913 -2305
rect 940 -2306 941 -2305
rect 947 -2306 948 -2305
rect 1332 -2306 1333 -2305
rect 352 -2308 353 -2307
rect 401 -2308 402 -2307
rect 940 -2308 941 -2307
rect 1087 -2308 1088 -2307
rect 1143 -2308 1144 -2307
rect 1325 -2308 1326 -2307
rect 352 -2310 353 -2309
rect 576 -2310 577 -2309
rect 1087 -2310 1088 -2309
rect 1178 -2310 1179 -2309
rect 359 -2312 360 -2311
rect 387 -2312 388 -2311
rect 576 -2312 577 -2311
rect 667 -2312 668 -2311
rect 996 -2312 997 -2311
rect 1178 -2312 1179 -2311
rect 387 -2314 388 -2313
rect 527 -2314 528 -2313
rect 667 -2314 668 -2313
rect 765 -2314 766 -2313
rect 996 -2314 997 -2313
rect 1269 -2314 1270 -2313
rect 443 -2316 444 -2315
rect 765 -2316 766 -2315
rect 443 -2318 444 -2317
rect 583 -2318 584 -2317
rect 471 -2320 472 -2319
rect 583 -2320 584 -2319
rect 527 -2322 528 -2321
rect 870 -2322 871 -2321
rect 51 -2333 52 -2332
rect 180 -2333 181 -2332
rect 215 -2333 216 -2332
rect 975 -2333 976 -2332
rect 982 -2333 983 -2332
rect 996 -2333 997 -2332
rect 999 -2333 1000 -2332
rect 1486 -2333 1487 -2332
rect 1514 -2333 1515 -2332
rect 1538 -2333 1539 -2332
rect 1605 -2333 1606 -2332
rect 1706 -2333 1707 -2332
rect 51 -2335 52 -2334
rect 226 -2335 227 -2334
rect 443 -2335 444 -2334
rect 824 -2335 825 -2334
rect 856 -2335 857 -2334
rect 971 -2335 972 -2334
rect 982 -2335 983 -2334
rect 1045 -2335 1046 -2334
rect 1076 -2335 1077 -2334
rect 1437 -2335 1438 -2334
rect 1493 -2335 1494 -2334
rect 1514 -2335 1515 -2334
rect 1605 -2335 1606 -2334
rect 1675 -2335 1676 -2334
rect 79 -2337 80 -2336
rect 702 -2337 703 -2336
rect 733 -2337 734 -2336
rect 1122 -2337 1123 -2336
rect 1171 -2337 1172 -2336
rect 1451 -2337 1452 -2336
rect 1612 -2337 1613 -2336
rect 1675 -2337 1676 -2336
rect 79 -2339 80 -2338
rect 93 -2339 94 -2338
rect 100 -2339 101 -2338
rect 1125 -2339 1126 -2338
rect 1171 -2339 1172 -2338
rect 1178 -2339 1179 -2338
rect 1244 -2339 1245 -2338
rect 1668 -2339 1669 -2338
rect 86 -2341 87 -2340
rect 1689 -2341 1690 -2340
rect 86 -2343 87 -2342
rect 128 -2343 129 -2342
rect 135 -2343 136 -2342
rect 380 -2343 381 -2342
rect 415 -2343 416 -2342
rect 443 -2343 444 -2342
rect 450 -2343 451 -2342
rect 583 -2343 584 -2342
rect 597 -2343 598 -2342
rect 656 -2343 657 -2342
rect 660 -2343 661 -2342
rect 677 -2343 678 -2342
rect 684 -2343 685 -2342
rect 1584 -2343 1585 -2342
rect 93 -2345 94 -2344
rect 422 -2345 423 -2344
rect 464 -2345 465 -2344
rect 467 -2345 468 -2344
rect 492 -2345 493 -2344
rect 730 -2345 731 -2344
rect 775 -2345 776 -2344
rect 1395 -2345 1396 -2344
rect 1437 -2345 1438 -2344
rect 1472 -2345 1473 -2344
rect 100 -2347 101 -2346
rect 261 -2347 262 -2346
rect 345 -2347 346 -2346
rect 450 -2347 451 -2346
rect 457 -2347 458 -2346
rect 492 -2347 493 -2346
rect 502 -2347 503 -2346
rect 534 -2347 535 -2346
rect 548 -2347 549 -2346
rect 583 -2347 584 -2346
rect 597 -2347 598 -2346
rect 642 -2347 643 -2346
rect 691 -2347 692 -2346
rect 1563 -2347 1564 -2346
rect 65 -2349 66 -2348
rect 457 -2349 458 -2348
rect 464 -2349 465 -2348
rect 485 -2349 486 -2348
rect 527 -2349 528 -2348
rect 1045 -2349 1046 -2348
rect 1080 -2349 1081 -2348
rect 1528 -2349 1529 -2348
rect 1556 -2349 1557 -2348
rect 1563 -2349 1564 -2348
rect 65 -2351 66 -2350
rect 149 -2351 150 -2350
rect 163 -2351 164 -2350
rect 236 -2351 237 -2350
rect 240 -2351 241 -2350
rect 380 -2351 381 -2350
rect 422 -2351 423 -2350
rect 730 -2351 731 -2350
rect 733 -2351 734 -2350
rect 1472 -2351 1473 -2350
rect 1521 -2351 1522 -2350
rect 1556 -2351 1557 -2350
rect 96 -2353 97 -2352
rect 1528 -2353 1529 -2352
rect 107 -2355 108 -2354
rect 534 -2355 535 -2354
rect 548 -2355 549 -2354
rect 562 -2355 563 -2354
rect 569 -2355 570 -2354
rect 653 -2355 654 -2354
rect 800 -2355 801 -2354
rect 1195 -2355 1196 -2354
rect 1304 -2355 1305 -2354
rect 1626 -2355 1627 -2354
rect 107 -2357 108 -2356
rect 138 -2357 139 -2356
rect 149 -2357 150 -2356
rect 205 -2357 206 -2356
rect 212 -2357 213 -2356
rect 415 -2357 416 -2356
rect 467 -2357 468 -2356
rect 485 -2357 486 -2356
rect 530 -2357 531 -2356
rect 975 -2357 976 -2356
rect 989 -2357 990 -2356
rect 1584 -2357 1585 -2356
rect 58 -2359 59 -2358
rect 205 -2359 206 -2358
rect 212 -2359 213 -2358
rect 1192 -2359 1193 -2358
rect 1304 -2359 1305 -2358
rect 1353 -2359 1354 -2358
rect 1384 -2359 1385 -2358
rect 1570 -2359 1571 -2358
rect 114 -2361 115 -2360
rect 499 -2361 500 -2360
rect 576 -2361 577 -2360
rect 660 -2361 661 -2360
rect 779 -2361 780 -2360
rect 800 -2361 801 -2360
rect 856 -2361 857 -2360
rect 1633 -2361 1634 -2360
rect 44 -2363 45 -2362
rect 576 -2363 577 -2362
rect 618 -2363 619 -2362
rect 688 -2363 689 -2362
rect 695 -2363 696 -2362
rect 779 -2363 780 -2362
rect 863 -2363 864 -2362
rect 1146 -2363 1147 -2362
rect 1178 -2363 1179 -2362
rect 1307 -2363 1308 -2362
rect 1314 -2363 1315 -2362
rect 1696 -2363 1697 -2362
rect 114 -2365 115 -2364
rect 359 -2365 360 -2364
rect 432 -2365 433 -2364
rect 618 -2365 619 -2364
rect 625 -2365 626 -2364
rect 1486 -2365 1487 -2364
rect 1521 -2365 1522 -2364
rect 1654 -2365 1655 -2364
rect 117 -2367 118 -2366
rect 233 -2367 234 -2366
rect 240 -2367 241 -2366
rect 387 -2367 388 -2366
rect 471 -2367 472 -2366
rect 562 -2367 563 -2366
rect 590 -2367 591 -2366
rect 625 -2367 626 -2366
rect 632 -2367 633 -2366
rect 747 -2367 748 -2366
rect 863 -2367 864 -2366
rect 1143 -2367 1144 -2366
rect 1283 -2367 1284 -2366
rect 1353 -2367 1354 -2366
rect 1388 -2367 1389 -2366
rect 1493 -2367 1494 -2366
rect 1570 -2367 1571 -2366
rect 1598 -2367 1599 -2366
rect 128 -2369 129 -2368
rect 156 -2369 157 -2368
rect 163 -2369 164 -2368
rect 835 -2369 836 -2368
rect 870 -2369 871 -2368
rect 877 -2369 878 -2368
rect 898 -2369 899 -2368
rect 1682 -2369 1683 -2368
rect 135 -2371 136 -2370
rect 604 -2371 605 -2370
rect 632 -2371 633 -2370
rect 947 -2371 948 -2370
rect 954 -2371 955 -2370
rect 1661 -2371 1662 -2370
rect 142 -2373 143 -2372
rect 877 -2373 878 -2372
rect 898 -2373 899 -2372
rect 1311 -2373 1312 -2372
rect 1332 -2373 1333 -2372
rect 1647 -2373 1648 -2372
rect 142 -2375 143 -2374
rect 478 -2375 479 -2374
rect 499 -2375 500 -2374
rect 1083 -2375 1084 -2374
rect 1097 -2375 1098 -2374
rect 1255 -2375 1256 -2374
rect 1388 -2375 1389 -2374
rect 1409 -2375 1410 -2374
rect 1451 -2375 1452 -2374
rect 1549 -2375 1550 -2374
rect 1598 -2375 1599 -2374
rect 1703 -2375 1704 -2374
rect 170 -2377 171 -2376
rect 520 -2377 521 -2376
rect 541 -2377 542 -2376
rect 747 -2377 748 -2376
rect 828 -2377 829 -2376
rect 835 -2377 836 -2376
rect 873 -2377 874 -2376
rect 1500 -2377 1501 -2376
rect 170 -2379 171 -2378
rect 198 -2379 199 -2378
rect 215 -2379 216 -2378
rect 674 -2379 675 -2378
rect 688 -2379 689 -2378
rect 723 -2379 724 -2378
rect 828 -2379 829 -2378
rect 1066 -2379 1067 -2378
rect 1080 -2379 1081 -2378
rect 1101 -2379 1102 -2378
rect 1108 -2379 1109 -2378
rect 1500 -2379 1501 -2378
rect 156 -2381 157 -2380
rect 674 -2381 675 -2380
rect 695 -2381 696 -2380
rect 709 -2381 710 -2380
rect 723 -2381 724 -2380
rect 814 -2381 815 -2380
rect 919 -2381 920 -2380
rect 989 -2381 990 -2380
rect 996 -2381 997 -2380
rect 1031 -2381 1032 -2380
rect 1066 -2381 1067 -2380
rect 1150 -2381 1151 -2380
rect 1192 -2381 1193 -2380
rect 1283 -2381 1284 -2380
rect 1395 -2381 1396 -2380
rect 1423 -2381 1424 -2380
rect 198 -2383 199 -2382
rect 296 -2383 297 -2382
rect 345 -2383 346 -2382
rect 373 -2383 374 -2382
rect 387 -2383 388 -2382
rect 474 -2383 475 -2382
rect 478 -2383 479 -2382
rect 681 -2383 682 -2382
rect 709 -2383 710 -2382
rect 716 -2383 717 -2382
rect 793 -2383 794 -2382
rect 1101 -2383 1102 -2382
rect 1122 -2383 1123 -2382
rect 1129 -2383 1130 -2382
rect 1143 -2383 1144 -2382
rect 1199 -2383 1200 -2382
rect 1255 -2383 1256 -2382
rect 1339 -2383 1340 -2382
rect 1374 -2383 1375 -2382
rect 1423 -2383 1424 -2382
rect 226 -2385 227 -2384
rect 247 -2385 248 -2384
rect 254 -2385 255 -2384
rect 261 -2385 262 -2384
rect 268 -2385 269 -2384
rect 569 -2385 570 -2384
rect 590 -2385 591 -2384
rect 611 -2385 612 -2384
rect 639 -2385 640 -2384
rect 1619 -2385 1620 -2384
rect 184 -2387 185 -2386
rect 247 -2387 248 -2386
rect 254 -2387 255 -2386
rect 401 -2387 402 -2386
rect 471 -2387 472 -2386
rect 765 -2387 766 -2386
rect 786 -2387 787 -2386
rect 793 -2387 794 -2386
rect 919 -2387 920 -2386
rect 1213 -2387 1214 -2386
rect 1339 -2387 1340 -2386
rect 1360 -2387 1361 -2386
rect 1374 -2387 1375 -2386
rect 1444 -2387 1445 -2386
rect 184 -2389 185 -2388
rect 849 -2389 850 -2388
rect 901 -2389 902 -2388
rect 1444 -2389 1445 -2388
rect 268 -2391 269 -2390
rect 429 -2391 430 -2390
rect 513 -2391 514 -2390
rect 1150 -2391 1151 -2390
rect 1185 -2391 1186 -2390
rect 1213 -2391 1214 -2390
rect 1360 -2391 1361 -2390
rect 1402 -2391 1403 -2390
rect 1409 -2391 1410 -2390
rect 1479 -2391 1480 -2390
rect 282 -2393 283 -2392
rect 513 -2393 514 -2392
rect 520 -2393 521 -2392
rect 744 -2393 745 -2392
rect 786 -2393 787 -2392
rect 821 -2393 822 -2392
rect 901 -2393 902 -2392
rect 1430 -2393 1431 -2392
rect 1479 -2393 1480 -2392
rect 1577 -2393 1578 -2392
rect 282 -2395 283 -2394
rect 289 -2395 290 -2394
rect 296 -2395 297 -2394
rect 772 -2395 773 -2394
rect 814 -2395 815 -2394
rect 849 -2395 850 -2394
rect 926 -2395 927 -2394
rect 954 -2395 955 -2394
rect 957 -2395 958 -2394
rect 1332 -2395 1333 -2394
rect 1346 -2395 1347 -2394
rect 1402 -2395 1403 -2394
rect 1430 -2395 1431 -2394
rect 1591 -2395 1592 -2394
rect 173 -2397 174 -2396
rect 289 -2397 290 -2396
rect 303 -2397 304 -2396
rect 401 -2397 402 -2396
rect 555 -2397 556 -2396
rect 611 -2397 612 -2396
rect 646 -2397 647 -2396
rect 765 -2397 766 -2396
rect 772 -2397 773 -2396
rect 852 -2397 853 -2396
rect 884 -2397 885 -2396
rect 926 -2397 927 -2396
rect 933 -2397 934 -2396
rect 947 -2397 948 -2396
rect 971 -2397 972 -2396
rect 1458 -2397 1459 -2396
rect 1577 -2397 1578 -2396
rect 1738 -2397 1739 -2396
rect 177 -2399 178 -2398
rect 303 -2399 304 -2398
rect 310 -2399 311 -2398
rect 555 -2399 556 -2398
rect 604 -2399 605 -2398
rect 751 -2399 752 -2398
rect 821 -2399 822 -2398
rect 1731 -2399 1732 -2398
rect 58 -2401 59 -2400
rect 310 -2401 311 -2400
rect 338 -2401 339 -2400
rect 373 -2401 374 -2400
rect 653 -2401 654 -2400
rect 667 -2401 668 -2400
rect 716 -2401 717 -2400
rect 737 -2401 738 -2400
rect 744 -2401 745 -2400
rect 912 -2401 913 -2400
rect 1024 -2401 1025 -2400
rect 1108 -2401 1109 -2400
rect 1115 -2401 1116 -2400
rect 1591 -2401 1592 -2400
rect 177 -2403 178 -2402
rect 436 -2403 437 -2402
rect 667 -2403 668 -2402
rect 807 -2403 808 -2402
rect 842 -2403 843 -2402
rect 884 -2403 885 -2402
rect 891 -2403 892 -2402
rect 912 -2403 913 -2402
rect 1017 -2403 1018 -2402
rect 1024 -2403 1025 -2402
rect 1031 -2403 1032 -2402
rect 1227 -2403 1228 -2402
rect 1318 -2403 1319 -2402
rect 1346 -2403 1347 -2402
rect 1458 -2403 1459 -2402
rect 1542 -2403 1543 -2402
rect 191 -2405 192 -2404
rect 338 -2405 339 -2404
rect 352 -2405 353 -2404
rect 646 -2405 647 -2404
rect 737 -2405 738 -2404
rect 810 -2405 811 -2404
rect 842 -2405 843 -2404
rect 1003 -2405 1004 -2404
rect 1038 -2405 1039 -2404
rect 1129 -2405 1130 -2404
rect 1136 -2405 1137 -2404
rect 1227 -2405 1228 -2404
rect 1535 -2405 1536 -2404
rect 1542 -2405 1543 -2404
rect 191 -2407 192 -2406
rect 331 -2407 332 -2406
rect 359 -2407 360 -2406
rect 366 -2407 367 -2406
rect 436 -2407 437 -2406
rect 506 -2407 507 -2406
rect 751 -2407 752 -2406
rect 968 -2407 969 -2406
rect 1003 -2407 1004 -2406
rect 1290 -2407 1291 -2406
rect 219 -2409 220 -2408
rect 352 -2409 353 -2408
rect 506 -2409 507 -2408
rect 541 -2409 542 -2408
rect 758 -2409 759 -2408
rect 1017 -2409 1018 -2408
rect 1038 -2409 1039 -2408
rect 1059 -2409 1060 -2408
rect 1115 -2409 1116 -2408
rect 1157 -2409 1158 -2408
rect 1185 -2409 1186 -2408
rect 1325 -2409 1326 -2408
rect 219 -2411 220 -2410
rect 317 -2411 318 -2410
rect 324 -2411 325 -2410
rect 366 -2411 367 -2410
rect 758 -2411 759 -2410
rect 1234 -2411 1235 -2410
rect 1290 -2411 1291 -2410
rect 1381 -2411 1382 -2410
rect 121 -2413 122 -2412
rect 317 -2413 318 -2412
rect 324 -2413 325 -2412
rect 807 -2413 808 -2412
rect 891 -2413 892 -2412
rect 1010 -2413 1011 -2412
rect 1059 -2413 1060 -2412
rect 1087 -2413 1088 -2412
rect 1136 -2413 1137 -2412
rect 1717 -2413 1718 -2412
rect 72 -2415 73 -2414
rect 121 -2415 122 -2414
rect 331 -2415 332 -2414
rect 614 -2415 615 -2414
rect 961 -2415 962 -2414
rect 1010 -2415 1011 -2414
rect 1073 -2415 1074 -2414
rect 1087 -2415 1088 -2414
rect 1157 -2415 1158 -2414
rect 1164 -2415 1165 -2414
rect 1199 -2415 1200 -2414
rect 1206 -2415 1207 -2414
rect 1220 -2415 1221 -2414
rect 1318 -2415 1319 -2414
rect 1325 -2415 1326 -2414
rect 1335 -2415 1336 -2414
rect 1381 -2415 1382 -2414
rect 1416 -2415 1417 -2414
rect 72 -2417 73 -2416
rect 1094 -2417 1095 -2416
rect 1164 -2417 1165 -2416
rect 1724 -2417 1725 -2416
rect 537 -2419 538 -2418
rect 1220 -2419 1221 -2418
rect 1234 -2419 1235 -2418
rect 1241 -2419 1242 -2418
rect 1276 -2419 1277 -2418
rect 1416 -2419 1417 -2418
rect 933 -2421 934 -2420
rect 1073 -2421 1074 -2420
rect 1206 -2421 1207 -2420
rect 1297 -2421 1298 -2420
rect 940 -2423 941 -2422
rect 1094 -2423 1095 -2422
rect 1241 -2423 1242 -2422
rect 1549 -2423 1550 -2422
rect 940 -2425 941 -2424
rect 1710 -2425 1711 -2424
rect 961 -2427 962 -2426
rect 1052 -2427 1053 -2426
rect 1262 -2427 1263 -2426
rect 1276 -2427 1277 -2426
rect 705 -2429 706 -2428
rect 1052 -2429 1053 -2428
rect 1262 -2429 1263 -2428
rect 1269 -2429 1270 -2428
rect 408 -2431 409 -2430
rect 705 -2431 706 -2430
rect 1269 -2431 1270 -2430
rect 1367 -2431 1368 -2430
rect 275 -2433 276 -2432
rect 408 -2433 409 -2432
rect 1367 -2433 1368 -2432
rect 1465 -2433 1466 -2432
rect 275 -2435 276 -2434
rect 394 -2435 395 -2434
rect 1465 -2435 1466 -2434
rect 1507 -2435 1508 -2434
rect 394 -2437 395 -2436
rect 845 -2437 846 -2436
rect 1507 -2437 1508 -2436
rect 1640 -2437 1641 -2436
rect 44 -2448 45 -2447
rect 163 -2448 164 -2447
rect 184 -2448 185 -2447
rect 649 -2448 650 -2447
rect 681 -2448 682 -2447
rect 744 -2448 745 -2447
rect 754 -2448 755 -2447
rect 779 -2448 780 -2447
rect 786 -2448 787 -2447
rect 873 -2448 874 -2447
rect 912 -2448 913 -2447
rect 1696 -2448 1697 -2447
rect 86 -2450 87 -2449
rect 177 -2450 178 -2449
rect 240 -2450 241 -2449
rect 859 -2450 860 -2449
rect 870 -2450 871 -2449
rect 912 -2450 913 -2449
rect 957 -2450 958 -2449
rect 996 -2450 997 -2449
rect 1062 -2450 1063 -2449
rect 1612 -2450 1613 -2449
rect 1675 -2450 1676 -2449
rect 1731 -2450 1732 -2449
rect 86 -2452 87 -2451
rect 597 -2452 598 -2451
rect 611 -2452 612 -2451
rect 1521 -2452 1522 -2451
rect 1528 -2452 1529 -2451
rect 1678 -2452 1679 -2451
rect 100 -2454 101 -2453
rect 240 -2454 241 -2453
rect 257 -2454 258 -2453
rect 681 -2454 682 -2453
rect 688 -2454 689 -2453
rect 740 -2454 741 -2453
rect 779 -2454 780 -2453
rect 800 -2454 801 -2453
rect 807 -2454 808 -2453
rect 954 -2454 955 -2453
rect 971 -2454 972 -2453
rect 1584 -2454 1585 -2453
rect 1605 -2454 1606 -2453
rect 1724 -2454 1725 -2453
rect 107 -2456 108 -2455
rect 870 -2456 871 -2455
rect 891 -2456 892 -2455
rect 996 -2456 997 -2455
rect 1076 -2456 1077 -2455
rect 1346 -2456 1347 -2455
rect 1367 -2456 1368 -2455
rect 1521 -2456 1522 -2455
rect 1538 -2456 1539 -2455
rect 1563 -2456 1564 -2455
rect 1577 -2456 1578 -2455
rect 1738 -2456 1739 -2455
rect 72 -2458 73 -2457
rect 107 -2458 108 -2457
rect 142 -2458 143 -2457
rect 166 -2458 167 -2457
rect 180 -2458 181 -2457
rect 800 -2458 801 -2457
rect 821 -2458 822 -2457
rect 1605 -2458 1606 -2457
rect 142 -2460 143 -2459
rect 628 -2460 629 -2459
rect 642 -2460 643 -2459
rect 1192 -2460 1193 -2459
rect 1227 -2460 1228 -2459
rect 1367 -2460 1368 -2459
rect 1381 -2460 1382 -2459
rect 1479 -2460 1480 -2459
rect 1500 -2460 1501 -2459
rect 1577 -2460 1578 -2459
rect 152 -2462 153 -2461
rect 1290 -2462 1291 -2461
rect 1300 -2462 1301 -2461
rect 1430 -2462 1431 -2461
rect 1458 -2462 1459 -2461
rect 1619 -2462 1620 -2461
rect 282 -2464 283 -2463
rect 551 -2464 552 -2463
rect 562 -2464 563 -2463
rect 611 -2464 612 -2463
rect 702 -2464 703 -2463
rect 828 -2464 829 -2463
rect 842 -2464 843 -2463
rect 1073 -2464 1074 -2463
rect 1115 -2464 1116 -2463
rect 1227 -2464 1228 -2463
rect 1244 -2464 1245 -2463
rect 1304 -2464 1305 -2463
rect 1311 -2464 1312 -2463
rect 1528 -2464 1529 -2463
rect 1556 -2464 1557 -2463
rect 1710 -2464 1711 -2463
rect 261 -2466 262 -2465
rect 282 -2466 283 -2465
rect 296 -2466 297 -2465
rect 471 -2466 472 -2465
rect 492 -2466 493 -2465
rect 562 -2466 563 -2465
rect 593 -2466 594 -2465
rect 1136 -2466 1137 -2465
rect 1157 -2466 1158 -2465
rect 1640 -2466 1641 -2465
rect 226 -2468 227 -2467
rect 261 -2468 262 -2467
rect 296 -2468 297 -2467
rect 352 -2468 353 -2467
rect 411 -2468 412 -2467
rect 464 -2468 465 -2467
rect 502 -2468 503 -2467
rect 1661 -2468 1662 -2467
rect 93 -2470 94 -2469
rect 352 -2470 353 -2469
rect 422 -2470 423 -2469
rect 464 -2470 465 -2469
rect 506 -2470 507 -2469
rect 688 -2470 689 -2469
rect 716 -2470 717 -2469
rect 828 -2470 829 -2469
rect 845 -2470 846 -2469
rect 1269 -2470 1270 -2469
rect 1276 -2470 1277 -2469
rect 1346 -2470 1347 -2469
rect 1395 -2470 1396 -2469
rect 1682 -2470 1683 -2469
rect 65 -2472 66 -2471
rect 93 -2472 94 -2471
rect 226 -2472 227 -2471
rect 317 -2472 318 -2471
rect 324 -2472 325 -2471
rect 499 -2472 500 -2471
rect 506 -2472 507 -2471
rect 684 -2472 685 -2471
rect 730 -2472 731 -2471
rect 1094 -2472 1095 -2471
rect 1129 -2472 1130 -2471
rect 1192 -2472 1193 -2471
rect 1199 -2472 1200 -2471
rect 1311 -2472 1312 -2471
rect 1314 -2472 1315 -2471
rect 1486 -2472 1487 -2471
rect 1507 -2472 1508 -2471
rect 1689 -2472 1690 -2471
rect 65 -2474 66 -2473
rect 79 -2474 80 -2473
rect 100 -2474 101 -2473
rect 317 -2474 318 -2473
rect 324 -2474 325 -2473
rect 408 -2474 409 -2473
rect 422 -2474 423 -2473
rect 485 -2474 486 -2473
rect 513 -2474 514 -2473
rect 541 -2474 542 -2473
rect 583 -2474 584 -2473
rect 716 -2474 717 -2473
rect 751 -2474 752 -2473
rect 1458 -2474 1459 -2473
rect 1465 -2474 1466 -2473
rect 1584 -2474 1585 -2473
rect 58 -2476 59 -2475
rect 485 -2476 486 -2475
rect 513 -2476 514 -2475
rect 590 -2476 591 -2475
rect 597 -2476 598 -2475
rect 653 -2476 654 -2475
rect 751 -2476 752 -2475
rect 1563 -2476 1564 -2475
rect 58 -2478 59 -2477
rect 632 -2478 633 -2477
rect 765 -2478 766 -2477
rect 891 -2478 892 -2477
rect 919 -2478 920 -2477
rect 1269 -2478 1270 -2477
rect 1276 -2478 1277 -2477
rect 1451 -2478 1452 -2477
rect 1507 -2478 1508 -2477
rect 1570 -2478 1571 -2477
rect 79 -2480 80 -2479
rect 345 -2480 346 -2479
rect 401 -2480 402 -2479
rect 765 -2480 766 -2479
rect 793 -2480 794 -2479
rect 807 -2480 808 -2479
rect 852 -2480 853 -2479
rect 1122 -2480 1123 -2479
rect 1129 -2480 1130 -2479
rect 1598 -2480 1599 -2479
rect 121 -2482 122 -2481
rect 401 -2482 402 -2481
rect 408 -2482 409 -2481
rect 898 -2482 899 -2481
rect 929 -2482 930 -2481
rect 1500 -2482 1501 -2481
rect 1514 -2482 1515 -2481
rect 1668 -2482 1669 -2481
rect 121 -2484 122 -2483
rect 128 -2484 129 -2483
rect 215 -2484 216 -2483
rect 1486 -2484 1487 -2483
rect 128 -2486 129 -2485
rect 149 -2486 150 -2485
rect 303 -2486 304 -2485
rect 432 -2486 433 -2485
rect 436 -2486 437 -2485
rect 492 -2486 493 -2485
rect 520 -2486 521 -2485
rect 674 -2486 675 -2485
rect 677 -2486 678 -2485
rect 1570 -2486 1571 -2485
rect 75 -2488 76 -2487
rect 436 -2488 437 -2487
rect 450 -2488 451 -2487
rect 653 -2488 654 -2487
rect 674 -2488 675 -2487
rect 786 -2488 787 -2487
rect 877 -2488 878 -2487
rect 898 -2488 899 -2487
rect 1024 -2488 1025 -2487
rect 1094 -2488 1095 -2487
rect 1167 -2488 1168 -2487
rect 1409 -2488 1410 -2487
rect 1416 -2488 1417 -2487
rect 1514 -2488 1515 -2487
rect 149 -2490 150 -2489
rect 184 -2490 185 -2489
rect 303 -2490 304 -2489
rect 387 -2490 388 -2489
rect 429 -2490 430 -2489
rect 1626 -2490 1627 -2489
rect 310 -2492 311 -2491
rect 373 -2492 374 -2491
rect 387 -2492 388 -2491
rect 457 -2492 458 -2491
rect 474 -2492 475 -2491
rect 499 -2492 500 -2491
rect 520 -2492 521 -2491
rect 961 -2492 962 -2491
rect 982 -2492 983 -2491
rect 1024 -2492 1025 -2491
rect 1031 -2492 1032 -2491
rect 1304 -2492 1305 -2491
rect 1332 -2492 1333 -2491
rect 1409 -2492 1410 -2491
rect 1472 -2492 1473 -2491
rect 1598 -2492 1599 -2491
rect 103 -2494 104 -2493
rect 373 -2494 374 -2493
rect 432 -2494 433 -2493
rect 1717 -2494 1718 -2493
rect 313 -2496 314 -2495
rect 359 -2496 360 -2495
rect 443 -2496 444 -2495
rect 450 -2496 451 -2495
rect 527 -2496 528 -2495
rect 569 -2496 570 -2495
rect 576 -2496 577 -2495
rect 1416 -2496 1417 -2495
rect 247 -2498 248 -2497
rect 359 -2498 360 -2497
rect 366 -2498 367 -2497
rect 527 -2498 528 -2497
rect 541 -2498 542 -2497
rect 723 -2498 724 -2497
rect 877 -2498 878 -2497
rect 894 -2498 895 -2497
rect 933 -2498 934 -2497
rect 961 -2498 962 -2497
rect 1031 -2498 1032 -2497
rect 1188 -2498 1189 -2497
rect 1199 -2498 1200 -2497
rect 1255 -2498 1256 -2497
rect 1290 -2498 1291 -2497
rect 1388 -2498 1389 -2497
rect 1395 -2498 1396 -2497
rect 1549 -2498 1550 -2497
rect 219 -2500 220 -2499
rect 247 -2500 248 -2499
rect 275 -2500 276 -2499
rect 366 -2500 367 -2499
rect 415 -2500 416 -2499
rect 443 -2500 444 -2499
rect 534 -2500 535 -2499
rect 723 -2500 724 -2499
rect 810 -2500 811 -2499
rect 1388 -2500 1389 -2499
rect 1542 -2500 1543 -2499
rect 1549 -2500 1550 -2499
rect 198 -2502 199 -2501
rect 219 -2502 220 -2501
rect 275 -2502 276 -2501
rect 733 -2502 734 -2501
rect 884 -2502 885 -2501
rect 919 -2502 920 -2501
rect 933 -2502 934 -2501
rect 1297 -2502 1298 -2501
rect 1325 -2502 1326 -2501
rect 1332 -2502 1333 -2501
rect 1339 -2502 1340 -2501
rect 1654 -2502 1655 -2501
rect 173 -2504 174 -2503
rect 198 -2504 199 -2503
rect 331 -2504 332 -2503
rect 457 -2504 458 -2503
rect 534 -2504 535 -2503
rect 849 -2504 850 -2503
rect 1038 -2504 1039 -2503
rect 1157 -2504 1158 -2503
rect 1178 -2504 1179 -2503
rect 1297 -2504 1298 -2503
rect 1339 -2504 1340 -2503
rect 1580 -2504 1581 -2503
rect 51 -2506 52 -2505
rect 849 -2506 850 -2505
rect 1003 -2506 1004 -2505
rect 1038 -2506 1039 -2505
rect 1052 -2506 1053 -2505
rect 1136 -2506 1137 -2505
rect 1185 -2506 1186 -2505
rect 1381 -2506 1382 -2505
rect 1444 -2506 1445 -2505
rect 1542 -2506 1543 -2505
rect 51 -2508 52 -2507
rect 170 -2508 171 -2507
rect 268 -2508 269 -2507
rect 331 -2508 332 -2507
rect 338 -2508 339 -2507
rect 341 -2508 342 -2507
rect 415 -2508 416 -2507
rect 530 -2508 531 -2507
rect 548 -2508 549 -2507
rect 583 -2508 584 -2507
rect 590 -2508 591 -2507
rect 639 -2508 640 -2507
rect 663 -2508 664 -2507
rect 1178 -2508 1179 -2507
rect 1185 -2508 1186 -2507
rect 1423 -2508 1424 -2507
rect 268 -2510 269 -2509
rect 289 -2510 290 -2509
rect 338 -2510 339 -2509
rect 380 -2510 381 -2509
rect 548 -2510 549 -2509
rect 1115 -2510 1116 -2509
rect 1206 -2510 1207 -2509
rect 1444 -2510 1445 -2509
rect 163 -2512 164 -2511
rect 1206 -2512 1207 -2511
rect 1209 -2512 1210 -2511
rect 1451 -2512 1452 -2511
rect 289 -2514 290 -2513
rect 446 -2514 447 -2513
rect 569 -2514 570 -2513
rect 604 -2514 605 -2513
rect 625 -2514 626 -2513
rect 632 -2514 633 -2513
rect 695 -2514 696 -2513
rect 793 -2514 794 -2513
rect 821 -2514 822 -2513
rect 1423 -2514 1424 -2513
rect 156 -2516 157 -2515
rect 625 -2516 626 -2515
rect 733 -2516 734 -2515
rect 1706 -2516 1707 -2515
rect 156 -2518 157 -2517
rect 747 -2518 748 -2517
rect 835 -2518 836 -2517
rect 884 -2518 885 -2517
rect 926 -2518 927 -2517
rect 1003 -2518 1004 -2517
rect 1010 -2518 1011 -2517
rect 1052 -2518 1053 -2517
rect 1059 -2518 1060 -2517
rect 1073 -2518 1074 -2517
rect 1083 -2518 1084 -2517
rect 1122 -2518 1123 -2517
rect 1213 -2518 1214 -2517
rect 1472 -2518 1473 -2517
rect 341 -2520 342 -2519
rect 380 -2520 381 -2519
rect 555 -2520 556 -2519
rect 695 -2520 696 -2519
rect 709 -2520 710 -2519
rect 835 -2520 836 -2519
rect 926 -2520 927 -2519
rect 982 -2520 983 -2519
rect 1059 -2520 1060 -2519
rect 1150 -2520 1151 -2519
rect 1213 -2520 1214 -2519
rect 1318 -2520 1319 -2519
rect 1360 -2520 1361 -2519
rect 1465 -2520 1466 -2519
rect 576 -2522 577 -2521
rect 737 -2522 738 -2521
rect 863 -2522 864 -2521
rect 1318 -2522 1319 -2521
rect 135 -2524 136 -2523
rect 737 -2524 738 -2523
rect 863 -2524 864 -2523
rect 905 -2524 906 -2523
rect 975 -2524 976 -2523
rect 1010 -2524 1011 -2523
rect 1066 -2524 1067 -2523
rect 1430 -2524 1431 -2523
rect 135 -2526 136 -2525
rect 191 -2526 192 -2525
rect 394 -2526 395 -2525
rect 1066 -2526 1067 -2525
rect 1087 -2526 1088 -2525
rect 1150 -2526 1151 -2525
rect 1220 -2526 1221 -2525
rect 1325 -2526 1326 -2525
rect 114 -2528 115 -2527
rect 191 -2528 192 -2527
rect 394 -2528 395 -2527
rect 667 -2528 668 -2527
rect 705 -2528 706 -2527
rect 905 -2528 906 -2527
rect 1087 -2528 1088 -2527
rect 1633 -2528 1634 -2527
rect 114 -2530 115 -2529
rect 618 -2530 619 -2529
rect 660 -2530 661 -2529
rect 747 -2530 748 -2529
rect 814 -2530 815 -2529
rect 975 -2530 976 -2529
rect 1090 -2530 1091 -2529
rect 1556 -2530 1557 -2529
rect 68 -2532 69 -2531
rect 618 -2532 619 -2531
rect 660 -2532 661 -2531
rect 1374 -2532 1375 -2531
rect 604 -2534 605 -2533
rect 940 -2534 941 -2533
rect 1220 -2534 1221 -2533
rect 1591 -2534 1592 -2533
rect 478 -2536 479 -2535
rect 940 -2536 941 -2535
rect 1248 -2536 1249 -2535
rect 1647 -2536 1648 -2535
rect 205 -2538 206 -2537
rect 478 -2538 479 -2537
rect 667 -2538 668 -2537
rect 901 -2538 902 -2537
rect 1143 -2538 1144 -2537
rect 1248 -2538 1249 -2537
rect 1255 -2538 1256 -2537
rect 1353 -2538 1354 -2537
rect 1374 -2538 1375 -2537
rect 1493 -2538 1494 -2537
rect 1535 -2538 1536 -2537
rect 1591 -2538 1592 -2537
rect 205 -2540 206 -2539
rect 968 -2540 969 -2539
rect 1045 -2540 1046 -2539
rect 1143 -2540 1144 -2539
rect 1234 -2540 1235 -2539
rect 1353 -2540 1354 -2539
rect 1402 -2540 1403 -2539
rect 1493 -2540 1494 -2539
rect 709 -2542 710 -2541
rect 789 -2542 790 -2541
rect 814 -2542 815 -2541
rect 824 -2542 825 -2541
rect 856 -2542 857 -2541
rect 968 -2542 969 -2541
rect 989 -2542 990 -2541
rect 1045 -2542 1046 -2541
rect 1171 -2542 1172 -2541
rect 1234 -2542 1235 -2541
rect 1262 -2542 1263 -2541
rect 1360 -2542 1361 -2541
rect 1437 -2542 1438 -2541
rect 1535 -2542 1536 -2541
rect 555 -2544 556 -2543
rect 824 -2544 825 -2543
rect 856 -2544 857 -2543
rect 954 -2544 955 -2543
rect 989 -2544 990 -2543
rect 1108 -2544 1109 -2543
rect 1164 -2544 1165 -2543
rect 1262 -2544 1263 -2543
rect 1283 -2544 1284 -2543
rect 1402 -2544 1403 -2543
rect 758 -2546 759 -2545
rect 1283 -2546 1284 -2545
rect 730 -2548 731 -2547
rect 758 -2548 759 -2547
rect 1017 -2548 1018 -2547
rect 1108 -2548 1109 -2547
rect 1164 -2548 1165 -2547
rect 1479 -2548 1480 -2547
rect 772 -2550 773 -2549
rect 1017 -2550 1018 -2549
rect 1101 -2550 1102 -2549
rect 1171 -2550 1172 -2549
rect 1195 -2550 1196 -2549
rect 1437 -2550 1438 -2549
rect 646 -2552 647 -2551
rect 772 -2552 773 -2551
rect 1080 -2552 1081 -2551
rect 1101 -2552 1102 -2551
rect 345 -2554 346 -2553
rect 646 -2554 647 -2553
rect 1080 -2554 1081 -2553
rect 1241 -2554 1242 -2553
rect 72 -2565 73 -2564
rect 478 -2565 479 -2564
rect 513 -2565 514 -2564
rect 786 -2565 787 -2564
rect 789 -2565 790 -2564
rect 1430 -2565 1431 -2564
rect 1678 -2565 1679 -2564
rect 1731 -2565 1732 -2564
rect 75 -2567 76 -2566
rect 1563 -2567 1564 -2566
rect 1703 -2567 1704 -2566
rect 1738 -2567 1739 -2566
rect 79 -2569 80 -2568
rect 446 -2569 447 -2568
rect 460 -2569 461 -2568
rect 604 -2569 605 -2568
rect 618 -2569 619 -2568
rect 1185 -2569 1186 -2568
rect 1430 -2569 1431 -2568
rect 1500 -2569 1501 -2568
rect 1563 -2569 1564 -2568
rect 1626 -2569 1627 -2568
rect 1703 -2569 1704 -2568
rect 1717 -2569 1718 -2568
rect 100 -2571 101 -2570
rect 849 -2571 850 -2570
rect 873 -2571 874 -2570
rect 1241 -2571 1242 -2570
rect 1500 -2571 1501 -2570
rect 1584 -2571 1585 -2570
rect 1626 -2571 1627 -2570
rect 1661 -2571 1662 -2570
rect 100 -2573 101 -2572
rect 135 -2573 136 -2572
rect 149 -2573 150 -2572
rect 1066 -2573 1067 -2572
rect 1080 -2573 1081 -2572
rect 1129 -2573 1130 -2572
rect 1178 -2573 1179 -2572
rect 1185 -2573 1186 -2572
rect 1374 -2573 1375 -2572
rect 1584 -2573 1585 -2572
rect 128 -2575 129 -2574
rect 149 -2575 150 -2574
rect 170 -2575 171 -2574
rect 401 -2575 402 -2574
rect 429 -2575 430 -2574
rect 856 -2575 857 -2574
rect 873 -2575 874 -2574
rect 1262 -2575 1263 -2574
rect 1374 -2575 1375 -2574
rect 1423 -2575 1424 -2574
rect 58 -2577 59 -2576
rect 429 -2577 430 -2576
rect 432 -2577 433 -2576
rect 527 -2577 528 -2576
rect 548 -2577 549 -2576
rect 1458 -2577 1459 -2576
rect 58 -2579 59 -2578
rect 324 -2579 325 -2578
rect 373 -2579 374 -2578
rect 376 -2579 377 -2578
rect 436 -2579 437 -2578
rect 548 -2579 549 -2578
rect 555 -2579 556 -2578
rect 786 -2579 787 -2578
rect 800 -2579 801 -2578
rect 1423 -2579 1424 -2578
rect 1458 -2579 1459 -2578
rect 1689 -2579 1690 -2578
rect 44 -2581 45 -2580
rect 555 -2581 556 -2580
rect 576 -2581 577 -2580
rect 824 -2581 825 -2580
rect 845 -2581 846 -2580
rect 1654 -2581 1655 -2580
rect 44 -2583 45 -2582
rect 89 -2583 90 -2582
rect 121 -2583 122 -2582
rect 170 -2583 171 -2582
rect 201 -2583 202 -2582
rect 1416 -2583 1417 -2582
rect 1542 -2583 1543 -2582
rect 1654 -2583 1655 -2582
rect 128 -2585 129 -2584
rect 394 -2585 395 -2584
rect 436 -2585 437 -2584
rect 478 -2585 479 -2584
rect 506 -2585 507 -2584
rect 849 -2585 850 -2584
rect 856 -2585 857 -2584
rect 891 -2585 892 -2584
rect 926 -2585 927 -2584
rect 1647 -2585 1648 -2584
rect 135 -2587 136 -2586
rect 663 -2587 664 -2586
rect 670 -2587 671 -2586
rect 1682 -2587 1683 -2586
rect 152 -2589 153 -2588
rect 1689 -2589 1690 -2588
rect 240 -2591 241 -2590
rect 576 -2591 577 -2590
rect 593 -2591 594 -2590
rect 611 -2591 612 -2590
rect 625 -2591 626 -2590
rect 1696 -2591 1697 -2590
rect 240 -2593 241 -2592
rect 261 -2593 262 -2592
rect 268 -2593 269 -2592
rect 527 -2593 528 -2592
rect 600 -2593 601 -2592
rect 1143 -2593 1144 -2592
rect 1178 -2593 1179 -2592
rect 1227 -2593 1228 -2592
rect 1262 -2593 1263 -2592
rect 1304 -2593 1305 -2592
rect 1395 -2593 1396 -2592
rect 1661 -2593 1662 -2592
rect 1696 -2593 1697 -2592
rect 1724 -2593 1725 -2592
rect 226 -2595 227 -2594
rect 268 -2595 269 -2594
rect 303 -2595 304 -2594
rect 394 -2595 395 -2594
rect 401 -2595 402 -2594
rect 891 -2595 892 -2594
rect 905 -2595 906 -2594
rect 926 -2595 927 -2594
rect 954 -2595 955 -2594
rect 1451 -2595 1452 -2594
rect 212 -2597 213 -2596
rect 226 -2597 227 -2596
rect 233 -2597 234 -2596
rect 303 -2597 304 -2596
rect 324 -2597 325 -2596
rect 380 -2597 381 -2596
rect 506 -2597 507 -2596
rect 590 -2597 591 -2596
rect 604 -2597 605 -2596
rect 674 -2597 675 -2596
rect 730 -2597 731 -2596
rect 940 -2597 941 -2596
rect 1034 -2597 1035 -2596
rect 1129 -2597 1130 -2596
rect 1213 -2597 1214 -2596
rect 1304 -2597 1305 -2596
rect 1395 -2597 1396 -2596
rect 1437 -2597 1438 -2596
rect 1451 -2597 1452 -2596
rect 1521 -2597 1522 -2596
rect 117 -2599 118 -2598
rect 940 -2599 941 -2598
rect 1038 -2599 1039 -2598
rect 1083 -2599 1084 -2598
rect 1087 -2599 1088 -2598
rect 1283 -2599 1284 -2598
rect 1416 -2599 1417 -2598
rect 1493 -2599 1494 -2598
rect 163 -2601 164 -2600
rect 590 -2601 591 -2600
rect 611 -2601 612 -2600
rect 695 -2601 696 -2600
rect 733 -2601 734 -2600
rect 1682 -2601 1683 -2600
rect 163 -2603 164 -2602
rect 551 -2603 552 -2602
rect 632 -2603 633 -2602
rect 646 -2603 647 -2602
rect 649 -2603 650 -2602
rect 1353 -2603 1354 -2602
rect 1437 -2603 1438 -2602
rect 1514 -2603 1515 -2602
rect 68 -2605 69 -2604
rect 1353 -2605 1354 -2604
rect 1493 -2605 1494 -2604
rect 1549 -2605 1550 -2604
rect 166 -2607 167 -2606
rect 674 -2607 675 -2606
rect 695 -2607 696 -2606
rect 838 -2607 839 -2606
rect 884 -2607 885 -2606
rect 929 -2607 930 -2606
rect 1010 -2607 1011 -2606
rect 1038 -2607 1039 -2606
rect 1059 -2607 1060 -2606
rect 1640 -2607 1641 -2606
rect 166 -2609 167 -2608
rect 1570 -2609 1571 -2608
rect 198 -2611 199 -2610
rect 233 -2611 234 -2610
rect 254 -2611 255 -2610
rect 282 -2611 283 -2610
rect 296 -2611 297 -2610
rect 905 -2611 906 -2610
rect 1003 -2611 1004 -2610
rect 1010 -2611 1011 -2610
rect 1059 -2611 1060 -2610
rect 1101 -2611 1102 -2610
rect 1122 -2611 1123 -2610
rect 1167 -2611 1168 -2610
rect 1227 -2611 1228 -2610
rect 1248 -2611 1249 -2610
rect 1276 -2611 1277 -2610
rect 1570 -2611 1571 -2610
rect 65 -2613 66 -2612
rect 1003 -2613 1004 -2612
rect 1066 -2613 1067 -2612
rect 1339 -2613 1340 -2612
rect 1507 -2613 1508 -2612
rect 1640 -2613 1641 -2612
rect 156 -2615 157 -2614
rect 296 -2615 297 -2614
rect 373 -2615 374 -2614
rect 422 -2615 423 -2614
rect 520 -2615 521 -2614
rect 1090 -2615 1091 -2614
rect 1094 -2615 1095 -2614
rect 1241 -2615 1242 -2614
rect 1276 -2615 1277 -2614
rect 1325 -2615 1326 -2614
rect 1507 -2615 1508 -2614
rect 1710 -2615 1711 -2614
rect 156 -2617 157 -2616
rect 345 -2617 346 -2616
rect 376 -2617 377 -2616
rect 422 -2617 423 -2616
rect 520 -2617 521 -2616
rect 562 -2617 563 -2616
rect 632 -2617 633 -2616
rect 716 -2617 717 -2616
rect 733 -2617 734 -2616
rect 758 -2617 759 -2616
rect 772 -2617 773 -2616
rect 954 -2617 955 -2616
rect 957 -2617 958 -2616
rect 1248 -2617 1249 -2616
rect 1283 -2617 1284 -2616
rect 1318 -2617 1319 -2616
rect 1325 -2617 1326 -2616
rect 1381 -2617 1382 -2616
rect 1514 -2617 1515 -2616
rect 1591 -2617 1592 -2616
rect 212 -2619 213 -2618
rect 359 -2619 360 -2618
rect 380 -2619 381 -2618
rect 387 -2619 388 -2618
rect 464 -2619 465 -2618
rect 758 -2619 759 -2618
rect 772 -2619 773 -2618
rect 807 -2619 808 -2618
rect 821 -2619 822 -2618
rect 1220 -2619 1221 -2618
rect 1255 -2619 1256 -2618
rect 1381 -2619 1382 -2618
rect 1549 -2619 1550 -2618
rect 1612 -2619 1613 -2618
rect 191 -2621 192 -2620
rect 359 -2621 360 -2620
rect 492 -2621 493 -2620
rect 562 -2621 563 -2620
rect 639 -2621 640 -2620
rect 691 -2621 692 -2620
rect 716 -2621 717 -2620
rect 1108 -2621 1109 -2620
rect 1122 -2621 1123 -2620
rect 1150 -2621 1151 -2620
rect 1157 -2621 1158 -2620
rect 1220 -2621 1221 -2620
rect 1255 -2621 1256 -2620
rect 1297 -2621 1298 -2620
rect 1318 -2621 1319 -2620
rect 1360 -2621 1361 -2620
rect 1612 -2621 1613 -2620
rect 1633 -2621 1634 -2620
rect 184 -2623 185 -2622
rect 191 -2623 192 -2622
rect 254 -2623 255 -2622
rect 257 -2623 258 -2622
rect 261 -2623 262 -2622
rect 275 -2623 276 -2622
rect 282 -2623 283 -2622
rect 499 -2623 500 -2622
rect 646 -2623 647 -2622
rect 1164 -2623 1165 -2622
rect 1199 -2623 1200 -2622
rect 1339 -2623 1340 -2622
rect 142 -2625 143 -2624
rect 184 -2625 185 -2624
rect 275 -2625 276 -2624
rect 408 -2625 409 -2624
rect 418 -2625 419 -2624
rect 499 -2625 500 -2624
rect 660 -2625 661 -2624
rect 814 -2625 815 -2624
rect 821 -2625 822 -2624
rect 828 -2625 829 -2624
rect 884 -2625 885 -2624
rect 933 -2625 934 -2624
rect 957 -2625 958 -2624
rect 1542 -2625 1543 -2624
rect 107 -2627 108 -2626
rect 408 -2627 409 -2626
rect 457 -2627 458 -2626
rect 492 -2627 493 -2626
rect 569 -2627 570 -2626
rect 828 -2627 829 -2626
rect 894 -2627 895 -2626
rect 1521 -2627 1522 -2626
rect 107 -2629 108 -2628
rect 205 -2629 206 -2628
rect 310 -2629 311 -2628
rect 457 -2629 458 -2628
rect 471 -2629 472 -2628
rect 569 -2629 570 -2628
rect 744 -2629 745 -2628
rect 765 -2629 766 -2628
rect 779 -2629 780 -2628
rect 814 -2629 815 -2628
rect 933 -2629 934 -2628
rect 961 -2629 962 -2628
rect 989 -2629 990 -2628
rect 1164 -2629 1165 -2628
rect 1199 -2629 1200 -2628
rect 1206 -2629 1207 -2628
rect 1269 -2629 1270 -2628
rect 1633 -2629 1634 -2628
rect 72 -2631 73 -2630
rect 765 -2631 766 -2630
rect 803 -2631 804 -2630
rect 989 -2631 990 -2630
rect 1024 -2631 1025 -2630
rect 1108 -2631 1109 -2630
rect 1150 -2631 1151 -2630
rect 1675 -2631 1676 -2630
rect 142 -2633 143 -2632
rect 667 -2633 668 -2632
rect 747 -2633 748 -2632
rect 1647 -2633 1648 -2632
rect 177 -2635 178 -2634
rect 471 -2635 472 -2634
rect 485 -2635 486 -2634
rect 639 -2635 640 -2634
rect 653 -2635 654 -2634
rect 667 -2635 668 -2634
rect 751 -2635 752 -2634
rect 1486 -2635 1487 -2634
rect 1556 -2635 1557 -2634
rect 1675 -2635 1676 -2634
rect 51 -2637 52 -2636
rect 177 -2637 178 -2636
rect 205 -2637 206 -2636
rect 289 -2637 290 -2636
rect 317 -2637 318 -2636
rect 660 -2637 661 -2636
rect 751 -2637 752 -2636
rect 1143 -2637 1144 -2636
rect 1157 -2637 1158 -2636
rect 1171 -2637 1172 -2636
rect 1206 -2637 1207 -2636
rect 1234 -2637 1235 -2636
rect 1269 -2637 1270 -2636
rect 1311 -2637 1312 -2636
rect 1486 -2637 1487 -2636
rect 1668 -2637 1669 -2636
rect 51 -2639 52 -2638
rect 541 -2639 542 -2638
rect 597 -2639 598 -2638
rect 779 -2639 780 -2638
rect 807 -2639 808 -2638
rect 835 -2639 836 -2638
rect 947 -2639 948 -2638
rect 961 -2639 962 -2638
rect 982 -2639 983 -2638
rect 1171 -2639 1172 -2638
rect 1297 -2639 1298 -2638
rect 1402 -2639 1403 -2638
rect 1556 -2639 1557 -2638
rect 1619 -2639 1620 -2638
rect 121 -2641 122 -2640
rect 597 -2641 598 -2640
rect 625 -2641 626 -2640
rect 1619 -2641 1620 -2640
rect 247 -2643 248 -2642
rect 310 -2643 311 -2642
rect 317 -2643 318 -2642
rect 450 -2643 451 -2642
rect 534 -2643 535 -2642
rect 653 -2643 654 -2642
rect 702 -2643 703 -2642
rect 982 -2643 983 -2642
rect 1017 -2643 1018 -2642
rect 1024 -2643 1025 -2642
rect 1062 -2643 1063 -2642
rect 1591 -2643 1592 -2642
rect 86 -2645 87 -2644
rect 702 -2645 703 -2644
rect 737 -2645 738 -2644
rect 1668 -2645 1669 -2644
rect 86 -2647 87 -2646
rect 1577 -2647 1578 -2646
rect 289 -2649 290 -2648
rect 464 -2649 465 -2648
rect 534 -2649 535 -2648
rect 800 -2649 801 -2648
rect 1017 -2649 1018 -2648
rect 1031 -2649 1032 -2648
rect 1094 -2649 1095 -2648
rect 1234 -2649 1235 -2648
rect 1290 -2649 1291 -2648
rect 1402 -2649 1403 -2648
rect 338 -2651 339 -2650
rect 387 -2651 388 -2650
rect 411 -2651 412 -2650
rect 485 -2651 486 -2650
rect 541 -2651 542 -2650
rect 863 -2651 864 -2650
rect 1031 -2651 1032 -2650
rect 1360 -2651 1361 -2650
rect 219 -2653 220 -2652
rect 338 -2653 339 -2652
rect 345 -2653 346 -2652
rect 709 -2653 710 -2652
rect 737 -2653 738 -2652
rect 877 -2653 878 -2652
rect 1097 -2653 1098 -2652
rect 1472 -2653 1473 -2652
rect 82 -2655 83 -2654
rect 219 -2655 220 -2654
rect 450 -2655 451 -2654
rect 1213 -2655 1214 -2654
rect 1290 -2655 1291 -2654
rect 1332 -2655 1333 -2654
rect 1472 -2655 1473 -2654
rect 1535 -2655 1536 -2654
rect 628 -2657 629 -2656
rect 947 -2657 948 -2656
rect 1101 -2657 1102 -2656
rect 1115 -2657 1116 -2656
rect 1311 -2657 1312 -2656
rect 1367 -2657 1368 -2656
rect 1535 -2657 1536 -2656
rect 1605 -2657 1606 -2656
rect 443 -2659 444 -2658
rect 1605 -2659 1606 -2658
rect 331 -2661 332 -2660
rect 443 -2661 444 -2660
rect 709 -2661 710 -2660
rect 723 -2661 724 -2660
rect 754 -2661 755 -2660
rect 1577 -2661 1578 -2660
rect 331 -2663 332 -2662
rect 352 -2663 353 -2662
rect 723 -2663 724 -2662
rect 842 -2663 843 -2662
rect 863 -2663 864 -2662
rect 1045 -2663 1046 -2662
rect 1115 -2663 1116 -2662
rect 1136 -2663 1137 -2662
rect 1332 -2663 1333 -2662
rect 1388 -2663 1389 -2662
rect 114 -2665 115 -2664
rect 352 -2665 353 -2664
rect 366 -2665 367 -2664
rect 1045 -2665 1046 -2664
rect 1073 -2665 1074 -2664
rect 1136 -2665 1137 -2664
rect 1367 -2665 1368 -2664
rect 1409 -2665 1410 -2664
rect 366 -2667 367 -2666
rect 583 -2667 584 -2666
rect 768 -2667 769 -2666
rect 1073 -2667 1074 -2666
rect 1388 -2667 1389 -2666
rect 1465 -2667 1466 -2666
rect 415 -2669 416 -2668
rect 583 -2669 584 -2668
rect 877 -2669 878 -2668
rect 912 -2669 913 -2668
rect 1409 -2669 1410 -2668
rect 1479 -2669 1480 -2668
rect 513 -2671 514 -2670
rect 842 -2671 843 -2670
rect 912 -2671 913 -2670
rect 919 -2671 920 -2670
rect 1465 -2671 1466 -2670
rect 1528 -2671 1529 -2670
rect 740 -2673 741 -2672
rect 1479 -2673 1480 -2672
rect 1528 -2673 1529 -2672
rect 1598 -2673 1599 -2672
rect 919 -2675 920 -2674
rect 968 -2675 969 -2674
rect 1444 -2675 1445 -2674
rect 1598 -2675 1599 -2674
rect 870 -2677 871 -2676
rect 1444 -2677 1445 -2676
rect 688 -2679 689 -2678
rect 870 -2679 871 -2678
rect 968 -2679 969 -2678
rect 996 -2679 997 -2678
rect 618 -2681 619 -2680
rect 688 -2681 689 -2680
rect 677 -2683 678 -2682
rect 996 -2683 997 -2682
rect 37 -2694 38 -2693
rect 569 -2694 570 -2693
rect 579 -2694 580 -2693
rect 793 -2694 794 -2693
rect 803 -2694 804 -2693
rect 1395 -2694 1396 -2693
rect 51 -2696 52 -2695
rect 901 -2696 902 -2695
rect 926 -2696 927 -2695
rect 1097 -2696 1098 -2695
rect 1395 -2696 1396 -2695
rect 1486 -2696 1487 -2695
rect 51 -2698 52 -2697
rect 212 -2698 213 -2697
rect 250 -2698 251 -2697
rect 702 -2698 703 -2697
rect 733 -2698 734 -2697
rect 1066 -2698 1067 -2697
rect 1094 -2698 1095 -2697
rect 1703 -2698 1704 -2697
rect 58 -2700 59 -2699
rect 628 -2700 629 -2699
rect 649 -2700 650 -2699
rect 849 -2700 850 -2699
rect 954 -2700 955 -2699
rect 1241 -2700 1242 -2699
rect 1486 -2700 1487 -2699
rect 1696 -2700 1697 -2699
rect 58 -2702 59 -2701
rect 240 -2702 241 -2701
rect 250 -2702 251 -2701
rect 632 -2702 633 -2701
rect 660 -2702 661 -2701
rect 702 -2702 703 -2701
rect 758 -2702 759 -2701
rect 1048 -2702 1049 -2701
rect 1066 -2702 1067 -2701
rect 1122 -2702 1123 -2701
rect 1241 -2702 1242 -2701
rect 1290 -2702 1291 -2701
rect 65 -2704 66 -2703
rect 653 -2704 654 -2703
rect 660 -2704 661 -2703
rect 670 -2704 671 -2703
rect 674 -2704 675 -2703
rect 1297 -2704 1298 -2703
rect 65 -2706 66 -2705
rect 887 -2706 888 -2705
rect 954 -2706 955 -2705
rect 1101 -2706 1102 -2705
rect 1290 -2706 1291 -2705
rect 1430 -2706 1431 -2705
rect 68 -2708 69 -2707
rect 1045 -2708 1046 -2707
rect 1094 -2708 1095 -2707
rect 1668 -2708 1669 -2707
rect 72 -2710 73 -2709
rect 418 -2710 419 -2709
rect 453 -2710 454 -2709
rect 520 -2710 521 -2709
rect 523 -2710 524 -2709
rect 1185 -2710 1186 -2709
rect 1297 -2710 1298 -2709
rect 1416 -2710 1417 -2709
rect 1430 -2710 1431 -2709
rect 1556 -2710 1557 -2709
rect 82 -2712 83 -2711
rect 786 -2712 787 -2711
rect 793 -2712 794 -2711
rect 947 -2712 948 -2711
rect 957 -2712 958 -2711
rect 1549 -2712 1550 -2711
rect 1556 -2712 1557 -2711
rect 1577 -2712 1578 -2711
rect 110 -2714 111 -2713
rect 1283 -2714 1284 -2713
rect 1416 -2714 1417 -2713
rect 1619 -2714 1620 -2713
rect 114 -2716 115 -2715
rect 555 -2716 556 -2715
rect 583 -2716 584 -2715
rect 1510 -2716 1511 -2715
rect 1549 -2716 1550 -2715
rect 1598 -2716 1599 -2715
rect 114 -2718 115 -2717
rect 639 -2718 640 -2717
rect 653 -2718 654 -2717
rect 1122 -2718 1123 -2717
rect 1283 -2718 1284 -2717
rect 1423 -2718 1424 -2717
rect 117 -2720 118 -2719
rect 618 -2720 619 -2719
rect 625 -2720 626 -2719
rect 884 -2720 885 -2719
rect 947 -2720 948 -2719
rect 1150 -2720 1151 -2719
rect 1423 -2720 1424 -2719
rect 1626 -2720 1627 -2719
rect 121 -2722 122 -2721
rect 800 -2722 801 -2721
rect 814 -2722 815 -2721
rect 845 -2722 846 -2721
rect 849 -2722 850 -2721
rect 1003 -2722 1004 -2721
rect 1034 -2722 1035 -2721
rect 1381 -2722 1382 -2721
rect 121 -2724 122 -2723
rect 247 -2724 248 -2723
rect 275 -2724 276 -2723
rect 278 -2724 279 -2723
rect 289 -2724 290 -2723
rect 478 -2724 479 -2723
rect 481 -2724 482 -2723
rect 562 -2724 563 -2723
rect 583 -2724 584 -2723
rect 982 -2724 983 -2723
rect 989 -2724 990 -2723
rect 1654 -2724 1655 -2723
rect 107 -2726 108 -2725
rect 289 -2726 290 -2725
rect 331 -2726 332 -2725
rect 775 -2726 776 -2725
rect 786 -2726 787 -2725
rect 940 -2726 941 -2725
rect 989 -2726 990 -2725
rect 1227 -2726 1228 -2725
rect 1381 -2726 1382 -2725
rect 1612 -2726 1613 -2725
rect 86 -2728 87 -2727
rect 107 -2728 108 -2727
rect 128 -2728 129 -2727
rect 754 -2728 755 -2727
rect 758 -2728 759 -2727
rect 933 -2728 934 -2727
rect 940 -2728 941 -2727
rect 1129 -2728 1130 -2727
rect 1150 -2728 1151 -2727
rect 1276 -2728 1277 -2727
rect 86 -2730 87 -2729
rect 1675 -2730 1676 -2729
rect 93 -2732 94 -2731
rect 128 -2732 129 -2731
rect 142 -2732 143 -2731
rect 677 -2732 678 -2731
rect 688 -2732 689 -2731
rect 1199 -2732 1200 -2731
rect 1227 -2732 1228 -2731
rect 1409 -2732 1410 -2731
rect 72 -2734 73 -2733
rect 93 -2734 94 -2733
rect 149 -2734 150 -2733
rect 152 -2734 153 -2733
rect 166 -2734 167 -2733
rect 331 -2734 332 -2733
rect 352 -2734 353 -2733
rect 639 -2734 640 -2733
rect 667 -2734 668 -2733
rect 681 -2734 682 -2733
rect 765 -2734 766 -2733
rect 1192 -2734 1193 -2733
rect 1199 -2734 1200 -2733
rect 1325 -2734 1326 -2733
rect 89 -2736 90 -2735
rect 142 -2736 143 -2735
rect 149 -2736 150 -2735
rect 198 -2736 199 -2735
rect 201 -2736 202 -2735
rect 730 -2736 731 -2735
rect 814 -2736 815 -2735
rect 863 -2736 864 -2735
rect 873 -2736 874 -2735
rect 1129 -2736 1130 -2735
rect 1192 -2736 1193 -2735
rect 1339 -2736 1340 -2735
rect 89 -2738 90 -2737
rect 338 -2738 339 -2737
rect 373 -2738 374 -2737
rect 415 -2738 416 -2737
rect 429 -2738 430 -2737
rect 800 -2738 801 -2737
rect 835 -2738 836 -2737
rect 898 -2738 899 -2737
rect 933 -2738 934 -2737
rect 1073 -2738 1074 -2737
rect 1101 -2738 1102 -2737
rect 1311 -2738 1312 -2737
rect 1325 -2738 1326 -2737
rect 1500 -2738 1501 -2737
rect 166 -2740 167 -2739
rect 576 -2740 577 -2739
rect 593 -2740 594 -2739
rect 1185 -2740 1186 -2739
rect 1311 -2740 1312 -2739
rect 1605 -2740 1606 -2739
rect 180 -2742 181 -2741
rect 1633 -2742 1634 -2741
rect 184 -2744 185 -2743
rect 198 -2744 199 -2743
rect 205 -2744 206 -2743
rect 338 -2744 339 -2743
rect 359 -2744 360 -2743
rect 373 -2744 374 -2743
rect 401 -2744 402 -2743
rect 569 -2744 570 -2743
rect 597 -2744 598 -2743
rect 1689 -2744 1690 -2743
rect 156 -2746 157 -2745
rect 205 -2746 206 -2745
rect 212 -2746 213 -2745
rect 226 -2746 227 -2745
rect 240 -2746 241 -2745
rect 261 -2746 262 -2745
rect 268 -2746 269 -2745
rect 352 -2746 353 -2745
rect 359 -2746 360 -2745
rect 485 -2746 486 -2745
rect 506 -2746 507 -2745
rect 632 -2746 633 -2745
rect 667 -2746 668 -2745
rect 1017 -2746 1018 -2745
rect 1045 -2746 1046 -2745
rect 1584 -2746 1585 -2745
rect 44 -2748 45 -2747
rect 226 -2748 227 -2747
rect 254 -2748 255 -2747
rect 261 -2748 262 -2747
rect 268 -2748 269 -2747
rect 467 -2748 468 -2747
rect 485 -2748 486 -2747
rect 723 -2748 724 -2747
rect 730 -2748 731 -2747
rect 856 -2748 857 -2747
rect 863 -2748 864 -2747
rect 1188 -2748 1189 -2747
rect 1339 -2748 1340 -2747
rect 1542 -2748 1543 -2747
rect 44 -2750 45 -2749
rect 100 -2750 101 -2749
rect 131 -2750 132 -2749
rect 723 -2750 724 -2749
rect 835 -2750 836 -2749
rect 996 -2750 997 -2749
rect 1003 -2750 1004 -2749
rect 1136 -2750 1137 -2749
rect 1374 -2750 1375 -2749
rect 1542 -2750 1543 -2749
rect 96 -2752 97 -2751
rect 156 -2752 157 -2751
rect 184 -2752 185 -2751
rect 191 -2752 192 -2751
rect 254 -2752 255 -2751
rect 383 -2752 384 -2751
rect 401 -2752 402 -2751
rect 436 -2752 437 -2751
rect 450 -2752 451 -2751
rect 982 -2752 983 -2751
rect 1017 -2752 1018 -2751
rect 1171 -2752 1172 -2751
rect 1374 -2752 1375 -2751
rect 1437 -2752 1438 -2751
rect 1458 -2752 1459 -2751
rect 1500 -2752 1501 -2751
rect 100 -2754 101 -2753
rect 282 -2754 283 -2753
rect 345 -2754 346 -2753
rect 996 -2754 997 -2753
rect 1073 -2754 1074 -2753
rect 1255 -2754 1256 -2753
rect 1437 -2754 1438 -2753
rect 1563 -2754 1564 -2753
rect 275 -2756 276 -2755
rect 324 -2756 325 -2755
rect 345 -2756 346 -2755
rect 492 -2756 493 -2755
rect 520 -2756 521 -2755
rect 688 -2756 689 -2755
rect 716 -2756 717 -2755
rect 856 -2756 857 -2755
rect 884 -2756 885 -2755
rect 1255 -2756 1256 -2755
rect 1458 -2756 1459 -2755
rect 1661 -2756 1662 -2755
rect 233 -2758 234 -2757
rect 492 -2758 493 -2757
rect 534 -2758 535 -2757
rect 1031 -2758 1032 -2757
rect 1136 -2758 1137 -2757
rect 1269 -2758 1270 -2757
rect 177 -2760 178 -2759
rect 233 -2760 234 -2759
rect 282 -2760 283 -2759
rect 450 -2760 451 -2759
rect 457 -2760 458 -2759
rect 1409 -2760 1410 -2759
rect 229 -2762 230 -2761
rect 457 -2762 458 -2761
rect 534 -2762 535 -2761
rect 975 -2762 976 -2761
rect 1031 -2762 1032 -2761
rect 1087 -2762 1088 -2761
rect 1171 -2762 1172 -2761
rect 1360 -2762 1361 -2761
rect 317 -2764 318 -2763
rect 324 -2764 325 -2763
rect 366 -2764 367 -2763
rect 506 -2764 507 -2763
rect 541 -2764 542 -2763
rect 894 -2764 895 -2763
rect 898 -2764 899 -2763
rect 926 -2764 927 -2763
rect 975 -2764 976 -2763
rect 1052 -2764 1053 -2763
rect 1269 -2764 1270 -2763
rect 1451 -2764 1452 -2763
rect 296 -2766 297 -2765
rect 366 -2766 367 -2765
rect 408 -2766 409 -2765
rect 1279 -2766 1280 -2765
rect 1360 -2766 1361 -2765
rect 1591 -2766 1592 -2765
rect 296 -2768 297 -2767
rect 422 -2768 423 -2767
rect 429 -2768 430 -2767
rect 611 -2768 612 -2767
rect 618 -2768 619 -2767
rect 1108 -2768 1109 -2767
rect 1451 -2768 1452 -2767
rect 1640 -2768 1641 -2767
rect 317 -2770 318 -2769
rect 443 -2770 444 -2769
rect 499 -2770 500 -2769
rect 611 -2770 612 -2769
rect 625 -2770 626 -2769
rect 709 -2770 710 -2769
rect 716 -2770 717 -2769
rect 751 -2770 752 -2769
rect 870 -2770 871 -2769
rect 1087 -2770 1088 -2769
rect 1108 -2770 1109 -2769
rect 1262 -2770 1263 -2769
rect 278 -2772 279 -2771
rect 443 -2772 444 -2771
rect 499 -2772 500 -2771
rect 744 -2772 745 -2771
rect 751 -2772 752 -2771
rect 772 -2772 773 -2771
rect 870 -2772 871 -2771
rect 1164 -2772 1165 -2771
rect 1262 -2772 1263 -2771
rect 1472 -2772 1473 -2771
rect 411 -2774 412 -2773
rect 527 -2774 528 -2773
rect 541 -2774 542 -2773
rect 590 -2774 591 -2773
rect 597 -2774 598 -2773
rect 919 -2774 920 -2773
rect 1052 -2774 1053 -2773
rect 1332 -2774 1333 -2773
rect 1472 -2774 1473 -2773
rect 1507 -2774 1508 -2773
rect 415 -2776 416 -2775
rect 684 -2776 685 -2775
rect 709 -2776 710 -2775
rect 877 -2776 878 -2775
rect 894 -2776 895 -2775
rect 1682 -2776 1683 -2775
rect 247 -2778 248 -2777
rect 877 -2778 878 -2777
rect 919 -2778 920 -2777
rect 1213 -2778 1214 -2777
rect 1332 -2778 1333 -2777
rect 1535 -2778 1536 -2777
rect 422 -2780 423 -2779
rect 803 -2780 804 -2779
rect 1164 -2780 1165 -2779
rect 1367 -2780 1368 -2779
rect 1493 -2780 1494 -2779
rect 1507 -2780 1508 -2779
rect 436 -2782 437 -2781
rect 548 -2782 549 -2781
rect 555 -2782 556 -2781
rect 807 -2782 808 -2781
rect 1213 -2782 1214 -2781
rect 1444 -2782 1445 -2781
rect 1493 -2782 1494 -2781
rect 1647 -2782 1648 -2781
rect 219 -2784 220 -2783
rect 548 -2784 549 -2783
rect 562 -2784 563 -2783
rect 779 -2784 780 -2783
rect 807 -2784 808 -2783
rect 961 -2784 962 -2783
rect 1248 -2784 1249 -2783
rect 1444 -2784 1445 -2783
rect 170 -2786 171 -2785
rect 219 -2786 220 -2785
rect 527 -2786 528 -2785
rect 985 -2786 986 -2785
rect 1206 -2786 1207 -2785
rect 1248 -2786 1249 -2785
rect 1346 -2786 1347 -2785
rect 1535 -2786 1536 -2785
rect 170 -2788 171 -2787
rect 768 -2788 769 -2787
rect 842 -2788 843 -2787
rect 1206 -2788 1207 -2787
rect 1346 -2788 1347 -2787
rect 1514 -2788 1515 -2787
rect 79 -2790 80 -2789
rect 1514 -2790 1515 -2789
rect 79 -2792 80 -2791
rect 394 -2792 395 -2791
rect 590 -2792 591 -2791
rect 821 -2792 822 -2791
rect 842 -2792 843 -2791
rect 912 -2792 913 -2791
rect 961 -2792 962 -2791
rect 1115 -2792 1116 -2791
rect 1367 -2792 1368 -2791
rect 1388 -2792 1389 -2791
rect 394 -2794 395 -2793
rect 471 -2794 472 -2793
rect 600 -2794 601 -2793
rect 737 -2794 738 -2793
rect 744 -2794 745 -2793
rect 828 -2794 829 -2793
rect 912 -2794 913 -2793
rect 968 -2794 969 -2793
rect 1115 -2794 1116 -2793
rect 1388 -2794 1389 -2793
rect 135 -2796 136 -2795
rect 471 -2796 472 -2795
rect 674 -2796 675 -2795
rect 1080 -2796 1081 -2795
rect 135 -2798 136 -2797
rect 646 -2798 647 -2797
rect 681 -2798 682 -2797
rect 1318 -2798 1319 -2797
rect 464 -2800 465 -2799
rect 737 -2800 738 -2799
rect 761 -2800 762 -2799
rect 779 -2800 780 -2799
rect 821 -2800 822 -2799
rect 1010 -2800 1011 -2799
rect 1318 -2800 1319 -2799
rect 1479 -2800 1480 -2799
rect 163 -2802 164 -2801
rect 1479 -2802 1480 -2801
rect 163 -2804 164 -2803
rect 905 -2804 906 -2803
rect 999 -2804 1000 -2803
rect 1080 -2804 1081 -2803
rect 310 -2806 311 -2805
rect 464 -2806 465 -2805
rect 765 -2806 766 -2805
rect 968 -2806 969 -2805
rect 303 -2808 304 -2807
rect 310 -2808 311 -2807
rect 768 -2808 769 -2807
rect 1024 -2808 1025 -2807
rect 303 -2810 304 -2809
rect 513 -2810 514 -2809
rect 772 -2810 773 -2809
rect 828 -2810 829 -2809
rect 838 -2810 839 -2809
rect 905 -2810 906 -2809
rect 1024 -2810 1025 -2809
rect 1157 -2810 1158 -2809
rect 513 -2812 514 -2811
rect 604 -2812 605 -2811
rect 891 -2812 892 -2811
rect 1010 -2812 1011 -2811
rect 1157 -2812 1158 -2811
rect 1178 -2812 1179 -2811
rect 604 -2814 605 -2813
rect 695 -2814 696 -2813
rect 1178 -2814 1179 -2813
rect 1220 -2814 1221 -2813
rect 695 -2816 696 -2815
rect 1038 -2816 1039 -2815
rect 1220 -2816 1221 -2815
rect 1465 -2816 1466 -2815
rect 1038 -2818 1039 -2817
rect 1059 -2818 1060 -2817
rect 1465 -2818 1466 -2817
rect 1521 -2818 1522 -2817
rect 1059 -2820 1060 -2819
rect 1353 -2820 1354 -2819
rect 1304 -2822 1305 -2821
rect 1521 -2822 1522 -2821
rect 1234 -2824 1235 -2823
rect 1304 -2824 1305 -2823
rect 1353 -2824 1354 -2823
rect 1570 -2824 1571 -2823
rect 1234 -2826 1235 -2825
rect 1402 -2826 1403 -2825
rect 1402 -2828 1403 -2827
rect 1528 -2828 1529 -2827
rect 1143 -2830 1144 -2829
rect 1528 -2830 1529 -2829
rect 1143 -2832 1144 -2831
rect 1276 -2832 1277 -2831
rect 30 -2843 31 -2842
rect 457 -2843 458 -2842
rect 506 -2843 507 -2842
rect 656 -2843 657 -2842
rect 765 -2843 766 -2842
rect 842 -2843 843 -2842
rect 887 -2843 888 -2842
rect 929 -2843 930 -2842
rect 982 -2843 983 -2842
rect 1402 -2843 1403 -2842
rect 1514 -2843 1515 -2842
rect 1556 -2843 1557 -2842
rect 37 -2845 38 -2844
rect 502 -2845 503 -2844
rect 583 -2845 584 -2844
rect 653 -2845 654 -2844
rect 702 -2845 703 -2844
rect 842 -2845 843 -2844
rect 898 -2845 899 -2844
rect 1374 -2845 1375 -2844
rect 1395 -2845 1396 -2844
rect 1402 -2845 1403 -2844
rect 37 -2847 38 -2846
rect 499 -2847 500 -2846
rect 569 -2847 570 -2846
rect 583 -2847 584 -2846
rect 593 -2847 594 -2846
rect 793 -2847 794 -2846
rect 803 -2847 804 -2846
rect 961 -2847 962 -2846
rect 996 -2847 997 -2846
rect 1192 -2847 1193 -2846
rect 1202 -2847 1203 -2846
rect 1367 -2847 1368 -2846
rect 44 -2849 45 -2848
rect 117 -2849 118 -2848
rect 121 -2849 122 -2848
rect 565 -2849 566 -2848
rect 607 -2849 608 -2848
rect 681 -2849 682 -2848
rect 751 -2849 752 -2848
rect 765 -2849 766 -2848
rect 775 -2849 776 -2848
rect 1199 -2849 1200 -2848
rect 1276 -2849 1277 -2848
rect 1332 -2849 1333 -2848
rect 1367 -2849 1368 -2848
rect 1388 -2849 1389 -2848
rect 51 -2851 52 -2850
rect 226 -2851 227 -2850
rect 250 -2851 251 -2850
rect 1374 -2851 1375 -2850
rect 1388 -2851 1389 -2850
rect 1444 -2851 1445 -2850
rect 51 -2853 52 -2852
rect 625 -2853 626 -2852
rect 653 -2853 654 -2852
rect 828 -2853 829 -2852
rect 877 -2853 878 -2852
rect 1395 -2853 1396 -2852
rect 72 -2855 73 -2854
rect 1115 -2855 1116 -2854
rect 1118 -2855 1119 -2854
rect 1500 -2855 1501 -2854
rect 75 -2857 76 -2856
rect 527 -2857 528 -2856
rect 618 -2857 619 -2856
rect 884 -2857 885 -2856
rect 898 -2857 899 -2856
rect 1507 -2857 1508 -2856
rect 86 -2859 87 -2858
rect 303 -2859 304 -2858
rect 345 -2859 346 -2858
rect 684 -2859 685 -2858
rect 751 -2859 752 -2858
rect 786 -2859 787 -2858
rect 807 -2859 808 -2858
rect 915 -2859 916 -2858
rect 947 -2859 948 -2858
rect 982 -2859 983 -2858
rect 996 -2859 997 -2858
rect 1066 -2859 1067 -2858
rect 1097 -2859 1098 -2858
rect 1437 -2859 1438 -2858
rect 1500 -2859 1501 -2858
rect 1549 -2859 1550 -2858
rect 93 -2861 94 -2860
rect 107 -2861 108 -2860
rect 121 -2861 122 -2860
rect 264 -2861 265 -2860
rect 268 -2861 269 -2860
rect 758 -2861 759 -2860
rect 828 -2861 829 -2860
rect 1031 -2861 1032 -2860
rect 1038 -2861 1039 -2860
rect 1094 -2861 1095 -2860
rect 1164 -2861 1165 -2860
rect 1185 -2861 1186 -2860
rect 1188 -2861 1189 -2860
rect 1430 -2861 1431 -2860
rect 93 -2863 94 -2862
rect 604 -2863 605 -2862
rect 618 -2863 619 -2862
rect 716 -2863 717 -2862
rect 779 -2863 780 -2862
rect 1038 -2863 1039 -2862
rect 1048 -2863 1049 -2862
rect 1136 -2863 1137 -2862
rect 1185 -2863 1186 -2862
rect 1206 -2863 1207 -2862
rect 1279 -2863 1280 -2862
rect 1451 -2863 1452 -2862
rect 96 -2865 97 -2864
rect 534 -2865 535 -2864
rect 625 -2865 626 -2864
rect 688 -2865 689 -2864
rect 695 -2865 696 -2864
rect 807 -2865 808 -2864
rect 856 -2865 857 -2864
rect 877 -2865 878 -2864
rect 905 -2865 906 -2864
rect 1066 -2865 1067 -2864
rect 1192 -2865 1193 -2864
rect 1213 -2865 1214 -2864
rect 1248 -2865 1249 -2864
rect 1451 -2865 1452 -2864
rect 100 -2867 101 -2866
rect 177 -2867 178 -2866
rect 226 -2867 227 -2866
rect 261 -2867 262 -2866
rect 268 -2867 269 -2866
rect 394 -2867 395 -2866
rect 411 -2867 412 -2866
rect 1206 -2867 1207 -2866
rect 1213 -2867 1214 -2866
rect 1283 -2867 1284 -2866
rect 1318 -2867 1319 -2866
rect 1332 -2867 1333 -2866
rect 1430 -2867 1431 -2866
rect 1458 -2867 1459 -2866
rect 100 -2869 101 -2868
rect 229 -2869 230 -2868
rect 275 -2869 276 -2868
rect 303 -2869 304 -2868
rect 345 -2869 346 -2868
rect 387 -2869 388 -2868
rect 429 -2869 430 -2868
rect 569 -2869 570 -2868
rect 576 -2869 577 -2868
rect 695 -2869 696 -2868
rect 709 -2869 710 -2868
rect 786 -2869 787 -2868
rect 800 -2869 801 -2868
rect 1164 -2869 1165 -2868
rect 1283 -2869 1284 -2868
rect 1510 -2869 1511 -2868
rect 107 -2871 108 -2870
rect 541 -2871 542 -2870
rect 646 -2871 647 -2870
rect 1437 -2871 1438 -2870
rect 1458 -2871 1459 -2870
rect 1535 -2871 1536 -2870
rect 128 -2873 129 -2872
rect 793 -2873 794 -2872
rect 800 -2873 801 -2872
rect 849 -2873 850 -2872
rect 866 -2873 867 -2872
rect 884 -2873 885 -2872
rect 905 -2873 906 -2872
rect 933 -2873 934 -2872
rect 940 -2873 941 -2872
rect 1031 -2873 1032 -2872
rect 1129 -2873 1130 -2872
rect 1248 -2873 1249 -2872
rect 1311 -2873 1312 -2872
rect 1318 -2873 1319 -2872
rect 128 -2875 129 -2874
rect 240 -2875 241 -2874
rect 275 -2875 276 -2874
rect 310 -2875 311 -2874
rect 359 -2875 360 -2874
rect 387 -2875 388 -2874
rect 450 -2875 451 -2874
rect 1409 -2875 1410 -2874
rect 135 -2877 136 -2876
rect 534 -2877 535 -2876
rect 541 -2877 542 -2876
rect 639 -2877 640 -2876
rect 646 -2877 647 -2876
rect 989 -2877 990 -2876
rect 1003 -2877 1004 -2876
rect 1136 -2877 1137 -2876
rect 1311 -2877 1312 -2876
rect 1360 -2877 1361 -2876
rect 1409 -2877 1410 -2876
rect 1423 -2877 1424 -2876
rect 135 -2879 136 -2878
rect 180 -2879 181 -2878
rect 191 -2879 192 -2878
rect 310 -2879 311 -2878
rect 331 -2879 332 -2878
rect 450 -2879 451 -2878
rect 457 -2879 458 -2878
rect 590 -2879 591 -2878
rect 660 -2879 661 -2878
rect 709 -2879 710 -2878
rect 716 -2879 717 -2878
rect 768 -2879 769 -2878
rect 779 -2879 780 -2878
rect 863 -2879 864 -2878
rect 912 -2879 913 -2878
rect 1045 -2879 1046 -2878
rect 1080 -2879 1081 -2878
rect 1129 -2879 1130 -2878
rect 1360 -2879 1361 -2878
rect 1381 -2879 1382 -2878
rect 1423 -2879 1424 -2878
rect 1486 -2879 1487 -2878
rect 142 -2881 143 -2880
rect 772 -2881 773 -2880
rect 863 -2881 864 -2880
rect 1150 -2881 1151 -2880
rect 1381 -2881 1382 -2880
rect 1416 -2881 1417 -2880
rect 1486 -2881 1487 -2880
rect 1521 -2881 1522 -2880
rect 142 -2883 143 -2882
rect 212 -2883 213 -2882
rect 219 -2883 220 -2882
rect 394 -2883 395 -2882
rect 474 -2883 475 -2882
rect 1115 -2883 1116 -2882
rect 1150 -2883 1151 -2882
rect 1227 -2883 1228 -2882
rect 1416 -2883 1417 -2882
rect 1447 -2883 1448 -2882
rect 72 -2885 73 -2884
rect 212 -2885 213 -2884
rect 219 -2885 220 -2884
rect 999 -2885 1000 -2884
rect 1003 -2885 1004 -2884
rect 1073 -2885 1074 -2884
rect 1080 -2885 1081 -2884
rect 1241 -2885 1242 -2884
rect 170 -2887 171 -2886
rect 499 -2887 500 -2886
rect 523 -2887 524 -2886
rect 940 -2887 941 -2886
rect 961 -2887 962 -2886
rect 975 -2887 976 -2886
rect 1010 -2887 1011 -2886
rect 1045 -2887 1046 -2886
rect 1122 -2887 1123 -2886
rect 1227 -2887 1228 -2886
rect 1241 -2887 1242 -2886
rect 1262 -2887 1263 -2886
rect 170 -2889 171 -2888
rect 1199 -2889 1200 -2888
rect 177 -2891 178 -2890
rect 240 -2891 241 -2890
rect 282 -2891 283 -2890
rect 576 -2891 577 -2890
rect 660 -2891 661 -2890
rect 744 -2891 745 -2890
rect 870 -2891 871 -2890
rect 1073 -2891 1074 -2890
rect 1087 -2891 1088 -2890
rect 1262 -2891 1263 -2890
rect 163 -2893 164 -2892
rect 282 -2893 283 -2892
rect 331 -2893 332 -2892
rect 366 -2893 367 -2892
rect 373 -2893 374 -2892
rect 520 -2893 521 -2892
rect 527 -2893 528 -2892
rect 548 -2893 549 -2892
rect 555 -2893 556 -2892
rect 639 -2893 640 -2892
rect 667 -2893 668 -2892
rect 849 -2893 850 -2892
rect 912 -2893 913 -2892
rect 1493 -2893 1494 -2892
rect 114 -2895 115 -2894
rect 520 -2895 521 -2894
rect 548 -2895 549 -2894
rect 611 -2895 612 -2894
rect 667 -2895 668 -2894
rect 744 -2895 745 -2894
rect 926 -2895 927 -2894
rect 989 -2895 990 -2894
rect 1010 -2895 1011 -2894
rect 1178 -2895 1179 -2894
rect 1493 -2895 1494 -2894
rect 1528 -2895 1529 -2894
rect 163 -2897 164 -2896
rect 247 -2897 248 -2896
rect 250 -2897 251 -2896
rect 870 -2897 871 -2896
rect 926 -2897 927 -2896
rect 1304 -2897 1305 -2896
rect 191 -2899 192 -2898
rect 205 -2899 206 -2898
rect 359 -2899 360 -2898
rect 936 -2899 937 -2898
rect 975 -2899 976 -2898
rect 1157 -2899 1158 -2898
rect 1178 -2899 1179 -2898
rect 1290 -2899 1291 -2898
rect 1304 -2899 1305 -2898
rect 1353 -2899 1354 -2898
rect 205 -2901 206 -2900
rect 254 -2901 255 -2900
rect 366 -2901 367 -2900
rect 649 -2901 650 -2900
rect 674 -2901 675 -2900
rect 702 -2901 703 -2900
rect 737 -2901 738 -2900
rect 856 -2901 857 -2900
rect 968 -2901 969 -2900
rect 1353 -2901 1354 -2900
rect 254 -2903 255 -2902
rect 338 -2903 339 -2902
rect 380 -2903 381 -2902
rect 429 -2903 430 -2902
rect 485 -2903 486 -2902
rect 590 -2903 591 -2902
rect 597 -2903 598 -2902
rect 674 -2903 675 -2902
rect 761 -2903 762 -2902
rect 968 -2903 969 -2902
rect 1027 -2903 1028 -2902
rect 1479 -2903 1480 -2902
rect 289 -2905 290 -2904
rect 338 -2905 339 -2904
rect 380 -2905 381 -2904
rect 478 -2905 479 -2904
rect 485 -2905 486 -2904
rect 562 -2905 563 -2904
rect 611 -2905 612 -2904
rect 814 -2905 815 -2904
rect 1052 -2905 1053 -2904
rect 1122 -2905 1123 -2904
rect 1157 -2905 1158 -2904
rect 1339 -2905 1340 -2904
rect 1479 -2905 1480 -2904
rect 1542 -2905 1543 -2904
rect 44 -2907 45 -2906
rect 562 -2907 563 -2906
rect 761 -2907 762 -2906
rect 947 -2907 948 -2906
rect 1052 -2907 1053 -2906
rect 1101 -2907 1102 -2906
rect 1255 -2907 1256 -2906
rect 1339 -2907 1340 -2906
rect 65 -2909 66 -2908
rect 289 -2909 290 -2908
rect 408 -2909 409 -2908
rect 737 -2909 738 -2908
rect 814 -2909 815 -2908
rect 835 -2909 836 -2908
rect 1059 -2909 1060 -2908
rect 1087 -2909 1088 -2908
rect 1101 -2909 1102 -2908
rect 1143 -2909 1144 -2908
rect 1255 -2909 1256 -2908
rect 1297 -2909 1298 -2908
rect 65 -2911 66 -2910
rect 415 -2911 416 -2910
rect 436 -2911 437 -2910
rect 597 -2911 598 -2910
rect 733 -2911 734 -2910
rect 1297 -2911 1298 -2910
rect 110 -2913 111 -2912
rect 835 -2913 836 -2912
rect 1059 -2913 1060 -2912
rect 1108 -2913 1109 -2912
rect 1143 -2913 1144 -2912
rect 1171 -2913 1172 -2912
rect 1290 -2913 1291 -2912
rect 1346 -2913 1347 -2912
rect 401 -2915 402 -2914
rect 415 -2915 416 -2914
rect 436 -2915 437 -2914
rect 492 -2915 493 -2914
rect 555 -2915 556 -2914
rect 919 -2915 920 -2914
rect 1171 -2915 1172 -2914
rect 1234 -2915 1235 -2914
rect 58 -2917 59 -2916
rect 401 -2917 402 -2916
rect 408 -2917 409 -2916
rect 464 -2917 465 -2916
rect 478 -2917 479 -2916
rect 901 -2917 902 -2916
rect 919 -2917 920 -2916
rect 954 -2917 955 -2916
rect 1220 -2917 1221 -2916
rect 1234 -2917 1235 -2916
rect 58 -2919 59 -2918
rect 632 -2919 633 -2918
rect 723 -2919 724 -2918
rect 1108 -2919 1109 -2918
rect 1220 -2919 1221 -2918
rect 1269 -2919 1270 -2918
rect 114 -2921 115 -2920
rect 632 -2921 633 -2920
rect 723 -2921 724 -2920
rect 730 -2921 731 -2920
rect 891 -2921 892 -2920
rect 1346 -2921 1347 -2920
rect 149 -2923 150 -2922
rect 891 -2923 892 -2922
rect 954 -2923 955 -2922
rect 1017 -2923 1018 -2922
rect 1269 -2923 1270 -2922
rect 1325 -2923 1326 -2922
rect 149 -2925 150 -2924
rect 184 -2925 185 -2924
rect 317 -2925 318 -2924
rect 464 -2925 465 -2924
rect 471 -2925 472 -2924
rect 730 -2925 731 -2924
rect 1017 -2925 1018 -2924
rect 1024 -2925 1025 -2924
rect 184 -2927 185 -2926
rect 198 -2927 199 -2926
rect 257 -2927 258 -2926
rect 317 -2927 318 -2926
rect 404 -2927 405 -2926
rect 1325 -2927 1326 -2926
rect 198 -2929 199 -2928
rect 296 -2929 297 -2928
rect 422 -2929 423 -2928
rect 492 -2929 493 -2928
rect 1024 -2929 1025 -2928
rect 1465 -2929 1466 -2928
rect 79 -2931 80 -2930
rect 296 -2931 297 -2930
rect 422 -2931 423 -2930
rect 670 -2931 671 -2930
rect 1465 -2931 1466 -2930
rect 1472 -2931 1473 -2930
rect 79 -2933 80 -2932
rect 324 -2933 325 -2932
rect 471 -2933 472 -2932
rect 506 -2933 507 -2932
rect 233 -2935 234 -2934
rect 324 -2935 325 -2934
rect 233 -2937 234 -2936
rect 352 -2937 353 -2936
rect 352 -2939 353 -2938
rect 513 -2939 514 -2938
rect 443 -2941 444 -2940
rect 513 -2941 514 -2940
rect 156 -2943 157 -2942
rect 443 -2943 444 -2942
rect 30 -2954 31 -2953
rect 72 -2954 73 -2953
rect 79 -2954 80 -2953
rect 474 -2954 475 -2953
rect 523 -2954 524 -2953
rect 632 -2954 633 -2953
rect 635 -2954 636 -2953
rect 968 -2954 969 -2953
rect 982 -2954 983 -2953
rect 1024 -2954 1025 -2953
rect 1038 -2954 1039 -2953
rect 1041 -2954 1042 -2953
rect 1062 -2954 1063 -2953
rect 1430 -2954 1431 -2953
rect 1444 -2954 1445 -2953
rect 1486 -2954 1487 -2953
rect 37 -2956 38 -2955
rect 96 -2956 97 -2955
rect 100 -2956 101 -2955
rect 702 -2956 703 -2955
rect 758 -2956 759 -2955
rect 765 -2956 766 -2955
rect 828 -2956 829 -2955
rect 863 -2956 864 -2955
rect 870 -2956 871 -2955
rect 999 -2956 1000 -2955
rect 1020 -2956 1021 -2955
rect 1150 -2956 1151 -2955
rect 1199 -2956 1200 -2955
rect 1276 -2956 1277 -2955
rect 1447 -2956 1448 -2955
rect 1500 -2956 1501 -2955
rect 37 -2958 38 -2957
rect 121 -2958 122 -2957
rect 124 -2958 125 -2957
rect 310 -2958 311 -2957
rect 366 -2958 367 -2957
rect 852 -2958 853 -2957
rect 870 -2958 871 -2957
rect 1437 -2958 1438 -2957
rect 1472 -2958 1473 -2957
rect 1493 -2958 1494 -2957
rect 44 -2960 45 -2959
rect 250 -2960 251 -2959
rect 254 -2960 255 -2959
rect 324 -2960 325 -2959
rect 373 -2960 374 -2959
rect 450 -2960 451 -2959
rect 464 -2960 465 -2959
rect 670 -2960 671 -2959
rect 684 -2960 685 -2959
rect 1283 -2960 1284 -2959
rect 44 -2962 45 -2961
rect 149 -2962 150 -2961
rect 156 -2962 157 -2961
rect 380 -2962 381 -2961
rect 429 -2962 430 -2961
rect 478 -2962 479 -2961
rect 534 -2962 535 -2961
rect 642 -2962 643 -2961
rect 646 -2962 647 -2961
rect 933 -2962 934 -2961
rect 936 -2962 937 -2961
rect 982 -2962 983 -2961
rect 996 -2962 997 -2961
rect 1185 -2962 1186 -2961
rect 1255 -2962 1256 -2961
rect 1283 -2962 1284 -2961
rect 51 -2964 52 -2963
rect 607 -2964 608 -2963
rect 611 -2964 612 -2963
rect 730 -2964 731 -2963
rect 758 -2964 759 -2963
rect 835 -2964 836 -2963
rect 877 -2964 878 -2963
rect 1024 -2964 1025 -2963
rect 1038 -2964 1039 -2963
rect 1122 -2964 1123 -2963
rect 1143 -2964 1144 -2963
rect 1185 -2964 1186 -2963
rect 1255 -2964 1256 -2963
rect 1395 -2964 1396 -2963
rect 51 -2966 52 -2965
rect 408 -2966 409 -2965
rect 429 -2966 430 -2965
rect 796 -2966 797 -2965
rect 828 -2966 829 -2965
rect 1374 -2966 1375 -2965
rect 65 -2968 66 -2967
rect 79 -2968 80 -2967
rect 93 -2968 94 -2967
rect 621 -2968 622 -2967
rect 625 -2968 626 -2967
rect 765 -2968 766 -2967
rect 793 -2968 794 -2967
rect 877 -2968 878 -2967
rect 922 -2968 923 -2967
rect 1052 -2968 1053 -2967
rect 1073 -2968 1074 -2967
rect 1122 -2968 1123 -2967
rect 1143 -2968 1144 -2967
rect 1241 -2968 1242 -2967
rect 1276 -2968 1277 -2967
rect 1318 -2968 1319 -2967
rect 1374 -2968 1375 -2967
rect 1458 -2968 1459 -2967
rect 65 -2970 66 -2969
rect 250 -2970 251 -2969
rect 254 -2970 255 -2969
rect 275 -2970 276 -2969
rect 289 -2970 290 -2969
rect 366 -2970 367 -2969
rect 373 -2970 374 -2969
rect 597 -2970 598 -2969
rect 632 -2970 633 -2969
rect 723 -2970 724 -2969
rect 933 -2970 934 -2969
rect 989 -2970 990 -2969
rect 996 -2970 997 -2969
rect 1332 -2970 1333 -2969
rect 1458 -2970 1459 -2969
rect 1465 -2970 1466 -2969
rect 100 -2972 101 -2971
rect 541 -2972 542 -2971
rect 555 -2972 556 -2971
rect 863 -2972 864 -2971
rect 954 -2972 955 -2971
rect 968 -2972 969 -2971
rect 1041 -2972 1042 -2971
rect 1073 -2972 1074 -2971
rect 1090 -2972 1091 -2971
rect 1409 -2972 1410 -2971
rect 1465 -2972 1466 -2971
rect 1479 -2972 1480 -2971
rect 114 -2974 115 -2973
rect 149 -2974 150 -2973
rect 159 -2974 160 -2973
rect 520 -2974 521 -2973
rect 527 -2974 528 -2973
rect 541 -2974 542 -2973
rect 555 -2974 556 -2973
rect 873 -2974 874 -2973
rect 954 -2974 955 -2973
rect 1003 -2974 1004 -2973
rect 1052 -2974 1053 -2973
rect 1129 -2974 1130 -2973
rect 1136 -2974 1137 -2973
rect 1318 -2974 1319 -2973
rect 1332 -2974 1333 -2973
rect 1451 -2974 1452 -2973
rect 114 -2976 115 -2975
rect 135 -2976 136 -2975
rect 177 -2976 178 -2975
rect 289 -2976 290 -2975
rect 352 -2976 353 -2975
rect 607 -2976 608 -2975
rect 646 -2976 647 -2975
rect 695 -2976 696 -2975
rect 723 -2976 724 -2975
rect 912 -2976 913 -2975
rect 1003 -2976 1004 -2975
rect 1059 -2976 1060 -2975
rect 1129 -2976 1130 -2975
rect 1171 -2976 1172 -2975
rect 121 -2978 122 -2977
rect 135 -2978 136 -2977
rect 177 -2978 178 -2977
rect 1325 -2978 1326 -2977
rect 180 -2980 181 -2979
rect 394 -2980 395 -2979
rect 408 -2980 409 -2979
rect 464 -2980 465 -2979
rect 534 -2980 535 -2979
rect 744 -2980 745 -2979
rect 912 -2980 913 -2979
rect 975 -2980 976 -2979
rect 1080 -2980 1081 -2979
rect 1171 -2980 1172 -2979
rect 198 -2982 199 -2981
rect 604 -2982 605 -2981
rect 653 -2982 654 -2981
rect 989 -2982 990 -2981
rect 1080 -2982 1081 -2981
rect 1108 -2982 1109 -2981
rect 1136 -2982 1137 -2981
rect 1227 -2982 1228 -2981
rect 201 -2984 202 -2983
rect 513 -2984 514 -2983
rect 562 -2984 563 -2983
rect 800 -2984 801 -2983
rect 1108 -2984 1109 -2983
rect 1269 -2984 1270 -2983
rect 219 -2986 220 -2985
rect 380 -2986 381 -2985
rect 394 -2986 395 -2985
rect 866 -2986 867 -2985
rect 1150 -2986 1151 -2985
rect 1262 -2986 1263 -2985
rect 226 -2988 227 -2987
rect 324 -2988 325 -2987
rect 352 -2988 353 -2987
rect 415 -2988 416 -2987
rect 422 -2988 423 -2987
rect 527 -2988 528 -2987
rect 565 -2988 566 -2987
rect 737 -2988 738 -2987
rect 800 -2988 801 -2987
rect 814 -2988 815 -2987
rect 1094 -2988 1095 -2987
rect 1262 -2988 1263 -2987
rect 170 -2990 171 -2989
rect 226 -2990 227 -2989
rect 233 -2990 234 -2989
rect 310 -2990 311 -2989
rect 355 -2990 356 -2989
rect 478 -2990 479 -2989
rect 506 -2990 507 -2989
rect 814 -2990 815 -2989
rect 1094 -2990 1095 -2989
rect 1192 -2990 1193 -2989
rect 1213 -2990 1214 -2989
rect 1269 -2990 1270 -2989
rect 128 -2992 129 -2991
rect 233 -2992 234 -2991
rect 243 -2992 244 -2991
rect 761 -2992 762 -2991
rect 1157 -2992 1158 -2991
rect 1213 -2992 1214 -2991
rect 1227 -2992 1228 -2991
rect 1304 -2992 1305 -2991
rect 58 -2994 59 -2993
rect 128 -2994 129 -2993
rect 170 -2994 171 -2993
rect 205 -2994 206 -2993
rect 257 -2994 258 -2993
rect 422 -2994 423 -2993
rect 443 -2994 444 -2993
rect 499 -2994 500 -2993
rect 506 -2994 507 -2993
rect 716 -2994 717 -2993
rect 1031 -2994 1032 -2993
rect 1304 -2994 1305 -2993
rect 58 -2996 59 -2995
rect 163 -2996 164 -2995
rect 205 -2996 206 -2995
rect 520 -2996 521 -2995
rect 569 -2996 570 -2995
rect 688 -2996 689 -2995
rect 691 -2996 692 -2995
rect 1087 -2996 1088 -2995
rect 1157 -2996 1158 -2995
rect 1178 -2996 1179 -2995
rect 1192 -2996 1193 -2995
rect 1234 -2996 1235 -2995
rect 86 -2998 87 -2997
rect 443 -2998 444 -2997
rect 450 -2998 451 -2997
rect 548 -2998 549 -2997
rect 569 -2998 570 -2997
rect 583 -2998 584 -2997
rect 590 -2998 591 -2997
rect 740 -2998 741 -2997
rect 1031 -2998 1032 -2997
rect 1066 -2998 1067 -2997
rect 1087 -2998 1088 -2997
rect 1325 -2998 1326 -2997
rect 86 -3000 87 -2999
rect 376 -3000 377 -2999
rect 401 -3000 402 -2999
rect 744 -3000 745 -2999
rect 1066 -3000 1067 -2999
rect 1101 -3000 1102 -2999
rect 1178 -3000 1179 -2999
rect 1381 -3000 1382 -2999
rect 163 -3002 164 -3001
rect 618 -3002 619 -3001
rect 639 -3002 640 -3001
rect 653 -3002 654 -3001
rect 667 -3002 668 -3001
rect 1353 -3002 1354 -3001
rect 1381 -3002 1382 -3001
rect 1416 -3002 1417 -3001
rect 261 -3004 262 -3003
rect 548 -3004 549 -3003
rect 590 -3004 591 -3003
rect 898 -3004 899 -3003
rect 926 -3004 927 -3003
rect 1101 -3004 1102 -3003
rect 1234 -3004 1235 -3003
rect 1339 -3004 1340 -3003
rect 1416 -3004 1417 -3003
rect 1423 -3004 1424 -3003
rect 142 -3006 143 -3005
rect 261 -3006 262 -3005
rect 264 -3006 265 -3005
rect 268 -3006 269 -3005
rect 275 -3006 276 -3005
rect 457 -3006 458 -3005
rect 502 -3006 503 -3005
rect 583 -3006 584 -3005
rect 597 -3006 598 -3005
rect 849 -3006 850 -3005
rect 898 -3006 899 -3005
rect 1223 -3006 1224 -3005
rect 1311 -3006 1312 -3005
rect 1339 -3006 1340 -3005
rect 107 -3008 108 -3007
rect 457 -3008 458 -3007
rect 604 -3008 605 -3007
rect 891 -3008 892 -3007
rect 1311 -3008 1312 -3007
rect 1388 -3008 1389 -3007
rect 107 -3010 108 -3009
rect 492 -3010 493 -3009
rect 611 -3010 612 -3009
rect 926 -3010 927 -3009
rect 142 -3012 143 -3011
rect 184 -3012 185 -3011
rect 264 -3012 265 -3011
rect 772 -3012 773 -3011
rect 891 -3012 892 -3011
rect 919 -3012 920 -3011
rect 184 -3014 185 -3013
rect 191 -3014 192 -3013
rect 268 -3014 269 -3013
rect 338 -3014 339 -3013
rect 359 -3014 360 -3013
rect 625 -3014 626 -3013
rect 639 -3014 640 -3013
rect 1346 -3014 1347 -3013
rect 191 -3016 192 -3015
rect 485 -3016 486 -3015
rect 492 -3016 493 -3015
rect 660 -3016 661 -3015
rect 667 -3016 668 -3015
rect 940 -3016 941 -3015
rect 1346 -3016 1347 -3015
rect 1402 -3016 1403 -3015
rect 282 -3018 283 -3017
rect 772 -3018 773 -3017
rect 940 -3018 941 -3017
rect 961 -3018 962 -3017
rect 282 -3020 283 -3019
rect 331 -3020 332 -3019
rect 338 -3020 339 -3019
rect 345 -3020 346 -3019
rect 401 -3020 402 -3019
rect 471 -3020 472 -3019
rect 485 -3020 486 -3019
rect 733 -3020 734 -3019
rect 807 -3020 808 -3019
rect 961 -3020 962 -3019
rect 296 -3022 297 -3021
rect 359 -3022 360 -3021
rect 404 -3022 405 -3021
rect 513 -3022 514 -3021
rect 576 -3022 577 -3021
rect 919 -3022 920 -3021
rect 296 -3024 297 -3023
rect 835 -3024 836 -3023
rect 317 -3026 318 -3025
rect 576 -3026 577 -3025
rect 618 -3026 619 -3025
rect 975 -3026 976 -3025
rect 303 -3028 304 -3027
rect 317 -3028 318 -3027
rect 331 -3028 332 -3027
rect 481 -3028 482 -3027
rect 660 -3028 661 -3027
rect 709 -3028 710 -3027
rect 716 -3028 717 -3027
rect 779 -3028 780 -3027
rect 303 -3030 304 -3029
rect 999 -3030 1000 -3029
rect 345 -3032 346 -3031
rect 436 -3032 437 -3031
rect 471 -3032 472 -3031
rect 705 -3032 706 -3031
rect 779 -3032 780 -3031
rect 786 -3032 787 -3031
rect 212 -3034 213 -3033
rect 436 -3034 437 -3033
rect 674 -3034 675 -3033
rect 730 -3034 731 -3033
rect 786 -3034 787 -3033
rect 849 -3034 850 -3033
rect 212 -3036 213 -3035
rect 240 -3036 241 -3035
rect 247 -3036 248 -3035
rect 674 -3036 675 -3035
rect 681 -3036 682 -3035
rect 709 -3036 710 -3035
rect 411 -3038 412 -3037
rect 415 -3038 416 -3037
rect 681 -3038 682 -3037
rect 884 -3038 885 -3037
rect 688 -3040 689 -3039
rect 842 -3040 843 -3039
rect 856 -3040 857 -3039
rect 884 -3040 885 -3039
rect 695 -3042 696 -3041
rect 751 -3042 752 -3041
rect 842 -3042 843 -3041
rect 947 -3042 948 -3041
rect 702 -3044 703 -3043
rect 807 -3044 808 -3043
rect 856 -3044 857 -3043
rect 1017 -3044 1018 -3043
rect 705 -3046 706 -3045
rect 1241 -3046 1242 -3045
rect 751 -3048 752 -3047
rect 929 -3048 930 -3047
rect 947 -3048 948 -3047
rect 1010 -3048 1011 -3047
rect 1017 -3048 1018 -3047
rect 1115 -3048 1116 -3047
rect 1010 -3050 1011 -3049
rect 1045 -3050 1046 -3049
rect 1115 -3050 1116 -3049
rect 1206 -3050 1207 -3049
rect 1045 -3052 1046 -3051
rect 1164 -3052 1165 -3051
rect 1206 -3052 1207 -3051
rect 1367 -3052 1368 -3051
rect 1164 -3054 1165 -3053
rect 1220 -3054 1221 -3053
rect 1220 -3056 1221 -3055
rect 1248 -3056 1249 -3055
rect 1248 -3058 1249 -3057
rect 1297 -3058 1298 -3057
rect 1290 -3060 1291 -3059
rect 1297 -3060 1298 -3059
rect 1290 -3062 1291 -3061
rect 1360 -3062 1361 -3061
rect 37 -3073 38 -3072
rect 96 -3073 97 -3072
rect 100 -3073 101 -3072
rect 579 -3073 580 -3072
rect 621 -3073 622 -3072
rect 744 -3073 745 -3072
rect 775 -3073 776 -3072
rect 1248 -3073 1249 -3072
rect 1262 -3073 1263 -3072
rect 1286 -3073 1287 -3072
rect 1293 -3073 1294 -3072
rect 1297 -3073 1298 -3072
rect 1339 -3073 1340 -3072
rect 1353 -3073 1354 -3072
rect 1367 -3073 1368 -3072
rect 1381 -3073 1382 -3072
rect 1409 -3073 1410 -3072
rect 1416 -3073 1417 -3072
rect 1451 -3073 1452 -3072
rect 1458 -3073 1459 -3072
rect 44 -3075 45 -3074
rect 219 -3075 220 -3074
rect 240 -3075 241 -3074
rect 982 -3075 983 -3074
rect 1010 -3075 1011 -3074
rect 1087 -3075 1088 -3074
rect 1090 -3075 1091 -3074
rect 1269 -3075 1270 -3074
rect 1283 -3075 1284 -3074
rect 1346 -3075 1347 -3074
rect 1458 -3075 1459 -3074
rect 1465 -3075 1466 -3074
rect 51 -3077 52 -3076
rect 215 -3077 216 -3076
rect 226 -3077 227 -3076
rect 240 -3077 241 -3076
rect 243 -3077 244 -3076
rect 338 -3077 339 -3076
rect 373 -3077 374 -3076
rect 621 -3077 622 -3076
rect 639 -3077 640 -3076
rect 807 -3077 808 -3076
rect 849 -3077 850 -3076
rect 968 -3077 969 -3076
rect 982 -3077 983 -3076
rect 1115 -3077 1116 -3076
rect 1220 -3077 1221 -3076
rect 1290 -3077 1291 -3076
rect 1346 -3077 1347 -3076
rect 1374 -3077 1375 -3076
rect 1465 -3077 1466 -3076
rect 1472 -3077 1473 -3076
rect 58 -3079 59 -3078
rect 180 -3079 181 -3078
rect 191 -3079 192 -3078
rect 250 -3079 251 -3078
rect 289 -3079 290 -3078
rect 607 -3079 608 -3078
rect 653 -3079 654 -3078
rect 705 -3079 706 -3078
rect 740 -3079 741 -3078
rect 968 -3079 969 -3078
rect 1010 -3079 1011 -3078
rect 1052 -3079 1053 -3078
rect 1059 -3079 1060 -3078
rect 1241 -3079 1242 -3078
rect 1262 -3079 1263 -3078
rect 1332 -3079 1333 -3078
rect 72 -3081 73 -3080
rect 187 -3081 188 -3080
rect 191 -3081 192 -3080
rect 268 -3081 269 -3080
rect 299 -3081 300 -3080
rect 324 -3081 325 -3080
rect 338 -3081 339 -3080
rect 464 -3081 465 -3080
rect 513 -3081 514 -3080
rect 737 -3081 738 -3080
rect 744 -3081 745 -3080
rect 800 -3081 801 -3080
rect 807 -3081 808 -3080
rect 856 -3081 857 -3080
rect 870 -3081 871 -3080
rect 947 -3081 948 -3080
rect 961 -3081 962 -3080
rect 1136 -3081 1137 -3080
rect 1164 -3081 1165 -3080
rect 1220 -3081 1221 -3080
rect 1230 -3081 1231 -3080
rect 1311 -3081 1312 -3080
rect 79 -3083 80 -3082
rect 408 -3083 409 -3082
rect 436 -3083 437 -3082
rect 1062 -3083 1063 -3082
rect 1066 -3083 1067 -3082
rect 1115 -3083 1116 -3082
rect 1136 -3083 1137 -3082
rect 1234 -3083 1235 -3082
rect 79 -3085 80 -3084
rect 93 -3085 94 -3084
rect 100 -3085 101 -3084
rect 114 -3085 115 -3084
rect 121 -3085 122 -3084
rect 737 -3085 738 -3084
rect 782 -3085 783 -3084
rect 1038 -3085 1039 -3084
rect 1052 -3085 1053 -3084
rect 1255 -3085 1256 -3084
rect 86 -3087 87 -3086
rect 355 -3087 356 -3086
rect 373 -3087 374 -3086
rect 471 -3087 472 -3086
rect 478 -3087 479 -3086
rect 800 -3087 801 -3086
rect 873 -3087 874 -3086
rect 905 -3087 906 -3086
rect 929 -3087 930 -3086
rect 1276 -3087 1277 -3086
rect 65 -3089 66 -3088
rect 86 -3089 87 -3088
rect 93 -3089 94 -3088
rect 163 -3089 164 -3088
rect 177 -3089 178 -3088
rect 415 -3089 416 -3088
rect 436 -3089 437 -3088
rect 520 -3089 521 -3088
rect 523 -3089 524 -3088
rect 877 -3089 878 -3088
rect 884 -3089 885 -3088
rect 919 -3089 920 -3088
rect 933 -3089 934 -3088
rect 947 -3089 948 -3088
rect 964 -3089 965 -3088
rect 1185 -3089 1186 -3088
rect 1276 -3089 1277 -3088
rect 1325 -3089 1326 -3088
rect 114 -3091 115 -3090
rect 128 -3091 129 -3090
rect 142 -3091 143 -3090
rect 222 -3091 223 -3090
rect 226 -3091 227 -3090
rect 635 -3091 636 -3090
rect 656 -3091 657 -3090
rect 828 -3091 829 -3090
rect 884 -3091 885 -3090
rect 891 -3091 892 -3090
rect 905 -3091 906 -3090
rect 964 -3091 965 -3090
rect 996 -3091 997 -3090
rect 1038 -3091 1039 -3090
rect 1066 -3091 1067 -3090
rect 1094 -3091 1095 -3090
rect 1101 -3091 1102 -3090
rect 1290 -3091 1291 -3090
rect 121 -3093 122 -3092
rect 156 -3093 157 -3092
rect 163 -3093 164 -3092
rect 205 -3093 206 -3092
rect 247 -3093 248 -3092
rect 362 -3093 363 -3092
rect 366 -3093 367 -3092
rect 478 -3093 479 -3092
rect 520 -3093 521 -3092
rect 611 -3093 612 -3092
rect 618 -3093 619 -3092
rect 877 -3093 878 -3092
rect 912 -3093 913 -3092
rect 933 -3093 934 -3092
rect 940 -3093 941 -3092
rect 961 -3093 962 -3092
rect 975 -3093 976 -3092
rect 1094 -3093 1095 -3092
rect 1101 -3093 1102 -3092
rect 1199 -3093 1200 -3092
rect 142 -3095 143 -3094
rect 170 -3095 171 -3094
rect 177 -3095 178 -3094
rect 184 -3095 185 -3094
rect 198 -3095 199 -3094
rect 688 -3095 689 -3094
rect 702 -3095 703 -3094
rect 1073 -3095 1074 -3094
rect 1129 -3095 1130 -3094
rect 1199 -3095 1200 -3094
rect 156 -3097 157 -3096
rect 296 -3097 297 -3096
rect 303 -3097 304 -3096
rect 513 -3097 514 -3096
rect 527 -3097 528 -3096
rect 919 -3097 920 -3096
rect 940 -3097 941 -3096
rect 954 -3097 955 -3096
rect 1073 -3097 1074 -3096
rect 1206 -3097 1207 -3096
rect 128 -3099 129 -3098
rect 303 -3099 304 -3098
rect 366 -3099 367 -3098
rect 856 -3099 857 -3098
rect 898 -3099 899 -3098
rect 954 -3099 955 -3098
rect 1164 -3099 1165 -3098
rect 1223 -3099 1224 -3098
rect 170 -3101 171 -3100
rect 275 -3101 276 -3100
rect 296 -3101 297 -3100
rect 387 -3101 388 -3100
rect 394 -3101 395 -3100
rect 415 -3101 416 -3100
rect 464 -3101 465 -3100
rect 642 -3101 643 -3100
rect 674 -3101 675 -3100
rect 870 -3101 871 -3100
rect 898 -3101 899 -3100
rect 1031 -3101 1032 -3100
rect 1206 -3101 1207 -3100
rect 1304 -3101 1305 -3100
rect 198 -3103 199 -3102
rect 282 -3103 283 -3102
rect 352 -3103 353 -3102
rect 674 -3103 675 -3102
rect 684 -3103 685 -3102
rect 772 -3103 773 -3102
rect 786 -3103 787 -3102
rect 849 -3103 850 -3102
rect 912 -3103 913 -3102
rect 1080 -3103 1081 -3102
rect 201 -3105 202 -3104
rect 324 -3105 325 -3104
rect 352 -3105 353 -3104
rect 429 -3105 430 -3104
rect 471 -3105 472 -3104
rect 597 -3105 598 -3104
rect 765 -3105 766 -3104
rect 786 -3105 787 -3104
rect 793 -3105 794 -3104
rect 1024 -3105 1025 -3104
rect 1031 -3105 1032 -3104
rect 1108 -3105 1109 -3104
rect 233 -3107 234 -3106
rect 247 -3107 248 -3106
rect 261 -3107 262 -3106
rect 394 -3107 395 -3106
rect 401 -3107 402 -3106
rect 845 -3107 846 -3106
rect 1024 -3107 1025 -3106
rect 1122 -3107 1123 -3106
rect 212 -3109 213 -3108
rect 261 -3109 262 -3108
rect 268 -3109 269 -3108
rect 310 -3109 311 -3108
rect 380 -3109 381 -3108
rect 383 -3109 384 -3108
rect 387 -3109 388 -3108
rect 681 -3109 682 -3108
rect 723 -3109 724 -3108
rect 765 -3109 766 -3108
rect 796 -3109 797 -3108
rect 880 -3109 881 -3108
rect 1080 -3109 1081 -3108
rect 1227 -3109 1228 -3108
rect 222 -3111 223 -3110
rect 401 -3111 402 -3110
rect 408 -3111 409 -3110
rect 485 -3111 486 -3110
rect 506 -3111 507 -3110
rect 597 -3111 598 -3110
rect 681 -3111 682 -3110
rect 695 -3111 696 -3110
rect 723 -3111 724 -3110
rect 758 -3111 759 -3110
rect 835 -3111 836 -3110
rect 891 -3111 892 -3110
rect 1108 -3111 1109 -3110
rect 1150 -3111 1151 -3110
rect 233 -3113 234 -3112
rect 331 -3113 332 -3112
rect 380 -3113 381 -3112
rect 604 -3113 605 -3112
rect 695 -3113 696 -3112
rect 709 -3113 710 -3112
rect 758 -3113 759 -3112
rect 842 -3113 843 -3112
rect 1122 -3113 1123 -3112
rect 1178 -3113 1179 -3112
rect 275 -3115 276 -3114
rect 345 -3115 346 -3114
rect 485 -3115 486 -3114
rect 653 -3115 654 -3114
rect 709 -3115 710 -3114
rect 730 -3115 731 -3114
rect 828 -3115 829 -3114
rect 842 -3115 843 -3114
rect 1129 -3115 1130 -3114
rect 1227 -3115 1228 -3114
rect 282 -3117 283 -3116
rect 555 -3117 556 -3116
rect 576 -3117 577 -3116
rect 611 -3117 612 -3116
rect 835 -3117 836 -3116
rect 926 -3117 927 -3116
rect 1150 -3117 1151 -3116
rect 1188 -3117 1189 -3116
rect 289 -3119 290 -3118
rect 730 -3119 731 -3118
rect 814 -3119 815 -3118
rect 926 -3119 927 -3118
rect 1178 -3119 1179 -3118
rect 1192 -3119 1193 -3118
rect 310 -3121 311 -3120
rect 457 -3121 458 -3120
rect 506 -3121 507 -3120
rect 632 -3121 633 -3120
rect 814 -3121 815 -3120
rect 821 -3121 822 -3120
rect 1192 -3121 1193 -3120
rect 1318 -3121 1319 -3120
rect 317 -3123 318 -3122
rect 331 -3123 332 -3122
rect 345 -3123 346 -3122
rect 359 -3123 360 -3122
rect 457 -3123 458 -3122
rect 772 -3123 773 -3122
rect 821 -3123 822 -3122
rect 1045 -3123 1046 -3122
rect 135 -3125 136 -3124
rect 317 -3125 318 -3124
rect 527 -3125 528 -3124
rect 625 -3125 626 -3124
rect 1045 -3125 1046 -3124
rect 1213 -3125 1214 -3124
rect 205 -3127 206 -3126
rect 359 -3127 360 -3126
rect 534 -3127 535 -3126
rect 632 -3127 633 -3126
rect 1157 -3127 1158 -3126
rect 1213 -3127 1214 -3126
rect 450 -3129 451 -3128
rect 534 -3129 535 -3128
rect 541 -3129 542 -3128
rect 555 -3129 556 -3128
rect 583 -3129 584 -3128
rect 793 -3129 794 -3128
rect 1157 -3129 1158 -3128
rect 1241 -3129 1242 -3128
rect 450 -3131 451 -3130
rect 548 -3131 549 -3130
rect 604 -3131 605 -3130
rect 863 -3131 864 -3130
rect 422 -3133 423 -3132
rect 548 -3133 549 -3132
rect 625 -3133 626 -3132
rect 716 -3133 717 -3132
rect 863 -3133 864 -3132
rect 989 -3133 990 -3132
rect 422 -3135 423 -3134
rect 576 -3135 577 -3134
rect 716 -3135 717 -3134
rect 779 -3135 780 -3134
rect 989 -3135 990 -3134
rect 1003 -3135 1004 -3134
rect 492 -3137 493 -3136
rect 1003 -3137 1004 -3136
rect 443 -3139 444 -3138
rect 492 -3139 493 -3138
rect 499 -3139 500 -3138
rect 583 -3139 584 -3138
rect 779 -3139 780 -3138
rect 975 -3139 976 -3138
rect 383 -3141 384 -3140
rect 443 -3141 444 -3140
rect 499 -3141 500 -3140
rect 569 -3141 570 -3140
rect 541 -3143 542 -3142
rect 646 -3143 647 -3142
rect 562 -3145 563 -3144
rect 646 -3145 647 -3144
rect 562 -3147 563 -3146
rect 751 -3147 752 -3146
rect 569 -3149 570 -3148
rect 660 -3149 661 -3148
rect 667 -3149 668 -3148
rect 751 -3149 752 -3148
rect 135 -3151 136 -3150
rect 660 -3151 661 -3150
rect 667 -3151 668 -3150
rect 705 -3151 706 -3150
rect 58 -3162 59 -3161
rect 198 -3162 199 -3161
rect 219 -3162 220 -3161
rect 352 -3162 353 -3161
rect 373 -3162 374 -3161
rect 429 -3162 430 -3161
rect 432 -3162 433 -3161
rect 555 -3162 556 -3161
rect 569 -3162 570 -3161
rect 579 -3162 580 -3161
rect 611 -3162 612 -3161
rect 663 -3162 664 -3161
rect 667 -3162 668 -3161
rect 779 -3162 780 -3161
rect 793 -3162 794 -3161
rect 842 -3162 843 -3161
rect 845 -3162 846 -3161
rect 1017 -3162 1018 -3161
rect 1080 -3162 1081 -3161
rect 1087 -3162 1088 -3161
rect 1094 -3162 1095 -3161
rect 1097 -3162 1098 -3161
rect 1188 -3162 1189 -3161
rect 1262 -3162 1263 -3161
rect 1332 -3162 1333 -3161
rect 1346 -3162 1347 -3161
rect 1353 -3162 1354 -3161
rect 1360 -3162 1361 -3161
rect 65 -3164 66 -3163
rect 135 -3164 136 -3163
rect 145 -3164 146 -3163
rect 187 -3164 188 -3163
rect 306 -3164 307 -3163
rect 338 -3164 339 -3163
rect 352 -3164 353 -3163
rect 387 -3164 388 -3163
rect 415 -3164 416 -3163
rect 418 -3164 419 -3163
rect 471 -3164 472 -3163
rect 635 -3164 636 -3163
rect 653 -3164 654 -3163
rect 737 -3164 738 -3163
rect 751 -3164 752 -3163
rect 793 -3164 794 -3163
rect 856 -3164 857 -3163
rect 1052 -3164 1053 -3163
rect 1080 -3164 1081 -3163
rect 1108 -3164 1109 -3163
rect 1220 -3164 1221 -3163
rect 1241 -3164 1242 -3163
rect 72 -3166 73 -3165
rect 205 -3166 206 -3165
rect 296 -3166 297 -3165
rect 338 -3166 339 -3165
rect 373 -3166 374 -3165
rect 499 -3166 500 -3165
rect 513 -3166 514 -3165
rect 611 -3166 612 -3165
rect 618 -3166 619 -3165
rect 709 -3166 710 -3165
rect 716 -3166 717 -3165
rect 737 -3166 738 -3165
rect 761 -3166 762 -3165
rect 772 -3166 773 -3165
rect 775 -3166 776 -3165
rect 835 -3166 836 -3165
rect 856 -3166 857 -3165
rect 870 -3166 871 -3165
rect 877 -3166 878 -3165
rect 968 -3166 969 -3165
rect 985 -3166 986 -3165
rect 1122 -3166 1123 -3165
rect 1227 -3166 1228 -3165
rect 1234 -3166 1235 -3165
rect 1237 -3166 1238 -3165
rect 1276 -3166 1277 -3165
rect 79 -3168 80 -3167
rect 215 -3168 216 -3167
rect 250 -3168 251 -3167
rect 716 -3168 717 -3167
rect 733 -3168 734 -3167
rect 912 -3168 913 -3167
rect 919 -3168 920 -3167
rect 1052 -3168 1053 -3167
rect 1094 -3168 1095 -3167
rect 1129 -3168 1130 -3167
rect 79 -3170 80 -3169
rect 156 -3170 157 -3169
rect 180 -3170 181 -3169
rect 667 -3170 668 -3169
rect 688 -3170 689 -3169
rect 891 -3170 892 -3169
rect 912 -3170 913 -3169
rect 947 -3170 948 -3169
rect 964 -3170 965 -3169
rect 989 -3170 990 -3169
rect 999 -3170 1000 -3169
rect 1038 -3170 1039 -3169
rect 1122 -3170 1123 -3169
rect 1192 -3170 1193 -3169
rect 93 -3172 94 -3171
rect 205 -3172 206 -3171
rect 327 -3172 328 -3171
rect 362 -3172 363 -3171
rect 387 -3172 388 -3171
rect 656 -3172 657 -3171
rect 660 -3172 661 -3171
rect 821 -3172 822 -3171
rect 835 -3172 836 -3171
rect 954 -3172 955 -3171
rect 968 -3172 969 -3171
rect 1059 -3172 1060 -3171
rect 1129 -3172 1130 -3171
rect 1136 -3172 1137 -3171
rect 1192 -3172 1193 -3171
rect 1293 -3172 1294 -3171
rect 93 -3174 94 -3173
rect 170 -3174 171 -3173
rect 201 -3174 202 -3173
rect 296 -3174 297 -3173
rect 401 -3174 402 -3173
rect 471 -3174 472 -3173
rect 492 -3174 493 -3173
rect 499 -3174 500 -3173
rect 534 -3174 535 -3173
rect 537 -3174 538 -3173
rect 541 -3174 542 -3173
rect 866 -3174 867 -3173
rect 870 -3174 871 -3173
rect 898 -3174 899 -3173
rect 933 -3174 934 -3173
rect 947 -3174 948 -3173
rect 989 -3174 990 -3173
rect 1045 -3174 1046 -3173
rect 100 -3176 101 -3175
rect 152 -3176 153 -3175
rect 156 -3176 157 -3175
rect 191 -3176 192 -3175
rect 324 -3176 325 -3175
rect 401 -3176 402 -3175
rect 415 -3176 416 -3175
rect 464 -3176 465 -3175
rect 534 -3176 535 -3175
rect 548 -3176 549 -3175
rect 569 -3176 570 -3175
rect 807 -3176 808 -3175
rect 863 -3176 864 -3175
rect 919 -3176 920 -3175
rect 933 -3176 934 -3175
rect 1031 -3176 1032 -3175
rect 1045 -3176 1046 -3175
rect 1073 -3176 1074 -3175
rect 100 -3178 101 -3177
rect 264 -3178 265 -3177
rect 268 -3178 269 -3177
rect 324 -3178 325 -3177
rect 422 -3178 423 -3177
rect 513 -3178 514 -3177
rect 541 -3178 542 -3177
rect 646 -3178 647 -3177
rect 660 -3178 661 -3177
rect 1024 -3178 1025 -3177
rect 1031 -3178 1032 -3177
rect 1244 -3178 1245 -3177
rect 114 -3180 115 -3179
rect 208 -3180 209 -3179
rect 247 -3180 248 -3179
rect 268 -3180 269 -3179
rect 422 -3180 423 -3179
rect 443 -3180 444 -3179
rect 464 -3180 465 -3179
rect 485 -3180 486 -3179
rect 492 -3180 493 -3179
rect 863 -3180 864 -3179
rect 880 -3180 881 -3179
rect 898 -3180 899 -3179
rect 940 -3180 941 -3179
rect 954 -3180 955 -3179
rect 1006 -3180 1007 -3179
rect 1066 -3180 1067 -3179
rect 1073 -3180 1074 -3179
rect 1150 -3180 1151 -3179
rect 121 -3182 122 -3181
rect 198 -3182 199 -3181
rect 436 -3182 437 -3181
rect 772 -3182 773 -3181
rect 779 -3182 780 -3181
rect 926 -3182 927 -3181
rect 1010 -3182 1011 -3181
rect 1038 -3182 1039 -3181
rect 1115 -3182 1116 -3181
rect 1150 -3182 1151 -3181
rect 121 -3184 122 -3183
rect 226 -3184 227 -3183
rect 282 -3184 283 -3183
rect 436 -3184 437 -3183
rect 443 -3184 444 -3183
rect 702 -3184 703 -3183
rect 705 -3184 706 -3183
rect 1017 -3184 1018 -3183
rect 1024 -3184 1025 -3183
rect 1157 -3184 1158 -3183
rect 131 -3186 132 -3185
rect 184 -3186 185 -3185
rect 282 -3186 283 -3185
rect 345 -3186 346 -3185
rect 485 -3186 486 -3185
rect 520 -3186 521 -3185
rect 548 -3186 549 -3185
rect 674 -3186 675 -3185
rect 681 -3186 682 -3185
rect 688 -3186 689 -3185
rect 695 -3186 696 -3185
rect 709 -3186 710 -3185
rect 765 -3186 766 -3185
rect 821 -3186 822 -3185
rect 884 -3186 885 -3185
rect 996 -3186 997 -3185
rect 1115 -3186 1116 -3185
rect 1185 -3186 1186 -3185
rect 135 -3188 136 -3187
rect 457 -3188 458 -3187
rect 506 -3188 507 -3187
rect 681 -3188 682 -3187
rect 800 -3188 801 -3187
rect 891 -3188 892 -3187
rect 905 -3188 906 -3187
rect 940 -3188 941 -3187
rect 1097 -3188 1098 -3187
rect 1136 -3188 1137 -3187
rect 1143 -3188 1144 -3187
rect 1185 -3188 1186 -3187
rect 142 -3190 143 -3189
rect 191 -3190 192 -3189
rect 331 -3190 332 -3189
rect 345 -3190 346 -3189
rect 359 -3190 360 -3189
rect 996 -3190 997 -3189
rect 1143 -3190 1144 -3189
rect 1164 -3190 1165 -3189
rect 86 -3192 87 -3191
rect 142 -3192 143 -3191
rect 149 -3192 150 -3191
rect 194 -3192 195 -3191
rect 359 -3192 360 -3191
rect 394 -3192 395 -3191
rect 408 -3192 409 -3191
rect 457 -3192 458 -3191
rect 506 -3192 507 -3191
rect 583 -3192 584 -3191
rect 597 -3192 598 -3191
rect 618 -3192 619 -3191
rect 625 -3192 626 -3191
rect 695 -3192 696 -3191
rect 786 -3192 787 -3191
rect 800 -3192 801 -3191
rect 807 -3192 808 -3191
rect 814 -3192 815 -3191
rect 884 -3192 885 -3191
rect 961 -3192 962 -3191
rect 1157 -3192 1158 -3191
rect 1171 -3192 1172 -3191
rect 86 -3194 87 -3193
rect 107 -3194 108 -3193
rect 163 -3194 164 -3193
rect 331 -3194 332 -3193
rect 380 -3194 381 -3193
rect 394 -3194 395 -3193
rect 478 -3194 479 -3193
rect 597 -3194 598 -3193
rect 607 -3194 608 -3193
rect 1010 -3194 1011 -3193
rect 1164 -3194 1165 -3193
rect 1178 -3194 1179 -3193
rect 107 -3196 108 -3195
rect 233 -3196 234 -3195
rect 303 -3196 304 -3195
rect 625 -3196 626 -3195
rect 632 -3196 633 -3195
rect 1003 -3196 1004 -3195
rect 1171 -3196 1172 -3195
rect 1206 -3196 1207 -3195
rect 163 -3198 164 -3197
rect 254 -3198 255 -3197
rect 317 -3198 318 -3197
rect 408 -3198 409 -3197
rect 562 -3198 563 -3197
rect 702 -3198 703 -3197
rect 730 -3198 731 -3197
rect 786 -3198 787 -3197
rect 814 -3198 815 -3197
rect 849 -3198 850 -3197
rect 905 -3198 906 -3197
rect 1111 -3198 1112 -3197
rect 1167 -3198 1168 -3197
rect 1206 -3198 1207 -3197
rect 173 -3200 174 -3199
rect 226 -3200 227 -3199
rect 254 -3200 255 -3199
rect 261 -3200 262 -3199
rect 366 -3200 367 -3199
rect 380 -3200 381 -3199
rect 527 -3200 528 -3199
rect 562 -3200 563 -3199
rect 583 -3200 584 -3199
rect 590 -3200 591 -3199
rect 639 -3200 640 -3199
rect 751 -3200 752 -3199
rect 828 -3200 829 -3199
rect 849 -3200 850 -3199
rect 926 -3200 927 -3199
rect 982 -3200 983 -3199
rect 212 -3202 213 -3201
rect 317 -3202 318 -3201
rect 366 -3202 367 -3201
rect 604 -3202 605 -3201
rect 632 -3202 633 -3201
rect 639 -3202 640 -3201
rect 646 -3202 647 -3201
rect 782 -3202 783 -3201
rect 828 -3202 829 -3201
rect 1003 -3202 1004 -3201
rect 177 -3204 178 -3203
rect 212 -3204 213 -3203
rect 222 -3204 223 -3203
rect 233 -3204 234 -3203
rect 310 -3204 311 -3203
rect 604 -3204 605 -3203
rect 730 -3204 731 -3203
rect 744 -3204 745 -3203
rect 961 -3204 962 -3203
rect 1059 -3204 1060 -3203
rect 240 -3206 241 -3205
rect 310 -3206 311 -3205
rect 450 -3206 451 -3205
rect 527 -3206 528 -3205
rect 555 -3206 556 -3205
rect 590 -3206 591 -3205
rect 744 -3206 745 -3205
rect 758 -3206 759 -3205
rect 240 -3208 241 -3207
rect 275 -3208 276 -3207
rect 289 -3208 290 -3207
rect 450 -3208 451 -3207
rect 478 -3208 479 -3207
rect 982 -3208 983 -3207
rect 247 -3210 248 -3209
rect 289 -3210 290 -3209
rect 758 -3210 759 -3209
rect 765 -3210 766 -3209
rect 261 -3212 262 -3211
rect 275 -3212 276 -3211
rect 58 -3223 59 -3222
rect 247 -3223 248 -3222
rect 338 -3223 339 -3222
rect 341 -3223 342 -3222
rect 359 -3223 360 -3222
rect 362 -3223 363 -3222
rect 380 -3223 381 -3222
rect 397 -3223 398 -3222
rect 408 -3223 409 -3222
rect 663 -3223 664 -3222
rect 702 -3223 703 -3222
rect 758 -3223 759 -3222
rect 782 -3223 783 -3222
rect 1031 -3223 1032 -3222
rect 1038 -3223 1039 -3222
rect 1062 -3223 1063 -3222
rect 1066 -3223 1067 -3222
rect 1080 -3223 1081 -3222
rect 1101 -3223 1102 -3222
rect 1111 -3223 1112 -3222
rect 1136 -3223 1137 -3222
rect 1157 -3223 1158 -3222
rect 1206 -3223 1207 -3222
rect 1251 -3223 1252 -3222
rect 1290 -3223 1291 -3222
rect 1325 -3223 1326 -3222
rect 1328 -3223 1329 -3222
rect 1332 -3223 1333 -3222
rect 1451 -3223 1452 -3222
rect 1454 -3223 1455 -3222
rect 65 -3225 66 -3224
rect 261 -3225 262 -3224
rect 338 -3225 339 -3224
rect 345 -3225 346 -3224
rect 359 -3225 360 -3224
rect 443 -3225 444 -3224
rect 464 -3225 465 -3224
rect 579 -3225 580 -3224
rect 604 -3225 605 -3224
rect 919 -3225 920 -3224
rect 982 -3225 983 -3224
rect 1216 -3225 1217 -3224
rect 1451 -3225 1452 -3224
rect 1458 -3225 1459 -3224
rect 72 -3227 73 -3226
rect 117 -3227 118 -3226
rect 121 -3227 122 -3226
rect 324 -3227 325 -3226
rect 380 -3227 381 -3226
rect 415 -3227 416 -3226
rect 429 -3227 430 -3226
rect 488 -3227 489 -3226
rect 534 -3227 535 -3226
rect 537 -3227 538 -3226
rect 548 -3227 549 -3226
rect 726 -3227 727 -3226
rect 737 -3227 738 -3226
rect 863 -3227 864 -3226
rect 866 -3227 867 -3226
rect 933 -3227 934 -3226
rect 982 -3227 983 -3226
rect 989 -3227 990 -3226
rect 992 -3227 993 -3226
rect 1045 -3227 1046 -3226
rect 1052 -3227 1053 -3226
rect 1101 -3227 1102 -3226
rect 1125 -3227 1126 -3226
rect 1136 -3227 1137 -3226
rect 1150 -3227 1151 -3226
rect 1188 -3227 1189 -3226
rect 1213 -3227 1214 -3226
rect 1220 -3227 1221 -3226
rect 79 -3229 80 -3228
rect 173 -3229 174 -3228
rect 177 -3229 178 -3228
rect 191 -3229 192 -3228
rect 201 -3229 202 -3228
rect 387 -3229 388 -3228
rect 422 -3229 423 -3228
rect 429 -3229 430 -3228
rect 443 -3229 444 -3228
rect 457 -3229 458 -3228
rect 534 -3229 535 -3228
rect 646 -3229 647 -3228
rect 730 -3229 731 -3228
rect 737 -3229 738 -3228
rect 758 -3229 759 -3228
rect 765 -3229 766 -3228
rect 786 -3229 787 -3228
rect 1003 -3229 1004 -3228
rect 1017 -3229 1018 -3228
rect 1167 -3229 1168 -3228
rect 1185 -3229 1186 -3228
rect 1206 -3229 1207 -3228
rect 86 -3231 87 -3230
rect 128 -3231 129 -3230
rect 131 -3231 132 -3230
rect 324 -3231 325 -3230
rect 352 -3231 353 -3230
rect 415 -3231 416 -3230
rect 450 -3231 451 -3230
rect 457 -3231 458 -3230
rect 541 -3231 542 -3230
rect 646 -3231 647 -3230
rect 733 -3231 734 -3230
rect 786 -3231 787 -3230
rect 849 -3231 850 -3230
rect 985 -3231 986 -3230
rect 996 -3231 997 -3230
rect 1108 -3231 1109 -3230
rect 1150 -3231 1151 -3230
rect 1171 -3231 1172 -3230
rect 1185 -3231 1186 -3230
rect 1199 -3231 1200 -3230
rect 93 -3233 94 -3232
rect 180 -3233 181 -3232
rect 187 -3233 188 -3232
rect 366 -3233 367 -3232
rect 387 -3233 388 -3232
rect 401 -3233 402 -3232
rect 450 -3233 451 -3232
rect 471 -3233 472 -3232
rect 548 -3233 549 -3232
rect 597 -3233 598 -3232
rect 604 -3233 605 -3232
rect 632 -3233 633 -3232
rect 639 -3233 640 -3232
rect 702 -3233 703 -3232
rect 765 -3233 766 -3232
rect 828 -3233 829 -3232
rect 880 -3233 881 -3232
rect 926 -3233 927 -3232
rect 933 -3233 934 -3232
rect 968 -3233 969 -3232
rect 996 -3233 997 -3232
rect 1164 -3233 1165 -3232
rect 100 -3235 101 -3234
rect 243 -3235 244 -3234
rect 247 -3235 248 -3234
rect 275 -3235 276 -3234
rect 282 -3235 283 -3234
rect 352 -3235 353 -3234
rect 366 -3235 367 -3234
rect 404 -3235 405 -3234
rect 474 -3235 475 -3234
rect 597 -3235 598 -3234
rect 611 -3235 612 -3234
rect 639 -3235 640 -3234
rect 807 -3235 808 -3234
rect 828 -3235 829 -3234
rect 898 -3235 899 -3234
rect 926 -3235 927 -3234
rect 940 -3235 941 -3234
rect 1003 -3235 1004 -3234
rect 1059 -3235 1060 -3234
rect 1122 -3235 1123 -3234
rect 1160 -3235 1161 -3234
rect 1171 -3235 1172 -3234
rect 114 -3237 115 -3236
rect 492 -3237 493 -3236
rect 555 -3237 556 -3236
rect 891 -3237 892 -3236
rect 898 -3237 899 -3236
rect 912 -3237 913 -3236
rect 919 -3237 920 -3236
rect 1122 -3237 1123 -3236
rect 1164 -3237 1165 -3236
rect 1192 -3237 1193 -3236
rect 135 -3239 136 -3238
rect 170 -3239 171 -3238
rect 191 -3239 192 -3238
rect 401 -3239 402 -3238
rect 555 -3239 556 -3238
rect 562 -3239 563 -3238
rect 569 -3239 570 -3238
rect 576 -3239 577 -3238
rect 611 -3239 612 -3238
rect 653 -3239 654 -3238
rect 800 -3239 801 -3238
rect 807 -3239 808 -3238
rect 856 -3239 857 -3238
rect 891 -3239 892 -3238
rect 940 -3239 941 -3238
rect 954 -3239 955 -3238
rect 1080 -3239 1081 -3238
rect 1115 -3239 1116 -3238
rect 149 -3241 150 -3240
rect 464 -3241 465 -3240
rect 527 -3241 528 -3240
rect 569 -3241 570 -3240
rect 618 -3241 619 -3240
rect 625 -3241 626 -3240
rect 628 -3241 629 -3240
rect 744 -3241 745 -3240
rect 793 -3241 794 -3240
rect 800 -3241 801 -3240
rect 884 -3241 885 -3240
rect 912 -3241 913 -3240
rect 947 -3241 948 -3240
rect 954 -3241 955 -3240
rect 1087 -3241 1088 -3240
rect 1108 -3241 1109 -3240
rect 152 -3243 153 -3242
rect 576 -3243 577 -3242
rect 618 -3243 619 -3242
rect 635 -3243 636 -3242
rect 653 -3243 654 -3242
rect 688 -3243 689 -3242
rect 744 -3243 745 -3242
rect 751 -3243 752 -3242
rect 793 -3243 794 -3242
rect 821 -3243 822 -3242
rect 842 -3243 843 -3242
rect 947 -3243 948 -3242
rect 226 -3245 227 -3244
rect 229 -3245 230 -3244
rect 264 -3245 265 -3244
rect 275 -3245 276 -3244
rect 296 -3245 297 -3244
rect 422 -3245 423 -3244
rect 513 -3245 514 -3244
rect 527 -3245 528 -3244
rect 558 -3245 559 -3244
rect 674 -3245 675 -3244
rect 751 -3245 752 -3244
rect 779 -3245 780 -3244
rect 821 -3245 822 -3244
rect 961 -3245 962 -3244
rect 107 -3247 108 -3246
rect 264 -3247 265 -3246
rect 268 -3247 269 -3246
rect 282 -3247 283 -3246
rect 296 -3247 297 -3246
rect 303 -3247 304 -3246
rect 394 -3247 395 -3246
rect 632 -3247 633 -3246
rect 635 -3247 636 -3246
rect 772 -3247 773 -3246
rect 842 -3247 843 -3246
rect 870 -3247 871 -3246
rect 884 -3247 885 -3246
rect 905 -3247 906 -3246
rect 961 -3247 962 -3246
rect 1024 -3247 1025 -3246
rect 156 -3249 157 -3248
rect 394 -3249 395 -3248
rect 506 -3249 507 -3248
rect 513 -3249 514 -3248
rect 562 -3249 563 -3248
rect 583 -3249 584 -3248
rect 660 -3249 661 -3248
rect 688 -3249 689 -3248
rect 772 -3249 773 -3248
rect 814 -3249 815 -3248
rect 870 -3249 871 -3248
rect 877 -3249 878 -3248
rect 905 -3249 906 -3248
rect 975 -3249 976 -3248
rect 156 -3251 157 -3250
rect 261 -3251 262 -3250
rect 268 -3251 269 -3250
rect 289 -3251 290 -3250
rect 436 -3251 437 -3250
rect 583 -3251 584 -3250
rect 660 -3251 661 -3250
rect 695 -3251 696 -3250
rect 877 -3251 878 -3250
rect 1010 -3251 1011 -3250
rect 198 -3253 199 -3252
rect 289 -3253 290 -3252
rect 373 -3253 374 -3252
rect 436 -3253 437 -3252
rect 506 -3253 507 -3252
rect 607 -3253 608 -3252
rect 667 -3253 668 -3252
rect 814 -3253 815 -3252
rect 184 -3255 185 -3254
rect 198 -3255 199 -3254
rect 219 -3255 220 -3254
rect 303 -3255 304 -3254
rect 331 -3255 332 -3254
rect 373 -3255 374 -3254
rect 590 -3255 591 -3254
rect 695 -3255 696 -3254
rect 212 -3257 213 -3256
rect 219 -3257 220 -3256
rect 226 -3257 227 -3256
rect 254 -3257 255 -3256
rect 310 -3257 311 -3256
rect 331 -3257 332 -3256
rect 667 -3257 668 -3256
rect 716 -3257 717 -3256
rect 212 -3259 213 -3258
rect 233 -3259 234 -3258
rect 310 -3259 311 -3258
rect 478 -3259 479 -3258
rect 674 -3259 675 -3258
rect 681 -3259 682 -3258
rect 709 -3259 710 -3258
rect 716 -3259 717 -3258
rect 1454 -3259 1455 -3258
rect 1458 -3259 1459 -3258
rect 163 -3261 164 -3260
rect 233 -3261 234 -3260
rect 478 -3261 479 -3260
rect 485 -3261 486 -3260
rect 681 -3261 682 -3260
rect 723 -3261 724 -3260
rect 163 -3263 164 -3262
rect 208 -3263 209 -3262
rect 408 -3263 409 -3262
rect 485 -3263 486 -3262
rect 709 -3263 710 -3262
rect 835 -3263 836 -3262
rect 208 -3265 209 -3264
rect 240 -3265 241 -3264
rect 240 -3267 241 -3266
rect 492 -3267 493 -3266
rect 163 -3278 164 -3277
rect 229 -3278 230 -3277
rect 243 -3278 244 -3277
rect 534 -3278 535 -3277
rect 593 -3278 594 -3277
rect 646 -3278 647 -3277
rect 670 -3278 671 -3277
rect 674 -3278 675 -3277
rect 684 -3278 685 -3277
rect 702 -3278 703 -3277
rect 723 -3278 724 -3277
rect 919 -3278 920 -3277
rect 936 -3278 937 -3277
rect 940 -3278 941 -3277
rect 947 -3278 948 -3277
rect 975 -3278 976 -3277
rect 982 -3278 983 -3277
rect 989 -3278 990 -3277
rect 1003 -3278 1004 -3277
rect 1059 -3278 1060 -3277
rect 1073 -3278 1074 -3277
rect 1076 -3278 1077 -3277
rect 1108 -3278 1109 -3277
rect 1115 -3278 1116 -3277
rect 1122 -3278 1123 -3277
rect 1129 -3278 1130 -3277
rect 1136 -3278 1137 -3277
rect 1157 -3278 1158 -3277
rect 1171 -3278 1172 -3277
rect 1185 -3278 1186 -3277
rect 1206 -3278 1207 -3277
rect 1213 -3278 1214 -3277
rect 1216 -3278 1217 -3277
rect 1220 -3278 1221 -3277
rect 1251 -3278 1252 -3277
rect 1290 -3278 1291 -3277
rect 1451 -3278 1452 -3277
rect 1461 -3278 1462 -3277
rect 177 -3280 178 -3279
rect 205 -3280 206 -3279
rect 208 -3280 209 -3279
rect 240 -3280 241 -3279
rect 289 -3280 290 -3279
rect 411 -3280 412 -3279
rect 415 -3280 416 -3279
rect 646 -3280 647 -3279
rect 688 -3280 689 -3279
rect 702 -3280 703 -3279
rect 730 -3280 731 -3279
rect 751 -3280 752 -3279
rect 779 -3280 780 -3279
rect 800 -3280 801 -3279
rect 807 -3280 808 -3279
rect 835 -3280 836 -3279
rect 838 -3280 839 -3279
rect 996 -3280 997 -3279
rect 1073 -3280 1074 -3279
rect 1080 -3280 1081 -3279
rect 1097 -3280 1098 -3279
rect 1290 -3280 1291 -3279
rect 1458 -3280 1459 -3279
rect 1465 -3280 1466 -3279
rect 177 -3282 178 -3281
rect 268 -3282 269 -3281
rect 282 -3282 283 -3281
rect 289 -3282 290 -3281
rect 331 -3282 332 -3281
rect 383 -3282 384 -3281
rect 394 -3282 395 -3281
rect 618 -3282 619 -3281
rect 639 -3282 640 -3281
rect 674 -3282 675 -3281
rect 681 -3282 682 -3281
rect 688 -3282 689 -3281
rect 751 -3282 752 -3281
rect 758 -3282 759 -3281
rect 779 -3282 780 -3281
rect 786 -3282 787 -3281
rect 793 -3282 794 -3281
rect 800 -3282 801 -3281
rect 814 -3282 815 -3281
rect 849 -3282 850 -3281
rect 856 -3282 857 -3281
rect 877 -3282 878 -3281
rect 912 -3282 913 -3281
rect 919 -3282 920 -3281
rect 940 -3282 941 -3281
rect 954 -3282 955 -3281
rect 1076 -3282 1077 -3281
rect 1080 -3282 1081 -3281
rect 1101 -3282 1102 -3281
rect 1108 -3282 1109 -3281
rect 1125 -3282 1126 -3281
rect 1164 -3282 1165 -3281
rect 184 -3284 185 -3283
rect 191 -3284 192 -3283
rect 226 -3284 227 -3283
rect 247 -3284 248 -3283
rect 282 -3284 283 -3283
rect 296 -3284 297 -3283
rect 324 -3284 325 -3283
rect 394 -3284 395 -3283
rect 415 -3284 416 -3283
rect 429 -3284 430 -3283
rect 457 -3284 458 -3283
rect 590 -3284 591 -3283
rect 593 -3284 594 -3283
rect 709 -3284 710 -3283
rect 712 -3284 713 -3283
rect 814 -3284 815 -3283
rect 863 -3284 864 -3283
rect 884 -3284 885 -3283
rect 912 -3284 913 -3283
rect 933 -3284 934 -3283
rect 954 -3284 955 -3283
rect 961 -3284 962 -3283
rect 1136 -3284 1137 -3283
rect 1150 -3284 1151 -3283
rect 156 -3286 157 -3285
rect 191 -3286 192 -3285
rect 226 -3286 227 -3285
rect 618 -3286 619 -3285
rect 639 -3286 640 -3285
rect 660 -3286 661 -3285
rect 681 -3286 682 -3285
rect 807 -3286 808 -3285
rect 870 -3286 871 -3285
rect 884 -3286 885 -3285
rect 926 -3286 927 -3285
rect 961 -3286 962 -3285
rect 184 -3288 185 -3287
rect 198 -3288 199 -3287
rect 296 -3288 297 -3287
rect 572 -3288 573 -3287
rect 576 -3288 577 -3287
rect 933 -3288 934 -3287
rect 187 -3290 188 -3289
rect 268 -3290 269 -3289
rect 331 -3290 332 -3289
rect 345 -3290 346 -3289
rect 366 -3290 367 -3289
rect 590 -3290 591 -3289
rect 597 -3290 598 -3289
rect 723 -3290 724 -3289
rect 744 -3290 745 -3289
rect 786 -3290 787 -3289
rect 793 -3290 794 -3289
rect 821 -3290 822 -3289
rect 877 -3290 878 -3289
rect 898 -3290 899 -3289
rect 198 -3292 199 -3291
rect 219 -3292 220 -3291
rect 338 -3292 339 -3291
rect 345 -3292 346 -3291
rect 366 -3292 367 -3291
rect 387 -3292 388 -3291
rect 422 -3292 423 -3291
rect 457 -3292 458 -3291
rect 471 -3292 472 -3291
rect 478 -3292 479 -3291
rect 488 -3292 489 -3291
rect 583 -3292 584 -3291
rect 635 -3292 636 -3291
rect 870 -3292 871 -3291
rect 891 -3292 892 -3291
rect 926 -3292 927 -3291
rect 170 -3294 171 -3293
rect 338 -3294 339 -3293
rect 373 -3294 374 -3293
rect 429 -3294 430 -3293
rect 446 -3294 447 -3293
rect 744 -3294 745 -3293
rect 758 -3294 759 -3293
rect 765 -3294 766 -3293
rect 821 -3294 822 -3293
rect 842 -3294 843 -3293
rect 898 -3294 899 -3293
rect 905 -3294 906 -3293
rect 219 -3296 220 -3295
rect 233 -3296 234 -3295
rect 275 -3296 276 -3295
rect 387 -3296 388 -3295
rect 422 -3296 423 -3295
rect 506 -3296 507 -3295
rect 534 -3296 535 -3295
rect 541 -3296 542 -3295
rect 555 -3296 556 -3295
rect 597 -3296 598 -3295
rect 660 -3296 661 -3295
rect 716 -3296 717 -3295
rect 765 -3296 766 -3295
rect 772 -3296 773 -3295
rect 842 -3296 843 -3295
rect 845 -3296 846 -3295
rect 880 -3296 881 -3295
rect 905 -3296 906 -3295
rect 233 -3298 234 -3297
rect 408 -3298 409 -3297
rect 464 -3298 465 -3297
rect 555 -3298 556 -3297
rect 576 -3298 577 -3297
rect 709 -3298 710 -3297
rect 716 -3298 717 -3297
rect 737 -3298 738 -3297
rect 254 -3300 255 -3299
rect 275 -3300 276 -3299
rect 317 -3300 318 -3299
rect 373 -3300 374 -3299
rect 464 -3300 465 -3299
rect 604 -3300 605 -3299
rect 695 -3300 696 -3299
rect 772 -3300 773 -3299
rect 254 -3302 255 -3301
rect 352 -3302 353 -3301
rect 401 -3302 402 -3301
rect 695 -3302 696 -3301
rect 737 -3302 738 -3301
rect 891 -3302 892 -3301
rect 310 -3304 311 -3303
rect 317 -3304 318 -3303
rect 352 -3304 353 -3303
rect 485 -3304 486 -3303
rect 492 -3304 493 -3303
rect 541 -3304 542 -3303
rect 583 -3304 584 -3303
rect 632 -3304 633 -3303
rect 303 -3306 304 -3305
rect 310 -3306 311 -3305
rect 380 -3306 381 -3305
rect 485 -3306 486 -3305
rect 604 -3306 605 -3305
rect 782 -3306 783 -3305
rect 303 -3308 304 -3307
rect 992 -3308 993 -3307
rect 380 -3310 381 -3309
rect 730 -3310 731 -3309
rect 401 -3312 402 -3311
rect 450 -3312 451 -3311
rect 467 -3312 468 -3311
rect 632 -3312 633 -3311
rect 436 -3314 437 -3313
rect 492 -3314 493 -3313
rect 436 -3316 437 -3315
rect 443 -3316 444 -3315
rect 450 -3316 451 -3315
rect 625 -3316 626 -3315
rect 324 -3318 325 -3317
rect 443 -3318 444 -3317
rect 474 -3318 475 -3317
rect 513 -3318 514 -3317
rect 625 -3318 626 -3317
rect 653 -3318 654 -3317
rect 478 -3320 479 -3319
rect 499 -3320 500 -3319
rect 513 -3320 514 -3319
rect 667 -3320 668 -3319
rect 499 -3322 500 -3321
rect 520 -3322 521 -3321
rect 548 -3322 549 -3321
rect 653 -3322 654 -3321
rect 506 -3324 507 -3323
rect 667 -3324 668 -3323
rect 520 -3326 521 -3325
rect 527 -3326 528 -3325
rect 548 -3326 549 -3325
rect 562 -3326 563 -3325
rect 408 -3328 409 -3327
rect 562 -3328 563 -3327
rect 527 -3330 528 -3329
rect 569 -3330 570 -3329
rect 191 -3341 192 -3340
rect 194 -3341 195 -3340
rect 261 -3341 262 -3340
rect 618 -3341 619 -3340
rect 621 -3341 622 -3340
rect 786 -3341 787 -3340
rect 807 -3341 808 -3340
rect 866 -3341 867 -3340
rect 870 -3341 871 -3340
rect 1097 -3341 1098 -3340
rect 1115 -3341 1116 -3340
rect 1122 -3341 1123 -3340
rect 1139 -3341 1140 -3340
rect 1143 -3341 1144 -3340
rect 1353 -3341 1354 -3340
rect 1367 -3341 1368 -3340
rect 191 -3343 192 -3342
rect 233 -3343 234 -3342
rect 240 -3343 241 -3342
rect 261 -3343 262 -3342
rect 264 -3343 265 -3342
rect 275 -3343 276 -3342
rect 282 -3343 283 -3342
rect 411 -3343 412 -3342
rect 471 -3343 472 -3342
rect 569 -3343 570 -3342
rect 576 -3343 577 -3342
rect 590 -3343 591 -3342
rect 604 -3343 605 -3342
rect 618 -3343 619 -3342
rect 709 -3343 710 -3342
rect 740 -3343 741 -3342
rect 821 -3343 822 -3342
rect 835 -3343 836 -3342
rect 842 -3343 843 -3342
rect 884 -3343 885 -3342
rect 894 -3343 895 -3342
rect 926 -3343 927 -3342
rect 947 -3343 948 -3342
rect 961 -3343 962 -3342
rect 975 -3343 976 -3342
rect 996 -3343 997 -3342
rect 1059 -3343 1060 -3342
rect 1073 -3343 1074 -3342
rect 1108 -3343 1109 -3342
rect 1115 -3343 1116 -3342
rect 1290 -3343 1291 -3342
rect 1367 -3343 1368 -3342
rect 198 -3345 199 -3344
rect 240 -3345 241 -3344
rect 254 -3345 255 -3344
rect 275 -3345 276 -3344
rect 282 -3345 283 -3344
rect 289 -3345 290 -3344
rect 303 -3345 304 -3344
rect 306 -3345 307 -3344
rect 338 -3345 339 -3344
rect 464 -3345 465 -3344
rect 471 -3345 472 -3344
rect 520 -3345 521 -3344
rect 541 -3345 542 -3344
rect 933 -3345 934 -3344
rect 1062 -3345 1063 -3344
rect 1066 -3345 1067 -3344
rect 1073 -3345 1074 -3344
rect 1080 -3345 1081 -3344
rect 198 -3347 199 -3346
rect 352 -3347 353 -3346
rect 355 -3347 356 -3346
rect 506 -3347 507 -3346
rect 520 -3347 521 -3346
rect 527 -3347 528 -3346
rect 558 -3347 559 -3346
rect 569 -3347 570 -3346
rect 604 -3347 605 -3346
rect 646 -3347 647 -3346
rect 660 -3347 661 -3346
rect 709 -3347 710 -3346
rect 712 -3347 713 -3346
rect 793 -3347 794 -3346
rect 828 -3347 829 -3346
rect 831 -3347 832 -3346
rect 870 -3347 871 -3346
rect 905 -3347 906 -3346
rect 926 -3347 927 -3346
rect 954 -3347 955 -3346
rect 226 -3349 227 -3348
rect 646 -3349 647 -3348
rect 737 -3349 738 -3348
rect 800 -3349 801 -3348
rect 884 -3349 885 -3348
rect 891 -3349 892 -3348
rect 905 -3349 906 -3348
rect 912 -3349 913 -3348
rect 247 -3351 248 -3350
rect 254 -3351 255 -3350
rect 268 -3351 269 -3350
rect 443 -3351 444 -3350
rect 492 -3351 493 -3350
rect 544 -3351 545 -3350
rect 555 -3351 556 -3350
rect 660 -3351 661 -3350
rect 737 -3351 738 -3350
rect 758 -3351 759 -3350
rect 775 -3351 776 -3350
rect 821 -3351 822 -3350
rect 877 -3351 878 -3350
rect 912 -3351 913 -3350
rect 212 -3353 213 -3352
rect 268 -3353 269 -3352
rect 289 -3353 290 -3352
rect 317 -3353 318 -3352
rect 366 -3353 367 -3352
rect 380 -3353 381 -3352
rect 383 -3353 384 -3352
rect 387 -3353 388 -3352
rect 394 -3353 395 -3352
rect 467 -3353 468 -3352
rect 495 -3353 496 -3352
rect 527 -3353 528 -3352
rect 744 -3353 745 -3352
rect 828 -3353 829 -3352
rect 863 -3353 864 -3352
rect 877 -3353 878 -3352
rect 177 -3355 178 -3354
rect 394 -3355 395 -3354
rect 397 -3355 398 -3354
rect 681 -3355 682 -3354
rect 744 -3355 745 -3354
rect 772 -3355 773 -3354
rect 863 -3355 864 -3354
rect 898 -3355 899 -3354
rect 177 -3357 178 -3356
rect 229 -3357 230 -3356
rect 296 -3357 297 -3356
rect 366 -3357 367 -3356
rect 373 -3357 374 -3356
rect 387 -3357 388 -3356
rect 443 -3357 444 -3356
rect 572 -3357 573 -3356
rect 576 -3357 577 -3356
rect 681 -3357 682 -3356
rect 758 -3357 759 -3356
rect 765 -3357 766 -3356
rect 205 -3359 206 -3358
rect 212 -3359 213 -3358
rect 219 -3359 220 -3358
rect 247 -3359 248 -3358
rect 296 -3359 297 -3358
rect 359 -3359 360 -3358
rect 373 -3359 374 -3358
rect 457 -3359 458 -3358
rect 499 -3359 500 -3358
rect 593 -3359 594 -3358
rect 751 -3359 752 -3358
rect 765 -3359 766 -3358
rect 205 -3361 206 -3360
rect 324 -3361 325 -3360
rect 359 -3361 360 -3360
rect 488 -3361 489 -3360
rect 499 -3361 500 -3360
rect 562 -3361 563 -3360
rect 730 -3361 731 -3360
rect 751 -3361 752 -3360
rect 219 -3363 220 -3362
rect 331 -3363 332 -3362
rect 415 -3363 416 -3362
rect 457 -3363 458 -3362
rect 716 -3363 717 -3362
rect 730 -3363 731 -3362
rect 303 -3365 304 -3364
rect 310 -3365 311 -3364
rect 317 -3365 318 -3364
rect 408 -3365 409 -3364
rect 450 -3365 451 -3364
rect 562 -3365 563 -3364
rect 639 -3365 640 -3364
rect 716 -3365 717 -3364
rect 310 -3367 311 -3366
rect 422 -3367 423 -3366
rect 450 -3367 451 -3366
rect 478 -3367 479 -3366
rect 639 -3367 640 -3366
rect 674 -3367 675 -3366
rect 306 -3369 307 -3368
rect 422 -3369 423 -3368
rect 478 -3369 479 -3368
rect 534 -3369 535 -3368
rect 667 -3369 668 -3368
rect 674 -3369 675 -3368
rect 324 -3371 325 -3370
rect 345 -3371 346 -3370
rect 352 -3371 353 -3370
rect 415 -3371 416 -3370
rect 625 -3371 626 -3370
rect 667 -3371 668 -3370
rect 331 -3373 332 -3372
rect 436 -3373 437 -3372
rect 611 -3373 612 -3372
rect 625 -3373 626 -3372
rect 345 -3375 346 -3374
rect 537 -3375 538 -3374
rect 611 -3375 612 -3374
rect 723 -3375 724 -3374
rect 401 -3377 402 -3376
rect 436 -3377 437 -3376
rect 723 -3377 724 -3376
rect 845 -3377 846 -3376
rect 401 -3379 402 -3378
rect 534 -3379 535 -3378
rect 814 -3379 815 -3378
rect 845 -3379 846 -3378
rect 408 -3381 409 -3380
rect 485 -3381 486 -3380
rect 814 -3381 815 -3380
rect 936 -3381 937 -3380
rect 485 -3383 486 -3382
rect 653 -3383 654 -3382
rect 653 -3385 654 -3384
rect 688 -3385 689 -3384
rect 583 -3387 584 -3386
rect 688 -3387 689 -3386
rect 583 -3389 584 -3388
rect 632 -3389 633 -3388
rect 548 -3391 549 -3390
rect 632 -3391 633 -3390
rect 548 -3393 549 -3392
rect 597 -3393 598 -3392
rect 446 -3395 447 -3394
rect 597 -3395 598 -3394
rect 177 -3406 178 -3405
rect 226 -3406 227 -3405
rect 247 -3406 248 -3405
rect 355 -3406 356 -3405
rect 366 -3406 367 -3405
rect 383 -3406 384 -3405
rect 457 -3406 458 -3405
rect 495 -3406 496 -3405
rect 499 -3406 500 -3405
rect 506 -3406 507 -3405
rect 513 -3406 514 -3405
rect 576 -3406 577 -3405
rect 632 -3406 633 -3405
rect 635 -3406 636 -3405
rect 695 -3406 696 -3405
rect 702 -3406 703 -3405
rect 719 -3406 720 -3405
rect 737 -3406 738 -3405
rect 765 -3406 766 -3405
rect 772 -3406 773 -3405
rect 782 -3406 783 -3405
rect 982 -3406 983 -3405
rect 1367 -3406 1368 -3405
rect 1395 -3406 1396 -3405
rect 184 -3408 185 -3407
rect 229 -3408 230 -3407
rect 264 -3408 265 -3407
rect 268 -3408 269 -3407
rect 275 -3408 276 -3407
rect 394 -3408 395 -3407
rect 467 -3408 468 -3407
rect 604 -3408 605 -3407
rect 632 -3408 633 -3407
rect 653 -3408 654 -3407
rect 681 -3408 682 -3407
rect 765 -3408 766 -3407
rect 772 -3408 773 -3407
rect 779 -3408 780 -3407
rect 831 -3408 832 -3407
rect 856 -3408 857 -3407
rect 891 -3408 892 -3407
rect 926 -3408 927 -3407
rect 947 -3408 948 -3407
rect 964 -3408 965 -3407
rect 968 -3408 969 -3407
rect 975 -3408 976 -3407
rect 212 -3410 213 -3409
rect 222 -3410 223 -3409
rect 233 -3410 234 -3409
rect 275 -3410 276 -3409
rect 310 -3410 311 -3409
rect 394 -3410 395 -3409
rect 471 -3410 472 -3409
rect 485 -3410 486 -3409
rect 499 -3410 500 -3409
rect 555 -3410 556 -3409
rect 558 -3410 559 -3409
rect 625 -3410 626 -3409
rect 653 -3410 654 -3409
rect 667 -3410 668 -3409
rect 688 -3410 689 -3409
rect 779 -3410 780 -3409
rect 842 -3410 843 -3409
rect 870 -3410 871 -3409
rect 912 -3410 913 -3409
rect 926 -3410 927 -3409
rect 954 -3410 955 -3409
rect 1010 -3410 1011 -3409
rect 254 -3412 255 -3411
rect 310 -3412 311 -3411
rect 317 -3412 318 -3411
rect 338 -3412 339 -3411
rect 341 -3412 342 -3411
rect 387 -3412 388 -3411
rect 408 -3412 409 -3411
rect 471 -3412 472 -3411
rect 478 -3412 479 -3411
rect 492 -3412 493 -3411
rect 520 -3412 521 -3411
rect 541 -3412 542 -3411
rect 569 -3412 570 -3411
rect 576 -3412 577 -3411
rect 625 -3412 626 -3411
rect 639 -3412 640 -3411
rect 660 -3412 661 -3411
rect 681 -3412 682 -3411
rect 688 -3412 689 -3411
rect 723 -3412 724 -3411
rect 730 -3412 731 -3411
rect 733 -3412 734 -3411
rect 842 -3412 843 -3411
rect 845 -3412 846 -3411
rect 856 -3412 857 -3411
rect 884 -3412 885 -3411
rect 905 -3412 906 -3411
rect 912 -3412 913 -3411
rect 961 -3412 962 -3411
rect 1094 -3412 1095 -3411
rect 191 -3414 192 -3413
rect 341 -3414 342 -3413
rect 352 -3414 353 -3413
rect 401 -3414 402 -3413
rect 534 -3414 535 -3413
rect 548 -3414 549 -3413
rect 569 -3414 570 -3413
rect 590 -3414 591 -3413
rect 597 -3414 598 -3413
rect 660 -3414 661 -3413
rect 695 -3414 696 -3413
rect 716 -3414 717 -3413
rect 723 -3414 724 -3413
rect 814 -3414 815 -3413
rect 863 -3414 864 -3413
rect 870 -3414 871 -3413
rect 877 -3414 878 -3413
rect 884 -3414 885 -3413
rect 240 -3416 241 -3415
rect 254 -3416 255 -3415
rect 261 -3416 262 -3415
rect 268 -3416 269 -3415
rect 289 -3416 290 -3415
rect 317 -3416 318 -3415
rect 327 -3416 328 -3415
rect 415 -3416 416 -3415
rect 488 -3416 489 -3415
rect 534 -3416 535 -3415
rect 541 -3416 542 -3415
rect 642 -3416 643 -3415
rect 730 -3416 731 -3415
rect 758 -3416 759 -3415
rect 821 -3416 822 -3415
rect 863 -3416 864 -3415
rect 198 -3418 199 -3417
rect 240 -3418 241 -3417
rect 331 -3418 332 -3417
rect 401 -3418 402 -3417
rect 527 -3418 528 -3417
rect 548 -3418 549 -3417
rect 562 -3418 563 -3417
rect 597 -3418 598 -3417
rect 639 -3418 640 -3417
rect 775 -3418 776 -3417
rect 821 -3418 822 -3417
rect 835 -3418 836 -3417
rect 359 -3420 360 -3419
rect 387 -3420 388 -3419
rect 562 -3420 563 -3419
rect 583 -3420 584 -3419
rect 646 -3420 647 -3419
rect 835 -3420 836 -3419
rect 296 -3422 297 -3421
rect 359 -3422 360 -3421
rect 373 -3422 374 -3421
rect 408 -3422 409 -3421
rect 583 -3422 584 -3421
rect 611 -3422 612 -3421
rect 618 -3422 619 -3421
rect 646 -3422 647 -3421
rect 733 -3422 734 -3421
rect 758 -3422 759 -3421
rect 219 -3424 220 -3423
rect 296 -3424 297 -3423
rect 303 -3424 304 -3423
rect 373 -3424 374 -3423
rect 303 -3426 304 -3425
rect 429 -3426 430 -3425
rect 429 -3428 430 -3427
rect 436 -3428 437 -3427
rect 436 -3430 437 -3429
rect 450 -3430 451 -3429
rect 422 -3432 423 -3431
rect 450 -3432 451 -3431
rect 345 -3434 346 -3433
rect 422 -3434 423 -3433
rect 324 -3436 325 -3435
rect 345 -3436 346 -3435
rect 205 -3438 206 -3437
rect 324 -3438 325 -3437
rect 222 -3449 223 -3448
rect 327 -3449 328 -3448
rect 338 -3449 339 -3448
rect 352 -3449 353 -3448
rect 359 -3449 360 -3448
rect 380 -3449 381 -3448
rect 401 -3449 402 -3448
rect 464 -3449 465 -3448
rect 478 -3449 479 -3448
rect 485 -3449 486 -3448
rect 506 -3449 507 -3448
rect 541 -3449 542 -3448
rect 597 -3449 598 -3448
rect 604 -3449 605 -3448
rect 614 -3449 615 -3448
rect 625 -3449 626 -3448
rect 642 -3449 643 -3448
rect 688 -3449 689 -3448
rect 698 -3449 699 -3448
rect 702 -3449 703 -3448
rect 709 -3449 710 -3448
rect 737 -3449 738 -3448
rect 740 -3449 741 -3448
rect 758 -3449 759 -3448
rect 765 -3449 766 -3448
rect 779 -3449 780 -3448
rect 782 -3449 783 -3448
rect 964 -3449 965 -3448
rect 982 -3449 983 -3448
rect 1066 -3449 1067 -3448
rect 1073 -3449 1074 -3448
rect 1076 -3449 1077 -3448
rect 1094 -3449 1095 -3448
rect 1220 -3449 1221 -3448
rect 1223 -3449 1224 -3448
rect 1227 -3449 1228 -3448
rect 1409 -3449 1410 -3448
rect 1416 -3449 1417 -3448
rect 254 -3451 255 -3450
rect 261 -3451 262 -3450
rect 264 -3451 265 -3450
rect 460 -3451 461 -3450
rect 471 -3451 472 -3450
rect 485 -3451 486 -3450
rect 520 -3451 521 -3450
rect 572 -3451 573 -3450
rect 621 -3451 622 -3450
rect 723 -3451 724 -3450
rect 737 -3451 738 -3450
rect 751 -3451 752 -3450
rect 821 -3451 822 -3450
rect 828 -3451 829 -3450
rect 831 -3451 832 -3450
rect 849 -3451 850 -3450
rect 933 -3451 934 -3450
rect 954 -3451 955 -3450
rect 957 -3451 958 -3450
rect 968 -3451 969 -3450
rect 1010 -3451 1011 -3450
rect 1073 -3451 1074 -3450
rect 1395 -3451 1396 -3450
rect 1409 -3451 1410 -3450
rect 240 -3453 241 -3452
rect 254 -3453 255 -3452
rect 268 -3453 269 -3452
rect 289 -3453 290 -3452
rect 292 -3453 293 -3452
rect 359 -3453 360 -3452
rect 373 -3453 374 -3452
rect 401 -3453 402 -3452
rect 408 -3453 409 -3452
rect 415 -3453 416 -3452
rect 422 -3453 423 -3452
rect 502 -3453 503 -3452
rect 541 -3453 542 -3452
rect 569 -3453 570 -3452
rect 625 -3453 626 -3452
rect 632 -3453 633 -3452
rect 674 -3453 675 -3452
rect 691 -3453 692 -3452
rect 695 -3453 696 -3452
rect 709 -3453 710 -3452
rect 719 -3453 720 -3452
rect 730 -3453 731 -3452
rect 824 -3453 825 -3452
rect 961 -3453 962 -3452
rect 275 -3455 276 -3454
rect 306 -3455 307 -3454
rect 317 -3455 318 -3454
rect 327 -3455 328 -3454
rect 345 -3455 346 -3454
rect 352 -3455 353 -3454
rect 394 -3455 395 -3454
rect 471 -3455 472 -3454
rect 569 -3455 570 -3454
rect 583 -3455 584 -3454
rect 667 -3455 668 -3454
rect 674 -3455 675 -3454
rect 681 -3455 682 -3454
rect 716 -3455 717 -3454
rect 835 -3455 836 -3454
rect 891 -3455 892 -3454
rect 947 -3455 948 -3454
rect 975 -3455 976 -3454
rect 282 -3457 283 -3456
rect 303 -3457 304 -3456
rect 310 -3457 311 -3456
rect 317 -3457 318 -3456
rect 387 -3457 388 -3456
rect 394 -3457 395 -3456
rect 422 -3457 423 -3456
rect 429 -3457 430 -3456
rect 450 -3457 451 -3456
rect 457 -3457 458 -3456
rect 576 -3457 577 -3456
rect 583 -3457 584 -3456
rect 660 -3457 661 -3456
rect 681 -3457 682 -3456
rect 688 -3457 689 -3456
rect 744 -3457 745 -3456
rect 821 -3457 822 -3456
rect 835 -3457 836 -3456
rect 849 -3457 850 -3456
rect 870 -3457 871 -3456
rect 296 -3459 297 -3458
rect 331 -3459 332 -3458
rect 425 -3459 426 -3458
rect 639 -3459 640 -3458
rect 660 -3459 661 -3458
rect 726 -3459 727 -3458
rect 863 -3459 864 -3458
rect 870 -3459 871 -3458
rect 429 -3461 430 -3460
rect 436 -3461 437 -3460
rect 555 -3461 556 -3460
rect 576 -3461 577 -3460
rect 695 -3461 696 -3460
rect 758 -3461 759 -3460
rect 555 -3463 556 -3462
rect 562 -3463 563 -3462
rect 534 -3465 535 -3464
rect 562 -3465 563 -3464
rect 261 -3476 262 -3475
rect 268 -3476 269 -3475
rect 303 -3476 304 -3475
rect 310 -3476 311 -3475
rect 317 -3476 318 -3475
rect 327 -3476 328 -3475
rect 380 -3476 381 -3475
rect 411 -3476 412 -3475
rect 415 -3476 416 -3475
rect 436 -3476 437 -3475
rect 467 -3476 468 -3475
rect 520 -3476 521 -3475
rect 548 -3476 549 -3475
rect 551 -3476 552 -3475
rect 583 -3476 584 -3475
rect 590 -3476 591 -3475
rect 597 -3476 598 -3475
rect 660 -3476 661 -3475
rect 681 -3476 682 -3475
rect 688 -3476 689 -3475
rect 695 -3476 696 -3475
rect 828 -3476 829 -3475
rect 842 -3476 843 -3475
rect 849 -3476 850 -3475
rect 852 -3476 853 -3475
rect 856 -3476 857 -3475
rect 870 -3476 871 -3475
rect 887 -3476 888 -3475
rect 891 -3476 892 -3475
rect 950 -3476 951 -3475
rect 989 -3476 990 -3475
rect 992 -3476 993 -3475
rect 1066 -3476 1067 -3475
rect 1094 -3476 1095 -3475
rect 1115 -3476 1116 -3475
rect 1118 -3476 1119 -3475
rect 1213 -3476 1214 -3475
rect 1220 -3476 1221 -3475
rect 1409 -3476 1410 -3475
rect 1412 -3476 1413 -3475
rect 254 -3478 255 -3477
rect 261 -3478 262 -3477
rect 394 -3478 395 -3477
rect 408 -3478 409 -3477
rect 418 -3478 419 -3477
rect 698 -3478 699 -3477
rect 709 -3478 710 -3477
rect 716 -3478 717 -3477
rect 726 -3478 727 -3477
rect 737 -3478 738 -3477
rect 758 -3478 759 -3477
rect 821 -3478 822 -3477
rect 877 -3478 878 -3477
rect 898 -3478 899 -3477
rect 905 -3478 906 -3477
rect 933 -3478 934 -3477
rect 1115 -3478 1116 -3477
rect 1122 -3478 1123 -3477
rect 1220 -3478 1221 -3477
rect 1227 -3478 1228 -3477
rect 1409 -3478 1410 -3477
rect 1416 -3478 1417 -3477
rect 401 -3480 402 -3479
rect 408 -3480 409 -3479
rect 429 -3480 430 -3479
rect 439 -3480 440 -3479
rect 471 -3480 472 -3479
rect 506 -3480 507 -3479
rect 548 -3480 549 -3479
rect 555 -3480 556 -3479
rect 576 -3480 577 -3479
rect 583 -3480 584 -3479
rect 604 -3480 605 -3479
rect 621 -3480 622 -3479
rect 646 -3480 647 -3479
rect 660 -3480 661 -3479
rect 674 -3480 675 -3479
rect 681 -3480 682 -3479
rect 359 -3482 360 -3481
rect 429 -3482 430 -3481
rect 436 -3482 437 -3481
rect 443 -3482 444 -3481
rect 478 -3482 479 -3481
rect 502 -3482 503 -3481
rect 513 -3482 514 -3481
rect 646 -3482 647 -3481
rect 1412 -3482 1413 -3481
rect 1416 -3482 1417 -3481
rect 478 -3484 479 -3483
rect 614 -3484 615 -3483
rect 485 -3486 486 -3485
rect 516 -3486 517 -3485
rect 562 -3486 563 -3485
rect 576 -3486 577 -3485
rect 611 -3486 612 -3485
rect 625 -3486 626 -3485
rect 492 -3488 493 -3487
rect 499 -3488 500 -3487
rect 261 -3499 262 -3498
rect 271 -3499 272 -3498
rect 310 -3499 311 -3498
rect 324 -3499 325 -3498
rect 331 -3499 332 -3498
rect 345 -3499 346 -3498
rect 352 -3499 353 -3498
rect 359 -3499 360 -3498
rect 408 -3499 409 -3498
rect 418 -3499 419 -3498
rect 429 -3499 430 -3498
rect 436 -3499 437 -3498
rect 541 -3499 542 -3498
rect 551 -3499 552 -3498
rect 555 -3499 556 -3498
rect 565 -3499 566 -3498
rect 583 -3499 584 -3498
rect 597 -3499 598 -3498
rect 646 -3499 647 -3498
rect 653 -3499 654 -3498
rect 660 -3499 661 -3498
rect 667 -3499 668 -3498
rect 681 -3499 682 -3498
rect 691 -3499 692 -3498
rect 716 -3499 717 -3498
rect 723 -3499 724 -3498
rect 828 -3499 829 -3498
rect 870 -3499 871 -3498
rect 898 -3499 899 -3498
rect 905 -3499 906 -3498
rect 922 -3499 923 -3498
rect 926 -3499 927 -3498
rect 940 -3499 941 -3498
rect 950 -3499 951 -3498
rect 989 -3499 990 -3498
rect 996 -3499 997 -3498
rect 1094 -3499 1095 -3498
rect 1115 -3499 1116 -3498
rect 1118 -3499 1119 -3498
rect 1122 -3499 1123 -3498
rect 1360 -3499 1361 -3498
rect 1367 -3499 1368 -3498
rect 1412 -3499 1413 -3498
rect 1416 -3499 1417 -3498
rect 268 -3501 269 -3500
rect 275 -3501 276 -3500
rect 331 -3501 332 -3500
rect 338 -3501 339 -3500
rect 355 -3501 356 -3500
rect 478 -3501 479 -3500
rect 541 -3501 542 -3500
rect 548 -3501 549 -3500
rect 576 -3501 577 -3500
rect 583 -3501 584 -3500
rect 835 -3501 836 -3500
rect 859 -3501 860 -3500
rect 576 -3503 577 -3502
rect 590 -3503 591 -3502
rect 842 -3503 843 -3502
rect 849 -3503 850 -3502
rect 271 -3514 272 -3513
rect 275 -3514 276 -3513
rect 327 -3514 328 -3513
rect 331 -3514 332 -3513
rect 355 -3514 356 -3513
rect 359 -3514 360 -3513
rect 541 -3514 542 -3513
rect 555 -3514 556 -3513
rect 565 -3514 566 -3513
rect 569 -3514 570 -3513
rect 579 -3514 580 -3513
rect 583 -3514 584 -3513
rect 660 -3514 661 -3513
rect 667 -3514 668 -3513
rect 856 -3514 857 -3513
rect 877 -3514 878 -3513
rect 1353 -3514 1354 -3513
rect 1360 -3514 1361 -3513
rect 1363 -3514 1364 -3513
rect 1367 -3514 1368 -3513
rect 870 -3516 871 -3515
rect 915 -3516 916 -3515
<< metal2 >>
rect 282 -5 283 1
rect 345 -5 346 1
rect 425 -5 426 1
rect 450 -5 451 1
rect 464 -5 465 1
rect 478 -5 479 1
rect 905 -5 906 1
rect 950 -5 951 1
rect 317 -5 318 -1
rect 352 -5 353 -1
rect 436 -5 437 -1
rect 513 -5 514 -1
rect 947 -5 948 -1
rect 989 -5 990 -1
rect 443 -5 444 -3
rect 457 -5 458 -3
rect 226 -24 227 -14
rect 285 -15 286 -13
rect 303 -24 304 -14
rect 317 -15 318 -13
rect 338 -24 339 -14
rect 359 -24 360 -14
rect 366 -24 367 -14
rect 436 -15 437 -13
rect 450 -15 451 -13
rect 457 -24 458 -14
rect 478 -15 479 -13
rect 499 -24 500 -14
rect 506 -15 507 -13
rect 611 -24 612 -14
rect 618 -24 619 -14
rect 625 -24 626 -14
rect 891 -24 892 -14
rect 905 -15 906 -13
rect 989 -15 990 -13
rect 1003 -24 1004 -14
rect 345 -17 346 -13
rect 373 -24 374 -16
rect 380 -24 381 -16
rect 425 -17 426 -13
rect 436 -24 437 -16
rect 443 -17 444 -13
rect 450 -24 451 -16
rect 464 -17 465 -13
rect 513 -17 514 -13
rect 548 -24 549 -16
rect 579 -24 580 -16
rect 590 -24 591 -16
rect 597 -24 598 -16
rect 639 -24 640 -16
rect 289 -24 290 -18
rect 345 -24 346 -18
rect 348 -24 349 -18
rect 408 -24 409 -18
rect 422 -24 423 -18
rect 509 -19 510 -13
rect 527 -24 528 -18
rect 541 -24 542 -18
rect 583 -24 584 -18
rect 604 -24 605 -18
rect 352 -21 353 -13
rect 387 -24 388 -20
rect 394 -24 395 -20
rect 418 -24 419 -20
rect 460 -21 461 -13
rect 464 -24 465 -20
rect 509 -24 510 -20
rect 513 -24 514 -20
rect 537 -24 538 -20
rect 674 -24 675 -20
rect 352 -24 353 -22
rect 362 -24 363 -22
rect 219 -47 220 -33
rect 226 -34 227 -32
rect 275 -47 276 -33
rect 289 -34 290 -32
rect 303 -34 304 -32
rect 303 -47 304 -33
rect 303 -34 304 -32
rect 303 -47 304 -33
rect 324 -47 325 -33
rect 366 -34 367 -32
rect 373 -34 374 -32
rect 373 -47 374 -33
rect 373 -34 374 -32
rect 373 -47 374 -33
rect 387 -34 388 -32
rect 401 -47 402 -33
rect 415 -47 416 -33
rect 436 -34 437 -32
rect 443 -47 444 -33
rect 457 -34 458 -32
rect 464 -34 465 -32
rect 471 -47 472 -33
rect 492 -47 493 -33
rect 565 -47 566 -33
rect 576 -47 577 -33
rect 597 -34 598 -32
rect 604 -34 605 -32
rect 604 -47 605 -33
rect 604 -34 605 -32
rect 604 -47 605 -33
rect 611 -34 612 -32
rect 653 -47 654 -33
rect 674 -34 675 -32
rect 723 -47 724 -33
rect 758 -47 759 -33
rect 828 -47 829 -33
rect 884 -47 885 -33
rect 891 -34 892 -32
rect 1003 -34 1004 -32
rect 1010 -47 1011 -33
rect 282 -47 283 -35
rect 296 -47 297 -35
rect 331 -47 332 -35
rect 341 -47 342 -35
rect 352 -36 353 -32
rect 352 -47 353 -35
rect 352 -36 353 -32
rect 352 -47 353 -35
rect 359 -47 360 -35
rect 432 -47 433 -35
rect 436 -47 437 -35
rect 457 -47 458 -35
rect 499 -36 500 -32
rect 502 -40 503 -35
rect 513 -36 514 -32
rect 520 -36 521 -32
rect 541 -36 542 -32
rect 555 -47 556 -35
rect 583 -47 584 -35
rect 621 -47 622 -35
rect 625 -36 626 -32
rect 632 -47 633 -35
rect 639 -36 640 -32
rect 674 -47 675 -35
rect 338 -38 339 -32
rect 345 -47 346 -37
rect 366 -47 367 -37
rect 380 -38 381 -32
rect 387 -47 388 -37
rect 485 -47 486 -37
rect 499 -47 500 -37
rect 506 -38 507 -32
rect 520 -47 521 -37
rect 527 -38 528 -32
rect 551 -47 552 -37
rect 730 -47 731 -37
rect 338 -47 339 -39
rect 422 -40 423 -32
rect 450 -40 451 -32
rect 464 -47 465 -39
rect 506 -47 507 -39
rect 523 -40 524 -32
rect 541 -47 542 -39
rect 590 -40 591 -32
rect 597 -47 598 -39
rect 625 -47 626 -39
rect 681 -47 682 -39
rect 380 -47 381 -41
rect 394 -42 395 -32
rect 408 -42 409 -32
rect 450 -47 451 -41
rect 548 -42 549 -32
rect 590 -47 591 -41
rect 635 -42 636 -32
rect 639 -47 640 -41
rect 394 -47 395 -43
rect 537 -44 538 -32
rect 408 -47 409 -45
rect 418 -46 419 -32
rect 422 -47 423 -45
rect 429 -47 430 -45
rect 191 -98 192 -56
rect 254 -98 255 -56
rect 278 -98 279 -56
rect 282 -57 283 -55
rect 289 -98 290 -56
rect 464 -57 465 -55
rect 506 -57 507 -55
rect 516 -98 517 -56
rect 523 -98 524 -56
rect 737 -98 738 -56
rect 789 -98 790 -56
rect 863 -98 864 -56
rect 884 -57 885 -55
rect 891 -98 892 -56
rect 1010 -57 1011 -55
rect 1017 -98 1018 -56
rect 205 -98 206 -58
rect 240 -98 241 -58
rect 243 -98 244 -58
rect 261 -98 262 -58
rect 275 -59 276 -55
rect 282 -98 283 -58
rect 296 -98 297 -58
rect 303 -59 304 -55
rect 317 -98 318 -58
rect 390 -59 391 -55
rect 401 -59 402 -55
rect 401 -98 402 -58
rect 401 -59 402 -55
rect 401 -98 402 -58
rect 408 -59 409 -55
rect 408 -98 409 -58
rect 408 -59 409 -55
rect 408 -98 409 -58
rect 464 -98 465 -58
rect 499 -59 500 -55
rect 513 -98 514 -58
rect 520 -59 521 -55
rect 527 -98 528 -58
rect 586 -98 587 -58
rect 597 -59 598 -55
rect 660 -98 661 -58
rect 709 -98 710 -58
rect 758 -59 759 -55
rect 793 -98 794 -58
rect 800 -98 801 -58
rect 828 -59 829 -55
rect 898 -98 899 -58
rect 219 -61 220 -55
rect 247 -98 248 -60
rect 275 -98 276 -60
rect 310 -98 311 -60
rect 341 -61 342 -55
rect 345 -61 346 -55
rect 390 -98 391 -60
rect 478 -98 479 -60
rect 562 -61 563 -55
rect 779 -98 780 -60
rect 233 -98 234 -62
rect 320 -63 321 -55
rect 345 -98 346 -62
rect 380 -63 381 -55
rect 471 -63 472 -55
rect 499 -98 500 -62
rect 569 -63 570 -55
rect 625 -63 626 -55
rect 632 -63 633 -55
rect 646 -98 647 -62
rect 653 -63 654 -55
rect 702 -98 703 -62
rect 730 -63 731 -55
rect 807 -98 808 -62
rect 299 -65 300 -55
rect 338 -65 339 -55
rect 373 -65 374 -55
rect 380 -98 381 -64
rect 471 -98 472 -64
rect 509 -98 510 -64
rect 569 -98 570 -64
rect 583 -65 584 -55
rect 590 -65 591 -55
rect 597 -98 598 -64
rect 604 -65 605 -55
rect 632 -98 633 -64
rect 639 -65 640 -55
rect 653 -98 654 -64
rect 723 -65 724 -55
rect 730 -98 731 -64
rect 219 -98 220 -66
rect 299 -98 300 -66
rect 303 -98 304 -66
rect 324 -67 325 -55
rect 338 -98 339 -66
rect 548 -67 549 -55
rect 576 -67 577 -55
rect 590 -98 591 -66
rect 604 -98 605 -66
rect 628 -98 629 -66
rect 681 -67 682 -55
rect 723 -98 724 -66
rect 324 -98 325 -68
rect 534 -98 535 -68
rect 555 -69 556 -55
rect 576 -98 577 -68
rect 611 -69 612 -55
rect 618 -98 619 -68
rect 621 -69 622 -55
rect 688 -98 689 -68
rect 373 -98 374 -70
rect 443 -71 444 -55
rect 485 -71 486 -55
rect 548 -98 549 -70
rect 572 -71 573 -55
rect 611 -98 612 -70
rect 614 -71 615 -55
rect 667 -98 668 -70
rect 674 -71 675 -55
rect 681 -98 682 -70
rect 436 -73 437 -55
rect 443 -98 444 -72
rect 457 -73 458 -55
rect 485 -98 486 -72
rect 520 -98 521 -72
rect 639 -98 640 -72
rect 383 -98 384 -74
rect 457 -98 458 -74
rect 541 -75 542 -55
rect 555 -98 556 -74
rect 422 -77 423 -55
rect 436 -98 437 -76
rect 422 -98 423 -78
rect 492 -79 493 -55
rect 429 -81 430 -55
rect 492 -98 493 -80
rect 415 -83 416 -55
rect 429 -98 430 -82
rect 415 -98 416 -84
rect 450 -85 451 -55
rect 331 -87 332 -55
rect 450 -98 451 -86
rect 331 -98 332 -88
rect 359 -89 360 -55
rect 352 -91 353 -55
rect 359 -98 360 -90
rect 352 -98 353 -92
rect 366 -93 367 -55
rect 366 -98 367 -94
rect 394 -95 395 -55
rect 394 -98 395 -96
rect 782 -98 783 -96
rect 114 -165 115 -107
rect 191 -108 192 -106
rect 198 -165 199 -107
rect 296 -165 297 -107
rect 299 -108 300 -106
rect 390 -108 391 -106
rect 471 -108 472 -106
rect 562 -108 563 -106
rect 565 -108 566 -106
rect 695 -165 696 -107
rect 723 -108 724 -106
rect 786 -108 787 -106
rect 793 -108 794 -106
rect 856 -165 857 -107
rect 891 -108 892 -106
rect 919 -165 920 -107
rect 1010 -165 1011 -107
rect 1136 -165 1137 -107
rect 121 -165 122 -109
rect 383 -110 384 -106
rect 387 -110 388 -106
rect 450 -110 451 -106
rect 509 -110 510 -106
rect 562 -165 563 -109
rect 569 -110 570 -106
rect 569 -165 570 -109
rect 569 -110 570 -106
rect 569 -165 570 -109
rect 572 -165 573 -109
rect 744 -165 745 -109
rect 782 -110 783 -106
rect 1171 -165 1172 -109
rect 135 -165 136 -111
rect 299 -165 300 -111
rect 334 -165 335 -111
rect 723 -165 724 -111
rect 737 -112 738 -106
rect 842 -165 843 -111
rect 898 -112 899 -106
rect 940 -165 941 -111
rect 1017 -112 1018 -106
rect 1024 -165 1025 -111
rect 142 -165 143 -113
rect 520 -114 521 -106
rect 537 -114 538 -106
rect 821 -165 822 -113
rect 863 -114 864 -106
rect 898 -165 899 -113
rect 149 -165 150 -115
rect 373 -116 374 -106
rect 380 -165 381 -115
rect 541 -116 542 -106
rect 558 -165 559 -115
rect 604 -116 605 -106
rect 611 -116 612 -106
rect 772 -165 773 -115
rect 800 -116 801 -106
rect 877 -165 878 -115
rect 156 -165 157 -117
rect 310 -118 311 -106
rect 369 -165 370 -117
rect 534 -165 535 -117
rect 583 -118 584 -106
rect 590 -118 591 -106
rect 593 -165 594 -117
rect 758 -165 759 -117
rect 807 -118 808 -106
rect 870 -165 871 -117
rect 163 -165 164 -119
rect 205 -120 206 -106
rect 212 -165 213 -119
rect 453 -165 454 -119
rect 516 -120 517 -106
rect 800 -165 801 -119
rect 863 -165 864 -119
rect 1013 -165 1014 -119
rect 170 -165 171 -121
rect 289 -122 290 -106
rect 310 -165 311 -121
rect 408 -122 409 -106
rect 443 -122 444 -106
rect 471 -165 472 -121
rect 614 -165 615 -121
rect 737 -165 738 -121
rect 177 -165 178 -123
rect 229 -165 230 -123
rect 240 -165 241 -123
rect 303 -124 304 -106
rect 408 -165 409 -123
rect 604 -165 605 -123
rect 618 -124 619 -106
rect 793 -165 794 -123
rect 184 -165 185 -125
rect 219 -126 220 -106
rect 226 -165 227 -125
rect 513 -126 514 -106
rect 586 -126 587 -106
rect 618 -165 619 -125
rect 625 -126 626 -106
rect 849 -165 850 -125
rect 191 -165 192 -127
rect 394 -128 395 -106
rect 415 -128 416 -106
rect 443 -165 444 -127
rect 450 -165 451 -127
rect 499 -128 500 -106
rect 513 -165 514 -127
rect 541 -165 542 -127
rect 576 -128 577 -106
rect 625 -165 626 -127
rect 628 -128 629 -106
rect 716 -165 717 -127
rect 205 -165 206 -129
rect 233 -130 234 -106
rect 247 -130 248 -106
rect 373 -165 374 -129
rect 394 -165 395 -129
rect 548 -130 549 -106
rect 639 -130 640 -106
rect 779 -165 780 -129
rect 219 -165 220 -131
rect 324 -132 325 -106
rect 415 -165 416 -131
rect 506 -132 507 -106
rect 639 -165 640 -131
rect 646 -132 647 -106
rect 660 -132 661 -106
rect 765 -165 766 -131
rect 233 -165 234 -133
rect 611 -165 612 -133
rect 667 -134 668 -106
rect 751 -165 752 -133
rect 247 -165 248 -135
rect 257 -136 258 -106
rect 261 -136 262 -106
rect 261 -165 262 -135
rect 261 -136 262 -106
rect 261 -165 262 -135
rect 268 -165 269 -135
rect 422 -136 423 -106
rect 464 -136 465 -106
rect 516 -165 517 -135
rect 597 -136 598 -106
rect 646 -165 647 -135
rect 681 -136 682 -106
rect 681 -165 682 -135
rect 681 -136 682 -106
rect 681 -165 682 -135
rect 688 -136 689 -106
rect 814 -165 815 -135
rect 271 -138 272 -106
rect 275 -138 276 -106
rect 282 -138 283 -106
rect 282 -165 283 -137
rect 282 -138 283 -106
rect 282 -165 283 -137
rect 289 -165 290 -137
rect 530 -165 531 -137
rect 555 -138 556 -106
rect 597 -165 598 -137
rect 632 -138 633 -106
rect 667 -165 668 -137
rect 702 -138 703 -106
rect 807 -165 808 -137
rect 275 -165 276 -139
rect 338 -140 339 -106
rect 390 -165 391 -139
rect 422 -165 423 -139
rect 464 -165 465 -139
rect 527 -140 528 -106
rect 555 -165 556 -139
rect 674 -165 675 -139
rect 702 -165 703 -139
rect 730 -140 731 -106
rect 303 -165 304 -141
rect 523 -165 524 -141
rect 527 -165 528 -141
rect 828 -165 829 -141
rect 324 -165 325 -143
rect 352 -144 353 -106
rect 478 -144 479 -106
rect 660 -165 661 -143
rect 730 -165 731 -143
rect 835 -165 836 -143
rect 338 -165 339 -145
rect 366 -146 367 -106
rect 478 -165 479 -145
rect 485 -146 486 -106
rect 492 -146 493 -106
rect 548 -165 549 -145
rect 632 -165 633 -145
rect 709 -146 710 -106
rect 128 -165 129 -147
rect 366 -165 367 -147
rect 457 -148 458 -106
rect 485 -165 486 -147
rect 492 -165 493 -147
rect 502 -165 503 -147
rect 653 -148 654 -106
rect 688 -165 689 -147
rect 345 -150 346 -106
rect 352 -165 353 -149
rect 436 -150 437 -106
rect 457 -165 458 -149
rect 499 -165 500 -149
rect 576 -165 577 -149
rect 583 -165 584 -149
rect 653 -165 654 -149
rect 656 -165 657 -149
rect 709 -165 710 -149
rect 345 -165 346 -151
rect 401 -152 402 -106
rect 359 -154 360 -106
rect 436 -165 437 -153
rect 359 -165 360 -155
rect 429 -156 430 -106
rect 317 -158 318 -106
rect 429 -165 430 -157
rect 254 -160 255 -106
rect 317 -165 318 -159
rect 401 -165 402 -159
rect 786 -165 787 -159
rect 254 -165 255 -161
rect 331 -162 332 -106
rect 331 -165 332 -163
rect 506 -165 507 -163
rect 72 -232 73 -174
rect 569 -175 570 -173
rect 597 -175 598 -173
rect 600 -191 601 -174
rect 709 -175 710 -173
rect 884 -232 885 -174
rect 898 -175 899 -173
rect 933 -232 934 -174
rect 940 -175 941 -173
rect 989 -232 990 -174
rect 1024 -175 1025 -173
rect 1038 -232 1039 -174
rect 1136 -175 1137 -173
rect 1185 -232 1186 -174
rect 86 -232 87 -176
rect 656 -177 657 -173
rect 751 -177 752 -173
rect 1017 -232 1018 -176
rect 1171 -177 1172 -173
rect 1325 -232 1326 -176
rect 93 -232 94 -178
rect 268 -179 269 -173
rect 275 -179 276 -173
rect 296 -179 297 -173
rect 310 -179 311 -173
rect 453 -232 454 -178
rect 457 -179 458 -173
rect 457 -232 458 -178
rect 457 -179 458 -173
rect 457 -232 458 -178
rect 478 -179 479 -173
rect 530 -179 531 -173
rect 548 -179 549 -173
rect 590 -232 591 -178
rect 597 -232 598 -178
rect 632 -179 633 -173
rect 772 -179 773 -173
rect 912 -232 913 -178
rect 919 -179 920 -173
rect 982 -232 983 -178
rect 100 -232 101 -180
rect 198 -181 199 -173
rect 205 -181 206 -173
rect 401 -181 402 -173
rect 446 -232 447 -180
rect 940 -232 941 -180
rect 107 -232 108 -182
rect 415 -183 416 -173
rect 513 -183 514 -173
rect 772 -232 773 -182
rect 793 -183 794 -173
rect 1003 -232 1004 -182
rect 114 -185 115 -173
rect 208 -232 209 -184
rect 222 -232 223 -184
rect 891 -232 892 -184
rect 121 -187 122 -173
rect 236 -232 237 -186
rect 240 -187 241 -173
rect 334 -187 335 -173
rect 401 -232 402 -186
rect 478 -232 479 -186
rect 520 -187 521 -173
rect 730 -232 731 -186
rect 800 -187 801 -173
rect 898 -232 899 -186
rect 121 -232 122 -188
rect 142 -189 143 -173
rect 149 -189 150 -173
rect 569 -232 570 -188
rect 576 -189 577 -173
rect 709 -232 710 -188
rect 716 -189 717 -173
rect 793 -232 794 -188
rect 807 -189 808 -173
rect 926 -232 927 -188
rect 142 -232 143 -190
rect 506 -191 507 -173
rect 523 -191 524 -173
rect 593 -191 594 -173
rect 632 -232 633 -190
rect 674 -191 675 -173
rect 919 -232 920 -190
rect 149 -232 150 -192
rect 184 -193 185 -173
rect 191 -193 192 -173
rect 527 -232 528 -192
rect 534 -193 535 -173
rect 576 -232 577 -192
rect 625 -193 626 -173
rect 674 -232 675 -192
rect 681 -193 682 -173
rect 716 -232 717 -192
rect 737 -193 738 -173
rect 800 -232 801 -192
rect 814 -193 815 -173
rect 1010 -232 1011 -192
rect 79 -232 80 -194
rect 625 -232 626 -194
rect 681 -232 682 -194
rect 688 -195 689 -173
rect 702 -195 703 -173
rect 737 -232 738 -194
rect 744 -195 745 -173
rect 814 -232 815 -194
rect 821 -195 822 -173
rect 961 -232 962 -194
rect 163 -197 164 -173
rect 275 -232 276 -196
rect 282 -197 283 -173
rect 282 -232 283 -196
rect 282 -197 283 -173
rect 282 -232 283 -196
rect 289 -197 290 -173
rect 296 -232 297 -196
rect 310 -232 311 -196
rect 390 -197 391 -173
rect 422 -197 423 -173
rect 513 -232 514 -196
rect 555 -232 556 -196
rect 614 -232 615 -196
rect 667 -197 668 -173
rect 744 -232 745 -196
rect 828 -197 829 -173
rect 947 -232 948 -196
rect 163 -232 164 -198
rect 177 -199 178 -173
rect 184 -232 185 -198
rect 219 -199 220 -173
rect 233 -199 234 -173
rect 415 -232 416 -198
rect 432 -232 433 -198
rect 807 -232 808 -198
rect 835 -199 836 -173
rect 905 -232 906 -198
rect 114 -232 115 -200
rect 219 -232 220 -200
rect 233 -232 234 -200
rect 369 -201 370 -173
rect 436 -201 437 -173
rect 520 -232 521 -200
rect 558 -201 559 -173
rect 653 -232 654 -200
rect 688 -232 689 -200
rect 751 -232 752 -200
rect 765 -201 766 -173
rect 835 -232 836 -200
rect 856 -201 857 -173
rect 968 -232 969 -200
rect 170 -203 171 -173
rect 198 -232 199 -202
rect 243 -232 244 -202
rect 422 -232 423 -202
rect 464 -203 465 -173
rect 534 -232 535 -202
rect 562 -203 563 -173
rect 604 -232 605 -202
rect 618 -203 619 -173
rect 765 -232 766 -202
rect 870 -203 871 -173
rect 975 -232 976 -202
rect 156 -205 157 -173
rect 170 -232 171 -204
rect 177 -232 178 -204
rect 404 -205 405 -173
rect 443 -205 444 -173
rect 464 -232 465 -204
rect 471 -205 472 -173
rect 667 -232 668 -204
rect 702 -232 703 -204
rect 758 -205 759 -173
rect 786 -205 787 -173
rect 870 -232 871 -204
rect 877 -205 878 -173
rect 1024 -232 1025 -204
rect 128 -207 129 -173
rect 443 -232 444 -206
rect 471 -232 472 -206
rect 492 -207 493 -173
rect 607 -207 608 -173
rect 758 -232 759 -206
rect 842 -207 843 -173
rect 877 -232 878 -206
rect 128 -232 129 -208
rect 226 -209 227 -173
rect 229 -232 230 -208
rect 842 -232 843 -208
rect 191 -232 192 -210
rect 205 -232 206 -210
rect 261 -211 262 -173
rect 268 -232 269 -210
rect 289 -232 290 -210
rect 352 -211 353 -173
rect 387 -211 388 -173
rect 786 -232 787 -210
rect 247 -213 248 -173
rect 261 -232 262 -212
rect 331 -213 332 -173
rect 338 -213 339 -173
rect 352 -232 353 -212
rect 366 -232 367 -212
rect 380 -213 381 -173
rect 387 -232 388 -212
rect 394 -213 395 -173
rect 436 -232 437 -212
rect 485 -213 486 -173
rect 506 -232 507 -212
rect 618 -232 619 -212
rect 646 -213 647 -173
rect 660 -213 661 -173
rect 856 -232 857 -212
rect 212 -215 213 -173
rect 338 -232 339 -214
rect 373 -215 374 -173
rect 380 -232 381 -214
rect 394 -232 395 -214
rect 551 -232 552 -214
rect 611 -215 612 -173
rect 660 -232 661 -214
rect 723 -215 724 -173
rect 821 -232 822 -214
rect 212 -232 213 -216
rect 499 -217 500 -173
rect 611 -232 612 -216
rect 954 -232 955 -216
rect 247 -232 248 -218
rect 324 -219 325 -173
rect 359 -219 360 -173
rect 373 -232 374 -218
rect 429 -219 430 -173
rect 646 -232 647 -218
rect 723 -232 724 -218
rect 863 -219 864 -173
rect 135 -221 136 -173
rect 429 -232 430 -220
rect 492 -232 493 -220
rect 541 -221 542 -173
rect 779 -221 780 -173
rect 863 -232 864 -220
rect 135 -232 136 -222
rect 254 -223 255 -173
rect 317 -223 318 -173
rect 331 -232 332 -222
rect 345 -223 346 -173
rect 359 -232 360 -222
rect 499 -232 500 -222
rect 562 -232 563 -222
rect 695 -223 696 -173
rect 779 -232 780 -222
rect 254 -232 255 -224
rect 303 -225 304 -173
rect 317 -232 318 -224
rect 408 -225 409 -173
rect 541 -232 542 -224
rect 639 -225 640 -173
rect 695 -232 696 -224
rect 831 -232 832 -224
rect 303 -232 304 -226
rect 450 -227 451 -173
rect 583 -227 584 -173
rect 639 -232 640 -226
rect 324 -232 325 -228
rect 485 -232 486 -228
rect 583 -232 584 -228
rect 849 -229 850 -173
rect 345 -232 346 -230
rect 408 -232 409 -230
rect 450 -232 451 -230
rect 628 -232 629 -230
rect 849 -232 850 -230
rect 996 -232 997 -230
rect 93 -242 94 -240
rect 485 -242 486 -240
rect 488 -242 489 -240
rect 856 -242 857 -240
rect 884 -242 885 -240
rect 1115 -315 1116 -241
rect 1185 -242 1186 -240
rect 1206 -315 1207 -241
rect 1307 -315 1308 -241
rect 1458 -315 1459 -241
rect 93 -315 94 -243
rect 142 -244 143 -240
rect 145 -315 146 -243
rect 401 -244 402 -240
rect 446 -244 447 -240
rect 492 -244 493 -240
rect 502 -244 503 -240
rect 912 -244 913 -240
rect 919 -244 920 -240
rect 1052 -315 1053 -243
rect 1325 -244 1326 -240
rect 1381 -315 1382 -243
rect 100 -246 101 -240
rect 173 -315 174 -245
rect 177 -246 178 -240
rect 478 -246 479 -240
rect 485 -315 486 -245
rect 747 -315 748 -245
rect 754 -246 755 -240
rect 1080 -315 1081 -245
rect 100 -315 101 -247
rect 236 -248 237 -240
rect 247 -248 248 -240
rect 401 -315 402 -247
rect 453 -248 454 -240
rect 1003 -248 1004 -240
rect 1038 -248 1039 -240
rect 1066 -315 1067 -247
rect 107 -250 108 -240
rect 443 -315 444 -249
rect 492 -315 493 -249
rect 506 -250 507 -240
rect 537 -315 538 -249
rect 1101 -315 1102 -249
rect 107 -315 108 -251
rect 142 -315 143 -251
rect 159 -252 160 -240
rect 257 -252 258 -240
rect 268 -252 269 -240
rect 268 -315 269 -251
rect 268 -252 269 -240
rect 268 -315 269 -251
rect 303 -252 304 -240
rect 551 -252 552 -240
rect 600 -315 601 -251
rect 912 -315 913 -251
rect 954 -252 955 -240
rect 1108 -315 1109 -251
rect 128 -254 129 -240
rect 240 -315 241 -253
rect 247 -315 248 -253
rect 366 -254 367 -240
rect 369 -254 370 -240
rect 457 -254 458 -240
rect 506 -315 507 -253
rect 527 -254 528 -240
rect 551 -315 552 -253
rect 618 -254 619 -240
rect 628 -254 629 -240
rect 919 -315 920 -253
rect 968 -254 969 -240
rect 1031 -315 1032 -253
rect 79 -256 80 -240
rect 128 -315 129 -255
rect 138 -315 139 -255
rect 688 -256 689 -240
rect 737 -256 738 -240
rect 751 -315 752 -255
rect 765 -256 766 -240
rect 1094 -315 1095 -255
rect 79 -315 80 -257
rect 149 -258 150 -240
rect 163 -258 164 -240
rect 177 -315 178 -257
rect 191 -258 192 -240
rect 194 -266 195 -257
rect 205 -258 206 -240
rect 226 -258 227 -240
rect 233 -315 234 -257
rect 289 -258 290 -240
rect 303 -315 304 -257
rect 576 -258 577 -240
rect 618 -315 619 -257
rect 628 -315 629 -257
rect 632 -258 633 -240
rect 688 -315 689 -257
rect 716 -258 717 -240
rect 737 -315 738 -257
rect 786 -258 787 -240
rect 856 -315 857 -257
rect 877 -258 878 -240
rect 954 -315 955 -257
rect 975 -258 976 -240
rect 1073 -315 1074 -257
rect 114 -260 115 -240
rect 149 -315 150 -259
rect 163 -315 164 -259
rect 184 -260 185 -240
rect 191 -315 192 -259
rect 219 -260 220 -240
rect 226 -315 227 -259
rect 562 -260 563 -240
rect 632 -315 633 -259
rect 1017 -260 1018 -240
rect 114 -315 115 -261
rect 121 -262 122 -240
rect 170 -262 171 -240
rect 499 -262 500 -240
rect 541 -262 542 -240
rect 562 -315 563 -261
rect 670 -315 671 -261
rect 807 -262 808 -240
rect 821 -262 822 -240
rect 884 -315 885 -261
rect 891 -262 892 -240
rect 1045 -315 1046 -261
rect 121 -315 122 -263
rect 352 -264 353 -240
rect 366 -315 367 -263
rect 373 -264 374 -240
rect 376 -315 377 -263
rect 520 -264 521 -240
rect 541 -315 542 -263
rect 555 -264 556 -240
rect 674 -264 675 -240
rect 968 -315 969 -263
rect 982 -264 983 -240
rect 1038 -315 1039 -263
rect 219 -315 220 -265
rect 289 -315 290 -265
rect 394 -266 395 -240
rect 450 -266 451 -240
rect 527 -315 528 -265
rect 646 -266 647 -240
rect 674 -315 675 -265
rect 695 -266 696 -240
rect 716 -315 717 -265
rect 779 -266 780 -240
rect 821 -315 822 -265
rect 835 -266 836 -240
rect 891 -315 892 -265
rect 905 -266 906 -240
rect 1003 -315 1004 -265
rect 198 -268 199 -240
rect 576 -315 577 -267
rect 625 -315 626 -267
rect 779 -315 780 -267
rect 793 -268 794 -240
rect 877 -315 878 -267
rect 905 -315 906 -267
rect 1024 -268 1025 -240
rect 198 -315 199 -269
rect 261 -270 262 -240
rect 331 -270 332 -240
rect 352 -315 353 -269
rect 380 -270 381 -240
rect 555 -315 556 -269
rect 646 -315 647 -269
rect 982 -315 983 -269
rect 989 -270 990 -240
rect 1059 -315 1060 -269
rect 208 -272 209 -240
rect 261 -315 262 -271
rect 380 -315 381 -271
rect 1122 -315 1123 -271
rect 86 -274 87 -240
rect 208 -315 209 -273
rect 212 -274 213 -240
rect 331 -315 332 -273
rect 383 -315 384 -273
rect 604 -274 605 -240
rect 709 -274 710 -240
rect 786 -315 787 -273
rect 898 -274 899 -240
rect 989 -315 990 -273
rect 996 -274 997 -240
rect 1087 -315 1088 -273
rect 86 -315 87 -275
rect 429 -276 430 -240
rect 450 -315 451 -275
rect 548 -315 549 -275
rect 604 -315 605 -275
rect 1010 -276 1011 -240
rect 184 -315 185 -277
rect 212 -315 213 -277
rect 387 -278 388 -240
rect 408 -315 409 -277
rect 415 -278 416 -240
rect 429 -315 430 -277
rect 457 -315 458 -277
rect 464 -278 465 -240
rect 478 -315 479 -277
rect 765 -315 766 -277
rect 926 -278 927 -240
rect 1010 -315 1011 -277
rect 187 -315 188 -279
rect 464 -315 465 -279
rect 499 -315 500 -279
rect 597 -280 598 -240
rect 607 -315 608 -279
rect 926 -315 927 -279
rect 933 -280 934 -240
rect 975 -315 976 -279
rect 317 -282 318 -240
rect 415 -315 416 -281
rect 513 -282 514 -240
rect 520 -315 521 -281
rect 534 -282 535 -240
rect 597 -315 598 -281
rect 611 -282 612 -240
rect 709 -315 710 -281
rect 723 -282 724 -240
rect 793 -315 794 -281
rect 842 -282 843 -240
rect 933 -315 934 -281
rect 940 -282 941 -240
rect 1017 -315 1018 -281
rect 65 -315 66 -283
rect 534 -315 535 -283
rect 590 -284 591 -240
rect 611 -315 612 -283
rect 660 -284 661 -240
rect 723 -315 724 -283
rect 744 -284 745 -240
rect 898 -315 899 -283
rect 947 -284 948 -240
rect 996 -315 997 -283
rect 317 -315 318 -285
rect 324 -286 325 -240
rect 387 -315 388 -285
rect 849 -286 850 -240
rect 863 -286 864 -240
rect 940 -315 941 -285
rect 961 -286 962 -240
rect 1024 -315 1025 -285
rect 324 -315 325 -287
rect 345 -288 346 -240
rect 390 -315 391 -287
rect 667 -288 668 -240
rect 744 -315 745 -287
rect 835 -315 836 -287
rect 870 -288 871 -240
rect 947 -315 948 -287
rect 72 -290 73 -240
rect 345 -315 346 -289
rect 394 -315 395 -289
rect 471 -290 472 -240
rect 590 -315 591 -289
rect 870 -315 871 -289
rect 72 -315 73 -291
rect 156 -292 157 -240
rect 275 -292 276 -240
rect 471 -315 472 -291
rect 653 -292 654 -240
rect 660 -315 661 -291
rect 667 -315 668 -291
rect 772 -292 773 -240
rect 800 -292 801 -240
rect 842 -315 843 -291
rect 156 -315 157 -293
rect 254 -294 255 -240
rect 275 -315 276 -293
rect 296 -294 297 -240
rect 411 -294 412 -240
rect 849 -315 850 -293
rect 170 -315 171 -295
rect 800 -315 801 -295
rect 814 -296 815 -240
rect 863 -315 864 -295
rect 254 -315 255 -297
rect 373 -315 374 -297
rect 422 -298 423 -240
rect 513 -315 514 -297
rect 639 -298 640 -240
rect 653 -315 654 -297
rect 730 -298 731 -240
rect 814 -315 815 -297
rect 828 -298 829 -240
rect 961 -315 962 -297
rect 282 -300 283 -240
rect 296 -315 297 -299
rect 422 -315 423 -299
rect 436 -300 437 -240
rect 481 -300 482 -240
rect 772 -315 773 -299
rect 135 -302 136 -240
rect 282 -315 283 -301
rect 583 -302 584 -240
rect 639 -315 640 -301
rect 681 -302 682 -240
rect 730 -315 731 -301
rect 758 -302 759 -240
rect 828 -315 829 -301
rect 243 -304 244 -240
rect 436 -315 437 -303
rect 446 -315 447 -303
rect 758 -315 759 -303
rect 569 -306 570 -240
rect 583 -315 584 -305
rect 681 -315 682 -305
rect 702 -306 703 -240
rect 338 -308 339 -240
rect 569 -315 570 -307
rect 695 -315 696 -307
rect 702 -315 703 -307
rect 338 -315 339 -309
rect 359 -310 360 -240
rect 310 -312 311 -240
rect 359 -315 360 -311
rect 310 -315 311 -313
rect 807 -315 808 -313
rect 65 -325 66 -323
rect 380 -414 381 -324
rect 446 -325 447 -323
rect 576 -325 577 -323
rect 590 -325 591 -323
rect 1094 -325 1095 -323
rect 1101 -325 1102 -323
rect 1213 -414 1214 -324
rect 1381 -325 1382 -323
rect 1409 -414 1410 -324
rect 1458 -325 1459 -323
rect 1521 -414 1522 -324
rect 72 -327 73 -323
rect 362 -414 363 -326
rect 369 -414 370 -326
rect 569 -327 570 -323
rect 597 -327 598 -323
rect 898 -327 899 -323
rect 912 -327 913 -323
rect 1150 -414 1151 -326
rect 1171 -414 1172 -326
rect 1223 -414 1224 -326
rect 72 -414 73 -328
rect 121 -329 122 -323
rect 135 -414 136 -328
rect 289 -329 290 -323
rect 345 -329 346 -323
rect 534 -329 535 -323
rect 548 -329 549 -323
rect 1052 -329 1053 -323
rect 1059 -329 1060 -323
rect 1164 -414 1165 -328
rect 1199 -414 1200 -328
rect 1307 -329 1308 -323
rect 79 -331 80 -323
rect 187 -331 188 -323
rect 205 -331 206 -323
rect 1108 -331 1109 -323
rect 1122 -331 1123 -323
rect 1388 -414 1389 -330
rect 58 -414 59 -332
rect 205 -414 206 -332
rect 250 -414 251 -332
rect 534 -414 535 -332
rect 541 -333 542 -323
rect 548 -414 549 -332
rect 551 -333 552 -323
rect 968 -333 969 -323
rect 989 -333 990 -323
rect 1122 -414 1123 -332
rect 1206 -333 1207 -323
rect 1206 -414 1207 -332
rect 1206 -333 1207 -323
rect 1206 -414 1207 -332
rect 79 -414 80 -334
rect 149 -335 150 -323
rect 166 -414 167 -334
rect 576 -414 577 -334
rect 597 -414 598 -334
rect 789 -414 790 -334
rect 807 -335 808 -323
rect 898 -414 899 -334
rect 926 -335 927 -323
rect 989 -414 990 -334
rect 1003 -335 1004 -323
rect 1129 -414 1130 -334
rect 86 -337 87 -323
rect 383 -337 384 -323
rect 478 -414 479 -336
rect 541 -414 542 -336
rect 565 -414 566 -336
rect 1178 -414 1179 -336
rect 86 -414 87 -338
rect 593 -339 594 -323
rect 604 -339 605 -323
rect 618 -339 619 -323
rect 625 -339 626 -323
rect 1045 -339 1046 -323
rect 1066 -339 1067 -323
rect 1108 -414 1109 -338
rect 93 -341 94 -323
rect 537 -341 538 -323
rect 618 -414 619 -340
rect 660 -341 661 -323
rect 667 -414 668 -340
rect 688 -341 689 -323
rect 702 -341 703 -323
rect 744 -414 745 -340
rect 821 -341 822 -323
rect 968 -414 969 -340
rect 975 -341 976 -323
rect 1045 -414 1046 -340
rect 1073 -341 1074 -323
rect 1185 -414 1186 -340
rect 93 -414 94 -342
rect 418 -414 419 -342
rect 464 -343 465 -323
rect 604 -414 605 -342
rect 625 -414 626 -342
rect 807 -414 808 -342
rect 835 -343 836 -323
rect 912 -414 913 -342
rect 961 -343 962 -323
rect 1003 -414 1004 -342
rect 1017 -343 1018 -323
rect 1143 -414 1144 -342
rect 100 -345 101 -323
rect 187 -414 188 -344
rect 191 -345 192 -323
rect 383 -414 384 -344
rect 464 -414 465 -344
rect 555 -345 556 -323
rect 583 -345 584 -323
rect 660 -414 661 -344
rect 702 -414 703 -344
rect 786 -345 787 -323
rect 856 -345 857 -323
rect 926 -414 927 -344
rect 947 -345 948 -323
rect 1017 -414 1018 -344
rect 1024 -345 1025 -323
rect 1094 -414 1095 -344
rect 100 -414 101 -346
rect 156 -347 157 -323
rect 170 -347 171 -323
rect 849 -347 850 -323
rect 856 -414 857 -346
rect 905 -347 906 -323
rect 947 -414 948 -346
rect 1010 -347 1011 -323
rect 1031 -347 1032 -323
rect 1136 -414 1137 -346
rect 121 -414 122 -348
rect 128 -349 129 -323
rect 149 -414 150 -348
rect 310 -349 311 -323
rect 345 -414 346 -348
rect 450 -349 451 -323
rect 495 -414 496 -348
rect 513 -349 514 -323
rect 555 -414 556 -348
rect 653 -349 654 -323
rect 758 -349 759 -323
rect 849 -414 850 -348
rect 870 -349 871 -323
rect 1052 -414 1053 -348
rect 1080 -349 1081 -323
rect 1192 -414 1193 -348
rect 128 -414 129 -350
rect 303 -351 304 -323
rect 310 -414 311 -350
rect 359 -351 360 -323
rect 373 -414 374 -350
rect 485 -351 486 -323
rect 506 -351 507 -323
rect 590 -414 591 -350
rect 628 -351 629 -323
rect 730 -351 731 -323
rect 765 -351 766 -323
rect 821 -414 822 -350
rect 884 -351 885 -323
rect 961 -414 962 -350
rect 982 -351 983 -323
rect 1066 -414 1067 -350
rect 1080 -414 1081 -350
rect 1115 -351 1116 -323
rect 173 -353 174 -323
rect 569 -414 570 -352
rect 583 -414 584 -352
rect 765 -414 766 -352
rect 772 -353 773 -323
rect 1031 -414 1032 -352
rect 1038 -353 1039 -323
rect 1059 -414 1060 -352
rect 1087 -353 1088 -323
rect 1157 -414 1158 -352
rect 107 -355 108 -323
rect 1087 -414 1088 -354
rect 107 -414 108 -356
rect 114 -357 115 -323
rect 173 -414 174 -356
rect 506 -414 507 -356
rect 513 -414 514 -356
rect 527 -357 528 -323
rect 632 -357 633 -323
rect 649 -357 650 -323
rect 709 -357 710 -323
rect 772 -414 773 -356
rect 786 -414 787 -356
rect 1101 -414 1102 -356
rect 114 -414 115 -358
rect 471 -359 472 -323
rect 481 -359 482 -323
rect 653 -414 654 -358
rect 730 -414 731 -358
rect 800 -359 801 -323
rect 814 -359 815 -323
rect 905 -414 906 -358
rect 919 -359 920 -323
rect 982 -414 983 -358
rect 996 -359 997 -323
rect 1024 -414 1025 -358
rect 184 -361 185 -323
rect 1073 -414 1074 -360
rect 138 -363 139 -323
rect 184 -414 185 -362
rect 194 -414 195 -362
rect 485 -414 486 -362
rect 520 -363 521 -323
rect 527 -414 528 -362
rect 572 -414 573 -362
rect 814 -414 815 -362
rect 828 -363 829 -323
rect 884 -414 885 -362
rect 891 -363 892 -323
rect 975 -414 976 -362
rect 247 -365 248 -323
rect 758 -414 759 -364
rect 793 -365 794 -323
rect 828 -414 829 -364
rect 842 -365 843 -323
rect 891 -414 892 -364
rect 940 -365 941 -323
rect 1010 -414 1011 -364
rect 156 -414 157 -366
rect 247 -414 248 -366
rect 282 -367 283 -323
rect 390 -367 391 -323
rect 415 -367 416 -323
rect 520 -414 521 -366
rect 646 -414 647 -366
rect 835 -414 836 -366
rect 842 -414 843 -366
rect 933 -367 934 -323
rect 954 -367 955 -323
rect 1038 -414 1039 -366
rect 142 -369 143 -323
rect 415 -414 416 -368
rect 436 -369 437 -323
rect 450 -414 451 -368
rect 586 -414 587 -368
rect 933 -414 934 -368
rect 142 -414 143 -370
rect 163 -371 164 -323
rect 233 -371 234 -323
rect 282 -414 283 -370
rect 289 -414 290 -370
rect 691 -414 692 -370
rect 723 -371 724 -323
rect 793 -414 794 -370
rect 863 -371 864 -323
rect 940 -414 941 -370
rect 233 -414 234 -372
rect 635 -414 636 -372
rect 670 -373 671 -323
rect 996 -414 997 -372
rect 303 -414 304 -374
rect 338 -375 339 -323
rect 376 -375 377 -323
rect 471 -414 472 -374
rect 737 -375 738 -323
rect 919 -414 920 -374
rect 261 -377 262 -323
rect 338 -414 339 -376
rect 387 -377 388 -323
rect 800 -414 801 -376
rect 877 -377 878 -323
rect 954 -414 955 -376
rect 212 -379 213 -323
rect 261 -414 262 -378
rect 313 -379 314 -323
rect 387 -414 388 -378
rect 408 -379 409 -323
rect 723 -414 724 -378
rect 747 -379 748 -323
rect 1115 -414 1116 -378
rect 212 -414 213 -380
rect 219 -381 220 -323
rect 366 -381 367 -323
rect 408 -414 409 -380
rect 436 -414 437 -380
rect 611 -381 612 -323
rect 716 -381 717 -323
rect 737 -414 738 -380
rect 779 -381 780 -323
rect 863 -414 864 -380
rect 177 -383 178 -323
rect 219 -414 220 -382
rect 443 -383 444 -323
rect 709 -414 710 -382
rect 716 -414 717 -382
rect 870 -414 871 -382
rect 177 -414 178 -384
rect 254 -385 255 -323
rect 422 -385 423 -323
rect 443 -414 444 -384
rect 562 -385 563 -323
rect 611 -414 612 -384
rect 751 -385 752 -323
rect 779 -414 780 -384
rect 240 -387 241 -323
rect 422 -414 423 -386
rect 600 -387 601 -323
rect 877 -414 878 -386
rect 240 -414 241 -388
rect 394 -389 395 -323
rect 632 -414 633 -388
rect 751 -414 752 -388
rect 254 -414 255 -390
rect 268 -391 269 -323
rect 394 -414 395 -390
rect 401 -391 402 -323
rect 198 -393 199 -323
rect 268 -414 269 -392
rect 401 -414 402 -392
rect 695 -393 696 -323
rect 198 -414 199 -394
rect 492 -395 493 -323
rect 681 -395 682 -323
rect 695 -414 696 -394
rect 275 -397 276 -323
rect 492 -414 493 -396
rect 639 -397 640 -323
rect 681 -414 682 -396
rect 275 -414 276 -398
rect 324 -399 325 -323
rect 639 -414 640 -398
rect 674 -399 675 -323
rect 324 -414 325 -400
rect 331 -401 332 -323
rect 499 -401 500 -323
rect 674 -414 675 -400
rect 226 -403 227 -323
rect 499 -414 500 -402
rect 226 -414 227 -404
rect 317 -405 318 -323
rect 331 -414 332 -404
rect 352 -405 353 -323
rect 296 -407 297 -323
rect 317 -414 318 -406
rect 352 -414 353 -406
rect 457 -407 458 -323
rect 208 -409 209 -323
rect 457 -414 458 -408
rect 296 -414 297 -410
rect 429 -411 430 -323
rect 429 -414 430 -412
rect 688 -414 689 -412
rect 51 -503 52 -423
rect 187 -424 188 -422
rect 194 -424 195 -422
rect 758 -424 759 -422
rect 838 -424 839 -422
rect 1213 -424 1214 -422
rect 1388 -424 1389 -422
rect 1486 -503 1487 -423
rect 1521 -424 1522 -422
rect 1542 -503 1543 -423
rect 58 -503 59 -425
rect 145 -503 146 -425
rect 149 -426 150 -422
rect 212 -426 213 -422
rect 250 -426 251 -422
rect 317 -426 318 -422
rect 359 -426 360 -422
rect 590 -426 591 -422
rect 611 -426 612 -422
rect 621 -503 622 -425
rect 656 -503 657 -425
rect 730 -426 731 -422
rect 754 -503 755 -425
rect 1122 -426 1123 -422
rect 1157 -426 1158 -422
rect 1227 -503 1228 -425
rect 1409 -426 1410 -422
rect 1430 -503 1431 -425
rect 65 -503 66 -427
rect 121 -428 122 -422
rect 124 -503 125 -427
rect 1143 -428 1144 -422
rect 1185 -428 1186 -422
rect 1213 -503 1214 -427
rect 72 -430 73 -422
rect 425 -503 426 -429
rect 450 -430 451 -422
rect 541 -430 542 -422
rect 544 -430 545 -422
rect 793 -430 794 -422
rect 856 -430 857 -422
rect 856 -503 857 -429
rect 856 -430 857 -422
rect 856 -503 857 -429
rect 891 -430 892 -422
rect 891 -503 892 -429
rect 891 -430 892 -422
rect 891 -503 892 -429
rect 919 -430 920 -422
rect 1234 -503 1235 -429
rect 72 -503 73 -431
rect 562 -432 563 -422
rect 572 -432 573 -422
rect 702 -432 703 -422
rect 737 -432 738 -422
rect 793 -503 794 -431
rect 870 -432 871 -422
rect 919 -503 920 -431
rect 996 -432 997 -422
rect 996 -503 997 -431
rect 996 -432 997 -422
rect 996 -503 997 -431
rect 1073 -432 1074 -422
rect 1157 -503 1158 -431
rect 1192 -432 1193 -422
rect 1241 -503 1242 -431
rect 79 -434 80 -422
rect 79 -503 80 -433
rect 79 -434 80 -422
rect 79 -503 80 -433
rect 86 -434 87 -422
rect 173 -434 174 -422
rect 177 -434 178 -422
rect 390 -503 391 -433
rect 415 -434 416 -422
rect 520 -434 521 -422
rect 541 -503 542 -433
rect 674 -434 675 -422
rect 688 -434 689 -422
rect 842 -434 843 -422
rect 1031 -434 1032 -422
rect 1073 -503 1074 -433
rect 1080 -434 1081 -422
rect 1255 -503 1256 -433
rect 86 -503 87 -435
rect 107 -436 108 -422
rect 114 -436 115 -422
rect 149 -503 150 -435
rect 163 -436 164 -422
rect 422 -436 423 -422
rect 450 -503 451 -435
rect 551 -503 552 -435
rect 558 -503 559 -435
rect 618 -436 619 -422
rect 628 -436 629 -422
rect 702 -503 703 -435
rect 821 -436 822 -422
rect 870 -503 871 -435
rect 1108 -436 1109 -422
rect 1185 -503 1186 -435
rect 1206 -436 1207 -422
rect 1223 -436 1224 -422
rect 93 -438 94 -422
rect 684 -503 685 -437
rect 691 -438 692 -422
rect 1129 -438 1130 -422
rect 1136 -438 1137 -422
rect 1143 -503 1144 -437
rect 1164 -438 1165 -422
rect 1192 -503 1193 -437
rect 93 -503 94 -439
rect 100 -440 101 -422
rect 114 -503 115 -439
rect 436 -440 437 -422
rect 464 -440 465 -422
rect 520 -503 521 -439
rect 548 -440 549 -422
rect 562 -503 563 -439
rect 583 -440 584 -422
rect 968 -440 969 -422
rect 1101 -440 1102 -422
rect 1129 -503 1130 -439
rect 1164 -503 1165 -439
rect 1199 -440 1200 -422
rect 100 -503 101 -441
rect 198 -442 199 -422
rect 212 -503 213 -441
rect 275 -442 276 -422
rect 296 -442 297 -422
rect 586 -442 587 -422
rect 590 -503 591 -441
rect 646 -442 647 -422
rect 663 -503 664 -441
rect 786 -503 787 -441
rect 824 -503 825 -441
rect 1080 -503 1081 -441
rect 1115 -442 1116 -422
rect 1122 -503 1123 -441
rect 1171 -442 1172 -422
rect 1206 -503 1207 -441
rect 121 -503 122 -443
rect 1087 -444 1088 -422
rect 1094 -444 1095 -422
rect 1115 -503 1116 -443
rect 1150 -444 1151 -422
rect 1171 -503 1172 -443
rect 135 -446 136 -422
rect 492 -503 493 -445
rect 495 -446 496 -422
rect 1108 -503 1109 -445
rect 107 -503 108 -447
rect 135 -503 136 -447
rect 138 -503 139 -447
rect 845 -503 846 -447
rect 852 -503 853 -447
rect 1031 -503 1032 -447
rect 1045 -448 1046 -422
rect 1087 -503 1088 -447
rect 142 -450 143 -422
rect 163 -503 164 -449
rect 166 -450 167 -422
rect 247 -450 248 -422
rect 257 -503 258 -449
rect 338 -450 339 -422
rect 359 -503 360 -449
rect 513 -450 514 -422
rect 548 -503 549 -449
rect 604 -450 605 -422
rect 632 -450 633 -422
rect 1150 -503 1151 -449
rect 152 -452 153 -422
rect 338 -503 339 -451
rect 366 -452 367 -422
rect 730 -503 731 -451
rect 947 -452 948 -422
rect 1094 -503 1095 -451
rect 166 -503 167 -453
rect 1220 -454 1221 -422
rect 170 -503 171 -455
rect 299 -503 300 -455
rect 317 -503 318 -455
rect 324 -456 325 -422
rect 366 -503 367 -455
rect 569 -456 570 -422
rect 632 -503 633 -455
rect 1251 -503 1252 -455
rect 177 -503 178 -457
rect 625 -458 626 -422
rect 667 -458 668 -422
rect 758 -503 759 -457
rect 905 -458 906 -422
rect 947 -503 948 -457
rect 968 -503 969 -457
rect 982 -458 983 -422
rect 1024 -458 1025 -422
rect 1101 -503 1102 -457
rect 184 -503 185 -459
rect 219 -460 220 -422
rect 247 -503 248 -459
rect 593 -503 594 -459
rect 667 -503 668 -459
rect 751 -460 752 -422
rect 835 -460 836 -422
rect 905 -503 906 -459
rect 961 -460 962 -422
rect 982 -503 983 -459
rect 989 -460 990 -422
rect 1024 -503 1025 -459
rect 1038 -460 1039 -422
rect 1045 -503 1046 -459
rect 191 -462 192 -422
rect 194 -503 195 -461
rect 219 -503 220 -461
rect 352 -462 353 -422
rect 380 -462 381 -422
rect 604 -503 605 -461
rect 695 -462 696 -422
rect 737 -503 738 -461
rect 779 -462 780 -422
rect 835 -503 836 -461
rect 898 -462 899 -422
rect 989 -503 990 -461
rect 1017 -462 1018 -422
rect 1038 -503 1039 -461
rect 142 -503 143 -463
rect 779 -503 780 -463
rect 814 -464 815 -422
rect 898 -503 899 -463
rect 954 -464 955 -422
rect 961 -503 962 -463
rect 1010 -464 1011 -422
rect 1017 -503 1018 -463
rect 191 -503 192 -465
rect 674 -503 675 -465
rect 698 -503 699 -465
rect 1052 -466 1053 -422
rect 261 -468 262 -422
rect 324 -503 325 -467
rect 331 -468 332 -422
rect 352 -503 353 -467
rect 383 -468 384 -422
rect 394 -468 395 -422
rect 401 -468 402 -422
rect 436 -503 437 -467
rect 464 -503 465 -467
rect 660 -468 661 -422
rect 723 -468 724 -422
rect 1199 -503 1200 -467
rect 261 -503 262 -469
rect 310 -470 311 -422
rect 345 -470 346 -422
rect 380 -503 381 -469
rect 394 -503 395 -469
rect 408 -470 409 -422
rect 415 -503 416 -469
rect 618 -503 619 -469
rect 726 -470 727 -422
rect 1136 -503 1137 -469
rect 275 -503 276 -471
rect 282 -472 283 -422
rect 296 -503 297 -471
rect 387 -472 388 -422
rect 408 -503 409 -471
rect 821 -503 822 -471
rect 877 -472 878 -422
rect 1010 -503 1011 -471
rect 156 -474 157 -422
rect 282 -503 283 -473
rect 303 -474 304 -422
rect 331 -503 332 -473
rect 345 -503 346 -473
rect 467 -503 468 -473
rect 471 -474 472 -422
rect 513 -503 514 -473
rect 569 -503 570 -473
rect 751 -503 752 -473
rect 765 -474 766 -422
rect 814 -503 815 -473
rect 940 -474 941 -422
rect 954 -503 955 -473
rect 1003 -474 1004 -422
rect 1052 -503 1053 -473
rect 198 -503 199 -475
rect 387 -503 388 -475
rect 418 -476 419 -422
rect 716 -503 717 -475
rect 744 -476 745 -422
rect 765 -503 766 -475
rect 800 -476 801 -422
rect 877 -503 878 -475
rect 912 -476 913 -422
rect 1003 -503 1004 -475
rect 303 -503 304 -477
rect 649 -503 650 -477
rect 653 -478 654 -422
rect 744 -503 745 -477
rect 772 -478 773 -422
rect 800 -503 801 -477
rect 863 -478 864 -422
rect 940 -503 941 -477
rect 310 -503 311 -479
rect 404 -503 405 -479
rect 422 -503 423 -479
rect 681 -480 682 -422
rect 807 -480 808 -422
rect 863 -503 864 -479
rect 884 -480 885 -422
rect 912 -503 913 -479
rect 429 -482 430 -422
rect 471 -503 472 -481
rect 478 -482 479 -422
rect 611 -503 612 -481
rect 653 -503 654 -481
rect 688 -503 689 -481
rect 709 -482 710 -422
rect 807 -503 808 -481
rect 828 -482 829 -422
rect 884 -503 885 -481
rect 226 -484 227 -422
rect 429 -503 430 -483
rect 478 -503 479 -483
rect 499 -484 500 -422
rect 506 -484 507 -422
rect 583 -503 584 -483
rect 597 -484 598 -422
rect 828 -503 829 -483
rect 226 -503 227 -485
rect 240 -486 241 -422
rect 373 -486 374 -422
rect 506 -503 507 -485
rect 534 -486 535 -422
rect 709 -503 710 -485
rect 205 -488 206 -422
rect 240 -503 241 -487
rect 373 -503 374 -487
rect 443 -488 444 -422
rect 485 -488 486 -422
rect 597 -503 598 -487
rect 681 -503 682 -487
rect 1178 -488 1179 -422
rect 128 -490 129 -422
rect 485 -503 486 -489
rect 499 -503 500 -489
rect 719 -490 720 -422
rect 1059 -490 1060 -422
rect 1178 -503 1179 -489
rect 128 -503 129 -491
rect 362 -492 363 -422
rect 443 -503 444 -491
rect 457 -492 458 -422
rect 527 -492 528 -422
rect 534 -503 535 -491
rect 555 -492 556 -422
rect 772 -503 773 -491
rect 1059 -503 1060 -491
rect 1066 -492 1067 -422
rect 205 -503 206 -493
rect 233 -494 234 -422
rect 289 -494 290 -422
rect 527 -503 528 -493
rect 555 -503 556 -493
rect 625 -503 626 -493
rect 975 -494 976 -422
rect 1066 -503 1067 -493
rect 268 -496 269 -422
rect 289 -503 290 -495
rect 457 -503 458 -495
rect 789 -496 790 -422
rect 933 -496 934 -422
rect 975 -503 976 -495
rect 254 -498 255 -422
rect 268 -503 269 -497
rect 576 -498 577 -422
rect 723 -503 724 -497
rect 926 -498 927 -422
rect 933 -503 934 -497
rect 156 -503 157 -499
rect 254 -503 255 -499
rect 576 -503 577 -499
rect 639 -500 640 -422
rect 849 -500 850 -422
rect 926 -503 927 -499
rect 369 -502 370 -422
rect 639 -503 640 -501
rect 44 -624 45 -512
rect 86 -513 87 -511
rect 93 -513 94 -511
rect 1388 -624 1389 -512
rect 1419 -624 1420 -512
rect 1619 -624 1620 -512
rect 58 -515 59 -511
rect 646 -515 647 -511
rect 649 -515 650 -511
rect 1262 -624 1263 -514
rect 1430 -515 1431 -511
rect 1458 -624 1459 -514
rect 1486 -515 1487 -511
rect 1528 -624 1529 -514
rect 1542 -515 1543 -511
rect 1549 -624 1550 -514
rect 58 -624 59 -516
rect 747 -624 748 -516
rect 751 -517 752 -511
rect 1073 -517 1074 -511
rect 1087 -517 1088 -511
rect 1220 -624 1221 -516
rect 1227 -517 1228 -511
rect 1437 -624 1438 -516
rect 65 -519 66 -511
rect 191 -519 192 -511
rect 254 -624 255 -518
rect 380 -519 381 -511
rect 387 -519 388 -511
rect 1157 -519 1158 -511
rect 1178 -519 1179 -511
rect 1360 -624 1361 -518
rect 65 -624 66 -520
rect 236 -624 237 -520
rect 264 -624 265 -520
rect 1318 -624 1319 -520
rect 72 -523 73 -511
rect 327 -624 328 -522
rect 401 -624 402 -522
rect 569 -523 570 -511
rect 590 -523 591 -511
rect 849 -624 850 -522
rect 863 -523 864 -511
rect 1451 -624 1452 -522
rect 72 -624 73 -524
rect 660 -525 661 -511
rect 663 -525 664 -511
rect 898 -525 899 -511
rect 905 -525 906 -511
rect 1332 -624 1333 -524
rect 86 -624 87 -526
rect 149 -527 150 -511
rect 156 -527 157 -511
rect 380 -624 381 -526
rect 425 -527 426 -511
rect 569 -624 570 -526
rect 593 -527 594 -511
rect 1066 -527 1067 -511
rect 1115 -527 1116 -511
rect 1304 -624 1305 -526
rect 93 -624 94 -528
rect 233 -529 234 -511
rect 268 -529 269 -511
rect 292 -624 293 -528
rect 296 -529 297 -511
rect 425 -624 426 -528
rect 450 -529 451 -511
rect 590 -624 591 -528
rect 618 -529 619 -511
rect 1444 -624 1445 -528
rect 121 -624 122 -530
rect 390 -531 391 -511
rect 429 -531 430 -511
rect 450 -624 451 -530
rect 520 -531 521 -511
rect 520 -624 521 -530
rect 520 -531 521 -511
rect 520 -624 521 -530
rect 527 -531 528 -511
rect 618 -624 619 -530
rect 621 -531 622 -511
rect 1374 -624 1375 -530
rect 128 -533 129 -511
rect 698 -533 699 -511
rect 730 -533 731 -511
rect 803 -624 804 -532
rect 821 -533 822 -511
rect 1465 -624 1466 -532
rect 128 -624 129 -534
rect 205 -535 206 -511
rect 296 -624 297 -534
rect 642 -624 643 -534
rect 646 -624 647 -534
rect 1017 -535 1018 -511
rect 1024 -535 1025 -511
rect 1430 -624 1431 -534
rect 124 -537 125 -511
rect 205 -624 206 -536
rect 299 -537 300 -511
rect 506 -537 507 -511
rect 534 -537 535 -511
rect 548 -624 549 -536
rect 555 -537 556 -511
rect 765 -537 766 -511
rect 789 -624 790 -536
rect 1283 -624 1284 -536
rect 135 -624 136 -538
rect 656 -539 657 -511
rect 660 -624 661 -538
rect 1223 -539 1224 -511
rect 1241 -539 1242 -511
rect 1251 -539 1252 -511
rect 142 -541 143 -511
rect 184 -541 185 -511
rect 191 -624 192 -540
rect 226 -541 227 -511
rect 359 -541 360 -511
rect 527 -624 528 -540
rect 555 -624 556 -540
rect 709 -541 710 -511
rect 716 -541 717 -511
rect 821 -624 822 -540
rect 856 -541 857 -511
rect 898 -624 899 -540
rect 933 -541 934 -511
rect 1290 -624 1291 -540
rect 142 -624 143 -542
rect 457 -543 458 -511
rect 471 -543 472 -511
rect 534 -624 535 -542
rect 625 -543 626 -511
rect 716 -624 717 -542
rect 744 -543 745 -511
rect 863 -624 864 -542
rect 873 -624 874 -542
rect 989 -543 990 -511
rect 1010 -543 1011 -511
rect 1087 -624 1088 -542
rect 1122 -543 1123 -511
rect 1353 -624 1354 -542
rect 114 -545 115 -511
rect 625 -624 626 -544
rect 653 -545 654 -511
rect 1094 -545 1095 -511
rect 1129 -545 1130 -511
rect 1241 -624 1242 -544
rect 100 -547 101 -511
rect 114 -624 115 -546
rect 145 -547 146 -511
rect 1423 -624 1424 -546
rect 100 -624 101 -548
rect 107 -549 108 -511
rect 149 -624 150 -548
rect 289 -549 290 -511
rect 359 -624 360 -548
rect 394 -549 395 -511
rect 471 -624 472 -548
rect 583 -549 584 -511
rect 632 -549 633 -511
rect 653 -624 654 -548
rect 667 -549 668 -511
rect 905 -624 906 -548
rect 919 -549 920 -511
rect 989 -624 990 -548
rect 1017 -624 1018 -548
rect 1164 -549 1165 -511
rect 1185 -549 1186 -511
rect 1311 -624 1312 -548
rect 156 -624 157 -550
rect 649 -624 650 -550
rect 674 -551 675 -511
rect 751 -624 752 -550
rect 754 -551 755 -511
rect 1269 -624 1270 -550
rect 110 -624 111 -552
rect 674 -624 675 -552
rect 684 -553 685 -511
rect 1248 -624 1249 -552
rect 163 -555 164 -511
rect 1339 -624 1340 -554
rect 163 -624 164 -556
rect 233 -624 234 -556
rect 268 -624 269 -556
rect 457 -624 458 -556
rect 478 -557 479 -511
rect 632 -624 633 -556
rect 684 -624 685 -556
rect 1003 -557 1004 -511
rect 1024 -624 1025 -556
rect 1255 -557 1256 -511
rect 166 -559 167 -511
rect 247 -559 248 -511
rect 355 -624 356 -558
rect 583 -624 584 -558
rect 611 -559 612 -511
rect 667 -624 668 -558
rect 688 -559 689 -511
rect 765 -624 766 -558
rect 800 -559 801 -511
rect 1115 -624 1116 -558
rect 1143 -559 1144 -511
rect 1367 -624 1368 -558
rect 177 -561 178 -511
rect 177 -624 178 -560
rect 177 -561 178 -511
rect 177 -624 178 -560
rect 184 -624 185 -560
rect 303 -561 304 -511
rect 373 -561 374 -511
rect 429 -624 430 -560
rect 443 -561 444 -511
rect 611 -624 612 -560
rect 698 -624 699 -560
rect 1234 -561 1235 -511
rect 194 -563 195 -511
rect 1234 -624 1235 -562
rect 219 -565 220 -511
rect 373 -624 374 -564
rect 394 -624 395 -564
rect 597 -565 598 -511
rect 702 -565 703 -511
rect 709 -624 710 -564
rect 744 -624 745 -564
rect 1276 -624 1277 -564
rect 219 -624 220 -566
rect 345 -567 346 -511
rect 366 -567 367 -511
rect 443 -624 444 -566
rect 478 -624 479 -566
rect 1227 -624 1228 -566
rect 198 -569 199 -511
rect 345 -624 346 -568
rect 366 -624 367 -568
rect 415 -569 416 -511
rect 485 -569 486 -511
rect 702 -624 703 -568
rect 758 -569 759 -511
rect 856 -624 857 -568
rect 884 -569 885 -511
rect 933 -624 934 -568
rect 954 -569 955 -511
rect 1003 -624 1004 -568
rect 1034 -624 1035 -568
rect 1094 -624 1095 -568
rect 1108 -569 1109 -511
rect 1164 -624 1165 -568
rect 1171 -569 1172 -511
rect 1185 -624 1186 -568
rect 1192 -569 1193 -511
rect 1381 -624 1382 -568
rect 226 -624 227 -570
rect 324 -571 325 -511
rect 495 -624 496 -570
rect 688 -624 689 -570
rect 761 -624 762 -570
rect 1192 -624 1193 -570
rect 1199 -571 1200 -511
rect 1395 -624 1396 -570
rect 247 -624 248 -572
rect 331 -573 332 -511
rect 506 -624 507 -572
rect 513 -573 514 -511
rect 562 -573 563 -511
rect 597 -624 598 -572
rect 828 -573 829 -511
rect 884 -624 885 -572
rect 891 -573 892 -511
rect 1010 -624 1011 -572
rect 1031 -573 1032 -511
rect 1199 -624 1200 -572
rect 1206 -573 1207 -511
rect 1325 -624 1326 -572
rect 303 -624 304 -574
rect 758 -624 759 -574
rect 786 -575 787 -511
rect 828 -624 829 -574
rect 835 -575 836 -511
rect 891 -624 892 -574
rect 926 -575 927 -511
rect 954 -624 955 -574
rect 961 -575 962 -511
rect 1073 -624 1074 -574
rect 1080 -575 1081 -511
rect 1255 -624 1256 -574
rect 310 -577 311 -511
rect 415 -624 416 -576
rect 481 -624 482 -576
rect 926 -624 927 -576
rect 968 -577 969 -511
rect 1157 -624 1158 -576
rect 1213 -577 1214 -511
rect 1409 -624 1410 -576
rect 240 -579 241 -511
rect 310 -624 311 -578
rect 324 -624 325 -578
rect 1122 -624 1123 -578
rect 1136 -579 1137 -511
rect 1206 -624 1207 -578
rect 240 -624 241 -580
rect 282 -581 283 -511
rect 331 -624 332 -580
rect 460 -624 461 -580
rect 492 -581 493 -511
rect 513 -624 514 -580
rect 723 -581 724 -511
rect 835 -624 836 -580
rect 842 -581 843 -511
rect 919 -624 920 -580
rect 940 -581 941 -511
rect 968 -624 969 -580
rect 975 -581 976 -511
rect 1143 -624 1144 -580
rect 1150 -581 1151 -511
rect 1346 -624 1347 -580
rect 261 -583 262 -511
rect 282 -624 283 -582
rect 317 -583 318 -511
rect 492 -624 493 -582
rect 499 -583 500 -511
rect 1213 -624 1214 -582
rect 79 -585 80 -511
rect 261 -624 262 -584
rect 275 -585 276 -511
rect 317 -624 318 -584
rect 576 -585 577 -511
rect 975 -624 976 -584
rect 982 -585 983 -511
rect 1402 -624 1403 -584
rect 79 -624 80 -586
rect 485 -624 486 -586
rect 639 -587 640 -511
rect 723 -624 724 -586
rect 824 -587 825 -511
rect 1080 -624 1081 -586
rect 1101 -587 1102 -511
rect 1150 -624 1151 -586
rect 275 -624 276 -588
rect 422 -589 423 -511
rect 436 -589 437 -511
rect 576 -624 577 -588
rect 639 -624 640 -588
rect 772 -589 773 -511
rect 870 -589 871 -511
rect 961 -624 962 -588
rect 996 -589 997 -511
rect 1108 -624 1109 -588
rect 51 -591 52 -511
rect 422 -624 423 -590
rect 467 -591 468 -511
rect 1101 -624 1102 -590
rect 51 -624 52 -592
rect 170 -593 171 -511
rect 289 -624 290 -592
rect 499 -624 500 -592
rect 562 -624 563 -592
rect 870 -624 871 -592
rect 912 -593 913 -511
rect 996 -624 997 -592
rect 1038 -593 1039 -511
rect 1129 -624 1130 -592
rect 107 -624 108 -594
rect 436 -624 437 -594
rect 681 -624 682 -594
rect 940 -624 941 -594
rect 1045 -595 1046 -511
rect 1171 -624 1172 -594
rect 170 -624 171 -596
rect 198 -624 199 -596
rect 390 -624 391 -596
rect 982 -624 983 -596
rect 1052 -597 1053 -511
rect 1178 -624 1179 -596
rect 772 -624 773 -598
rect 807 -599 808 -511
rect 814 -599 815 -511
rect 912 -624 913 -598
rect 947 -599 948 -511
rect 1045 -624 1046 -598
rect 1059 -599 1060 -511
rect 1136 -624 1137 -598
rect 607 -624 608 -600
rect 807 -624 808 -600
rect 845 -601 846 -511
rect 1052 -624 1053 -600
rect 695 -603 696 -511
rect 1059 -624 1060 -602
rect 695 -624 696 -604
rect 1066 -624 1067 -604
rect 737 -607 738 -511
rect 814 -624 815 -606
rect 845 -624 846 -606
rect 1297 -624 1298 -606
rect 604 -609 605 -511
rect 737 -624 738 -608
rect 779 -609 780 -511
rect 1038 -624 1039 -608
rect 464 -611 465 -511
rect 604 -624 605 -610
rect 779 -624 780 -610
rect 852 -611 853 -511
rect 877 -611 878 -511
rect 947 -624 948 -610
rect 408 -613 409 -511
rect 464 -624 465 -612
rect 793 -613 794 -511
rect 877 -624 878 -612
rect 338 -615 339 -511
rect 408 -624 409 -614
rect 338 -624 339 -616
rect 352 -617 353 -511
rect 404 -617 405 -511
rect 793 -624 794 -616
rect 212 -619 213 -511
rect 352 -624 353 -618
rect 212 -624 213 -620
rect 541 -621 542 -511
rect 387 -624 388 -622
rect 541 -624 542 -622
rect 65 -634 66 -632
rect 264 -634 265 -632
rect 310 -634 311 -632
rect 324 -634 325 -632
rect 334 -757 335 -633
rect 422 -634 423 -632
rect 523 -757 524 -633
rect 611 -634 612 -632
rect 618 -634 619 -632
rect 681 -634 682 -632
rect 691 -757 692 -633
rect 779 -634 780 -632
rect 786 -634 787 -632
rect 1339 -634 1340 -632
rect 1419 -634 1420 -632
rect 1458 -634 1459 -632
rect 1549 -634 1550 -632
rect 1556 -757 1557 -633
rect 1619 -634 1620 -632
rect 1696 -757 1697 -633
rect 72 -636 73 -632
rect 639 -757 640 -635
rect 646 -757 647 -635
rect 1479 -757 1480 -635
rect 1528 -636 1529 -632
rect 1549 -757 1550 -635
rect 68 -757 69 -637
rect 72 -757 73 -637
rect 100 -638 101 -632
rect 100 -757 101 -637
rect 100 -638 101 -632
rect 100 -757 101 -637
rect 121 -638 122 -632
rect 635 -757 636 -637
rect 649 -757 650 -637
rect 772 -638 773 -632
rect 831 -757 832 -637
rect 1409 -638 1410 -632
rect 1444 -638 1445 -632
rect 1458 -757 1459 -637
rect 1465 -638 1466 -632
rect 1528 -757 1529 -637
rect 121 -757 122 -639
rect 212 -640 213 -632
rect 222 -757 223 -639
rect 1227 -640 1228 -632
rect 1276 -640 1277 -632
rect 1486 -757 1487 -639
rect 128 -642 129 -632
rect 233 -642 234 -632
rect 240 -642 241 -632
rect 481 -642 482 -632
rect 485 -642 486 -632
rect 772 -757 773 -641
rect 838 -757 839 -641
rect 1143 -642 1144 -632
rect 1360 -642 1361 -632
rect 1409 -757 1410 -641
rect 1437 -642 1438 -632
rect 1444 -757 1445 -641
rect 128 -757 129 -643
rect 282 -644 283 -632
rect 296 -644 297 -632
rect 422 -757 423 -643
rect 429 -644 430 -632
rect 485 -757 486 -643
rect 548 -644 549 -632
rect 548 -757 549 -643
rect 548 -644 549 -632
rect 548 -757 549 -643
rect 555 -644 556 -632
rect 607 -644 608 -632
rect 674 -644 675 -632
rect 1227 -757 1228 -643
rect 1423 -644 1424 -632
rect 1437 -757 1438 -643
rect 159 -757 160 -645
rect 975 -646 976 -632
rect 982 -646 983 -632
rect 1143 -757 1144 -645
rect 1164 -646 1165 -632
rect 1360 -757 1361 -645
rect 117 -757 118 -647
rect 982 -757 983 -647
rect 1017 -648 1018 -632
rect 1374 -648 1375 -632
rect 79 -650 80 -632
rect 1017 -757 1018 -649
rect 1052 -650 1053 -632
rect 1276 -757 1277 -649
rect 1318 -650 1319 -632
rect 1423 -757 1424 -649
rect 58 -652 59 -632
rect 79 -757 80 -651
rect 191 -652 192 -632
rect 618 -757 619 -651
rect 674 -757 675 -651
rect 1297 -652 1298 -632
rect 93 -654 94 -632
rect 191 -757 192 -653
rect 198 -654 199 -632
rect 1269 -654 1270 -632
rect 93 -757 94 -655
rect 156 -656 157 -632
rect 198 -757 199 -655
rect 359 -656 360 -632
rect 394 -656 395 -632
rect 457 -656 458 -632
rect 492 -656 493 -632
rect 975 -757 976 -655
rect 1066 -656 1067 -632
rect 1164 -757 1165 -655
rect 1192 -656 1193 -632
rect 1269 -757 1270 -655
rect 114 -658 115 -632
rect 492 -757 493 -657
rect 555 -757 556 -657
rect 856 -658 857 -632
rect 870 -757 871 -657
rect 1430 -658 1431 -632
rect 44 -660 45 -632
rect 114 -757 115 -659
rect 201 -660 202 -632
rect 1234 -660 1235 -632
rect 1255 -660 1256 -632
rect 1297 -757 1298 -659
rect 44 -757 45 -661
rect 373 -662 374 -632
rect 457 -757 458 -661
rect 842 -662 843 -632
rect 845 -662 846 -632
rect 1325 -662 1326 -632
rect 205 -664 206 -632
rect 240 -757 241 -663
rect 247 -664 248 -632
rect 324 -757 325 -663
rect 345 -664 346 -632
rect 572 -757 573 -663
rect 590 -664 591 -632
rect 695 -757 696 -663
rect 709 -664 710 -632
rect 779 -757 780 -663
rect 800 -664 801 -632
rect 1318 -757 1319 -663
rect 149 -666 150 -632
rect 247 -757 248 -665
rect 282 -757 283 -665
rect 289 -666 290 -632
rect 296 -757 297 -665
rect 331 -666 332 -632
rect 345 -757 346 -665
rect 607 -757 608 -665
rect 677 -757 678 -665
rect 1290 -666 1291 -632
rect 149 -757 150 -667
rect 751 -668 752 -632
rect 758 -668 759 -632
rect 1451 -668 1452 -632
rect 212 -757 213 -669
rect 219 -670 220 -632
rect 226 -670 227 -632
rect 478 -670 479 -632
rect 495 -757 496 -669
rect 842 -757 843 -669
rect 926 -670 927 -632
rect 1066 -757 1067 -669
rect 1108 -670 1109 -632
rect 1465 -757 1466 -669
rect 219 -757 220 -671
rect 800 -757 801 -671
rect 803 -757 804 -671
rect 1374 -757 1375 -671
rect 1395 -672 1396 -632
rect 1451 -757 1452 -671
rect 226 -757 227 -673
rect 261 -674 262 -632
rect 275 -674 276 -632
rect 289 -757 290 -673
rect 310 -757 311 -673
rect 366 -674 367 -632
rect 478 -757 479 -673
rect 534 -674 535 -632
rect 569 -674 570 -632
rect 611 -757 612 -673
rect 653 -674 654 -632
rect 758 -757 759 -673
rect 828 -674 829 -632
rect 856 -757 857 -673
rect 933 -674 934 -632
rect 1031 -757 1032 -673
rect 1038 -674 1039 -632
rect 1192 -757 1193 -673
rect 1206 -674 1207 -632
rect 1255 -757 1256 -673
rect 1283 -674 1284 -632
rect 1290 -757 1291 -673
rect 1304 -674 1305 -632
rect 1395 -757 1396 -673
rect 170 -676 171 -632
rect 366 -757 367 -675
rect 471 -676 472 -632
rect 653 -757 654 -675
rect 681 -757 682 -675
rect 737 -676 738 -632
rect 744 -676 745 -632
rect 1157 -676 1158 -632
rect 1220 -676 1221 -632
rect 1325 -757 1326 -675
rect 142 -678 143 -632
rect 471 -757 472 -677
rect 527 -678 528 -632
rect 534 -757 535 -677
rect 590 -757 591 -677
rect 625 -678 626 -632
rect 632 -678 633 -632
rect 744 -757 745 -677
rect 751 -757 752 -677
rect 905 -678 906 -632
rect 912 -678 913 -632
rect 933 -757 934 -677
rect 961 -678 962 -632
rect 1108 -757 1109 -677
rect 1122 -678 1123 -632
rect 1430 -757 1431 -677
rect 142 -757 143 -679
rect 436 -680 437 -632
rect 527 -757 528 -679
rect 940 -680 941 -632
rect 1059 -680 1060 -632
rect 1157 -757 1158 -679
rect 1248 -680 1249 -632
rect 1283 -757 1284 -679
rect 156 -757 157 -681
rect 1059 -757 1060 -681
rect 1080 -682 1081 -632
rect 1206 -757 1207 -681
rect 1262 -682 1263 -632
rect 1304 -757 1305 -681
rect 170 -757 171 -683
rect 450 -684 451 -632
rect 597 -684 598 -632
rect 625 -757 626 -683
rect 632 -757 633 -683
rect 1115 -684 1116 -632
rect 1129 -684 1130 -632
rect 1220 -757 1221 -683
rect 184 -686 185 -632
rect 569 -757 570 -685
rect 604 -686 605 -632
rect 1213 -686 1214 -632
rect 184 -757 185 -687
rect 303 -688 304 -632
rect 317 -688 318 -632
rect 387 -688 388 -632
rect 425 -688 426 -632
rect 737 -757 738 -687
rect 761 -688 762 -632
rect 1080 -757 1081 -687
rect 1087 -688 1088 -632
rect 1122 -757 1123 -687
rect 1136 -688 1137 -632
rect 1339 -757 1340 -687
rect 86 -690 87 -632
rect 387 -757 388 -689
rect 558 -757 559 -689
rect 597 -757 598 -689
rect 604 -757 605 -689
rect 1332 -690 1333 -632
rect 86 -757 87 -691
rect 107 -692 108 -632
rect 233 -757 234 -691
rect 352 -692 353 -632
rect 355 -692 356 -632
rect 394 -757 395 -691
rect 530 -757 531 -691
rect 1332 -757 1333 -691
rect 107 -757 108 -693
rect 789 -694 790 -632
rect 821 -694 822 -632
rect 1038 -757 1039 -693
rect 1094 -694 1095 -632
rect 1213 -757 1214 -693
rect 254 -696 255 -632
rect 352 -757 353 -695
rect 359 -757 360 -695
rect 464 -696 465 -632
rect 688 -696 689 -632
rect 786 -757 787 -695
rect 814 -696 815 -632
rect 821 -757 822 -695
rect 828 -757 829 -695
rect 1472 -757 1473 -695
rect 177 -698 178 -632
rect 814 -757 815 -697
rect 849 -698 850 -632
rect 940 -757 941 -697
rect 954 -698 955 -632
rect 1087 -757 1088 -697
rect 1150 -698 1151 -632
rect 1234 -757 1235 -697
rect 177 -757 178 -699
rect 327 -700 328 -632
rect 380 -700 381 -632
rect 450 -757 451 -699
rect 464 -757 465 -699
rect 1416 -700 1417 -632
rect 254 -757 255 -701
rect 373 -757 374 -701
rect 429 -757 430 -701
rect 954 -757 955 -701
rect 968 -702 969 -632
rect 1115 -757 1116 -701
rect 1178 -702 1179 -632
rect 1262 -757 1263 -701
rect 1388 -702 1389 -632
rect 1416 -757 1417 -701
rect 261 -757 262 -703
rect 338 -704 339 -632
rect 467 -757 468 -703
rect 968 -757 969 -703
rect 989 -704 990 -632
rect 1129 -757 1130 -703
rect 1178 -757 1179 -703
rect 1381 -704 1382 -632
rect 268 -706 269 -632
rect 338 -757 339 -705
rect 702 -706 703 -632
rect 709 -757 710 -705
rect 719 -757 720 -705
rect 1367 -706 1368 -632
rect 268 -757 269 -707
rect 401 -708 402 -632
rect 460 -708 461 -632
rect 702 -757 703 -707
rect 730 -708 731 -632
rect 1052 -757 1053 -707
rect 1185 -708 1186 -632
rect 1388 -757 1389 -707
rect 135 -710 136 -632
rect 401 -757 402 -709
rect 684 -710 685 -632
rect 1185 -757 1186 -709
rect 1311 -710 1312 -632
rect 1367 -757 1368 -709
rect 135 -757 136 -711
rect 205 -757 206 -711
rect 303 -757 304 -711
rect 415 -712 416 -632
rect 733 -712 734 -632
rect 1101 -712 1102 -632
rect 1346 -712 1347 -632
rect 1381 -757 1382 -711
rect 317 -757 318 -713
rect 408 -714 409 -632
rect 415 -757 416 -713
rect 499 -714 500 -632
rect 733 -757 734 -713
rect 1402 -714 1403 -632
rect 163 -716 164 -632
rect 408 -757 409 -715
rect 499 -757 500 -715
rect 576 -716 577 -632
rect 793 -716 794 -632
rect 849 -757 850 -715
rect 873 -716 874 -632
rect 1311 -757 1312 -715
rect 58 -757 59 -717
rect 163 -757 164 -717
rect 331 -757 332 -717
rect 380 -757 381 -717
rect 576 -757 577 -717
rect 716 -718 717 -632
rect 884 -718 885 -632
rect 912 -757 913 -717
rect 919 -718 920 -632
rect 961 -757 962 -717
rect 989 -757 990 -717
rect 1024 -718 1025 -632
rect 1045 -718 1046 -632
rect 1150 -757 1151 -717
rect 1171 -718 1172 -632
rect 1402 -757 1403 -717
rect 275 -757 276 -719
rect 716 -757 717 -719
rect 877 -720 878 -632
rect 1045 -757 1046 -719
rect 432 -757 433 -721
rect 884 -757 885 -721
rect 891 -722 892 -632
rect 919 -757 920 -721
rect 929 -757 930 -721
rect 1094 -757 1095 -721
rect 51 -724 52 -632
rect 891 -757 892 -723
rect 905 -757 906 -723
rect 1199 -724 1200 -632
rect 51 -757 52 -725
rect 243 -726 244 -632
rect 436 -757 437 -725
rect 1024 -757 1025 -725
rect 1073 -726 1074 -632
rect 1199 -757 1200 -725
rect 642 -728 643 -632
rect 1073 -757 1074 -727
rect 807 -730 808 -632
rect 877 -757 878 -729
rect 908 -757 909 -729
rect 1346 -757 1347 -729
rect 723 -732 724 -632
rect 807 -757 808 -731
rect 996 -732 997 -632
rect 1136 -757 1137 -731
rect 506 -734 507 -632
rect 723 -757 724 -733
rect 947 -734 948 -632
rect 996 -757 997 -733
rect 1003 -734 1004 -632
rect 1171 -757 1172 -733
rect 257 -757 258 -735
rect 506 -757 507 -735
rect 520 -736 521 -632
rect 1003 -757 1004 -735
rect 1010 -736 1011 -632
rect 1101 -757 1102 -735
rect 863 -738 864 -632
rect 947 -757 948 -737
rect 1020 -738 1021 -632
rect 1248 -757 1249 -737
rect 765 -740 766 -632
rect 863 -757 864 -739
rect 898 -740 899 -632
rect 1010 -757 1011 -739
rect 443 -742 444 -632
rect 765 -757 766 -741
rect 835 -742 836 -632
rect 898 -757 899 -741
rect 443 -757 444 -743
rect 660 -744 661 -632
rect 835 -757 836 -743
rect 1353 -744 1354 -632
rect 660 -757 661 -745
rect 667 -746 668 -632
rect 1241 -746 1242 -632
rect 1353 -757 1354 -745
rect 583 -748 584 -632
rect 667 -757 668 -747
rect 698 -748 699 -632
rect 1241 -757 1242 -747
rect 541 -750 542 -632
rect 583 -757 584 -749
rect 513 -752 514 -632
rect 541 -757 542 -751
rect 513 -757 514 -753
rect 562 -754 563 -632
rect 562 -757 563 -755
rect 796 -757 797 -755
rect 37 -870 38 -766
rect 51 -767 52 -765
rect 58 -870 59 -766
rect 562 -767 563 -765
rect 572 -767 573 -765
rect 1423 -767 1424 -765
rect 1430 -767 1431 -765
rect 1584 -870 1585 -766
rect 1696 -767 1697 -765
rect 1724 -870 1725 -766
rect 44 -769 45 -765
rect 432 -769 433 -765
rect 485 -769 486 -765
rect 530 -769 531 -765
rect 551 -870 552 -768
rect 737 -769 738 -765
rect 793 -769 794 -765
rect 1192 -769 1193 -765
rect 1255 -769 1256 -765
rect 1535 -870 1536 -768
rect 1549 -769 1550 -765
rect 1577 -870 1578 -768
rect 44 -870 45 -770
rect 61 -771 62 -765
rect 65 -771 66 -765
rect 345 -771 346 -765
rect 366 -771 367 -765
rect 646 -771 647 -765
rect 667 -771 668 -765
rect 716 -771 717 -765
rect 737 -870 738 -770
rect 947 -771 948 -765
rect 954 -771 955 -765
rect 954 -870 955 -770
rect 954 -771 955 -765
rect 954 -870 955 -770
rect 961 -771 962 -765
rect 1192 -870 1193 -770
rect 1297 -771 1298 -765
rect 1297 -870 1298 -770
rect 1297 -771 1298 -765
rect 1297 -870 1298 -770
rect 1332 -771 1333 -765
rect 1332 -870 1333 -770
rect 1332 -771 1333 -765
rect 1332 -870 1333 -770
rect 1353 -771 1354 -765
rect 1430 -870 1431 -770
rect 1437 -771 1438 -765
rect 1507 -870 1508 -770
rect 1528 -771 1529 -765
rect 1570 -870 1571 -770
rect 65 -870 66 -772
rect 72 -773 73 -765
rect 114 -870 115 -772
rect 359 -773 360 -765
rect 366 -870 367 -772
rect 513 -773 514 -765
rect 530 -870 531 -772
rect 548 -773 549 -765
rect 558 -773 559 -765
rect 1038 -773 1039 -765
rect 1108 -773 1109 -765
rect 1108 -870 1109 -772
rect 1108 -773 1109 -765
rect 1108 -870 1109 -772
rect 1115 -773 1116 -765
rect 1255 -870 1256 -772
rect 1262 -773 1263 -765
rect 1353 -870 1354 -772
rect 1409 -773 1410 -765
rect 1528 -870 1529 -772
rect 1556 -773 1557 -765
rect 1556 -870 1557 -772
rect 1556 -773 1557 -765
rect 1556 -870 1557 -772
rect 72 -870 73 -774
rect 93 -775 94 -765
rect 124 -870 125 -774
rect 289 -775 290 -765
rect 296 -775 297 -765
rect 555 -775 556 -765
rect 607 -775 608 -765
rect 772 -775 773 -765
rect 793 -870 794 -774
rect 877 -775 878 -765
rect 905 -775 906 -765
rect 1437 -870 1438 -774
rect 1444 -775 1445 -765
rect 1549 -870 1550 -774
rect 93 -870 94 -776
rect 184 -777 185 -765
rect 187 -870 188 -776
rect 310 -777 311 -765
rect 324 -777 325 -765
rect 359 -870 360 -776
rect 380 -777 381 -765
rect 555 -870 556 -776
rect 604 -777 605 -765
rect 905 -870 906 -776
rect 908 -777 909 -765
rect 1325 -777 1326 -765
rect 1367 -777 1368 -765
rect 1444 -870 1445 -776
rect 1458 -777 1459 -765
rect 1514 -870 1515 -776
rect 135 -779 136 -765
rect 331 -779 332 -765
rect 345 -870 346 -778
rect 352 -779 353 -765
rect 380 -870 381 -778
rect 457 -779 458 -765
rect 478 -779 479 -765
rect 513 -870 514 -778
rect 534 -779 535 -765
rect 604 -870 605 -778
rect 611 -779 612 -765
rect 677 -779 678 -765
rect 684 -870 685 -778
rect 922 -870 923 -778
rect 926 -779 927 -765
rect 1178 -779 1179 -765
rect 1220 -779 1221 -765
rect 1262 -870 1263 -778
rect 1290 -779 1291 -765
rect 1409 -870 1410 -778
rect 1416 -779 1417 -765
rect 1500 -870 1501 -778
rect 135 -870 136 -780
rect 156 -781 157 -765
rect 163 -781 164 -765
rect 331 -870 332 -780
rect 394 -781 395 -765
rect 478 -870 479 -780
rect 506 -781 507 -765
rect 828 -781 829 -765
rect 835 -781 836 -765
rect 856 -781 857 -765
rect 926 -870 927 -780
rect 989 -781 990 -765
rect 1017 -781 1018 -765
rect 1038 -870 1039 -780
rect 1115 -870 1116 -780
rect 1241 -781 1242 -765
rect 1346 -781 1347 -765
rect 1367 -870 1368 -780
rect 1374 -781 1375 -765
rect 1416 -870 1417 -780
rect 1472 -781 1473 -765
rect 1521 -870 1522 -780
rect 163 -870 164 -782
rect 782 -870 783 -782
rect 796 -783 797 -765
rect 1101 -783 1102 -765
rect 1150 -783 1151 -765
rect 1150 -870 1151 -782
rect 1150 -783 1151 -765
rect 1150 -870 1151 -782
rect 1157 -783 1158 -765
rect 1157 -870 1158 -782
rect 1157 -783 1158 -765
rect 1157 -870 1158 -782
rect 1171 -783 1172 -765
rect 1171 -870 1172 -782
rect 1171 -783 1172 -765
rect 1171 -870 1172 -782
rect 1178 -870 1179 -782
rect 1206 -783 1207 -765
rect 1213 -783 1214 -765
rect 1220 -870 1221 -782
rect 1227 -783 1228 -765
rect 1325 -870 1326 -782
rect 1479 -783 1480 -765
rect 1559 -870 1560 -782
rect 117 -785 118 -765
rect 1213 -870 1214 -784
rect 1241 -870 1242 -784
rect 1276 -785 1277 -765
rect 1311 -785 1312 -765
rect 1479 -870 1480 -784
rect 1486 -785 1487 -765
rect 1542 -870 1543 -784
rect 166 -870 167 -786
rect 674 -787 675 -765
rect 688 -787 689 -765
rect 1045 -787 1046 -765
rect 1059 -787 1060 -765
rect 1346 -870 1347 -786
rect 184 -870 185 -788
rect 1003 -789 1004 -765
rect 1024 -789 1025 -765
rect 1374 -870 1375 -788
rect 191 -791 192 -765
rect 464 -791 465 -765
rect 485 -870 486 -790
rect 835 -870 836 -790
rect 849 -791 850 -765
rect 856 -870 857 -790
rect 929 -791 930 -765
rect 1066 -791 1067 -765
rect 1094 -791 1095 -765
rect 1206 -870 1207 -790
rect 1248 -791 1249 -765
rect 1311 -870 1312 -790
rect 191 -870 192 -792
rect 548 -870 549 -792
rect 569 -870 570 -792
rect 1066 -870 1067 -792
rect 1080 -793 1081 -765
rect 1094 -870 1095 -792
rect 1199 -793 1200 -765
rect 1276 -870 1277 -792
rect 205 -795 206 -765
rect 765 -795 766 -765
rect 772 -870 773 -794
rect 807 -795 808 -765
rect 828 -870 829 -794
rect 1493 -870 1494 -794
rect 208 -797 209 -765
rect 1227 -870 1228 -796
rect 1248 -870 1249 -796
rect 1304 -797 1305 -765
rect 208 -870 209 -798
rect 723 -799 724 -765
rect 751 -799 752 -765
rect 1003 -870 1004 -798
rect 1027 -799 1028 -765
rect 1472 -870 1473 -798
rect 226 -801 227 -765
rect 310 -870 311 -800
rect 352 -870 353 -800
rect 506 -870 507 -800
rect 527 -801 528 -765
rect 1199 -870 1200 -800
rect 212 -803 213 -765
rect 226 -870 227 -802
rect 240 -803 241 -765
rect 289 -870 290 -802
rect 296 -870 297 -802
rect 492 -803 493 -765
rect 534 -870 535 -802
rect 758 -803 759 -765
rect 800 -803 801 -765
rect 1101 -870 1102 -802
rect 212 -870 213 -804
rect 436 -805 437 -765
rect 457 -870 458 -804
rect 527 -870 528 -804
rect 541 -805 542 -765
rect 1017 -870 1018 -804
rect 1045 -870 1046 -804
rect 1087 -805 1088 -765
rect 233 -807 234 -765
rect 436 -870 437 -806
rect 464 -870 465 -806
rect 471 -807 472 -765
rect 576 -807 577 -765
rect 765 -870 766 -806
rect 786 -807 787 -765
rect 800 -870 801 -806
rect 807 -870 808 -806
rect 863 -807 864 -765
rect 940 -807 941 -765
rect 947 -870 948 -806
rect 961 -870 962 -806
rect 1339 -807 1340 -765
rect 121 -809 122 -765
rect 786 -870 787 -808
rect 821 -809 822 -765
rect 940 -870 941 -808
rect 975 -809 976 -765
rect 1024 -870 1025 -808
rect 1059 -870 1060 -808
rect 1129 -809 1130 -765
rect 233 -870 234 -810
rect 411 -870 412 -810
rect 415 -811 416 -765
rect 523 -811 524 -765
rect 583 -811 584 -765
rect 611 -870 612 -810
rect 632 -870 633 -810
rect 667 -870 668 -810
rect 702 -811 703 -765
rect 723 -870 724 -810
rect 814 -811 815 -765
rect 821 -870 822 -810
rect 838 -811 839 -765
rect 1304 -870 1305 -810
rect 142 -813 143 -765
rect 523 -870 524 -812
rect 583 -870 584 -812
rect 681 -813 682 -765
rect 709 -813 710 -765
rect 758 -870 759 -812
rect 814 -870 815 -812
rect 1458 -870 1459 -812
rect 142 -870 143 -814
rect 891 -815 892 -765
rect 968 -815 969 -765
rect 975 -870 976 -814
rect 982 -815 983 -765
rect 989 -870 990 -814
rect 996 -815 997 -765
rect 1087 -870 1088 -814
rect 1122 -815 1123 -765
rect 1129 -870 1130 -814
rect 79 -817 80 -765
rect 891 -870 892 -816
rect 919 -817 920 -765
rect 996 -870 997 -816
rect 1073 -817 1074 -765
rect 1080 -870 1081 -816
rect 1122 -870 1123 -816
rect 1136 -817 1137 -765
rect 79 -870 80 -818
rect 86 -819 87 -765
rect 156 -870 157 -818
rect 681 -870 682 -818
rect 716 -870 717 -818
rect 964 -870 965 -818
rect 982 -870 983 -818
rect 1010 -819 1011 -765
rect 1052 -819 1053 -765
rect 1073 -870 1074 -818
rect 1136 -870 1137 -818
rect 1143 -819 1144 -765
rect 86 -870 87 -820
rect 100 -821 101 -765
rect 240 -870 241 -820
rect 387 -821 388 -765
rect 401 -821 402 -765
rect 576 -870 577 -820
rect 590 -821 591 -765
rect 849 -870 850 -820
rect 863 -870 864 -820
rect 884 -821 885 -765
rect 933 -821 934 -765
rect 1010 -870 1011 -820
rect 1031 -821 1032 -765
rect 1052 -870 1053 -820
rect 100 -870 101 -822
rect 443 -823 444 -765
rect 509 -870 510 -822
rect 1339 -870 1340 -822
rect 152 -870 153 -824
rect 443 -870 444 -824
rect 590 -870 591 -824
rect 639 -825 640 -765
rect 646 -870 647 -824
rect 1465 -825 1466 -765
rect 149 -827 150 -765
rect 639 -870 640 -826
rect 649 -827 650 -765
rect 1486 -870 1487 -826
rect 51 -870 52 -828
rect 149 -870 150 -828
rect 261 -829 262 -765
rect 324 -870 325 -828
rect 338 -829 339 -765
rect 387 -870 388 -828
rect 401 -870 402 -828
rect 422 -829 423 -765
rect 429 -829 430 -765
rect 719 -829 720 -765
rect 744 -829 745 -765
rect 884 -870 885 -828
rect 912 -829 913 -765
rect 933 -870 934 -828
rect 1381 -829 1382 -765
rect 1465 -870 1466 -828
rect 170 -831 171 -765
rect 338 -870 339 -830
rect 373 -831 374 -765
rect 492 -870 493 -830
rect 499 -831 500 -765
rect 744 -870 745 -830
rect 838 -870 839 -830
rect 1402 -831 1403 -765
rect 170 -870 171 -832
rect 198 -833 199 -765
rect 247 -833 248 -765
rect 261 -870 262 -832
rect 282 -833 283 -765
rect 394 -870 395 -832
rect 408 -833 409 -765
rect 562 -870 563 -832
rect 625 -833 626 -765
rect 968 -870 969 -832
rect 1283 -833 1284 -765
rect 1381 -870 1382 -832
rect 121 -870 122 -834
rect 282 -870 283 -834
rect 303 -835 304 -765
rect 415 -870 416 -834
rect 422 -870 423 -834
rect 873 -835 874 -765
rect 877 -870 878 -834
rect 1143 -870 1144 -834
rect 1269 -835 1270 -765
rect 1283 -870 1284 -834
rect 1360 -835 1361 -765
rect 1402 -870 1403 -834
rect 128 -837 129 -765
rect 247 -870 248 -836
rect 268 -837 269 -765
rect 303 -870 304 -836
rect 317 -837 318 -765
rect 429 -870 430 -836
rect 499 -870 500 -836
rect 1290 -870 1291 -836
rect 128 -870 129 -838
rect 177 -839 178 -765
rect 198 -870 199 -838
rect 205 -870 206 -838
rect 268 -870 269 -838
rect 831 -839 832 -765
rect 873 -870 874 -838
rect 1451 -839 1452 -765
rect 177 -870 178 -840
rect 275 -841 276 -765
rect 317 -870 318 -840
rect 450 -841 451 -765
rect 635 -841 636 -765
rect 709 -870 710 -840
rect 831 -870 832 -840
rect 1395 -841 1396 -765
rect 107 -843 108 -765
rect 450 -870 451 -842
rect 649 -870 650 -842
rect 702 -870 703 -842
rect 880 -870 881 -842
rect 1395 -870 1396 -842
rect 107 -870 108 -844
rect 1423 -870 1424 -844
rect 254 -870 255 -846
rect 275 -870 276 -846
rect 373 -870 374 -846
rect 730 -847 731 -765
rect 898 -847 899 -765
rect 912 -870 913 -846
rect 919 -870 920 -846
rect 1031 -870 1032 -846
rect 1164 -847 1165 -765
rect 1360 -870 1361 -846
rect 1388 -847 1389 -765
rect 1451 -870 1452 -846
rect 159 -849 160 -765
rect 898 -870 899 -848
rect 1185 -849 1186 -765
rect 1388 -870 1389 -848
rect 520 -851 521 -765
rect 1185 -870 1186 -850
rect 1234 -851 1235 -765
rect 1269 -870 1270 -850
rect 520 -870 521 -852
rect 541 -870 542 -852
rect 653 -853 654 -765
rect 730 -870 731 -852
rect 870 -853 871 -765
rect 1164 -870 1165 -852
rect 1234 -870 1235 -852
rect 1318 -853 1319 -765
rect 653 -870 654 -854
rect 674 -870 675 -854
rect 691 -855 692 -765
rect 1318 -870 1319 -854
rect 660 -857 661 -765
rect 688 -870 689 -856
rect 751 -870 752 -856
rect 870 -870 871 -856
rect 660 -870 661 -858
rect 695 -859 696 -765
rect 618 -861 619 -765
rect 695 -870 696 -860
rect 597 -863 598 -765
rect 618 -870 619 -862
rect 597 -870 598 -864
rect 842 -865 843 -765
rect 779 -867 780 -765
rect 842 -870 843 -866
rect 471 -870 472 -868
rect 779 -870 780 -868
rect 30 -997 31 -879
rect 142 -880 143 -878
rect 149 -880 150 -878
rect 891 -880 892 -878
rect 919 -880 920 -878
rect 1451 -880 1452 -878
rect 1458 -880 1459 -878
rect 1458 -997 1459 -879
rect 1458 -880 1459 -878
rect 1458 -997 1459 -879
rect 1500 -880 1501 -878
rect 1500 -997 1501 -879
rect 1500 -880 1501 -878
rect 1500 -997 1501 -879
rect 1542 -880 1543 -878
rect 1566 -997 1567 -879
rect 1570 -880 1571 -878
rect 1626 -997 1627 -879
rect 1724 -880 1725 -878
rect 1738 -997 1739 -879
rect 44 -882 45 -878
rect 628 -882 629 -878
rect 656 -997 657 -881
rect 1570 -997 1571 -881
rect 1577 -882 1578 -878
rect 1612 -997 1613 -881
rect 44 -997 45 -883
rect 51 -884 52 -878
rect 79 -884 80 -878
rect 649 -884 650 -878
rect 660 -884 661 -878
rect 831 -884 832 -878
rect 838 -884 839 -878
rect 870 -884 871 -878
rect 873 -884 874 -878
rect 1255 -884 1256 -878
rect 1318 -884 1319 -878
rect 1633 -997 1634 -883
rect 51 -997 52 -885
rect 65 -886 66 -878
rect 79 -997 80 -885
rect 128 -886 129 -878
rect 135 -886 136 -878
rect 142 -997 143 -885
rect 166 -886 167 -878
rect 1360 -886 1361 -878
rect 1521 -886 1522 -878
rect 1542 -997 1543 -885
rect 1573 -997 1574 -885
rect 1577 -997 1578 -885
rect 1584 -886 1585 -878
rect 1619 -997 1620 -885
rect 65 -997 66 -887
rect 72 -888 73 -878
rect 82 -997 83 -887
rect 233 -888 234 -878
rect 257 -888 258 -878
rect 1437 -888 1438 -878
rect 1479 -888 1480 -878
rect 1584 -997 1585 -887
rect 72 -997 73 -889
rect 86 -890 87 -878
rect 93 -890 94 -878
rect 152 -997 153 -889
rect 208 -890 209 -878
rect 352 -890 353 -878
rect 408 -890 409 -878
rect 551 -890 552 -878
rect 660 -997 661 -889
rect 856 -890 857 -878
rect 880 -890 881 -878
rect 1528 -890 1529 -878
rect 58 -892 59 -878
rect 86 -997 87 -891
rect 93 -997 94 -891
rect 569 -892 570 -878
rect 667 -892 668 -878
rect 940 -892 941 -878
rect 964 -892 965 -878
rect 1416 -892 1417 -878
rect 1437 -997 1438 -891
rect 1444 -892 1445 -878
rect 1479 -997 1480 -891
rect 1486 -892 1487 -878
rect 1493 -892 1494 -878
rect 1521 -997 1522 -891
rect 58 -997 59 -893
rect 422 -894 423 -878
rect 436 -894 437 -878
rect 642 -997 643 -893
rect 667 -997 668 -893
rect 688 -894 689 -878
rect 775 -997 776 -893
rect 1206 -894 1207 -878
rect 1346 -894 1347 -878
rect 1556 -894 1557 -878
rect 100 -896 101 -878
rect 964 -997 965 -895
rect 985 -997 986 -895
rect 1381 -896 1382 -878
rect 1388 -896 1389 -878
rect 1444 -997 1445 -895
rect 1465 -896 1466 -878
rect 1493 -997 1494 -895
rect 1514 -896 1515 -878
rect 1528 -997 1529 -895
rect 100 -997 101 -897
rect 877 -898 878 -878
rect 891 -997 892 -897
rect 954 -898 955 -878
rect 961 -997 962 -897
rect 1556 -997 1557 -897
rect 107 -900 108 -878
rect 296 -900 297 -878
rect 317 -900 318 -878
rect 320 -954 321 -899
rect 331 -900 332 -878
rect 331 -997 332 -899
rect 331 -900 332 -878
rect 331 -997 332 -899
rect 338 -900 339 -878
rect 499 -900 500 -878
rect 502 -900 503 -878
rect 968 -900 969 -878
rect 992 -997 993 -899
rect 1451 -997 1452 -899
rect 1465 -997 1466 -899
rect 1507 -900 1508 -878
rect 107 -997 108 -901
rect 212 -902 213 -878
rect 219 -997 220 -901
rect 534 -902 535 -878
rect 548 -902 549 -878
rect 590 -902 591 -878
rect 674 -902 675 -878
rect 884 -902 885 -878
rect 905 -902 906 -878
rect 919 -997 920 -901
rect 926 -902 927 -878
rect 929 -902 930 -878
rect 940 -997 941 -901
rect 1010 -902 1011 -878
rect 1069 -902 1070 -878
rect 1549 -902 1550 -878
rect 110 -904 111 -878
rect 310 -904 311 -878
rect 317 -997 318 -903
rect 352 -997 353 -903
rect 450 -904 451 -878
rect 502 -997 503 -903
rect 1423 -904 1424 -878
rect 1472 -904 1473 -878
rect 1514 -997 1515 -903
rect 1549 -997 1550 -903
rect 1563 -904 1564 -878
rect 121 -906 122 -878
rect 366 -906 367 -878
rect 408 -997 409 -905
rect 723 -906 724 -878
rect 779 -997 780 -905
rect 842 -906 843 -878
rect 856 -997 857 -905
rect 975 -906 976 -878
rect 1111 -997 1112 -905
rect 1486 -997 1487 -905
rect 1563 -997 1564 -905
rect 1605 -997 1606 -905
rect 121 -997 122 -907
rect 124 -908 125 -878
rect 128 -997 129 -907
rect 275 -908 276 -878
rect 289 -908 290 -878
rect 296 -997 297 -907
rect 310 -997 311 -907
rect 394 -908 395 -878
rect 411 -908 412 -878
rect 922 -908 923 -878
rect 926 -997 927 -907
rect 933 -908 934 -878
rect 968 -997 969 -907
rect 989 -908 990 -878
rect 1129 -908 1130 -878
rect 1129 -997 1130 -907
rect 1129 -908 1130 -878
rect 1129 -997 1130 -907
rect 1171 -908 1172 -878
rect 1206 -997 1207 -907
rect 1248 -908 1249 -878
rect 1381 -997 1382 -907
rect 1409 -908 1410 -878
rect 1416 -997 1417 -907
rect 138 -997 139 -909
rect 380 -910 381 -878
rect 394 -997 395 -909
rect 702 -910 703 -878
rect 723 -997 724 -909
rect 758 -910 759 -878
rect 782 -910 783 -878
rect 1395 -910 1396 -878
rect 163 -912 164 -878
rect 212 -997 213 -911
rect 222 -912 223 -878
rect 254 -912 255 -878
rect 268 -912 269 -878
rect 436 -997 437 -911
rect 446 -997 447 -911
rect 870 -997 871 -911
rect 877 -997 878 -911
rect 1192 -912 1193 -878
rect 1248 -997 1249 -911
rect 1262 -912 1263 -878
rect 1290 -912 1291 -878
rect 1346 -997 1347 -911
rect 1367 -912 1368 -878
rect 1409 -997 1410 -911
rect 163 -997 164 -913
rect 177 -914 178 -878
rect 191 -914 192 -878
rect 289 -997 290 -913
rect 380 -997 381 -913
rect 772 -914 773 -878
rect 828 -914 829 -878
rect 1360 -997 1361 -913
rect 1374 -914 1375 -878
rect 1507 -997 1508 -913
rect 177 -997 178 -915
rect 387 -916 388 -878
rect 450 -997 451 -915
rect 492 -916 493 -878
rect 506 -916 507 -878
rect 1017 -916 1018 -878
rect 1164 -916 1165 -878
rect 1192 -997 1193 -915
rect 1241 -916 1242 -878
rect 1262 -997 1263 -915
rect 1269 -916 1270 -878
rect 1290 -997 1291 -915
rect 1297 -916 1298 -878
rect 1367 -997 1368 -915
rect 1395 -997 1396 -915
rect 1430 -916 1431 -878
rect 191 -997 192 -917
rect 513 -918 514 -878
rect 520 -918 521 -878
rect 1318 -997 1319 -917
rect 135 -997 136 -919
rect 513 -997 514 -919
rect 523 -920 524 -878
rect 695 -920 696 -878
rect 698 -997 699 -919
rect 954 -997 955 -919
rect 975 -997 976 -919
rect 1255 -997 1256 -919
rect 1304 -920 1305 -878
rect 1388 -997 1389 -919
rect 198 -922 199 -878
rect 422 -997 423 -921
rect 425 -997 426 -921
rect 520 -997 521 -921
rect 530 -922 531 -878
rect 1024 -922 1025 -878
rect 1115 -922 1116 -878
rect 1297 -997 1298 -921
rect 198 -997 199 -923
rect 261 -924 262 -878
rect 268 -997 269 -923
rect 303 -924 304 -878
rect 387 -997 388 -923
rect 632 -924 633 -878
rect 670 -924 671 -878
rect 828 -997 829 -923
rect 845 -997 846 -923
rect 1374 -997 1375 -923
rect 205 -926 206 -878
rect 338 -997 339 -925
rect 492 -997 493 -925
rect 684 -926 685 -878
rect 688 -997 689 -925
rect 1311 -926 1312 -878
rect 205 -997 206 -927
rect 373 -928 374 -878
rect 509 -928 510 -878
rect 516 -954 517 -927
rect 534 -997 535 -927
rect 555 -928 556 -878
rect 569 -997 570 -927
rect 618 -928 619 -878
rect 625 -928 626 -878
rect 1423 -997 1424 -927
rect 184 -930 185 -878
rect 555 -997 556 -929
rect 586 -997 587 -929
rect 1115 -997 1116 -929
rect 1157 -930 1158 -878
rect 1164 -997 1165 -929
rect 1171 -997 1172 -929
rect 1178 -930 1179 -878
rect 1227 -930 1228 -878
rect 1269 -997 1270 -929
rect 1283 -930 1284 -878
rect 1304 -997 1305 -929
rect 149 -997 150 -931
rect 184 -997 185 -931
rect 226 -932 227 -878
rect 366 -997 367 -931
rect 373 -997 374 -931
rect 401 -932 402 -878
rect 506 -997 507 -931
rect 1283 -997 1284 -931
rect 233 -997 234 -933
rect 478 -934 479 -878
rect 509 -997 510 -933
rect 527 -934 528 -878
rect 590 -997 591 -933
rect 821 -934 822 -878
rect 898 -934 899 -878
rect 905 -997 906 -933
rect 933 -997 934 -933
rect 947 -934 948 -878
rect 999 -997 1000 -933
rect 1157 -997 1158 -933
rect 1234 -934 1235 -878
rect 1241 -997 1242 -933
rect 250 -997 251 -935
rect 548 -997 549 -935
rect 611 -936 612 -878
rect 632 -997 633 -935
rect 674 -997 675 -935
rect 730 -936 731 -878
rect 758 -997 759 -935
rect 786 -936 787 -878
rect 898 -997 899 -935
rect 1353 -936 1354 -878
rect 254 -997 255 -937
rect 282 -938 283 -878
rect 303 -997 304 -937
rect 415 -938 416 -878
rect 478 -997 479 -937
rect 485 -938 486 -878
rect 527 -997 528 -937
rect 814 -938 815 -878
rect 835 -938 836 -878
rect 1353 -997 1354 -937
rect 170 -940 171 -878
rect 282 -997 283 -939
rect 401 -997 402 -939
rect 429 -940 430 -878
rect 485 -997 486 -939
rect 653 -940 654 -878
rect 677 -940 678 -878
rect 1325 -940 1326 -878
rect 156 -942 157 -878
rect 170 -997 171 -941
rect 261 -997 262 -941
rect 345 -942 346 -878
rect 415 -997 416 -941
rect 541 -942 542 -878
rect 604 -942 605 -878
rect 611 -997 612 -941
rect 625 -997 626 -941
rect 649 -997 650 -941
rect 684 -997 685 -941
rect 786 -997 787 -941
rect 800 -942 801 -878
rect 814 -997 815 -941
rect 901 -997 902 -941
rect 1311 -997 1312 -941
rect 1325 -997 1326 -941
rect 1339 -942 1340 -878
rect 156 -997 157 -943
rect 247 -944 248 -878
rect 275 -997 276 -943
rect 471 -944 472 -878
rect 541 -997 542 -943
rect 562 -944 563 -878
rect 695 -997 696 -943
rect 744 -944 745 -878
rect 768 -997 769 -943
rect 1339 -997 1340 -943
rect 345 -997 346 -945
rect 359 -946 360 -878
rect 429 -997 430 -945
rect 576 -946 577 -878
rect 597 -946 598 -878
rect 744 -997 745 -945
rect 772 -997 773 -945
rect 1591 -997 1592 -945
rect 114 -948 115 -878
rect 359 -997 360 -947
rect 457 -948 458 -878
rect 604 -997 605 -947
rect 702 -997 703 -947
rect 751 -948 752 -878
rect 793 -948 794 -878
rect 800 -997 801 -947
rect 1017 -997 1018 -947
rect 1038 -948 1039 -878
rect 1150 -948 1151 -878
rect 1178 -997 1179 -947
rect 1220 -948 1221 -878
rect 1234 -997 1235 -947
rect 114 -997 115 -949
rect 240 -950 241 -878
rect 443 -950 444 -878
rect 457 -997 458 -949
rect 464 -950 465 -878
rect 471 -997 472 -949
rect 562 -997 563 -949
rect 765 -950 766 -878
rect 793 -997 794 -949
rect 807 -950 808 -878
rect 1024 -997 1025 -949
rect 1052 -950 1053 -878
rect 1108 -950 1109 -878
rect 1220 -997 1221 -949
rect 37 -952 38 -878
rect 240 -997 241 -951
rect 443 -997 444 -951
rect 1472 -997 1473 -951
rect 37 -997 38 -953
rect 863 -954 864 -878
rect 929 -997 930 -953
rect 947 -997 948 -953
rect 1038 -997 1039 -953
rect 1094 -954 1095 -878
rect 1150 -997 1151 -953
rect 1332 -954 1333 -878
rect 464 -997 465 -955
rect 1010 -997 1011 -955
rect 1052 -997 1053 -955
rect 1101 -956 1102 -878
rect 1332 -997 1333 -955
rect 1402 -956 1403 -878
rect 576 -997 577 -957
rect 737 -958 738 -878
rect 765 -997 766 -957
rect 1598 -997 1599 -957
rect 583 -960 584 -878
rect 751 -997 752 -959
rect 842 -997 843 -959
rect 1402 -997 1403 -959
rect 583 -997 584 -961
rect 849 -962 850 -878
rect 1059 -962 1060 -878
rect 1101 -997 1102 -961
rect 597 -997 598 -963
rect 1003 -964 1004 -878
rect 1031 -964 1032 -878
rect 1059 -997 1060 -963
rect 1094 -997 1095 -963
rect 1185 -964 1186 -878
rect 639 -966 640 -878
rect 1185 -997 1186 -965
rect 639 -997 640 -967
rect 1430 -997 1431 -967
rect 646 -970 647 -878
rect 863 -997 864 -969
rect 982 -970 983 -878
rect 1003 -997 1004 -969
rect 1031 -997 1032 -969
rect 1073 -970 1074 -878
rect 646 -997 647 -971
rect 1276 -972 1277 -878
rect 716 -974 717 -878
rect 821 -997 822 -973
rect 849 -997 850 -973
rect 912 -974 913 -878
rect 978 -997 979 -973
rect 1276 -997 1277 -973
rect 681 -976 682 -878
rect 912 -997 913 -975
rect 982 -997 983 -975
rect 1213 -976 1214 -878
rect 226 -997 227 -977
rect 681 -997 682 -977
rect 709 -978 710 -878
rect 716 -997 717 -977
rect 730 -997 731 -977
rect 1227 -997 1228 -977
rect 499 -997 500 -979
rect 709 -997 710 -979
rect 733 -997 734 -979
rect 835 -997 836 -979
rect 1073 -997 1074 -979
rect 1080 -980 1081 -878
rect 1199 -980 1200 -878
rect 1213 -997 1214 -979
rect 737 -997 738 -981
rect 996 -982 997 -878
rect 1045 -982 1046 -878
rect 1199 -997 1200 -981
rect 996 -997 997 -983
rect 1535 -984 1536 -878
rect 653 -997 654 -985
rect 1535 -997 1536 -985
rect 1045 -997 1046 -987
rect 1143 -988 1144 -878
rect 1080 -997 1081 -989
rect 1087 -990 1088 -878
rect 1136 -990 1137 -878
rect 1143 -997 1144 -989
rect 884 -997 885 -991
rect 1087 -997 1088 -991
rect 1122 -992 1123 -878
rect 1136 -997 1137 -991
rect 1066 -994 1067 -878
rect 1122 -997 1123 -993
rect 537 -996 538 -878
rect 1066 -997 1067 -995
rect 23 -1098 24 -1006
rect 618 -1007 619 -1005
rect 628 -1098 629 -1006
rect 723 -1007 724 -1005
rect 751 -1007 752 -1005
rect 751 -1098 752 -1006
rect 751 -1007 752 -1005
rect 751 -1098 752 -1006
rect 768 -1007 769 -1005
rect 940 -1007 941 -1005
rect 961 -1007 962 -1005
rect 1332 -1007 1333 -1005
rect 1339 -1007 1340 -1005
rect 1339 -1098 1340 -1006
rect 1339 -1007 1340 -1005
rect 1339 -1098 1340 -1006
rect 1374 -1007 1375 -1005
rect 1566 -1007 1567 -1005
rect 1570 -1007 1571 -1005
rect 1675 -1098 1676 -1006
rect 1738 -1007 1739 -1005
rect 1745 -1098 1746 -1006
rect 30 -1009 31 -1005
rect 135 -1098 136 -1008
rect 149 -1098 150 -1008
rect 205 -1009 206 -1005
rect 250 -1009 251 -1005
rect 296 -1009 297 -1005
rect 310 -1009 311 -1005
rect 516 -1098 517 -1008
rect 555 -1009 556 -1005
rect 723 -1098 724 -1008
rect 786 -1009 787 -1005
rect 901 -1009 902 -1005
rect 919 -1009 920 -1005
rect 1384 -1098 1385 -1008
rect 1528 -1009 1529 -1005
rect 1570 -1098 1571 -1008
rect 1591 -1009 1592 -1005
rect 1682 -1098 1683 -1008
rect 30 -1098 31 -1010
rect 597 -1011 598 -1005
rect 611 -1011 612 -1005
rect 656 -1011 657 -1005
rect 667 -1011 668 -1005
rect 730 -1011 731 -1005
rect 786 -1098 787 -1010
rect 800 -1011 801 -1005
rect 845 -1011 846 -1005
rect 1199 -1011 1200 -1005
rect 1241 -1011 1242 -1005
rect 1374 -1098 1375 -1010
rect 1486 -1011 1487 -1005
rect 1528 -1098 1529 -1010
rect 1535 -1011 1536 -1005
rect 1640 -1098 1641 -1010
rect 37 -1013 38 -1005
rect 695 -1013 696 -1005
rect 698 -1013 699 -1005
rect 1591 -1098 1592 -1012
rect 1626 -1013 1627 -1005
rect 1654 -1098 1655 -1012
rect 44 -1015 45 -1005
rect 75 -1098 76 -1014
rect 82 -1015 83 -1005
rect 107 -1015 108 -1005
rect 114 -1015 115 -1005
rect 215 -1098 216 -1014
rect 275 -1015 276 -1005
rect 999 -1015 1000 -1005
rect 1010 -1015 1011 -1005
rect 1521 -1015 1522 -1005
rect 1552 -1015 1553 -1005
rect 1612 -1015 1613 -1005
rect 1633 -1015 1634 -1005
rect 1633 -1098 1634 -1014
rect 1633 -1015 1634 -1005
rect 1633 -1098 1634 -1014
rect 44 -1098 45 -1016
rect 86 -1017 87 -1005
rect 89 -1098 90 -1016
rect 408 -1017 409 -1005
rect 422 -1017 423 -1005
rect 1605 -1017 1606 -1005
rect 58 -1019 59 -1005
rect 61 -1077 62 -1018
rect 72 -1019 73 -1005
rect 86 -1098 87 -1018
rect 100 -1019 101 -1005
rect 425 -1019 426 -1005
rect 485 -1019 486 -1005
rect 611 -1098 612 -1018
rect 618 -1098 619 -1018
rect 632 -1019 633 -1005
rect 684 -1019 685 -1005
rect 1220 -1019 1221 -1005
rect 1241 -1098 1242 -1018
rect 1297 -1019 1298 -1005
rect 1360 -1019 1361 -1005
rect 1486 -1098 1487 -1018
rect 1500 -1019 1501 -1005
rect 1535 -1098 1536 -1018
rect 1556 -1019 1557 -1005
rect 1612 -1098 1613 -1018
rect 51 -1021 52 -1005
rect 72 -1098 73 -1020
rect 100 -1098 101 -1020
rect 436 -1021 437 -1005
rect 492 -1021 493 -1005
rect 775 -1021 776 -1005
rect 800 -1098 801 -1020
rect 1248 -1021 1249 -1005
rect 1269 -1021 1270 -1005
rect 1269 -1098 1270 -1020
rect 1269 -1021 1270 -1005
rect 1269 -1098 1270 -1020
rect 1297 -1098 1298 -1020
rect 1311 -1021 1312 -1005
rect 1395 -1021 1396 -1005
rect 1500 -1098 1501 -1020
rect 1563 -1021 1564 -1005
rect 1647 -1098 1648 -1020
rect 51 -1098 52 -1022
rect 121 -1023 122 -1005
rect 128 -1023 129 -1005
rect 236 -1098 237 -1022
rect 268 -1023 269 -1005
rect 408 -1098 409 -1022
rect 492 -1098 493 -1022
rect 992 -1023 993 -1005
rect 996 -1023 997 -1005
rect 1325 -1023 1326 -1005
rect 1381 -1023 1382 -1005
rect 1395 -1098 1396 -1022
rect 1423 -1023 1424 -1005
rect 1521 -1098 1522 -1022
rect 1577 -1023 1578 -1005
rect 1626 -1098 1627 -1022
rect 58 -1098 59 -1024
rect 107 -1098 108 -1024
rect 481 -1098 482 -1024
rect 499 -1025 500 -1005
rect 604 -1025 605 -1005
rect 632 -1098 633 -1024
rect 702 -1025 703 -1005
rect 730 -1098 731 -1024
rect 758 -1025 759 -1005
rect 835 -1025 836 -1005
rect 996 -1098 997 -1024
rect 1003 -1025 1004 -1005
rect 1010 -1098 1011 -1024
rect 1013 -1025 1014 -1005
rect 1031 -1025 1032 -1005
rect 1108 -1025 1109 -1005
rect 1556 -1098 1557 -1024
rect 1584 -1025 1585 -1005
rect 1605 -1098 1606 -1024
rect 114 -1098 115 -1026
rect 212 -1027 213 -1005
rect 275 -1098 276 -1026
rect 842 -1027 843 -1005
rect 849 -1027 850 -1005
rect 849 -1098 850 -1026
rect 849 -1027 850 -1005
rect 849 -1098 850 -1026
rect 856 -1027 857 -1005
rect 919 -1098 920 -1026
rect 933 -1027 934 -1005
rect 961 -1098 962 -1026
rect 975 -1098 976 -1026
rect 1066 -1027 1067 -1005
rect 1111 -1027 1112 -1005
rect 1493 -1027 1494 -1005
rect 1507 -1027 1508 -1005
rect 1584 -1098 1585 -1026
rect 121 -1098 122 -1028
rect 317 -1029 318 -1005
rect 324 -1029 325 -1005
rect 509 -1029 510 -1005
rect 520 -1029 521 -1005
rect 702 -1098 703 -1028
rect 733 -1029 734 -1005
rect 1360 -1098 1361 -1028
rect 1409 -1029 1410 -1005
rect 1423 -1098 1424 -1028
rect 1430 -1029 1431 -1005
rect 1507 -1098 1508 -1028
rect 1542 -1029 1543 -1005
rect 1577 -1098 1578 -1028
rect 128 -1098 129 -1030
rect 233 -1031 234 -1005
rect 282 -1031 283 -1005
rect 443 -1031 444 -1005
rect 541 -1031 542 -1005
rect 667 -1098 668 -1030
rect 688 -1098 689 -1030
rect 1185 -1031 1186 -1005
rect 1220 -1098 1221 -1030
rect 1255 -1031 1256 -1005
rect 1318 -1031 1319 -1005
rect 1325 -1098 1326 -1030
rect 1409 -1098 1410 -1030
rect 1437 -1031 1438 -1005
rect 1444 -1031 1445 -1005
rect 1563 -1098 1564 -1030
rect 138 -1033 139 -1005
rect 485 -1098 486 -1032
rect 506 -1033 507 -1005
rect 1318 -1098 1319 -1032
rect 1416 -1033 1417 -1005
rect 1437 -1098 1438 -1032
rect 1444 -1098 1445 -1032
rect 1451 -1033 1452 -1005
rect 138 -1098 139 -1034
rect 1472 -1035 1473 -1005
rect 156 -1037 157 -1005
rect 317 -1098 318 -1036
rect 331 -1037 332 -1005
rect 502 -1037 503 -1005
rect 541 -1098 542 -1036
rect 569 -1037 570 -1005
rect 576 -1037 577 -1005
rect 695 -1098 696 -1036
rect 737 -1037 738 -1005
rect 842 -1098 843 -1036
rect 863 -1037 864 -1005
rect 887 -1037 888 -1005
rect 891 -1037 892 -1005
rect 940 -1098 941 -1036
rect 954 -1037 955 -1005
rect 1031 -1098 1032 -1036
rect 1066 -1098 1067 -1036
rect 1101 -1037 1102 -1005
rect 1115 -1037 1116 -1005
rect 1332 -1098 1333 -1036
rect 1402 -1037 1403 -1005
rect 1416 -1098 1417 -1036
rect 1472 -1098 1473 -1036
rect 1619 -1037 1620 -1005
rect 156 -1098 157 -1038
rect 387 -1039 388 -1005
rect 394 -1039 395 -1005
rect 520 -1098 521 -1038
rect 548 -1039 549 -1005
rect 555 -1098 556 -1038
rect 562 -1039 563 -1005
rect 604 -1098 605 -1038
rect 660 -1039 661 -1005
rect 758 -1098 759 -1038
rect 793 -1039 794 -1005
rect 835 -1098 836 -1038
rect 866 -1098 867 -1038
rect 1150 -1039 1151 -1005
rect 1157 -1039 1158 -1005
rect 1311 -1098 1312 -1038
rect 1388 -1039 1389 -1005
rect 1402 -1098 1403 -1038
rect 1598 -1039 1599 -1005
rect 1619 -1098 1620 -1038
rect 170 -1041 171 -1005
rect 173 -1077 174 -1040
rect 177 -1041 178 -1005
rect 268 -1098 269 -1040
rect 296 -1098 297 -1040
rect 880 -1098 881 -1040
rect 891 -1098 892 -1040
rect 1115 -1098 1116 -1040
rect 1129 -1041 1130 -1005
rect 1132 -1041 1133 -1005
rect 1157 -1098 1158 -1040
rect 1381 -1098 1382 -1040
rect 1388 -1098 1389 -1040
rect 1475 -1098 1476 -1040
rect 170 -1098 171 -1042
rect 310 -1098 311 -1042
rect 397 -1098 398 -1042
rect 401 -1043 402 -1005
rect 436 -1098 437 -1042
rect 457 -1043 458 -1005
rect 506 -1098 507 -1042
rect 548 -1098 549 -1042
rect 677 -1098 678 -1042
rect 691 -1043 692 -1005
rect 772 -1098 773 -1042
rect 894 -1098 895 -1042
rect 1080 -1043 1081 -1005
rect 1090 -1098 1091 -1042
rect 1430 -1098 1431 -1042
rect 177 -1098 178 -1044
rect 212 -1098 213 -1044
rect 219 -1045 220 -1005
rect 282 -1098 283 -1044
rect 331 -1098 332 -1044
rect 450 -1045 451 -1005
rect 457 -1098 458 -1044
rect 471 -1045 472 -1005
rect 562 -1098 563 -1044
rect 1493 -1098 1494 -1044
rect 184 -1047 185 -1005
rect 205 -1098 206 -1046
rect 219 -1098 220 -1046
rect 534 -1047 535 -1005
rect 569 -1098 570 -1046
rect 674 -1047 675 -1005
rect 716 -1047 717 -1005
rect 737 -1098 738 -1046
rect 870 -1047 871 -1005
rect 1080 -1098 1081 -1046
rect 1129 -1098 1130 -1046
rect 1164 -1047 1165 -1005
rect 1185 -1098 1186 -1046
rect 1206 -1047 1207 -1005
rect 1234 -1047 1235 -1005
rect 1248 -1098 1249 -1046
rect 1255 -1098 1256 -1046
rect 1304 -1047 1305 -1005
rect 142 -1049 143 -1005
rect 184 -1098 185 -1048
rect 191 -1049 192 -1005
rect 646 -1049 647 -1005
rect 660 -1098 661 -1048
rect 803 -1098 804 -1048
rect 821 -1049 822 -1005
rect 870 -1098 871 -1048
rect 877 -1049 878 -1005
rect 1304 -1098 1305 -1048
rect 142 -1098 143 -1050
rect 646 -1098 647 -1050
rect 733 -1098 734 -1050
rect 1598 -1098 1599 -1050
rect 191 -1098 192 -1052
rect 254 -1053 255 -1005
rect 338 -1053 339 -1005
rect 387 -1098 388 -1052
rect 394 -1098 395 -1052
rect 1353 -1053 1354 -1005
rect 198 -1055 199 -1005
rect 324 -1098 325 -1054
rect 345 -1055 346 -1005
rect 345 -1098 346 -1054
rect 345 -1055 346 -1005
rect 345 -1098 346 -1054
rect 352 -1055 353 -1005
rect 621 -1055 622 -1005
rect 625 -1055 626 -1005
rect 716 -1098 717 -1054
rect 744 -1055 745 -1005
rect 821 -1098 822 -1054
rect 877 -1098 878 -1054
rect 1199 -1098 1200 -1054
rect 1206 -1098 1207 -1054
rect 1549 -1055 1550 -1005
rect 163 -1057 164 -1005
rect 198 -1098 199 -1056
rect 254 -1098 255 -1056
rect 415 -1057 416 -1005
rect 446 -1057 447 -1005
rect 625 -1098 626 -1056
rect 744 -1098 745 -1056
rect 779 -1057 780 -1005
rect 912 -1057 913 -1005
rect 1542 -1098 1543 -1056
rect 163 -1098 164 -1058
rect 380 -1059 381 -1005
rect 401 -1098 402 -1058
rect 590 -1059 591 -1005
rect 597 -1098 598 -1058
rect 1055 -1098 1056 -1058
rect 1073 -1059 1074 -1005
rect 1101 -1098 1102 -1058
rect 1227 -1059 1228 -1005
rect 1234 -1098 1235 -1058
rect 1353 -1098 1354 -1058
rect 1367 -1059 1368 -1005
rect 1465 -1059 1466 -1005
rect 1549 -1098 1550 -1058
rect 261 -1061 262 -1005
rect 352 -1098 353 -1060
rect 359 -1061 360 -1005
rect 415 -1098 416 -1060
rect 450 -1098 451 -1060
rect 649 -1061 650 -1005
rect 653 -1061 654 -1005
rect 779 -1098 780 -1060
rect 926 -1061 927 -1005
rect 954 -1098 955 -1060
rect 982 -1061 983 -1005
rect 1108 -1098 1109 -1060
rect 1213 -1061 1214 -1005
rect 1227 -1098 1228 -1060
rect 1346 -1061 1347 -1005
rect 1367 -1098 1368 -1060
rect 1465 -1098 1466 -1060
rect 1479 -1061 1480 -1005
rect 359 -1098 360 -1062
rect 887 -1098 888 -1062
rect 905 -1063 906 -1005
rect 982 -1098 983 -1062
rect 985 -1063 986 -1005
rect 1514 -1063 1515 -1005
rect 366 -1065 367 -1005
rect 366 -1098 367 -1064
rect 366 -1065 367 -1005
rect 366 -1098 367 -1064
rect 373 -1065 374 -1005
rect 443 -1098 444 -1064
rect 464 -1065 465 -1005
rect 590 -1098 591 -1064
rect 649 -1098 650 -1064
rect 926 -1098 927 -1064
rect 933 -1098 934 -1064
rect 1017 -1065 1018 -1005
rect 1024 -1065 1025 -1005
rect 1027 -1065 1028 -1005
rect 1073 -1098 1074 -1064
rect 1136 -1065 1137 -1005
rect 1171 -1065 1172 -1005
rect 1213 -1098 1214 -1064
rect 1458 -1065 1459 -1005
rect 1514 -1098 1515 -1064
rect 226 -1067 227 -1005
rect 373 -1098 374 -1066
rect 380 -1098 381 -1066
rect 429 -1067 430 -1005
rect 471 -1098 472 -1066
rect 912 -1098 913 -1066
rect 968 -1067 969 -1005
rect 1017 -1098 1018 -1066
rect 1024 -1098 1025 -1066
rect 1038 -1067 1039 -1005
rect 1136 -1098 1137 -1066
rect 1178 -1067 1179 -1005
rect 226 -1098 227 -1068
rect 303 -1069 304 -1005
rect 429 -1098 430 -1068
rect 478 -1069 479 -1005
rect 534 -1098 535 -1068
rect 698 -1098 699 -1068
rect 863 -1098 864 -1068
rect 1479 -1098 1480 -1068
rect 289 -1071 290 -1005
rect 464 -1098 465 -1070
rect 576 -1098 577 -1070
rect 1451 -1098 1452 -1070
rect 289 -1098 290 -1072
rect 527 -1073 528 -1005
rect 583 -1073 584 -1005
rect 856 -1098 857 -1072
rect 905 -1098 906 -1072
rect 1003 -1098 1004 -1072
rect 1122 -1073 1123 -1005
rect 1178 -1098 1179 -1072
rect 250 -1098 251 -1074
rect 527 -1098 528 -1074
rect 586 -1075 587 -1005
rect 793 -1098 794 -1074
rect 947 -1075 948 -1005
rect 968 -1098 969 -1074
rect 989 -1075 990 -1005
rect 1262 -1075 1263 -1005
rect 303 -1098 304 -1076
rect 765 -1077 766 -1005
rect 947 -1098 948 -1076
rect 1052 -1077 1053 -1005
rect 1132 -1098 1133 -1076
rect 1164 -1098 1165 -1076
rect 1171 -1098 1172 -1076
rect 1192 -1077 1193 -1005
rect 1262 -1098 1263 -1076
rect 1290 -1077 1291 -1005
rect 131 -1079 132 -1005
rect 765 -1098 766 -1078
rect 1045 -1079 1046 -1005
rect 1122 -1098 1123 -1078
rect 1143 -1079 1144 -1005
rect 1192 -1098 1193 -1078
rect 1283 -1079 1284 -1005
rect 1290 -1098 1291 -1078
rect 338 -1098 339 -1080
rect 989 -1098 990 -1080
rect 1045 -1098 1046 -1080
rect 1059 -1081 1060 -1005
rect 1094 -1081 1095 -1005
rect 1143 -1098 1144 -1080
rect 1276 -1081 1277 -1005
rect 1283 -1098 1284 -1080
rect 513 -1083 514 -1005
rect 583 -1098 584 -1082
rect 642 -1098 643 -1082
rect 1458 -1098 1459 -1082
rect 513 -1098 514 -1084
rect 681 -1085 682 -1005
rect 828 -1085 829 -1005
rect 1094 -1098 1095 -1084
rect 79 -1087 80 -1005
rect 681 -1098 682 -1086
rect 814 -1087 815 -1005
rect 828 -1098 829 -1086
rect 978 -1087 979 -1005
rect 1059 -1098 1060 -1086
rect 79 -1098 80 -1088
rect 93 -1089 94 -1005
rect 653 -1098 654 -1088
rect 709 -1089 710 -1005
rect 807 -1089 808 -1005
rect 814 -1098 815 -1088
rect 1006 -1098 1007 -1088
rect 1276 -1098 1277 -1088
rect 93 -1098 94 -1090
rect 639 -1091 640 -1005
rect 674 -1098 675 -1090
rect 1346 -1098 1347 -1090
rect 499 -1098 500 -1092
rect 639 -1098 640 -1092
rect 709 -1098 710 -1092
rect 898 -1093 899 -1005
rect 807 -1098 808 -1094
rect 884 -1098 885 -1094
rect 898 -1098 899 -1094
rect 1087 -1095 1088 -1005
rect 1087 -1098 1088 -1096
rect 1150 -1098 1151 -1096
rect 23 -1108 24 -1106
rect 439 -1217 440 -1107
rect 471 -1108 472 -1106
rect 702 -1108 703 -1106
rect 730 -1108 731 -1106
rect 1241 -1108 1242 -1106
rect 1255 -1108 1256 -1106
rect 1381 -1108 1382 -1106
rect 1384 -1108 1385 -1106
rect 1626 -1108 1627 -1106
rect 1640 -1108 1641 -1106
rect 1724 -1217 1725 -1107
rect 1745 -1108 1746 -1106
rect 1759 -1217 1760 -1107
rect 23 -1217 24 -1109
rect 243 -1217 244 -1109
rect 275 -1110 276 -1106
rect 478 -1217 479 -1109
rect 499 -1110 500 -1106
rect 625 -1110 626 -1106
rect 649 -1110 650 -1106
rect 744 -1110 745 -1106
rect 765 -1110 766 -1106
rect 866 -1110 867 -1106
rect 887 -1110 888 -1106
rect 1374 -1110 1375 -1106
rect 1423 -1110 1424 -1106
rect 1423 -1217 1424 -1109
rect 1423 -1110 1424 -1106
rect 1423 -1217 1424 -1109
rect 1444 -1110 1445 -1106
rect 1661 -1217 1662 -1109
rect 1675 -1110 1676 -1106
rect 1703 -1217 1704 -1109
rect 37 -1217 38 -1111
rect 212 -1112 213 -1106
rect 219 -1112 220 -1106
rect 250 -1112 251 -1106
rect 275 -1217 276 -1111
rect 303 -1112 304 -1106
rect 324 -1112 325 -1106
rect 341 -1112 342 -1106
rect 366 -1112 367 -1106
rect 366 -1217 367 -1111
rect 366 -1112 367 -1106
rect 366 -1217 367 -1111
rect 401 -1112 402 -1106
rect 677 -1112 678 -1106
rect 681 -1112 682 -1106
rect 800 -1217 801 -1111
rect 817 -1217 818 -1111
rect 1185 -1112 1186 -1106
rect 1213 -1112 1214 -1106
rect 1381 -1217 1382 -1111
rect 1444 -1217 1445 -1111
rect 1766 -1217 1767 -1111
rect 72 -1217 73 -1113
rect 541 -1114 542 -1106
rect 656 -1217 657 -1113
rect 1346 -1114 1347 -1106
rect 1451 -1114 1452 -1106
rect 1563 -1114 1564 -1106
rect 1570 -1114 1571 -1106
rect 1717 -1217 1718 -1113
rect 75 -1116 76 -1106
rect 1675 -1217 1676 -1115
rect 1682 -1116 1683 -1106
rect 1769 -1217 1770 -1115
rect 89 -1118 90 -1106
rect 513 -1217 514 -1117
rect 516 -1118 517 -1106
rect 597 -1118 598 -1106
rect 681 -1217 682 -1117
rect 772 -1118 773 -1106
rect 835 -1118 836 -1106
rect 877 -1118 878 -1106
rect 929 -1217 930 -1117
rect 1297 -1118 1298 -1106
rect 1318 -1118 1319 -1106
rect 1451 -1217 1452 -1117
rect 1465 -1118 1466 -1106
rect 1682 -1217 1683 -1117
rect 93 -1120 94 -1106
rect 544 -1217 545 -1119
rect 548 -1120 549 -1106
rect 877 -1217 878 -1119
rect 933 -1120 934 -1106
rect 1374 -1217 1375 -1119
rect 1437 -1120 1438 -1106
rect 1563 -1217 1564 -1119
rect 1570 -1217 1571 -1119
rect 1605 -1120 1606 -1106
rect 1612 -1120 1613 -1106
rect 1752 -1217 1753 -1119
rect 93 -1217 94 -1121
rect 138 -1122 139 -1106
rect 173 -1217 174 -1121
rect 667 -1122 668 -1106
rect 688 -1122 689 -1106
rect 824 -1217 825 -1121
rect 859 -1217 860 -1121
rect 898 -1122 899 -1106
rect 912 -1122 913 -1106
rect 933 -1217 934 -1121
rect 950 -1217 951 -1121
rect 1304 -1122 1305 -1106
rect 1311 -1122 1312 -1106
rect 1437 -1217 1438 -1121
rect 1479 -1122 1480 -1106
rect 1605 -1217 1606 -1121
rect 1654 -1122 1655 -1106
rect 1780 -1217 1781 -1121
rect 100 -1124 101 -1106
rect 422 -1217 423 -1123
rect 506 -1124 507 -1106
rect 730 -1217 731 -1123
rect 737 -1124 738 -1106
rect 744 -1217 745 -1123
rect 758 -1124 759 -1106
rect 912 -1217 913 -1123
rect 1045 -1124 1046 -1106
rect 1234 -1124 1235 -1106
rect 1248 -1124 1249 -1106
rect 1612 -1217 1613 -1123
rect 58 -1126 59 -1106
rect 100 -1217 101 -1125
rect 107 -1126 108 -1106
rect 233 -1126 234 -1106
rect 236 -1126 237 -1106
rect 1472 -1217 1473 -1125
rect 1493 -1126 1494 -1106
rect 1619 -1126 1620 -1106
rect 58 -1217 59 -1127
rect 170 -1128 171 -1106
rect 177 -1128 178 -1106
rect 625 -1217 626 -1127
rect 653 -1128 654 -1106
rect 772 -1217 773 -1127
rect 891 -1128 892 -1106
rect 1311 -1217 1312 -1127
rect 1332 -1128 1333 -1106
rect 1454 -1128 1455 -1106
rect 1496 -1128 1497 -1106
rect 1647 -1128 1648 -1106
rect 68 -1217 69 -1129
rect 1248 -1217 1249 -1129
rect 1290 -1130 1291 -1106
rect 1619 -1217 1620 -1129
rect 89 -1217 90 -1131
rect 1493 -1217 1494 -1131
rect 1500 -1132 1501 -1106
rect 1640 -1217 1641 -1131
rect 110 -1217 111 -1133
rect 324 -1217 325 -1133
rect 380 -1134 381 -1106
rect 548 -1217 549 -1133
rect 698 -1134 699 -1106
rect 786 -1134 787 -1106
rect 891 -1217 892 -1133
rect 1290 -1217 1291 -1133
rect 1325 -1134 1326 -1106
rect 1500 -1217 1501 -1133
rect 1507 -1134 1508 -1106
rect 1647 -1217 1648 -1133
rect 114 -1136 115 -1106
rect 114 -1217 115 -1135
rect 114 -1136 115 -1106
rect 114 -1217 115 -1135
rect 121 -1136 122 -1106
rect 397 -1136 398 -1106
rect 401 -1217 402 -1135
rect 408 -1136 409 -1106
rect 415 -1136 416 -1106
rect 635 -1217 636 -1135
rect 716 -1136 717 -1106
rect 1213 -1217 1214 -1135
rect 1220 -1136 1221 -1106
rect 1710 -1217 1711 -1135
rect 121 -1217 122 -1137
rect 1626 -1217 1627 -1137
rect 128 -1140 129 -1106
rect 135 -1217 136 -1139
rect 180 -1217 181 -1139
rect 310 -1140 311 -1106
rect 380 -1217 381 -1139
rect 569 -1140 570 -1106
rect 649 -1217 650 -1139
rect 1220 -1217 1221 -1139
rect 1325 -1217 1326 -1139
rect 1430 -1140 1431 -1106
rect 1514 -1140 1515 -1106
rect 1668 -1217 1669 -1139
rect 128 -1217 129 -1141
rect 229 -1217 230 -1141
rect 233 -1217 234 -1141
rect 429 -1142 430 -1106
rect 485 -1142 486 -1106
rect 786 -1217 787 -1141
rect 919 -1142 920 -1106
rect 1045 -1217 1046 -1141
rect 1048 -1142 1049 -1106
rect 1199 -1142 1200 -1106
rect 1339 -1142 1340 -1106
rect 1507 -1217 1508 -1141
rect 1528 -1142 1529 -1106
rect 1689 -1217 1690 -1141
rect 184 -1144 185 -1106
rect 303 -1217 304 -1143
rect 387 -1144 388 -1106
rect 408 -1217 409 -1143
rect 415 -1217 416 -1143
rect 450 -1144 451 -1106
rect 492 -1144 493 -1106
rect 716 -1217 717 -1143
rect 723 -1144 724 -1106
rect 835 -1217 836 -1143
rect 968 -1144 969 -1106
rect 1332 -1217 1333 -1143
rect 1367 -1144 1368 -1106
rect 1514 -1217 1515 -1143
rect 1549 -1144 1550 -1106
rect 1696 -1217 1697 -1143
rect 79 -1146 80 -1106
rect 387 -1217 388 -1145
rect 443 -1146 444 -1106
rect 450 -1217 451 -1145
rect 499 -1217 500 -1145
rect 737 -1217 738 -1145
rect 758 -1217 759 -1145
rect 831 -1217 832 -1145
rect 1055 -1146 1056 -1106
rect 1353 -1146 1354 -1106
rect 1402 -1146 1403 -1106
rect 1528 -1217 1529 -1145
rect 1556 -1146 1557 -1106
rect 1738 -1217 1739 -1145
rect 51 -1148 52 -1106
rect 1353 -1217 1354 -1147
rect 1409 -1148 1410 -1106
rect 1654 -1217 1655 -1147
rect 51 -1217 52 -1149
rect 597 -1217 598 -1149
rect 611 -1150 612 -1106
rect 723 -1217 724 -1149
rect 765 -1217 766 -1149
rect 884 -1217 885 -1149
rect 1055 -1217 1056 -1149
rect 1185 -1217 1186 -1149
rect 1269 -1150 1270 -1106
rect 1367 -1217 1368 -1149
rect 1416 -1150 1417 -1106
rect 1549 -1217 1550 -1149
rect 1577 -1150 1578 -1106
rect 1731 -1217 1732 -1149
rect 65 -1152 66 -1106
rect 79 -1217 80 -1151
rect 124 -1217 125 -1151
rect 968 -1217 969 -1151
rect 1066 -1152 1067 -1106
rect 1255 -1217 1256 -1151
rect 1276 -1152 1277 -1106
rect 1402 -1217 1403 -1151
rect 1416 -1217 1417 -1151
rect 1745 -1217 1746 -1151
rect 65 -1217 66 -1153
rect 1479 -1217 1480 -1153
rect 1535 -1154 1536 -1106
rect 1556 -1217 1557 -1153
rect 1577 -1217 1578 -1153
rect 1633 -1154 1634 -1106
rect 142 -1156 143 -1106
rect 492 -1217 493 -1155
rect 520 -1156 521 -1106
rect 667 -1217 668 -1155
rect 768 -1217 769 -1155
rect 842 -1156 843 -1106
rect 905 -1156 906 -1106
rect 1269 -1217 1270 -1155
rect 1283 -1156 1284 -1106
rect 1409 -1217 1410 -1155
rect 1486 -1156 1487 -1106
rect 1633 -1217 1634 -1155
rect 184 -1217 185 -1157
rect 583 -1158 584 -1106
rect 779 -1158 780 -1106
rect 1430 -1217 1431 -1157
rect 1598 -1158 1599 -1106
rect 1787 -1217 1788 -1157
rect 191 -1160 192 -1106
rect 191 -1217 192 -1159
rect 191 -1160 192 -1106
rect 191 -1217 192 -1159
rect 198 -1160 199 -1106
rect 310 -1217 311 -1159
rect 338 -1160 339 -1106
rect 842 -1217 843 -1159
rect 880 -1160 881 -1106
rect 1283 -1217 1284 -1159
rect 1388 -1160 1389 -1106
rect 1535 -1217 1536 -1159
rect 198 -1217 199 -1161
rect 254 -1162 255 -1106
rect 282 -1162 283 -1106
rect 646 -1217 647 -1161
rect 793 -1162 794 -1106
rect 919 -1217 920 -1161
rect 1003 -1162 1004 -1106
rect 1276 -1217 1277 -1161
rect 1458 -1162 1459 -1106
rect 1598 -1217 1599 -1161
rect 177 -1217 178 -1163
rect 254 -1217 255 -1163
rect 261 -1164 262 -1106
rect 1003 -1217 1004 -1163
rect 1052 -1164 1053 -1106
rect 1486 -1217 1487 -1163
rect 212 -1217 213 -1165
rect 803 -1166 804 -1106
rect 821 -1166 822 -1106
rect 905 -1217 906 -1165
rect 1066 -1217 1067 -1165
rect 1542 -1166 1543 -1106
rect 219 -1217 220 -1167
rect 264 -1217 265 -1167
rect 282 -1217 283 -1167
rect 425 -1168 426 -1106
rect 443 -1217 444 -1167
rect 695 -1168 696 -1106
rect 793 -1217 794 -1167
rect 1073 -1168 1074 -1106
rect 1087 -1168 1088 -1106
rect 1129 -1168 1130 -1106
rect 1143 -1168 1144 -1106
rect 1388 -1217 1389 -1167
rect 1458 -1217 1459 -1167
rect 1591 -1168 1592 -1106
rect 226 -1170 227 -1106
rect 639 -1170 640 -1106
rect 688 -1217 689 -1169
rect 821 -1217 822 -1169
rect 961 -1170 962 -1106
rect 1073 -1217 1074 -1169
rect 1094 -1170 1095 -1106
rect 1346 -1217 1347 -1169
rect 1521 -1170 1522 -1106
rect 1542 -1217 1543 -1169
rect 1584 -1170 1585 -1106
rect 1591 -1217 1592 -1169
rect 30 -1172 31 -1106
rect 226 -1217 227 -1171
rect 247 -1172 248 -1106
rect 485 -1217 486 -1171
rect 520 -1217 521 -1171
rect 894 -1172 895 -1106
rect 996 -1172 997 -1106
rect 1094 -1217 1095 -1171
rect 1101 -1172 1102 -1106
rect 1199 -1217 1200 -1171
rect 1395 -1172 1396 -1106
rect 1521 -1217 1522 -1171
rect 30 -1217 31 -1173
rect 86 -1174 87 -1106
rect 205 -1174 206 -1106
rect 247 -1217 248 -1173
rect 296 -1174 297 -1106
rect 429 -1217 430 -1173
rect 471 -1217 472 -1173
rect 894 -1217 895 -1173
rect 1010 -1174 1011 -1106
rect 1129 -1217 1130 -1173
rect 1150 -1174 1151 -1106
rect 1241 -1217 1242 -1173
rect 86 -1217 87 -1175
rect 163 -1176 164 -1106
rect 205 -1217 206 -1175
rect 457 -1176 458 -1106
rect 527 -1176 528 -1106
rect 611 -1217 612 -1175
rect 618 -1176 619 -1106
rect 639 -1217 640 -1175
rect 695 -1217 696 -1175
rect 1360 -1176 1361 -1106
rect 149 -1178 150 -1106
rect 163 -1217 164 -1177
rect 289 -1178 290 -1106
rect 296 -1217 297 -1177
rect 338 -1217 339 -1177
rect 436 -1178 437 -1106
rect 457 -1217 458 -1177
rect 534 -1178 535 -1106
rect 569 -1217 570 -1177
rect 709 -1178 710 -1106
rect 828 -1178 829 -1106
rect 961 -1217 962 -1177
rect 982 -1178 983 -1106
rect 1010 -1217 1011 -1177
rect 1017 -1178 1018 -1106
rect 1087 -1217 1088 -1177
rect 1101 -1217 1102 -1177
rect 1136 -1178 1137 -1106
rect 1157 -1178 1158 -1106
rect 1234 -1217 1235 -1177
rect 1360 -1217 1361 -1177
rect 1748 -1217 1749 -1177
rect 145 -1217 146 -1179
rect 149 -1217 150 -1179
rect 170 -1217 171 -1179
rect 1136 -1217 1137 -1179
rect 1164 -1180 1165 -1106
rect 1465 -1217 1466 -1179
rect 268 -1182 269 -1106
rect 436 -1217 437 -1181
rect 464 -1182 465 -1106
rect 534 -1217 535 -1181
rect 562 -1182 563 -1106
rect 709 -1217 710 -1181
rect 740 -1217 741 -1181
rect 1164 -1217 1165 -1181
rect 1171 -1182 1172 -1106
rect 1318 -1217 1319 -1181
rect 142 -1217 143 -1183
rect 268 -1217 269 -1183
rect 331 -1184 332 -1106
rect 464 -1217 465 -1183
rect 562 -1217 563 -1183
rect 674 -1184 675 -1106
rect 849 -1184 850 -1106
rect 1017 -1217 1018 -1183
rect 1038 -1184 1039 -1106
rect 1171 -1217 1172 -1183
rect 1178 -1184 1179 -1106
rect 1339 -1217 1340 -1183
rect 331 -1217 332 -1185
rect 359 -1186 360 -1106
rect 576 -1186 577 -1106
rect 779 -1217 780 -1185
rect 856 -1186 857 -1106
rect 982 -1217 983 -1185
rect 1059 -1186 1060 -1106
rect 1143 -1217 1144 -1185
rect 1178 -1217 1179 -1185
rect 1206 -1186 1207 -1106
rect 1227 -1186 1228 -1106
rect 1395 -1217 1396 -1185
rect 345 -1188 346 -1106
rect 359 -1217 360 -1187
rect 555 -1188 556 -1106
rect 576 -1217 577 -1187
rect 583 -1217 584 -1187
rect 733 -1188 734 -1106
rect 751 -1188 752 -1106
rect 849 -1217 850 -1187
rect 856 -1217 857 -1187
rect 996 -1217 997 -1187
rect 1080 -1188 1081 -1106
rect 1206 -1217 1207 -1187
rect 1227 -1217 1228 -1187
rect 1262 -1188 1263 -1106
rect 345 -1217 346 -1189
rect 481 -1190 482 -1106
rect 555 -1217 556 -1189
rect 632 -1190 633 -1106
rect 674 -1217 675 -1189
rect 807 -1190 808 -1106
rect 926 -1190 927 -1106
rect 1059 -1217 1060 -1189
rect 1108 -1190 1109 -1106
rect 1150 -1217 1151 -1189
rect 1192 -1190 1193 -1106
rect 1584 -1217 1585 -1189
rect 394 -1192 395 -1106
rect 1080 -1217 1081 -1191
rect 1115 -1192 1116 -1106
rect 1297 -1217 1298 -1191
rect 352 -1194 353 -1106
rect 394 -1217 395 -1193
rect 618 -1217 619 -1193
rect 828 -1217 829 -1193
rect 898 -1217 899 -1193
rect 926 -1217 927 -1193
rect 940 -1194 941 -1106
rect 1038 -1217 1039 -1193
rect 1122 -1194 1123 -1106
rect 1304 -1217 1305 -1193
rect 352 -1217 353 -1195
rect 373 -1196 374 -1106
rect 691 -1196 692 -1106
rect 1108 -1217 1109 -1195
rect 1262 -1217 1263 -1195
rect 1475 -1196 1476 -1106
rect 317 -1198 318 -1106
rect 373 -1217 374 -1197
rect 702 -1217 703 -1197
rect 1115 -1217 1116 -1197
rect 44 -1200 45 -1106
rect 317 -1217 318 -1199
rect 751 -1217 752 -1199
rect 863 -1200 864 -1106
rect 947 -1200 948 -1106
rect 1157 -1217 1158 -1199
rect 44 -1217 45 -1201
rect 156 -1202 157 -1106
rect 541 -1217 542 -1201
rect 863 -1217 864 -1201
rect 947 -1217 948 -1201
rect 1024 -1202 1025 -1106
rect 1031 -1202 1032 -1106
rect 1122 -1217 1123 -1201
rect 156 -1217 157 -1203
rect 590 -1204 591 -1106
rect 796 -1217 797 -1203
rect 807 -1217 808 -1203
rect 954 -1204 955 -1106
rect 1031 -1217 1032 -1203
rect 590 -1217 591 -1205
rect 660 -1206 661 -1106
rect 698 -1217 699 -1205
rect 954 -1217 955 -1205
rect 975 -1206 976 -1106
rect 1024 -1217 1025 -1205
rect 604 -1208 605 -1106
rect 660 -1217 661 -1207
rect 814 -1208 815 -1106
rect 975 -1217 976 -1207
rect 989 -1208 990 -1106
rect 1192 -1217 1193 -1207
rect 527 -1217 528 -1209
rect 604 -1217 605 -1209
rect 814 -1217 815 -1209
rect 940 -1217 941 -1209
rect 870 -1212 871 -1106
rect 989 -1217 990 -1211
rect 240 -1214 241 -1106
rect 870 -1217 871 -1213
rect 240 -1217 241 -1215
rect 289 -1217 290 -1215
rect 16 -1360 17 -1226
rect 446 -1360 447 -1226
rect 471 -1227 472 -1225
rect 471 -1360 472 -1226
rect 471 -1227 472 -1225
rect 471 -1360 472 -1226
rect 506 -1227 507 -1225
rect 863 -1227 864 -1225
rect 891 -1227 892 -1225
rect 1087 -1227 1088 -1225
rect 1094 -1227 1095 -1225
rect 1202 -1360 1203 -1226
rect 1276 -1227 1277 -1225
rect 1276 -1360 1277 -1226
rect 1276 -1227 1277 -1225
rect 1276 -1360 1277 -1226
rect 1283 -1227 1284 -1225
rect 1283 -1360 1284 -1226
rect 1283 -1227 1284 -1225
rect 1283 -1360 1284 -1226
rect 1290 -1227 1291 -1225
rect 1293 -1243 1294 -1226
rect 1311 -1227 1312 -1225
rect 1314 -1227 1315 -1225
rect 1451 -1227 1452 -1225
rect 1451 -1360 1452 -1226
rect 1451 -1227 1452 -1225
rect 1451 -1360 1452 -1226
rect 1661 -1227 1662 -1225
rect 1661 -1360 1662 -1226
rect 1661 -1227 1662 -1225
rect 1661 -1360 1662 -1226
rect 1703 -1227 1704 -1225
rect 1748 -1227 1749 -1225
rect 1766 -1227 1767 -1225
rect 1787 -1227 1788 -1225
rect 44 -1229 45 -1225
rect 264 -1229 265 -1225
rect 289 -1229 290 -1225
rect 509 -1229 510 -1225
rect 548 -1229 549 -1225
rect 565 -1229 566 -1225
rect 590 -1229 591 -1225
rect 597 -1229 598 -1225
rect 607 -1229 608 -1225
rect 1269 -1229 1270 -1225
rect 1290 -1360 1291 -1228
rect 1311 -1360 1312 -1228
rect 1318 -1229 1319 -1225
rect 1696 -1229 1697 -1225
rect 1703 -1360 1704 -1228
rect 1745 -1229 1746 -1225
rect 1759 -1229 1760 -1225
rect 44 -1360 45 -1230
rect 89 -1231 90 -1225
rect 93 -1231 94 -1225
rect 93 -1360 94 -1230
rect 93 -1231 94 -1225
rect 93 -1360 94 -1230
rect 103 -1360 104 -1230
rect 303 -1231 304 -1225
rect 345 -1231 346 -1225
rect 796 -1231 797 -1225
rect 800 -1231 801 -1225
rect 863 -1360 864 -1230
rect 894 -1231 895 -1225
rect 1612 -1231 1613 -1225
rect 1745 -1360 1746 -1230
rect 1776 -1231 1777 -1225
rect 65 -1233 66 -1225
rect 1353 -1233 1354 -1225
rect 1612 -1360 1613 -1232
rect 1717 -1233 1718 -1225
rect 54 -1360 55 -1234
rect 65 -1360 66 -1234
rect 68 -1235 69 -1225
rect 79 -1235 80 -1225
rect 107 -1235 108 -1225
rect 114 -1235 115 -1225
rect 121 -1235 122 -1225
rect 1374 -1235 1375 -1225
rect 1717 -1360 1718 -1234
rect 1731 -1235 1732 -1225
rect 72 -1237 73 -1225
rect 653 -1360 654 -1236
rect 709 -1237 710 -1225
rect 793 -1237 794 -1225
rect 817 -1237 818 -1225
rect 961 -1237 962 -1225
rect 1010 -1237 1011 -1225
rect 1094 -1360 1095 -1236
rect 1146 -1360 1147 -1236
rect 1465 -1237 1466 -1225
rect 51 -1239 52 -1225
rect 72 -1360 73 -1238
rect 110 -1239 111 -1225
rect 660 -1239 661 -1225
rect 667 -1239 668 -1225
rect 793 -1360 794 -1238
rect 821 -1239 822 -1225
rect 1619 -1239 1620 -1225
rect 114 -1360 115 -1240
rect 940 -1241 941 -1225
rect 947 -1360 948 -1240
rect 1535 -1241 1536 -1225
rect 121 -1360 122 -1242
rect 453 -1360 454 -1242
rect 551 -1360 552 -1242
rect 1136 -1243 1137 -1225
rect 1178 -1243 1179 -1225
rect 1178 -1360 1179 -1242
rect 1178 -1243 1179 -1225
rect 1178 -1360 1179 -1242
rect 1248 -1243 1249 -1225
rect 1269 -1360 1270 -1242
rect 1314 -1360 1315 -1242
rect 1318 -1360 1319 -1242
rect 1353 -1360 1354 -1242
rect 1479 -1243 1480 -1225
rect 1486 -1243 1487 -1225
rect 1535 -1360 1536 -1242
rect 124 -1245 125 -1225
rect 478 -1245 479 -1225
rect 565 -1360 566 -1244
rect 716 -1245 717 -1225
rect 737 -1245 738 -1225
rect 744 -1245 745 -1225
rect 751 -1245 752 -1225
rect 765 -1360 766 -1244
rect 779 -1245 780 -1225
rect 800 -1360 801 -1244
rect 821 -1360 822 -1244
rect 1542 -1245 1543 -1225
rect 61 -1360 62 -1246
rect 737 -1360 738 -1246
rect 740 -1247 741 -1225
rect 1332 -1247 1333 -1225
rect 1360 -1247 1361 -1225
rect 1374 -1360 1375 -1246
rect 1458 -1247 1459 -1225
rect 1731 -1360 1732 -1246
rect 145 -1249 146 -1225
rect 1556 -1249 1557 -1225
rect 170 -1251 171 -1225
rect 177 -1251 178 -1225
rect 180 -1251 181 -1225
rect 1738 -1251 1739 -1225
rect 142 -1253 143 -1225
rect 170 -1360 171 -1252
rect 177 -1360 178 -1252
rect 198 -1253 199 -1225
rect 208 -1360 209 -1252
rect 240 -1360 241 -1252
rect 243 -1253 244 -1225
rect 1157 -1253 1158 -1225
rect 1220 -1253 1221 -1225
rect 1248 -1360 1249 -1252
rect 1325 -1253 1326 -1225
rect 1556 -1360 1557 -1252
rect 142 -1360 143 -1254
rect 212 -1255 213 -1225
rect 226 -1255 227 -1225
rect 1003 -1255 1004 -1225
rect 1010 -1360 1011 -1254
rect 1045 -1255 1046 -1225
rect 1052 -1255 1053 -1225
rect 1584 -1255 1585 -1225
rect 128 -1257 129 -1225
rect 212 -1360 213 -1256
rect 226 -1360 227 -1256
rect 254 -1257 255 -1225
rect 261 -1360 262 -1256
rect 436 -1257 437 -1225
rect 443 -1257 444 -1225
rect 1020 -1360 1021 -1256
rect 1059 -1257 1060 -1225
rect 1157 -1360 1158 -1256
rect 1171 -1257 1172 -1225
rect 1220 -1360 1221 -1256
rect 1325 -1360 1326 -1256
rect 1769 -1257 1770 -1225
rect 163 -1259 164 -1225
rect 254 -1360 255 -1258
rect 292 -1360 293 -1258
rect 870 -1259 871 -1225
rect 933 -1259 934 -1225
rect 1059 -1360 1060 -1258
rect 1087 -1360 1088 -1258
rect 1500 -1259 1501 -1225
rect 1542 -1360 1543 -1258
rect 1549 -1259 1550 -1225
rect 1584 -1360 1585 -1258
rect 1591 -1259 1592 -1225
rect 163 -1360 164 -1260
rect 705 -1261 706 -1225
rect 723 -1261 724 -1225
rect 744 -1360 745 -1260
rect 751 -1360 752 -1260
rect 768 -1261 769 -1225
rect 824 -1360 825 -1260
rect 1055 -1261 1056 -1225
rect 1101 -1261 1102 -1225
rect 1332 -1360 1333 -1260
rect 1402 -1261 1403 -1225
rect 1458 -1360 1459 -1260
rect 1465 -1360 1466 -1260
rect 1507 -1261 1508 -1225
rect 1549 -1360 1550 -1260
rect 1598 -1261 1599 -1225
rect 184 -1263 185 -1225
rect 709 -1360 710 -1262
rect 740 -1360 741 -1262
rect 1430 -1263 1431 -1225
rect 1479 -1360 1480 -1262
rect 1640 -1263 1641 -1225
rect 184 -1360 185 -1264
rect 618 -1265 619 -1225
rect 632 -1265 633 -1225
rect 1346 -1265 1347 -1225
rect 1402 -1360 1403 -1264
rect 1444 -1265 1445 -1225
rect 1486 -1360 1487 -1264
rect 1528 -1265 1529 -1225
rect 1570 -1265 1571 -1225
rect 1591 -1360 1592 -1264
rect 1598 -1360 1599 -1264
rect 1633 -1265 1634 -1225
rect 1640 -1360 1641 -1264
rect 1654 -1265 1655 -1225
rect 198 -1360 199 -1266
rect 779 -1360 780 -1266
rect 828 -1267 829 -1225
rect 1360 -1360 1361 -1266
rect 1423 -1267 1424 -1225
rect 1507 -1360 1508 -1266
rect 1528 -1360 1529 -1266
rect 1577 -1267 1578 -1225
rect 1633 -1360 1634 -1266
rect 1647 -1267 1648 -1225
rect 1654 -1360 1655 -1266
rect 1675 -1267 1676 -1225
rect 296 -1269 297 -1225
rect 604 -1269 605 -1225
rect 611 -1269 612 -1225
rect 632 -1360 633 -1268
rect 639 -1269 640 -1225
rect 660 -1360 661 -1268
rect 831 -1269 832 -1225
rect 1255 -1269 1256 -1225
rect 1339 -1269 1340 -1225
rect 1346 -1360 1347 -1268
rect 1423 -1360 1424 -1268
rect 1514 -1269 1515 -1225
rect 1577 -1360 1578 -1268
rect 1626 -1269 1627 -1225
rect 1647 -1360 1648 -1268
rect 1668 -1269 1669 -1225
rect 1675 -1360 1676 -1268
rect 1689 -1269 1690 -1225
rect 58 -1271 59 -1225
rect 604 -1360 605 -1270
rect 611 -1360 612 -1270
rect 912 -1271 913 -1225
rect 922 -1360 923 -1270
rect 1570 -1360 1571 -1270
rect 1682 -1271 1683 -1225
rect 1689 -1360 1690 -1270
rect 58 -1360 59 -1272
rect 100 -1273 101 -1225
rect 296 -1360 297 -1272
rect 352 -1273 353 -1225
rect 380 -1273 381 -1225
rect 695 -1273 696 -1225
rect 702 -1273 703 -1225
rect 1339 -1360 1340 -1272
rect 1500 -1360 1501 -1272
rect 1521 -1273 1522 -1225
rect 1682 -1360 1683 -1272
rect 1710 -1273 1711 -1225
rect 205 -1275 206 -1225
rect 352 -1360 353 -1274
rect 380 -1360 381 -1274
rect 597 -1360 598 -1274
rect 600 -1360 601 -1274
rect 639 -1360 640 -1274
rect 688 -1275 689 -1225
rect 702 -1360 703 -1274
rect 831 -1360 832 -1274
rect 1262 -1275 1263 -1225
rect 1710 -1360 1711 -1274
rect 1724 -1275 1725 -1225
rect 23 -1277 24 -1225
rect 205 -1360 206 -1276
rect 303 -1360 304 -1276
rect 331 -1277 332 -1225
rect 345 -1360 346 -1276
rect 373 -1277 374 -1225
rect 387 -1277 388 -1225
rect 590 -1360 591 -1276
rect 681 -1277 682 -1225
rect 688 -1360 689 -1276
rect 835 -1277 836 -1225
rect 891 -1360 892 -1276
rect 912 -1360 913 -1276
rect 982 -1277 983 -1225
rect 996 -1277 997 -1225
rect 1045 -1360 1046 -1276
rect 1101 -1360 1102 -1276
rect 1472 -1277 1473 -1225
rect 1724 -1360 1725 -1276
rect 1752 -1277 1753 -1225
rect 23 -1360 24 -1278
rect 541 -1279 542 -1225
rect 548 -1360 549 -1278
rect 1255 -1360 1256 -1278
rect 1752 -1360 1753 -1278
rect 1780 -1279 1781 -1225
rect 310 -1281 311 -1225
rect 716 -1360 717 -1280
rect 852 -1360 853 -1280
rect 919 -1281 920 -1225
rect 929 -1281 930 -1225
rect 1668 -1360 1669 -1280
rect 156 -1283 157 -1225
rect 310 -1360 311 -1282
rect 317 -1283 318 -1225
rect 387 -1360 388 -1282
rect 415 -1283 416 -1225
rect 506 -1360 507 -1282
rect 513 -1283 514 -1225
rect 870 -1360 871 -1282
rect 933 -1360 934 -1282
rect 1696 -1360 1697 -1282
rect 149 -1285 150 -1225
rect 156 -1360 157 -1284
rect 317 -1360 318 -1284
rect 789 -1360 790 -1284
rect 856 -1285 857 -1225
rect 1493 -1285 1494 -1225
rect 100 -1360 101 -1286
rect 1493 -1360 1494 -1286
rect 149 -1360 150 -1288
rect 877 -1289 878 -1225
rect 936 -1360 937 -1288
rect 1297 -1289 1298 -1225
rect 331 -1360 332 -1290
rect 359 -1291 360 -1225
rect 366 -1291 367 -1225
rect 541 -1360 542 -1290
rect 625 -1291 626 -1225
rect 681 -1360 682 -1290
rect 807 -1291 808 -1225
rect 877 -1360 878 -1290
rect 940 -1360 941 -1290
rect 1006 -1360 1007 -1290
rect 1017 -1291 1018 -1225
rect 1052 -1360 1053 -1290
rect 1104 -1360 1105 -1290
rect 1619 -1360 1620 -1290
rect 275 -1293 276 -1225
rect 625 -1360 626 -1292
rect 667 -1360 668 -1292
rect 982 -1360 983 -1292
rect 1038 -1293 1039 -1225
rect 1626 -1360 1627 -1292
rect 135 -1295 136 -1225
rect 275 -1360 276 -1294
rect 282 -1295 283 -1225
rect 366 -1360 367 -1294
rect 373 -1360 374 -1294
rect 464 -1295 465 -1225
rect 499 -1295 500 -1225
rect 723 -1360 724 -1294
rect 772 -1295 773 -1225
rect 807 -1360 808 -1294
rect 842 -1295 843 -1225
rect 856 -1360 857 -1294
rect 859 -1295 860 -1225
rect 1073 -1295 1074 -1225
rect 1115 -1295 1116 -1225
rect 1738 -1360 1739 -1294
rect 82 -1360 83 -1296
rect 135 -1360 136 -1296
rect 187 -1360 188 -1296
rect 499 -1360 500 -1296
rect 635 -1297 636 -1225
rect 1038 -1360 1039 -1296
rect 1108 -1297 1109 -1225
rect 1115 -1360 1116 -1296
rect 1129 -1297 1130 -1225
rect 1136 -1360 1137 -1296
rect 1150 -1297 1151 -1225
rect 1297 -1360 1298 -1296
rect 191 -1299 192 -1225
rect 464 -1360 465 -1298
rect 558 -1360 559 -1298
rect 1129 -1360 1130 -1298
rect 1143 -1299 1144 -1225
rect 1150 -1360 1151 -1298
rect 1164 -1299 1165 -1225
rect 1171 -1360 1172 -1298
rect 1192 -1299 1193 -1225
rect 1521 -1360 1522 -1298
rect 191 -1360 192 -1300
rect 975 -1301 976 -1225
rect 1031 -1301 1032 -1225
rect 1073 -1360 1074 -1300
rect 1080 -1301 1081 -1225
rect 1108 -1360 1109 -1300
rect 1164 -1360 1165 -1300
rect 1206 -1301 1207 -1225
rect 1227 -1301 1228 -1225
rect 1472 -1360 1473 -1300
rect 247 -1303 248 -1225
rect 282 -1360 283 -1302
rect 338 -1303 339 -1225
rect 415 -1360 416 -1302
rect 422 -1303 423 -1225
rect 835 -1360 836 -1302
rect 950 -1303 951 -1225
rect 1514 -1360 1515 -1302
rect 173 -1305 174 -1225
rect 338 -1360 339 -1304
rect 359 -1360 360 -1304
rect 656 -1305 657 -1225
rect 674 -1305 675 -1225
rect 772 -1360 773 -1304
rect 950 -1360 951 -1304
rect 961 -1360 962 -1304
rect 989 -1305 990 -1225
rect 1031 -1360 1032 -1304
rect 1080 -1360 1081 -1304
rect 1185 -1305 1186 -1225
rect 1206 -1360 1207 -1304
rect 1213 -1305 1214 -1225
rect 1234 -1305 1235 -1225
rect 1430 -1360 1431 -1304
rect 86 -1307 87 -1225
rect 674 -1360 675 -1306
rect 695 -1360 696 -1306
rect 1213 -1360 1214 -1306
rect 1241 -1307 1242 -1225
rect 1262 -1360 1263 -1306
rect 86 -1360 87 -1308
rect 527 -1309 528 -1225
rect 562 -1309 563 -1225
rect 1192 -1360 1193 -1308
rect 247 -1360 248 -1310
rect 268 -1311 269 -1225
rect 408 -1311 409 -1225
rect 842 -1360 843 -1310
rect 926 -1311 927 -1225
rect 1234 -1360 1235 -1310
rect 222 -1360 223 -1312
rect 268 -1360 269 -1312
rect 324 -1313 325 -1225
rect 408 -1360 409 -1312
rect 422 -1360 423 -1312
rect 754 -1360 755 -1312
rect 898 -1313 899 -1225
rect 926 -1360 927 -1312
rect 954 -1313 955 -1225
rect 989 -1360 990 -1312
rect 1003 -1360 1004 -1312
rect 1185 -1360 1186 -1312
rect 324 -1360 325 -1314
rect 968 -1315 969 -1225
rect 1024 -1315 1025 -1225
rect 1241 -1360 1242 -1314
rect 436 -1360 437 -1316
rect 758 -1317 759 -1225
rect 849 -1317 850 -1225
rect 1024 -1360 1025 -1316
rect 450 -1319 451 -1225
rect 478 -1360 479 -1318
rect 485 -1319 486 -1225
rect 562 -1360 563 -1318
rect 572 -1360 573 -1318
rect 1227 -1360 1228 -1318
rect 450 -1360 451 -1320
rect 996 -1360 997 -1320
rect 457 -1323 458 -1225
rect 513 -1360 514 -1322
rect 555 -1323 556 -1225
rect 758 -1360 759 -1322
rect 884 -1323 885 -1225
rect 968 -1360 969 -1322
rect 401 -1325 402 -1225
rect 555 -1360 556 -1324
rect 583 -1325 584 -1225
rect 898 -1360 899 -1324
rect 905 -1325 906 -1225
rect 954 -1360 955 -1324
rect 394 -1327 395 -1225
rect 401 -1360 402 -1326
rect 429 -1327 430 -1225
rect 884 -1360 885 -1326
rect 219 -1329 220 -1225
rect 429 -1360 430 -1328
rect 457 -1360 458 -1328
rect 534 -1329 535 -1225
rect 618 -1360 619 -1328
rect 849 -1360 850 -1328
rect 394 -1360 395 -1330
rect 576 -1331 577 -1225
rect 698 -1331 699 -1225
rect 975 -1360 976 -1330
rect 37 -1333 38 -1225
rect 576 -1360 577 -1332
rect 786 -1333 787 -1225
rect 905 -1360 906 -1332
rect 492 -1335 493 -1225
rect 527 -1360 528 -1334
rect 534 -1360 535 -1334
rect 814 -1335 815 -1225
rect 233 -1337 234 -1225
rect 492 -1360 493 -1336
rect 520 -1337 521 -1225
rect 583 -1360 584 -1336
rect 646 -1360 647 -1336
rect 814 -1360 815 -1336
rect 30 -1339 31 -1225
rect 233 -1360 234 -1338
rect 520 -1360 521 -1338
rect 730 -1339 731 -1225
rect 786 -1360 787 -1338
rect 1367 -1339 1368 -1225
rect 30 -1360 31 -1340
rect 569 -1341 570 -1225
rect 730 -1360 731 -1340
rect 1066 -1341 1067 -1225
rect 1367 -1360 1368 -1340
rect 1381 -1341 1382 -1225
rect 485 -1360 486 -1342
rect 569 -1360 570 -1342
rect 1066 -1360 1067 -1342
rect 1122 -1343 1123 -1225
rect 1381 -1360 1382 -1342
rect 1388 -1343 1389 -1225
rect 1122 -1360 1123 -1344
rect 1199 -1345 1200 -1225
rect 1388 -1360 1389 -1344
rect 1395 -1345 1396 -1225
rect 1199 -1360 1200 -1346
rect 1444 -1360 1445 -1346
rect 1395 -1360 1396 -1348
rect 1409 -1349 1410 -1225
rect 1409 -1360 1410 -1350
rect 1416 -1351 1417 -1225
rect 1416 -1360 1417 -1352
rect 1437 -1353 1438 -1225
rect 1437 -1360 1438 -1354
rect 1563 -1355 1564 -1225
rect 1563 -1360 1564 -1356
rect 1605 -1357 1606 -1225
rect 817 -1360 818 -1358
rect 1605 -1360 1606 -1358
rect 16 -1370 17 -1368
rect 110 -1370 111 -1368
rect 121 -1370 122 -1368
rect 208 -1370 209 -1368
rect 219 -1370 220 -1368
rect 1038 -1370 1039 -1368
rect 1048 -1501 1049 -1369
rect 1094 -1370 1095 -1368
rect 1104 -1370 1105 -1368
rect 1689 -1370 1690 -1368
rect 1738 -1370 1739 -1368
rect 1801 -1501 1802 -1369
rect 51 -1372 52 -1368
rect 93 -1372 94 -1368
rect 100 -1372 101 -1368
rect 100 -1501 101 -1371
rect 100 -1372 101 -1368
rect 100 -1501 101 -1371
rect 107 -1501 108 -1371
rect 646 -1372 647 -1368
rect 688 -1372 689 -1368
rect 688 -1501 689 -1371
rect 688 -1372 689 -1368
rect 688 -1501 689 -1371
rect 719 -1501 720 -1371
rect 1024 -1372 1025 -1368
rect 1038 -1501 1039 -1371
rect 1108 -1372 1109 -1368
rect 1146 -1372 1147 -1368
rect 1661 -1372 1662 -1368
rect 1689 -1501 1690 -1371
rect 1696 -1372 1697 -1368
rect 51 -1501 52 -1373
rect 149 -1374 150 -1368
rect 159 -1501 160 -1373
rect 177 -1374 178 -1368
rect 187 -1501 188 -1373
rect 765 -1374 766 -1368
rect 814 -1374 815 -1368
rect 1136 -1374 1137 -1368
rect 1164 -1374 1165 -1368
rect 1164 -1501 1165 -1373
rect 1164 -1374 1165 -1368
rect 1164 -1501 1165 -1373
rect 1199 -1501 1200 -1373
rect 1346 -1374 1347 -1368
rect 1591 -1374 1592 -1368
rect 1696 -1501 1697 -1373
rect 58 -1501 59 -1375
rect 618 -1376 619 -1368
rect 646 -1501 647 -1375
rect 660 -1376 661 -1368
rect 744 -1376 745 -1368
rect 744 -1501 745 -1375
rect 744 -1376 745 -1368
rect 744 -1501 745 -1375
rect 751 -1376 752 -1368
rect 1290 -1376 1291 -1368
rect 1346 -1501 1347 -1375
rect 1395 -1376 1396 -1368
rect 1591 -1501 1592 -1375
rect 1633 -1376 1634 -1368
rect 65 -1378 66 -1368
rect 79 -1378 80 -1368
rect 82 -1378 83 -1368
rect 1374 -1378 1375 -1368
rect 1395 -1501 1396 -1377
rect 1402 -1378 1403 -1368
rect 1528 -1378 1529 -1368
rect 1633 -1501 1634 -1377
rect 79 -1501 80 -1379
rect 940 -1380 941 -1368
rect 978 -1501 979 -1379
rect 1500 -1380 1501 -1368
rect 1612 -1380 1613 -1368
rect 1661 -1501 1662 -1379
rect 93 -1501 94 -1381
rect 520 -1382 521 -1368
rect 551 -1382 552 -1368
rect 835 -1382 836 -1368
rect 849 -1382 850 -1368
rect 1325 -1382 1326 -1368
rect 1374 -1501 1375 -1381
rect 1409 -1382 1410 -1368
rect 1437 -1382 1438 -1368
rect 1528 -1501 1529 -1381
rect 1612 -1501 1613 -1381
rect 1647 -1382 1648 -1368
rect 124 -1501 125 -1383
rect 716 -1384 717 -1368
rect 751 -1501 752 -1383
rect 758 -1384 759 -1368
rect 761 -1501 762 -1383
rect 1626 -1384 1627 -1368
rect 1647 -1501 1648 -1383
rect 1682 -1384 1683 -1368
rect 149 -1501 150 -1385
rect 824 -1386 825 -1368
rect 831 -1501 832 -1385
rect 1220 -1386 1221 -1368
rect 1227 -1386 1228 -1368
rect 1409 -1501 1410 -1385
rect 1500 -1501 1501 -1385
rect 1556 -1386 1557 -1368
rect 1626 -1501 1627 -1385
rect 1675 -1386 1676 -1368
rect 156 -1388 157 -1368
rect 177 -1501 178 -1387
rect 194 -1501 195 -1387
rect 282 -1388 283 -1368
rect 289 -1501 290 -1387
rect 471 -1388 472 -1368
rect 478 -1388 479 -1368
rect 516 -1501 517 -1387
rect 520 -1501 521 -1387
rect 1031 -1388 1032 -1368
rect 1034 -1501 1035 -1387
rect 1682 -1501 1683 -1387
rect 103 -1390 104 -1368
rect 1031 -1501 1032 -1389
rect 1066 -1390 1067 -1368
rect 1094 -1501 1095 -1389
rect 1108 -1501 1109 -1389
rect 1248 -1390 1249 -1368
rect 1402 -1501 1403 -1389
rect 1587 -1501 1588 -1389
rect 156 -1501 157 -1391
rect 292 -1392 293 -1368
rect 317 -1392 318 -1368
rect 618 -1501 619 -1391
rect 625 -1392 626 -1368
rect 660 -1501 661 -1391
rect 758 -1501 759 -1391
rect 1325 -1501 1326 -1391
rect 1556 -1501 1557 -1391
rect 1563 -1392 1564 -1368
rect 170 -1394 171 -1368
rect 205 -1394 206 -1368
rect 219 -1501 220 -1393
rect 310 -1394 311 -1368
rect 324 -1394 325 -1368
rect 670 -1501 671 -1393
rect 786 -1501 787 -1393
rect 1136 -1501 1137 -1393
rect 1202 -1394 1203 -1368
rect 1703 -1394 1704 -1368
rect 114 -1396 115 -1368
rect 205 -1501 206 -1395
rect 222 -1396 223 -1368
rect 1339 -1396 1340 -1368
rect 1563 -1501 1564 -1395
rect 1668 -1396 1669 -1368
rect 114 -1501 115 -1397
rect 716 -1501 717 -1397
rect 789 -1398 790 -1368
rect 940 -1501 941 -1397
rect 982 -1398 983 -1368
rect 1731 -1398 1732 -1368
rect 170 -1501 171 -1399
rect 639 -1400 640 -1368
rect 817 -1400 818 -1368
rect 1220 -1501 1221 -1399
rect 1227 -1501 1228 -1399
rect 1255 -1400 1256 -1368
rect 1339 -1501 1340 -1399
rect 1381 -1400 1382 -1368
rect 1584 -1400 1585 -1368
rect 1668 -1501 1669 -1399
rect 1731 -1501 1732 -1399
rect 1745 -1400 1746 -1368
rect 163 -1402 164 -1368
rect 639 -1501 640 -1401
rect 821 -1501 822 -1401
rect 1332 -1402 1333 -1368
rect 1381 -1501 1382 -1401
rect 1430 -1402 1431 -1368
rect 1584 -1501 1585 -1401
rect 1703 -1501 1704 -1401
rect 163 -1501 164 -1403
rect 254 -1404 255 -1368
rect 257 -1501 258 -1403
rect 611 -1404 612 -1368
rect 849 -1501 850 -1403
rect 891 -1404 892 -1368
rect 919 -1404 920 -1368
rect 1608 -1501 1609 -1403
rect 198 -1406 199 -1368
rect 541 -1406 542 -1368
rect 555 -1406 556 -1368
rect 905 -1406 906 -1368
rect 919 -1501 920 -1405
rect 926 -1406 927 -1368
rect 982 -1501 983 -1405
rect 996 -1406 997 -1368
rect 1003 -1501 1004 -1405
rect 1213 -1406 1214 -1368
rect 1216 -1406 1217 -1368
rect 1507 -1406 1508 -1368
rect 54 -1408 55 -1368
rect 996 -1501 997 -1407
rect 1006 -1408 1007 -1368
rect 1472 -1408 1473 -1368
rect 1507 -1501 1508 -1407
rect 1598 -1408 1599 -1368
rect 135 -1410 136 -1368
rect 198 -1501 199 -1409
rect 201 -1410 202 -1368
rect 1437 -1501 1438 -1409
rect 1472 -1501 1473 -1409
rect 1605 -1410 1606 -1368
rect 135 -1501 136 -1411
rect 142 -1412 143 -1368
rect 226 -1412 227 -1368
rect 282 -1501 283 -1411
rect 310 -1501 311 -1411
rect 457 -1412 458 -1368
rect 471 -1501 472 -1411
rect 485 -1412 486 -1368
rect 506 -1412 507 -1368
rect 555 -1501 556 -1411
rect 558 -1412 559 -1368
rect 1570 -1412 1571 -1368
rect 1598 -1501 1599 -1411
rect 1724 -1412 1725 -1368
rect 142 -1501 143 -1413
rect 212 -1414 213 -1368
rect 229 -1501 230 -1413
rect 303 -1414 304 -1368
rect 366 -1414 367 -1368
rect 485 -1501 486 -1413
rect 541 -1501 542 -1413
rect 933 -1414 934 -1368
rect 1010 -1414 1011 -1368
rect 1024 -1501 1025 -1413
rect 1066 -1501 1067 -1413
rect 1115 -1414 1116 -1368
rect 1157 -1414 1158 -1368
rect 1605 -1501 1606 -1413
rect 191 -1416 192 -1368
rect 212 -1501 213 -1415
rect 215 -1501 216 -1415
rect 366 -1501 367 -1415
rect 380 -1416 381 -1368
rect 506 -1501 507 -1415
rect 562 -1416 563 -1368
rect 835 -1501 836 -1415
rect 891 -1501 892 -1415
rect 954 -1416 955 -1368
rect 1010 -1501 1011 -1415
rect 1059 -1416 1060 -1368
rect 1115 -1501 1116 -1415
rect 1150 -1416 1151 -1368
rect 1157 -1501 1158 -1415
rect 1192 -1416 1193 -1368
rect 1213 -1501 1214 -1415
rect 1262 -1416 1263 -1368
rect 1332 -1501 1333 -1415
rect 1535 -1416 1536 -1368
rect 37 -1501 38 -1417
rect 191 -1501 192 -1417
rect 240 -1418 241 -1368
rect 324 -1501 325 -1417
rect 380 -1501 381 -1417
rect 513 -1418 514 -1368
rect 562 -1501 563 -1417
rect 681 -1418 682 -1368
rect 730 -1418 731 -1368
rect 926 -1501 927 -1417
rect 933 -1501 934 -1417
rect 1290 -1501 1291 -1417
rect 1318 -1418 1319 -1368
rect 1535 -1501 1536 -1417
rect 86 -1420 87 -1368
rect 730 -1501 731 -1419
rect 922 -1420 923 -1368
rect 1234 -1420 1235 -1368
rect 1248 -1501 1249 -1419
rect 1276 -1420 1277 -1368
rect 1318 -1501 1319 -1419
rect 1416 -1420 1417 -1368
rect 1430 -1501 1431 -1419
rect 1451 -1420 1452 -1368
rect 1479 -1420 1480 -1368
rect 1570 -1501 1571 -1419
rect 86 -1501 87 -1421
rect 793 -1422 794 -1368
rect 950 -1422 951 -1368
rect 1451 -1501 1452 -1421
rect 1479 -1501 1480 -1421
rect 1654 -1422 1655 -1368
rect 254 -1501 255 -1423
rect 303 -1501 304 -1423
rect 387 -1424 388 -1368
rect 814 -1501 815 -1423
rect 954 -1501 955 -1423
rect 968 -1424 969 -1368
rect 1017 -1424 1018 -1368
rect 1675 -1501 1676 -1423
rect 61 -1426 62 -1368
rect 387 -1501 388 -1425
rect 408 -1426 409 -1368
rect 765 -1501 766 -1425
rect 793 -1501 794 -1425
rect 800 -1426 801 -1368
rect 968 -1501 969 -1425
rect 1045 -1426 1046 -1368
rect 1059 -1501 1060 -1425
rect 1129 -1426 1130 -1368
rect 1192 -1501 1193 -1425
rect 1269 -1426 1270 -1368
rect 1276 -1501 1277 -1425
rect 1577 -1426 1578 -1368
rect 268 -1428 269 -1368
rect 1101 -1428 1102 -1368
rect 1129 -1501 1130 -1427
rect 1171 -1428 1172 -1368
rect 1255 -1501 1256 -1427
rect 1297 -1428 1298 -1368
rect 1416 -1501 1417 -1427
rect 1514 -1428 1515 -1368
rect 1538 -1501 1539 -1427
rect 1654 -1501 1655 -1427
rect 268 -1501 269 -1429
rect 296 -1430 297 -1368
rect 408 -1501 409 -1429
rect 604 -1430 605 -1368
rect 611 -1501 612 -1429
rect 740 -1430 741 -1368
rect 1017 -1501 1018 -1429
rect 1073 -1430 1074 -1368
rect 1080 -1430 1081 -1368
rect 1150 -1501 1151 -1429
rect 1171 -1501 1172 -1429
rect 1206 -1430 1207 -1368
rect 1262 -1501 1263 -1429
rect 1304 -1430 1305 -1368
rect 1577 -1501 1578 -1429
rect 1619 -1430 1620 -1368
rect 184 -1501 185 -1431
rect 1619 -1501 1620 -1431
rect 275 -1434 276 -1368
rect 481 -1501 482 -1433
rect 499 -1434 500 -1368
rect 800 -1501 801 -1433
rect 975 -1434 976 -1368
rect 1073 -1501 1074 -1433
rect 1143 -1434 1144 -1368
rect 1514 -1501 1515 -1433
rect 275 -1501 276 -1435
rect 828 -1436 829 -1368
rect 1020 -1436 1021 -1368
rect 1122 -1436 1123 -1368
rect 1143 -1501 1144 -1435
rect 1178 -1436 1179 -1368
rect 1297 -1501 1298 -1435
rect 1493 -1436 1494 -1368
rect 296 -1501 297 -1437
rect 464 -1438 465 -1368
rect 478 -1501 479 -1437
rect 1206 -1501 1207 -1437
rect 1304 -1501 1305 -1437
rect 1353 -1438 1354 -1368
rect 1360 -1438 1361 -1368
rect 1493 -1501 1494 -1437
rect 44 -1440 45 -1368
rect 464 -1501 465 -1439
rect 499 -1501 500 -1439
rect 534 -1440 535 -1368
rect 569 -1440 570 -1368
rect 1052 -1440 1053 -1368
rect 1178 -1501 1179 -1439
rect 1185 -1440 1186 -1368
rect 1353 -1501 1354 -1439
rect 1444 -1440 1445 -1368
rect 44 -1501 45 -1441
rect 72 -1442 73 -1368
rect 415 -1442 416 -1368
rect 572 -1442 573 -1368
rect 597 -1442 598 -1368
rect 737 -1442 738 -1368
rect 779 -1442 780 -1368
rect 1080 -1501 1081 -1441
rect 1185 -1501 1186 -1441
rect 1311 -1442 1312 -1368
rect 1360 -1501 1361 -1441
rect 1465 -1442 1466 -1368
rect 72 -1501 73 -1443
rect 226 -1501 227 -1443
rect 240 -1501 241 -1443
rect 737 -1501 738 -1443
rect 1045 -1501 1046 -1443
rect 1458 -1444 1459 -1368
rect 1465 -1501 1466 -1443
rect 1640 -1444 1641 -1368
rect 247 -1446 248 -1368
rect 415 -1501 416 -1445
rect 436 -1446 437 -1368
rect 947 -1446 948 -1368
rect 1052 -1501 1053 -1445
rect 1241 -1446 1242 -1368
rect 1444 -1501 1445 -1445
rect 1486 -1446 1487 -1368
rect 247 -1501 248 -1447
rect 338 -1448 339 -1368
rect 436 -1501 437 -1447
rect 936 -1448 937 -1368
rect 947 -1501 948 -1447
rect 1717 -1448 1718 -1368
rect 261 -1450 262 -1368
rect 338 -1501 339 -1449
rect 450 -1501 451 -1449
rect 667 -1450 668 -1368
rect 674 -1450 675 -1368
rect 1724 -1501 1725 -1449
rect 261 -1501 262 -1451
rect 331 -1452 332 -1368
rect 453 -1452 454 -1368
rect 842 -1452 843 -1368
rect 1241 -1501 1242 -1451
rect 1283 -1452 1284 -1368
rect 1458 -1501 1459 -1451
rect 1542 -1452 1543 -1368
rect 1710 -1452 1711 -1368
rect 1717 -1501 1718 -1451
rect 233 -1454 234 -1368
rect 842 -1501 843 -1453
rect 1283 -1501 1284 -1453
rect 1367 -1454 1368 -1368
rect 1486 -1501 1487 -1453
rect 1521 -1454 1522 -1368
rect 1542 -1501 1543 -1453
rect 1549 -1454 1550 -1368
rect 1643 -1501 1644 -1453
rect 1710 -1501 1711 -1453
rect 233 -1501 234 -1455
rect 422 -1456 423 -1368
rect 457 -1501 458 -1455
rect 905 -1501 906 -1455
rect 1367 -1501 1368 -1455
rect 1423 -1456 1424 -1368
rect 1549 -1501 1550 -1455
rect 1752 -1456 1753 -1368
rect 331 -1501 332 -1457
rect 548 -1458 549 -1368
rect 569 -1501 570 -1457
rect 590 -1458 591 -1368
rect 604 -1501 605 -1457
rect 870 -1458 871 -1368
rect 1388 -1458 1389 -1368
rect 1423 -1501 1424 -1457
rect 422 -1501 423 -1459
rect 936 -1501 937 -1459
rect 460 -1501 461 -1461
rect 1234 -1501 1235 -1461
rect 513 -1501 514 -1463
rect 1269 -1501 1270 -1463
rect 527 -1466 528 -1368
rect 597 -1501 598 -1465
rect 653 -1466 654 -1368
rect 674 -1501 675 -1465
rect 681 -1501 682 -1465
rect 807 -1466 808 -1368
rect 852 -1466 853 -1368
rect 1521 -1501 1522 -1465
rect 373 -1468 374 -1368
rect 527 -1501 528 -1467
rect 534 -1501 535 -1467
rect 824 -1501 825 -1467
rect 870 -1501 871 -1467
rect 877 -1468 878 -1368
rect 373 -1501 374 -1469
rect 492 -1470 493 -1368
rect 548 -1501 549 -1469
rect 950 -1501 951 -1469
rect 30 -1472 31 -1368
rect 492 -1501 493 -1471
rect 576 -1472 577 -1368
rect 779 -1501 780 -1471
rect 877 -1501 878 -1471
rect 884 -1472 885 -1368
rect 30 -1501 31 -1473
rect 131 -1474 132 -1368
rect 576 -1501 577 -1473
rect 632 -1474 633 -1368
rect 653 -1501 654 -1473
rect 1087 -1474 1088 -1368
rect 131 -1501 132 -1475
rect 583 -1476 584 -1368
rect 590 -1501 591 -1475
rect 985 -1476 986 -1368
rect 394 -1478 395 -1368
rect 583 -1501 584 -1477
rect 632 -1501 633 -1477
rect 989 -1478 990 -1368
rect 394 -1501 395 -1479
rect 429 -1480 430 -1368
rect 443 -1480 444 -1368
rect 1087 -1501 1088 -1479
rect 359 -1482 360 -1368
rect 429 -1501 430 -1481
rect 443 -1501 444 -1481
rect 702 -1482 703 -1368
rect 726 -1501 727 -1481
rect 1122 -1501 1123 -1481
rect 352 -1484 353 -1368
rect 359 -1501 360 -1483
rect 695 -1484 696 -1368
rect 1101 -1501 1102 -1483
rect 352 -1501 353 -1485
rect 401 -1486 402 -1368
rect 695 -1501 696 -1485
rect 723 -1486 724 -1368
rect 740 -1501 741 -1485
rect 1388 -1501 1389 -1485
rect 345 -1488 346 -1368
rect 401 -1501 402 -1487
rect 702 -1501 703 -1487
rect 828 -1501 829 -1487
rect 884 -1501 885 -1487
rect 898 -1488 899 -1368
rect 912 -1488 913 -1368
rect 989 -1501 990 -1487
rect 23 -1490 24 -1368
rect 345 -1501 346 -1489
rect 754 -1490 755 -1368
rect 807 -1501 808 -1489
rect 856 -1490 857 -1368
rect 898 -1501 899 -1489
rect 912 -1501 913 -1489
rect 961 -1490 962 -1368
rect 23 -1501 24 -1491
rect 128 -1492 129 -1368
rect 856 -1501 857 -1491
rect 863 -1492 864 -1368
rect 961 -1501 962 -1491
rect 1552 -1501 1553 -1491
rect 128 -1501 129 -1493
rect 1311 -1501 1312 -1493
rect 772 -1496 773 -1368
rect 863 -1501 864 -1495
rect 709 -1498 710 -1368
rect 772 -1501 773 -1497
rect 709 -1501 710 -1499
rect 866 -1501 867 -1499
rect 23 -1511 24 -1509
rect 229 -1511 230 -1509
rect 240 -1511 241 -1509
rect 320 -1511 321 -1509
rect 352 -1511 353 -1509
rect 352 -1636 353 -1510
rect 352 -1511 353 -1509
rect 352 -1636 353 -1510
rect 373 -1511 374 -1509
rect 376 -1519 377 -1510
rect 401 -1511 402 -1509
rect 457 -1511 458 -1509
rect 460 -1511 461 -1509
rect 1227 -1511 1228 -1509
rect 1248 -1511 1249 -1509
rect 1248 -1636 1249 -1510
rect 1248 -1511 1249 -1509
rect 1248 -1636 1249 -1510
rect 1374 -1511 1375 -1509
rect 1374 -1636 1375 -1510
rect 1374 -1511 1375 -1509
rect 1374 -1636 1375 -1510
rect 1437 -1511 1438 -1509
rect 1437 -1636 1438 -1510
rect 1437 -1511 1438 -1509
rect 1437 -1636 1438 -1510
rect 1451 -1511 1452 -1509
rect 1454 -1511 1455 -1509
rect 1486 -1511 1487 -1509
rect 1486 -1636 1487 -1510
rect 1486 -1511 1487 -1509
rect 1486 -1636 1487 -1510
rect 1521 -1511 1522 -1509
rect 1549 -1511 1550 -1509
rect 1584 -1511 1585 -1509
rect 1668 -1511 1669 -1509
rect 1706 -1636 1707 -1510
rect 1710 -1511 1711 -1509
rect 1801 -1511 1802 -1509
rect 1822 -1636 1823 -1510
rect 23 -1636 24 -1512
rect 418 -1513 419 -1509
rect 436 -1513 437 -1509
rect 761 -1513 762 -1509
rect 779 -1513 780 -1509
rect 828 -1636 829 -1512
rect 866 -1513 867 -1509
rect 1423 -1513 1424 -1509
rect 1451 -1636 1452 -1512
rect 1472 -1513 1473 -1509
rect 1521 -1636 1522 -1512
rect 1605 -1513 1606 -1509
rect 1619 -1513 1620 -1509
rect 1619 -1636 1620 -1512
rect 1619 -1513 1620 -1509
rect 1619 -1636 1620 -1512
rect 1640 -1513 1641 -1509
rect 1731 -1513 1732 -1509
rect 37 -1515 38 -1509
rect 726 -1515 727 -1509
rect 737 -1515 738 -1509
rect 1220 -1515 1221 -1509
rect 1227 -1636 1228 -1514
rect 1255 -1515 1256 -1509
rect 1304 -1515 1305 -1509
rect 1423 -1636 1424 -1514
rect 1528 -1515 1529 -1509
rect 1528 -1636 1529 -1514
rect 1528 -1515 1529 -1509
rect 1528 -1636 1529 -1514
rect 1535 -1515 1536 -1509
rect 1696 -1515 1697 -1509
rect 37 -1636 38 -1516
rect 65 -1517 66 -1509
rect 93 -1517 94 -1509
rect 317 -1636 318 -1516
rect 373 -1636 374 -1516
rect 492 -1517 493 -1509
rect 670 -1517 671 -1509
rect 681 -1517 682 -1509
rect 978 -1517 979 -1509
rect 1020 -1636 1021 -1516
rect 1465 -1517 1466 -1509
rect 1535 -1636 1536 -1516
rect 1542 -1517 1543 -1509
rect 1577 -1517 1578 -1509
rect 1584 -1636 1585 -1516
rect 1598 -1517 1599 -1509
rect 1696 -1636 1697 -1516
rect 51 -1519 52 -1509
rect 625 -1519 626 -1509
rect 646 -1519 647 -1509
rect 646 -1636 647 -1518
rect 646 -1519 647 -1509
rect 646 -1636 647 -1518
rect 688 -1519 689 -1509
rect 950 -1519 951 -1509
rect 961 -1519 962 -1509
rect 961 -1636 962 -1518
rect 961 -1519 962 -1509
rect 961 -1636 962 -1518
rect 1031 -1519 1032 -1509
rect 1199 -1519 1200 -1509
rect 1255 -1636 1256 -1518
rect 1262 -1519 1263 -1509
rect 1454 -1636 1455 -1518
rect 1472 -1636 1473 -1518
rect 1507 -1519 1508 -1509
rect 1542 -1636 1543 -1518
rect 1577 -1636 1578 -1518
rect 1612 -1519 1613 -1509
rect 1640 -1636 1641 -1518
rect 1647 -1519 1648 -1509
rect 1650 -1636 1651 -1518
rect 1724 -1519 1725 -1509
rect 51 -1636 52 -1520
rect 261 -1521 262 -1509
rect 264 -1636 265 -1520
rect 520 -1521 521 -1509
rect 527 -1521 528 -1509
rect 656 -1521 657 -1509
rect 695 -1521 696 -1509
rect 695 -1636 696 -1520
rect 695 -1521 696 -1509
rect 695 -1636 696 -1520
rect 716 -1521 717 -1509
rect 1262 -1636 1263 -1520
rect 1311 -1521 1312 -1509
rect 1507 -1636 1508 -1520
rect 1591 -1521 1592 -1509
rect 1598 -1636 1599 -1520
rect 1612 -1636 1613 -1520
rect 1626 -1521 1627 -1509
rect 1643 -1521 1644 -1509
rect 1710 -1636 1711 -1520
rect 1717 -1521 1718 -1509
rect 1724 -1636 1725 -1520
rect 58 -1523 59 -1509
rect 957 -1636 958 -1522
rect 989 -1523 990 -1509
rect 1031 -1636 1032 -1522
rect 1034 -1523 1035 -1509
rect 1108 -1523 1109 -1509
rect 1157 -1523 1158 -1509
rect 1199 -1636 1200 -1522
rect 1311 -1636 1312 -1522
rect 1318 -1523 1319 -1509
rect 1479 -1523 1480 -1509
rect 1591 -1636 1592 -1522
rect 1668 -1636 1669 -1522
rect 1682 -1523 1683 -1509
rect 1703 -1523 1704 -1509
rect 1717 -1636 1718 -1522
rect 65 -1636 66 -1524
rect 870 -1525 871 -1509
rect 880 -1636 881 -1524
rect 1017 -1525 1018 -1509
rect 1045 -1636 1046 -1524
rect 1066 -1525 1067 -1509
rect 1171 -1525 1172 -1509
rect 1171 -1636 1172 -1524
rect 1171 -1525 1172 -1509
rect 1171 -1636 1172 -1524
rect 1188 -1636 1189 -1524
rect 1458 -1525 1459 -1509
rect 1514 -1525 1515 -1509
rect 1626 -1636 1627 -1524
rect 1633 -1525 1634 -1509
rect 1682 -1636 1683 -1524
rect 93 -1636 94 -1526
rect 541 -1527 542 -1509
rect 607 -1636 608 -1526
rect 919 -1527 920 -1509
rect 936 -1527 937 -1509
rect 1185 -1527 1186 -1509
rect 1192 -1527 1193 -1509
rect 1220 -1636 1221 -1526
rect 1318 -1636 1319 -1526
rect 1647 -1636 1648 -1526
rect 124 -1529 125 -1509
rect 313 -1636 314 -1528
rect 380 -1529 381 -1509
rect 457 -1636 458 -1528
rect 481 -1529 482 -1509
rect 1608 -1529 1609 -1509
rect 44 -1531 45 -1509
rect 124 -1636 125 -1530
rect 128 -1531 129 -1509
rect 198 -1531 199 -1509
rect 212 -1531 213 -1509
rect 240 -1636 241 -1530
rect 303 -1531 304 -1509
rect 303 -1636 304 -1530
rect 303 -1531 304 -1509
rect 303 -1636 304 -1530
rect 310 -1531 311 -1509
rect 726 -1636 727 -1530
rect 737 -1636 738 -1530
rect 744 -1531 745 -1509
rect 747 -1636 748 -1530
rect 933 -1531 934 -1509
rect 947 -1531 948 -1509
rect 1234 -1531 1235 -1509
rect 1332 -1531 1333 -1509
rect 1514 -1636 1515 -1530
rect 1563 -1531 1564 -1509
rect 1633 -1636 1634 -1530
rect 44 -1636 45 -1532
rect 61 -1636 62 -1532
rect 79 -1533 80 -1509
rect 128 -1636 129 -1532
rect 131 -1533 132 -1509
rect 296 -1533 297 -1509
rect 415 -1533 416 -1509
rect 569 -1533 570 -1509
rect 611 -1533 612 -1509
rect 681 -1636 682 -1532
rect 702 -1533 703 -1509
rect 716 -1636 717 -1532
rect 723 -1636 724 -1532
rect 1360 -1533 1361 -1509
rect 1416 -1533 1417 -1509
rect 1479 -1636 1480 -1532
rect 1556 -1533 1557 -1509
rect 1563 -1636 1564 -1532
rect 79 -1636 80 -1534
rect 1006 -1636 1007 -1534
rect 1048 -1535 1049 -1509
rect 1283 -1535 1284 -1509
rect 1325 -1535 1326 -1509
rect 1332 -1636 1333 -1534
rect 1395 -1535 1396 -1509
rect 1416 -1636 1417 -1534
rect 1430 -1535 1431 -1509
rect 1458 -1636 1459 -1534
rect 1556 -1636 1557 -1534
rect 1570 -1535 1571 -1509
rect 149 -1537 150 -1509
rect 611 -1636 612 -1536
rect 625 -1636 626 -1536
rect 821 -1537 822 -1509
rect 831 -1537 832 -1509
rect 1605 -1636 1606 -1536
rect 135 -1539 136 -1509
rect 149 -1636 150 -1538
rect 156 -1539 157 -1509
rect 1549 -1636 1550 -1538
rect 159 -1541 160 -1509
rect 380 -1636 381 -1540
rect 415 -1636 416 -1540
rect 471 -1541 472 -1509
rect 506 -1541 507 -1509
rect 527 -1636 528 -1540
rect 569 -1636 570 -1540
rect 1654 -1541 1655 -1509
rect 177 -1543 178 -1509
rect 177 -1636 178 -1542
rect 177 -1543 178 -1509
rect 177 -1636 178 -1542
rect 184 -1543 185 -1509
rect 443 -1543 444 -1509
rect 506 -1636 507 -1542
rect 555 -1543 556 -1509
rect 604 -1543 605 -1509
rect 702 -1636 703 -1542
rect 709 -1543 710 -1509
rect 1066 -1636 1067 -1542
rect 1073 -1543 1074 -1509
rect 1192 -1636 1193 -1542
rect 1206 -1543 1207 -1509
rect 1283 -1636 1284 -1542
rect 1290 -1543 1291 -1509
rect 1325 -1636 1326 -1542
rect 1381 -1543 1382 -1509
rect 1395 -1636 1396 -1542
rect 1493 -1543 1494 -1509
rect 1570 -1636 1571 -1542
rect 1654 -1636 1655 -1542
rect 1661 -1543 1662 -1509
rect 184 -1636 185 -1544
rect 1430 -1636 1431 -1544
rect 1661 -1636 1662 -1544
rect 1675 -1545 1676 -1509
rect 191 -1547 192 -1509
rect 401 -1636 402 -1546
rect 422 -1547 423 -1509
rect 520 -1636 521 -1546
rect 544 -1636 545 -1546
rect 1381 -1636 1382 -1546
rect 1675 -1636 1676 -1546
rect 1689 -1547 1690 -1509
rect 86 -1549 87 -1509
rect 422 -1636 423 -1548
rect 436 -1636 437 -1548
rect 996 -1549 997 -1509
rect 1059 -1549 1060 -1509
rect 1073 -1636 1074 -1548
rect 1164 -1549 1165 -1509
rect 1234 -1636 1235 -1548
rect 1269 -1549 1270 -1509
rect 1290 -1636 1291 -1548
rect 1685 -1636 1686 -1548
rect 1689 -1636 1690 -1548
rect 68 -1551 69 -1509
rect 86 -1636 87 -1550
rect 191 -1636 192 -1550
rect 247 -1551 248 -1509
rect 387 -1551 388 -1509
rect 471 -1636 472 -1550
rect 478 -1551 479 -1509
rect 1493 -1636 1494 -1550
rect 194 -1553 195 -1509
rect 1465 -1636 1466 -1552
rect 198 -1636 199 -1554
rect 450 -1555 451 -1509
rect 653 -1555 654 -1509
rect 919 -1636 920 -1554
rect 947 -1636 948 -1554
rect 1538 -1555 1539 -1509
rect 205 -1557 206 -1509
rect 933 -1636 934 -1556
rect 968 -1557 969 -1509
rect 989 -1636 990 -1556
rect 996 -1636 997 -1556
rect 1122 -1557 1123 -1509
rect 1178 -1557 1179 -1509
rect 1269 -1636 1270 -1556
rect 121 -1559 122 -1509
rect 205 -1636 206 -1558
rect 212 -1636 213 -1558
rect 324 -1559 325 -1509
rect 387 -1636 388 -1558
rect 464 -1559 465 -1509
rect 541 -1636 542 -1558
rect 1122 -1636 1123 -1558
rect 1136 -1559 1137 -1509
rect 1178 -1636 1179 -1558
rect 1185 -1636 1186 -1558
rect 1304 -1636 1305 -1558
rect 121 -1636 122 -1560
rect 156 -1636 157 -1560
rect 215 -1561 216 -1509
rect 408 -1561 409 -1509
rect 443 -1636 444 -1560
rect 562 -1561 563 -1509
rect 632 -1561 633 -1509
rect 968 -1636 969 -1560
rect 1062 -1636 1063 -1560
rect 1444 -1561 1445 -1509
rect 219 -1563 220 -1509
rect 688 -1636 689 -1562
rect 709 -1636 710 -1562
rect 835 -1563 836 -1509
rect 863 -1563 864 -1509
rect 1360 -1636 1361 -1562
rect 1367 -1563 1368 -1509
rect 1444 -1636 1445 -1562
rect 30 -1565 31 -1509
rect 219 -1636 220 -1564
rect 222 -1636 223 -1564
rect 733 -1636 734 -1564
rect 740 -1565 741 -1509
rect 1101 -1565 1102 -1509
rect 1136 -1636 1137 -1564
rect 1143 -1565 1144 -1509
rect 1346 -1565 1347 -1509
rect 1367 -1636 1368 -1564
rect 30 -1636 31 -1566
rect 628 -1567 629 -1509
rect 653 -1636 654 -1566
rect 674 -1567 675 -1509
rect 754 -1636 755 -1566
rect 1052 -1567 1053 -1509
rect 1101 -1636 1102 -1566
rect 1150 -1567 1151 -1509
rect 1346 -1636 1347 -1566
rect 1402 -1567 1403 -1509
rect 233 -1569 234 -1509
rect 296 -1636 297 -1568
rect 324 -1636 325 -1568
rect 817 -1636 818 -1568
rect 863 -1636 864 -1568
rect 1157 -1636 1158 -1568
rect 1388 -1569 1389 -1509
rect 1402 -1636 1403 -1568
rect 233 -1636 234 -1570
rect 429 -1571 430 -1509
rect 446 -1636 447 -1570
rect 478 -1636 479 -1570
rect 499 -1571 500 -1509
rect 632 -1636 633 -1570
rect 667 -1571 668 -1509
rect 1164 -1636 1165 -1570
rect 1388 -1636 1389 -1570
rect 1500 -1571 1501 -1509
rect 247 -1636 248 -1572
rect 310 -1636 311 -1572
rect 429 -1636 430 -1572
rect 821 -1636 822 -1572
rect 870 -1636 871 -1572
rect 1003 -1573 1004 -1509
rect 1094 -1573 1095 -1509
rect 1150 -1636 1151 -1572
rect 1409 -1573 1410 -1509
rect 1500 -1636 1501 -1572
rect 275 -1575 276 -1509
rect 408 -1636 409 -1574
rect 464 -1636 465 -1574
rect 604 -1636 605 -1574
rect 758 -1575 759 -1509
rect 856 -1575 857 -1509
rect 894 -1636 895 -1574
rect 1241 -1575 1242 -1509
rect 1353 -1575 1354 -1509
rect 1409 -1636 1410 -1574
rect 142 -1577 143 -1509
rect 275 -1636 276 -1576
rect 499 -1636 500 -1576
rect 639 -1577 640 -1509
rect 730 -1577 731 -1509
rect 758 -1636 759 -1576
rect 779 -1636 780 -1576
rect 1017 -1636 1018 -1576
rect 1094 -1636 1095 -1576
rect 1129 -1577 1130 -1509
rect 1297 -1577 1298 -1509
rect 1353 -1636 1354 -1576
rect 142 -1636 143 -1578
rect 163 -1579 164 -1509
rect 548 -1579 549 -1509
rect 667 -1636 668 -1578
rect 730 -1636 731 -1578
rect 1339 -1579 1340 -1509
rect 163 -1636 164 -1580
rect 1241 -1636 1242 -1580
rect 1297 -1636 1298 -1580
rect 1339 -1636 1340 -1580
rect 548 -1636 549 -1582
rect 583 -1583 584 -1509
rect 590 -1583 591 -1509
rect 674 -1636 675 -1582
rect 786 -1583 787 -1509
rect 926 -1583 927 -1509
rect 940 -1583 941 -1509
rect 1003 -1636 1004 -1582
rect 1115 -1583 1116 -1509
rect 1129 -1636 1130 -1582
rect 187 -1636 188 -1584
rect 590 -1636 591 -1584
rect 639 -1636 640 -1584
rect 891 -1585 892 -1509
rect 905 -1585 906 -1509
rect 905 -1636 906 -1584
rect 905 -1585 906 -1509
rect 905 -1636 906 -1584
rect 912 -1585 913 -1509
rect 926 -1636 927 -1584
rect 940 -1636 941 -1584
rect 1080 -1585 1081 -1509
rect 1087 -1585 1088 -1509
rect 1115 -1636 1116 -1584
rect 1125 -1636 1126 -1584
rect 1143 -1636 1144 -1584
rect 492 -1636 493 -1586
rect 891 -1636 892 -1586
rect 898 -1587 899 -1509
rect 912 -1636 913 -1586
rect 975 -1587 976 -1509
rect 1052 -1636 1053 -1586
rect 1080 -1636 1081 -1586
rect 1206 -1636 1207 -1586
rect 562 -1636 563 -1588
rect 576 -1589 577 -1509
rect 583 -1636 584 -1588
rect 660 -1589 661 -1509
rect 786 -1636 787 -1588
rect 824 -1589 825 -1509
rect 884 -1589 885 -1509
rect 898 -1636 899 -1588
rect 954 -1589 955 -1509
rect 975 -1636 976 -1588
rect 1024 -1589 1025 -1509
rect 1087 -1636 1088 -1588
rect 135 -1636 136 -1590
rect 824 -1636 825 -1590
rect 849 -1591 850 -1509
rect 884 -1636 885 -1590
rect 954 -1636 955 -1590
rect 1276 -1591 1277 -1509
rect 450 -1636 451 -1592
rect 849 -1636 850 -1592
rect 1010 -1593 1011 -1509
rect 1024 -1636 1025 -1592
rect 1213 -1593 1214 -1509
rect 1276 -1636 1277 -1592
rect 551 -1636 552 -1594
rect 1213 -1636 1214 -1594
rect 576 -1636 577 -1596
rect 765 -1597 766 -1509
rect 789 -1597 790 -1509
rect 842 -1597 843 -1509
rect 982 -1597 983 -1509
rect 1010 -1636 1011 -1596
rect 597 -1599 598 -1509
rect 660 -1636 661 -1598
rect 800 -1599 801 -1509
rect 835 -1636 836 -1598
rect 982 -1636 983 -1598
rect 1038 -1599 1039 -1509
rect 72 -1601 73 -1509
rect 1038 -1636 1039 -1600
rect 72 -1636 73 -1602
rect 254 -1603 255 -1509
rect 618 -1603 619 -1509
rect 765 -1636 766 -1602
rect 793 -1603 794 -1509
rect 800 -1636 801 -1602
rect 807 -1603 808 -1509
rect 866 -1636 867 -1602
rect 100 -1605 101 -1509
rect 618 -1636 619 -1604
rect 772 -1605 773 -1509
rect 793 -1636 794 -1604
rect 814 -1605 815 -1509
rect 842 -1636 843 -1604
rect 100 -1636 101 -1606
rect 226 -1607 227 -1509
rect 513 -1607 514 -1509
rect 807 -1636 808 -1606
rect 114 -1609 115 -1509
rect 226 -1636 227 -1608
rect 359 -1609 360 -1509
rect 513 -1636 514 -1608
rect 555 -1636 556 -1608
rect 814 -1636 815 -1608
rect 114 -1636 115 -1610
rect 331 -1611 332 -1509
rect 359 -1636 360 -1610
rect 366 -1611 367 -1509
rect 751 -1611 752 -1509
rect 772 -1636 773 -1610
rect 166 -1636 167 -1612
rect 254 -1636 255 -1612
rect 366 -1636 367 -1612
rect 751 -1636 752 -1612
rect 170 -1615 171 -1509
rect 597 -1636 598 -1614
rect 170 -1636 171 -1616
rect 289 -1617 290 -1509
rect 107 -1619 108 -1509
rect 289 -1636 290 -1618
rect 107 -1636 108 -1620
rect 394 -1621 395 -1509
rect 268 -1623 269 -1509
rect 394 -1636 395 -1622
rect 268 -1636 269 -1624
rect 282 -1625 283 -1509
rect 282 -1636 283 -1626
rect 338 -1627 339 -1509
rect 338 -1636 339 -1628
rect 345 -1629 346 -1509
rect 345 -1636 346 -1630
rect 534 -1631 535 -1509
rect 534 -1636 535 -1632
rect 877 -1633 878 -1509
rect 331 -1636 332 -1634
rect 877 -1636 878 -1634
rect 30 -1646 31 -1644
rect 310 -1646 311 -1644
rect 324 -1646 325 -1644
rect 383 -1783 384 -1645
rect 387 -1646 388 -1644
rect 607 -1646 608 -1644
rect 660 -1646 661 -1644
rect 733 -1646 734 -1644
rect 789 -1783 790 -1645
rect 1297 -1783 1298 -1645
rect 1300 -1646 1301 -1644
rect 1458 -1646 1459 -1644
rect 1549 -1646 1550 -1644
rect 1703 -1783 1704 -1645
rect 1822 -1646 1823 -1644
rect 1839 -1783 1840 -1645
rect 30 -1783 31 -1647
rect 198 -1648 199 -1644
rect 219 -1648 220 -1644
rect 502 -1783 503 -1647
rect 548 -1648 549 -1644
rect 1710 -1648 1711 -1644
rect 23 -1650 24 -1644
rect 198 -1783 199 -1649
rect 236 -1783 237 -1649
rect 1794 -1783 1795 -1649
rect 23 -1783 24 -1651
rect 233 -1652 234 -1644
rect 275 -1652 276 -1644
rect 310 -1783 311 -1651
rect 338 -1652 339 -1644
rect 338 -1783 339 -1651
rect 338 -1652 339 -1644
rect 338 -1783 339 -1651
rect 345 -1652 346 -1644
rect 345 -1783 346 -1651
rect 345 -1652 346 -1644
rect 345 -1783 346 -1651
rect 352 -1652 353 -1644
rect 450 -1652 451 -1644
rect 551 -1652 552 -1644
rect 1115 -1652 1116 -1644
rect 1122 -1652 1123 -1644
rect 1458 -1783 1459 -1651
rect 1598 -1652 1599 -1644
rect 1731 -1783 1732 -1651
rect 58 -1783 59 -1653
rect 730 -1654 731 -1644
rect 800 -1654 801 -1644
rect 817 -1654 818 -1644
rect 856 -1783 857 -1653
rect 884 -1654 885 -1644
rect 891 -1654 892 -1644
rect 1787 -1783 1788 -1653
rect 107 -1656 108 -1644
rect 891 -1783 892 -1655
rect 954 -1783 955 -1655
rect 1111 -1656 1112 -1644
rect 1125 -1656 1126 -1644
rect 1255 -1656 1256 -1644
rect 1423 -1656 1424 -1644
rect 1549 -1783 1550 -1655
rect 1605 -1656 1606 -1644
rect 1745 -1783 1746 -1655
rect 93 -1658 94 -1644
rect 107 -1783 108 -1657
rect 121 -1658 122 -1644
rect 1171 -1658 1172 -1644
rect 1185 -1658 1186 -1644
rect 1836 -1783 1837 -1657
rect 93 -1783 94 -1659
rect 537 -1783 538 -1659
rect 576 -1660 577 -1644
rect 800 -1783 801 -1659
rect 814 -1660 815 -1644
rect 1640 -1660 1641 -1644
rect 1647 -1660 1648 -1644
rect 1780 -1783 1781 -1659
rect 121 -1783 122 -1661
rect 719 -1783 720 -1661
rect 782 -1783 783 -1661
rect 1605 -1783 1606 -1661
rect 1619 -1662 1620 -1644
rect 1752 -1783 1753 -1661
rect 124 -1664 125 -1644
rect 887 -1783 888 -1663
rect 957 -1664 958 -1644
rect 1738 -1783 1739 -1663
rect 135 -1666 136 -1644
rect 677 -1783 678 -1665
rect 681 -1666 682 -1644
rect 751 -1666 752 -1644
rect 835 -1666 836 -1644
rect 1171 -1783 1172 -1665
rect 1185 -1783 1186 -1665
rect 1234 -1666 1235 -1644
rect 1304 -1666 1305 -1644
rect 1423 -1783 1424 -1665
rect 1451 -1666 1452 -1644
rect 1710 -1783 1711 -1665
rect 135 -1783 136 -1667
rect 1062 -1668 1063 -1644
rect 1066 -1668 1067 -1644
rect 1083 -1668 1084 -1644
rect 1101 -1668 1102 -1644
rect 1255 -1783 1256 -1667
rect 1332 -1668 1333 -1644
rect 1451 -1783 1452 -1667
rect 1479 -1668 1480 -1644
rect 1619 -1783 1620 -1667
rect 1626 -1668 1627 -1644
rect 1759 -1783 1760 -1667
rect 159 -1783 160 -1669
rect 579 -1783 580 -1669
rect 590 -1670 591 -1644
rect 751 -1783 752 -1669
rect 835 -1783 836 -1669
rect 849 -1670 850 -1644
rect 859 -1670 860 -1644
rect 996 -1670 997 -1644
rect 1003 -1670 1004 -1644
rect 1563 -1670 1564 -1644
rect 1633 -1670 1634 -1644
rect 1766 -1783 1767 -1669
rect 184 -1672 185 -1644
rect 212 -1672 213 -1644
rect 275 -1783 276 -1671
rect 520 -1672 521 -1644
rect 604 -1783 605 -1671
rect 726 -1672 727 -1644
rect 863 -1672 864 -1644
rect 1087 -1672 1088 -1644
rect 1101 -1783 1102 -1671
rect 1689 -1672 1690 -1644
rect 1696 -1672 1697 -1644
rect 1829 -1783 1830 -1671
rect 145 -1783 146 -1673
rect 184 -1783 185 -1673
rect 187 -1674 188 -1644
rect 534 -1674 535 -1644
rect 611 -1674 612 -1644
rect 660 -1783 661 -1673
rect 674 -1674 675 -1644
rect 814 -1783 815 -1673
rect 828 -1674 829 -1644
rect 863 -1783 864 -1673
rect 877 -1674 878 -1644
rect 1360 -1674 1361 -1644
rect 1374 -1674 1375 -1644
rect 1479 -1783 1480 -1673
rect 1521 -1674 1522 -1644
rect 1640 -1783 1641 -1673
rect 1650 -1674 1651 -1644
rect 1724 -1674 1725 -1644
rect 44 -1676 45 -1644
rect 674 -1783 675 -1675
rect 681 -1783 682 -1675
rect 779 -1676 780 -1644
rect 786 -1676 787 -1644
rect 828 -1783 829 -1675
rect 877 -1783 878 -1675
rect 905 -1676 906 -1644
rect 950 -1783 951 -1675
rect 1633 -1783 1634 -1675
rect 1654 -1676 1655 -1644
rect 1808 -1783 1809 -1675
rect 44 -1783 45 -1677
rect 639 -1678 640 -1644
rect 716 -1678 717 -1644
rect 730 -1783 731 -1677
rect 779 -1783 780 -1677
rect 824 -1678 825 -1644
rect 880 -1678 881 -1644
rect 1325 -1678 1326 -1644
rect 1395 -1678 1396 -1644
rect 1521 -1783 1522 -1677
rect 1528 -1678 1529 -1644
rect 1689 -1783 1690 -1677
rect 212 -1783 213 -1679
rect 555 -1680 556 -1644
rect 611 -1783 612 -1679
rect 842 -1680 843 -1644
rect 901 -1783 902 -1679
rect 996 -1783 997 -1679
rect 1017 -1680 1018 -1644
rect 1129 -1680 1130 -1644
rect 1146 -1783 1147 -1679
rect 1577 -1680 1578 -1644
rect 1584 -1680 1585 -1644
rect 1724 -1783 1725 -1679
rect 282 -1682 283 -1644
rect 282 -1783 283 -1681
rect 282 -1682 283 -1644
rect 282 -1783 283 -1681
rect 303 -1682 304 -1644
rect 324 -1783 325 -1681
rect 352 -1783 353 -1681
rect 544 -1682 545 -1644
rect 618 -1682 619 -1644
rect 905 -1783 906 -1681
rect 947 -1682 948 -1644
rect 1017 -1783 1018 -1681
rect 1020 -1682 1021 -1644
rect 1234 -1783 1235 -1681
rect 1262 -1682 1263 -1644
rect 1325 -1783 1326 -1681
rect 1402 -1682 1403 -1644
rect 1528 -1783 1529 -1681
rect 1542 -1682 1543 -1644
rect 1696 -1783 1697 -1681
rect 205 -1684 206 -1644
rect 1402 -1783 1403 -1683
rect 1416 -1684 1417 -1644
rect 1542 -1783 1543 -1683
rect 1661 -1684 1662 -1644
rect 1801 -1783 1802 -1683
rect 37 -1686 38 -1644
rect 1661 -1783 1662 -1685
rect 1668 -1686 1669 -1644
rect 1815 -1783 1816 -1685
rect 37 -1783 38 -1687
rect 506 -1688 507 -1644
rect 534 -1783 535 -1687
rect 1087 -1783 1088 -1687
rect 1108 -1688 1109 -1644
rect 1591 -1688 1592 -1644
rect 1675 -1688 1676 -1644
rect 1822 -1783 1823 -1687
rect 79 -1690 80 -1644
rect 205 -1783 206 -1689
rect 254 -1690 255 -1644
rect 303 -1783 304 -1689
rect 331 -1690 332 -1644
rect 618 -1783 619 -1689
rect 639 -1783 640 -1689
rect 646 -1690 647 -1644
rect 716 -1783 717 -1689
rect 1031 -1690 1032 -1644
rect 1038 -1690 1039 -1644
rect 1598 -1783 1599 -1689
rect 1682 -1690 1683 -1644
rect 1717 -1690 1718 -1644
rect 79 -1783 80 -1691
rect 366 -1692 367 -1644
rect 387 -1783 388 -1691
rect 492 -1692 493 -1644
rect 499 -1692 500 -1644
rect 520 -1783 521 -1691
rect 646 -1783 647 -1691
rect 653 -1692 654 -1644
rect 723 -1783 724 -1691
rect 1066 -1783 1067 -1691
rect 1080 -1692 1081 -1644
rect 1416 -1783 1417 -1691
rect 1437 -1692 1438 -1644
rect 1563 -1783 1564 -1691
rect 1570 -1692 1571 -1644
rect 1591 -1783 1592 -1691
rect 254 -1783 255 -1693
rect 464 -1694 465 -1644
rect 485 -1694 486 -1644
rect 544 -1783 545 -1693
rect 632 -1694 633 -1644
rect 653 -1783 654 -1693
rect 747 -1694 748 -1644
rect 1395 -1783 1396 -1693
rect 1444 -1694 1445 -1644
rect 1584 -1783 1585 -1693
rect 331 -1783 332 -1695
rect 359 -1696 360 -1644
rect 362 -1783 363 -1695
rect 1003 -1783 1004 -1695
rect 1010 -1696 1011 -1644
rect 1080 -1783 1081 -1695
rect 1129 -1783 1130 -1695
rect 1248 -1696 1249 -1644
rect 1269 -1696 1270 -1644
rect 1332 -1783 1333 -1695
rect 1388 -1696 1389 -1644
rect 1675 -1783 1676 -1695
rect 366 -1783 367 -1697
rect 380 -1698 381 -1644
rect 394 -1698 395 -1644
rect 593 -1783 594 -1697
rect 807 -1698 808 -1644
rect 842 -1783 843 -1697
rect 975 -1698 976 -1644
rect 1031 -1783 1032 -1697
rect 1038 -1783 1039 -1697
rect 1059 -1698 1060 -1644
rect 1136 -1698 1137 -1644
rect 1269 -1783 1270 -1697
rect 1290 -1698 1291 -1644
rect 1388 -1783 1389 -1697
rect 1472 -1698 1473 -1644
rect 1626 -1783 1627 -1697
rect 394 -1783 395 -1699
rect 597 -1700 598 -1644
rect 754 -1700 755 -1644
rect 1136 -1783 1137 -1699
rect 1157 -1700 1158 -1644
rect 1444 -1783 1445 -1699
rect 1493 -1700 1494 -1644
rect 1654 -1783 1655 -1699
rect 401 -1702 402 -1644
rect 597 -1783 598 -1701
rect 726 -1783 727 -1701
rect 1493 -1783 1494 -1701
rect 1500 -1702 1501 -1644
rect 1577 -1783 1578 -1701
rect 240 -1704 241 -1644
rect 401 -1783 402 -1703
rect 408 -1704 409 -1644
rect 551 -1783 552 -1703
rect 765 -1704 766 -1644
rect 807 -1783 808 -1703
rect 824 -1783 825 -1703
rect 968 -1704 969 -1644
rect 978 -1783 979 -1703
rect 1647 -1783 1648 -1703
rect 114 -1706 115 -1644
rect 240 -1783 241 -1705
rect 408 -1783 409 -1705
rect 884 -1783 885 -1705
rect 898 -1706 899 -1644
rect 968 -1783 969 -1705
rect 989 -1706 990 -1644
rect 1108 -1783 1109 -1705
rect 1157 -1783 1158 -1705
rect 1318 -1706 1319 -1644
rect 1339 -1706 1340 -1644
rect 1472 -1783 1473 -1705
rect 1507 -1706 1508 -1644
rect 1570 -1783 1571 -1705
rect 415 -1708 416 -1644
rect 450 -1783 451 -1707
rect 457 -1708 458 -1644
rect 492 -1783 493 -1707
rect 506 -1783 507 -1707
rect 541 -1708 542 -1644
rect 758 -1708 759 -1644
rect 765 -1783 766 -1707
rect 919 -1708 920 -1644
rect 989 -1783 990 -1707
rect 1010 -1783 1011 -1707
rect 1143 -1708 1144 -1644
rect 1164 -1708 1165 -1644
rect 1248 -1783 1249 -1707
rect 1276 -1708 1277 -1644
rect 1339 -1783 1340 -1707
rect 1381 -1708 1382 -1644
rect 1500 -1783 1501 -1707
rect 1514 -1708 1515 -1644
rect 1668 -1783 1669 -1707
rect 219 -1783 220 -1709
rect 1514 -1783 1515 -1709
rect 1535 -1710 1536 -1644
rect 1682 -1783 1683 -1709
rect 415 -1783 416 -1711
rect 576 -1783 577 -1711
rect 635 -1783 636 -1711
rect 1381 -1783 1382 -1711
rect 1409 -1712 1410 -1644
rect 1535 -1783 1536 -1711
rect 1556 -1712 1557 -1644
rect 1717 -1783 1718 -1711
rect 429 -1714 430 -1644
rect 1304 -1783 1305 -1713
rect 1311 -1714 1312 -1644
rect 1507 -1783 1508 -1713
rect 436 -1716 437 -1644
rect 744 -1716 745 -1644
rect 758 -1783 759 -1715
rect 772 -1716 773 -1644
rect 786 -1783 787 -1715
rect 1276 -1783 1277 -1715
rect 1430 -1716 1431 -1644
rect 1556 -1783 1557 -1715
rect 114 -1783 115 -1717
rect 772 -1783 773 -1717
rect 849 -1783 850 -1717
rect 1143 -1783 1144 -1717
rect 1178 -1718 1179 -1644
rect 1311 -1783 1312 -1717
rect 1367 -1718 1368 -1644
rect 1430 -1783 1431 -1717
rect 436 -1783 437 -1719
rect 569 -1720 570 -1644
rect 695 -1720 696 -1644
rect 744 -1783 745 -1719
rect 870 -1720 871 -1644
rect 919 -1783 920 -1719
rect 933 -1720 934 -1644
rect 1059 -1783 1060 -1719
rect 1206 -1720 1207 -1644
rect 1612 -1720 1613 -1644
rect 89 -1783 90 -1721
rect 1206 -1783 1207 -1721
rect 1220 -1722 1221 -1644
rect 1318 -1783 1319 -1721
rect 1353 -1722 1354 -1644
rect 1612 -1783 1613 -1721
rect 443 -1724 444 -1644
rect 443 -1783 444 -1723
rect 443 -1724 444 -1644
rect 443 -1783 444 -1723
rect 446 -1724 447 -1644
rect 513 -1724 514 -1644
rect 541 -1783 542 -1723
rect 555 -1783 556 -1723
rect 562 -1724 563 -1644
rect 569 -1783 570 -1723
rect 695 -1783 696 -1723
rect 793 -1724 794 -1644
rect 870 -1783 871 -1723
rect 947 -1783 948 -1723
rect 1006 -1724 1007 -1644
rect 1409 -1783 1410 -1723
rect 317 -1726 318 -1644
rect 793 -1783 794 -1725
rect 933 -1783 934 -1725
rect 961 -1726 962 -1644
rect 1024 -1726 1025 -1644
rect 1374 -1783 1375 -1725
rect 268 -1728 269 -1644
rect 1024 -1783 1025 -1727
rect 1027 -1783 1028 -1727
rect 1122 -1783 1123 -1727
rect 1227 -1728 1228 -1644
rect 1367 -1783 1368 -1727
rect 268 -1783 269 -1729
rect 548 -1783 549 -1729
rect 562 -1783 563 -1729
rect 898 -1783 899 -1729
rect 940 -1730 941 -1644
rect 1178 -1783 1179 -1729
rect 1241 -1730 1242 -1644
rect 1262 -1783 1263 -1729
rect 1283 -1730 1284 -1644
rect 1353 -1783 1354 -1729
rect 100 -1732 101 -1644
rect 1241 -1783 1242 -1731
rect 100 -1783 101 -1733
rect 170 -1734 171 -1644
rect 261 -1734 262 -1644
rect 940 -1783 941 -1733
rect 1045 -1734 1046 -1644
rect 1164 -1783 1165 -1733
rect 1213 -1734 1214 -1644
rect 1283 -1783 1284 -1733
rect 317 -1783 318 -1735
rect 1209 -1736 1210 -1644
rect 453 -1738 454 -1644
rect 1220 -1783 1221 -1737
rect 457 -1783 458 -1739
rect 478 -1740 479 -1644
rect 485 -1783 486 -1739
rect 527 -1740 528 -1644
rect 1045 -1783 1046 -1739
rect 1199 -1740 1200 -1644
rect 163 -1742 164 -1644
rect 1199 -1783 1200 -1741
rect 163 -1783 164 -1743
rect 191 -1744 192 -1644
rect 289 -1744 290 -1644
rect 527 -1783 528 -1743
rect 1052 -1744 1053 -1644
rect 1115 -1783 1116 -1743
rect 1150 -1744 1151 -1644
rect 1213 -1783 1214 -1743
rect 156 -1746 157 -1644
rect 191 -1783 192 -1745
rect 222 -1746 223 -1644
rect 289 -1783 290 -1745
rect 464 -1783 465 -1745
rect 471 -1746 472 -1644
rect 478 -1783 479 -1745
rect 583 -1746 584 -1644
rect 982 -1746 983 -1644
rect 1150 -1783 1151 -1745
rect 156 -1783 157 -1747
rect 429 -1783 430 -1747
rect 471 -1783 472 -1747
rect 625 -1748 626 -1644
rect 912 -1748 913 -1644
rect 982 -1783 983 -1747
rect 1052 -1783 1053 -1747
rect 1486 -1748 1487 -1644
rect 170 -1783 171 -1749
rect 222 -1783 223 -1749
rect 499 -1783 500 -1749
rect 961 -1783 962 -1749
rect 1055 -1783 1056 -1749
rect 1360 -1783 1361 -1749
rect 1465 -1750 1466 -1644
rect 1486 -1783 1487 -1749
rect 513 -1783 514 -1751
rect 667 -1752 668 -1644
rect 702 -1752 703 -1644
rect 912 -1783 913 -1751
rect 1094 -1752 1095 -1644
rect 1227 -1783 1228 -1751
rect 1346 -1752 1347 -1644
rect 1465 -1783 1466 -1751
rect 296 -1754 297 -1644
rect 1094 -1783 1095 -1753
rect 1192 -1754 1193 -1644
rect 1346 -1783 1347 -1753
rect 226 -1756 227 -1644
rect 296 -1783 297 -1755
rect 422 -1756 423 -1644
rect 702 -1783 703 -1755
rect 1073 -1756 1074 -1644
rect 1192 -1783 1193 -1755
rect 51 -1758 52 -1644
rect 226 -1783 227 -1757
rect 422 -1783 423 -1757
rect 737 -1758 738 -1644
rect 51 -1783 52 -1759
rect 926 -1760 927 -1644
rect 65 -1762 66 -1644
rect 926 -1783 927 -1761
rect 65 -1783 66 -1763
rect 373 -1764 374 -1644
rect 583 -1783 584 -1763
rect 1437 -1783 1438 -1763
rect 247 -1766 248 -1644
rect 373 -1783 374 -1765
rect 625 -1783 626 -1765
rect 1685 -1766 1686 -1644
rect 72 -1768 73 -1644
rect 247 -1783 248 -1767
rect 667 -1783 668 -1767
rect 705 -1783 706 -1767
rect 709 -1768 710 -1644
rect 1073 -1783 1074 -1767
rect 72 -1783 73 -1769
rect 1773 -1783 1774 -1769
rect 688 -1772 689 -1644
rect 737 -1783 738 -1771
rect 128 -1774 129 -1644
rect 688 -1783 689 -1773
rect 709 -1783 710 -1773
rect 866 -1774 867 -1644
rect 86 -1776 87 -1644
rect 128 -1783 129 -1775
rect 86 -1783 87 -1777
rect 149 -1778 150 -1644
rect 149 -1783 150 -1779
rect 177 -1780 178 -1644
rect 142 -1782 143 -1644
rect 177 -1783 178 -1781
rect 37 -1793 38 -1791
rect 537 -1793 538 -1791
rect 541 -1922 542 -1792
rect 684 -1922 685 -1792
rect 695 -1793 696 -1791
rect 915 -1922 916 -1792
rect 947 -1793 948 -1791
rect 1206 -1793 1207 -1791
rect 1230 -1922 1231 -1792
rect 1640 -1793 1641 -1791
rect 37 -1922 38 -1794
rect 611 -1795 612 -1791
rect 621 -1922 622 -1794
rect 1087 -1795 1088 -1791
rect 1143 -1922 1144 -1794
rect 1192 -1795 1193 -1791
rect 1395 -1795 1396 -1791
rect 1755 -1922 1756 -1794
rect 30 -1797 31 -1791
rect 611 -1922 612 -1796
rect 635 -1797 636 -1791
rect 646 -1797 647 -1791
rect 656 -1922 657 -1796
rect 891 -1797 892 -1791
rect 898 -1797 899 -1791
rect 1213 -1797 1214 -1791
rect 1423 -1797 1424 -1791
rect 1426 -1797 1427 -1791
rect 1451 -1797 1452 -1791
rect 1451 -1922 1452 -1796
rect 1451 -1797 1452 -1791
rect 1451 -1922 1452 -1796
rect 1563 -1797 1564 -1791
rect 1563 -1922 1564 -1796
rect 1563 -1797 1564 -1791
rect 1563 -1922 1564 -1796
rect 1640 -1922 1641 -1796
rect 1829 -1797 1830 -1791
rect 30 -1922 31 -1798
rect 93 -1799 94 -1791
rect 100 -1799 101 -1791
rect 117 -1799 118 -1791
rect 142 -1922 143 -1798
rect 1052 -1799 1053 -1791
rect 1192 -1922 1193 -1798
rect 1325 -1799 1326 -1791
rect 1423 -1922 1424 -1798
rect 1535 -1799 1536 -1791
rect 65 -1801 66 -1791
rect 264 -1801 265 -1791
rect 268 -1801 269 -1791
rect 646 -1922 647 -1800
rect 674 -1801 675 -1791
rect 695 -1922 696 -1800
rect 716 -1801 717 -1791
rect 1444 -1801 1445 -1791
rect 68 -1922 69 -1802
rect 373 -1803 374 -1791
rect 387 -1803 388 -1791
rect 387 -1922 388 -1802
rect 387 -1803 388 -1791
rect 387 -1922 388 -1802
rect 394 -1803 395 -1791
rect 502 -1803 503 -1791
rect 548 -1803 549 -1791
rect 1178 -1803 1179 -1791
rect 1213 -1922 1214 -1802
rect 1283 -1803 1284 -1791
rect 1325 -1922 1326 -1802
rect 1493 -1803 1494 -1791
rect 72 -1805 73 -1791
rect 128 -1805 129 -1791
rect 145 -1805 146 -1791
rect 359 -1805 360 -1791
rect 373 -1922 374 -1804
rect 709 -1805 710 -1791
rect 723 -1922 724 -1804
rect 992 -1922 993 -1804
rect 1024 -1805 1025 -1791
rect 1689 -1805 1690 -1791
rect 72 -1922 73 -1806
rect 457 -1807 458 -1791
rect 499 -1807 500 -1791
rect 1101 -1807 1102 -1791
rect 1178 -1922 1179 -1806
rect 1227 -1807 1228 -1791
rect 1234 -1807 1235 -1791
rect 1493 -1922 1494 -1806
rect 1689 -1922 1690 -1806
rect 1787 -1807 1788 -1791
rect 75 -1809 76 -1791
rect 814 -1809 815 -1791
rect 821 -1809 822 -1791
rect 835 -1809 836 -1791
rect 884 -1809 885 -1791
rect 1668 -1809 1669 -1791
rect 79 -1811 80 -1791
rect 82 -1833 83 -1810
rect 89 -1811 90 -1791
rect 177 -1811 178 -1791
rect 184 -1811 185 -1791
rect 236 -1811 237 -1791
rect 250 -1922 251 -1810
rect 457 -1922 458 -1810
rect 548 -1922 549 -1810
rect 597 -1811 598 -1791
rect 674 -1922 675 -1810
rect 772 -1811 773 -1791
rect 782 -1811 783 -1791
rect 1794 -1811 1795 -1791
rect 58 -1813 59 -1791
rect 177 -1922 178 -1812
rect 184 -1922 185 -1812
rect 317 -1813 318 -1791
rect 338 -1813 339 -1791
rect 432 -1922 433 -1812
rect 576 -1922 577 -1812
rect 667 -1813 668 -1791
rect 677 -1813 678 -1791
rect 1066 -1813 1067 -1791
rect 1101 -1922 1102 -1812
rect 1164 -1813 1165 -1791
rect 1283 -1922 1284 -1812
rect 1332 -1813 1333 -1791
rect 1444 -1922 1445 -1812
rect 1724 -1813 1725 -1791
rect 1794 -1922 1795 -1812
rect 1836 -1813 1837 -1791
rect 58 -1922 59 -1814
rect 1661 -1815 1662 -1791
rect 1668 -1922 1669 -1814
rect 1745 -1815 1746 -1791
rect 79 -1922 80 -1816
rect 443 -1817 444 -1791
rect 583 -1817 584 -1791
rect 625 -1817 626 -1791
rect 726 -1817 727 -1791
rect 1227 -1922 1228 -1816
rect 1332 -1922 1333 -1816
rect 1381 -1817 1382 -1791
rect 1661 -1922 1662 -1816
rect 1738 -1817 1739 -1791
rect 1745 -1922 1746 -1816
rect 1815 -1817 1816 -1791
rect 93 -1922 94 -1818
rect 478 -1819 479 -1791
rect 534 -1819 535 -1791
rect 583 -1922 584 -1818
rect 597 -1922 598 -1818
rect 772 -1922 773 -1818
rect 786 -1819 787 -1791
rect 1374 -1819 1375 -1791
rect 1381 -1922 1382 -1818
rect 1808 -1819 1809 -1791
rect 100 -1922 101 -1820
rect 415 -1821 416 -1791
rect 422 -1821 423 -1791
rect 670 -1922 671 -1820
rect 726 -1922 727 -1820
rect 1027 -1821 1028 -1791
rect 1052 -1922 1053 -1820
rect 1150 -1821 1151 -1791
rect 1374 -1922 1375 -1820
rect 1416 -1821 1417 -1791
rect 1577 -1821 1578 -1791
rect 1738 -1922 1739 -1820
rect 110 -1922 111 -1822
rect 1234 -1922 1235 -1822
rect 1416 -1922 1417 -1822
rect 1584 -1823 1585 -1791
rect 128 -1922 129 -1824
rect 149 -1825 150 -1791
rect 159 -1825 160 -1791
rect 1839 -1825 1840 -1791
rect 149 -1922 150 -1826
rect 520 -1827 521 -1791
rect 527 -1827 528 -1791
rect 534 -1922 535 -1826
rect 730 -1922 731 -1826
rect 758 -1827 759 -1791
rect 765 -1827 766 -1791
rect 887 -1827 888 -1791
rect 891 -1922 892 -1826
rect 954 -1827 955 -1791
rect 975 -1827 976 -1791
rect 1269 -1827 1270 -1791
rect 1293 -1827 1294 -1791
rect 1584 -1922 1585 -1826
rect 170 -1829 171 -1791
rect 1125 -1922 1126 -1828
rect 1150 -1922 1151 -1828
rect 1164 -1922 1165 -1828
rect 1269 -1922 1270 -1828
rect 1458 -1829 1459 -1791
rect 1577 -1922 1578 -1828
rect 1619 -1829 1620 -1791
rect 443 -1922 444 -1830
rect 471 -1831 472 -1791
rect 625 -1922 626 -1830
rect 733 -1831 734 -1791
rect 828 -1831 829 -1791
rect 831 -1922 832 -1830
rect 1780 -1831 1781 -1791
rect 114 -1922 115 -1832
rect 828 -1922 829 -1832
rect 856 -1833 857 -1791
rect 884 -1922 885 -1832
rect 898 -1922 899 -1832
rect 919 -1833 920 -1791
rect 947 -1922 948 -1832
rect 1384 -1922 1385 -1832
rect 1426 -1922 1427 -1832
rect 1535 -1922 1536 -1832
rect 219 -1835 220 -1791
rect 324 -1835 325 -1791
rect 341 -1922 342 -1834
rect 1094 -1835 1095 -1791
rect 1290 -1835 1291 -1791
rect 1619 -1922 1620 -1834
rect 135 -1837 136 -1791
rect 324 -1922 325 -1836
rect 352 -1837 353 -1791
rect 352 -1922 353 -1836
rect 352 -1837 353 -1791
rect 352 -1922 353 -1836
rect 359 -1922 360 -1836
rect 562 -1837 563 -1791
rect 758 -1922 759 -1836
rect 793 -1837 794 -1791
rect 810 -1922 811 -1836
rect 1311 -1837 1312 -1791
rect 1458 -1922 1459 -1836
rect 1465 -1837 1466 -1791
rect 135 -1922 136 -1838
rect 163 -1839 164 -1791
rect 222 -1839 223 -1791
rect 716 -1922 717 -1838
rect 765 -1922 766 -1838
rect 1059 -1839 1060 -1791
rect 1066 -1922 1067 -1838
rect 1157 -1839 1158 -1791
rect 1311 -1922 1312 -1838
rect 1353 -1839 1354 -1791
rect 1465 -1922 1466 -1838
rect 1472 -1839 1473 -1791
rect 163 -1922 164 -1840
rect 191 -1841 192 -1791
rect 222 -1922 223 -1840
rect 1598 -1841 1599 -1791
rect 191 -1922 192 -1842
rect 254 -1843 255 -1791
rect 261 -1843 262 -1791
rect 499 -1922 500 -1842
rect 527 -1922 528 -1842
rect 1206 -1922 1207 -1842
rect 1353 -1922 1354 -1842
rect 1402 -1843 1403 -1791
rect 1430 -1843 1431 -1791
rect 1472 -1922 1473 -1842
rect 1570 -1843 1571 -1791
rect 1598 -1922 1599 -1842
rect 61 -1922 62 -1844
rect 261 -1922 262 -1844
rect 268 -1922 269 -1844
rect 485 -1845 486 -1791
rect 544 -1845 545 -1791
rect 1290 -1922 1291 -1844
rect 1297 -1845 1298 -1791
rect 1430 -1922 1431 -1844
rect 1570 -1922 1571 -1844
rect 1822 -1845 1823 -1791
rect 173 -1922 174 -1846
rect 1402 -1922 1403 -1846
rect 226 -1849 227 -1791
rect 404 -1922 405 -1848
rect 415 -1922 416 -1848
rect 593 -1849 594 -1791
rect 786 -1922 787 -1848
rect 1647 -1849 1648 -1791
rect 23 -1851 24 -1791
rect 593 -1922 594 -1850
rect 793 -1922 794 -1850
rect 842 -1851 843 -1791
rect 856 -1922 857 -1850
rect 1097 -1922 1098 -1850
rect 1157 -1922 1158 -1850
rect 1717 -1851 1718 -1791
rect 226 -1922 227 -1852
rect 632 -1853 633 -1791
rect 814 -1922 815 -1852
rect 870 -1853 871 -1791
rect 901 -1853 902 -1791
rect 1654 -1853 1655 -1791
rect 233 -1855 234 -1791
rect 289 -1855 290 -1791
rect 303 -1855 304 -1791
rect 380 -1855 381 -1791
rect 394 -1922 395 -1854
rect 789 -1855 790 -1791
rect 821 -1922 822 -1854
rect 1136 -1855 1137 -1791
rect 1297 -1922 1298 -1854
rect 1339 -1855 1340 -1791
rect 1605 -1855 1606 -1791
rect 1717 -1922 1718 -1854
rect 44 -1857 45 -1791
rect 789 -1922 790 -1856
rect 824 -1857 825 -1791
rect 1059 -1922 1060 -1856
rect 1080 -1857 1081 -1791
rect 1136 -1922 1137 -1856
rect 1605 -1922 1606 -1856
rect 1766 -1857 1767 -1791
rect 44 -1922 45 -1858
rect 744 -1859 745 -1791
rect 842 -1922 843 -1858
rect 905 -1859 906 -1791
rect 919 -1922 920 -1858
rect 968 -1859 969 -1791
rect 975 -1922 976 -1858
rect 1017 -1859 1018 -1791
rect 1024 -1922 1025 -1858
rect 1409 -1859 1410 -1791
rect 1647 -1922 1648 -1858
rect 1710 -1859 1711 -1791
rect 219 -1922 220 -1860
rect 303 -1922 304 -1860
rect 317 -1922 318 -1860
rect 506 -1861 507 -1791
rect 562 -1922 563 -1860
rect 800 -1861 801 -1791
rect 870 -1922 871 -1860
rect 1087 -1922 1088 -1860
rect 1094 -1922 1095 -1860
rect 1626 -1861 1627 -1791
rect 1654 -1922 1655 -1860
rect 1703 -1861 1704 -1791
rect 1710 -1922 1711 -1860
rect 1773 -1861 1774 -1791
rect 198 -1863 199 -1791
rect 506 -1922 507 -1862
rect 632 -1922 633 -1862
rect 639 -1863 640 -1791
rect 702 -1863 703 -1791
rect 744 -1922 745 -1862
rect 800 -1922 801 -1862
rect 849 -1863 850 -1791
rect 877 -1863 878 -1791
rect 968 -1922 969 -1862
rect 1017 -1922 1018 -1862
rect 1073 -1863 1074 -1791
rect 1080 -1922 1081 -1862
rect 1115 -1863 1116 -1791
rect 1346 -1863 1347 -1791
rect 1766 -1922 1767 -1862
rect 86 -1865 87 -1791
rect 1073 -1922 1074 -1864
rect 1409 -1922 1410 -1864
rect 1437 -1865 1438 -1791
rect 1626 -1922 1627 -1864
rect 1682 -1865 1683 -1791
rect 1703 -1922 1704 -1864
rect 1759 -1865 1760 -1791
rect 86 -1922 87 -1866
rect 408 -1867 409 -1791
rect 422 -1922 423 -1866
rect 450 -1867 451 -1791
rect 471 -1922 472 -1866
rect 985 -1922 986 -1866
rect 1045 -1867 1046 -1791
rect 1115 -1922 1116 -1866
rect 1437 -1922 1438 -1866
rect 1521 -1867 1522 -1791
rect 1591 -1867 1592 -1791
rect 1682 -1922 1683 -1866
rect 156 -1869 157 -1791
rect 1346 -1922 1347 -1868
rect 1521 -1922 1522 -1868
rect 1542 -1869 1543 -1791
rect 1591 -1922 1592 -1868
rect 1612 -1869 1613 -1791
rect 1633 -1869 1634 -1791
rect 1759 -1922 1760 -1868
rect 156 -1922 157 -1870
rect 247 -1871 248 -1791
rect 254 -1922 255 -1870
rect 719 -1871 720 -1791
rect 849 -1922 850 -1870
rect 1304 -1871 1305 -1791
rect 1542 -1922 1543 -1870
rect 1549 -1871 1550 -1791
rect 1612 -1922 1613 -1870
rect 1675 -1871 1676 -1791
rect 198 -1922 199 -1872
rect 345 -1873 346 -1791
rect 366 -1873 367 -1791
rect 835 -1922 836 -1872
rect 877 -1922 878 -1872
rect 1010 -1873 1011 -1791
rect 1045 -1922 1046 -1872
rect 1171 -1873 1172 -1791
rect 1304 -1922 1305 -1872
rect 1318 -1873 1319 -1791
rect 1549 -1922 1550 -1872
rect 1556 -1873 1557 -1791
rect 1633 -1922 1634 -1872
rect 1696 -1873 1697 -1791
rect 240 -1875 241 -1791
rect 289 -1922 290 -1874
rect 296 -1875 297 -1791
rect 408 -1922 409 -1874
rect 429 -1875 430 -1791
rect 709 -1922 710 -1874
rect 905 -1922 906 -1874
rect 1146 -1875 1147 -1791
rect 1171 -1922 1172 -1874
rect 1220 -1875 1221 -1791
rect 1318 -1922 1319 -1874
rect 1367 -1875 1368 -1791
rect 1675 -1922 1676 -1874
rect 1731 -1875 1732 -1791
rect 275 -1877 276 -1791
rect 520 -1922 521 -1876
rect 618 -1877 619 -1791
rect 639 -1922 640 -1876
rect 702 -1922 703 -1876
rect 961 -1877 962 -1791
rect 1010 -1922 1011 -1876
rect 1031 -1877 1032 -1791
rect 1360 -1877 1361 -1791
rect 1556 -1922 1557 -1876
rect 1696 -1922 1697 -1876
rect 1752 -1877 1753 -1791
rect 275 -1922 276 -1878
rect 660 -1879 661 -1791
rect 688 -1879 689 -1791
rect 961 -1922 962 -1878
rect 1360 -1922 1361 -1878
rect 1388 -1879 1389 -1791
rect 1731 -1922 1732 -1878
rect 1801 -1879 1802 -1791
rect 282 -1881 283 -1791
rect 362 -1881 363 -1791
rect 366 -1922 367 -1880
rect 604 -1881 605 -1791
rect 618 -1922 619 -1880
rect 1339 -1922 1340 -1880
rect 1367 -1922 1368 -1880
rect 1479 -1881 1480 -1791
rect 282 -1922 283 -1882
rect 310 -1883 311 -1791
rect 331 -1883 332 -1791
rect 450 -1922 451 -1882
rect 478 -1922 479 -1882
rect 492 -1883 493 -1791
rect 579 -1883 580 -1791
rect 1388 -1922 1389 -1882
rect 1479 -1922 1480 -1882
rect 1500 -1883 1501 -1791
rect 205 -1885 206 -1791
rect 310 -1922 311 -1884
rect 331 -1922 332 -1884
rect 338 -1922 339 -1884
rect 345 -1922 346 -1884
rect 1160 -1922 1161 -1884
rect 1500 -1922 1501 -1884
rect 1507 -1885 1508 -1791
rect 205 -1922 206 -1886
rect 940 -1887 941 -1791
rect 954 -1922 955 -1886
rect 1003 -1887 1004 -1791
rect 1507 -1922 1508 -1886
rect 1514 -1887 1515 -1791
rect 296 -1922 297 -1888
rect 464 -1889 465 -1791
rect 485 -1922 486 -1888
rect 653 -1889 654 -1791
rect 660 -1922 661 -1888
rect 681 -1889 682 -1791
rect 688 -1922 689 -1888
rect 978 -1889 979 -1791
rect 1514 -1922 1515 -1888
rect 1528 -1889 1529 -1791
rect 121 -1891 122 -1791
rect 653 -1922 654 -1890
rect 681 -1922 682 -1890
rect 1038 -1891 1039 -1791
rect 1486 -1891 1487 -1791
rect 1528 -1922 1529 -1890
rect 121 -1922 122 -1892
rect 737 -1893 738 -1791
rect 779 -1893 780 -1791
rect 1220 -1922 1221 -1892
rect 380 -1922 381 -1894
rect 383 -1895 384 -1791
rect 401 -1895 402 -1791
rect 464 -1922 465 -1894
rect 492 -1922 493 -1894
rect 912 -1895 913 -1791
rect 933 -1895 934 -1791
rect 1031 -1922 1032 -1894
rect 1038 -1922 1039 -1894
rect 1108 -1895 1109 -1791
rect 1129 -1895 1130 -1791
rect 1486 -1922 1487 -1894
rect 401 -1922 402 -1896
rect 1724 -1922 1725 -1896
rect 436 -1899 437 -1791
rect 604 -1922 605 -1898
rect 737 -1922 738 -1898
rect 807 -1899 808 -1791
rect 912 -1922 913 -1898
rect 1395 -1922 1396 -1898
rect 51 -1901 52 -1791
rect 807 -1922 808 -1900
rect 933 -1922 934 -1900
rect 982 -1901 983 -1791
rect 1108 -1922 1109 -1900
rect 1276 -1901 1277 -1791
rect 51 -1922 52 -1902
rect 243 -1922 244 -1902
rect 436 -1922 437 -1902
rect 555 -1903 556 -1791
rect 751 -1903 752 -1791
rect 779 -1922 780 -1902
rect 940 -1922 941 -1902
rect 996 -1903 997 -1791
rect 1122 -1903 1123 -1791
rect 1276 -1922 1277 -1902
rect 551 -1905 552 -1791
rect 1003 -1922 1004 -1904
rect 1129 -1922 1130 -1904
rect 1199 -1905 1200 -1791
rect 555 -1922 556 -1906
rect 569 -1907 570 -1791
rect 751 -1922 752 -1906
rect 926 -1907 927 -1791
rect 1199 -1922 1200 -1906
rect 1255 -1907 1256 -1791
rect 513 -1909 514 -1791
rect 569 -1922 570 -1908
rect 926 -1922 927 -1908
rect 989 -1909 990 -1791
rect 1241 -1909 1242 -1791
rect 1255 -1922 1256 -1908
rect 107 -1911 108 -1791
rect 513 -1922 514 -1910
rect 1185 -1911 1186 -1791
rect 1241 -1922 1242 -1910
rect 107 -1922 108 -1912
rect 863 -1913 864 -1791
rect 1185 -1922 1186 -1912
rect 1248 -1913 1249 -1791
rect 233 -1922 234 -1914
rect 989 -1922 990 -1914
rect 1248 -1922 1249 -1914
rect 1262 -1915 1263 -1791
rect 590 -1917 591 -1791
rect 1262 -1922 1263 -1916
rect 590 -1922 591 -1918
rect 996 -1922 997 -1918
rect 863 -1922 864 -1920
rect 1167 -1922 1168 -1920
rect 23 -2049 24 -1931
rect 936 -2049 937 -1931
rect 950 -2049 951 -1931
rect 1136 -1932 1137 -1930
rect 1143 -1932 1144 -1930
rect 1143 -2049 1144 -1931
rect 1143 -1932 1144 -1930
rect 1143 -2049 1144 -1931
rect 1157 -1932 1158 -1930
rect 1766 -1932 1767 -1930
rect 30 -1934 31 -1930
rect 61 -1934 62 -1930
rect 65 -1934 66 -1930
rect 506 -1934 507 -1930
rect 534 -1934 535 -1930
rect 607 -2049 608 -1933
rect 618 -1934 619 -1930
rect 1290 -1934 1291 -1930
rect 1297 -1934 1298 -1930
rect 1297 -2049 1298 -1933
rect 1297 -1934 1298 -1930
rect 1297 -2049 1298 -1933
rect 1304 -1934 1305 -1930
rect 1304 -2049 1305 -1933
rect 1304 -1934 1305 -1930
rect 1304 -2049 1305 -1933
rect 1318 -1934 1319 -1930
rect 1318 -2049 1319 -1933
rect 1318 -1934 1319 -1930
rect 1318 -2049 1319 -1933
rect 1381 -1934 1382 -1930
rect 1675 -1934 1676 -1930
rect 1738 -1934 1739 -1930
rect 1773 -2049 1774 -1933
rect 37 -1936 38 -1930
rect 170 -1936 171 -1930
rect 219 -1936 220 -1930
rect 394 -1936 395 -1930
rect 408 -1936 409 -1930
rect 600 -2049 601 -1935
rect 656 -1936 657 -1930
rect 1717 -1936 1718 -1930
rect 37 -2049 38 -1937
rect 86 -1938 87 -1930
rect 93 -1938 94 -1930
rect 768 -2049 769 -1937
rect 772 -1938 773 -1930
rect 933 -1938 934 -1930
rect 968 -1938 969 -1930
rect 968 -2049 969 -1937
rect 968 -1938 969 -1930
rect 968 -2049 969 -1937
rect 985 -1938 986 -1930
rect 1360 -1938 1361 -1930
rect 1381 -2049 1382 -1937
rect 1395 -1938 1396 -1930
rect 1619 -1938 1620 -1930
rect 1619 -2049 1620 -1937
rect 1619 -1938 1620 -1930
rect 1619 -2049 1620 -1937
rect 1626 -1938 1627 -1930
rect 1626 -2049 1627 -1937
rect 1626 -1938 1627 -1930
rect 1626 -2049 1627 -1937
rect 1633 -1938 1634 -1930
rect 1633 -2049 1634 -1937
rect 1633 -1938 1634 -1930
rect 1633 -2049 1634 -1937
rect 1640 -1938 1641 -1930
rect 1738 -2049 1739 -1937
rect 58 -2049 59 -1939
rect 604 -1940 605 -1930
rect 716 -1940 717 -1930
rect 803 -2049 804 -1939
rect 849 -2049 850 -1939
rect 898 -1940 899 -1930
rect 912 -1940 913 -1930
rect 1591 -1940 1592 -1930
rect 1640 -2049 1641 -1939
rect 1654 -1940 1655 -1930
rect 1675 -2049 1676 -1939
rect 1710 -1940 1711 -1930
rect 1717 -2049 1718 -1939
rect 1745 -1940 1746 -1930
rect 68 -1942 69 -1930
rect 1689 -1942 1690 -1930
rect 1710 -2049 1711 -1941
rect 1724 -1942 1725 -1930
rect 79 -1944 80 -1930
rect 93 -2049 94 -1943
rect 100 -1944 101 -1930
rect 534 -2049 535 -1943
rect 583 -1944 584 -1930
rect 583 -2049 584 -1943
rect 583 -1944 584 -1930
rect 583 -2049 584 -1943
rect 604 -2049 605 -1943
rect 681 -1944 682 -1930
rect 716 -2049 717 -1943
rect 730 -1944 731 -1930
rect 744 -1944 745 -1930
rect 744 -2049 745 -1943
rect 744 -1944 745 -1930
rect 744 -2049 745 -1943
rect 754 -2049 755 -1943
rect 821 -1944 822 -1930
rect 873 -1944 874 -1930
rect 1108 -1944 1109 -1930
rect 1122 -1944 1123 -1930
rect 1493 -1944 1494 -1930
rect 1500 -1944 1501 -1930
rect 1689 -2049 1690 -1943
rect 79 -2049 80 -1945
rect 135 -1946 136 -1930
rect 138 -2049 139 -1945
rect 639 -1946 640 -1930
rect 646 -1946 647 -1930
rect 681 -2049 682 -1945
rect 723 -2049 724 -1945
rect 933 -2049 934 -1945
rect 989 -1946 990 -1930
rect 1367 -1946 1368 -1930
rect 1384 -1946 1385 -1930
rect 1528 -1946 1529 -1930
rect 1549 -1946 1550 -1930
rect 1591 -2049 1592 -1945
rect 1654 -2049 1655 -1945
rect 1661 -1946 1662 -1930
rect 1682 -1946 1683 -1930
rect 1745 -2049 1746 -1945
rect 100 -2049 101 -1947
rect 142 -1948 143 -1930
rect 149 -1948 150 -1930
rect 908 -2049 909 -1947
rect 912 -2049 913 -1947
rect 954 -1948 955 -1930
rect 1059 -1948 1060 -1930
rect 1766 -2049 1767 -1947
rect 107 -1950 108 -1930
rect 317 -1950 318 -1930
rect 359 -1950 360 -1930
rect 870 -1950 871 -1930
rect 884 -1950 885 -1930
rect 884 -2049 885 -1949
rect 884 -1950 885 -1930
rect 884 -2049 885 -1949
rect 898 -2049 899 -1949
rect 940 -1950 941 -1930
rect 947 -1950 948 -1930
rect 989 -2049 990 -1949
rect 1080 -1950 1081 -1930
rect 1108 -2049 1109 -1949
rect 1157 -2049 1158 -1949
rect 1171 -1950 1172 -1930
rect 1185 -1950 1186 -1930
rect 1188 -1990 1189 -1949
rect 1199 -1950 1200 -1930
rect 1199 -2049 1200 -1949
rect 1199 -1950 1200 -1930
rect 1199 -2049 1200 -1949
rect 1227 -1950 1228 -1930
rect 1416 -1950 1417 -1930
rect 1423 -1950 1424 -1930
rect 1500 -2049 1501 -1949
rect 1528 -2049 1529 -1949
rect 1762 -2049 1763 -1949
rect 135 -2049 136 -1951
rect 1220 -1952 1221 -1930
rect 1234 -1952 1235 -1930
rect 1234 -2049 1235 -1951
rect 1234 -1952 1235 -1930
rect 1234 -2049 1235 -1951
rect 1269 -1952 1270 -1930
rect 1269 -2049 1270 -1951
rect 1269 -1952 1270 -1930
rect 1269 -2049 1270 -1951
rect 1290 -2049 1291 -1951
rect 1472 -1952 1473 -1930
rect 1570 -1952 1571 -1930
rect 1724 -2049 1725 -1951
rect 142 -2049 143 -1953
rect 541 -1954 542 -1930
rect 597 -1954 598 -1930
rect 954 -2049 955 -1953
rect 1066 -1954 1067 -1930
rect 1080 -2049 1081 -1953
rect 1087 -1954 1088 -1930
rect 1122 -2049 1123 -1953
rect 1160 -1954 1161 -1930
rect 1759 -1954 1760 -1930
rect 149 -2049 150 -1955
rect 163 -1956 164 -1930
rect 166 -2049 167 -1955
rect 709 -1956 710 -1930
rect 730 -2049 731 -1955
rect 1020 -2049 1021 -1955
rect 1097 -1956 1098 -1930
rect 1437 -1956 1438 -1930
rect 1661 -2049 1662 -1955
rect 1668 -1956 1669 -1930
rect 1682 -2049 1683 -1955
rect 1752 -2049 1753 -1955
rect 1759 -2049 1760 -1955
rect 1794 -1956 1795 -1930
rect 65 -2049 66 -1957
rect 163 -2049 164 -1957
rect 170 -2049 171 -1957
rect 415 -1958 416 -1930
rect 432 -1958 433 -1930
rect 1136 -2049 1137 -1957
rect 1167 -1958 1168 -1930
rect 1647 -1958 1648 -1930
rect 1668 -2049 1669 -1957
rect 1703 -1958 1704 -1930
rect 159 -2049 160 -1959
rect 352 -1960 353 -1930
rect 359 -2049 360 -1959
rect 527 -1960 528 -1930
rect 639 -2049 640 -1959
rect 919 -1960 920 -1930
rect 929 -2049 930 -1959
rect 1570 -2049 1571 -1959
rect 1696 -1960 1697 -1930
rect 1703 -2049 1704 -1959
rect 72 -1962 73 -1930
rect 352 -2049 353 -1961
rect 380 -1962 381 -1930
rect 621 -1962 622 -1930
rect 646 -2049 647 -1961
rect 660 -1962 661 -1930
rect 670 -1962 671 -1930
rect 1696 -2049 1697 -1961
rect 72 -2049 73 -1963
rect 131 -2049 132 -1963
rect 219 -2049 220 -1963
rect 373 -1964 374 -1930
rect 394 -2049 395 -1963
rect 436 -1964 437 -1930
rect 471 -1964 472 -1930
rect 541 -2049 542 -1963
rect 621 -2049 622 -1963
rect 1535 -1964 1536 -1930
rect 51 -1966 52 -1930
rect 471 -2049 472 -1965
rect 492 -1966 493 -1930
rect 593 -1966 594 -1930
rect 660 -2049 661 -1965
rect 1150 -1966 1151 -1930
rect 1171 -2049 1172 -1965
rect 1178 -1966 1179 -1930
rect 1185 -2049 1186 -1965
rect 1241 -1966 1242 -1930
rect 1325 -1966 1326 -1930
rect 1472 -2049 1473 -1965
rect 51 -2049 52 -1967
rect 345 -1968 346 -1930
rect 373 -2049 374 -1967
rect 817 -2049 818 -1967
rect 821 -2049 822 -1967
rect 856 -1968 857 -1930
rect 877 -1968 878 -1930
rect 1150 -2049 1151 -1967
rect 1178 -2049 1179 -1967
rect 1563 -1968 1564 -1930
rect 117 -2049 118 -1969
rect 436 -2049 437 -1969
rect 450 -1970 451 -1930
rect 492 -2049 493 -1969
rect 506 -2049 507 -1969
rect 569 -1970 570 -1930
rect 593 -2049 594 -1969
rect 1395 -2049 1396 -1969
rect 1444 -1970 1445 -1930
rect 1647 -2049 1648 -1969
rect 226 -1972 227 -1930
rect 310 -1972 311 -1930
rect 324 -1972 325 -1930
rect 380 -2049 381 -1971
rect 401 -1972 402 -1930
rect 1066 -2049 1067 -1971
rect 1101 -1972 1102 -1930
rect 1416 -2049 1417 -1971
rect 1444 -2049 1445 -1971
rect 1465 -1972 1466 -1930
rect 1514 -1972 1515 -1930
rect 1563 -2049 1564 -1971
rect 177 -1974 178 -1930
rect 226 -2049 227 -1973
rect 240 -1974 241 -1930
rect 338 -1974 339 -1930
rect 345 -2049 346 -1973
rect 513 -1974 514 -1930
rect 555 -1974 556 -1930
rect 569 -2049 570 -1973
rect 670 -2049 671 -1973
rect 905 -1974 906 -1930
rect 915 -1974 916 -1930
rect 1248 -1974 1249 -1930
rect 1353 -1974 1354 -1930
rect 1549 -2049 1550 -1973
rect 156 -1976 157 -1930
rect 513 -2049 514 -1975
rect 691 -2049 692 -1975
rect 1514 -2049 1515 -1975
rect 156 -2049 157 -1977
rect 726 -1978 727 -1930
rect 765 -1978 766 -1930
rect 1493 -2049 1494 -1977
rect 177 -2049 178 -1979
rect 985 -2049 986 -1979
rect 1024 -1980 1025 -1930
rect 1353 -2049 1354 -1979
rect 1360 -2049 1361 -1979
rect 1374 -1980 1375 -1930
rect 1388 -1980 1389 -1930
rect 1423 -2049 1424 -1979
rect 184 -1982 185 -1930
rect 338 -2049 339 -1981
rect 401 -2049 402 -1981
rect 684 -1982 685 -1930
rect 695 -1982 696 -1930
rect 709 -2049 710 -1981
rect 765 -2049 766 -1981
rect 1059 -2049 1060 -1981
rect 1073 -1982 1074 -1930
rect 1101 -2049 1102 -1981
rect 1115 -1982 1116 -1930
rect 1220 -2049 1221 -1981
rect 1230 -1982 1231 -1930
rect 1248 -2049 1249 -1981
rect 1367 -2049 1368 -1981
rect 1451 -1982 1452 -1930
rect 184 -2049 185 -1983
rect 835 -1984 836 -1930
rect 856 -2049 857 -1983
rect 1206 -1984 1207 -1930
rect 1213 -1984 1214 -1930
rect 1227 -2049 1228 -1983
rect 1374 -2049 1375 -1983
rect 1479 -1984 1480 -1930
rect 205 -1986 206 -1930
rect 835 -2049 836 -1985
rect 905 -2049 906 -1985
rect 1612 -1986 1613 -1930
rect 205 -2049 206 -1987
rect 208 -2049 209 -1987
rect 233 -1988 234 -1930
rect 695 -2049 696 -1987
rect 702 -1988 703 -1930
rect 870 -2049 871 -1987
rect 940 -2049 941 -1987
rect 975 -1988 976 -1930
rect 1038 -1988 1039 -1930
rect 1073 -2049 1074 -1987
rect 1087 -2049 1088 -1987
rect 1115 -2049 1116 -1987
rect 1192 -1988 1193 -1930
rect 1241 -2049 1242 -1987
rect 1388 -2049 1389 -1987
rect 1402 -1988 1403 -1930
rect 1409 -1988 1410 -1930
rect 1465 -2049 1466 -1987
rect 1584 -1988 1585 -1930
rect 1612 -2049 1613 -1987
rect 233 -2049 234 -1989
rect 597 -2049 598 -1989
rect 702 -2049 703 -1989
rect 996 -1990 997 -1930
rect 1017 -1990 1018 -1930
rect 1038 -2049 1039 -1989
rect 1192 -2049 1193 -1989
rect 1213 -2049 1214 -1989
rect 1339 -1990 1340 -1930
rect 1402 -2049 1403 -1989
rect 1542 -1990 1543 -1930
rect 240 -2049 241 -1991
rect 387 -1992 388 -1930
rect 408 -2049 409 -1991
rect 653 -1992 654 -1930
rect 688 -1992 689 -1930
rect 996 -2049 997 -1991
rect 1017 -2049 1018 -1991
rect 1283 -1992 1284 -1930
rect 1409 -2049 1410 -1991
rect 1458 -1992 1459 -1930
rect 1542 -2049 1543 -1991
rect 1605 -1992 1606 -1930
rect 247 -1994 248 -1930
rect 310 -2049 311 -1993
rect 324 -2049 325 -1993
rect 674 -1994 675 -1930
rect 772 -2049 773 -1993
rect 842 -1994 843 -1930
rect 975 -2049 976 -1993
rect 1003 -1994 1004 -1930
rect 1129 -1994 1130 -1930
rect 1339 -2049 1340 -1993
rect 1430 -1994 1431 -1930
rect 1479 -2049 1480 -1993
rect 1598 -1994 1599 -1930
rect 1605 -2049 1606 -1993
rect 107 -2049 108 -1995
rect 674 -2049 675 -1995
rect 789 -1996 790 -1930
rect 1024 -2049 1025 -1995
rect 1052 -1996 1053 -1930
rect 1129 -2049 1130 -1995
rect 1276 -1996 1277 -1930
rect 1283 -2049 1284 -1995
rect 1332 -1996 1333 -1930
rect 1430 -2049 1431 -1995
rect 1556 -1996 1557 -1930
rect 1598 -2049 1599 -1995
rect 243 -1998 244 -1930
rect 247 -2049 248 -1997
rect 250 -1998 251 -1930
rect 1255 -1998 1256 -1930
rect 1332 -2049 1333 -1997
rect 1346 -1998 1347 -1930
rect 1556 -2049 1557 -1997
rect 1577 -1998 1578 -1930
rect 254 -2000 255 -1930
rect 415 -2049 416 -1999
rect 450 -2049 451 -1999
rect 635 -2049 636 -1999
rect 667 -2000 668 -1930
rect 1052 -2049 1053 -1999
rect 1255 -2049 1256 -1999
rect 1437 -2049 1438 -1999
rect 1577 -2049 1578 -1999
rect 1731 -2000 1732 -1930
rect 254 -2049 255 -2001
rect 289 -2002 290 -1930
rect 303 -2002 304 -1930
rect 317 -2049 318 -2001
rect 387 -2049 388 -2001
rect 548 -2002 549 -1930
rect 576 -2002 577 -1930
rect 653 -2049 654 -2001
rect 667 -2049 668 -2001
rect 1325 -2049 1326 -2001
rect 1346 -2049 1347 -2001
rect 1507 -2002 1508 -1930
rect 1521 -2002 1522 -1930
rect 1731 -2049 1732 -2001
rect 268 -2004 269 -1930
rect 618 -2049 619 -2003
rect 800 -2004 801 -1930
rect 982 -2004 983 -1930
rect 1003 -2049 1004 -2003
rect 1010 -2004 1011 -1930
rect 1262 -2004 1263 -1930
rect 1507 -2049 1508 -2003
rect 198 -2006 199 -1930
rect 268 -2049 269 -2005
rect 275 -2006 276 -1930
rect 530 -2006 531 -1930
rect 548 -2049 549 -2005
rect 688 -2049 689 -2005
rect 800 -2049 801 -2005
rect 877 -2049 878 -2005
rect 1010 -2049 1011 -2005
rect 1164 -2006 1165 -1930
rect 1311 -2006 1312 -1930
rect 1521 -2049 1522 -2005
rect 110 -2049 111 -2007
rect 275 -2049 276 -2007
rect 282 -2008 283 -1930
rect 369 -2049 370 -2007
rect 457 -2008 458 -1930
rect 576 -2049 577 -2007
rect 590 -2008 591 -1930
rect 1584 -2049 1585 -2007
rect 114 -2010 115 -1930
rect 198 -2049 199 -2009
rect 229 -2010 230 -1930
rect 1311 -2049 1312 -2009
rect 114 -2049 115 -2011
rect 1276 -2049 1277 -2011
rect 282 -2049 283 -2013
rect 782 -2049 783 -2013
rect 807 -2014 808 -1930
rect 919 -2049 920 -2013
rect 1045 -2014 1046 -1930
rect 1262 -2049 1263 -2013
rect 289 -2049 290 -2015
rect 429 -2016 430 -1930
rect 457 -2049 458 -2015
rect 625 -2016 626 -1930
rect 793 -2016 794 -1930
rect 807 -2049 808 -2015
rect 810 -2016 811 -1930
rect 1535 -2049 1536 -2015
rect 303 -2049 304 -2017
rect 331 -2018 332 -1930
rect 404 -2018 405 -1930
rect 1045 -2049 1046 -2017
rect 1164 -2049 1165 -2017
rect 1258 -2049 1259 -2017
rect 331 -2049 332 -2019
rect 366 -2020 367 -1930
rect 429 -2049 430 -2019
rect 611 -2020 612 -1930
rect 625 -2049 626 -2019
rect 863 -2020 864 -1930
rect 485 -2022 486 -1930
rect 611 -2049 612 -2021
rect 814 -2022 815 -1930
rect 842 -2049 843 -2021
rect 863 -2049 864 -2021
rect 891 -2022 892 -1930
rect 443 -2024 444 -1930
rect 485 -2049 486 -2023
rect 499 -2024 500 -1930
rect 1206 -2049 1207 -2023
rect 422 -2026 423 -1930
rect 443 -2049 444 -2025
rect 478 -2026 479 -1930
rect 499 -2049 500 -2025
rect 530 -2049 531 -2025
rect 555 -2049 556 -2025
rect 562 -2026 563 -1930
rect 793 -2049 794 -2025
rect 814 -2049 815 -2025
rect 1486 -2026 1487 -1930
rect 44 -2028 45 -1930
rect 422 -2049 423 -2027
rect 562 -2049 563 -2027
rect 961 -2028 962 -1930
rect 1125 -2028 1126 -1930
rect 1486 -2049 1487 -2027
rect 44 -2049 45 -2029
rect 128 -2030 129 -1930
rect 212 -2030 213 -1930
rect 478 -2049 479 -2029
rect 590 -2049 591 -2029
rect 758 -2030 759 -1930
rect 891 -2049 892 -2029
rect 926 -2030 927 -1930
rect 961 -2049 962 -2029
rect 1031 -2030 1032 -1930
rect 128 -2049 129 -2031
rect 191 -2032 192 -1930
rect 212 -2049 213 -2031
rect 261 -2032 262 -1930
rect 737 -2032 738 -1930
rect 926 -2049 927 -2031
rect 121 -2034 122 -1930
rect 737 -2049 738 -2033
rect 758 -2049 759 -2033
rect 779 -2034 780 -1930
rect 828 -2034 829 -1930
rect 1031 -2049 1032 -2033
rect 121 -2049 122 -2035
rect 1094 -2036 1095 -1930
rect 173 -2038 174 -1930
rect 1094 -2049 1095 -2037
rect 191 -2049 192 -2039
rect 296 -2040 297 -1930
rect 786 -2040 787 -1930
rect 828 -2049 829 -2039
rect 261 -2049 262 -2041
rect 520 -2042 521 -1930
rect 751 -2042 752 -1930
rect 786 -2049 787 -2041
rect 296 -2049 297 -2043
rect 464 -2044 465 -1930
rect 520 -2049 521 -2043
rect 663 -2049 664 -2043
rect 751 -2049 752 -2043
rect 1458 -2049 1459 -2043
rect 464 -2049 465 -2045
rect 632 -2046 633 -1930
rect 86 -2049 87 -2047
rect 632 -2049 633 -2047
rect 40 -2188 41 -2058
rect 1549 -2059 1550 -2057
rect 1626 -2059 1627 -2057
rect 1629 -2059 1630 -2057
rect 1661 -2059 1662 -2057
rect 1661 -2188 1662 -2058
rect 1661 -2059 1662 -2057
rect 1661 -2188 1662 -2058
rect 1675 -2059 1676 -2057
rect 1675 -2188 1676 -2058
rect 1675 -2059 1676 -2057
rect 1675 -2188 1676 -2058
rect 1738 -2059 1739 -2057
rect 1738 -2188 1739 -2058
rect 1738 -2059 1739 -2057
rect 1738 -2188 1739 -2058
rect 1759 -2188 1760 -2058
rect 1766 -2059 1767 -2057
rect 44 -2061 45 -2057
rect 152 -2188 153 -2060
rect 163 -2061 164 -2057
rect 562 -2061 563 -2057
rect 611 -2061 612 -2057
rect 611 -2188 612 -2060
rect 611 -2061 612 -2057
rect 611 -2188 612 -2060
rect 632 -2061 633 -2057
rect 1521 -2061 1522 -2057
rect 1626 -2188 1627 -2060
rect 1654 -2061 1655 -2057
rect 1766 -2188 1767 -2060
rect 1773 -2061 1774 -2057
rect 23 -2063 24 -2057
rect 562 -2188 563 -2062
rect 663 -2063 664 -2057
rect 716 -2063 717 -2057
rect 726 -2188 727 -2062
rect 1017 -2063 1018 -2057
rect 1066 -2063 1067 -2057
rect 1066 -2188 1067 -2062
rect 1066 -2063 1067 -2057
rect 1066 -2188 1067 -2062
rect 1080 -2063 1081 -2057
rect 1080 -2188 1081 -2062
rect 1080 -2063 1081 -2057
rect 1080 -2188 1081 -2062
rect 1090 -2063 1091 -2057
rect 1290 -2063 1291 -2057
rect 1346 -2063 1347 -2057
rect 1521 -2188 1522 -2062
rect 47 -2188 48 -2064
rect 681 -2065 682 -2057
rect 688 -2065 689 -2057
rect 737 -2065 738 -2057
rect 782 -2065 783 -2057
rect 1178 -2065 1179 -2057
rect 1206 -2065 1207 -2057
rect 1752 -2065 1753 -2057
rect 68 -2188 69 -2066
rect 135 -2188 136 -2066
rect 142 -2067 143 -2057
rect 800 -2067 801 -2057
rect 803 -2067 804 -2057
rect 1563 -2067 1564 -2057
rect 100 -2069 101 -2057
rect 779 -2069 780 -2057
rect 786 -2069 787 -2057
rect 800 -2188 801 -2068
rect 835 -2069 836 -2057
rect 835 -2188 836 -2068
rect 835 -2069 836 -2057
rect 835 -2188 836 -2068
rect 873 -2188 874 -2068
rect 1762 -2069 1763 -2057
rect 100 -2188 101 -2070
rect 856 -2071 857 -2057
rect 919 -2071 920 -2057
rect 922 -2083 923 -2070
rect 926 -2071 927 -2057
rect 1416 -2071 1417 -2057
rect 1451 -2071 1452 -2057
rect 1598 -2071 1599 -2057
rect 107 -2073 108 -2057
rect 705 -2188 706 -2072
rect 716 -2188 717 -2072
rect 744 -2073 745 -2057
rect 758 -2073 759 -2057
rect 786 -2188 787 -2072
rect 856 -2188 857 -2072
rect 877 -2073 878 -2057
rect 912 -2073 913 -2057
rect 926 -2188 927 -2072
rect 936 -2073 937 -2057
rect 1703 -2073 1704 -2057
rect 107 -2188 108 -2074
rect 369 -2075 370 -2057
rect 436 -2075 437 -2057
rect 761 -2188 762 -2074
rect 779 -2188 780 -2074
rect 870 -2075 871 -2057
rect 877 -2188 878 -2074
rect 954 -2075 955 -2057
rect 985 -2075 986 -2057
rect 1549 -2188 1550 -2074
rect 1703 -2188 1704 -2074
rect 1710 -2075 1711 -2057
rect 114 -2077 115 -2057
rect 296 -2077 297 -2057
rect 352 -2077 353 -2057
rect 436 -2188 437 -2076
rect 453 -2188 454 -2076
rect 499 -2077 500 -2057
rect 506 -2077 507 -2057
rect 681 -2188 682 -2076
rect 744 -2188 745 -2076
rect 1591 -2077 1592 -2057
rect 1696 -2077 1697 -2057
rect 1710 -2188 1711 -2076
rect 54 -2188 55 -2078
rect 114 -2188 115 -2078
rect 128 -2079 129 -2057
rect 1465 -2079 1466 -2057
rect 1570 -2079 1571 -2057
rect 1591 -2188 1592 -2078
rect 1682 -2079 1683 -2057
rect 1696 -2188 1697 -2078
rect 128 -2188 129 -2080
rect 275 -2081 276 -2057
rect 289 -2081 290 -2057
rect 352 -2188 353 -2080
rect 359 -2081 360 -2057
rect 621 -2081 622 -2057
rect 667 -2081 668 -2057
rect 807 -2081 808 -2057
rect 898 -2081 899 -2057
rect 912 -2188 913 -2080
rect 919 -2188 920 -2080
rect 947 -2081 948 -2057
rect 1339 -2081 1340 -2057
rect 1395 -2081 1396 -2057
rect 1416 -2188 1417 -2080
rect 1451 -2188 1452 -2080
rect 1556 -2081 1557 -2057
rect 1605 -2081 1606 -2057
rect 1682 -2188 1683 -2080
rect 121 -2083 122 -2057
rect 667 -2188 668 -2082
rect 674 -2083 675 -2057
rect 754 -2083 755 -2057
rect 758 -2188 759 -2082
rect 1262 -2083 1263 -2057
rect 1269 -2083 1270 -2057
rect 1465 -2188 1466 -2082
rect 1528 -2083 1529 -2057
rect 1556 -2188 1557 -2082
rect 1605 -2188 1606 -2082
rect 1612 -2083 1613 -2057
rect 1629 -2188 1630 -2082
rect 1654 -2188 1655 -2082
rect 121 -2188 122 -2084
rect 149 -2085 150 -2057
rect 163 -2188 164 -2084
rect 821 -2085 822 -2057
rect 884 -2085 885 -2057
rect 947 -2188 948 -2084
rect 989 -2085 990 -2057
rect 1020 -2085 1021 -2057
rect 1104 -2188 1105 -2084
rect 1689 -2085 1690 -2057
rect 173 -2188 174 -2086
rect 1423 -2087 1424 -2057
rect 1500 -2087 1501 -2057
rect 1528 -2188 1529 -2086
rect 1535 -2087 1536 -2057
rect 1570 -2188 1571 -2086
rect 1612 -2188 1613 -2086
rect 1633 -2087 1634 -2057
rect 177 -2089 178 -2057
rect 817 -2089 818 -2057
rect 821 -2188 822 -2088
rect 842 -2089 843 -2057
rect 936 -2188 937 -2088
rect 1262 -2188 1263 -2088
rect 1311 -2089 1312 -2057
rect 1346 -2188 1347 -2088
rect 1353 -2089 1354 -2057
rect 1395 -2188 1396 -2088
rect 1402 -2089 1403 -2057
rect 1563 -2188 1564 -2088
rect 1619 -2089 1620 -2057
rect 1633 -2188 1634 -2088
rect 177 -2188 178 -2090
rect 324 -2091 325 -2057
rect 331 -2091 332 -2057
rect 506 -2188 507 -2090
rect 534 -2091 535 -2057
rect 747 -2188 748 -2090
rect 989 -2188 990 -2090
rect 1038 -2091 1039 -2057
rect 1157 -2091 1158 -2057
rect 1178 -2188 1179 -2090
rect 1199 -2091 1200 -2057
rect 1206 -2188 1207 -2090
rect 1227 -2091 1228 -2057
rect 1290 -2188 1291 -2090
rect 1325 -2091 1326 -2057
rect 1353 -2188 1354 -2090
rect 1402 -2188 1403 -2090
rect 1444 -2091 1445 -2057
rect 1584 -2091 1585 -2057
rect 1619 -2188 1620 -2090
rect 51 -2093 52 -2057
rect 534 -2188 535 -2092
rect 555 -2093 556 -2057
rect 954 -2188 955 -2092
rect 1010 -2093 1011 -2057
rect 1038 -2188 1039 -2092
rect 1073 -2093 1074 -2057
rect 1227 -2188 1228 -2092
rect 1255 -2093 1256 -2057
rect 1598 -2188 1599 -2092
rect 184 -2095 185 -2057
rect 737 -2188 738 -2094
rect 950 -2095 951 -2057
rect 1199 -2188 1200 -2094
rect 1258 -2095 1259 -2057
rect 1731 -2095 1732 -2057
rect 184 -2188 185 -2096
rect 373 -2097 374 -2057
rect 408 -2097 409 -2057
rect 842 -2188 843 -2096
rect 1017 -2188 1018 -2096
rect 1031 -2097 1032 -2057
rect 1073 -2188 1074 -2096
rect 1220 -2097 1221 -2057
rect 1339 -2188 1340 -2096
rect 1367 -2097 1368 -2057
rect 1423 -2188 1424 -2096
rect 1647 -2097 1648 -2057
rect 1717 -2097 1718 -2057
rect 1731 -2188 1732 -2096
rect 191 -2099 192 -2057
rect 635 -2099 636 -2057
rect 674 -2188 675 -2098
rect 723 -2099 724 -2057
rect 817 -2188 818 -2098
rect 1717 -2188 1718 -2098
rect 142 -2188 143 -2100
rect 723 -2188 724 -2100
rect 1031 -2188 1032 -2100
rect 1045 -2101 1046 -2057
rect 1118 -2188 1119 -2100
rect 1325 -2188 1326 -2100
rect 1444 -2188 1445 -2100
rect 1748 -2101 1749 -2057
rect 191 -2188 192 -2102
rect 261 -2103 262 -2057
rect 289 -2188 290 -2102
rect 814 -2103 815 -2057
rect 1045 -2188 1046 -2102
rect 1052 -2103 1053 -2057
rect 1129 -2103 1130 -2057
rect 1367 -2188 1368 -2102
rect 1542 -2103 1543 -2057
rect 1647 -2188 1648 -2102
rect 205 -2105 206 -2057
rect 1514 -2105 1515 -2057
rect 1584 -2188 1585 -2104
rect 1668 -2105 1669 -2057
rect 96 -2188 97 -2106
rect 1668 -2188 1669 -2106
rect 205 -2188 206 -2108
rect 268 -2109 269 -2057
rect 296 -2188 297 -2108
rect 303 -2109 304 -2057
rect 310 -2109 311 -2057
rect 331 -2188 332 -2108
rect 345 -2109 346 -2057
rect 359 -2188 360 -2108
rect 366 -2109 367 -2057
rect 1255 -2188 1256 -2108
rect 1374 -2109 1375 -2057
rect 1514 -2188 1515 -2108
rect 208 -2111 209 -2057
rect 632 -2188 633 -2110
rect 691 -2111 692 -2057
rect 898 -2188 899 -2110
rect 1052 -2188 1053 -2110
rect 1108 -2111 1109 -2057
rect 1115 -2111 1116 -2057
rect 1129 -2188 1130 -2110
rect 1157 -2188 1158 -2110
rect 1213 -2111 1214 -2057
rect 1220 -2188 1221 -2110
rect 1234 -2111 1235 -2057
rect 1332 -2111 1333 -2057
rect 1374 -2188 1375 -2110
rect 1507 -2111 1508 -2057
rect 1542 -2188 1543 -2110
rect 212 -2113 213 -2057
rect 303 -2188 304 -2112
rect 310 -2188 311 -2112
rect 317 -2113 318 -2057
rect 324 -2188 325 -2112
rect 1013 -2188 1014 -2112
rect 1101 -2113 1102 -2057
rect 1108 -2188 1109 -2112
rect 1115 -2188 1116 -2112
rect 1500 -2188 1501 -2112
rect 79 -2115 80 -2057
rect 317 -2188 318 -2114
rect 338 -2115 339 -2057
rect 366 -2188 367 -2114
rect 373 -2188 374 -2114
rect 394 -2115 395 -2057
rect 408 -2188 409 -2114
rect 548 -2115 549 -2057
rect 555 -2188 556 -2114
rect 569 -2115 570 -2057
rect 576 -2115 577 -2057
rect 688 -2188 689 -2114
rect 1171 -2115 1172 -2057
rect 1311 -2188 1312 -2114
rect 1472 -2115 1473 -2057
rect 1507 -2188 1508 -2114
rect 79 -2188 80 -2116
rect 1745 -2117 1746 -2057
rect 156 -2119 157 -2057
rect 394 -2188 395 -2118
rect 422 -2119 423 -2057
rect 807 -2188 808 -2118
rect 1192 -2119 1193 -2057
rect 1213 -2188 1214 -2118
rect 1234 -2188 1235 -2118
rect 1248 -2119 1249 -2057
rect 1437 -2119 1438 -2057
rect 1472 -2188 1473 -2118
rect 1724 -2119 1725 -2057
rect 1745 -2188 1746 -2118
rect 131 -2188 132 -2120
rect 156 -2188 157 -2120
rect 166 -2121 167 -2057
rect 576 -2188 577 -2120
rect 593 -2121 594 -2057
rect 1332 -2188 1333 -2120
rect 1409 -2121 1410 -2057
rect 1437 -2188 1438 -2120
rect 1577 -2121 1578 -2057
rect 1724 -2188 1725 -2120
rect 212 -2188 213 -2122
rect 831 -2188 832 -2122
rect 905 -2123 906 -2057
rect 1577 -2188 1578 -2122
rect 233 -2125 234 -2057
rect 527 -2188 528 -2124
rect 541 -2125 542 -2057
rect 548 -2188 549 -2124
rect 569 -2188 570 -2124
rect 772 -2125 773 -2057
rect 1192 -2188 1193 -2124
rect 1276 -2125 1277 -2057
rect 1388 -2125 1389 -2057
rect 1409 -2188 1410 -2124
rect 233 -2188 234 -2126
rect 254 -2127 255 -2057
rect 338 -2188 339 -2126
rect 415 -2127 416 -2057
rect 429 -2127 430 -2057
rect 499 -2188 500 -2126
rect 530 -2127 531 -2057
rect 541 -2188 542 -2126
rect 607 -2127 608 -2057
rect 1535 -2188 1536 -2126
rect 86 -2129 87 -2057
rect 254 -2188 255 -2128
rect 345 -2188 346 -2128
rect 733 -2188 734 -2128
rect 765 -2129 766 -2057
rect 1171 -2188 1172 -2128
rect 1276 -2188 1277 -2128
rect 1640 -2129 1641 -2057
rect 37 -2131 38 -2057
rect 765 -2188 766 -2130
rect 772 -2188 773 -2130
rect 1493 -2131 1494 -2057
rect 86 -2188 87 -2132
rect 478 -2133 479 -2057
rect 485 -2133 486 -2057
rect 597 -2188 598 -2132
rect 618 -2133 619 -2057
rect 905 -2188 906 -2132
rect 1381 -2133 1382 -2057
rect 1388 -2188 1389 -2132
rect 1479 -2133 1480 -2057
rect 1493 -2188 1494 -2132
rect 30 -2188 31 -2134
rect 618 -2188 619 -2134
rect 621 -2188 622 -2134
rect 646 -2135 647 -2057
rect 660 -2135 661 -2057
rect 1248 -2188 1249 -2134
rect 1360 -2135 1361 -2057
rect 1381 -2188 1382 -2134
rect 1458 -2135 1459 -2057
rect 1479 -2188 1480 -2134
rect 1486 -2135 1487 -2057
rect 1640 -2188 1641 -2134
rect 51 -2188 52 -2136
rect 478 -2188 479 -2136
rect 485 -2188 486 -2136
rect 730 -2137 731 -2057
rect 1059 -2137 1060 -2057
rect 1486 -2188 1487 -2136
rect 240 -2139 241 -2057
rect 275 -2188 276 -2138
rect 387 -2139 388 -2057
rect 422 -2188 423 -2138
rect 429 -2188 430 -2138
rect 968 -2139 969 -2057
rect 1059 -2188 1060 -2138
rect 1087 -2139 1088 -2057
rect 1318 -2139 1319 -2057
rect 1360 -2188 1361 -2138
rect 170 -2141 171 -2057
rect 240 -2188 241 -2140
rect 247 -2141 248 -2057
rect 261 -2188 262 -2140
rect 387 -2188 388 -2140
rect 443 -2141 444 -2057
rect 457 -2141 458 -2057
rect 884 -2188 885 -2140
rect 968 -2188 969 -2140
rect 1003 -2141 1004 -2057
rect 1087 -2188 1088 -2140
rect 1094 -2141 1095 -2057
rect 1304 -2141 1305 -2057
rect 1318 -2188 1319 -2140
rect 93 -2143 94 -2057
rect 457 -2188 458 -2142
rect 464 -2143 465 -2057
rect 590 -2188 591 -2142
rect 653 -2143 654 -2057
rect 730 -2188 731 -2142
rect 814 -2188 815 -2142
rect 1003 -2188 1004 -2142
rect 1094 -2188 1095 -2142
rect 1143 -2143 1144 -2057
rect 1297 -2143 1298 -2057
rect 1304 -2188 1305 -2142
rect 93 -2188 94 -2144
rect 996 -2145 997 -2057
rect 1122 -2145 1123 -2057
rect 1143 -2188 1144 -2144
rect 1283 -2145 1284 -2057
rect 1297 -2188 1298 -2144
rect 58 -2147 59 -2057
rect 996 -2188 997 -2146
rect 1241 -2147 1242 -2057
rect 1283 -2188 1284 -2146
rect 58 -2188 59 -2148
rect 625 -2149 626 -2057
rect 670 -2149 671 -2057
rect 1458 -2188 1459 -2148
rect 170 -2188 171 -2150
rect 1689 -2188 1690 -2150
rect 219 -2153 220 -2057
rect 443 -2188 444 -2152
rect 471 -2153 472 -2057
rect 908 -2153 909 -2057
rect 1185 -2153 1186 -2057
rect 1241 -2188 1242 -2152
rect 198 -2155 199 -2057
rect 219 -2188 220 -2154
rect 226 -2155 227 -2057
rect 247 -2188 248 -2154
rect 362 -2188 363 -2154
rect 464 -2188 465 -2154
rect 492 -2155 493 -2057
rect 492 -2188 493 -2154
rect 492 -2155 493 -2057
rect 492 -2188 493 -2154
rect 520 -2155 521 -2057
rect 646 -2188 647 -2154
rect 751 -2155 752 -2057
rect 1122 -2188 1123 -2154
rect 1164 -2155 1165 -2057
rect 1185 -2188 1186 -2154
rect 198 -2188 199 -2156
rect 1755 -2188 1756 -2156
rect 226 -2188 227 -2158
rect 1430 -2159 1431 -2057
rect 229 -2188 230 -2160
rect 471 -2188 472 -2160
rect 513 -2161 514 -2057
rect 520 -2188 521 -2160
rect 583 -2161 584 -2057
rect 653 -2188 654 -2160
rect 751 -2188 752 -2160
rect 828 -2161 829 -2057
rect 1150 -2161 1151 -2057
rect 1164 -2188 1165 -2160
rect 65 -2163 66 -2057
rect 513 -2188 514 -2162
rect 583 -2188 584 -2162
rect 695 -2163 696 -2057
rect 1136 -2163 1137 -2057
rect 1150 -2188 1151 -2162
rect 65 -2188 66 -2164
rect 1024 -2165 1025 -2057
rect 415 -2188 416 -2166
rect 978 -2188 979 -2166
rect 982 -2167 983 -2057
rect 1136 -2188 1137 -2166
rect 600 -2169 601 -2057
rect 1430 -2188 1431 -2168
rect 625 -2188 626 -2170
rect 891 -2171 892 -2057
rect 961 -2171 962 -2057
rect 1024 -2188 1025 -2170
rect 695 -2188 696 -2172
rect 709 -2173 710 -2057
rect 849 -2173 850 -2057
rect 891 -2188 892 -2172
rect 975 -2173 976 -2057
rect 982 -2188 983 -2172
rect 282 -2175 283 -2057
rect 709 -2188 710 -2174
rect 849 -2188 850 -2174
rect 863 -2175 864 -2057
rect 282 -2188 283 -2176
rect 401 -2177 402 -2057
rect 639 -2177 640 -2057
rect 863 -2188 864 -2176
rect 72 -2179 73 -2057
rect 639 -2188 640 -2178
rect 702 -2179 703 -2057
rect 961 -2188 962 -2178
rect 72 -2188 73 -2180
rect 933 -2181 934 -2057
rect 380 -2183 381 -2057
rect 401 -2188 402 -2182
rect 702 -2188 703 -2182
rect 793 -2183 794 -2057
rect 933 -2188 934 -2182
rect 1269 -2188 1270 -2182
rect 380 -2188 381 -2184
rect 450 -2185 451 -2057
rect 450 -2188 451 -2186
rect 660 -2188 661 -2186
rect 30 -2198 31 -2196
rect 450 -2198 451 -2196
rect 453 -2198 454 -2196
rect 653 -2198 654 -2196
rect 688 -2198 689 -2196
rect 793 -2198 794 -2196
rect 796 -2198 797 -2196
rect 1395 -2198 1396 -2196
rect 1437 -2198 1438 -2196
rect 1437 -2323 1438 -2197
rect 1437 -2198 1438 -2196
rect 1437 -2323 1438 -2197
rect 1500 -2198 1501 -2196
rect 1500 -2323 1501 -2197
rect 1500 -2198 1501 -2196
rect 1500 -2323 1501 -2197
rect 1535 -2198 1536 -2196
rect 1535 -2323 1536 -2197
rect 1535 -2198 1536 -2196
rect 1535 -2323 1536 -2197
rect 1570 -2198 1571 -2196
rect 1570 -2323 1571 -2197
rect 1570 -2198 1571 -2196
rect 1570 -2323 1571 -2197
rect 1640 -2198 1641 -2196
rect 1706 -2323 1707 -2197
rect 1752 -2198 1753 -2196
rect 1766 -2198 1767 -2196
rect 44 -2200 45 -2196
rect 870 -2200 871 -2196
rect 873 -2200 874 -2196
rect 1465 -2200 1466 -2196
rect 1640 -2323 1641 -2199
rect 1696 -2200 1697 -2196
rect 51 -2202 52 -2196
rect 72 -2202 73 -2196
rect 89 -2202 90 -2196
rect 103 -2280 104 -2201
rect 117 -2323 118 -2201
rect 1444 -2202 1445 -2196
rect 1465 -2323 1466 -2201
rect 1514 -2202 1515 -2196
rect 1647 -2202 1648 -2196
rect 1647 -2323 1648 -2201
rect 1647 -2202 1648 -2196
rect 1647 -2323 1648 -2201
rect 1682 -2202 1683 -2196
rect 1713 -2323 1714 -2201
rect 51 -2323 52 -2203
rect 394 -2204 395 -2196
rect 408 -2323 409 -2203
rect 779 -2204 780 -2196
rect 786 -2204 787 -2196
rect 814 -2204 815 -2196
rect 828 -2204 829 -2196
rect 1367 -2204 1368 -2196
rect 1514 -2323 1515 -2203
rect 1549 -2204 1550 -2196
rect 1682 -2323 1683 -2203
rect 1717 -2204 1718 -2196
rect 58 -2206 59 -2196
rect 957 -2323 958 -2205
rect 978 -2206 979 -2196
rect 1423 -2206 1424 -2196
rect 1549 -2323 1550 -2205
rect 1591 -2206 1592 -2196
rect 1696 -2323 1697 -2205
rect 1738 -2206 1739 -2196
rect 58 -2323 59 -2207
rect 639 -2208 640 -2196
rect 691 -2323 692 -2207
rect 716 -2208 717 -2196
rect 723 -2208 724 -2196
rect 1346 -2208 1347 -2196
rect 1423 -2323 1424 -2207
rect 1472 -2208 1473 -2196
rect 1738 -2323 1739 -2207
rect 1759 -2208 1760 -2196
rect 65 -2323 66 -2209
rect 604 -2210 605 -2196
rect 607 -2210 608 -2196
rect 807 -2210 808 -2196
rect 814 -2323 815 -2209
rect 821 -2210 822 -2196
rect 828 -2323 829 -2209
rect 842 -2210 843 -2196
rect 852 -2323 853 -2209
rect 1031 -2210 1032 -2196
rect 1118 -2210 1119 -2196
rect 1661 -2210 1662 -2196
rect 68 -2212 69 -2196
rect 562 -2212 563 -2196
rect 590 -2212 591 -2196
rect 590 -2323 591 -2211
rect 590 -2212 591 -2196
rect 590 -2323 591 -2211
rect 611 -2212 612 -2196
rect 747 -2212 748 -2196
rect 758 -2323 759 -2211
rect 1129 -2212 1130 -2196
rect 1146 -2323 1147 -2211
rect 1731 -2212 1732 -2196
rect 72 -2323 73 -2213
rect 121 -2214 122 -2196
rect 131 -2214 132 -2196
rect 1017 -2214 1018 -2196
rect 1031 -2323 1032 -2213
rect 1101 -2214 1102 -2196
rect 1129 -2323 1130 -2213
rect 1206 -2214 1207 -2196
rect 1227 -2214 1228 -2196
rect 1731 -2323 1732 -2213
rect 89 -2323 90 -2215
rect 177 -2216 178 -2196
rect 184 -2216 185 -2196
rect 604 -2323 605 -2215
rect 618 -2216 619 -2196
rect 1367 -2323 1368 -2215
rect 1507 -2216 1508 -2196
rect 1661 -2323 1662 -2215
rect 93 -2323 94 -2217
rect 884 -2218 885 -2196
rect 891 -2218 892 -2196
rect 936 -2218 937 -2196
rect 999 -2218 1000 -2196
rect 1276 -2218 1277 -2196
rect 1335 -2323 1336 -2217
rect 1654 -2218 1655 -2196
rect 96 -2220 97 -2196
rect 1122 -2220 1123 -2196
rect 1192 -2220 1193 -2196
rect 1395 -2323 1396 -2219
rect 96 -2323 97 -2221
rect 184 -2323 185 -2221
rect 226 -2323 227 -2221
rect 415 -2222 416 -2196
rect 450 -2323 451 -2221
rect 646 -2222 647 -2196
rect 695 -2222 696 -2196
rect 730 -2222 731 -2196
rect 733 -2222 734 -2196
rect 1703 -2222 1704 -2196
rect 121 -2323 122 -2223
rect 233 -2224 234 -2196
rect 236 -2323 237 -2223
rect 793 -2323 794 -2223
rect 807 -2323 808 -2223
rect 835 -2224 836 -2196
rect 842 -2323 843 -2223
rect 877 -2224 878 -2196
rect 884 -2323 885 -2223
rect 1066 -2224 1067 -2196
rect 1122 -2323 1123 -2223
rect 1745 -2224 1746 -2196
rect 142 -2226 143 -2196
rect 145 -2280 146 -2225
rect 152 -2226 153 -2196
rect 1444 -2323 1445 -2225
rect 142 -2323 143 -2227
rect 625 -2228 626 -2196
rect 639 -2323 640 -2227
rect 1038 -2228 1039 -2196
rect 1066 -2323 1067 -2227
rect 1755 -2228 1756 -2196
rect 170 -2230 171 -2196
rect 317 -2230 318 -2196
rect 362 -2230 363 -2196
rect 873 -2323 874 -2229
rect 877 -2323 878 -2229
rect 905 -2230 906 -2196
rect 933 -2230 934 -2196
rect 1283 -2230 1284 -2196
rect 1346 -2323 1347 -2229
rect 1402 -2230 1403 -2196
rect 170 -2323 171 -2231
rect 523 -2232 524 -2196
rect 569 -2232 570 -2196
rect 695 -2323 696 -2231
rect 702 -2232 703 -2196
rect 1633 -2232 1634 -2196
rect 177 -2323 178 -2233
rect 205 -2234 206 -2196
rect 229 -2234 230 -2196
rect 954 -2234 955 -2196
rect 999 -2323 1000 -2233
rect 1717 -2323 1718 -2233
rect 205 -2323 206 -2235
rect 345 -2236 346 -2196
rect 464 -2236 465 -2196
rect 611 -2323 612 -2235
rect 618 -2323 619 -2235
rect 674 -2236 675 -2196
rect 702 -2323 703 -2235
rect 1213 -2236 1214 -2196
rect 1227 -2323 1228 -2235
rect 1297 -2236 1298 -2196
rect 1339 -2236 1340 -2196
rect 1402 -2323 1403 -2235
rect 1626 -2236 1627 -2196
rect 1633 -2323 1634 -2235
rect 100 -2238 101 -2196
rect 674 -2323 675 -2237
rect 716 -2323 717 -2237
rect 751 -2238 752 -2196
rect 772 -2238 773 -2196
rect 1507 -2323 1508 -2237
rect 1612 -2238 1613 -2196
rect 1626 -2323 1627 -2237
rect 44 -2323 45 -2239
rect 772 -2323 773 -2239
rect 786 -2323 787 -2239
rect 800 -2240 801 -2196
rect 821 -2323 822 -2239
rect 849 -2240 850 -2196
rect 891 -2323 892 -2239
rect 1045 -2240 1046 -2196
rect 1206 -2323 1207 -2239
rect 1318 -2240 1319 -2196
rect 1339 -2323 1340 -2239
rect 1388 -2240 1389 -2196
rect 1542 -2240 1543 -2196
rect 1612 -2323 1613 -2239
rect 100 -2323 101 -2241
rect 135 -2242 136 -2196
rect 191 -2242 192 -2196
rect 345 -2323 346 -2241
rect 422 -2242 423 -2196
rect 464 -2323 465 -2241
rect 471 -2242 472 -2196
rect 562 -2323 563 -2241
rect 569 -2323 570 -2241
rect 1059 -2242 1060 -2196
rect 1213 -2323 1214 -2241
rect 1255 -2242 1256 -2196
rect 1276 -2323 1277 -2241
rect 1486 -2242 1487 -2196
rect 1542 -2323 1543 -2241
rect 1577 -2242 1578 -2196
rect 135 -2323 136 -2243
rect 1619 -2244 1620 -2196
rect 191 -2323 192 -2245
rect 240 -2246 241 -2196
rect 268 -2323 269 -2245
rect 555 -2246 556 -2196
rect 586 -2323 587 -2245
rect 1192 -2323 1193 -2245
rect 1237 -2323 1238 -2245
rect 1675 -2246 1676 -2196
rect 107 -2248 108 -2196
rect 240 -2323 241 -2247
rect 271 -2248 272 -2196
rect 541 -2248 542 -2196
rect 548 -2248 549 -2196
rect 555 -2323 556 -2247
rect 646 -2323 647 -2247
rect 660 -2248 661 -2196
rect 730 -2323 731 -2247
rect 1472 -2323 1473 -2247
rect 1486 -2323 1487 -2247
rect 1521 -2248 1522 -2196
rect 1577 -2323 1578 -2247
rect 1703 -2323 1704 -2247
rect 107 -2323 108 -2249
rect 163 -2250 164 -2196
rect 233 -2323 234 -2249
rect 261 -2250 262 -2196
rect 282 -2250 283 -2196
rect 775 -2250 776 -2196
rect 800 -2323 801 -2249
rect 926 -2250 927 -2196
rect 933 -2323 934 -2249
rect 968 -2250 969 -2196
rect 1003 -2250 1004 -2196
rect 1101 -2323 1102 -2249
rect 1255 -2323 1256 -2249
rect 1430 -2250 1431 -2196
rect 1521 -2323 1522 -2249
rect 1724 -2250 1725 -2196
rect 114 -2252 115 -2196
rect 261 -2323 262 -2251
rect 282 -2323 283 -2251
rect 436 -2252 437 -2196
rect 506 -2252 507 -2196
rect 733 -2323 734 -2251
rect 737 -2252 738 -2196
rect 779 -2323 780 -2251
rect 835 -2323 836 -2251
rect 961 -2252 962 -2196
rect 1003 -2323 1004 -2251
rect 1150 -2252 1151 -2196
rect 1283 -2323 1284 -2251
rect 1416 -2252 1417 -2196
rect 163 -2323 164 -2253
rect 632 -2254 633 -2196
rect 656 -2323 657 -2253
rect 660 -2323 661 -2253
rect 747 -2323 748 -2253
rect 1675 -2323 1676 -2253
rect 215 -2323 216 -2255
rect 737 -2323 738 -2255
rect 751 -2323 752 -2255
rect 856 -2256 857 -2196
rect 898 -2256 899 -2196
rect 961 -2323 962 -2255
rect 1010 -2256 1011 -2196
rect 1360 -2256 1361 -2196
rect 1388 -2323 1389 -2255
rect 1598 -2256 1599 -2196
rect 156 -2258 157 -2196
rect 898 -2323 899 -2257
rect 905 -2323 906 -2257
rect 919 -2258 920 -2196
rect 926 -2323 927 -2257
rect 1024 -2258 1025 -2196
rect 1038 -2323 1039 -2257
rect 1199 -2258 1200 -2196
rect 1290 -2258 1291 -2196
rect 1724 -2323 1725 -2257
rect 156 -2323 157 -2259
rect 534 -2260 535 -2196
rect 541 -2323 542 -2259
rect 982 -2260 983 -2196
rect 1010 -2323 1011 -2259
rect 1108 -2260 1109 -2196
rect 1199 -2323 1200 -2259
rect 1234 -2260 1235 -2196
rect 1290 -2323 1291 -2259
rect 1374 -2260 1375 -2196
rect 1584 -2260 1585 -2196
rect 1598 -2323 1599 -2259
rect 128 -2262 129 -2196
rect 1584 -2323 1585 -2261
rect 40 -2264 41 -2196
rect 128 -2323 129 -2263
rect 289 -2264 290 -2196
rect 625 -2323 626 -2263
rect 761 -2264 762 -2196
rect 919 -2323 920 -2263
rect 982 -2323 983 -2263
rect 1136 -2264 1137 -2196
rect 1297 -2323 1298 -2263
rect 1381 -2264 1382 -2196
rect 173 -2266 174 -2196
rect 1381 -2323 1382 -2265
rect 173 -2323 174 -2267
rect 901 -2323 902 -2267
rect 1013 -2268 1014 -2196
rect 1024 -2323 1025 -2267
rect 1045 -2323 1046 -2267
rect 1094 -2268 1095 -2196
rect 1108 -2323 1109 -2267
rect 1668 -2268 1669 -2196
rect 289 -2323 290 -2269
rect 380 -2270 381 -2196
rect 436 -2323 437 -2269
rect 513 -2270 514 -2196
rect 520 -2270 521 -2196
rect 1619 -2323 1620 -2269
rect 1668 -2323 1669 -2269
rect 1710 -2270 1711 -2196
rect 114 -2323 115 -2271
rect 513 -2323 514 -2271
rect 548 -2323 549 -2271
rect 681 -2272 682 -2196
rect 849 -2323 850 -2271
rect 1654 -2323 1655 -2271
rect 149 -2274 150 -2196
rect 520 -2323 521 -2273
rect 681 -2323 682 -2273
rect 831 -2274 832 -2196
rect 1017 -2323 1018 -2273
rect 1052 -2274 1053 -2196
rect 1059 -2323 1060 -2273
rect 1185 -2274 1186 -2196
rect 1318 -2323 1319 -2273
rect 1458 -2274 1459 -2196
rect 1591 -2323 1592 -2273
rect 1710 -2323 1711 -2273
rect 149 -2323 150 -2275
rect 254 -2276 255 -2196
rect 296 -2276 297 -2196
rect 359 -2276 360 -2196
rect 478 -2276 479 -2196
rect 632 -2323 633 -2275
rect 1052 -2323 1053 -2275
rect 1080 -2276 1081 -2196
rect 1094 -2323 1095 -2275
rect 1563 -2276 1564 -2196
rect 219 -2278 220 -2196
rect 380 -2323 381 -2277
rect 478 -2323 479 -2277
rect 597 -2278 598 -2196
rect 1073 -2278 1074 -2196
rect 1150 -2323 1151 -2277
rect 1185 -2323 1186 -2277
rect 1248 -2278 1249 -2196
rect 1332 -2278 1333 -2196
rect 1416 -2323 1417 -2277
rect 1458 -2323 1459 -2277
rect 1479 -2278 1480 -2196
rect 1556 -2278 1557 -2196
rect 1563 -2323 1564 -2277
rect 219 -2323 220 -2279
rect 247 -2280 248 -2196
rect 254 -2323 255 -2279
rect 296 -2323 297 -2279
rect 709 -2280 710 -2196
rect 1073 -2323 1074 -2279
rect 1164 -2280 1165 -2196
rect 1353 -2280 1354 -2196
rect 1430 -2323 1431 -2279
rect 1479 -2323 1480 -2279
rect 1528 -2280 1529 -2196
rect 1556 -2323 1557 -2279
rect 1605 -2280 1606 -2196
rect 79 -2282 80 -2196
rect 247 -2323 248 -2281
rect 303 -2282 304 -2196
rect 394 -2323 395 -2281
rect 457 -2282 458 -2196
rect 709 -2323 710 -2281
rect 968 -2323 969 -2281
rect 1353 -2323 1354 -2281
rect 1360 -2323 1361 -2281
rect 1409 -2282 1410 -2196
rect 1493 -2282 1494 -2196
rect 1605 -2323 1606 -2281
rect 79 -2323 80 -2283
rect 198 -2284 199 -2196
rect 310 -2284 311 -2196
rect 975 -2284 976 -2196
rect 1136 -2323 1137 -2283
rect 1262 -2284 1263 -2196
rect 1304 -2284 1305 -2196
rect 1528 -2323 1529 -2283
rect 86 -2286 87 -2196
rect 457 -2323 458 -2285
rect 492 -2286 493 -2196
rect 534 -2323 535 -2285
rect 723 -2323 724 -2285
rect 1304 -2323 1305 -2285
rect 1374 -2323 1375 -2285
rect 1451 -2286 1452 -2196
rect 1493 -2323 1494 -2285
rect 1689 -2286 1690 -2196
rect 138 -2323 139 -2287
rect 303 -2323 304 -2287
rect 310 -2323 311 -2287
rect 485 -2288 486 -2196
rect 499 -2288 500 -2196
rect 506 -2323 507 -2287
rect 653 -2323 654 -2287
rect 1689 -2323 1690 -2287
rect 198 -2323 199 -2289
rect 1104 -2290 1105 -2196
rect 1157 -2290 1158 -2196
rect 1248 -2323 1249 -2289
rect 1269 -2290 1270 -2196
rect 1451 -2323 1452 -2289
rect 317 -2323 318 -2291
rect 688 -2323 689 -2291
rect 744 -2292 745 -2196
rect 1409 -2323 1410 -2291
rect 324 -2294 325 -2196
rect 856 -2323 857 -2293
rect 975 -2323 976 -2293
rect 989 -2294 990 -2196
rect 1083 -2323 1084 -2293
rect 1262 -2323 1263 -2293
rect 324 -2323 325 -2295
rect 366 -2296 367 -2196
rect 373 -2296 374 -2196
rect 485 -2323 486 -2295
rect 499 -2323 500 -2295
rect 863 -2296 864 -2196
rect 989 -2323 990 -2295
rect 1311 -2296 1312 -2196
rect 275 -2298 276 -2196
rect 366 -2323 367 -2297
rect 429 -2298 430 -2196
rect 492 -2323 493 -2297
rect 744 -2323 745 -2297
rect 947 -2298 948 -2196
rect 954 -2323 955 -2297
rect 1311 -2323 1312 -2297
rect 212 -2300 213 -2196
rect 275 -2323 276 -2299
rect 331 -2300 332 -2196
rect 422 -2323 423 -2299
rect 429 -2323 430 -2299
rect 705 -2300 706 -2196
rect 863 -2323 864 -2299
rect 1143 -2300 1144 -2196
rect 1157 -2323 1158 -2299
rect 1220 -2300 1221 -2196
rect 331 -2323 332 -2301
rect 1115 -2302 1116 -2196
rect 1164 -2323 1165 -2301
rect 1241 -2302 1242 -2196
rect 338 -2304 339 -2196
rect 373 -2323 374 -2303
rect 415 -2323 416 -2303
rect 705 -2323 706 -2303
rect 912 -2304 913 -2196
rect 1115 -2323 1116 -2303
rect 1171 -2304 1172 -2196
rect 1220 -2323 1221 -2303
rect 1241 -2323 1242 -2303
rect 1325 -2304 1326 -2196
rect 338 -2323 339 -2305
rect 401 -2306 402 -2196
rect 912 -2323 913 -2305
rect 940 -2306 941 -2196
rect 947 -2323 948 -2305
rect 1332 -2323 1333 -2305
rect 352 -2308 353 -2196
rect 401 -2323 402 -2307
rect 940 -2323 941 -2307
rect 1087 -2308 1088 -2196
rect 1143 -2323 1144 -2307
rect 1325 -2323 1326 -2307
rect 352 -2323 353 -2309
rect 576 -2310 577 -2196
rect 1087 -2323 1088 -2309
rect 1178 -2310 1179 -2196
rect 359 -2323 360 -2311
rect 387 -2312 388 -2196
rect 576 -2323 577 -2311
rect 667 -2312 668 -2196
rect 996 -2312 997 -2196
rect 1178 -2323 1179 -2311
rect 387 -2323 388 -2313
rect 527 -2314 528 -2196
rect 667 -2323 668 -2313
rect 765 -2314 766 -2196
rect 996 -2323 997 -2313
rect 1269 -2323 1270 -2313
rect 443 -2316 444 -2196
rect 765 -2323 766 -2315
rect 443 -2323 444 -2317
rect 583 -2318 584 -2196
rect 471 -2323 472 -2319
rect 583 -2323 584 -2319
rect 527 -2323 528 -2321
rect 870 -2323 871 -2321
rect 51 -2333 52 -2331
rect 180 -2438 181 -2332
rect 215 -2333 216 -2331
rect 975 -2333 976 -2331
rect 982 -2333 983 -2331
rect 996 -2333 997 -2331
rect 999 -2333 1000 -2331
rect 1486 -2333 1487 -2331
rect 1514 -2333 1515 -2331
rect 1538 -2438 1539 -2332
rect 1605 -2333 1606 -2331
rect 1706 -2333 1707 -2331
rect 51 -2438 52 -2334
rect 226 -2335 227 -2331
rect 443 -2335 444 -2331
rect 824 -2438 825 -2334
rect 856 -2335 857 -2331
rect 971 -2335 972 -2331
rect 982 -2438 983 -2334
rect 1045 -2335 1046 -2331
rect 1076 -2438 1077 -2334
rect 1437 -2335 1438 -2331
rect 1493 -2335 1494 -2331
rect 1514 -2438 1515 -2334
rect 1605 -2438 1606 -2334
rect 1675 -2335 1676 -2331
rect 79 -2337 80 -2331
rect 702 -2337 703 -2331
rect 733 -2337 734 -2331
rect 1122 -2337 1123 -2331
rect 1171 -2337 1172 -2331
rect 1451 -2337 1452 -2331
rect 1612 -2337 1613 -2331
rect 1675 -2438 1676 -2336
rect 79 -2438 80 -2338
rect 93 -2339 94 -2331
rect 100 -2339 101 -2331
rect 1125 -2339 1126 -2331
rect 1171 -2438 1172 -2338
rect 1178 -2339 1179 -2331
rect 1244 -2438 1245 -2338
rect 1668 -2339 1669 -2331
rect 86 -2341 87 -2331
rect 1689 -2341 1690 -2331
rect 86 -2438 87 -2342
rect 128 -2343 129 -2331
rect 135 -2343 136 -2331
rect 380 -2343 381 -2331
rect 415 -2343 416 -2331
rect 443 -2438 444 -2342
rect 450 -2343 451 -2331
rect 583 -2343 584 -2331
rect 597 -2343 598 -2331
rect 656 -2343 657 -2331
rect 660 -2343 661 -2331
rect 677 -2438 678 -2342
rect 684 -2438 685 -2342
rect 1584 -2343 1585 -2331
rect 93 -2438 94 -2344
rect 422 -2345 423 -2331
rect 464 -2345 465 -2331
rect 467 -2357 468 -2344
rect 492 -2345 493 -2331
rect 730 -2345 731 -2331
rect 775 -2345 776 -2331
rect 1395 -2345 1396 -2331
rect 1437 -2438 1438 -2344
rect 1472 -2345 1473 -2331
rect 100 -2438 101 -2346
rect 261 -2347 262 -2331
rect 345 -2347 346 -2331
rect 450 -2438 451 -2346
rect 457 -2347 458 -2331
rect 492 -2438 493 -2346
rect 502 -2438 503 -2346
rect 534 -2347 535 -2331
rect 548 -2347 549 -2331
rect 583 -2438 584 -2346
rect 597 -2438 598 -2346
rect 642 -2347 643 -2331
rect 691 -2347 692 -2331
rect 1563 -2347 1564 -2331
rect 65 -2349 66 -2331
rect 457 -2438 458 -2348
rect 464 -2438 465 -2348
rect 485 -2349 486 -2331
rect 527 -2349 528 -2331
rect 1045 -2438 1046 -2348
rect 1080 -2349 1081 -2331
rect 1528 -2349 1529 -2331
rect 1556 -2349 1557 -2331
rect 1563 -2438 1564 -2348
rect 65 -2438 66 -2350
rect 149 -2351 150 -2331
rect 163 -2351 164 -2331
rect 236 -2351 237 -2331
rect 240 -2351 241 -2331
rect 380 -2438 381 -2350
rect 422 -2438 423 -2350
rect 730 -2438 731 -2350
rect 733 -2438 734 -2350
rect 1472 -2438 1473 -2350
rect 1521 -2351 1522 -2331
rect 1556 -2438 1557 -2350
rect 96 -2353 97 -2331
rect 1528 -2438 1529 -2352
rect 107 -2355 108 -2331
rect 534 -2438 535 -2354
rect 548 -2438 549 -2354
rect 562 -2355 563 -2331
rect 569 -2355 570 -2331
rect 653 -2355 654 -2331
rect 800 -2355 801 -2331
rect 1195 -2438 1196 -2354
rect 1248 -2355 1249 -2331
rect 1248 -2438 1249 -2354
rect 1248 -2355 1249 -2331
rect 1248 -2438 1249 -2354
rect 1304 -2355 1305 -2331
rect 1626 -2355 1627 -2331
rect 107 -2438 108 -2356
rect 138 -2357 139 -2331
rect 149 -2438 150 -2356
rect 205 -2357 206 -2331
rect 212 -2357 213 -2331
rect 415 -2438 416 -2356
rect 485 -2438 486 -2356
rect 530 -2438 531 -2356
rect 975 -2438 976 -2356
rect 989 -2357 990 -2331
rect 1584 -2438 1585 -2356
rect 58 -2359 59 -2331
rect 205 -2438 206 -2358
rect 212 -2438 213 -2358
rect 1192 -2359 1193 -2331
rect 1304 -2438 1305 -2358
rect 1353 -2359 1354 -2331
rect 1384 -2438 1385 -2358
rect 1570 -2359 1571 -2331
rect 114 -2361 115 -2331
rect 499 -2361 500 -2331
rect 576 -2361 577 -2331
rect 660 -2438 661 -2360
rect 779 -2361 780 -2331
rect 800 -2438 801 -2360
rect 856 -2438 857 -2360
rect 1633 -2361 1634 -2331
rect 44 -2363 45 -2331
rect 576 -2438 577 -2362
rect 618 -2363 619 -2331
rect 688 -2363 689 -2331
rect 695 -2363 696 -2331
rect 779 -2438 780 -2362
rect 863 -2363 864 -2331
rect 1146 -2363 1147 -2331
rect 1178 -2438 1179 -2362
rect 1307 -2363 1308 -2331
rect 1314 -2438 1315 -2362
rect 1696 -2363 1697 -2331
rect 114 -2438 115 -2364
rect 359 -2365 360 -2331
rect 432 -2438 433 -2364
rect 618 -2438 619 -2364
rect 625 -2365 626 -2331
rect 1486 -2438 1487 -2364
rect 1521 -2438 1522 -2364
rect 1654 -2365 1655 -2331
rect 117 -2367 118 -2331
rect 233 -2438 234 -2366
rect 240 -2438 241 -2366
rect 387 -2367 388 -2331
rect 471 -2367 472 -2331
rect 562 -2438 563 -2366
rect 590 -2367 591 -2331
rect 625 -2438 626 -2366
rect 632 -2367 633 -2331
rect 747 -2367 748 -2331
rect 863 -2438 864 -2366
rect 1143 -2367 1144 -2331
rect 1283 -2367 1284 -2331
rect 1353 -2438 1354 -2366
rect 1388 -2367 1389 -2331
rect 1493 -2438 1494 -2366
rect 1570 -2438 1571 -2366
rect 1598 -2367 1599 -2331
rect 128 -2438 129 -2368
rect 156 -2369 157 -2331
rect 163 -2438 164 -2368
rect 835 -2369 836 -2331
rect 870 -2438 871 -2368
rect 877 -2369 878 -2331
rect 898 -2369 899 -2331
rect 1682 -2369 1683 -2331
rect 135 -2438 136 -2370
rect 604 -2371 605 -2331
rect 632 -2438 633 -2370
rect 947 -2371 948 -2331
rect 954 -2371 955 -2331
rect 1661 -2371 1662 -2331
rect 142 -2373 143 -2331
rect 877 -2438 878 -2372
rect 898 -2438 899 -2372
rect 1311 -2373 1312 -2331
rect 1332 -2373 1333 -2331
rect 1647 -2373 1648 -2331
rect 142 -2438 143 -2374
rect 478 -2375 479 -2331
rect 499 -2438 500 -2374
rect 1083 -2375 1084 -2331
rect 1097 -2375 1098 -2331
rect 1255 -2375 1256 -2331
rect 1388 -2438 1389 -2374
rect 1409 -2375 1410 -2331
rect 1451 -2438 1452 -2374
rect 1549 -2375 1550 -2331
rect 1598 -2438 1599 -2374
rect 1703 -2375 1704 -2331
rect 170 -2377 171 -2331
rect 520 -2377 521 -2331
rect 541 -2377 542 -2331
rect 747 -2438 748 -2376
rect 828 -2377 829 -2331
rect 835 -2438 836 -2376
rect 873 -2377 874 -2331
rect 1500 -2377 1501 -2331
rect 170 -2438 171 -2378
rect 198 -2379 199 -2331
rect 215 -2438 216 -2378
rect 674 -2379 675 -2331
rect 688 -2438 689 -2378
rect 723 -2379 724 -2331
rect 828 -2438 829 -2378
rect 1066 -2379 1067 -2331
rect 1080 -2438 1081 -2378
rect 1101 -2379 1102 -2331
rect 1108 -2379 1109 -2331
rect 1500 -2438 1501 -2378
rect 156 -2438 157 -2380
rect 674 -2438 675 -2380
rect 695 -2438 696 -2380
rect 709 -2381 710 -2331
rect 723 -2438 724 -2380
rect 814 -2381 815 -2331
rect 905 -2381 906 -2331
rect 905 -2438 906 -2380
rect 905 -2381 906 -2331
rect 905 -2438 906 -2380
rect 919 -2381 920 -2331
rect 989 -2438 990 -2380
rect 996 -2438 997 -2380
rect 1031 -2381 1032 -2331
rect 1066 -2438 1067 -2380
rect 1150 -2381 1151 -2331
rect 1192 -2438 1193 -2380
rect 1283 -2438 1284 -2380
rect 1395 -2438 1396 -2380
rect 1423 -2381 1424 -2331
rect 198 -2438 199 -2382
rect 296 -2383 297 -2331
rect 345 -2438 346 -2382
rect 373 -2383 374 -2331
rect 387 -2438 388 -2382
rect 474 -2438 475 -2382
rect 478 -2438 479 -2382
rect 681 -2383 682 -2331
rect 709 -2438 710 -2382
rect 716 -2383 717 -2331
rect 793 -2383 794 -2331
rect 1101 -2438 1102 -2382
rect 1122 -2438 1123 -2382
rect 1129 -2383 1130 -2331
rect 1143 -2438 1144 -2382
rect 1199 -2383 1200 -2331
rect 1255 -2438 1256 -2382
rect 1339 -2383 1340 -2331
rect 1374 -2383 1375 -2331
rect 1423 -2438 1424 -2382
rect 226 -2438 227 -2384
rect 247 -2385 248 -2331
rect 254 -2385 255 -2331
rect 261 -2438 262 -2384
rect 268 -2385 269 -2331
rect 569 -2438 570 -2384
rect 590 -2438 591 -2384
rect 611 -2385 612 -2331
rect 639 -2438 640 -2384
rect 1619 -2385 1620 -2331
rect 184 -2387 185 -2331
rect 247 -2438 248 -2386
rect 254 -2438 255 -2386
rect 401 -2387 402 -2331
rect 471 -2438 472 -2386
rect 765 -2387 766 -2331
rect 786 -2387 787 -2331
rect 793 -2438 794 -2386
rect 919 -2438 920 -2386
rect 1213 -2387 1214 -2331
rect 1339 -2438 1340 -2386
rect 1360 -2387 1361 -2331
rect 1374 -2438 1375 -2386
rect 1444 -2387 1445 -2331
rect 184 -2438 185 -2388
rect 849 -2389 850 -2331
rect 901 -2389 902 -2331
rect 1444 -2438 1445 -2388
rect 268 -2438 269 -2390
rect 429 -2391 430 -2331
rect 513 -2391 514 -2331
rect 1150 -2438 1151 -2390
rect 1185 -2391 1186 -2331
rect 1213 -2438 1214 -2390
rect 1360 -2438 1361 -2390
rect 1402 -2391 1403 -2331
rect 1409 -2438 1410 -2390
rect 1479 -2391 1480 -2331
rect 282 -2393 283 -2331
rect 513 -2438 514 -2392
rect 520 -2438 521 -2392
rect 744 -2393 745 -2331
rect 786 -2438 787 -2392
rect 821 -2393 822 -2331
rect 901 -2438 902 -2392
rect 1430 -2393 1431 -2331
rect 1479 -2438 1480 -2392
rect 1577 -2393 1578 -2331
rect 282 -2438 283 -2394
rect 289 -2395 290 -2331
rect 296 -2438 297 -2394
rect 772 -2395 773 -2331
rect 814 -2438 815 -2394
rect 849 -2438 850 -2394
rect 926 -2395 927 -2331
rect 954 -2438 955 -2394
rect 957 -2395 958 -2331
rect 1332 -2438 1333 -2394
rect 1346 -2395 1347 -2331
rect 1402 -2438 1403 -2394
rect 1430 -2438 1431 -2394
rect 1591 -2395 1592 -2331
rect 173 -2397 174 -2331
rect 289 -2438 290 -2396
rect 303 -2397 304 -2331
rect 401 -2438 402 -2396
rect 555 -2397 556 -2331
rect 611 -2438 612 -2396
rect 646 -2397 647 -2331
rect 765 -2438 766 -2396
rect 772 -2438 773 -2396
rect 852 -2438 853 -2396
rect 884 -2397 885 -2331
rect 926 -2438 927 -2396
rect 933 -2397 934 -2331
rect 947 -2438 948 -2396
rect 971 -2438 972 -2396
rect 1458 -2397 1459 -2331
rect 1577 -2438 1578 -2396
rect 1738 -2397 1739 -2331
rect 177 -2399 178 -2331
rect 303 -2438 304 -2398
rect 310 -2399 311 -2331
rect 555 -2438 556 -2398
rect 604 -2438 605 -2398
rect 751 -2399 752 -2331
rect 821 -2438 822 -2398
rect 1731 -2399 1732 -2331
rect 58 -2438 59 -2400
rect 310 -2438 311 -2400
rect 338 -2401 339 -2331
rect 373 -2438 374 -2400
rect 653 -2438 654 -2400
rect 667 -2401 668 -2331
rect 716 -2438 717 -2400
rect 737 -2401 738 -2331
rect 744 -2438 745 -2400
rect 912 -2401 913 -2331
rect 1024 -2401 1025 -2331
rect 1108 -2438 1109 -2400
rect 1115 -2401 1116 -2331
rect 1591 -2438 1592 -2400
rect 177 -2438 178 -2402
rect 436 -2403 437 -2331
rect 667 -2438 668 -2402
rect 807 -2403 808 -2331
rect 842 -2403 843 -2331
rect 884 -2438 885 -2402
rect 891 -2403 892 -2331
rect 912 -2438 913 -2402
rect 1017 -2403 1018 -2331
rect 1024 -2438 1025 -2402
rect 1031 -2438 1032 -2402
rect 1227 -2403 1228 -2331
rect 1318 -2403 1319 -2331
rect 1346 -2438 1347 -2402
rect 1458 -2438 1459 -2402
rect 1542 -2403 1543 -2331
rect 191 -2405 192 -2331
rect 338 -2438 339 -2404
rect 352 -2405 353 -2331
rect 646 -2438 647 -2404
rect 737 -2438 738 -2404
rect 810 -2438 811 -2404
rect 842 -2438 843 -2404
rect 1003 -2405 1004 -2331
rect 1038 -2405 1039 -2331
rect 1129 -2438 1130 -2404
rect 1136 -2405 1137 -2331
rect 1227 -2438 1228 -2404
rect 1535 -2405 1536 -2331
rect 1542 -2438 1543 -2404
rect 191 -2438 192 -2406
rect 331 -2407 332 -2331
rect 359 -2438 360 -2406
rect 366 -2407 367 -2331
rect 436 -2438 437 -2406
rect 506 -2407 507 -2331
rect 751 -2438 752 -2406
rect 968 -2438 969 -2406
rect 1003 -2438 1004 -2406
rect 1290 -2407 1291 -2331
rect 219 -2409 220 -2331
rect 352 -2438 353 -2408
rect 506 -2438 507 -2408
rect 541 -2438 542 -2408
rect 758 -2409 759 -2331
rect 1017 -2438 1018 -2408
rect 1038 -2438 1039 -2408
rect 1059 -2409 1060 -2331
rect 1115 -2438 1116 -2408
rect 1157 -2409 1158 -2331
rect 1185 -2438 1186 -2408
rect 1325 -2409 1326 -2331
rect 219 -2438 220 -2410
rect 317 -2411 318 -2331
rect 324 -2411 325 -2331
rect 366 -2438 367 -2410
rect 758 -2438 759 -2410
rect 1234 -2411 1235 -2331
rect 1290 -2438 1291 -2410
rect 1381 -2411 1382 -2331
rect 121 -2413 122 -2331
rect 317 -2438 318 -2412
rect 324 -2438 325 -2412
rect 807 -2438 808 -2412
rect 891 -2438 892 -2412
rect 1010 -2413 1011 -2331
rect 1059 -2438 1060 -2412
rect 1087 -2413 1088 -2331
rect 1136 -2438 1137 -2412
rect 1717 -2413 1718 -2331
rect 72 -2415 73 -2331
rect 121 -2438 122 -2414
rect 331 -2438 332 -2414
rect 614 -2438 615 -2414
rect 961 -2415 962 -2331
rect 1010 -2438 1011 -2414
rect 1073 -2415 1074 -2331
rect 1087 -2438 1088 -2414
rect 1157 -2438 1158 -2414
rect 1164 -2415 1165 -2331
rect 1199 -2438 1200 -2414
rect 1206 -2415 1207 -2331
rect 1220 -2415 1221 -2331
rect 1318 -2438 1319 -2414
rect 1325 -2438 1326 -2414
rect 1335 -2415 1336 -2331
rect 1381 -2438 1382 -2414
rect 1416 -2415 1417 -2331
rect 72 -2438 73 -2416
rect 1094 -2417 1095 -2331
rect 1164 -2438 1165 -2416
rect 1724 -2417 1725 -2331
rect 537 -2419 538 -2331
rect 1220 -2438 1221 -2418
rect 1234 -2438 1235 -2418
rect 1241 -2419 1242 -2331
rect 1276 -2419 1277 -2331
rect 1416 -2438 1417 -2418
rect 933 -2438 934 -2420
rect 1073 -2438 1074 -2420
rect 1206 -2438 1207 -2420
rect 1297 -2421 1298 -2331
rect 940 -2423 941 -2331
rect 1094 -2438 1095 -2422
rect 1241 -2438 1242 -2422
rect 1549 -2438 1550 -2422
rect 940 -2438 941 -2424
rect 1710 -2425 1711 -2331
rect 961 -2438 962 -2426
rect 1052 -2427 1053 -2331
rect 1262 -2427 1263 -2331
rect 1276 -2438 1277 -2426
rect 705 -2429 706 -2331
rect 1052 -2438 1053 -2428
rect 1262 -2438 1263 -2428
rect 1269 -2429 1270 -2331
rect 408 -2431 409 -2331
rect 705 -2438 706 -2430
rect 1269 -2438 1270 -2430
rect 1367 -2431 1368 -2331
rect 275 -2433 276 -2331
rect 408 -2438 409 -2432
rect 1367 -2438 1368 -2432
rect 1465 -2433 1466 -2331
rect 275 -2438 276 -2434
rect 394 -2435 395 -2331
rect 1465 -2438 1466 -2434
rect 1507 -2435 1508 -2331
rect 394 -2438 395 -2436
rect 845 -2438 846 -2436
rect 1507 -2438 1508 -2436
rect 1640 -2437 1641 -2331
rect 44 -2555 45 -2447
rect 163 -2448 164 -2446
rect 184 -2448 185 -2446
rect 649 -2555 650 -2447
rect 681 -2448 682 -2446
rect 744 -2555 745 -2447
rect 754 -2555 755 -2447
rect 779 -2448 780 -2446
rect 786 -2448 787 -2446
rect 873 -2555 874 -2447
rect 912 -2448 913 -2446
rect 1696 -2555 1697 -2447
rect 86 -2450 87 -2446
rect 177 -2555 178 -2449
rect 212 -2450 213 -2446
rect 212 -2555 213 -2449
rect 212 -2450 213 -2446
rect 212 -2555 213 -2449
rect 233 -2450 234 -2446
rect 233 -2555 234 -2449
rect 233 -2450 234 -2446
rect 233 -2555 234 -2449
rect 240 -2450 241 -2446
rect 859 -2450 860 -2446
rect 870 -2450 871 -2446
rect 912 -2555 913 -2449
rect 947 -2450 948 -2446
rect 947 -2555 948 -2449
rect 947 -2450 948 -2446
rect 947 -2555 948 -2449
rect 957 -2555 958 -2449
rect 996 -2450 997 -2446
rect 1062 -2555 1063 -2449
rect 1612 -2555 1613 -2449
rect 1675 -2450 1676 -2446
rect 1731 -2555 1732 -2449
rect 86 -2555 87 -2451
rect 597 -2452 598 -2446
rect 611 -2452 612 -2446
rect 1521 -2452 1522 -2446
rect 1528 -2452 1529 -2446
rect 1678 -2555 1679 -2451
rect 100 -2454 101 -2446
rect 240 -2555 241 -2453
rect 257 -2454 258 -2446
rect 681 -2555 682 -2453
rect 688 -2454 689 -2446
rect 740 -2555 741 -2453
rect 779 -2555 780 -2453
rect 800 -2454 801 -2446
rect 807 -2454 808 -2446
rect 954 -2454 955 -2446
rect 971 -2454 972 -2446
rect 1584 -2454 1585 -2446
rect 1605 -2454 1606 -2446
rect 1724 -2555 1725 -2453
rect 107 -2456 108 -2446
rect 870 -2555 871 -2455
rect 891 -2456 892 -2446
rect 996 -2555 997 -2455
rect 1076 -2456 1077 -2446
rect 1346 -2456 1347 -2446
rect 1367 -2456 1368 -2446
rect 1521 -2555 1522 -2455
rect 1538 -2456 1539 -2446
rect 1563 -2456 1564 -2446
rect 1577 -2456 1578 -2446
rect 1738 -2555 1739 -2455
rect 72 -2458 73 -2446
rect 107 -2555 108 -2457
rect 142 -2458 143 -2446
rect 166 -2555 167 -2457
rect 180 -2458 181 -2446
rect 800 -2555 801 -2457
rect 821 -2458 822 -2446
rect 1605 -2555 1606 -2457
rect 142 -2555 143 -2459
rect 628 -2555 629 -2459
rect 642 -2460 643 -2446
rect 1192 -2460 1193 -2446
rect 1227 -2460 1228 -2446
rect 1367 -2555 1368 -2459
rect 1381 -2460 1382 -2446
rect 1479 -2460 1480 -2446
rect 1500 -2460 1501 -2446
rect 1577 -2555 1578 -2459
rect 152 -2555 153 -2461
rect 1290 -2462 1291 -2446
rect 1300 -2462 1301 -2446
rect 1430 -2462 1431 -2446
rect 1458 -2462 1459 -2446
rect 1619 -2555 1620 -2461
rect 282 -2464 283 -2446
rect 551 -2555 552 -2463
rect 562 -2464 563 -2446
rect 611 -2555 612 -2463
rect 702 -2555 703 -2463
rect 828 -2464 829 -2446
rect 842 -2555 843 -2463
rect 1073 -2464 1074 -2446
rect 1115 -2464 1116 -2446
rect 1227 -2555 1228 -2463
rect 1244 -2464 1245 -2446
rect 1304 -2464 1305 -2446
rect 1311 -2464 1312 -2446
rect 1528 -2555 1529 -2463
rect 1556 -2464 1557 -2446
rect 1710 -2555 1711 -2463
rect 261 -2466 262 -2446
rect 282 -2555 283 -2465
rect 296 -2466 297 -2446
rect 471 -2555 472 -2465
rect 492 -2466 493 -2446
rect 562 -2555 563 -2465
rect 593 -2555 594 -2465
rect 1136 -2466 1137 -2446
rect 1157 -2466 1158 -2446
rect 1640 -2555 1641 -2465
rect 226 -2468 227 -2446
rect 261 -2555 262 -2467
rect 296 -2555 297 -2467
rect 352 -2468 353 -2446
rect 411 -2555 412 -2467
rect 464 -2468 465 -2446
rect 502 -2468 503 -2446
rect 1661 -2555 1662 -2467
rect 93 -2470 94 -2446
rect 352 -2555 353 -2469
rect 422 -2470 423 -2446
rect 464 -2555 465 -2469
rect 506 -2470 507 -2446
rect 688 -2555 689 -2469
rect 716 -2470 717 -2446
rect 828 -2555 829 -2469
rect 845 -2470 846 -2446
rect 1269 -2470 1270 -2446
rect 1276 -2470 1277 -2446
rect 1346 -2555 1347 -2469
rect 1395 -2470 1396 -2446
rect 1682 -2555 1683 -2469
rect 65 -2472 66 -2446
rect 93 -2555 94 -2471
rect 226 -2555 227 -2471
rect 317 -2472 318 -2446
rect 324 -2472 325 -2446
rect 499 -2472 500 -2446
rect 506 -2555 507 -2471
rect 684 -2472 685 -2446
rect 730 -2472 731 -2446
rect 1094 -2472 1095 -2446
rect 1129 -2472 1130 -2446
rect 1192 -2555 1193 -2471
rect 1199 -2472 1200 -2446
rect 1311 -2555 1312 -2471
rect 1314 -2472 1315 -2446
rect 1486 -2472 1487 -2446
rect 1507 -2472 1508 -2446
rect 1689 -2555 1690 -2471
rect 65 -2555 66 -2473
rect 79 -2474 80 -2446
rect 100 -2555 101 -2473
rect 317 -2555 318 -2473
rect 324 -2555 325 -2473
rect 408 -2474 409 -2446
rect 422 -2555 423 -2473
rect 485 -2474 486 -2446
rect 513 -2474 514 -2446
rect 541 -2474 542 -2446
rect 583 -2474 584 -2446
rect 716 -2555 717 -2473
rect 751 -2474 752 -2446
rect 1458 -2555 1459 -2473
rect 1465 -2474 1466 -2446
rect 1584 -2555 1585 -2473
rect 58 -2476 59 -2446
rect 485 -2555 486 -2475
rect 513 -2555 514 -2475
rect 590 -2476 591 -2446
rect 597 -2555 598 -2475
rect 653 -2476 654 -2446
rect 751 -2555 752 -2475
rect 1563 -2555 1564 -2475
rect 58 -2555 59 -2477
rect 632 -2478 633 -2446
rect 765 -2478 766 -2446
rect 891 -2555 892 -2477
rect 919 -2478 920 -2446
rect 1269 -2555 1270 -2477
rect 1276 -2555 1277 -2477
rect 1451 -2478 1452 -2446
rect 1507 -2555 1508 -2477
rect 1570 -2478 1571 -2446
rect 79 -2555 80 -2479
rect 345 -2480 346 -2446
rect 401 -2480 402 -2446
rect 765 -2555 766 -2479
rect 793 -2480 794 -2446
rect 807 -2555 808 -2479
rect 852 -2480 853 -2446
rect 1122 -2480 1123 -2446
rect 1129 -2555 1130 -2479
rect 1598 -2480 1599 -2446
rect 121 -2482 122 -2446
rect 401 -2555 402 -2481
rect 408 -2555 409 -2481
rect 898 -2482 899 -2446
rect 929 -2555 930 -2481
rect 1500 -2555 1501 -2481
rect 1514 -2482 1515 -2446
rect 1668 -2555 1669 -2481
rect 121 -2555 122 -2483
rect 128 -2484 129 -2446
rect 215 -2484 216 -2446
rect 1486 -2555 1487 -2483
rect 128 -2555 129 -2485
rect 149 -2486 150 -2446
rect 303 -2486 304 -2446
rect 432 -2486 433 -2446
rect 436 -2486 437 -2446
rect 492 -2555 493 -2485
rect 520 -2486 521 -2446
rect 674 -2486 675 -2446
rect 677 -2486 678 -2446
rect 1570 -2555 1571 -2485
rect 75 -2555 76 -2487
rect 436 -2555 437 -2487
rect 450 -2488 451 -2446
rect 653 -2555 654 -2487
rect 674 -2555 675 -2487
rect 786 -2555 787 -2487
rect 877 -2488 878 -2446
rect 898 -2555 899 -2487
rect 1024 -2488 1025 -2446
rect 1094 -2555 1095 -2487
rect 1167 -2555 1168 -2487
rect 1409 -2488 1410 -2446
rect 1416 -2488 1417 -2446
rect 1514 -2555 1515 -2487
rect 149 -2555 150 -2489
rect 184 -2555 185 -2489
rect 303 -2555 304 -2489
rect 387 -2490 388 -2446
rect 429 -2490 430 -2446
rect 1626 -2555 1627 -2489
rect 310 -2555 311 -2491
rect 373 -2492 374 -2446
rect 387 -2555 388 -2491
rect 457 -2492 458 -2446
rect 474 -2492 475 -2446
rect 499 -2555 500 -2491
rect 520 -2555 521 -2491
rect 961 -2492 962 -2446
rect 982 -2492 983 -2446
rect 1024 -2555 1025 -2491
rect 1031 -2492 1032 -2446
rect 1304 -2555 1305 -2491
rect 1332 -2492 1333 -2446
rect 1409 -2555 1410 -2491
rect 1472 -2492 1473 -2446
rect 1598 -2555 1599 -2491
rect 103 -2555 104 -2493
rect 373 -2555 374 -2493
rect 432 -2555 433 -2493
rect 1717 -2555 1718 -2493
rect 313 -2496 314 -2446
rect 359 -2496 360 -2446
rect 443 -2496 444 -2446
rect 450 -2555 451 -2495
rect 527 -2496 528 -2446
rect 569 -2496 570 -2446
rect 576 -2496 577 -2446
rect 1416 -2555 1417 -2495
rect 247 -2498 248 -2446
rect 359 -2555 360 -2497
rect 366 -2498 367 -2446
rect 527 -2555 528 -2497
rect 541 -2555 542 -2497
rect 723 -2498 724 -2446
rect 877 -2555 878 -2497
rect 894 -2498 895 -2446
rect 933 -2498 934 -2446
rect 961 -2555 962 -2497
rect 1031 -2555 1032 -2497
rect 1188 -2555 1189 -2497
rect 1199 -2555 1200 -2497
rect 1255 -2498 1256 -2446
rect 1290 -2555 1291 -2497
rect 1388 -2498 1389 -2446
rect 1395 -2555 1396 -2497
rect 1549 -2498 1550 -2446
rect 219 -2500 220 -2446
rect 247 -2555 248 -2499
rect 275 -2500 276 -2446
rect 366 -2555 367 -2499
rect 415 -2500 416 -2446
rect 443 -2555 444 -2499
rect 534 -2500 535 -2446
rect 723 -2555 724 -2499
rect 810 -2500 811 -2446
rect 1388 -2555 1389 -2499
rect 1542 -2500 1543 -2446
rect 1549 -2555 1550 -2499
rect 198 -2502 199 -2446
rect 219 -2555 220 -2501
rect 275 -2555 276 -2501
rect 733 -2502 734 -2446
rect 884 -2502 885 -2446
rect 919 -2555 920 -2501
rect 933 -2555 934 -2501
rect 1297 -2502 1298 -2446
rect 1325 -2502 1326 -2446
rect 1332 -2555 1333 -2501
rect 1339 -2502 1340 -2446
rect 1654 -2555 1655 -2501
rect 173 -2555 174 -2503
rect 198 -2555 199 -2503
rect 331 -2504 332 -2446
rect 457 -2555 458 -2503
rect 534 -2555 535 -2503
rect 849 -2504 850 -2446
rect 1038 -2504 1039 -2446
rect 1157 -2555 1158 -2503
rect 1178 -2504 1179 -2446
rect 1297 -2555 1298 -2503
rect 1339 -2555 1340 -2503
rect 1580 -2504 1581 -2446
rect 51 -2506 52 -2446
rect 849 -2555 850 -2505
rect 1003 -2506 1004 -2446
rect 1038 -2555 1039 -2505
rect 1052 -2506 1053 -2446
rect 1136 -2555 1137 -2505
rect 1185 -2506 1186 -2446
rect 1381 -2555 1382 -2505
rect 1444 -2506 1445 -2446
rect 1542 -2555 1543 -2505
rect 51 -2555 52 -2507
rect 170 -2508 171 -2446
rect 268 -2508 269 -2446
rect 331 -2555 332 -2507
rect 338 -2508 339 -2446
rect 341 -2520 342 -2507
rect 415 -2555 416 -2507
rect 530 -2508 531 -2446
rect 548 -2508 549 -2446
rect 583 -2555 584 -2507
rect 590 -2555 591 -2507
rect 639 -2555 640 -2507
rect 663 -2555 664 -2507
rect 1178 -2555 1179 -2507
rect 1185 -2555 1186 -2507
rect 1423 -2508 1424 -2446
rect 268 -2555 269 -2509
rect 289 -2510 290 -2446
rect 338 -2555 339 -2509
rect 380 -2510 381 -2446
rect 548 -2555 549 -2509
rect 1115 -2555 1116 -2509
rect 1206 -2510 1207 -2446
rect 1444 -2555 1445 -2509
rect 163 -2555 164 -2511
rect 1206 -2555 1207 -2511
rect 1209 -2512 1210 -2446
rect 1451 -2555 1452 -2511
rect 289 -2555 290 -2513
rect 446 -2555 447 -2513
rect 569 -2555 570 -2513
rect 604 -2514 605 -2446
rect 625 -2514 626 -2446
rect 632 -2555 633 -2513
rect 695 -2514 696 -2446
rect 793 -2555 794 -2513
rect 821 -2555 822 -2513
rect 1423 -2555 1424 -2513
rect 156 -2516 157 -2446
rect 625 -2555 626 -2515
rect 733 -2555 734 -2515
rect 1706 -2555 1707 -2515
rect 156 -2555 157 -2517
rect 747 -2518 748 -2446
rect 835 -2518 836 -2446
rect 884 -2555 885 -2517
rect 926 -2518 927 -2446
rect 1003 -2555 1004 -2517
rect 1010 -2518 1011 -2446
rect 1052 -2555 1053 -2517
rect 1059 -2518 1060 -2446
rect 1073 -2555 1074 -2517
rect 1083 -2555 1084 -2517
rect 1122 -2555 1123 -2517
rect 1213 -2518 1214 -2446
rect 1472 -2555 1473 -2517
rect 380 -2555 381 -2519
rect 555 -2520 556 -2446
rect 695 -2555 696 -2519
rect 709 -2520 710 -2446
rect 835 -2555 836 -2519
rect 926 -2555 927 -2519
rect 982 -2555 983 -2519
rect 1059 -2555 1060 -2519
rect 1150 -2520 1151 -2446
rect 1213 -2555 1214 -2519
rect 1318 -2520 1319 -2446
rect 1360 -2520 1361 -2446
rect 1465 -2555 1466 -2519
rect 576 -2555 577 -2521
rect 737 -2522 738 -2446
rect 863 -2522 864 -2446
rect 1318 -2555 1319 -2521
rect 135 -2524 136 -2446
rect 737 -2555 738 -2523
rect 863 -2555 864 -2523
rect 905 -2524 906 -2446
rect 975 -2524 976 -2446
rect 1010 -2555 1011 -2523
rect 1066 -2524 1067 -2446
rect 1430 -2555 1431 -2523
rect 135 -2555 136 -2525
rect 191 -2526 192 -2446
rect 394 -2526 395 -2446
rect 1066 -2555 1067 -2525
rect 1087 -2526 1088 -2446
rect 1150 -2555 1151 -2525
rect 1220 -2526 1221 -2446
rect 1325 -2555 1326 -2525
rect 114 -2528 115 -2446
rect 191 -2555 192 -2527
rect 394 -2555 395 -2527
rect 667 -2528 668 -2446
rect 705 -2528 706 -2446
rect 905 -2555 906 -2527
rect 1087 -2555 1088 -2527
rect 1633 -2555 1634 -2527
rect 114 -2555 115 -2529
rect 618 -2530 619 -2446
rect 660 -2530 661 -2446
rect 747 -2555 748 -2529
rect 814 -2530 815 -2446
rect 975 -2555 976 -2529
rect 1090 -2555 1091 -2529
rect 1556 -2555 1557 -2529
rect 68 -2555 69 -2531
rect 618 -2555 619 -2531
rect 660 -2555 661 -2531
rect 1374 -2532 1375 -2446
rect 604 -2555 605 -2533
rect 940 -2534 941 -2446
rect 1220 -2555 1221 -2533
rect 1591 -2534 1592 -2446
rect 478 -2536 479 -2446
rect 940 -2555 941 -2535
rect 1248 -2536 1249 -2446
rect 1647 -2555 1648 -2535
rect 205 -2538 206 -2446
rect 478 -2555 479 -2537
rect 667 -2555 668 -2537
rect 901 -2538 902 -2446
rect 1143 -2538 1144 -2446
rect 1248 -2555 1249 -2537
rect 1255 -2555 1256 -2537
rect 1353 -2538 1354 -2446
rect 1374 -2555 1375 -2537
rect 1493 -2538 1494 -2446
rect 1535 -2538 1536 -2446
rect 1591 -2555 1592 -2537
rect 205 -2555 206 -2539
rect 968 -2540 969 -2446
rect 1045 -2540 1046 -2446
rect 1143 -2555 1144 -2539
rect 1234 -2540 1235 -2446
rect 1353 -2555 1354 -2539
rect 1402 -2540 1403 -2446
rect 1493 -2555 1494 -2539
rect 709 -2555 710 -2541
rect 789 -2555 790 -2541
rect 814 -2555 815 -2541
rect 824 -2542 825 -2446
rect 856 -2542 857 -2446
rect 968 -2555 969 -2541
rect 989 -2542 990 -2446
rect 1045 -2555 1046 -2541
rect 1171 -2542 1172 -2446
rect 1234 -2555 1235 -2541
rect 1262 -2542 1263 -2446
rect 1360 -2555 1361 -2541
rect 1437 -2542 1438 -2446
rect 1535 -2555 1536 -2541
rect 555 -2555 556 -2543
rect 824 -2555 825 -2543
rect 856 -2555 857 -2543
rect 954 -2555 955 -2543
rect 989 -2555 990 -2543
rect 1108 -2544 1109 -2446
rect 1164 -2544 1165 -2446
rect 1262 -2555 1263 -2543
rect 1283 -2544 1284 -2446
rect 1402 -2555 1403 -2543
rect 758 -2546 759 -2446
rect 1283 -2555 1284 -2545
rect 730 -2555 731 -2547
rect 758 -2555 759 -2547
rect 1017 -2548 1018 -2446
rect 1108 -2555 1109 -2547
rect 1164 -2555 1165 -2547
rect 1479 -2555 1480 -2547
rect 772 -2550 773 -2446
rect 1017 -2555 1018 -2549
rect 1101 -2550 1102 -2446
rect 1171 -2555 1172 -2549
rect 1195 -2550 1196 -2446
rect 1437 -2555 1438 -2549
rect 646 -2552 647 -2446
rect 772 -2555 773 -2551
rect 1080 -2552 1081 -2446
rect 1101 -2555 1102 -2551
rect 345 -2555 346 -2553
rect 646 -2555 647 -2553
rect 1080 -2555 1081 -2553
rect 1241 -2555 1242 -2553
rect 72 -2565 73 -2563
rect 478 -2565 479 -2563
rect 513 -2565 514 -2563
rect 786 -2565 787 -2563
rect 789 -2565 790 -2563
rect 1430 -2565 1431 -2563
rect 1678 -2565 1679 -2563
rect 1731 -2565 1732 -2563
rect 75 -2567 76 -2563
rect 1563 -2567 1564 -2563
rect 1703 -2567 1704 -2563
rect 1738 -2567 1739 -2563
rect 79 -2569 80 -2563
rect 446 -2569 447 -2563
rect 460 -2684 461 -2568
rect 604 -2569 605 -2563
rect 618 -2569 619 -2563
rect 1185 -2569 1186 -2563
rect 1192 -2569 1193 -2563
rect 1192 -2684 1193 -2568
rect 1192 -2569 1193 -2563
rect 1192 -2684 1193 -2568
rect 1346 -2569 1347 -2563
rect 1346 -2684 1347 -2568
rect 1346 -2569 1347 -2563
rect 1346 -2684 1347 -2568
rect 1430 -2684 1431 -2568
rect 1500 -2569 1501 -2563
rect 1563 -2684 1564 -2568
rect 1626 -2569 1627 -2563
rect 1703 -2684 1704 -2568
rect 1717 -2569 1718 -2563
rect 93 -2571 94 -2563
rect 93 -2684 94 -2570
rect 93 -2571 94 -2563
rect 93 -2684 94 -2570
rect 100 -2571 101 -2563
rect 849 -2571 850 -2563
rect 873 -2571 874 -2563
rect 1241 -2571 1242 -2563
rect 1500 -2684 1501 -2570
rect 1584 -2571 1585 -2563
rect 1626 -2684 1627 -2570
rect 1661 -2571 1662 -2563
rect 100 -2684 101 -2572
rect 135 -2573 136 -2563
rect 149 -2573 150 -2563
rect 1066 -2573 1067 -2563
rect 1080 -2684 1081 -2572
rect 1129 -2573 1130 -2563
rect 1178 -2573 1179 -2563
rect 1185 -2684 1186 -2572
rect 1374 -2573 1375 -2563
rect 1584 -2684 1585 -2572
rect 128 -2575 129 -2563
rect 149 -2684 150 -2574
rect 170 -2575 171 -2563
rect 401 -2575 402 -2563
rect 429 -2575 430 -2563
rect 856 -2575 857 -2563
rect 873 -2684 874 -2574
rect 1262 -2575 1263 -2563
rect 1374 -2684 1375 -2574
rect 1423 -2575 1424 -2563
rect 58 -2577 59 -2563
rect 429 -2684 430 -2576
rect 432 -2577 433 -2563
rect 527 -2577 528 -2563
rect 548 -2577 549 -2563
rect 1458 -2577 1459 -2563
rect 58 -2684 59 -2578
rect 324 -2579 325 -2563
rect 373 -2579 374 -2563
rect 376 -2617 377 -2578
rect 436 -2579 437 -2563
rect 548 -2684 549 -2578
rect 555 -2579 556 -2563
rect 786 -2684 787 -2578
rect 793 -2579 794 -2563
rect 793 -2684 794 -2578
rect 793 -2579 794 -2563
rect 793 -2684 794 -2578
rect 800 -2579 801 -2563
rect 1423 -2684 1424 -2578
rect 1458 -2684 1459 -2578
rect 1689 -2579 1690 -2563
rect 44 -2581 45 -2563
rect 555 -2684 556 -2580
rect 576 -2581 577 -2563
rect 824 -2581 825 -2563
rect 845 -2684 846 -2580
rect 1654 -2581 1655 -2563
rect 44 -2684 45 -2582
rect 89 -2684 90 -2582
rect 121 -2583 122 -2563
rect 170 -2684 171 -2582
rect 201 -2684 202 -2582
rect 1416 -2583 1417 -2563
rect 1542 -2583 1543 -2563
rect 1654 -2684 1655 -2582
rect 128 -2684 129 -2584
rect 394 -2585 395 -2563
rect 436 -2684 437 -2584
rect 478 -2684 479 -2584
rect 506 -2585 507 -2563
rect 849 -2684 850 -2584
rect 856 -2684 857 -2584
rect 891 -2585 892 -2563
rect 898 -2585 899 -2563
rect 898 -2684 899 -2584
rect 898 -2585 899 -2563
rect 898 -2684 899 -2584
rect 926 -2585 927 -2563
rect 1647 -2585 1648 -2563
rect 135 -2684 136 -2586
rect 663 -2587 664 -2563
rect 670 -2684 671 -2586
rect 1682 -2587 1683 -2563
rect 152 -2589 153 -2563
rect 1689 -2684 1690 -2588
rect 240 -2591 241 -2563
rect 576 -2684 577 -2590
rect 593 -2591 594 -2563
rect 611 -2591 612 -2563
rect 625 -2591 626 -2563
rect 1696 -2591 1697 -2563
rect 240 -2684 241 -2592
rect 261 -2593 262 -2563
rect 268 -2593 269 -2563
rect 527 -2684 528 -2592
rect 600 -2684 601 -2592
rect 1143 -2593 1144 -2563
rect 1178 -2684 1179 -2592
rect 1227 -2593 1228 -2563
rect 1262 -2684 1263 -2592
rect 1304 -2593 1305 -2563
rect 1395 -2593 1396 -2563
rect 1661 -2684 1662 -2592
rect 1696 -2684 1697 -2592
rect 1724 -2593 1725 -2563
rect 226 -2595 227 -2563
rect 268 -2684 269 -2594
rect 303 -2595 304 -2563
rect 394 -2684 395 -2594
rect 401 -2684 402 -2594
rect 891 -2684 892 -2594
rect 905 -2595 906 -2563
rect 926 -2684 927 -2594
rect 954 -2595 955 -2563
rect 1451 -2595 1452 -2563
rect 212 -2597 213 -2563
rect 226 -2684 227 -2596
rect 233 -2597 234 -2563
rect 303 -2684 304 -2596
rect 324 -2684 325 -2596
rect 380 -2597 381 -2563
rect 506 -2684 507 -2596
rect 590 -2597 591 -2563
rect 604 -2684 605 -2596
rect 674 -2597 675 -2563
rect 681 -2597 682 -2563
rect 681 -2684 682 -2596
rect 681 -2597 682 -2563
rect 681 -2684 682 -2596
rect 730 -2597 731 -2563
rect 940 -2597 941 -2563
rect 975 -2597 976 -2563
rect 975 -2684 976 -2596
rect 975 -2597 976 -2563
rect 975 -2684 976 -2596
rect 1034 -2684 1035 -2596
rect 1129 -2684 1130 -2596
rect 1213 -2597 1214 -2563
rect 1304 -2684 1305 -2596
rect 1395 -2684 1396 -2596
rect 1437 -2597 1438 -2563
rect 1451 -2684 1452 -2596
rect 1521 -2597 1522 -2563
rect 117 -2684 118 -2598
rect 940 -2684 941 -2598
rect 1038 -2599 1039 -2563
rect 1083 -2599 1084 -2563
rect 1087 -2684 1088 -2598
rect 1283 -2599 1284 -2563
rect 1416 -2684 1417 -2598
rect 1493 -2599 1494 -2563
rect 163 -2601 164 -2563
rect 590 -2684 591 -2600
rect 611 -2684 612 -2600
rect 695 -2601 696 -2563
rect 733 -2601 734 -2563
rect 1682 -2684 1683 -2600
rect 163 -2684 164 -2602
rect 551 -2603 552 -2563
rect 632 -2603 633 -2563
rect 646 -2603 647 -2563
rect 649 -2603 650 -2563
rect 1353 -2603 1354 -2563
rect 1437 -2684 1438 -2602
rect 1514 -2603 1515 -2563
rect 68 -2684 69 -2604
rect 1353 -2684 1354 -2604
rect 1493 -2684 1494 -2604
rect 1549 -2605 1550 -2563
rect 166 -2607 167 -2563
rect 674 -2684 675 -2606
rect 695 -2684 696 -2606
rect 838 -2684 839 -2606
rect 884 -2607 885 -2563
rect 929 -2607 930 -2563
rect 1010 -2607 1011 -2563
rect 1038 -2684 1039 -2606
rect 1052 -2607 1053 -2563
rect 1052 -2684 1053 -2606
rect 1052 -2607 1053 -2563
rect 1052 -2684 1053 -2606
rect 1059 -2607 1060 -2563
rect 1640 -2607 1641 -2563
rect 166 -2684 167 -2608
rect 1570 -2609 1571 -2563
rect 198 -2611 199 -2563
rect 233 -2684 234 -2610
rect 254 -2611 255 -2563
rect 282 -2611 283 -2563
rect 296 -2611 297 -2563
rect 905 -2684 906 -2610
rect 1003 -2611 1004 -2563
rect 1010 -2684 1011 -2610
rect 1059 -2684 1060 -2610
rect 1101 -2611 1102 -2563
rect 1122 -2611 1123 -2563
rect 1167 -2611 1168 -2563
rect 1227 -2684 1228 -2610
rect 1248 -2611 1249 -2563
rect 1276 -2611 1277 -2563
rect 1570 -2684 1571 -2610
rect 65 -2684 66 -2612
rect 1003 -2684 1004 -2612
rect 1066 -2684 1067 -2612
rect 1339 -2613 1340 -2563
rect 1507 -2613 1508 -2563
rect 1640 -2684 1641 -2612
rect 156 -2615 157 -2563
rect 296 -2684 297 -2614
rect 373 -2684 374 -2614
rect 422 -2615 423 -2563
rect 520 -2615 521 -2563
rect 1090 -2615 1091 -2563
rect 1094 -2615 1095 -2563
rect 1241 -2684 1242 -2614
rect 1276 -2684 1277 -2614
rect 1325 -2615 1326 -2563
rect 1507 -2684 1508 -2614
rect 1710 -2615 1711 -2563
rect 156 -2684 157 -2616
rect 345 -2617 346 -2563
rect 422 -2684 423 -2616
rect 520 -2684 521 -2616
rect 562 -2617 563 -2563
rect 632 -2684 633 -2616
rect 716 -2617 717 -2563
rect 733 -2684 734 -2616
rect 758 -2617 759 -2563
rect 772 -2617 773 -2563
rect 954 -2684 955 -2616
rect 957 -2617 958 -2563
rect 1248 -2684 1249 -2616
rect 1283 -2684 1284 -2616
rect 1318 -2617 1319 -2563
rect 1325 -2684 1326 -2616
rect 1381 -2617 1382 -2563
rect 1514 -2684 1515 -2616
rect 1591 -2617 1592 -2563
rect 212 -2684 213 -2618
rect 359 -2619 360 -2563
rect 380 -2684 381 -2618
rect 387 -2619 388 -2563
rect 464 -2619 465 -2563
rect 758 -2684 759 -2618
rect 772 -2684 773 -2618
rect 807 -2619 808 -2563
rect 821 -2619 822 -2563
rect 1220 -2619 1221 -2563
rect 1255 -2619 1256 -2563
rect 1381 -2684 1382 -2618
rect 1549 -2684 1550 -2618
rect 1612 -2619 1613 -2563
rect 191 -2621 192 -2563
rect 359 -2684 360 -2620
rect 492 -2621 493 -2563
rect 562 -2684 563 -2620
rect 639 -2621 640 -2563
rect 691 -2684 692 -2620
rect 716 -2684 717 -2620
rect 1108 -2621 1109 -2563
rect 1122 -2684 1123 -2620
rect 1150 -2621 1151 -2563
rect 1157 -2621 1158 -2563
rect 1220 -2684 1221 -2620
rect 1255 -2684 1256 -2620
rect 1297 -2621 1298 -2563
rect 1318 -2684 1319 -2620
rect 1360 -2621 1361 -2563
rect 1612 -2684 1613 -2620
rect 1633 -2621 1634 -2563
rect 184 -2623 185 -2563
rect 191 -2684 192 -2622
rect 254 -2684 255 -2622
rect 257 -2623 258 -2563
rect 261 -2684 262 -2622
rect 275 -2623 276 -2563
rect 282 -2684 283 -2622
rect 499 -2623 500 -2563
rect 646 -2684 647 -2622
rect 1164 -2623 1165 -2563
rect 1199 -2623 1200 -2563
rect 1339 -2684 1340 -2622
rect 142 -2625 143 -2563
rect 184 -2684 185 -2624
rect 275 -2684 276 -2624
rect 408 -2625 409 -2563
rect 418 -2684 419 -2624
rect 499 -2684 500 -2624
rect 660 -2625 661 -2563
rect 814 -2625 815 -2563
rect 821 -2684 822 -2624
rect 828 -2625 829 -2563
rect 884 -2684 885 -2624
rect 933 -2625 934 -2563
rect 957 -2684 958 -2624
rect 1542 -2684 1543 -2624
rect 107 -2627 108 -2563
rect 408 -2684 409 -2626
rect 457 -2627 458 -2563
rect 492 -2684 493 -2626
rect 569 -2627 570 -2563
rect 828 -2684 829 -2626
rect 894 -2684 895 -2626
rect 1521 -2684 1522 -2626
rect 107 -2684 108 -2628
rect 205 -2629 206 -2563
rect 310 -2629 311 -2563
rect 457 -2684 458 -2628
rect 471 -2629 472 -2563
rect 569 -2684 570 -2628
rect 744 -2684 745 -2628
rect 765 -2629 766 -2563
rect 779 -2629 780 -2563
rect 814 -2684 815 -2628
rect 933 -2684 934 -2628
rect 961 -2629 962 -2563
rect 989 -2629 990 -2563
rect 1164 -2684 1165 -2628
rect 1199 -2684 1200 -2628
rect 1206 -2629 1207 -2563
rect 1269 -2629 1270 -2563
rect 1633 -2684 1634 -2628
rect 72 -2684 73 -2630
rect 765 -2684 766 -2630
rect 803 -2684 804 -2630
rect 989 -2684 990 -2630
rect 1024 -2631 1025 -2563
rect 1108 -2684 1109 -2630
rect 1150 -2684 1151 -2630
rect 1675 -2631 1676 -2563
rect 142 -2684 143 -2632
rect 667 -2633 668 -2563
rect 747 -2633 748 -2563
rect 1647 -2684 1648 -2632
rect 177 -2635 178 -2563
rect 471 -2684 472 -2634
rect 485 -2635 486 -2563
rect 639 -2684 640 -2634
rect 653 -2635 654 -2563
rect 667 -2684 668 -2634
rect 751 -2635 752 -2563
rect 1486 -2635 1487 -2563
rect 1556 -2635 1557 -2563
rect 1675 -2684 1676 -2634
rect 51 -2637 52 -2563
rect 177 -2684 178 -2636
rect 205 -2684 206 -2636
rect 289 -2637 290 -2563
rect 317 -2637 318 -2563
rect 660 -2684 661 -2636
rect 751 -2684 752 -2636
rect 1143 -2684 1144 -2636
rect 1157 -2684 1158 -2636
rect 1171 -2637 1172 -2563
rect 1206 -2684 1207 -2636
rect 1234 -2637 1235 -2563
rect 1269 -2684 1270 -2636
rect 1311 -2637 1312 -2563
rect 1486 -2684 1487 -2636
rect 1668 -2637 1669 -2563
rect 51 -2684 52 -2638
rect 541 -2639 542 -2563
rect 597 -2639 598 -2563
rect 779 -2684 780 -2638
rect 807 -2684 808 -2638
rect 835 -2639 836 -2563
rect 947 -2639 948 -2563
rect 961 -2684 962 -2638
rect 982 -2639 983 -2563
rect 1171 -2684 1172 -2638
rect 1297 -2684 1298 -2638
rect 1402 -2639 1403 -2563
rect 1556 -2684 1557 -2638
rect 1619 -2639 1620 -2563
rect 121 -2684 122 -2640
rect 597 -2684 598 -2640
rect 625 -2684 626 -2640
rect 1619 -2684 1620 -2640
rect 247 -2643 248 -2563
rect 310 -2684 311 -2642
rect 317 -2684 318 -2642
rect 450 -2643 451 -2563
rect 534 -2643 535 -2563
rect 653 -2684 654 -2642
rect 702 -2643 703 -2563
rect 982 -2684 983 -2642
rect 1017 -2643 1018 -2563
rect 1024 -2684 1025 -2642
rect 1062 -2643 1063 -2563
rect 1591 -2684 1592 -2642
rect 86 -2645 87 -2563
rect 702 -2684 703 -2644
rect 737 -2645 738 -2563
rect 1668 -2684 1669 -2644
rect 86 -2684 87 -2646
rect 1577 -2647 1578 -2563
rect 289 -2684 290 -2648
rect 464 -2684 465 -2648
rect 534 -2684 535 -2648
rect 800 -2684 801 -2648
rect 1017 -2684 1018 -2648
rect 1031 -2649 1032 -2563
rect 1094 -2684 1095 -2648
rect 1234 -2684 1235 -2648
rect 1290 -2649 1291 -2563
rect 1402 -2684 1403 -2648
rect 338 -2651 339 -2563
rect 387 -2684 388 -2650
rect 411 -2684 412 -2650
rect 485 -2684 486 -2650
rect 541 -2684 542 -2650
rect 863 -2651 864 -2563
rect 1031 -2684 1032 -2650
rect 1360 -2684 1361 -2650
rect 219 -2653 220 -2563
rect 338 -2684 339 -2652
rect 345 -2684 346 -2652
rect 709 -2653 710 -2563
rect 737 -2684 738 -2652
rect 877 -2653 878 -2563
rect 1097 -2684 1098 -2652
rect 1472 -2653 1473 -2563
rect 82 -2684 83 -2654
rect 219 -2684 220 -2654
rect 450 -2684 451 -2654
rect 1213 -2684 1214 -2654
rect 1290 -2684 1291 -2654
rect 1332 -2655 1333 -2563
rect 1472 -2684 1473 -2654
rect 1535 -2655 1536 -2563
rect 628 -2684 629 -2656
rect 947 -2684 948 -2656
rect 1101 -2684 1102 -2656
rect 1115 -2657 1116 -2563
rect 1311 -2684 1312 -2656
rect 1367 -2657 1368 -2563
rect 1535 -2684 1536 -2656
rect 1605 -2657 1606 -2563
rect 443 -2659 444 -2563
rect 1605 -2684 1606 -2658
rect 331 -2661 332 -2563
rect 443 -2684 444 -2660
rect 709 -2684 710 -2660
rect 723 -2661 724 -2563
rect 754 -2661 755 -2563
rect 1577 -2684 1578 -2660
rect 331 -2684 332 -2662
rect 352 -2663 353 -2563
rect 723 -2684 724 -2662
rect 842 -2663 843 -2563
rect 863 -2684 864 -2662
rect 1045 -2663 1046 -2563
rect 1115 -2684 1116 -2662
rect 1136 -2663 1137 -2563
rect 1332 -2684 1333 -2662
rect 1388 -2663 1389 -2563
rect 114 -2665 115 -2563
rect 352 -2684 353 -2664
rect 366 -2665 367 -2563
rect 1045 -2684 1046 -2664
rect 1073 -2665 1074 -2563
rect 1136 -2684 1137 -2664
rect 1367 -2684 1368 -2664
rect 1409 -2665 1410 -2563
rect 366 -2684 367 -2666
rect 583 -2667 584 -2563
rect 768 -2684 769 -2666
rect 1073 -2684 1074 -2666
rect 1388 -2684 1389 -2666
rect 1465 -2667 1466 -2563
rect 415 -2669 416 -2563
rect 583 -2684 584 -2668
rect 877 -2684 878 -2668
rect 912 -2669 913 -2563
rect 1409 -2684 1410 -2668
rect 1479 -2669 1480 -2563
rect 513 -2684 514 -2670
rect 842 -2684 843 -2670
rect 912 -2684 913 -2670
rect 919 -2671 920 -2563
rect 1465 -2684 1466 -2670
rect 1528 -2671 1529 -2563
rect 740 -2673 741 -2563
rect 1479 -2684 1480 -2672
rect 1528 -2684 1529 -2672
rect 1598 -2673 1599 -2563
rect 919 -2684 920 -2674
rect 968 -2675 969 -2563
rect 1444 -2675 1445 -2563
rect 1598 -2684 1599 -2674
rect 870 -2677 871 -2563
rect 1444 -2684 1445 -2676
rect 688 -2679 689 -2563
rect 870 -2684 871 -2678
rect 968 -2684 969 -2678
rect 996 -2679 997 -2563
rect 618 -2684 619 -2680
rect 688 -2684 689 -2680
rect 677 -2684 678 -2682
rect 996 -2684 997 -2682
rect 37 -2833 38 -2693
rect 569 -2694 570 -2692
rect 579 -2694 580 -2692
rect 793 -2694 794 -2692
rect 803 -2694 804 -2692
rect 1395 -2694 1396 -2692
rect 51 -2696 52 -2692
rect 901 -2833 902 -2695
rect 926 -2696 927 -2692
rect 1097 -2833 1098 -2695
rect 1395 -2833 1396 -2695
rect 1486 -2696 1487 -2692
rect 51 -2833 52 -2697
rect 212 -2698 213 -2692
rect 250 -2698 251 -2692
rect 702 -2698 703 -2692
rect 733 -2698 734 -2692
rect 1066 -2698 1067 -2692
rect 1094 -2698 1095 -2692
rect 1703 -2698 1704 -2692
rect 58 -2700 59 -2692
rect 628 -2700 629 -2692
rect 649 -2833 650 -2699
rect 849 -2700 850 -2692
rect 954 -2700 955 -2692
rect 1241 -2700 1242 -2692
rect 1486 -2833 1487 -2699
rect 1696 -2700 1697 -2692
rect 58 -2833 59 -2701
rect 240 -2702 241 -2692
rect 250 -2833 251 -2701
rect 632 -2702 633 -2692
rect 660 -2702 661 -2692
rect 702 -2833 703 -2701
rect 758 -2702 759 -2692
rect 1048 -2833 1049 -2701
rect 1066 -2833 1067 -2701
rect 1122 -2702 1123 -2692
rect 1241 -2833 1242 -2701
rect 1290 -2702 1291 -2692
rect 65 -2704 66 -2692
rect 653 -2704 654 -2692
rect 660 -2833 661 -2703
rect 670 -2704 671 -2692
rect 674 -2704 675 -2692
rect 1297 -2704 1298 -2692
rect 65 -2833 66 -2705
rect 887 -2833 888 -2705
rect 954 -2833 955 -2705
rect 1101 -2706 1102 -2692
rect 1290 -2833 1291 -2705
rect 1430 -2706 1431 -2692
rect 68 -2708 69 -2692
rect 1045 -2708 1046 -2692
rect 1094 -2833 1095 -2707
rect 1668 -2708 1669 -2692
rect 72 -2710 73 -2692
rect 418 -2710 419 -2692
rect 453 -2710 454 -2692
rect 520 -2710 521 -2692
rect 523 -2833 524 -2709
rect 1185 -2710 1186 -2692
rect 1297 -2833 1298 -2709
rect 1416 -2710 1417 -2692
rect 1430 -2833 1431 -2709
rect 1556 -2710 1557 -2692
rect 82 -2712 83 -2692
rect 786 -2712 787 -2692
rect 793 -2833 794 -2711
rect 947 -2712 948 -2692
rect 957 -2712 958 -2692
rect 1549 -2712 1550 -2692
rect 1556 -2833 1557 -2711
rect 1577 -2712 1578 -2692
rect 110 -2833 111 -2713
rect 1283 -2714 1284 -2692
rect 1416 -2833 1417 -2713
rect 1619 -2714 1620 -2692
rect 114 -2716 115 -2692
rect 555 -2716 556 -2692
rect 583 -2716 584 -2692
rect 1510 -2833 1511 -2715
rect 1549 -2833 1550 -2715
rect 1598 -2716 1599 -2692
rect 114 -2833 115 -2717
rect 639 -2718 640 -2692
rect 653 -2833 654 -2717
rect 1122 -2833 1123 -2717
rect 1283 -2833 1284 -2717
rect 1423 -2718 1424 -2692
rect 117 -2720 118 -2692
rect 618 -2720 619 -2692
rect 625 -2720 626 -2692
rect 884 -2720 885 -2692
rect 947 -2833 948 -2719
rect 1150 -2720 1151 -2692
rect 1423 -2833 1424 -2719
rect 1626 -2720 1627 -2692
rect 121 -2722 122 -2692
rect 800 -2722 801 -2692
rect 814 -2722 815 -2692
rect 845 -2722 846 -2692
rect 849 -2833 850 -2721
rect 1003 -2722 1004 -2692
rect 1034 -2722 1035 -2692
rect 1381 -2722 1382 -2692
rect 121 -2833 122 -2723
rect 247 -2724 248 -2692
rect 275 -2724 276 -2692
rect 278 -2724 279 -2692
rect 289 -2724 290 -2692
rect 478 -2833 479 -2723
rect 481 -2724 482 -2692
rect 562 -2724 563 -2692
rect 583 -2833 584 -2723
rect 982 -2724 983 -2692
rect 989 -2724 990 -2692
rect 1654 -2724 1655 -2692
rect 107 -2726 108 -2692
rect 289 -2833 290 -2725
rect 331 -2726 332 -2692
rect 775 -2833 776 -2725
rect 786 -2833 787 -2725
rect 940 -2726 941 -2692
rect 989 -2833 990 -2725
rect 1227 -2726 1228 -2692
rect 1381 -2833 1382 -2725
rect 1612 -2726 1613 -2692
rect 86 -2728 87 -2692
rect 107 -2833 108 -2727
rect 128 -2728 129 -2692
rect 754 -2728 755 -2692
rect 758 -2833 759 -2727
rect 933 -2728 934 -2692
rect 940 -2833 941 -2727
rect 1129 -2728 1130 -2692
rect 1150 -2833 1151 -2727
rect 1276 -2728 1277 -2692
rect 86 -2833 87 -2729
rect 1675 -2730 1676 -2692
rect 93 -2732 94 -2692
rect 128 -2833 129 -2731
rect 142 -2732 143 -2692
rect 677 -2732 678 -2692
rect 688 -2732 689 -2692
rect 1199 -2732 1200 -2692
rect 1227 -2833 1228 -2731
rect 1409 -2732 1410 -2692
rect 72 -2833 73 -2733
rect 93 -2833 94 -2733
rect 149 -2734 150 -2692
rect 152 -2772 153 -2733
rect 166 -2734 167 -2692
rect 331 -2833 332 -2733
rect 352 -2734 353 -2692
rect 639 -2833 640 -2733
rect 667 -2734 668 -2692
rect 681 -2734 682 -2692
rect 765 -2734 766 -2692
rect 1192 -2734 1193 -2692
rect 1199 -2833 1200 -2733
rect 1325 -2734 1326 -2692
rect 89 -2736 90 -2692
rect 142 -2833 143 -2735
rect 149 -2833 150 -2735
rect 198 -2736 199 -2692
rect 201 -2736 202 -2692
rect 730 -2736 731 -2692
rect 814 -2833 815 -2735
rect 863 -2736 864 -2692
rect 873 -2736 874 -2692
rect 1129 -2833 1130 -2735
rect 1192 -2833 1193 -2735
rect 1339 -2736 1340 -2692
rect 89 -2833 90 -2737
rect 338 -2738 339 -2692
rect 373 -2738 374 -2692
rect 415 -2738 416 -2692
rect 429 -2738 430 -2692
rect 800 -2833 801 -2737
rect 835 -2738 836 -2692
rect 898 -2738 899 -2692
rect 933 -2833 934 -2737
rect 1073 -2738 1074 -2692
rect 1101 -2833 1102 -2737
rect 1311 -2738 1312 -2692
rect 1325 -2833 1326 -2737
rect 1500 -2738 1501 -2692
rect 166 -2833 167 -2739
rect 576 -2833 577 -2739
rect 593 -2833 594 -2739
rect 1185 -2833 1186 -2739
rect 1311 -2833 1312 -2739
rect 1605 -2740 1606 -2692
rect 180 -2833 181 -2741
rect 1633 -2742 1634 -2692
rect 184 -2744 185 -2692
rect 198 -2833 199 -2743
rect 205 -2744 206 -2692
rect 338 -2833 339 -2743
rect 359 -2744 360 -2692
rect 373 -2833 374 -2743
rect 380 -2744 381 -2692
rect 380 -2833 381 -2743
rect 380 -2744 381 -2692
rect 380 -2833 381 -2743
rect 387 -2744 388 -2692
rect 387 -2833 388 -2743
rect 387 -2744 388 -2692
rect 387 -2833 388 -2743
rect 401 -2744 402 -2692
rect 569 -2833 570 -2743
rect 597 -2744 598 -2692
rect 1689 -2744 1690 -2692
rect 156 -2746 157 -2692
rect 205 -2833 206 -2745
rect 212 -2833 213 -2745
rect 226 -2746 227 -2692
rect 240 -2833 241 -2745
rect 261 -2746 262 -2692
rect 268 -2746 269 -2692
rect 352 -2833 353 -2745
rect 359 -2833 360 -2745
rect 485 -2746 486 -2692
rect 506 -2746 507 -2692
rect 632 -2833 633 -2745
rect 667 -2833 668 -2745
rect 1017 -2746 1018 -2692
rect 1045 -2833 1046 -2745
rect 1584 -2746 1585 -2692
rect 44 -2748 45 -2692
rect 226 -2833 227 -2747
rect 254 -2748 255 -2692
rect 261 -2833 262 -2747
rect 268 -2833 269 -2747
rect 467 -2748 468 -2692
rect 485 -2833 486 -2747
rect 723 -2748 724 -2692
rect 730 -2833 731 -2747
rect 856 -2748 857 -2692
rect 863 -2833 864 -2747
rect 1188 -2833 1189 -2747
rect 1339 -2833 1340 -2747
rect 1542 -2748 1543 -2692
rect 44 -2833 45 -2749
rect 100 -2750 101 -2692
rect 131 -2833 132 -2749
rect 723 -2833 724 -2749
rect 835 -2833 836 -2749
rect 996 -2750 997 -2692
rect 1003 -2833 1004 -2749
rect 1136 -2750 1137 -2692
rect 1374 -2750 1375 -2692
rect 1542 -2833 1543 -2749
rect 96 -2833 97 -2751
rect 156 -2833 157 -2751
rect 184 -2833 185 -2751
rect 254 -2833 255 -2751
rect 383 -2833 384 -2751
rect 401 -2833 402 -2751
rect 436 -2752 437 -2692
rect 450 -2752 451 -2692
rect 982 -2833 983 -2751
rect 1017 -2833 1018 -2751
rect 1171 -2752 1172 -2692
rect 1374 -2833 1375 -2751
rect 1437 -2752 1438 -2692
rect 1458 -2752 1459 -2692
rect 1500 -2833 1501 -2751
rect 100 -2833 101 -2753
rect 282 -2754 283 -2692
rect 345 -2754 346 -2692
rect 996 -2833 997 -2753
rect 1073 -2833 1074 -2753
rect 1255 -2754 1256 -2692
rect 1437 -2833 1438 -2753
rect 1563 -2754 1564 -2692
rect 275 -2833 276 -2755
rect 324 -2756 325 -2692
rect 345 -2833 346 -2755
rect 492 -2756 493 -2692
rect 520 -2833 521 -2755
rect 688 -2833 689 -2755
rect 716 -2756 717 -2692
rect 856 -2833 857 -2755
rect 884 -2833 885 -2755
rect 1255 -2833 1256 -2755
rect 1458 -2833 1459 -2755
rect 1661 -2756 1662 -2692
rect 233 -2758 234 -2692
rect 492 -2833 493 -2757
rect 534 -2758 535 -2692
rect 1031 -2758 1032 -2692
rect 1136 -2833 1137 -2757
rect 1269 -2758 1270 -2692
rect 177 -2760 178 -2692
rect 233 -2833 234 -2759
rect 282 -2833 283 -2759
rect 450 -2833 451 -2759
rect 457 -2760 458 -2692
rect 1409 -2833 1410 -2759
rect 229 -2833 230 -2761
rect 457 -2833 458 -2761
rect 534 -2833 535 -2761
rect 975 -2762 976 -2692
rect 1031 -2833 1032 -2761
rect 1087 -2762 1088 -2692
rect 1171 -2833 1172 -2761
rect 1360 -2762 1361 -2692
rect 317 -2764 318 -2692
rect 324 -2833 325 -2763
rect 366 -2764 367 -2692
rect 506 -2833 507 -2763
rect 541 -2764 542 -2692
rect 894 -2764 895 -2692
rect 898 -2833 899 -2763
rect 926 -2833 927 -2763
rect 975 -2833 976 -2763
rect 1052 -2764 1053 -2692
rect 1269 -2833 1270 -2763
rect 1451 -2764 1452 -2692
rect 296 -2766 297 -2692
rect 366 -2833 367 -2765
rect 408 -2833 409 -2765
rect 1279 -2833 1280 -2765
rect 1360 -2833 1361 -2765
rect 1591 -2766 1592 -2692
rect 296 -2833 297 -2767
rect 422 -2768 423 -2692
rect 429 -2833 430 -2767
rect 611 -2768 612 -2692
rect 618 -2833 619 -2767
rect 1108 -2768 1109 -2692
rect 1451 -2833 1452 -2767
rect 1640 -2768 1641 -2692
rect 317 -2833 318 -2769
rect 443 -2770 444 -2692
rect 499 -2770 500 -2692
rect 611 -2833 612 -2769
rect 625 -2833 626 -2769
rect 709 -2770 710 -2692
rect 716 -2833 717 -2769
rect 751 -2770 752 -2692
rect 870 -2770 871 -2692
rect 1087 -2833 1088 -2769
rect 1108 -2833 1109 -2769
rect 1262 -2770 1263 -2692
rect 278 -2833 279 -2771
rect 443 -2833 444 -2771
rect 499 -2833 500 -2771
rect 744 -2772 745 -2692
rect 751 -2833 752 -2771
rect 772 -2772 773 -2692
rect 870 -2833 871 -2771
rect 1164 -2772 1165 -2692
rect 1262 -2833 1263 -2771
rect 1472 -2772 1473 -2692
rect 411 -2774 412 -2692
rect 527 -2774 528 -2692
rect 541 -2833 542 -2773
rect 590 -2774 591 -2692
rect 597 -2833 598 -2773
rect 919 -2774 920 -2692
rect 1052 -2833 1053 -2773
rect 1332 -2774 1333 -2692
rect 1472 -2833 1473 -2773
rect 1507 -2774 1508 -2692
rect 415 -2833 416 -2775
rect 684 -2833 685 -2775
rect 709 -2833 710 -2775
rect 877 -2776 878 -2692
rect 894 -2833 895 -2775
rect 1682 -2776 1683 -2692
rect 247 -2833 248 -2777
rect 877 -2833 878 -2777
rect 919 -2833 920 -2777
rect 1213 -2778 1214 -2692
rect 1332 -2833 1333 -2777
rect 1535 -2778 1536 -2692
rect 422 -2833 423 -2779
rect 803 -2833 804 -2779
rect 1164 -2833 1165 -2779
rect 1367 -2780 1368 -2692
rect 1493 -2780 1494 -2692
rect 1507 -2833 1508 -2779
rect 436 -2833 437 -2781
rect 548 -2782 549 -2692
rect 555 -2833 556 -2781
rect 807 -2782 808 -2692
rect 1213 -2833 1214 -2781
rect 1444 -2782 1445 -2692
rect 1493 -2833 1494 -2781
rect 1647 -2782 1648 -2692
rect 219 -2784 220 -2692
rect 548 -2833 549 -2783
rect 562 -2833 563 -2783
rect 779 -2784 780 -2692
rect 807 -2833 808 -2783
rect 961 -2784 962 -2692
rect 1248 -2784 1249 -2692
rect 1444 -2833 1445 -2783
rect 170 -2786 171 -2692
rect 219 -2833 220 -2785
rect 527 -2833 528 -2785
rect 985 -2833 986 -2785
rect 1206 -2786 1207 -2692
rect 1248 -2833 1249 -2785
rect 1346 -2786 1347 -2692
rect 1535 -2833 1536 -2785
rect 170 -2833 171 -2787
rect 768 -2788 769 -2692
rect 842 -2788 843 -2692
rect 1206 -2833 1207 -2787
rect 1346 -2833 1347 -2787
rect 1514 -2788 1515 -2692
rect 79 -2790 80 -2692
rect 1514 -2833 1515 -2789
rect 79 -2833 80 -2791
rect 394 -2792 395 -2692
rect 590 -2833 591 -2791
rect 821 -2792 822 -2692
rect 842 -2833 843 -2791
rect 912 -2792 913 -2692
rect 961 -2833 962 -2791
rect 1115 -2792 1116 -2692
rect 1367 -2833 1368 -2791
rect 1388 -2792 1389 -2692
rect 394 -2833 395 -2793
rect 471 -2794 472 -2692
rect 600 -2794 601 -2692
rect 737 -2794 738 -2692
rect 744 -2833 745 -2793
rect 828 -2794 829 -2692
rect 912 -2833 913 -2793
rect 968 -2794 969 -2692
rect 1115 -2833 1116 -2793
rect 1388 -2833 1389 -2793
rect 135 -2796 136 -2692
rect 471 -2833 472 -2795
rect 674 -2833 675 -2795
rect 1080 -2796 1081 -2692
rect 135 -2833 136 -2797
rect 646 -2798 647 -2692
rect 681 -2833 682 -2797
rect 1318 -2798 1319 -2692
rect 464 -2800 465 -2692
rect 737 -2833 738 -2799
rect 761 -2833 762 -2799
rect 779 -2833 780 -2799
rect 821 -2833 822 -2799
rect 1010 -2800 1011 -2692
rect 1318 -2833 1319 -2799
rect 1479 -2800 1480 -2692
rect 163 -2802 164 -2692
rect 1479 -2833 1480 -2801
rect 163 -2833 164 -2803
rect 905 -2804 906 -2692
rect 999 -2833 1000 -2803
rect 1080 -2833 1081 -2803
rect 310 -2806 311 -2692
rect 464 -2833 465 -2805
rect 765 -2833 766 -2805
rect 968 -2833 969 -2805
rect 303 -2808 304 -2692
rect 310 -2833 311 -2807
rect 768 -2833 769 -2807
rect 1024 -2808 1025 -2692
rect 303 -2833 304 -2809
rect 513 -2810 514 -2692
rect 772 -2833 773 -2809
rect 828 -2833 829 -2809
rect 838 -2810 839 -2692
rect 905 -2833 906 -2809
rect 1024 -2833 1025 -2809
rect 1157 -2810 1158 -2692
rect 513 -2833 514 -2811
rect 604 -2812 605 -2692
rect 891 -2833 892 -2811
rect 1010 -2833 1011 -2811
rect 1157 -2833 1158 -2811
rect 1178 -2812 1179 -2692
rect 604 -2833 605 -2813
rect 695 -2814 696 -2692
rect 1178 -2833 1179 -2813
rect 1220 -2814 1221 -2692
rect 695 -2833 696 -2815
rect 1038 -2816 1039 -2692
rect 1220 -2833 1221 -2815
rect 1465 -2816 1466 -2692
rect 1038 -2833 1039 -2817
rect 1059 -2818 1060 -2692
rect 1465 -2833 1466 -2817
rect 1521 -2818 1522 -2692
rect 1059 -2833 1060 -2819
rect 1353 -2820 1354 -2692
rect 1304 -2822 1305 -2692
rect 1521 -2833 1522 -2821
rect 1234 -2824 1235 -2692
rect 1304 -2833 1305 -2823
rect 1353 -2833 1354 -2823
rect 1570 -2824 1571 -2692
rect 1234 -2833 1235 -2825
rect 1402 -2826 1403 -2692
rect 1402 -2833 1403 -2827
rect 1528 -2828 1529 -2692
rect 1143 -2830 1144 -2692
rect 1528 -2833 1529 -2829
rect 1143 -2833 1144 -2831
rect 1276 -2833 1277 -2831
rect 30 -2944 31 -2842
rect 457 -2843 458 -2841
rect 506 -2843 507 -2841
rect 656 -2843 657 -2841
rect 765 -2843 766 -2841
rect 842 -2843 843 -2841
rect 887 -2843 888 -2841
rect 929 -2944 930 -2842
rect 982 -2843 983 -2841
rect 1402 -2843 1403 -2841
rect 1514 -2843 1515 -2841
rect 1556 -2843 1557 -2841
rect 37 -2845 38 -2841
rect 502 -2944 503 -2844
rect 583 -2845 584 -2841
rect 653 -2845 654 -2841
rect 702 -2845 703 -2841
rect 842 -2944 843 -2844
rect 898 -2845 899 -2841
rect 1374 -2845 1375 -2841
rect 1395 -2845 1396 -2841
rect 1402 -2944 1403 -2844
rect 37 -2944 38 -2846
rect 499 -2847 500 -2841
rect 569 -2847 570 -2841
rect 583 -2944 584 -2846
rect 593 -2847 594 -2841
rect 793 -2847 794 -2841
rect 803 -2847 804 -2841
rect 961 -2847 962 -2841
rect 996 -2847 997 -2841
rect 1192 -2847 1193 -2841
rect 1202 -2944 1203 -2846
rect 1367 -2847 1368 -2841
rect 44 -2849 45 -2841
rect 117 -2944 118 -2848
rect 121 -2849 122 -2841
rect 565 -2944 566 -2848
rect 607 -2944 608 -2848
rect 681 -2944 682 -2848
rect 751 -2849 752 -2841
rect 765 -2944 766 -2848
rect 775 -2849 776 -2841
rect 1199 -2849 1200 -2841
rect 1276 -2944 1277 -2848
rect 1332 -2849 1333 -2841
rect 1367 -2944 1368 -2848
rect 1388 -2849 1389 -2841
rect 51 -2851 52 -2841
rect 226 -2851 227 -2841
rect 250 -2851 251 -2841
rect 1374 -2944 1375 -2850
rect 1388 -2944 1389 -2850
rect 1444 -2851 1445 -2841
rect 51 -2944 52 -2852
rect 625 -2853 626 -2841
rect 653 -2944 654 -2852
rect 828 -2853 829 -2841
rect 877 -2853 878 -2841
rect 1395 -2944 1396 -2852
rect 72 -2855 73 -2841
rect 1115 -2855 1116 -2841
rect 1118 -2855 1119 -2841
rect 1500 -2855 1501 -2841
rect 75 -2944 76 -2856
rect 527 -2857 528 -2841
rect 618 -2857 619 -2841
rect 884 -2857 885 -2841
rect 898 -2944 899 -2856
rect 1507 -2857 1508 -2841
rect 86 -2944 87 -2858
rect 303 -2859 304 -2841
rect 345 -2859 346 -2841
rect 684 -2859 685 -2841
rect 751 -2944 752 -2858
rect 786 -2859 787 -2841
rect 807 -2859 808 -2841
rect 915 -2944 916 -2858
rect 947 -2859 948 -2841
rect 982 -2944 983 -2858
rect 996 -2944 997 -2858
rect 1066 -2859 1067 -2841
rect 1097 -2859 1098 -2841
rect 1437 -2859 1438 -2841
rect 1500 -2944 1501 -2858
rect 1549 -2859 1550 -2841
rect 93 -2861 94 -2841
rect 107 -2861 108 -2841
rect 121 -2944 122 -2860
rect 264 -2944 265 -2860
rect 268 -2861 269 -2841
rect 758 -2861 759 -2841
rect 821 -2861 822 -2841
rect 821 -2944 822 -2860
rect 821 -2861 822 -2841
rect 821 -2944 822 -2860
rect 828 -2944 829 -2860
rect 1031 -2861 1032 -2841
rect 1038 -2861 1039 -2841
rect 1094 -2944 1095 -2860
rect 1164 -2861 1165 -2841
rect 1185 -2861 1186 -2841
rect 1188 -2861 1189 -2841
rect 1430 -2861 1431 -2841
rect 93 -2944 94 -2862
rect 604 -2863 605 -2841
rect 618 -2944 619 -2862
rect 716 -2863 717 -2841
rect 779 -2863 780 -2841
rect 1038 -2944 1039 -2862
rect 1048 -2863 1049 -2841
rect 1136 -2863 1137 -2841
rect 1185 -2944 1186 -2862
rect 1206 -2863 1207 -2841
rect 1279 -2863 1280 -2841
rect 1451 -2863 1452 -2841
rect 96 -2865 97 -2841
rect 534 -2865 535 -2841
rect 625 -2944 626 -2864
rect 688 -2865 689 -2841
rect 695 -2865 696 -2841
rect 807 -2944 808 -2864
rect 856 -2865 857 -2841
rect 877 -2944 878 -2864
rect 905 -2865 906 -2841
rect 1066 -2944 1067 -2864
rect 1192 -2944 1193 -2864
rect 1213 -2865 1214 -2841
rect 1248 -2865 1249 -2841
rect 1451 -2944 1452 -2864
rect 100 -2867 101 -2841
rect 177 -2867 178 -2841
rect 226 -2944 227 -2866
rect 261 -2867 262 -2841
rect 268 -2944 269 -2866
rect 394 -2867 395 -2841
rect 411 -2944 412 -2866
rect 1206 -2944 1207 -2866
rect 1213 -2944 1214 -2866
rect 1283 -2867 1284 -2841
rect 1318 -2867 1319 -2841
rect 1332 -2944 1333 -2866
rect 1430 -2944 1431 -2866
rect 1458 -2867 1459 -2841
rect 100 -2944 101 -2868
rect 229 -2869 230 -2841
rect 275 -2869 276 -2841
rect 303 -2944 304 -2868
rect 345 -2944 346 -2868
rect 387 -2869 388 -2841
rect 429 -2869 430 -2841
rect 569 -2944 570 -2868
rect 576 -2869 577 -2841
rect 695 -2944 696 -2868
rect 709 -2869 710 -2841
rect 786 -2944 787 -2868
rect 800 -2869 801 -2841
rect 1164 -2944 1165 -2868
rect 1283 -2944 1284 -2868
rect 1510 -2869 1511 -2841
rect 107 -2944 108 -2870
rect 541 -2871 542 -2841
rect 646 -2871 647 -2841
rect 1437 -2944 1438 -2870
rect 1458 -2944 1459 -2870
rect 1535 -2871 1536 -2841
rect 128 -2873 129 -2841
rect 793 -2944 794 -2872
rect 800 -2944 801 -2872
rect 849 -2873 850 -2841
rect 866 -2944 867 -2872
rect 884 -2944 885 -2872
rect 905 -2944 906 -2872
rect 933 -2873 934 -2841
rect 940 -2873 941 -2841
rect 1031 -2944 1032 -2872
rect 1129 -2873 1130 -2841
rect 1248 -2944 1249 -2872
rect 1311 -2873 1312 -2841
rect 1318 -2944 1319 -2872
rect 128 -2944 129 -2874
rect 240 -2875 241 -2841
rect 275 -2944 276 -2874
rect 310 -2875 311 -2841
rect 359 -2875 360 -2841
rect 387 -2944 388 -2874
rect 450 -2875 451 -2841
rect 1409 -2875 1410 -2841
rect 135 -2877 136 -2841
rect 534 -2944 535 -2876
rect 541 -2944 542 -2876
rect 639 -2877 640 -2841
rect 646 -2944 647 -2876
rect 989 -2877 990 -2841
rect 1003 -2877 1004 -2841
rect 1136 -2944 1137 -2876
rect 1311 -2944 1312 -2876
rect 1360 -2877 1361 -2841
rect 1409 -2944 1410 -2876
rect 1423 -2877 1424 -2841
rect 135 -2944 136 -2878
rect 180 -2879 181 -2841
rect 191 -2879 192 -2841
rect 310 -2944 311 -2878
rect 331 -2879 332 -2841
rect 450 -2944 451 -2878
rect 457 -2944 458 -2878
rect 590 -2879 591 -2841
rect 660 -2879 661 -2841
rect 709 -2944 710 -2878
rect 716 -2944 717 -2878
rect 768 -2879 769 -2841
rect 779 -2944 780 -2878
rect 863 -2879 864 -2841
rect 912 -2879 913 -2841
rect 1045 -2879 1046 -2841
rect 1080 -2879 1081 -2841
rect 1129 -2944 1130 -2878
rect 1360 -2944 1361 -2878
rect 1381 -2879 1382 -2841
rect 1423 -2944 1424 -2878
rect 1486 -2879 1487 -2841
rect 142 -2881 143 -2841
rect 772 -2944 773 -2880
rect 863 -2944 864 -2880
rect 1150 -2881 1151 -2841
rect 1381 -2944 1382 -2880
rect 1416 -2881 1417 -2841
rect 1486 -2944 1487 -2880
rect 1521 -2881 1522 -2841
rect 142 -2944 143 -2882
rect 212 -2883 213 -2841
rect 219 -2883 220 -2841
rect 394 -2944 395 -2882
rect 474 -2944 475 -2882
rect 1115 -2944 1116 -2882
rect 1150 -2944 1151 -2882
rect 1227 -2883 1228 -2841
rect 1416 -2944 1417 -2882
rect 1447 -2944 1448 -2882
rect 72 -2944 73 -2884
rect 212 -2944 213 -2884
rect 219 -2944 220 -2884
rect 999 -2885 1000 -2841
rect 1003 -2944 1004 -2884
rect 1073 -2885 1074 -2841
rect 1080 -2944 1081 -2884
rect 1241 -2885 1242 -2841
rect 170 -2887 171 -2841
rect 499 -2944 500 -2886
rect 523 -2887 524 -2841
rect 940 -2944 941 -2886
rect 961 -2944 962 -2886
rect 975 -2887 976 -2841
rect 1010 -2887 1011 -2841
rect 1045 -2944 1046 -2886
rect 1122 -2887 1123 -2841
rect 1227 -2944 1228 -2886
rect 1241 -2944 1242 -2886
rect 1262 -2887 1263 -2841
rect 170 -2944 171 -2888
rect 1199 -2944 1200 -2888
rect 177 -2944 178 -2890
rect 240 -2944 241 -2890
rect 282 -2891 283 -2841
rect 576 -2944 577 -2890
rect 660 -2944 661 -2890
rect 744 -2891 745 -2841
rect 870 -2891 871 -2841
rect 1073 -2944 1074 -2890
rect 1087 -2891 1088 -2841
rect 1262 -2944 1263 -2890
rect 163 -2893 164 -2841
rect 282 -2944 283 -2892
rect 331 -2944 332 -2892
rect 366 -2893 367 -2841
rect 373 -2893 374 -2841
rect 520 -2893 521 -2841
rect 527 -2944 528 -2892
rect 548 -2893 549 -2841
rect 555 -2893 556 -2841
rect 639 -2944 640 -2892
rect 667 -2893 668 -2841
rect 849 -2944 850 -2892
rect 912 -2944 913 -2892
rect 1493 -2893 1494 -2841
rect 114 -2895 115 -2841
rect 520 -2944 521 -2894
rect 548 -2944 549 -2894
rect 611 -2895 612 -2841
rect 667 -2944 668 -2894
rect 744 -2944 745 -2894
rect 926 -2895 927 -2841
rect 989 -2944 990 -2894
rect 1010 -2944 1011 -2894
rect 1178 -2895 1179 -2841
rect 1493 -2944 1494 -2894
rect 1528 -2895 1529 -2841
rect 163 -2944 164 -2896
rect 247 -2944 248 -2896
rect 250 -2944 251 -2896
rect 870 -2944 871 -2896
rect 926 -2944 927 -2896
rect 1304 -2897 1305 -2841
rect 191 -2944 192 -2898
rect 205 -2899 206 -2841
rect 359 -2944 360 -2898
rect 936 -2944 937 -2898
rect 975 -2944 976 -2898
rect 1157 -2899 1158 -2841
rect 1178 -2944 1179 -2898
rect 1290 -2899 1291 -2841
rect 1304 -2944 1305 -2898
rect 1353 -2899 1354 -2841
rect 205 -2944 206 -2900
rect 254 -2901 255 -2841
rect 366 -2944 367 -2900
rect 649 -2901 650 -2841
rect 674 -2901 675 -2841
rect 702 -2944 703 -2900
rect 737 -2901 738 -2841
rect 856 -2944 857 -2900
rect 968 -2901 969 -2841
rect 1353 -2944 1354 -2900
rect 254 -2944 255 -2902
rect 338 -2903 339 -2841
rect 380 -2903 381 -2841
rect 429 -2944 430 -2902
rect 485 -2903 486 -2841
rect 590 -2944 591 -2902
rect 597 -2903 598 -2841
rect 674 -2944 675 -2902
rect 761 -2903 762 -2841
rect 968 -2944 969 -2902
rect 1027 -2944 1028 -2902
rect 1479 -2903 1480 -2841
rect 289 -2905 290 -2841
rect 338 -2944 339 -2904
rect 380 -2944 381 -2904
rect 478 -2905 479 -2841
rect 485 -2944 486 -2904
rect 562 -2905 563 -2841
rect 611 -2944 612 -2904
rect 814 -2905 815 -2841
rect 1052 -2905 1053 -2841
rect 1122 -2944 1123 -2904
rect 1157 -2944 1158 -2904
rect 1339 -2905 1340 -2841
rect 1479 -2944 1480 -2904
rect 1542 -2905 1543 -2841
rect 44 -2944 45 -2906
rect 562 -2944 563 -2906
rect 761 -2944 762 -2906
rect 947 -2944 948 -2906
rect 1052 -2944 1053 -2906
rect 1101 -2907 1102 -2841
rect 1255 -2907 1256 -2841
rect 1339 -2944 1340 -2906
rect 65 -2909 66 -2841
rect 289 -2944 290 -2908
rect 408 -2909 409 -2841
rect 737 -2944 738 -2908
rect 814 -2944 815 -2908
rect 835 -2909 836 -2841
rect 1059 -2909 1060 -2841
rect 1087 -2944 1088 -2908
rect 1101 -2944 1102 -2908
rect 1143 -2909 1144 -2841
rect 1255 -2944 1256 -2908
rect 1297 -2909 1298 -2841
rect 65 -2944 66 -2910
rect 415 -2911 416 -2841
rect 436 -2911 437 -2841
rect 597 -2944 598 -2910
rect 733 -2944 734 -2910
rect 1297 -2944 1298 -2910
rect 110 -2913 111 -2841
rect 835 -2944 836 -2912
rect 1059 -2944 1060 -2912
rect 1108 -2913 1109 -2841
rect 1143 -2944 1144 -2912
rect 1171 -2913 1172 -2841
rect 1290 -2944 1291 -2912
rect 1346 -2913 1347 -2841
rect 401 -2915 402 -2841
rect 415 -2944 416 -2914
rect 436 -2944 437 -2914
rect 492 -2915 493 -2841
rect 555 -2944 556 -2914
rect 919 -2915 920 -2841
rect 1171 -2944 1172 -2914
rect 1234 -2915 1235 -2841
rect 58 -2917 59 -2841
rect 401 -2944 402 -2916
rect 408 -2944 409 -2916
rect 464 -2917 465 -2841
rect 478 -2944 479 -2916
rect 901 -2917 902 -2841
rect 919 -2944 920 -2916
rect 954 -2917 955 -2841
rect 1220 -2917 1221 -2841
rect 1234 -2944 1235 -2916
rect 58 -2944 59 -2918
rect 632 -2919 633 -2841
rect 723 -2919 724 -2841
rect 1108 -2944 1109 -2918
rect 1220 -2944 1221 -2918
rect 1269 -2919 1270 -2841
rect 114 -2944 115 -2920
rect 632 -2944 633 -2920
rect 723 -2944 724 -2920
rect 730 -2921 731 -2841
rect 891 -2921 892 -2841
rect 1346 -2944 1347 -2920
rect 149 -2923 150 -2841
rect 891 -2944 892 -2922
rect 954 -2944 955 -2922
rect 1017 -2923 1018 -2841
rect 1269 -2944 1270 -2922
rect 1325 -2923 1326 -2841
rect 149 -2944 150 -2924
rect 184 -2925 185 -2841
rect 317 -2925 318 -2841
rect 464 -2944 465 -2924
rect 471 -2925 472 -2841
rect 730 -2944 731 -2924
rect 1017 -2944 1018 -2924
rect 1024 -2925 1025 -2841
rect 184 -2944 185 -2926
rect 198 -2927 199 -2841
rect 257 -2944 258 -2926
rect 317 -2944 318 -2926
rect 404 -2944 405 -2926
rect 1325 -2944 1326 -2926
rect 198 -2944 199 -2928
rect 296 -2929 297 -2841
rect 422 -2929 423 -2841
rect 492 -2944 493 -2928
rect 1024 -2944 1025 -2928
rect 1465 -2929 1466 -2841
rect 79 -2931 80 -2841
rect 296 -2944 297 -2930
rect 422 -2944 423 -2930
rect 670 -2944 671 -2930
rect 1465 -2944 1466 -2930
rect 1472 -2931 1473 -2841
rect 79 -2944 80 -2932
rect 324 -2933 325 -2841
rect 471 -2944 472 -2932
rect 506 -2944 507 -2932
rect 233 -2935 234 -2841
rect 324 -2944 325 -2934
rect 233 -2944 234 -2936
rect 352 -2937 353 -2841
rect 352 -2944 353 -2938
rect 513 -2939 514 -2841
rect 443 -2941 444 -2841
rect 513 -2944 514 -2940
rect 156 -2943 157 -2841
rect 443 -2944 444 -2942
rect 30 -2954 31 -2952
rect 72 -3063 73 -2953
rect 79 -2954 80 -2952
rect 474 -2954 475 -2952
rect 523 -3063 524 -2953
rect 632 -2954 633 -2952
rect 635 -2954 636 -2952
rect 968 -2954 969 -2952
rect 982 -2954 983 -2952
rect 1024 -2954 1025 -2952
rect 1038 -2954 1039 -2952
rect 1041 -2972 1042 -2953
rect 1062 -3063 1063 -2953
rect 1430 -2954 1431 -2952
rect 1444 -2954 1445 -2952
rect 1486 -2954 1487 -2952
rect 37 -2956 38 -2952
rect 96 -3063 97 -2955
rect 100 -2956 101 -2952
rect 702 -2956 703 -2952
rect 758 -2956 759 -2952
rect 765 -2956 766 -2952
rect 821 -2956 822 -2952
rect 821 -3063 822 -2955
rect 821 -2956 822 -2952
rect 821 -3063 822 -2955
rect 828 -2956 829 -2952
rect 863 -2956 864 -2952
rect 870 -2956 871 -2952
rect 999 -2956 1000 -2952
rect 1020 -2956 1021 -2952
rect 1150 -2956 1151 -2952
rect 1199 -3063 1200 -2955
rect 1276 -2956 1277 -2952
rect 1447 -2956 1448 -2952
rect 1500 -2956 1501 -2952
rect 37 -3063 38 -2957
rect 121 -2958 122 -2952
rect 124 -3063 125 -2957
rect 310 -2958 311 -2952
rect 366 -2958 367 -2952
rect 852 -3063 853 -2957
rect 870 -3063 871 -2957
rect 1437 -2958 1438 -2952
rect 1472 -3063 1473 -2957
rect 1493 -2958 1494 -2952
rect 44 -2960 45 -2952
rect 250 -2960 251 -2952
rect 254 -2960 255 -2952
rect 324 -2960 325 -2952
rect 373 -2960 374 -2952
rect 450 -2960 451 -2952
rect 464 -2960 465 -2952
rect 670 -2960 671 -2952
rect 684 -3063 685 -2959
rect 1283 -2960 1284 -2952
rect 44 -3063 45 -2961
rect 149 -2962 150 -2952
rect 156 -3063 157 -2961
rect 380 -2962 381 -2952
rect 387 -2962 388 -2952
rect 387 -3063 388 -2961
rect 387 -2962 388 -2952
rect 387 -3063 388 -2961
rect 429 -2962 430 -2952
rect 478 -2962 479 -2952
rect 534 -2962 535 -2952
rect 642 -3063 643 -2961
rect 646 -2962 647 -2952
rect 933 -2962 934 -2952
rect 936 -2962 937 -2952
rect 982 -3063 983 -2961
rect 996 -2962 997 -2952
rect 1185 -2962 1186 -2952
rect 1255 -2962 1256 -2952
rect 1283 -3063 1284 -2961
rect 51 -2964 52 -2952
rect 607 -2964 608 -2952
rect 611 -2964 612 -2952
rect 730 -2964 731 -2952
rect 758 -3063 759 -2963
rect 835 -2964 836 -2952
rect 877 -2964 878 -2952
rect 1024 -3063 1025 -2963
rect 1038 -3063 1039 -2963
rect 1122 -2964 1123 -2952
rect 1143 -2964 1144 -2952
rect 1185 -3063 1186 -2963
rect 1255 -3063 1256 -2963
rect 1395 -2964 1396 -2952
rect 51 -3063 52 -2965
rect 408 -2966 409 -2952
rect 429 -3063 430 -2965
rect 796 -3063 797 -2965
rect 828 -3063 829 -2965
rect 1374 -2966 1375 -2952
rect 65 -2968 66 -2952
rect 79 -3063 80 -2967
rect 93 -2968 94 -2952
rect 621 -3063 622 -2967
rect 625 -2968 626 -2952
rect 765 -3063 766 -2967
rect 793 -2968 794 -2952
rect 877 -3063 878 -2967
rect 905 -2968 906 -2952
rect 905 -3063 906 -2967
rect 905 -2968 906 -2952
rect 905 -3063 906 -2967
rect 922 -3063 923 -2967
rect 1052 -2968 1053 -2952
rect 1073 -2968 1074 -2952
rect 1122 -3063 1123 -2967
rect 1143 -3063 1144 -2967
rect 1241 -2968 1242 -2952
rect 1276 -3063 1277 -2967
rect 1318 -2968 1319 -2952
rect 1374 -3063 1375 -2967
rect 1458 -2968 1459 -2952
rect 65 -3063 66 -2969
rect 250 -3063 251 -2969
rect 254 -3063 255 -2969
rect 275 -2970 276 -2952
rect 289 -2970 290 -2952
rect 366 -3063 367 -2969
rect 373 -3063 374 -2969
rect 597 -2970 598 -2952
rect 632 -3063 633 -2969
rect 723 -2970 724 -2952
rect 933 -3063 934 -2969
rect 989 -2970 990 -2952
rect 996 -3063 997 -2969
rect 1332 -2970 1333 -2952
rect 1458 -3063 1459 -2969
rect 1465 -2970 1466 -2952
rect 100 -3063 101 -2971
rect 541 -2972 542 -2952
rect 555 -2972 556 -2952
rect 863 -3063 864 -2971
rect 954 -2972 955 -2952
rect 968 -3063 969 -2971
rect 1073 -3063 1074 -2971
rect 1090 -3063 1091 -2971
rect 1409 -2972 1410 -2952
rect 1465 -3063 1466 -2971
rect 1479 -2972 1480 -2952
rect 114 -2974 115 -2952
rect 149 -3063 150 -2973
rect 159 -2974 160 -2952
rect 520 -2974 521 -2952
rect 527 -2974 528 -2952
rect 541 -3063 542 -2973
rect 555 -3063 556 -2973
rect 873 -3063 874 -2973
rect 954 -3063 955 -2973
rect 1003 -2974 1004 -2952
rect 1052 -3063 1053 -2973
rect 1129 -2974 1130 -2952
rect 1136 -2974 1137 -2952
rect 1318 -3063 1319 -2973
rect 1332 -3063 1333 -2973
rect 1451 -2974 1452 -2952
rect 114 -3063 115 -2975
rect 135 -2976 136 -2952
rect 177 -2976 178 -2952
rect 289 -3063 290 -2975
rect 352 -2976 353 -2952
rect 607 -3063 608 -2975
rect 646 -3063 647 -2975
rect 695 -2976 696 -2952
rect 723 -3063 724 -2975
rect 912 -2976 913 -2952
rect 1003 -3063 1004 -2975
rect 1059 -2976 1060 -2952
rect 1129 -3063 1130 -2975
rect 1171 -2976 1172 -2952
rect 121 -3063 122 -2977
rect 135 -3063 136 -2977
rect 177 -3063 178 -2977
rect 1325 -2978 1326 -2952
rect 180 -2980 181 -2952
rect 394 -2980 395 -2952
rect 408 -3063 409 -2979
rect 464 -3063 465 -2979
rect 534 -3063 535 -2979
rect 744 -2980 745 -2952
rect 912 -3063 913 -2979
rect 975 -2980 976 -2952
rect 1080 -2980 1081 -2952
rect 1171 -3063 1172 -2979
rect 198 -2982 199 -2952
rect 604 -2982 605 -2952
rect 653 -2982 654 -2952
rect 989 -3063 990 -2981
rect 1080 -3063 1081 -2981
rect 1108 -2982 1109 -2952
rect 1136 -3063 1137 -2981
rect 1227 -2982 1228 -2952
rect 201 -3063 202 -2983
rect 513 -2984 514 -2952
rect 562 -3063 563 -2983
rect 800 -2984 801 -2952
rect 1108 -3063 1109 -2983
rect 1269 -2984 1270 -2952
rect 219 -2986 220 -2952
rect 380 -3063 381 -2985
rect 394 -3063 395 -2985
rect 866 -2986 867 -2952
rect 1150 -3063 1151 -2985
rect 1262 -2986 1263 -2952
rect 226 -2988 227 -2952
rect 324 -3063 325 -2987
rect 352 -3063 353 -2987
rect 415 -2988 416 -2952
rect 422 -2988 423 -2952
rect 527 -3063 528 -2987
rect 565 -2988 566 -2952
rect 737 -2988 738 -2952
rect 800 -3063 801 -2987
rect 814 -2988 815 -2952
rect 1094 -2988 1095 -2952
rect 1262 -3063 1263 -2987
rect 170 -2990 171 -2952
rect 226 -3063 227 -2989
rect 233 -2990 234 -2952
rect 310 -3063 311 -2989
rect 355 -3063 356 -2989
rect 478 -3063 479 -2989
rect 506 -2990 507 -2952
rect 814 -3063 815 -2989
rect 1094 -3063 1095 -2989
rect 1192 -2990 1193 -2952
rect 1213 -2990 1214 -2952
rect 1269 -3063 1270 -2989
rect 128 -2992 129 -2952
rect 233 -3063 234 -2991
rect 243 -3063 244 -2991
rect 761 -2992 762 -2952
rect 1157 -2992 1158 -2952
rect 1213 -3063 1214 -2991
rect 1227 -3063 1228 -2991
rect 1304 -2992 1305 -2952
rect 58 -2994 59 -2952
rect 128 -3063 129 -2993
rect 170 -3063 171 -2993
rect 205 -2994 206 -2952
rect 257 -2994 258 -2952
rect 422 -3063 423 -2993
rect 443 -2994 444 -2952
rect 499 -3063 500 -2993
rect 506 -3063 507 -2993
rect 716 -2994 717 -2952
rect 1031 -2994 1032 -2952
rect 1304 -3063 1305 -2993
rect 58 -3063 59 -2995
rect 163 -2996 164 -2952
rect 205 -3063 206 -2995
rect 520 -3063 521 -2995
rect 569 -2996 570 -2952
rect 688 -2996 689 -2952
rect 691 -2996 692 -2952
rect 1087 -2996 1088 -2952
rect 1157 -3063 1158 -2995
rect 1178 -2996 1179 -2952
rect 1192 -3063 1193 -2995
rect 1234 -2996 1235 -2952
rect 86 -2998 87 -2952
rect 443 -3063 444 -2997
rect 450 -3063 451 -2997
rect 548 -2998 549 -2952
rect 569 -3063 570 -2997
rect 583 -2998 584 -2952
rect 590 -2998 591 -2952
rect 740 -3063 741 -2997
rect 1031 -3063 1032 -2997
rect 1066 -2998 1067 -2952
rect 1087 -3063 1088 -2997
rect 1325 -3063 1326 -2997
rect 86 -3063 87 -2999
rect 376 -3000 377 -2952
rect 401 -3000 402 -2952
rect 744 -3063 745 -2999
rect 1066 -3063 1067 -2999
rect 1101 -3000 1102 -2952
rect 1178 -3063 1179 -2999
rect 1381 -3000 1382 -2952
rect 163 -3063 164 -3001
rect 618 -3002 619 -2952
rect 639 -3002 640 -2952
rect 653 -3063 654 -3001
rect 667 -3002 668 -2952
rect 1353 -3002 1354 -2952
rect 1381 -3063 1382 -3001
rect 1416 -3002 1417 -2952
rect 261 -3004 262 -2952
rect 548 -3063 549 -3003
rect 590 -3063 591 -3003
rect 898 -3004 899 -2952
rect 926 -3004 927 -2952
rect 1101 -3063 1102 -3003
rect 1234 -3063 1235 -3003
rect 1339 -3004 1340 -2952
rect 1416 -3063 1417 -3003
rect 1423 -3004 1424 -2952
rect 142 -3006 143 -2952
rect 261 -3063 262 -3005
rect 264 -3006 265 -2952
rect 268 -3006 269 -2952
rect 275 -3063 276 -3005
rect 457 -3006 458 -2952
rect 502 -3006 503 -2952
rect 583 -3063 584 -3005
rect 597 -3063 598 -3005
rect 849 -3006 850 -2952
rect 898 -3063 899 -3005
rect 1223 -3063 1224 -3005
rect 1311 -3006 1312 -2952
rect 1339 -3063 1340 -3005
rect 107 -3008 108 -2952
rect 457 -3063 458 -3007
rect 604 -3063 605 -3007
rect 891 -3008 892 -2952
rect 1311 -3063 1312 -3007
rect 1388 -3008 1389 -2952
rect 107 -3063 108 -3009
rect 492 -3010 493 -2952
rect 611 -3063 612 -3009
rect 926 -3063 927 -3009
rect 142 -3063 143 -3011
rect 184 -3012 185 -2952
rect 264 -3063 265 -3011
rect 772 -3012 773 -2952
rect 891 -3063 892 -3011
rect 919 -3012 920 -2952
rect 184 -3063 185 -3013
rect 191 -3014 192 -2952
rect 268 -3063 269 -3013
rect 338 -3014 339 -2952
rect 359 -3014 360 -2952
rect 625 -3063 626 -3013
rect 639 -3063 640 -3013
rect 1346 -3014 1347 -2952
rect 191 -3063 192 -3015
rect 485 -3016 486 -2952
rect 492 -3063 493 -3015
rect 660 -3016 661 -2952
rect 667 -3063 668 -3015
rect 940 -3016 941 -2952
rect 1346 -3063 1347 -3015
rect 1402 -3016 1403 -2952
rect 282 -3018 283 -2952
rect 772 -3063 773 -3017
rect 940 -3063 941 -3017
rect 961 -3018 962 -2952
rect 282 -3063 283 -3019
rect 331 -3020 332 -2952
rect 338 -3063 339 -3019
rect 345 -3020 346 -2952
rect 401 -3063 402 -3019
rect 471 -3020 472 -2952
rect 485 -3063 486 -3019
rect 733 -3020 734 -2952
rect 807 -3020 808 -2952
rect 961 -3063 962 -3019
rect 296 -3022 297 -2952
rect 359 -3063 360 -3021
rect 404 -3022 405 -2952
rect 513 -3063 514 -3021
rect 576 -3022 577 -2952
rect 919 -3063 920 -3021
rect 296 -3063 297 -3023
rect 835 -3063 836 -3023
rect 317 -3026 318 -2952
rect 576 -3063 577 -3025
rect 618 -3063 619 -3025
rect 975 -3063 976 -3025
rect 303 -3028 304 -2952
rect 317 -3063 318 -3027
rect 331 -3063 332 -3027
rect 481 -3028 482 -2952
rect 660 -3063 661 -3027
rect 709 -3028 710 -2952
rect 716 -3063 717 -3027
rect 779 -3028 780 -2952
rect 303 -3063 304 -3029
rect 999 -3063 1000 -3029
rect 345 -3063 346 -3031
rect 436 -3032 437 -2952
rect 471 -3063 472 -3031
rect 705 -3032 706 -2952
rect 779 -3063 780 -3031
rect 786 -3032 787 -2952
rect 212 -3034 213 -2952
rect 436 -3063 437 -3033
rect 674 -3034 675 -2952
rect 730 -3063 731 -3033
rect 786 -3063 787 -3033
rect 849 -3063 850 -3033
rect 212 -3063 213 -3035
rect 240 -3036 241 -2952
rect 247 -3063 248 -3035
rect 674 -3063 675 -3035
rect 681 -3036 682 -2952
rect 709 -3063 710 -3035
rect 411 -3063 412 -3037
rect 415 -3063 416 -3037
rect 681 -3063 682 -3037
rect 884 -3038 885 -2952
rect 688 -3063 689 -3039
rect 842 -3040 843 -2952
rect 856 -3040 857 -2952
rect 884 -3063 885 -3039
rect 695 -3063 696 -3041
rect 751 -3042 752 -2952
rect 842 -3063 843 -3041
rect 947 -3042 948 -2952
rect 702 -3063 703 -3043
rect 807 -3063 808 -3043
rect 856 -3063 857 -3043
rect 1017 -3044 1018 -2952
rect 705 -3063 706 -3045
rect 1241 -3063 1242 -3045
rect 751 -3063 752 -3047
rect 929 -3048 930 -2952
rect 947 -3063 948 -3047
rect 1010 -3048 1011 -2952
rect 1017 -3063 1018 -3047
rect 1115 -3048 1116 -2952
rect 1010 -3063 1011 -3049
rect 1045 -3050 1046 -2952
rect 1115 -3063 1116 -3049
rect 1206 -3050 1207 -2952
rect 1045 -3063 1046 -3051
rect 1164 -3052 1165 -2952
rect 1206 -3063 1207 -3051
rect 1367 -3052 1368 -2952
rect 1164 -3063 1165 -3053
rect 1220 -3054 1221 -2952
rect 1220 -3063 1221 -3055
rect 1248 -3056 1249 -2952
rect 1248 -3063 1249 -3057
rect 1297 -3058 1298 -2952
rect 1290 -3060 1291 -2952
rect 1297 -3063 1298 -3059
rect 1290 -3063 1291 -3061
rect 1360 -3062 1361 -2952
rect 37 -3073 38 -3071
rect 96 -3073 97 -3071
rect 100 -3073 101 -3071
rect 579 -3152 580 -3072
rect 590 -3073 591 -3071
rect 590 -3152 591 -3072
rect 590 -3073 591 -3071
rect 590 -3152 591 -3072
rect 621 -3073 622 -3071
rect 744 -3073 745 -3071
rect 775 -3152 776 -3072
rect 1248 -3073 1249 -3071
rect 1262 -3073 1263 -3071
rect 1286 -3073 1287 -3071
rect 1293 -3152 1294 -3072
rect 1297 -3073 1298 -3071
rect 1339 -3073 1340 -3071
rect 1353 -3152 1354 -3072
rect 1367 -3152 1368 -3072
rect 1381 -3073 1382 -3071
rect 1409 -3152 1410 -3072
rect 1416 -3073 1417 -3071
rect 1451 -3152 1452 -3072
rect 1458 -3073 1459 -3071
rect 44 -3075 45 -3071
rect 219 -3152 220 -3074
rect 240 -3075 241 -3071
rect 982 -3075 983 -3071
rect 1010 -3075 1011 -3071
rect 1087 -3075 1088 -3071
rect 1090 -3152 1091 -3074
rect 1269 -3075 1270 -3071
rect 1283 -3075 1284 -3071
rect 1346 -3075 1347 -3071
rect 1458 -3152 1459 -3074
rect 1465 -3075 1466 -3071
rect 51 -3077 52 -3071
rect 215 -3152 216 -3076
rect 226 -3077 227 -3071
rect 240 -3152 241 -3076
rect 243 -3077 244 -3071
rect 338 -3077 339 -3071
rect 373 -3077 374 -3071
rect 621 -3152 622 -3076
rect 639 -3152 640 -3076
rect 807 -3077 808 -3071
rect 849 -3077 850 -3071
rect 968 -3077 969 -3071
rect 982 -3152 983 -3076
rect 1115 -3077 1116 -3071
rect 1143 -3077 1144 -3071
rect 1143 -3152 1144 -3076
rect 1143 -3077 1144 -3071
rect 1143 -3152 1144 -3076
rect 1171 -3077 1172 -3071
rect 1171 -3152 1172 -3076
rect 1171 -3077 1172 -3071
rect 1171 -3152 1172 -3076
rect 1220 -3077 1221 -3071
rect 1290 -3077 1291 -3071
rect 1346 -3152 1347 -3076
rect 1374 -3077 1375 -3071
rect 1465 -3152 1466 -3076
rect 1472 -3077 1473 -3071
rect 58 -3079 59 -3071
rect 180 -3079 181 -3071
rect 191 -3079 192 -3071
rect 250 -3079 251 -3071
rect 254 -3079 255 -3071
rect 254 -3152 255 -3078
rect 254 -3079 255 -3071
rect 254 -3152 255 -3078
rect 289 -3079 290 -3071
rect 607 -3152 608 -3078
rect 653 -3079 654 -3071
rect 705 -3079 706 -3071
rect 740 -3079 741 -3071
rect 968 -3152 969 -3078
rect 1010 -3152 1011 -3078
rect 1052 -3079 1053 -3071
rect 1059 -3152 1060 -3078
rect 1241 -3079 1242 -3071
rect 1262 -3152 1263 -3078
rect 1332 -3079 1333 -3071
rect 72 -3081 73 -3071
rect 187 -3152 188 -3080
rect 191 -3152 192 -3080
rect 268 -3081 269 -3071
rect 299 -3081 300 -3071
rect 324 -3081 325 -3071
rect 338 -3152 339 -3080
rect 464 -3081 465 -3071
rect 513 -3081 514 -3071
rect 737 -3081 738 -3071
rect 744 -3152 745 -3080
rect 800 -3081 801 -3071
rect 807 -3152 808 -3080
rect 856 -3081 857 -3071
rect 870 -3081 871 -3071
rect 947 -3081 948 -3071
rect 961 -3081 962 -3071
rect 1136 -3081 1137 -3071
rect 1164 -3081 1165 -3071
rect 1220 -3152 1221 -3080
rect 1230 -3152 1231 -3080
rect 1311 -3081 1312 -3071
rect 79 -3083 80 -3071
rect 408 -3083 409 -3071
rect 436 -3083 437 -3071
rect 1062 -3083 1063 -3071
rect 1066 -3083 1067 -3071
rect 1115 -3152 1116 -3082
rect 1136 -3152 1137 -3082
rect 1234 -3083 1235 -3071
rect 79 -3152 80 -3084
rect 93 -3085 94 -3071
rect 100 -3152 101 -3084
rect 114 -3085 115 -3071
rect 121 -3085 122 -3071
rect 737 -3152 738 -3084
rect 782 -3152 783 -3084
rect 1038 -3085 1039 -3071
rect 1052 -3152 1053 -3084
rect 1255 -3085 1256 -3071
rect 86 -3087 87 -3071
rect 355 -3087 356 -3071
rect 373 -3152 374 -3086
rect 471 -3087 472 -3071
rect 478 -3087 479 -3071
rect 800 -3152 801 -3086
rect 873 -3087 874 -3071
rect 905 -3087 906 -3071
rect 929 -3087 930 -3071
rect 1276 -3087 1277 -3071
rect 65 -3089 66 -3071
rect 86 -3152 87 -3088
rect 93 -3152 94 -3088
rect 163 -3089 164 -3071
rect 177 -3089 178 -3071
rect 415 -3089 416 -3071
rect 436 -3152 437 -3088
rect 520 -3089 521 -3071
rect 523 -3089 524 -3071
rect 877 -3089 878 -3071
rect 884 -3089 885 -3071
rect 919 -3089 920 -3071
rect 933 -3089 934 -3071
rect 947 -3152 948 -3088
rect 964 -3089 965 -3071
rect 1185 -3089 1186 -3071
rect 1276 -3152 1277 -3088
rect 1325 -3089 1326 -3071
rect 107 -3091 108 -3071
rect 107 -3152 108 -3090
rect 107 -3091 108 -3071
rect 107 -3152 108 -3090
rect 114 -3152 115 -3090
rect 128 -3091 129 -3071
rect 142 -3091 143 -3071
rect 222 -3091 223 -3071
rect 226 -3152 227 -3090
rect 635 -3152 636 -3090
rect 656 -3152 657 -3090
rect 828 -3091 829 -3071
rect 884 -3152 885 -3090
rect 891 -3091 892 -3071
rect 905 -3152 906 -3090
rect 964 -3152 965 -3090
rect 996 -3091 997 -3071
rect 1038 -3152 1039 -3090
rect 1066 -3152 1067 -3090
rect 1094 -3091 1095 -3071
rect 1101 -3091 1102 -3071
rect 1290 -3152 1291 -3090
rect 121 -3152 122 -3092
rect 156 -3093 157 -3071
rect 163 -3152 164 -3092
rect 205 -3093 206 -3071
rect 247 -3093 248 -3071
rect 362 -3152 363 -3092
rect 366 -3093 367 -3071
rect 478 -3152 479 -3092
rect 520 -3152 521 -3092
rect 611 -3093 612 -3071
rect 618 -3093 619 -3071
rect 877 -3152 878 -3092
rect 912 -3093 913 -3071
rect 933 -3152 934 -3092
rect 940 -3093 941 -3071
rect 961 -3152 962 -3092
rect 975 -3093 976 -3071
rect 1094 -3152 1095 -3092
rect 1101 -3152 1102 -3092
rect 1199 -3093 1200 -3071
rect 142 -3152 143 -3094
rect 170 -3095 171 -3071
rect 177 -3152 178 -3094
rect 184 -3095 185 -3071
rect 198 -3095 199 -3071
rect 688 -3095 689 -3071
rect 702 -3095 703 -3071
rect 1073 -3095 1074 -3071
rect 1129 -3095 1130 -3071
rect 1199 -3152 1200 -3094
rect 149 -3097 150 -3071
rect 149 -3152 150 -3096
rect 149 -3097 150 -3071
rect 149 -3152 150 -3096
rect 156 -3152 157 -3096
rect 296 -3097 297 -3071
rect 303 -3097 304 -3071
rect 513 -3152 514 -3096
rect 527 -3097 528 -3071
rect 919 -3152 920 -3096
rect 940 -3152 941 -3096
rect 954 -3097 955 -3071
rect 1017 -3097 1018 -3071
rect 1017 -3152 1018 -3096
rect 1017 -3097 1018 -3071
rect 1017 -3152 1018 -3096
rect 1073 -3152 1074 -3096
rect 1206 -3097 1207 -3071
rect 128 -3152 129 -3098
rect 303 -3152 304 -3098
rect 366 -3152 367 -3098
rect 856 -3152 857 -3098
rect 898 -3099 899 -3071
rect 954 -3152 955 -3098
rect 1164 -3152 1165 -3098
rect 1223 -3099 1224 -3071
rect 170 -3152 171 -3100
rect 275 -3101 276 -3071
rect 296 -3152 297 -3100
rect 387 -3101 388 -3071
rect 394 -3101 395 -3071
rect 415 -3152 416 -3100
rect 464 -3152 465 -3100
rect 642 -3101 643 -3071
rect 674 -3101 675 -3071
rect 870 -3152 871 -3100
rect 898 -3152 899 -3100
rect 1031 -3101 1032 -3071
rect 1206 -3152 1207 -3100
rect 1304 -3101 1305 -3071
rect 198 -3152 199 -3102
rect 282 -3103 283 -3071
rect 352 -3103 353 -3071
rect 674 -3152 675 -3102
rect 684 -3103 685 -3071
rect 772 -3103 773 -3071
rect 786 -3103 787 -3071
rect 849 -3152 850 -3102
rect 912 -3152 913 -3102
rect 1080 -3103 1081 -3071
rect 201 -3105 202 -3071
rect 324 -3152 325 -3104
rect 352 -3152 353 -3104
rect 429 -3105 430 -3071
rect 471 -3152 472 -3104
rect 597 -3105 598 -3071
rect 765 -3105 766 -3071
rect 786 -3152 787 -3104
rect 793 -3105 794 -3071
rect 1024 -3105 1025 -3071
rect 1031 -3152 1032 -3104
rect 1108 -3105 1109 -3071
rect 233 -3107 234 -3071
rect 247 -3152 248 -3106
rect 261 -3107 262 -3071
rect 394 -3152 395 -3106
rect 401 -3107 402 -3071
rect 845 -3152 846 -3106
rect 1024 -3152 1025 -3106
rect 1122 -3107 1123 -3071
rect 212 -3109 213 -3071
rect 261 -3152 262 -3108
rect 268 -3152 269 -3108
rect 310 -3109 311 -3071
rect 380 -3109 381 -3071
rect 383 -3141 384 -3108
rect 387 -3152 388 -3108
rect 681 -3109 682 -3071
rect 723 -3109 724 -3071
rect 765 -3152 766 -3108
rect 796 -3109 797 -3071
rect 880 -3152 881 -3108
rect 1080 -3152 1081 -3108
rect 1227 -3109 1228 -3071
rect 222 -3152 223 -3110
rect 401 -3152 402 -3110
rect 408 -3152 409 -3110
rect 485 -3111 486 -3071
rect 506 -3111 507 -3071
rect 597 -3152 598 -3110
rect 681 -3152 682 -3110
rect 695 -3111 696 -3071
rect 723 -3152 724 -3110
rect 758 -3111 759 -3071
rect 835 -3111 836 -3071
rect 891 -3152 892 -3110
rect 1108 -3152 1109 -3110
rect 1150 -3111 1151 -3071
rect 233 -3152 234 -3112
rect 331 -3113 332 -3071
rect 380 -3152 381 -3112
rect 604 -3113 605 -3071
rect 695 -3152 696 -3112
rect 709 -3113 710 -3071
rect 758 -3152 759 -3112
rect 842 -3113 843 -3071
rect 1122 -3152 1123 -3112
rect 1178 -3113 1179 -3071
rect 275 -3152 276 -3114
rect 345 -3115 346 -3071
rect 485 -3152 486 -3114
rect 653 -3152 654 -3114
rect 709 -3152 710 -3114
rect 730 -3115 731 -3071
rect 828 -3152 829 -3114
rect 842 -3152 843 -3114
rect 1129 -3152 1130 -3114
rect 1227 -3152 1228 -3114
rect 282 -3152 283 -3116
rect 555 -3117 556 -3071
rect 576 -3117 577 -3071
rect 611 -3152 612 -3116
rect 835 -3152 836 -3116
rect 926 -3117 927 -3071
rect 1150 -3152 1151 -3116
rect 1188 -3152 1189 -3116
rect 289 -3152 290 -3118
rect 730 -3152 731 -3118
rect 814 -3119 815 -3071
rect 926 -3152 927 -3118
rect 1178 -3152 1179 -3118
rect 1192 -3119 1193 -3071
rect 310 -3152 311 -3120
rect 457 -3121 458 -3071
rect 506 -3152 507 -3120
rect 632 -3121 633 -3071
rect 814 -3152 815 -3120
rect 821 -3121 822 -3071
rect 1192 -3152 1193 -3120
rect 1318 -3121 1319 -3071
rect 317 -3123 318 -3071
rect 331 -3152 332 -3122
rect 345 -3152 346 -3122
rect 359 -3123 360 -3071
rect 457 -3152 458 -3122
rect 772 -3152 773 -3122
rect 821 -3152 822 -3122
rect 1045 -3123 1046 -3071
rect 135 -3125 136 -3071
rect 317 -3152 318 -3124
rect 527 -3152 528 -3124
rect 625 -3125 626 -3071
rect 1045 -3152 1046 -3124
rect 1213 -3125 1214 -3071
rect 205 -3152 206 -3126
rect 359 -3152 360 -3126
rect 534 -3127 535 -3071
rect 632 -3152 633 -3126
rect 1157 -3127 1158 -3071
rect 1213 -3152 1214 -3126
rect 450 -3129 451 -3071
rect 534 -3152 535 -3128
rect 541 -3129 542 -3071
rect 555 -3152 556 -3128
rect 583 -3129 584 -3071
rect 793 -3152 794 -3128
rect 1157 -3152 1158 -3128
rect 1241 -3152 1242 -3128
rect 450 -3152 451 -3130
rect 548 -3131 549 -3071
rect 604 -3152 605 -3130
rect 863 -3131 864 -3071
rect 422 -3133 423 -3071
rect 548 -3152 549 -3132
rect 625 -3152 626 -3132
rect 716 -3133 717 -3071
rect 863 -3152 864 -3132
rect 989 -3133 990 -3071
rect 422 -3152 423 -3134
rect 576 -3152 577 -3134
rect 716 -3152 717 -3134
rect 779 -3135 780 -3071
rect 989 -3152 990 -3134
rect 1003 -3135 1004 -3071
rect 492 -3137 493 -3071
rect 1003 -3152 1004 -3136
rect 443 -3139 444 -3071
rect 492 -3152 493 -3138
rect 499 -3139 500 -3071
rect 583 -3152 584 -3138
rect 779 -3152 780 -3138
rect 975 -3152 976 -3138
rect 443 -3152 444 -3140
rect 499 -3152 500 -3140
rect 569 -3141 570 -3071
rect 541 -3152 542 -3142
rect 646 -3143 647 -3071
rect 562 -3145 563 -3071
rect 646 -3152 647 -3144
rect 562 -3152 563 -3146
rect 751 -3147 752 -3071
rect 569 -3152 570 -3148
rect 660 -3149 661 -3071
rect 667 -3149 668 -3071
rect 751 -3152 752 -3148
rect 135 -3152 136 -3150
rect 660 -3152 661 -3150
rect 667 -3152 668 -3150
rect 705 -3152 706 -3150
rect 58 -3213 59 -3161
rect 198 -3162 199 -3160
rect 219 -3213 220 -3161
rect 352 -3162 353 -3160
rect 373 -3162 374 -3160
rect 429 -3213 430 -3161
rect 432 -3162 433 -3160
rect 555 -3162 556 -3160
rect 569 -3162 570 -3160
rect 579 -3162 580 -3160
rect 611 -3162 612 -3160
rect 663 -3162 664 -3160
rect 667 -3162 668 -3160
rect 779 -3162 780 -3160
rect 793 -3162 794 -3160
rect 842 -3213 843 -3161
rect 845 -3162 846 -3160
rect 1017 -3162 1018 -3160
rect 1080 -3162 1081 -3160
rect 1087 -3213 1088 -3161
rect 1094 -3162 1095 -3160
rect 1097 -3162 1098 -3160
rect 1101 -3162 1102 -3160
rect 1101 -3213 1102 -3161
rect 1101 -3162 1102 -3160
rect 1101 -3213 1102 -3161
rect 1188 -3162 1189 -3160
rect 1262 -3162 1263 -3160
rect 1332 -3213 1333 -3161
rect 1346 -3162 1347 -3160
rect 1353 -3162 1354 -3160
rect 1360 -3213 1361 -3161
rect 1367 -3162 1368 -3160
rect 1367 -3213 1368 -3161
rect 1367 -3162 1368 -3160
rect 1367 -3213 1368 -3161
rect 1409 -3162 1410 -3160
rect 1409 -3213 1410 -3161
rect 1409 -3162 1410 -3160
rect 1409 -3213 1410 -3161
rect 1451 -3162 1452 -3160
rect 1451 -3213 1452 -3161
rect 1451 -3162 1452 -3160
rect 1451 -3213 1452 -3161
rect 1458 -3162 1459 -3160
rect 1458 -3213 1459 -3161
rect 1458 -3162 1459 -3160
rect 1458 -3213 1459 -3161
rect 1465 -3162 1466 -3160
rect 1465 -3213 1466 -3161
rect 1465 -3162 1466 -3160
rect 1465 -3213 1466 -3161
rect 65 -3213 66 -3163
rect 135 -3164 136 -3160
rect 145 -3213 146 -3163
rect 187 -3164 188 -3160
rect 306 -3164 307 -3160
rect 338 -3164 339 -3160
rect 352 -3213 353 -3163
rect 387 -3164 388 -3160
rect 415 -3164 416 -3160
rect 418 -3188 419 -3163
rect 471 -3164 472 -3160
rect 635 -3213 636 -3163
rect 653 -3213 654 -3163
rect 737 -3164 738 -3160
rect 751 -3164 752 -3160
rect 793 -3213 794 -3163
rect 856 -3164 857 -3160
rect 1052 -3164 1053 -3160
rect 1080 -3213 1081 -3163
rect 1108 -3164 1109 -3160
rect 1199 -3164 1200 -3160
rect 1199 -3213 1200 -3163
rect 1199 -3164 1200 -3160
rect 1199 -3213 1200 -3163
rect 1213 -3164 1214 -3160
rect 1213 -3213 1214 -3163
rect 1213 -3164 1214 -3160
rect 1213 -3213 1214 -3163
rect 1220 -3164 1221 -3160
rect 1241 -3164 1242 -3160
rect 72 -3213 73 -3165
rect 205 -3166 206 -3160
rect 296 -3166 297 -3160
rect 338 -3213 339 -3165
rect 373 -3213 374 -3165
rect 499 -3166 500 -3160
rect 513 -3166 514 -3160
rect 611 -3213 612 -3165
rect 618 -3166 619 -3160
rect 709 -3166 710 -3160
rect 716 -3166 717 -3160
rect 737 -3213 738 -3165
rect 761 -3213 762 -3165
rect 772 -3166 773 -3160
rect 775 -3166 776 -3160
rect 835 -3166 836 -3160
rect 856 -3213 857 -3165
rect 870 -3166 871 -3160
rect 877 -3213 878 -3165
rect 968 -3166 969 -3160
rect 975 -3166 976 -3160
rect 975 -3213 976 -3165
rect 975 -3166 976 -3160
rect 975 -3213 976 -3165
rect 985 -3213 986 -3165
rect 1122 -3166 1123 -3160
rect 1227 -3166 1228 -3160
rect 1234 -3213 1235 -3165
rect 1237 -3166 1238 -3160
rect 1276 -3166 1277 -3160
rect 79 -3168 80 -3160
rect 215 -3168 216 -3160
rect 250 -3213 251 -3167
rect 716 -3213 717 -3167
rect 723 -3168 724 -3160
rect 723 -3213 724 -3167
rect 723 -3168 724 -3160
rect 723 -3213 724 -3167
rect 733 -3168 734 -3160
rect 912 -3168 913 -3160
rect 919 -3168 920 -3160
rect 1052 -3213 1053 -3167
rect 1094 -3213 1095 -3167
rect 1129 -3168 1130 -3160
rect 79 -3213 80 -3169
rect 156 -3170 157 -3160
rect 180 -3213 181 -3169
rect 667 -3213 668 -3169
rect 688 -3170 689 -3160
rect 891 -3170 892 -3160
rect 912 -3213 913 -3169
rect 947 -3170 948 -3160
rect 964 -3170 965 -3160
rect 989 -3170 990 -3160
rect 999 -3170 1000 -3160
rect 1038 -3170 1039 -3160
rect 1122 -3213 1123 -3169
rect 1192 -3170 1193 -3160
rect 93 -3172 94 -3160
rect 205 -3213 206 -3171
rect 327 -3213 328 -3171
rect 362 -3172 363 -3160
rect 387 -3213 388 -3171
rect 656 -3172 657 -3160
rect 660 -3172 661 -3160
rect 821 -3172 822 -3160
rect 835 -3213 836 -3171
rect 954 -3172 955 -3160
rect 968 -3213 969 -3171
rect 1059 -3172 1060 -3160
rect 1129 -3213 1130 -3171
rect 1136 -3172 1137 -3160
rect 1192 -3213 1193 -3171
rect 1293 -3172 1294 -3160
rect 93 -3213 94 -3173
rect 170 -3174 171 -3160
rect 201 -3213 202 -3173
rect 296 -3213 297 -3173
rect 401 -3174 402 -3160
rect 471 -3213 472 -3173
rect 492 -3174 493 -3160
rect 499 -3213 500 -3173
rect 534 -3174 535 -3160
rect 537 -3188 538 -3173
rect 541 -3174 542 -3160
rect 866 -3213 867 -3173
rect 870 -3213 871 -3173
rect 898 -3174 899 -3160
rect 933 -3174 934 -3160
rect 947 -3213 948 -3173
rect 989 -3213 990 -3173
rect 1045 -3174 1046 -3160
rect 100 -3176 101 -3160
rect 152 -3213 153 -3175
rect 156 -3213 157 -3175
rect 191 -3176 192 -3160
rect 324 -3176 325 -3160
rect 401 -3213 402 -3175
rect 415 -3213 416 -3175
rect 464 -3176 465 -3160
rect 534 -3213 535 -3175
rect 548 -3176 549 -3160
rect 569 -3213 570 -3175
rect 807 -3176 808 -3160
rect 863 -3176 864 -3160
rect 919 -3213 920 -3175
rect 933 -3213 934 -3175
rect 1031 -3176 1032 -3160
rect 1045 -3213 1046 -3175
rect 1073 -3176 1074 -3160
rect 100 -3213 101 -3177
rect 264 -3213 265 -3177
rect 268 -3178 269 -3160
rect 324 -3213 325 -3177
rect 422 -3178 423 -3160
rect 513 -3213 514 -3177
rect 541 -3213 542 -3177
rect 646 -3178 647 -3160
rect 660 -3213 661 -3177
rect 1024 -3178 1025 -3160
rect 1031 -3213 1032 -3177
rect 1244 -3178 1245 -3160
rect 114 -3180 115 -3160
rect 208 -3213 209 -3179
rect 247 -3180 248 -3160
rect 268 -3213 269 -3179
rect 422 -3213 423 -3179
rect 443 -3180 444 -3160
rect 464 -3213 465 -3179
rect 485 -3180 486 -3160
rect 492 -3213 493 -3179
rect 863 -3213 864 -3179
rect 880 -3180 881 -3160
rect 898 -3213 899 -3179
rect 940 -3180 941 -3160
rect 954 -3213 955 -3179
rect 1006 -3213 1007 -3179
rect 1066 -3180 1067 -3160
rect 1073 -3213 1074 -3179
rect 1150 -3180 1151 -3160
rect 121 -3182 122 -3160
rect 198 -3213 199 -3181
rect 436 -3182 437 -3160
rect 772 -3213 773 -3181
rect 779 -3213 780 -3181
rect 926 -3182 927 -3160
rect 1010 -3182 1011 -3160
rect 1038 -3213 1039 -3181
rect 1115 -3182 1116 -3160
rect 1150 -3213 1151 -3181
rect 121 -3213 122 -3183
rect 226 -3184 227 -3160
rect 282 -3184 283 -3160
rect 436 -3213 437 -3183
rect 443 -3213 444 -3183
rect 702 -3184 703 -3160
rect 705 -3184 706 -3160
rect 1017 -3213 1018 -3183
rect 1024 -3213 1025 -3183
rect 1157 -3184 1158 -3160
rect 128 -3186 129 -3160
rect 128 -3213 129 -3185
rect 128 -3186 129 -3160
rect 128 -3213 129 -3185
rect 131 -3213 132 -3185
rect 184 -3213 185 -3185
rect 282 -3213 283 -3185
rect 345 -3186 346 -3160
rect 485 -3213 486 -3185
rect 548 -3213 549 -3185
rect 674 -3186 675 -3160
rect 681 -3186 682 -3160
rect 688 -3213 689 -3185
rect 695 -3186 696 -3160
rect 709 -3213 710 -3185
rect 765 -3186 766 -3160
rect 821 -3213 822 -3185
rect 884 -3186 885 -3160
rect 996 -3186 997 -3160
rect 1115 -3213 1116 -3185
rect 1185 -3186 1186 -3160
rect 135 -3213 136 -3187
rect 457 -3188 458 -3160
rect 506 -3188 507 -3160
rect 681 -3213 682 -3187
rect 800 -3188 801 -3160
rect 891 -3213 892 -3187
rect 905 -3188 906 -3160
rect 940 -3213 941 -3187
rect 1097 -3213 1098 -3187
rect 1136 -3213 1137 -3187
rect 1143 -3188 1144 -3160
rect 1185 -3213 1186 -3187
rect 142 -3190 143 -3160
rect 191 -3213 192 -3189
rect 331 -3190 332 -3160
rect 345 -3213 346 -3189
rect 359 -3190 360 -3160
rect 996 -3213 997 -3189
rect 1143 -3213 1144 -3189
rect 1164 -3190 1165 -3160
rect 86 -3192 87 -3160
rect 142 -3213 143 -3191
rect 149 -3192 150 -3160
rect 194 -3213 195 -3191
rect 359 -3213 360 -3191
rect 394 -3192 395 -3160
rect 408 -3192 409 -3160
rect 457 -3213 458 -3191
rect 506 -3213 507 -3191
rect 583 -3192 584 -3160
rect 597 -3192 598 -3160
rect 618 -3213 619 -3191
rect 625 -3192 626 -3160
rect 695 -3213 696 -3191
rect 786 -3192 787 -3160
rect 800 -3213 801 -3191
rect 807 -3213 808 -3191
rect 814 -3192 815 -3160
rect 884 -3213 885 -3191
rect 961 -3192 962 -3160
rect 1157 -3213 1158 -3191
rect 1171 -3192 1172 -3160
rect 86 -3213 87 -3193
rect 107 -3194 108 -3160
rect 163 -3194 164 -3160
rect 331 -3213 332 -3193
rect 380 -3194 381 -3160
rect 394 -3213 395 -3193
rect 478 -3194 479 -3160
rect 597 -3213 598 -3193
rect 607 -3213 608 -3193
rect 1010 -3213 1011 -3193
rect 1164 -3213 1165 -3193
rect 1178 -3194 1179 -3160
rect 107 -3213 108 -3195
rect 233 -3196 234 -3160
rect 303 -3213 304 -3195
rect 625 -3213 626 -3195
rect 632 -3196 633 -3160
rect 1003 -3196 1004 -3160
rect 1171 -3213 1172 -3195
rect 1206 -3196 1207 -3160
rect 163 -3213 164 -3197
rect 254 -3198 255 -3160
rect 317 -3198 318 -3160
rect 408 -3213 409 -3197
rect 562 -3198 563 -3160
rect 702 -3213 703 -3197
rect 730 -3198 731 -3160
rect 786 -3213 787 -3197
rect 814 -3213 815 -3197
rect 849 -3198 850 -3160
rect 905 -3213 906 -3197
rect 1111 -3213 1112 -3197
rect 1167 -3213 1168 -3197
rect 1206 -3213 1207 -3197
rect 173 -3213 174 -3199
rect 226 -3213 227 -3199
rect 254 -3213 255 -3199
rect 261 -3200 262 -3160
rect 366 -3200 367 -3160
rect 380 -3213 381 -3199
rect 527 -3200 528 -3160
rect 562 -3213 563 -3199
rect 583 -3213 584 -3199
rect 590 -3200 591 -3160
rect 639 -3200 640 -3160
rect 751 -3213 752 -3199
rect 828 -3200 829 -3160
rect 849 -3213 850 -3199
rect 926 -3213 927 -3199
rect 982 -3200 983 -3160
rect 212 -3202 213 -3160
rect 317 -3213 318 -3201
rect 366 -3213 367 -3201
rect 604 -3202 605 -3160
rect 632 -3213 633 -3201
rect 639 -3213 640 -3201
rect 646 -3213 647 -3201
rect 782 -3202 783 -3160
rect 828 -3213 829 -3201
rect 1003 -3213 1004 -3201
rect 177 -3204 178 -3160
rect 212 -3213 213 -3203
rect 222 -3204 223 -3160
rect 233 -3213 234 -3203
rect 310 -3204 311 -3160
rect 604 -3213 605 -3203
rect 730 -3213 731 -3203
rect 744 -3204 745 -3160
rect 961 -3213 962 -3203
rect 1059 -3213 1060 -3203
rect 240 -3206 241 -3160
rect 310 -3213 311 -3205
rect 450 -3206 451 -3160
rect 527 -3213 528 -3205
rect 555 -3213 556 -3205
rect 590 -3213 591 -3205
rect 744 -3213 745 -3205
rect 758 -3206 759 -3160
rect 240 -3213 241 -3207
rect 275 -3208 276 -3160
rect 289 -3208 290 -3160
rect 450 -3213 451 -3207
rect 478 -3213 479 -3207
rect 982 -3213 983 -3207
rect 247 -3213 248 -3209
rect 289 -3213 290 -3209
rect 758 -3213 759 -3209
rect 765 -3213 766 -3209
rect 261 -3213 262 -3211
rect 275 -3213 276 -3211
rect 58 -3223 59 -3221
rect 247 -3223 248 -3221
rect 250 -3223 251 -3221
rect 250 -3268 251 -3222
rect 250 -3223 251 -3221
rect 250 -3268 251 -3222
rect 317 -3223 318 -3221
rect 317 -3268 318 -3222
rect 317 -3223 318 -3221
rect 317 -3268 318 -3222
rect 338 -3223 339 -3221
rect 341 -3259 342 -3222
rect 359 -3223 360 -3221
rect 362 -3259 363 -3222
rect 380 -3223 381 -3221
rect 397 -3268 398 -3222
rect 408 -3223 409 -3221
rect 663 -3223 664 -3221
rect 702 -3223 703 -3221
rect 758 -3223 759 -3221
rect 782 -3268 783 -3222
rect 1031 -3223 1032 -3221
rect 1038 -3223 1039 -3221
rect 1062 -3223 1063 -3221
rect 1066 -3268 1067 -3222
rect 1080 -3223 1081 -3221
rect 1094 -3223 1095 -3221
rect 1094 -3268 1095 -3222
rect 1094 -3223 1095 -3221
rect 1094 -3268 1095 -3222
rect 1101 -3223 1102 -3221
rect 1111 -3223 1112 -3221
rect 1129 -3223 1130 -3221
rect 1129 -3268 1130 -3222
rect 1129 -3223 1130 -3221
rect 1129 -3268 1130 -3222
rect 1136 -3223 1137 -3221
rect 1157 -3223 1158 -3221
rect 1206 -3223 1207 -3221
rect 1251 -3268 1252 -3222
rect 1290 -3268 1291 -3222
rect 1325 -3268 1326 -3222
rect 1328 -3268 1329 -3222
rect 1332 -3223 1333 -3221
rect 1360 -3223 1361 -3221
rect 1360 -3268 1361 -3222
rect 1360 -3223 1361 -3221
rect 1360 -3268 1361 -3222
rect 1367 -3223 1368 -3221
rect 1367 -3268 1368 -3222
rect 1367 -3223 1368 -3221
rect 1367 -3268 1368 -3222
rect 1409 -3223 1410 -3221
rect 1409 -3268 1410 -3222
rect 1409 -3223 1410 -3221
rect 1409 -3268 1410 -3222
rect 1451 -3223 1452 -3221
rect 1454 -3223 1455 -3221
rect 1465 -3223 1466 -3221
rect 1465 -3268 1466 -3222
rect 1465 -3223 1466 -3221
rect 1465 -3268 1466 -3222
rect 65 -3225 66 -3221
rect 261 -3225 262 -3221
rect 338 -3268 339 -3224
rect 359 -3268 360 -3224
rect 443 -3225 444 -3221
rect 464 -3225 465 -3221
rect 579 -3225 580 -3221
rect 604 -3225 605 -3221
rect 919 -3225 920 -3221
rect 982 -3225 983 -3221
rect 1216 -3268 1217 -3224
rect 1234 -3225 1235 -3221
rect 1234 -3268 1235 -3224
rect 1234 -3225 1235 -3221
rect 1234 -3268 1235 -3224
rect 1451 -3268 1452 -3224
rect 1458 -3225 1459 -3221
rect 72 -3227 73 -3221
rect 117 -3227 118 -3221
rect 121 -3227 122 -3221
rect 324 -3227 325 -3221
rect 380 -3268 381 -3226
rect 415 -3227 416 -3221
rect 429 -3227 430 -3221
rect 488 -3268 489 -3226
rect 499 -3227 500 -3221
rect 499 -3268 500 -3226
rect 499 -3227 500 -3221
rect 499 -3268 500 -3226
rect 520 -3227 521 -3221
rect 520 -3268 521 -3226
rect 520 -3227 521 -3221
rect 520 -3268 521 -3226
rect 534 -3227 535 -3221
rect 537 -3227 538 -3221
rect 548 -3227 549 -3221
rect 726 -3268 727 -3226
rect 737 -3227 738 -3221
rect 863 -3227 864 -3221
rect 866 -3227 867 -3221
rect 933 -3227 934 -3221
rect 982 -3268 983 -3226
rect 989 -3227 990 -3221
rect 992 -3268 993 -3226
rect 1045 -3227 1046 -3221
rect 1052 -3227 1053 -3221
rect 1101 -3268 1102 -3226
rect 1125 -3268 1126 -3226
rect 1136 -3268 1137 -3226
rect 1143 -3227 1144 -3221
rect 1143 -3268 1144 -3226
rect 1143 -3227 1144 -3221
rect 1143 -3268 1144 -3226
rect 1150 -3227 1151 -3221
rect 1188 -3268 1189 -3226
rect 1213 -3227 1214 -3221
rect 1220 -3268 1221 -3226
rect 79 -3229 80 -3221
rect 173 -3229 174 -3221
rect 177 -3268 178 -3228
rect 191 -3229 192 -3221
rect 201 -3229 202 -3221
rect 387 -3229 388 -3221
rect 422 -3229 423 -3221
rect 429 -3268 430 -3228
rect 443 -3268 444 -3228
rect 457 -3229 458 -3221
rect 534 -3268 535 -3228
rect 646 -3229 647 -3221
rect 730 -3229 731 -3221
rect 737 -3268 738 -3228
rect 758 -3268 759 -3228
rect 765 -3229 766 -3221
rect 786 -3229 787 -3221
rect 1003 -3229 1004 -3221
rect 1017 -3229 1018 -3221
rect 1167 -3229 1168 -3221
rect 1185 -3229 1186 -3221
rect 1206 -3268 1207 -3228
rect 86 -3231 87 -3221
rect 128 -3231 129 -3221
rect 131 -3231 132 -3221
rect 324 -3268 325 -3230
rect 352 -3231 353 -3221
rect 415 -3268 416 -3230
rect 450 -3231 451 -3221
rect 457 -3268 458 -3230
rect 541 -3231 542 -3221
rect 646 -3268 647 -3230
rect 733 -3268 734 -3230
rect 786 -3268 787 -3230
rect 849 -3231 850 -3221
rect 985 -3231 986 -3221
rect 996 -3231 997 -3221
rect 1108 -3231 1109 -3221
rect 1150 -3268 1151 -3230
rect 1171 -3231 1172 -3221
rect 1185 -3268 1186 -3230
rect 1199 -3231 1200 -3221
rect 93 -3233 94 -3221
rect 180 -3233 181 -3221
rect 187 -3268 188 -3232
rect 366 -3233 367 -3221
rect 387 -3268 388 -3232
rect 401 -3233 402 -3221
rect 450 -3268 451 -3232
rect 471 -3233 472 -3221
rect 548 -3268 549 -3232
rect 597 -3233 598 -3221
rect 604 -3268 605 -3232
rect 632 -3233 633 -3221
rect 639 -3233 640 -3221
rect 702 -3268 703 -3232
rect 765 -3268 766 -3232
rect 828 -3233 829 -3221
rect 880 -3268 881 -3232
rect 926 -3233 927 -3221
rect 933 -3268 934 -3232
rect 968 -3233 969 -3221
rect 996 -3268 997 -3232
rect 1164 -3233 1165 -3221
rect 100 -3235 101 -3221
rect 243 -3268 244 -3234
rect 247 -3268 248 -3234
rect 275 -3235 276 -3221
rect 282 -3235 283 -3221
rect 352 -3268 353 -3234
rect 366 -3268 367 -3234
rect 404 -3268 405 -3234
rect 474 -3268 475 -3234
rect 597 -3268 598 -3234
rect 611 -3235 612 -3221
rect 639 -3268 640 -3234
rect 807 -3235 808 -3221
rect 828 -3268 829 -3234
rect 898 -3235 899 -3221
rect 926 -3268 927 -3234
rect 940 -3235 941 -3221
rect 1003 -3268 1004 -3234
rect 1059 -3235 1060 -3221
rect 1122 -3235 1123 -3221
rect 1160 -3268 1161 -3234
rect 1171 -3268 1172 -3234
rect 114 -3237 115 -3221
rect 492 -3237 493 -3221
rect 555 -3237 556 -3221
rect 891 -3237 892 -3221
rect 898 -3268 899 -3236
rect 912 -3237 913 -3221
rect 919 -3268 920 -3236
rect 1122 -3268 1123 -3236
rect 1164 -3268 1165 -3236
rect 1192 -3237 1193 -3221
rect 135 -3239 136 -3221
rect 170 -3268 171 -3238
rect 191 -3268 192 -3238
rect 401 -3268 402 -3238
rect 555 -3268 556 -3238
rect 562 -3239 563 -3221
rect 569 -3239 570 -3221
rect 576 -3239 577 -3221
rect 611 -3268 612 -3238
rect 653 -3239 654 -3221
rect 800 -3239 801 -3221
rect 807 -3268 808 -3238
rect 856 -3239 857 -3221
rect 891 -3268 892 -3238
rect 940 -3268 941 -3238
rect 954 -3239 955 -3221
rect 1073 -3239 1074 -3221
rect 1073 -3268 1074 -3238
rect 1073 -3239 1074 -3221
rect 1073 -3268 1074 -3238
rect 1080 -3268 1081 -3238
rect 1115 -3239 1116 -3221
rect 149 -3241 150 -3221
rect 464 -3268 465 -3240
rect 527 -3241 528 -3221
rect 569 -3268 570 -3240
rect 618 -3241 619 -3221
rect 625 -3268 626 -3240
rect 628 -3241 629 -3221
rect 744 -3241 745 -3221
rect 793 -3241 794 -3221
rect 800 -3268 801 -3240
rect 884 -3241 885 -3221
rect 912 -3268 913 -3240
rect 947 -3241 948 -3221
rect 954 -3268 955 -3240
rect 1087 -3241 1088 -3221
rect 1108 -3268 1109 -3240
rect 152 -3243 153 -3221
rect 576 -3268 577 -3242
rect 618 -3268 619 -3242
rect 635 -3243 636 -3221
rect 653 -3268 654 -3242
rect 688 -3243 689 -3221
rect 744 -3268 745 -3242
rect 751 -3243 752 -3221
rect 793 -3268 794 -3242
rect 821 -3243 822 -3221
rect 842 -3243 843 -3221
rect 947 -3268 948 -3242
rect 226 -3245 227 -3221
rect 229 -3259 230 -3244
rect 264 -3245 265 -3221
rect 275 -3268 276 -3244
rect 296 -3245 297 -3221
rect 422 -3268 423 -3244
rect 513 -3245 514 -3221
rect 527 -3268 528 -3244
rect 558 -3245 559 -3221
rect 674 -3245 675 -3221
rect 751 -3268 752 -3244
rect 779 -3245 780 -3221
rect 821 -3268 822 -3244
rect 961 -3245 962 -3221
rect 107 -3247 108 -3221
rect 264 -3268 265 -3246
rect 268 -3247 269 -3221
rect 282 -3268 283 -3246
rect 296 -3268 297 -3246
rect 303 -3247 304 -3221
rect 394 -3247 395 -3221
rect 632 -3268 633 -3246
rect 635 -3268 636 -3246
rect 772 -3247 773 -3221
rect 842 -3268 843 -3246
rect 870 -3247 871 -3221
rect 884 -3268 885 -3246
rect 905 -3247 906 -3221
rect 961 -3268 962 -3246
rect 1024 -3247 1025 -3221
rect 156 -3249 157 -3221
rect 394 -3268 395 -3248
rect 506 -3249 507 -3221
rect 513 -3268 514 -3248
rect 562 -3268 563 -3248
rect 583 -3249 584 -3221
rect 660 -3249 661 -3221
rect 688 -3268 689 -3248
rect 772 -3268 773 -3248
rect 814 -3249 815 -3221
rect 870 -3268 871 -3248
rect 877 -3249 878 -3221
rect 905 -3268 906 -3248
rect 975 -3249 976 -3221
rect 156 -3268 157 -3250
rect 261 -3268 262 -3250
rect 268 -3268 269 -3250
rect 289 -3251 290 -3221
rect 436 -3251 437 -3221
rect 583 -3268 584 -3250
rect 660 -3268 661 -3250
rect 695 -3251 696 -3221
rect 877 -3268 878 -3250
rect 1010 -3251 1011 -3221
rect 198 -3253 199 -3221
rect 289 -3268 290 -3252
rect 373 -3253 374 -3221
rect 436 -3268 437 -3252
rect 506 -3268 507 -3252
rect 607 -3253 608 -3221
rect 667 -3253 668 -3221
rect 814 -3268 815 -3252
rect 184 -3255 185 -3221
rect 198 -3268 199 -3254
rect 219 -3255 220 -3221
rect 303 -3268 304 -3254
rect 331 -3255 332 -3221
rect 373 -3268 374 -3254
rect 590 -3255 591 -3221
rect 695 -3268 696 -3254
rect 212 -3257 213 -3221
rect 219 -3268 220 -3256
rect 226 -3268 227 -3256
rect 310 -3257 311 -3221
rect 331 -3268 332 -3256
rect 667 -3268 668 -3256
rect 716 -3257 717 -3221
rect 212 -3268 213 -3258
rect 233 -3259 234 -3221
rect 310 -3268 311 -3258
rect 478 -3259 479 -3221
rect 674 -3268 675 -3258
rect 681 -3259 682 -3221
rect 709 -3259 710 -3221
rect 716 -3268 717 -3258
rect 1454 -3268 1455 -3258
rect 1458 -3268 1459 -3258
rect 163 -3261 164 -3221
rect 233 -3268 234 -3260
rect 478 -3268 479 -3260
rect 485 -3261 486 -3221
rect 681 -3268 682 -3260
rect 723 -3261 724 -3221
rect 163 -3268 164 -3262
rect 208 -3263 209 -3221
rect 408 -3268 409 -3262
rect 485 -3268 486 -3262
rect 709 -3268 710 -3262
rect 835 -3263 836 -3221
rect 208 -3268 209 -3264
rect 240 -3265 241 -3221
rect 240 -3268 241 -3266
rect 492 -3268 493 -3266
rect 163 -3278 164 -3276
rect 229 -3331 230 -3277
rect 243 -3278 244 -3276
rect 534 -3278 535 -3276
rect 593 -3278 594 -3276
rect 646 -3278 647 -3276
rect 670 -3331 671 -3277
rect 674 -3278 675 -3276
rect 684 -3331 685 -3277
rect 702 -3278 703 -3276
rect 723 -3278 724 -3276
rect 919 -3278 920 -3276
rect 936 -3331 937 -3277
rect 940 -3278 941 -3276
rect 947 -3278 948 -3276
rect 975 -3331 976 -3277
rect 982 -3278 983 -3276
rect 989 -3331 990 -3277
rect 1003 -3278 1004 -3276
rect 1059 -3331 1060 -3277
rect 1066 -3278 1067 -3276
rect 1066 -3331 1067 -3277
rect 1066 -3278 1067 -3276
rect 1066 -3331 1067 -3277
rect 1073 -3278 1074 -3276
rect 1076 -3282 1077 -3277
rect 1094 -3278 1095 -3276
rect 1094 -3331 1095 -3277
rect 1094 -3278 1095 -3276
rect 1094 -3331 1095 -3277
rect 1108 -3278 1109 -3276
rect 1115 -3331 1116 -3277
rect 1122 -3278 1123 -3276
rect 1129 -3278 1130 -3276
rect 1136 -3278 1137 -3276
rect 1157 -3278 1158 -3276
rect 1171 -3278 1172 -3276
rect 1185 -3278 1186 -3276
rect 1206 -3278 1207 -3276
rect 1213 -3331 1214 -3277
rect 1216 -3278 1217 -3276
rect 1220 -3278 1221 -3276
rect 1251 -3278 1252 -3276
rect 1290 -3278 1291 -3276
rect 1360 -3278 1361 -3276
rect 1360 -3331 1361 -3277
rect 1360 -3278 1361 -3276
rect 1360 -3331 1361 -3277
rect 1367 -3278 1368 -3276
rect 1367 -3331 1368 -3277
rect 1367 -3278 1368 -3276
rect 1367 -3331 1368 -3277
rect 1409 -3278 1410 -3276
rect 1409 -3331 1410 -3277
rect 1409 -3278 1410 -3276
rect 1409 -3331 1410 -3277
rect 1451 -3278 1452 -3276
rect 1461 -3278 1462 -3276
rect 177 -3280 178 -3276
rect 205 -3331 206 -3279
rect 208 -3280 209 -3276
rect 240 -3331 241 -3279
rect 289 -3280 290 -3276
rect 411 -3331 412 -3279
rect 415 -3280 416 -3276
rect 646 -3331 647 -3279
rect 688 -3280 689 -3276
rect 702 -3331 703 -3279
rect 730 -3280 731 -3276
rect 751 -3280 752 -3276
rect 779 -3280 780 -3276
rect 800 -3280 801 -3276
rect 807 -3280 808 -3276
rect 835 -3331 836 -3279
rect 838 -3331 839 -3279
rect 996 -3280 997 -3276
rect 1073 -3331 1074 -3279
rect 1080 -3280 1081 -3276
rect 1097 -3331 1098 -3279
rect 1290 -3331 1291 -3279
rect 1458 -3280 1459 -3276
rect 1465 -3280 1466 -3276
rect 177 -3331 178 -3281
rect 268 -3282 269 -3276
rect 282 -3282 283 -3276
rect 289 -3331 290 -3281
rect 331 -3282 332 -3276
rect 383 -3331 384 -3281
rect 394 -3282 395 -3276
rect 618 -3282 619 -3276
rect 639 -3282 640 -3276
rect 674 -3331 675 -3281
rect 681 -3282 682 -3276
rect 688 -3331 689 -3281
rect 751 -3331 752 -3281
rect 758 -3282 759 -3276
rect 779 -3331 780 -3281
rect 786 -3282 787 -3276
rect 793 -3282 794 -3276
rect 800 -3331 801 -3281
rect 814 -3282 815 -3276
rect 849 -3331 850 -3281
rect 856 -3331 857 -3281
rect 877 -3282 878 -3276
rect 912 -3282 913 -3276
rect 919 -3331 920 -3281
rect 940 -3331 941 -3281
rect 954 -3282 955 -3276
rect 1080 -3331 1081 -3281
rect 1101 -3282 1102 -3276
rect 1108 -3331 1109 -3281
rect 1125 -3282 1126 -3276
rect 1164 -3282 1165 -3276
rect 184 -3284 185 -3276
rect 191 -3284 192 -3276
rect 212 -3284 213 -3276
rect 212 -3331 213 -3283
rect 212 -3284 213 -3276
rect 212 -3331 213 -3283
rect 226 -3284 227 -3276
rect 247 -3331 248 -3283
rect 282 -3331 283 -3283
rect 296 -3284 297 -3276
rect 324 -3284 325 -3276
rect 394 -3331 395 -3283
rect 415 -3331 416 -3283
rect 429 -3284 430 -3276
rect 457 -3284 458 -3276
rect 590 -3284 591 -3276
rect 593 -3331 594 -3283
rect 709 -3284 710 -3276
rect 712 -3331 713 -3283
rect 814 -3331 815 -3283
rect 828 -3284 829 -3276
rect 828 -3331 829 -3283
rect 828 -3284 829 -3276
rect 828 -3331 829 -3283
rect 863 -3331 864 -3283
rect 884 -3284 885 -3276
rect 912 -3331 913 -3283
rect 933 -3284 934 -3276
rect 954 -3331 955 -3283
rect 961 -3284 962 -3276
rect 1136 -3331 1137 -3283
rect 1150 -3284 1151 -3276
rect 156 -3286 157 -3276
rect 191 -3331 192 -3285
rect 226 -3331 227 -3285
rect 618 -3331 619 -3285
rect 639 -3331 640 -3285
rect 660 -3286 661 -3276
rect 681 -3331 682 -3285
rect 807 -3331 808 -3285
rect 870 -3286 871 -3276
rect 884 -3331 885 -3285
rect 926 -3286 927 -3276
rect 961 -3331 962 -3285
rect 1143 -3286 1144 -3276
rect 1143 -3331 1144 -3285
rect 1143 -3286 1144 -3276
rect 1143 -3331 1144 -3285
rect 184 -3331 185 -3287
rect 198 -3288 199 -3276
rect 296 -3331 297 -3287
rect 572 -3331 573 -3287
rect 576 -3288 577 -3276
rect 933 -3331 934 -3287
rect 187 -3290 188 -3276
rect 268 -3331 269 -3289
rect 331 -3331 332 -3289
rect 345 -3290 346 -3276
rect 359 -3290 360 -3276
rect 359 -3331 360 -3289
rect 359 -3290 360 -3276
rect 359 -3331 360 -3289
rect 366 -3290 367 -3276
rect 590 -3331 591 -3289
rect 597 -3290 598 -3276
rect 723 -3331 724 -3289
rect 744 -3290 745 -3276
rect 786 -3331 787 -3289
rect 793 -3331 794 -3289
rect 821 -3290 822 -3276
rect 877 -3331 878 -3289
rect 898 -3290 899 -3276
rect 198 -3331 199 -3291
rect 219 -3292 220 -3276
rect 338 -3292 339 -3276
rect 345 -3331 346 -3291
rect 366 -3331 367 -3291
rect 387 -3292 388 -3276
rect 422 -3292 423 -3276
rect 457 -3331 458 -3291
rect 471 -3331 472 -3291
rect 478 -3292 479 -3276
rect 488 -3292 489 -3276
rect 583 -3292 584 -3276
rect 611 -3292 612 -3276
rect 611 -3331 612 -3291
rect 611 -3292 612 -3276
rect 611 -3331 612 -3291
rect 635 -3292 636 -3276
rect 870 -3331 871 -3291
rect 891 -3292 892 -3276
rect 926 -3331 927 -3291
rect 170 -3294 171 -3276
rect 338 -3331 339 -3293
rect 373 -3294 374 -3276
rect 429 -3331 430 -3293
rect 446 -3331 447 -3293
rect 744 -3331 745 -3293
rect 758 -3331 759 -3293
rect 765 -3294 766 -3276
rect 821 -3331 822 -3293
rect 842 -3294 843 -3276
rect 898 -3331 899 -3293
rect 905 -3294 906 -3276
rect 219 -3331 220 -3295
rect 233 -3296 234 -3276
rect 275 -3296 276 -3276
rect 387 -3331 388 -3295
rect 422 -3331 423 -3295
rect 506 -3296 507 -3276
rect 534 -3331 535 -3295
rect 541 -3296 542 -3276
rect 555 -3296 556 -3276
rect 597 -3331 598 -3295
rect 660 -3331 661 -3295
rect 716 -3296 717 -3276
rect 765 -3331 766 -3295
rect 772 -3296 773 -3276
rect 842 -3331 843 -3295
rect 845 -3331 846 -3295
rect 880 -3296 881 -3276
rect 905 -3331 906 -3295
rect 233 -3331 234 -3297
rect 408 -3298 409 -3276
rect 464 -3298 465 -3276
rect 555 -3331 556 -3297
rect 576 -3331 577 -3297
rect 709 -3331 710 -3297
rect 716 -3331 717 -3297
rect 737 -3298 738 -3276
rect 254 -3300 255 -3276
rect 275 -3331 276 -3299
rect 317 -3300 318 -3276
rect 373 -3331 374 -3299
rect 464 -3331 465 -3299
rect 604 -3300 605 -3276
rect 695 -3300 696 -3276
rect 772 -3331 773 -3299
rect 254 -3331 255 -3301
rect 352 -3302 353 -3276
rect 401 -3302 402 -3276
rect 695 -3331 696 -3301
rect 737 -3331 738 -3301
rect 891 -3331 892 -3301
rect 310 -3304 311 -3276
rect 317 -3331 318 -3303
rect 352 -3331 353 -3303
rect 485 -3304 486 -3276
rect 492 -3304 493 -3276
rect 541 -3331 542 -3303
rect 583 -3331 584 -3303
rect 632 -3304 633 -3276
rect 303 -3306 304 -3276
rect 310 -3331 311 -3305
rect 380 -3306 381 -3276
rect 485 -3331 486 -3305
rect 604 -3331 605 -3305
rect 782 -3306 783 -3276
rect 303 -3331 304 -3307
rect 992 -3308 993 -3276
rect 380 -3331 381 -3309
rect 730 -3331 731 -3309
rect 401 -3331 402 -3311
rect 450 -3312 451 -3276
rect 467 -3331 468 -3311
rect 632 -3331 633 -3311
rect 436 -3314 437 -3276
rect 492 -3331 493 -3313
rect 436 -3331 437 -3315
rect 443 -3316 444 -3276
rect 450 -3331 451 -3315
rect 625 -3316 626 -3276
rect 324 -3331 325 -3317
rect 443 -3331 444 -3317
rect 474 -3318 475 -3276
rect 513 -3318 514 -3276
rect 625 -3331 626 -3317
rect 653 -3318 654 -3276
rect 478 -3331 479 -3319
rect 499 -3320 500 -3276
rect 513 -3331 514 -3319
rect 667 -3320 668 -3276
rect 499 -3331 500 -3321
rect 520 -3322 521 -3276
rect 548 -3322 549 -3276
rect 653 -3331 654 -3321
rect 506 -3331 507 -3323
rect 667 -3331 668 -3323
rect 520 -3331 521 -3325
rect 527 -3326 528 -3276
rect 548 -3331 549 -3325
rect 562 -3326 563 -3276
rect 408 -3331 409 -3327
rect 562 -3331 563 -3327
rect 527 -3331 528 -3329
rect 569 -3330 570 -3276
rect 184 -3341 185 -3339
rect 184 -3396 185 -3340
rect 184 -3341 185 -3339
rect 184 -3396 185 -3340
rect 191 -3341 192 -3339
rect 194 -3369 195 -3340
rect 261 -3341 262 -3339
rect 618 -3341 619 -3339
rect 621 -3341 622 -3339
rect 786 -3341 787 -3339
rect 807 -3341 808 -3339
rect 866 -3396 867 -3340
rect 870 -3341 871 -3339
rect 1097 -3341 1098 -3339
rect 1115 -3341 1116 -3339
rect 1122 -3396 1123 -3340
rect 1139 -3341 1140 -3339
rect 1143 -3341 1144 -3339
rect 1213 -3341 1214 -3339
rect 1213 -3396 1214 -3340
rect 1213 -3341 1214 -3339
rect 1213 -3396 1214 -3340
rect 1353 -3396 1354 -3340
rect 1367 -3341 1368 -3339
rect 1409 -3341 1410 -3339
rect 1409 -3396 1410 -3340
rect 1409 -3341 1410 -3339
rect 1409 -3396 1410 -3340
rect 191 -3396 192 -3342
rect 240 -3343 241 -3339
rect 261 -3396 262 -3342
rect 264 -3343 265 -3339
rect 275 -3343 276 -3339
rect 282 -3343 283 -3339
rect 411 -3343 412 -3339
rect 429 -3343 430 -3339
rect 429 -3396 430 -3342
rect 429 -3343 430 -3339
rect 429 -3396 430 -3342
rect 471 -3343 472 -3339
rect 569 -3343 570 -3339
rect 576 -3343 577 -3339
rect 590 -3396 591 -3342
rect 604 -3343 605 -3339
rect 618 -3396 619 -3342
rect 695 -3343 696 -3339
rect 695 -3396 696 -3342
rect 695 -3343 696 -3339
rect 695 -3396 696 -3342
rect 702 -3343 703 -3339
rect 702 -3396 703 -3342
rect 702 -3343 703 -3339
rect 702 -3396 703 -3342
rect 709 -3343 710 -3339
rect 740 -3343 741 -3339
rect 779 -3343 780 -3339
rect 779 -3396 780 -3342
rect 779 -3343 780 -3339
rect 779 -3396 780 -3342
rect 821 -3343 822 -3339
rect 835 -3396 836 -3342
rect 842 -3343 843 -3339
rect 884 -3343 885 -3339
rect 894 -3396 895 -3342
rect 926 -3343 927 -3339
rect 940 -3343 941 -3339
rect 940 -3396 941 -3342
rect 940 -3343 941 -3339
rect 940 -3396 941 -3342
rect 947 -3343 948 -3339
rect 961 -3343 962 -3339
rect 975 -3343 976 -3339
rect 996 -3396 997 -3342
rect 1059 -3343 1060 -3339
rect 1073 -3343 1074 -3339
rect 1108 -3343 1109 -3339
rect 1115 -3396 1116 -3342
rect 1290 -3343 1291 -3339
rect 1367 -3396 1368 -3342
rect 198 -3345 199 -3339
rect 240 -3396 241 -3344
rect 254 -3345 255 -3339
rect 275 -3396 276 -3344
rect 282 -3396 283 -3344
rect 289 -3345 290 -3339
rect 303 -3345 304 -3339
rect 306 -3345 307 -3339
rect 338 -3345 339 -3339
rect 464 -3396 465 -3344
rect 471 -3396 472 -3344
rect 520 -3345 521 -3339
rect 541 -3396 542 -3344
rect 933 -3345 934 -3339
rect 989 -3345 990 -3339
rect 989 -3396 990 -3344
rect 989 -3345 990 -3339
rect 989 -3396 990 -3344
rect 1062 -3345 1063 -3339
rect 1066 -3345 1067 -3339
rect 1073 -3396 1074 -3344
rect 1080 -3345 1081 -3339
rect 1360 -3345 1361 -3339
rect 1360 -3396 1361 -3344
rect 1360 -3345 1361 -3339
rect 1360 -3396 1361 -3344
rect 198 -3396 199 -3346
rect 352 -3347 353 -3339
rect 355 -3396 356 -3346
rect 506 -3347 507 -3339
rect 513 -3347 514 -3339
rect 513 -3396 514 -3346
rect 513 -3347 514 -3339
rect 513 -3396 514 -3346
rect 520 -3396 521 -3346
rect 527 -3347 528 -3339
rect 558 -3396 559 -3346
rect 569 -3396 570 -3346
rect 604 -3396 605 -3346
rect 646 -3347 647 -3339
rect 660 -3347 661 -3339
rect 709 -3396 710 -3346
rect 712 -3347 713 -3339
rect 793 -3347 794 -3339
rect 828 -3347 829 -3339
rect 831 -3396 832 -3346
rect 849 -3347 850 -3339
rect 849 -3396 850 -3346
rect 849 -3347 850 -3339
rect 849 -3396 850 -3346
rect 856 -3347 857 -3339
rect 856 -3396 857 -3346
rect 856 -3347 857 -3339
rect 856 -3396 857 -3346
rect 870 -3396 871 -3346
rect 905 -3347 906 -3339
rect 919 -3347 920 -3339
rect 919 -3396 920 -3346
rect 919 -3347 920 -3339
rect 919 -3396 920 -3346
rect 926 -3396 927 -3346
rect 954 -3347 955 -3339
rect 226 -3396 227 -3348
rect 646 -3396 647 -3348
rect 737 -3349 738 -3339
rect 800 -3349 801 -3339
rect 884 -3396 885 -3348
rect 891 -3349 892 -3339
rect 905 -3396 906 -3348
rect 912 -3349 913 -3339
rect 247 -3351 248 -3339
rect 254 -3396 255 -3350
rect 268 -3351 269 -3339
rect 443 -3351 444 -3339
rect 492 -3351 493 -3339
rect 544 -3351 545 -3339
rect 555 -3351 556 -3339
rect 660 -3396 661 -3350
rect 737 -3396 738 -3350
rect 758 -3351 759 -3339
rect 775 -3396 776 -3350
rect 821 -3396 822 -3350
rect 877 -3351 878 -3339
rect 912 -3396 913 -3350
rect 212 -3353 213 -3339
rect 268 -3396 269 -3352
rect 289 -3396 290 -3352
rect 317 -3353 318 -3339
rect 366 -3353 367 -3339
rect 380 -3396 381 -3352
rect 383 -3353 384 -3339
rect 387 -3353 388 -3339
rect 394 -3353 395 -3339
rect 467 -3353 468 -3339
rect 495 -3396 496 -3352
rect 527 -3396 528 -3352
rect 744 -3353 745 -3339
rect 828 -3396 829 -3352
rect 863 -3353 864 -3339
rect 877 -3396 878 -3352
rect 177 -3355 178 -3339
rect 394 -3396 395 -3354
rect 397 -3396 398 -3354
rect 681 -3355 682 -3339
rect 744 -3396 745 -3354
rect 772 -3355 773 -3339
rect 863 -3396 864 -3354
rect 898 -3355 899 -3339
rect 177 -3396 178 -3356
rect 229 -3396 230 -3356
rect 296 -3357 297 -3339
rect 366 -3396 367 -3356
rect 373 -3357 374 -3339
rect 387 -3396 388 -3356
rect 443 -3396 444 -3356
rect 572 -3357 573 -3339
rect 576 -3396 577 -3356
rect 681 -3396 682 -3356
rect 758 -3396 759 -3356
rect 765 -3357 766 -3339
rect 205 -3359 206 -3339
rect 212 -3396 213 -3358
rect 219 -3359 220 -3339
rect 247 -3396 248 -3358
rect 296 -3396 297 -3358
rect 359 -3359 360 -3339
rect 373 -3396 374 -3358
rect 457 -3359 458 -3339
rect 499 -3359 500 -3339
rect 593 -3359 594 -3339
rect 751 -3359 752 -3339
rect 765 -3396 766 -3358
rect 205 -3396 206 -3360
rect 324 -3361 325 -3339
rect 359 -3396 360 -3360
rect 488 -3396 489 -3360
rect 499 -3396 500 -3360
rect 562 -3361 563 -3339
rect 730 -3361 731 -3339
rect 751 -3396 752 -3360
rect 219 -3396 220 -3362
rect 331 -3363 332 -3339
rect 415 -3363 416 -3339
rect 457 -3396 458 -3362
rect 716 -3363 717 -3339
rect 730 -3396 731 -3362
rect 303 -3396 304 -3364
rect 310 -3365 311 -3339
rect 317 -3396 318 -3364
rect 408 -3365 409 -3339
rect 450 -3365 451 -3339
rect 562 -3396 563 -3364
rect 639 -3365 640 -3339
rect 716 -3396 717 -3364
rect 310 -3396 311 -3366
rect 422 -3367 423 -3339
rect 450 -3396 451 -3366
rect 478 -3367 479 -3339
rect 639 -3396 640 -3366
rect 674 -3367 675 -3339
rect 306 -3396 307 -3368
rect 422 -3396 423 -3368
rect 478 -3396 479 -3368
rect 534 -3369 535 -3339
rect 667 -3369 668 -3339
rect 674 -3396 675 -3368
rect 324 -3396 325 -3370
rect 345 -3371 346 -3339
rect 352 -3396 353 -3370
rect 415 -3396 416 -3370
rect 625 -3371 626 -3339
rect 667 -3396 668 -3370
rect 331 -3396 332 -3372
rect 436 -3373 437 -3339
rect 611 -3373 612 -3339
rect 625 -3396 626 -3372
rect 345 -3396 346 -3374
rect 537 -3396 538 -3374
rect 611 -3396 612 -3374
rect 723 -3375 724 -3339
rect 401 -3377 402 -3339
rect 436 -3396 437 -3376
rect 723 -3396 724 -3376
rect 845 -3377 846 -3339
rect 401 -3396 402 -3378
rect 534 -3396 535 -3378
rect 814 -3379 815 -3339
rect 845 -3396 846 -3378
rect 408 -3396 409 -3380
rect 485 -3381 486 -3339
rect 814 -3396 815 -3380
rect 936 -3381 937 -3339
rect 485 -3396 486 -3382
rect 653 -3383 654 -3339
rect 653 -3396 654 -3384
rect 688 -3385 689 -3339
rect 583 -3387 584 -3339
rect 688 -3396 689 -3386
rect 583 -3396 584 -3388
rect 632 -3389 633 -3339
rect 548 -3391 549 -3339
rect 632 -3396 633 -3390
rect 548 -3396 549 -3392
rect 597 -3393 598 -3339
rect 446 -3395 447 -3339
rect 597 -3396 598 -3394
rect 177 -3406 178 -3404
rect 226 -3406 227 -3404
rect 247 -3406 248 -3404
rect 355 -3406 356 -3404
rect 366 -3406 367 -3404
rect 383 -3406 384 -3404
rect 443 -3406 444 -3404
rect 443 -3439 444 -3405
rect 443 -3406 444 -3404
rect 443 -3439 444 -3405
rect 457 -3406 458 -3404
rect 495 -3406 496 -3404
rect 499 -3406 500 -3404
rect 506 -3406 507 -3404
rect 513 -3406 514 -3404
rect 576 -3406 577 -3404
rect 632 -3406 633 -3404
rect 635 -3422 636 -3405
rect 674 -3406 675 -3404
rect 674 -3439 675 -3405
rect 674 -3406 675 -3404
rect 674 -3439 675 -3405
rect 695 -3406 696 -3404
rect 702 -3439 703 -3405
rect 709 -3406 710 -3404
rect 709 -3439 710 -3405
rect 709 -3406 710 -3404
rect 709 -3439 710 -3405
rect 719 -3439 720 -3405
rect 737 -3406 738 -3404
rect 744 -3406 745 -3404
rect 744 -3439 745 -3405
rect 744 -3406 745 -3404
rect 744 -3439 745 -3405
rect 751 -3406 752 -3404
rect 751 -3439 752 -3405
rect 751 -3406 752 -3404
rect 751 -3439 752 -3405
rect 765 -3406 766 -3404
rect 772 -3406 773 -3404
rect 782 -3439 783 -3405
rect 982 -3439 983 -3405
rect 989 -3406 990 -3404
rect 989 -3439 990 -3405
rect 989 -3406 990 -3404
rect 989 -3439 990 -3405
rect 996 -3406 997 -3404
rect 996 -3439 997 -3405
rect 996 -3406 997 -3404
rect 996 -3439 997 -3405
rect 1073 -3406 1074 -3404
rect 1073 -3439 1074 -3405
rect 1073 -3406 1074 -3404
rect 1073 -3439 1074 -3405
rect 1115 -3406 1116 -3404
rect 1115 -3439 1116 -3405
rect 1115 -3406 1116 -3404
rect 1115 -3439 1116 -3405
rect 1122 -3406 1123 -3404
rect 1122 -3439 1123 -3405
rect 1122 -3406 1123 -3404
rect 1122 -3439 1123 -3405
rect 1213 -3406 1214 -3404
rect 1213 -3439 1214 -3405
rect 1213 -3406 1214 -3404
rect 1213 -3439 1214 -3405
rect 1353 -3406 1354 -3404
rect 1353 -3439 1354 -3405
rect 1353 -3406 1354 -3404
rect 1353 -3439 1354 -3405
rect 1360 -3406 1361 -3404
rect 1360 -3439 1361 -3405
rect 1360 -3406 1361 -3404
rect 1360 -3439 1361 -3405
rect 1367 -3406 1368 -3404
rect 1395 -3439 1396 -3405
rect 1409 -3406 1410 -3404
rect 1409 -3439 1410 -3405
rect 1409 -3406 1410 -3404
rect 1409 -3439 1410 -3405
rect 184 -3408 185 -3404
rect 229 -3408 230 -3404
rect 264 -3439 265 -3407
rect 268 -3408 269 -3404
rect 275 -3408 276 -3404
rect 394 -3408 395 -3404
rect 467 -3408 468 -3404
rect 604 -3408 605 -3404
rect 632 -3439 633 -3407
rect 653 -3408 654 -3404
rect 681 -3408 682 -3404
rect 765 -3439 766 -3407
rect 772 -3439 773 -3407
rect 779 -3408 780 -3404
rect 831 -3439 832 -3407
rect 856 -3408 857 -3404
rect 891 -3408 892 -3404
rect 926 -3408 927 -3404
rect 940 -3408 941 -3404
rect 940 -3439 941 -3407
rect 940 -3408 941 -3404
rect 940 -3439 941 -3407
rect 947 -3439 948 -3407
rect 964 -3439 965 -3407
rect 968 -3439 969 -3407
rect 975 -3439 976 -3407
rect 212 -3410 213 -3404
rect 222 -3439 223 -3409
rect 233 -3410 234 -3404
rect 275 -3439 276 -3409
rect 282 -3410 283 -3404
rect 282 -3439 283 -3409
rect 282 -3410 283 -3404
rect 282 -3439 283 -3409
rect 310 -3410 311 -3404
rect 394 -3439 395 -3409
rect 471 -3410 472 -3404
rect 485 -3439 486 -3409
rect 499 -3439 500 -3409
rect 555 -3439 556 -3409
rect 558 -3410 559 -3404
rect 625 -3410 626 -3404
rect 653 -3439 654 -3409
rect 688 -3410 689 -3404
rect 779 -3439 780 -3409
rect 842 -3410 843 -3404
rect 870 -3410 871 -3404
rect 912 -3410 913 -3404
rect 926 -3439 927 -3409
rect 954 -3439 955 -3409
rect 1010 -3439 1011 -3409
rect 254 -3412 255 -3404
rect 310 -3439 311 -3411
rect 317 -3412 318 -3404
rect 338 -3439 339 -3411
rect 341 -3412 342 -3404
rect 387 -3412 388 -3404
rect 408 -3412 409 -3404
rect 471 -3439 472 -3411
rect 478 -3412 479 -3404
rect 492 -3439 493 -3411
rect 520 -3412 521 -3404
rect 541 -3412 542 -3404
rect 569 -3412 570 -3404
rect 576 -3439 577 -3411
rect 625 -3439 626 -3411
rect 639 -3412 640 -3404
rect 660 -3412 661 -3404
rect 681 -3439 682 -3411
rect 688 -3439 689 -3411
rect 723 -3412 724 -3404
rect 730 -3412 731 -3404
rect 733 -3412 734 -3404
rect 842 -3439 843 -3411
rect 845 -3412 846 -3404
rect 849 -3412 850 -3404
rect 849 -3439 850 -3411
rect 849 -3412 850 -3404
rect 849 -3439 850 -3411
rect 856 -3439 857 -3411
rect 884 -3412 885 -3404
rect 905 -3412 906 -3404
rect 912 -3439 913 -3411
rect 919 -3412 920 -3404
rect 919 -3439 920 -3411
rect 919 -3412 920 -3404
rect 919 -3439 920 -3411
rect 961 -3439 962 -3411
rect 1094 -3439 1095 -3411
rect 191 -3414 192 -3404
rect 341 -3439 342 -3413
rect 352 -3439 353 -3413
rect 401 -3414 402 -3404
rect 534 -3414 535 -3404
rect 548 -3414 549 -3404
rect 569 -3439 570 -3413
rect 590 -3414 591 -3404
rect 597 -3414 598 -3404
rect 660 -3439 661 -3413
rect 695 -3439 696 -3413
rect 716 -3414 717 -3404
rect 723 -3439 724 -3413
rect 814 -3414 815 -3404
rect 863 -3414 864 -3404
rect 870 -3439 871 -3413
rect 877 -3414 878 -3404
rect 884 -3439 885 -3413
rect 240 -3416 241 -3404
rect 254 -3439 255 -3415
rect 261 -3416 262 -3404
rect 268 -3439 269 -3415
rect 289 -3416 290 -3404
rect 317 -3439 318 -3415
rect 327 -3439 328 -3415
rect 415 -3416 416 -3404
rect 488 -3416 489 -3404
rect 534 -3439 535 -3415
rect 541 -3439 542 -3415
rect 642 -3439 643 -3415
rect 730 -3439 731 -3415
rect 758 -3416 759 -3404
rect 821 -3416 822 -3404
rect 863 -3439 864 -3415
rect 198 -3418 199 -3404
rect 240 -3439 241 -3417
rect 331 -3418 332 -3404
rect 401 -3439 402 -3417
rect 527 -3418 528 -3404
rect 548 -3439 549 -3417
rect 562 -3418 563 -3404
rect 597 -3439 598 -3417
rect 639 -3439 640 -3417
rect 775 -3418 776 -3404
rect 821 -3439 822 -3417
rect 835 -3418 836 -3404
rect 359 -3420 360 -3404
rect 387 -3439 388 -3419
rect 562 -3439 563 -3419
rect 583 -3420 584 -3404
rect 646 -3420 647 -3404
rect 835 -3439 836 -3419
rect 296 -3422 297 -3404
rect 359 -3439 360 -3421
rect 373 -3422 374 -3404
rect 408 -3439 409 -3421
rect 583 -3439 584 -3421
rect 611 -3422 612 -3404
rect 618 -3422 619 -3404
rect 646 -3439 647 -3421
rect 733 -3439 734 -3421
rect 758 -3439 759 -3421
rect 219 -3424 220 -3404
rect 296 -3439 297 -3423
rect 303 -3424 304 -3404
rect 373 -3439 374 -3423
rect 303 -3439 304 -3425
rect 429 -3426 430 -3404
rect 429 -3439 430 -3427
rect 436 -3428 437 -3404
rect 436 -3439 437 -3429
rect 450 -3430 451 -3404
rect 422 -3432 423 -3404
rect 450 -3439 451 -3431
rect 345 -3434 346 -3404
rect 422 -3439 423 -3433
rect 324 -3436 325 -3404
rect 345 -3439 346 -3435
rect 205 -3438 206 -3404
rect 324 -3439 325 -3437
rect 222 -3449 223 -3447
rect 327 -3449 328 -3447
rect 338 -3466 339 -3448
rect 352 -3449 353 -3447
rect 359 -3449 360 -3447
rect 380 -3466 381 -3448
rect 401 -3449 402 -3447
rect 464 -3466 465 -3448
rect 478 -3466 479 -3448
rect 485 -3449 486 -3447
rect 492 -3449 493 -3447
rect 492 -3466 493 -3448
rect 492 -3449 493 -3447
rect 492 -3466 493 -3448
rect 506 -3466 507 -3448
rect 541 -3449 542 -3447
rect 548 -3449 549 -3447
rect 548 -3466 549 -3448
rect 548 -3449 549 -3447
rect 548 -3466 549 -3448
rect 597 -3449 598 -3447
rect 604 -3466 605 -3448
rect 614 -3466 615 -3448
rect 625 -3449 626 -3447
rect 642 -3449 643 -3447
rect 688 -3449 689 -3447
rect 698 -3466 699 -3448
rect 702 -3449 703 -3447
rect 709 -3449 710 -3447
rect 737 -3449 738 -3447
rect 740 -3449 741 -3447
rect 758 -3449 759 -3447
rect 765 -3449 766 -3447
rect 779 -3449 780 -3447
rect 782 -3449 783 -3447
rect 964 -3449 965 -3447
rect 982 -3449 983 -3447
rect 1066 -3466 1067 -3448
rect 1073 -3449 1074 -3447
rect 1076 -3466 1077 -3448
rect 1094 -3449 1095 -3447
rect 1220 -3466 1221 -3448
rect 1223 -3466 1224 -3448
rect 1227 -3466 1228 -3448
rect 1353 -3449 1354 -3447
rect 1353 -3466 1354 -3448
rect 1353 -3449 1354 -3447
rect 1353 -3466 1354 -3448
rect 1360 -3449 1361 -3447
rect 1360 -3466 1361 -3448
rect 1360 -3449 1361 -3447
rect 1360 -3466 1361 -3448
rect 1409 -3449 1410 -3447
rect 1416 -3466 1417 -3448
rect 254 -3451 255 -3447
rect 261 -3466 262 -3450
rect 264 -3451 265 -3447
rect 460 -3466 461 -3450
rect 471 -3451 472 -3447
rect 485 -3466 486 -3450
rect 520 -3466 521 -3450
rect 572 -3451 573 -3447
rect 621 -3466 622 -3450
rect 723 -3451 724 -3447
rect 737 -3466 738 -3450
rect 751 -3451 752 -3447
rect 821 -3451 822 -3447
rect 828 -3451 829 -3447
rect 831 -3451 832 -3447
rect 849 -3451 850 -3447
rect 856 -3451 857 -3447
rect 856 -3466 857 -3450
rect 856 -3451 857 -3447
rect 856 -3466 857 -3450
rect 884 -3451 885 -3447
rect 884 -3466 885 -3450
rect 884 -3451 885 -3447
rect 884 -3466 885 -3450
rect 912 -3451 913 -3447
rect 912 -3466 913 -3450
rect 912 -3451 913 -3447
rect 912 -3466 913 -3450
rect 919 -3451 920 -3447
rect 919 -3466 920 -3450
rect 919 -3451 920 -3447
rect 919 -3466 920 -3450
rect 926 -3451 927 -3447
rect 926 -3466 927 -3450
rect 926 -3451 927 -3447
rect 926 -3466 927 -3450
rect 933 -3466 934 -3450
rect 954 -3451 955 -3447
rect 957 -3451 958 -3447
rect 968 -3451 969 -3447
rect 989 -3451 990 -3447
rect 989 -3466 990 -3450
rect 989 -3451 990 -3447
rect 989 -3466 990 -3450
rect 996 -3451 997 -3447
rect 996 -3466 997 -3450
rect 996 -3451 997 -3447
rect 996 -3466 997 -3450
rect 1010 -3451 1011 -3447
rect 1073 -3466 1074 -3450
rect 1115 -3451 1116 -3447
rect 1115 -3466 1116 -3450
rect 1115 -3451 1116 -3447
rect 1115 -3466 1116 -3450
rect 1122 -3451 1123 -3447
rect 1122 -3466 1123 -3450
rect 1122 -3451 1123 -3447
rect 1122 -3466 1123 -3450
rect 1213 -3451 1214 -3447
rect 1213 -3466 1214 -3450
rect 1213 -3451 1214 -3447
rect 1213 -3466 1214 -3450
rect 1395 -3451 1396 -3447
rect 1409 -3466 1410 -3450
rect 240 -3453 241 -3447
rect 254 -3466 255 -3452
rect 268 -3453 269 -3447
rect 289 -3453 290 -3447
rect 292 -3453 293 -3447
rect 359 -3466 360 -3452
rect 373 -3453 374 -3447
rect 401 -3466 402 -3452
rect 408 -3453 409 -3447
rect 415 -3466 416 -3452
rect 422 -3453 423 -3447
rect 502 -3453 503 -3447
rect 541 -3466 542 -3452
rect 569 -3453 570 -3447
rect 625 -3466 626 -3452
rect 632 -3453 633 -3447
rect 646 -3453 647 -3447
rect 646 -3466 647 -3452
rect 646 -3453 647 -3447
rect 646 -3466 647 -3452
rect 653 -3453 654 -3447
rect 653 -3466 654 -3452
rect 653 -3453 654 -3447
rect 653 -3466 654 -3452
rect 674 -3453 675 -3447
rect 691 -3466 692 -3452
rect 695 -3453 696 -3447
rect 709 -3466 710 -3452
rect 719 -3453 720 -3447
rect 730 -3453 731 -3447
rect 824 -3466 825 -3452
rect 961 -3453 962 -3447
rect 275 -3455 276 -3447
rect 306 -3455 307 -3447
rect 317 -3455 318 -3447
rect 327 -3466 328 -3454
rect 345 -3455 346 -3447
rect 352 -3466 353 -3454
rect 394 -3455 395 -3447
rect 471 -3466 472 -3454
rect 569 -3466 570 -3454
rect 583 -3455 584 -3447
rect 667 -3455 668 -3447
rect 674 -3466 675 -3454
rect 681 -3455 682 -3447
rect 716 -3455 717 -3447
rect 835 -3455 836 -3447
rect 891 -3466 892 -3454
rect 940 -3455 941 -3447
rect 940 -3466 941 -3454
rect 940 -3455 941 -3447
rect 940 -3466 941 -3454
rect 947 -3455 948 -3447
rect 975 -3455 976 -3447
rect 282 -3457 283 -3447
rect 303 -3466 304 -3456
rect 310 -3457 311 -3447
rect 317 -3466 318 -3456
rect 387 -3457 388 -3447
rect 394 -3466 395 -3456
rect 422 -3466 423 -3456
rect 429 -3457 430 -3447
rect 443 -3457 444 -3447
rect 443 -3466 444 -3456
rect 443 -3457 444 -3447
rect 443 -3466 444 -3456
rect 450 -3457 451 -3447
rect 457 -3466 458 -3456
rect 576 -3457 577 -3447
rect 583 -3466 584 -3456
rect 660 -3457 661 -3447
rect 681 -3466 682 -3456
rect 688 -3466 689 -3456
rect 744 -3457 745 -3447
rect 821 -3466 822 -3456
rect 835 -3466 836 -3456
rect 842 -3457 843 -3447
rect 842 -3466 843 -3456
rect 842 -3457 843 -3447
rect 842 -3466 843 -3456
rect 849 -3466 850 -3456
rect 870 -3457 871 -3447
rect 296 -3459 297 -3447
rect 331 -3466 332 -3458
rect 425 -3466 426 -3458
rect 639 -3459 640 -3447
rect 660 -3466 661 -3458
rect 726 -3459 727 -3447
rect 863 -3459 864 -3447
rect 870 -3466 871 -3458
rect 429 -3466 430 -3460
rect 436 -3461 437 -3447
rect 555 -3461 556 -3447
rect 576 -3466 577 -3460
rect 695 -3466 696 -3460
rect 758 -3466 759 -3460
rect 555 -3466 556 -3462
rect 562 -3463 563 -3447
rect 534 -3465 535 -3447
rect 562 -3466 563 -3464
rect 261 -3476 262 -3474
rect 268 -3489 269 -3475
rect 303 -3476 304 -3474
rect 310 -3489 311 -3475
rect 317 -3476 318 -3474
rect 327 -3476 328 -3474
rect 331 -3476 332 -3474
rect 331 -3489 332 -3475
rect 331 -3476 332 -3474
rect 331 -3489 332 -3475
rect 338 -3476 339 -3474
rect 338 -3489 339 -3475
rect 338 -3476 339 -3474
rect 338 -3489 339 -3475
rect 352 -3476 353 -3474
rect 352 -3489 353 -3475
rect 352 -3476 353 -3474
rect 352 -3489 353 -3475
rect 380 -3476 381 -3474
rect 411 -3476 412 -3474
rect 415 -3476 416 -3474
rect 436 -3476 437 -3474
rect 467 -3476 468 -3474
rect 520 -3476 521 -3474
rect 541 -3476 542 -3474
rect 541 -3489 542 -3475
rect 541 -3476 542 -3474
rect 541 -3489 542 -3475
rect 548 -3476 549 -3474
rect 551 -3482 552 -3475
rect 569 -3476 570 -3474
rect 569 -3489 570 -3475
rect 569 -3476 570 -3474
rect 569 -3489 570 -3475
rect 583 -3476 584 -3474
rect 590 -3489 591 -3475
rect 597 -3489 598 -3475
rect 660 -3476 661 -3474
rect 681 -3476 682 -3474
rect 688 -3489 689 -3475
rect 695 -3476 696 -3474
rect 828 -3489 829 -3475
rect 835 -3476 836 -3474
rect 835 -3489 836 -3475
rect 835 -3476 836 -3474
rect 835 -3489 836 -3475
rect 842 -3476 843 -3474
rect 849 -3489 850 -3475
rect 852 -3476 853 -3474
rect 856 -3476 857 -3474
rect 870 -3476 871 -3474
rect 887 -3489 888 -3475
rect 891 -3476 892 -3474
rect 950 -3489 951 -3475
rect 989 -3476 990 -3474
rect 992 -3489 993 -3475
rect 996 -3476 997 -3474
rect 996 -3489 997 -3475
rect 996 -3476 997 -3474
rect 996 -3489 997 -3475
rect 1066 -3476 1067 -3474
rect 1094 -3489 1095 -3475
rect 1115 -3476 1116 -3474
rect 1118 -3482 1119 -3475
rect 1213 -3476 1214 -3474
rect 1220 -3476 1221 -3474
rect 1353 -3476 1354 -3474
rect 1353 -3489 1354 -3475
rect 1353 -3476 1354 -3474
rect 1353 -3489 1354 -3475
rect 1360 -3476 1361 -3474
rect 1360 -3489 1361 -3475
rect 1360 -3476 1361 -3474
rect 1360 -3489 1361 -3475
rect 1409 -3476 1410 -3474
rect 1412 -3476 1413 -3474
rect 254 -3478 255 -3474
rect 261 -3489 262 -3477
rect 394 -3478 395 -3474
rect 408 -3478 409 -3474
rect 418 -3489 419 -3477
rect 698 -3478 699 -3474
rect 709 -3478 710 -3474
rect 716 -3489 717 -3477
rect 726 -3489 727 -3477
rect 737 -3478 738 -3474
rect 758 -3478 759 -3474
rect 821 -3478 822 -3474
rect 877 -3489 878 -3477
rect 898 -3489 899 -3477
rect 905 -3489 906 -3477
rect 933 -3478 934 -3474
rect 940 -3478 941 -3474
rect 940 -3489 941 -3477
rect 940 -3478 941 -3474
rect 940 -3489 941 -3477
rect 1115 -3489 1116 -3477
rect 1122 -3478 1123 -3474
rect 1220 -3489 1221 -3477
rect 1227 -3478 1228 -3474
rect 1409 -3489 1410 -3477
rect 1416 -3478 1417 -3474
rect 401 -3480 402 -3474
rect 408 -3489 409 -3479
rect 429 -3480 430 -3474
rect 439 -3480 440 -3474
rect 471 -3480 472 -3474
rect 506 -3480 507 -3474
rect 548 -3489 549 -3479
rect 576 -3480 577 -3474
rect 583 -3489 584 -3479
rect 604 -3480 605 -3474
rect 621 -3480 622 -3474
rect 646 -3480 647 -3474
rect 660 -3489 661 -3479
rect 674 -3480 675 -3474
rect 681 -3489 682 -3479
rect 884 -3480 885 -3474
rect 884 -3489 885 -3479
rect 884 -3480 885 -3474
rect 884 -3489 885 -3479
rect 912 -3480 913 -3474
rect 912 -3489 913 -3479
rect 912 -3480 913 -3474
rect 912 -3489 913 -3479
rect 919 -3480 920 -3474
rect 919 -3489 920 -3479
rect 919 -3480 920 -3474
rect 919 -3489 920 -3479
rect 926 -3480 927 -3474
rect 926 -3489 927 -3479
rect 926 -3480 927 -3474
rect 926 -3489 927 -3479
rect 359 -3482 360 -3474
rect 429 -3489 430 -3481
rect 436 -3489 437 -3481
rect 443 -3482 444 -3474
rect 478 -3482 479 -3474
rect 502 -3482 503 -3474
rect 513 -3482 514 -3474
rect 646 -3489 647 -3481
rect 653 -3482 654 -3474
rect 653 -3489 654 -3481
rect 653 -3482 654 -3474
rect 653 -3489 654 -3481
rect 1412 -3489 1413 -3481
rect 1416 -3489 1417 -3481
rect 478 -3489 479 -3483
rect 614 -3484 615 -3474
rect 485 -3486 486 -3474
rect 516 -3486 517 -3474
rect 562 -3486 563 -3474
rect 576 -3489 577 -3485
rect 611 -3486 612 -3474
rect 625 -3486 626 -3474
rect 492 -3488 493 -3474
rect 499 -3488 500 -3474
rect 261 -3499 262 -3497
rect 271 -3504 272 -3498
rect 310 -3499 311 -3497
rect 324 -3504 325 -3498
rect 331 -3499 332 -3497
rect 345 -3499 346 -3497
rect 352 -3499 353 -3497
rect 359 -3504 360 -3498
rect 408 -3499 409 -3497
rect 418 -3499 419 -3497
rect 429 -3499 430 -3497
rect 436 -3499 437 -3497
rect 541 -3499 542 -3497
rect 551 -3504 552 -3498
rect 555 -3499 556 -3497
rect 565 -3504 566 -3498
rect 569 -3499 570 -3497
rect 569 -3504 570 -3498
rect 569 -3499 570 -3497
rect 569 -3504 570 -3498
rect 583 -3499 584 -3497
rect 597 -3499 598 -3497
rect 646 -3499 647 -3497
rect 653 -3499 654 -3497
rect 660 -3499 661 -3497
rect 667 -3504 668 -3498
rect 681 -3499 682 -3497
rect 691 -3504 692 -3498
rect 716 -3499 717 -3497
rect 723 -3499 724 -3497
rect 828 -3499 829 -3497
rect 870 -3504 871 -3498
rect 877 -3499 878 -3497
rect 877 -3504 878 -3498
rect 877 -3499 878 -3497
rect 877 -3504 878 -3498
rect 898 -3499 899 -3497
rect 905 -3499 906 -3497
rect 912 -3499 913 -3497
rect 912 -3504 913 -3498
rect 912 -3499 913 -3497
rect 912 -3504 913 -3498
rect 919 -3499 920 -3497
rect 919 -3504 920 -3498
rect 919 -3499 920 -3497
rect 919 -3504 920 -3498
rect 922 -3504 923 -3498
rect 926 -3499 927 -3497
rect 940 -3499 941 -3497
rect 950 -3499 951 -3497
rect 989 -3499 990 -3497
rect 996 -3499 997 -3497
rect 1094 -3499 1095 -3497
rect 1115 -3499 1116 -3497
rect 1118 -3499 1119 -3497
rect 1122 -3499 1123 -3497
rect 1353 -3499 1354 -3497
rect 1353 -3504 1354 -3498
rect 1353 -3499 1354 -3497
rect 1353 -3504 1354 -3498
rect 1360 -3499 1361 -3497
rect 1367 -3504 1368 -3498
rect 1412 -3499 1413 -3497
rect 1416 -3499 1417 -3497
rect 268 -3501 269 -3497
rect 275 -3504 276 -3500
rect 331 -3504 332 -3500
rect 338 -3501 339 -3497
rect 355 -3504 356 -3500
rect 478 -3501 479 -3497
rect 541 -3504 542 -3500
rect 548 -3501 549 -3497
rect 576 -3501 577 -3497
rect 583 -3504 584 -3500
rect 688 -3501 689 -3497
rect 688 -3504 689 -3500
rect 688 -3501 689 -3497
rect 688 -3504 689 -3500
rect 835 -3501 836 -3497
rect 859 -3504 860 -3500
rect 576 -3504 577 -3502
rect 590 -3503 591 -3497
rect 842 -3503 843 -3497
rect 849 -3503 850 -3497
rect 271 -3514 272 -3512
rect 275 -3514 276 -3512
rect 327 -3514 328 -3512
rect 331 -3514 332 -3512
rect 355 -3514 356 -3512
rect 359 -3514 360 -3512
rect 541 -3514 542 -3512
rect 555 -3514 556 -3512
rect 565 -3514 566 -3512
rect 569 -3514 570 -3512
rect 579 -3514 580 -3512
rect 583 -3514 584 -3512
rect 660 -3514 661 -3512
rect 667 -3514 668 -3512
rect 856 -3514 857 -3512
rect 877 -3514 878 -3512
rect 1353 -3514 1354 -3512
rect 1360 -3514 1361 -3512
rect 1363 -3514 1364 -3512
rect 1367 -3514 1368 -3512
rect 870 -3516 871 -3512
rect 915 -3516 916 -3512
<< labels >>
rlabel pdiffusion 3 -10 3 -10 0 cellNo=156
rlabel pdiffusion 10 -10 10 -10 0 cellNo=1083
rlabel pdiffusion 17 -10 17 -10 0 cellNo=1007
rlabel pdiffusion 24 -10 24 -10 0 cellNo=1046
rlabel pdiffusion 31 -10 31 -10 0 cellNo=1087
rlabel pdiffusion 38 -10 38 -10 0 cellNo=1094
rlabel pdiffusion 45 -10 45 -10 0 cellNo=1010
rlabel pdiffusion 52 -10 52 -10 0 cellNo=1020
rlabel pdiffusion 59 -10 59 -10 0 cellNo=1036
rlabel pdiffusion 66 -10 66 -10 0 cellNo=1032
rlabel pdiffusion 73 -10 73 -10 0 cellNo=1042
rlabel pdiffusion 80 -10 80 -10 0 cellNo=1056
rlabel pdiffusion 87 -10 87 -10 0 cellNo=1068
rlabel pdiffusion 94 -10 94 -10 0 cellNo=1082
rlabel pdiffusion 101 -10 101 -10 0 cellNo=1099
rlabel pdiffusion 108 -10 108 -10 0 cellNo=1111
rlabel pdiffusion 115 -10 115 -10 0 cellNo=1143
rlabel pdiffusion 122 -10 122 -10 0 cellNo=1148
rlabel pdiffusion 129 -10 129 -10 0 cellNo=1154
rlabel pdiffusion 136 -10 136 -10 0 cellNo=1170
rlabel pdiffusion 143 -10 143 -10 0 cellNo=1180
rlabel pdiffusion 150 -10 150 -10 0 cellNo=1189
rlabel pdiffusion 283 -10 283 -10 0 cellNo=883
rlabel pdiffusion 318 -10 318 -10 0 feedthrough
rlabel pdiffusion 346 -10 346 -10 0 feedthrough
rlabel pdiffusion 353 -10 353 -10 0 cellNo=886
rlabel pdiffusion 423 -10 423 -10 0 cellNo=548
rlabel pdiffusion 437 -10 437 -10 0 cellNo=518
rlabel pdiffusion 444 -10 444 -10 0 feedthrough
rlabel pdiffusion 451 -10 451 -10 0 feedthrough
rlabel pdiffusion 458 -10 458 -10 0 cellNo=661
rlabel pdiffusion 465 -10 465 -10 0 feedthrough
rlabel pdiffusion 479 -10 479 -10 0 cellNo=342
rlabel pdiffusion 507 -10 507 -10 0 cellNo=972
rlabel pdiffusion 514 -10 514 -10 0 feedthrough
rlabel pdiffusion 906 -10 906 -10 0 feedthrough
rlabel pdiffusion 948 -10 948 -10 0 cellNo=682
rlabel pdiffusion 990 -10 990 -10 0 feedthrough
rlabel pdiffusion 3 -29 3 -29 0 cellNo=520
rlabel pdiffusion 10 -29 10 -29 0 cellNo=590
rlabel pdiffusion 17 -29 17 -29 0 cellNo=1017
rlabel pdiffusion 24 -29 24 -29 0 cellNo=1004
rlabel pdiffusion 31 -29 31 -29 0 cellNo=1005
rlabel pdiffusion 38 -29 38 -29 0 cellNo=1168
rlabel pdiffusion 45 -29 45 -29 0 cellNo=1019
rlabel pdiffusion 52 -29 52 -29 0 cellNo=1024
rlabel pdiffusion 59 -29 59 -29 0 cellNo=1164
rlabel pdiffusion 66 -29 66 -29 0 cellNo=1169
rlabel pdiffusion 73 -29 73 -29 0 cellNo=1055
rlabel pdiffusion 80 -29 80 -29 0 cellNo=1067
rlabel pdiffusion 87 -29 87 -29 0 cellNo=1081
rlabel pdiffusion 94 -29 94 -29 0 cellNo=1098
rlabel pdiffusion 101 -29 101 -29 0 cellNo=1179
rlabel pdiffusion 108 -29 108 -29 0 cellNo=1193
rlabel pdiffusion 115 -29 115 -29 0 cellNo=1188
rlabel pdiffusion 227 -29 227 -29 0 feedthrough
rlabel pdiffusion 290 -29 290 -29 0 feedthrough
rlabel pdiffusion 304 -29 304 -29 0 feedthrough
rlabel pdiffusion 339 -29 339 -29 0 feedthrough
rlabel pdiffusion 346 -29 346 -29 0 cellNo=846
rlabel pdiffusion 353 -29 353 -29 0 feedthrough
rlabel pdiffusion 360 -29 360 -29 0 cellNo=976
rlabel pdiffusion 367 -29 367 -29 0 feedthrough
rlabel pdiffusion 374 -29 374 -29 0 feedthrough
rlabel pdiffusion 381 -29 381 -29 0 feedthrough
rlabel pdiffusion 388 -29 388 -29 0 feedthrough
rlabel pdiffusion 395 -29 395 -29 0 feedthrough
rlabel pdiffusion 409 -29 409 -29 0 feedthrough
rlabel pdiffusion 416 -29 416 -29 0 cellNo=834
rlabel pdiffusion 423 -29 423 -29 0 feedthrough
rlabel pdiffusion 437 -29 437 -29 0 feedthrough
rlabel pdiffusion 451 -29 451 -29 0 feedthrough
rlabel pdiffusion 458 -29 458 -29 0 feedthrough
rlabel pdiffusion 465 -29 465 -29 0 feedthrough
rlabel pdiffusion 500 -29 500 -29 0 feedthrough
rlabel pdiffusion 507 -29 507 -29 0 cellNo=816
rlabel pdiffusion 514 -29 514 -29 0 feedthrough
rlabel pdiffusion 521 -29 521 -29 0 cellNo=634
rlabel pdiffusion 528 -29 528 -29 0 cellNo=612
rlabel pdiffusion 535 -29 535 -29 0 cellNo=756
rlabel pdiffusion 542 -29 542 -29 0 feedthrough
rlabel pdiffusion 549 -29 549 -29 0 feedthrough
rlabel pdiffusion 577 -29 577 -29 0 cellNo=118
rlabel pdiffusion 584 -29 584 -29 0 cellNo=833
rlabel pdiffusion 591 -29 591 -29 0 feedthrough
rlabel pdiffusion 598 -29 598 -29 0 feedthrough
rlabel pdiffusion 605 -29 605 -29 0 feedthrough
rlabel pdiffusion 612 -29 612 -29 0 feedthrough
rlabel pdiffusion 619 -29 619 -29 0 cellNo=475
rlabel pdiffusion 626 -29 626 -29 0 feedthrough
rlabel pdiffusion 633 -29 633 -29 0 cellNo=153
rlabel pdiffusion 640 -29 640 -29 0 cellNo=400
rlabel pdiffusion 675 -29 675 -29 0 feedthrough
rlabel pdiffusion 892 -29 892 -29 0 feedthrough
rlabel pdiffusion 1004 -29 1004 -29 0 feedthrough
rlabel pdiffusion 3 -52 3 -52 0 cellNo=1002
rlabel pdiffusion 10 -52 10 -52 0 cellNo=1075
rlabel pdiffusion 17 -52 17 -52 0 cellNo=1012
rlabel pdiffusion 24 -52 24 -52 0 cellNo=1187
rlabel pdiffusion 31 -52 31 -52 0 cellNo=1038
rlabel pdiffusion 38 -52 38 -52 0 cellNo=1018
rlabel pdiffusion 45 -52 45 -52 0 cellNo=1132
rlabel pdiffusion 52 -52 52 -52 0 cellNo=1031
rlabel pdiffusion 59 -52 59 -52 0 cellNo=1041
rlabel pdiffusion 66 -52 66 -52 0 cellNo=1054
rlabel pdiffusion 73 -52 73 -52 0 cellNo=1066
rlabel pdiffusion 80 -52 80 -52 0 cellNo=1080
rlabel pdiffusion 87 -52 87 -52 0 cellNo=1161
rlabel pdiffusion 94 -52 94 -52 0 cellNo=1178
rlabel pdiffusion 101 -52 101 -52 0 cellNo=1199
rlabel pdiffusion 108 -52 108 -52 0 cellNo=1085
rlabel pdiffusion 220 -52 220 -52 0 feedthrough
rlabel pdiffusion 276 -52 276 -52 0 feedthrough
rlabel pdiffusion 283 -52 283 -52 0 feedthrough
rlabel pdiffusion 297 -52 297 -52 0 cellNo=145
rlabel pdiffusion 304 -52 304 -52 0 feedthrough
rlabel pdiffusion 318 -52 318 -52 0 cellNo=151
rlabel pdiffusion 325 -52 325 -52 0 feedthrough
rlabel pdiffusion 332 -52 332 -52 0 feedthrough
rlabel pdiffusion 339 -52 339 -52 0 cellNo=623
rlabel pdiffusion 346 -52 346 -52 0 feedthrough
rlabel pdiffusion 353 -52 353 -52 0 feedthrough
rlabel pdiffusion 360 -52 360 -52 0 feedthrough
rlabel pdiffusion 367 -52 367 -52 0 feedthrough
rlabel pdiffusion 374 -52 374 -52 0 feedthrough
rlabel pdiffusion 381 -52 381 -52 0 feedthrough
rlabel pdiffusion 388 -52 388 -52 0 cellNo=396
rlabel pdiffusion 395 -52 395 -52 0 feedthrough
rlabel pdiffusion 402 -52 402 -52 0 feedthrough
rlabel pdiffusion 409 -52 409 -52 0 feedthrough
rlabel pdiffusion 416 -52 416 -52 0 feedthrough
rlabel pdiffusion 423 -52 423 -52 0 feedthrough
rlabel pdiffusion 430 -52 430 -52 0 cellNo=649
rlabel pdiffusion 437 -52 437 -52 0 feedthrough
rlabel pdiffusion 444 -52 444 -52 0 feedthrough
rlabel pdiffusion 451 -52 451 -52 0 feedthrough
rlabel pdiffusion 458 -52 458 -52 0 cellNo=221
rlabel pdiffusion 465 -52 465 -52 0 feedthrough
rlabel pdiffusion 472 -52 472 -52 0 feedthrough
rlabel pdiffusion 486 -52 486 -52 0 feedthrough
rlabel pdiffusion 493 -52 493 -52 0 feedthrough
rlabel pdiffusion 500 -52 500 -52 0 feedthrough
rlabel pdiffusion 507 -52 507 -52 0 feedthrough
rlabel pdiffusion 521 -52 521 -52 0 feedthrough
rlabel pdiffusion 542 -52 542 -52 0 feedthrough
rlabel pdiffusion 549 -52 549 -52 0 cellNo=896
rlabel pdiffusion 556 -52 556 -52 0 feedthrough
rlabel pdiffusion 563 -52 563 -52 0 cellNo=68
rlabel pdiffusion 570 -52 570 -52 0 cellNo=711
rlabel pdiffusion 577 -52 577 -52 0 feedthrough
rlabel pdiffusion 584 -52 584 -52 0 feedthrough
rlabel pdiffusion 591 -52 591 -52 0 feedthrough
rlabel pdiffusion 598 -52 598 -52 0 feedthrough
rlabel pdiffusion 605 -52 605 -52 0 feedthrough
rlabel pdiffusion 612 -52 612 -52 0 cellNo=785
rlabel pdiffusion 619 -52 619 -52 0 cellNo=25
rlabel pdiffusion 626 -52 626 -52 0 feedthrough
rlabel pdiffusion 633 -52 633 -52 0 feedthrough
rlabel pdiffusion 640 -52 640 -52 0 feedthrough
rlabel pdiffusion 654 -52 654 -52 0 feedthrough
rlabel pdiffusion 675 -52 675 -52 0 feedthrough
rlabel pdiffusion 682 -52 682 -52 0 cellNo=176
rlabel pdiffusion 724 -52 724 -52 0 feedthrough
rlabel pdiffusion 731 -52 731 -52 0 feedthrough
rlabel pdiffusion 759 -52 759 -52 0 feedthrough
rlabel pdiffusion 829 -52 829 -52 0 cellNo=116
rlabel pdiffusion 885 -52 885 -52 0 feedthrough
rlabel pdiffusion 1011 -52 1011 -52 0 feedthrough
rlabel pdiffusion 3 -103 3 -103 0 cellNo=443
rlabel pdiffusion 10 -103 10 -103 0 cellNo=1003
rlabel pdiffusion 17 -103 17 -103 0 cellNo=1166
rlabel pdiffusion 24 -103 24 -103 0 cellNo=1009
rlabel pdiffusion 31 -103 31 -103 0 cellNo=1016
rlabel pdiffusion 38 -103 38 -103 0 cellNo=1026
rlabel pdiffusion 45 -103 45 -103 0 cellNo=1062
rlabel pdiffusion 52 -103 52 -103 0 cellNo=1040
rlabel pdiffusion 59 -103 59 -103 0 cellNo=1052
rlabel pdiffusion 66 -103 66 -103 0 cellNo=1065
rlabel pdiffusion 73 -103 73 -103 0 cellNo=1079
rlabel pdiffusion 80 -103 80 -103 0 cellNo=1197
rlabel pdiffusion 192 -103 192 -103 0 feedthrough
rlabel pdiffusion 206 -103 206 -103 0 feedthrough
rlabel pdiffusion 220 -103 220 -103 0 feedthrough
rlabel pdiffusion 234 -103 234 -103 0 feedthrough
rlabel pdiffusion 241 -103 241 -103 0 cellNo=316
rlabel pdiffusion 248 -103 248 -103 0 feedthrough
rlabel pdiffusion 255 -103 255 -103 0 cellNo=843
rlabel pdiffusion 262 -103 262 -103 0 feedthrough
rlabel pdiffusion 269 -103 269 -103 0 cellNo=703
rlabel pdiffusion 276 -103 276 -103 0 cellNo=131
rlabel pdiffusion 283 -103 283 -103 0 feedthrough
rlabel pdiffusion 290 -103 290 -103 0 feedthrough
rlabel pdiffusion 297 -103 297 -103 0 cellNo=200
rlabel pdiffusion 304 -103 304 -103 0 feedthrough
rlabel pdiffusion 311 -103 311 -103 0 feedthrough
rlabel pdiffusion 318 -103 318 -103 0 feedthrough
rlabel pdiffusion 325 -103 325 -103 0 feedthrough
rlabel pdiffusion 332 -103 332 -103 0 feedthrough
rlabel pdiffusion 339 -103 339 -103 0 feedthrough
rlabel pdiffusion 346 -103 346 -103 0 feedthrough
rlabel pdiffusion 353 -103 353 -103 0 feedthrough
rlabel pdiffusion 360 -103 360 -103 0 feedthrough
rlabel pdiffusion 367 -103 367 -103 0 feedthrough
rlabel pdiffusion 374 -103 374 -103 0 feedthrough
rlabel pdiffusion 381 -103 381 -103 0 cellNo=602
rlabel pdiffusion 388 -103 388 -103 0 cellNo=867
rlabel pdiffusion 395 -103 395 -103 0 feedthrough
rlabel pdiffusion 402 -103 402 -103 0 feedthrough
rlabel pdiffusion 409 -103 409 -103 0 feedthrough
rlabel pdiffusion 416 -103 416 -103 0 feedthrough
rlabel pdiffusion 423 -103 423 -103 0 feedthrough
rlabel pdiffusion 430 -103 430 -103 0 feedthrough
rlabel pdiffusion 437 -103 437 -103 0 feedthrough
rlabel pdiffusion 444 -103 444 -103 0 feedthrough
rlabel pdiffusion 451 -103 451 -103 0 feedthrough
rlabel pdiffusion 458 -103 458 -103 0 feedthrough
rlabel pdiffusion 465 -103 465 -103 0 feedthrough
rlabel pdiffusion 472 -103 472 -103 0 feedthrough
rlabel pdiffusion 479 -103 479 -103 0 feedthrough
rlabel pdiffusion 486 -103 486 -103 0 feedthrough
rlabel pdiffusion 493 -103 493 -103 0 feedthrough
rlabel pdiffusion 500 -103 500 -103 0 feedthrough
rlabel pdiffusion 507 -103 507 -103 0 cellNo=849
rlabel pdiffusion 514 -103 514 -103 0 cellNo=747
rlabel pdiffusion 521 -103 521 -103 0 cellNo=624
rlabel pdiffusion 528 -103 528 -103 0 feedthrough
rlabel pdiffusion 535 -103 535 -103 0 cellNo=380
rlabel pdiffusion 542 -103 542 -103 0 cellNo=58
rlabel pdiffusion 549 -103 549 -103 0 feedthrough
rlabel pdiffusion 556 -103 556 -103 0 feedthrough
rlabel pdiffusion 563 -103 563 -103 0 cellNo=23
rlabel pdiffusion 570 -103 570 -103 0 feedthrough
rlabel pdiffusion 577 -103 577 -103 0 feedthrough
rlabel pdiffusion 584 -103 584 -103 0 cellNo=814
rlabel pdiffusion 591 -103 591 -103 0 feedthrough
rlabel pdiffusion 598 -103 598 -103 0 feedthrough
rlabel pdiffusion 605 -103 605 -103 0 feedthrough
rlabel pdiffusion 612 -103 612 -103 0 feedthrough
rlabel pdiffusion 619 -103 619 -103 0 feedthrough
rlabel pdiffusion 626 -103 626 -103 0 cellNo=782
rlabel pdiffusion 633 -103 633 -103 0 feedthrough
rlabel pdiffusion 640 -103 640 -103 0 feedthrough
rlabel pdiffusion 647 -103 647 -103 0 feedthrough
rlabel pdiffusion 654 -103 654 -103 0 feedthrough
rlabel pdiffusion 661 -103 661 -103 0 feedthrough
rlabel pdiffusion 668 -103 668 -103 0 feedthrough
rlabel pdiffusion 682 -103 682 -103 0 feedthrough
rlabel pdiffusion 689 -103 689 -103 0 feedthrough
rlabel pdiffusion 703 -103 703 -103 0 feedthrough
rlabel pdiffusion 710 -103 710 -103 0 feedthrough
rlabel pdiffusion 724 -103 724 -103 0 feedthrough
rlabel pdiffusion 731 -103 731 -103 0 feedthrough
rlabel pdiffusion 738 -103 738 -103 0 feedthrough
rlabel pdiffusion 780 -103 780 -103 0 cellNo=897
rlabel pdiffusion 787 -103 787 -103 0 cellNo=442
rlabel pdiffusion 794 -103 794 -103 0 feedthrough
rlabel pdiffusion 801 -103 801 -103 0 cellNo=290
rlabel pdiffusion 808 -103 808 -103 0 feedthrough
rlabel pdiffusion 864 -103 864 -103 0 feedthrough
rlabel pdiffusion 892 -103 892 -103 0 feedthrough
rlabel pdiffusion 899 -103 899 -103 0 feedthrough
rlabel pdiffusion 1018 -103 1018 -103 0 feedthrough
rlabel pdiffusion 3 -170 3 -170 0 cellNo=1001
rlabel pdiffusion 10 -170 10 -170 0 cellNo=1157
rlabel pdiffusion 17 -170 17 -170 0 cellNo=1008
rlabel pdiffusion 24 -170 24 -170 0 cellNo=1015
rlabel pdiffusion 31 -170 31 -170 0 cellNo=1025
rlabel pdiffusion 38 -170 38 -170 0 cellNo=1030
rlabel pdiffusion 45 -170 45 -170 0 cellNo=1039
rlabel pdiffusion 52 -170 52 -170 0 cellNo=1051
rlabel pdiffusion 59 -170 59 -170 0 cellNo=1064
rlabel pdiffusion 66 -170 66 -170 0 cellNo=1078
rlabel pdiffusion 73 -170 73 -170 0 cellNo=1097
rlabel pdiffusion 80 -170 80 -170 0 cellNo=1107
rlabel pdiffusion 115 -170 115 -170 0 feedthrough
rlabel pdiffusion 122 -170 122 -170 0 feedthrough
rlabel pdiffusion 129 -170 129 -170 0 feedthrough
rlabel pdiffusion 136 -170 136 -170 0 feedthrough
rlabel pdiffusion 143 -170 143 -170 0 feedthrough
rlabel pdiffusion 150 -170 150 -170 0 feedthrough
rlabel pdiffusion 157 -170 157 -170 0 feedthrough
rlabel pdiffusion 164 -170 164 -170 0 feedthrough
rlabel pdiffusion 171 -170 171 -170 0 feedthrough
rlabel pdiffusion 178 -170 178 -170 0 feedthrough
rlabel pdiffusion 185 -170 185 -170 0 feedthrough
rlabel pdiffusion 192 -170 192 -170 0 feedthrough
rlabel pdiffusion 199 -170 199 -170 0 feedthrough
rlabel pdiffusion 206 -170 206 -170 0 feedthrough
rlabel pdiffusion 213 -170 213 -170 0 feedthrough
rlabel pdiffusion 220 -170 220 -170 0 feedthrough
rlabel pdiffusion 227 -170 227 -170 0 cellNo=505
rlabel pdiffusion 234 -170 234 -170 0 feedthrough
rlabel pdiffusion 241 -170 241 -170 0 feedthrough
rlabel pdiffusion 248 -170 248 -170 0 feedthrough
rlabel pdiffusion 255 -170 255 -170 0 feedthrough
rlabel pdiffusion 262 -170 262 -170 0 feedthrough
rlabel pdiffusion 269 -170 269 -170 0 feedthrough
rlabel pdiffusion 276 -170 276 -170 0 feedthrough
rlabel pdiffusion 283 -170 283 -170 0 feedthrough
rlabel pdiffusion 290 -170 290 -170 0 feedthrough
rlabel pdiffusion 297 -170 297 -170 0 cellNo=84
rlabel pdiffusion 304 -170 304 -170 0 feedthrough
rlabel pdiffusion 311 -170 311 -170 0 feedthrough
rlabel pdiffusion 318 -170 318 -170 0 feedthrough
rlabel pdiffusion 325 -170 325 -170 0 feedthrough
rlabel pdiffusion 332 -170 332 -170 0 cellNo=82
rlabel pdiffusion 339 -170 339 -170 0 feedthrough
rlabel pdiffusion 346 -170 346 -170 0 feedthrough
rlabel pdiffusion 353 -170 353 -170 0 feedthrough
rlabel pdiffusion 360 -170 360 -170 0 feedthrough
rlabel pdiffusion 367 -170 367 -170 0 cellNo=306
rlabel pdiffusion 374 -170 374 -170 0 feedthrough
rlabel pdiffusion 381 -170 381 -170 0 feedthrough
rlabel pdiffusion 388 -170 388 -170 0 cellNo=383
rlabel pdiffusion 395 -170 395 -170 0 feedthrough
rlabel pdiffusion 402 -170 402 -170 0 cellNo=840
rlabel pdiffusion 409 -170 409 -170 0 feedthrough
rlabel pdiffusion 416 -170 416 -170 0 feedthrough
rlabel pdiffusion 423 -170 423 -170 0 feedthrough
rlabel pdiffusion 430 -170 430 -170 0 feedthrough
rlabel pdiffusion 437 -170 437 -170 0 feedthrough
rlabel pdiffusion 444 -170 444 -170 0 feedthrough
rlabel pdiffusion 451 -170 451 -170 0 cellNo=477
rlabel pdiffusion 458 -170 458 -170 0 feedthrough
rlabel pdiffusion 465 -170 465 -170 0 feedthrough
rlabel pdiffusion 472 -170 472 -170 0 feedthrough
rlabel pdiffusion 479 -170 479 -170 0 feedthrough
rlabel pdiffusion 486 -170 486 -170 0 feedthrough
rlabel pdiffusion 493 -170 493 -170 0 feedthrough
rlabel pdiffusion 500 -170 500 -170 0 cellNo=870
rlabel pdiffusion 507 -170 507 -170 0 feedthrough
rlabel pdiffusion 514 -170 514 -170 0 cellNo=296
rlabel pdiffusion 521 -170 521 -170 0 cellNo=605
rlabel pdiffusion 528 -170 528 -170 0 cellNo=781
rlabel pdiffusion 535 -170 535 -170 0 feedthrough
rlabel pdiffusion 542 -170 542 -170 0 feedthrough
rlabel pdiffusion 549 -170 549 -170 0 feedthrough
rlabel pdiffusion 556 -170 556 -170 0 cellNo=289
rlabel pdiffusion 563 -170 563 -170 0 feedthrough
rlabel pdiffusion 570 -170 570 -170 0 cellNo=70
rlabel pdiffusion 577 -170 577 -170 0 feedthrough
rlabel pdiffusion 584 -170 584 -170 0 feedthrough
rlabel pdiffusion 591 -170 591 -170 0 cellNo=618
rlabel pdiffusion 598 -170 598 -170 0 feedthrough
rlabel pdiffusion 605 -170 605 -170 0 cellNo=928
rlabel pdiffusion 612 -170 612 -170 0 cellNo=732
rlabel pdiffusion 619 -170 619 -170 0 feedthrough
rlabel pdiffusion 626 -170 626 -170 0 feedthrough
rlabel pdiffusion 633 -170 633 -170 0 feedthrough
rlabel pdiffusion 640 -170 640 -170 0 feedthrough
rlabel pdiffusion 647 -170 647 -170 0 feedthrough
rlabel pdiffusion 654 -170 654 -170 0 cellNo=774
rlabel pdiffusion 661 -170 661 -170 0 feedthrough
rlabel pdiffusion 668 -170 668 -170 0 feedthrough
rlabel pdiffusion 675 -170 675 -170 0 feedthrough
rlabel pdiffusion 682 -170 682 -170 0 feedthrough
rlabel pdiffusion 689 -170 689 -170 0 feedthrough
rlabel pdiffusion 696 -170 696 -170 0 feedthrough
rlabel pdiffusion 703 -170 703 -170 0 feedthrough
rlabel pdiffusion 710 -170 710 -170 0 feedthrough
rlabel pdiffusion 717 -170 717 -170 0 feedthrough
rlabel pdiffusion 724 -170 724 -170 0 feedthrough
rlabel pdiffusion 731 -170 731 -170 0 cellNo=324
rlabel pdiffusion 738 -170 738 -170 0 feedthrough
rlabel pdiffusion 745 -170 745 -170 0 feedthrough
rlabel pdiffusion 752 -170 752 -170 0 feedthrough
rlabel pdiffusion 759 -170 759 -170 0 feedthrough
rlabel pdiffusion 766 -170 766 -170 0 feedthrough
rlabel pdiffusion 773 -170 773 -170 0 feedthrough
rlabel pdiffusion 780 -170 780 -170 0 feedthrough
rlabel pdiffusion 787 -170 787 -170 0 feedthrough
rlabel pdiffusion 794 -170 794 -170 0 feedthrough
rlabel pdiffusion 801 -170 801 -170 0 feedthrough
rlabel pdiffusion 808 -170 808 -170 0 feedthrough
rlabel pdiffusion 815 -170 815 -170 0 feedthrough
rlabel pdiffusion 822 -170 822 -170 0 feedthrough
rlabel pdiffusion 829 -170 829 -170 0 feedthrough
rlabel pdiffusion 836 -170 836 -170 0 feedthrough
rlabel pdiffusion 843 -170 843 -170 0 feedthrough
rlabel pdiffusion 850 -170 850 -170 0 feedthrough
rlabel pdiffusion 857 -170 857 -170 0 feedthrough
rlabel pdiffusion 864 -170 864 -170 0 feedthrough
rlabel pdiffusion 871 -170 871 -170 0 feedthrough
rlabel pdiffusion 878 -170 878 -170 0 feedthrough
rlabel pdiffusion 899 -170 899 -170 0 feedthrough
rlabel pdiffusion 920 -170 920 -170 0 feedthrough
rlabel pdiffusion 941 -170 941 -170 0 feedthrough
rlabel pdiffusion 1011 -170 1011 -170 0 cellNo=651
rlabel pdiffusion 1025 -170 1025 -170 0 feedthrough
rlabel pdiffusion 1137 -170 1137 -170 0 feedthrough
rlabel pdiffusion 1172 -170 1172 -170 0 feedthrough
rlabel pdiffusion 3 -237 3 -237 0 cellNo=1006
rlabel pdiffusion 10 -237 10 -237 0 cellNo=1053
rlabel pdiffusion 17 -237 17 -237 0 cellNo=1014
rlabel pdiffusion 24 -237 24 -237 0 cellNo=1023
rlabel pdiffusion 31 -237 31 -237 0 cellNo=1029
rlabel pdiffusion 38 -237 38 -237 0 cellNo=1158
rlabel pdiffusion 45 -237 45 -237 0 cellNo=1050
rlabel pdiffusion 52 -237 52 -237 0 cellNo=1130
rlabel pdiffusion 59 -237 59 -237 0 cellNo=1077
rlabel pdiffusion 66 -237 66 -237 0 cellNo=1096
rlabel pdiffusion 73 -237 73 -237 0 feedthrough
rlabel pdiffusion 80 -237 80 -237 0 feedthrough
rlabel pdiffusion 87 -237 87 -237 0 feedthrough
rlabel pdiffusion 94 -237 94 -237 0 feedthrough
rlabel pdiffusion 101 -237 101 -237 0 feedthrough
rlabel pdiffusion 108 -237 108 -237 0 feedthrough
rlabel pdiffusion 115 -237 115 -237 0 feedthrough
rlabel pdiffusion 122 -237 122 -237 0 feedthrough
rlabel pdiffusion 129 -237 129 -237 0 feedthrough
rlabel pdiffusion 136 -237 136 -237 0 feedthrough
rlabel pdiffusion 143 -237 143 -237 0 feedthrough
rlabel pdiffusion 150 -237 150 -237 0 feedthrough
rlabel pdiffusion 157 -237 157 -237 0 cellNo=790
rlabel pdiffusion 164 -237 164 -237 0 feedthrough
rlabel pdiffusion 171 -237 171 -237 0 feedthrough
rlabel pdiffusion 178 -237 178 -237 0 feedthrough
rlabel pdiffusion 185 -237 185 -237 0 feedthrough
rlabel pdiffusion 192 -237 192 -237 0 feedthrough
rlabel pdiffusion 199 -237 199 -237 0 feedthrough
rlabel pdiffusion 206 -237 206 -237 0 cellNo=696
rlabel pdiffusion 213 -237 213 -237 0 feedthrough
rlabel pdiffusion 220 -237 220 -237 0 cellNo=64
rlabel pdiffusion 227 -237 227 -237 0 cellNo=8
rlabel pdiffusion 234 -237 234 -237 0 cellNo=359
rlabel pdiffusion 241 -237 241 -237 0 cellNo=1000
rlabel pdiffusion 248 -237 248 -237 0 feedthrough
rlabel pdiffusion 255 -237 255 -237 0 cellNo=544
rlabel pdiffusion 262 -237 262 -237 0 feedthrough
rlabel pdiffusion 269 -237 269 -237 0 feedthrough
rlabel pdiffusion 276 -237 276 -237 0 feedthrough
rlabel pdiffusion 283 -237 283 -237 0 feedthrough
rlabel pdiffusion 290 -237 290 -237 0 feedthrough
rlabel pdiffusion 297 -237 297 -237 0 feedthrough
rlabel pdiffusion 304 -237 304 -237 0 feedthrough
rlabel pdiffusion 311 -237 311 -237 0 feedthrough
rlabel pdiffusion 318 -237 318 -237 0 feedthrough
rlabel pdiffusion 325 -237 325 -237 0 feedthrough
rlabel pdiffusion 332 -237 332 -237 0 feedthrough
rlabel pdiffusion 339 -237 339 -237 0 feedthrough
rlabel pdiffusion 346 -237 346 -237 0 feedthrough
rlabel pdiffusion 353 -237 353 -237 0 feedthrough
rlabel pdiffusion 360 -237 360 -237 0 feedthrough
rlabel pdiffusion 367 -237 367 -237 0 cellNo=948
rlabel pdiffusion 374 -237 374 -237 0 feedthrough
rlabel pdiffusion 381 -237 381 -237 0 feedthrough
rlabel pdiffusion 388 -237 388 -237 0 feedthrough
rlabel pdiffusion 395 -237 395 -237 0 feedthrough
rlabel pdiffusion 402 -237 402 -237 0 feedthrough
rlabel pdiffusion 409 -237 409 -237 0 cellNo=155
rlabel pdiffusion 416 -237 416 -237 0 feedthrough
rlabel pdiffusion 423 -237 423 -237 0 feedthrough
rlabel pdiffusion 430 -237 430 -237 0 cellNo=613
rlabel pdiffusion 437 -237 437 -237 0 feedthrough
rlabel pdiffusion 444 -237 444 -237 0 cellNo=591
rlabel pdiffusion 451 -237 451 -237 0 cellNo=132
rlabel pdiffusion 458 -237 458 -237 0 feedthrough
rlabel pdiffusion 465 -237 465 -237 0 feedthrough
rlabel pdiffusion 472 -237 472 -237 0 feedthrough
rlabel pdiffusion 479 -237 479 -237 0 cellNo=228
rlabel pdiffusion 486 -237 486 -237 0 cellNo=424
rlabel pdiffusion 493 -237 493 -237 0 feedthrough
rlabel pdiffusion 500 -237 500 -237 0 cellNo=973
rlabel pdiffusion 507 -237 507 -237 0 feedthrough
rlabel pdiffusion 514 -237 514 -237 0 feedthrough
rlabel pdiffusion 521 -237 521 -237 0 feedthrough
rlabel pdiffusion 528 -237 528 -237 0 feedthrough
rlabel pdiffusion 535 -237 535 -237 0 feedthrough
rlabel pdiffusion 542 -237 542 -237 0 feedthrough
rlabel pdiffusion 549 -237 549 -237 0 cellNo=569
rlabel pdiffusion 556 -237 556 -237 0 feedthrough
rlabel pdiffusion 563 -237 563 -237 0 feedthrough
rlabel pdiffusion 570 -237 570 -237 0 feedthrough
rlabel pdiffusion 577 -237 577 -237 0 feedthrough
rlabel pdiffusion 584 -237 584 -237 0 feedthrough
rlabel pdiffusion 591 -237 591 -237 0 feedthrough
rlabel pdiffusion 598 -237 598 -237 0 feedthrough
rlabel pdiffusion 605 -237 605 -237 0 feedthrough
rlabel pdiffusion 612 -237 612 -237 0 cellNo=149
rlabel pdiffusion 619 -237 619 -237 0 feedthrough
rlabel pdiffusion 626 -237 626 -237 0 cellNo=804
rlabel pdiffusion 633 -237 633 -237 0 feedthrough
rlabel pdiffusion 640 -237 640 -237 0 feedthrough
rlabel pdiffusion 647 -237 647 -237 0 feedthrough
rlabel pdiffusion 654 -237 654 -237 0 feedthrough
rlabel pdiffusion 661 -237 661 -237 0 feedthrough
rlabel pdiffusion 668 -237 668 -237 0 feedthrough
rlabel pdiffusion 675 -237 675 -237 0 feedthrough
rlabel pdiffusion 682 -237 682 -237 0 feedthrough
rlabel pdiffusion 689 -237 689 -237 0 feedthrough
rlabel pdiffusion 696 -237 696 -237 0 feedthrough
rlabel pdiffusion 703 -237 703 -237 0 feedthrough
rlabel pdiffusion 710 -237 710 -237 0 feedthrough
rlabel pdiffusion 717 -237 717 -237 0 feedthrough
rlabel pdiffusion 724 -237 724 -237 0 feedthrough
rlabel pdiffusion 731 -237 731 -237 0 feedthrough
rlabel pdiffusion 738 -237 738 -237 0 feedthrough
rlabel pdiffusion 745 -237 745 -237 0 feedthrough
rlabel pdiffusion 752 -237 752 -237 0 cellNo=381
rlabel pdiffusion 759 -237 759 -237 0 feedthrough
rlabel pdiffusion 766 -237 766 -237 0 feedthrough
rlabel pdiffusion 773 -237 773 -237 0 feedthrough
rlabel pdiffusion 780 -237 780 -237 0 feedthrough
rlabel pdiffusion 787 -237 787 -237 0 feedthrough
rlabel pdiffusion 794 -237 794 -237 0 feedthrough
rlabel pdiffusion 801 -237 801 -237 0 feedthrough
rlabel pdiffusion 808 -237 808 -237 0 feedthrough
rlabel pdiffusion 815 -237 815 -237 0 feedthrough
rlabel pdiffusion 822 -237 822 -237 0 feedthrough
rlabel pdiffusion 829 -237 829 -237 0 cellNo=439
rlabel pdiffusion 836 -237 836 -237 0 feedthrough
rlabel pdiffusion 843 -237 843 -237 0 feedthrough
rlabel pdiffusion 850 -237 850 -237 0 cellNo=440
rlabel pdiffusion 857 -237 857 -237 0 feedthrough
rlabel pdiffusion 864 -237 864 -237 0 feedthrough
rlabel pdiffusion 871 -237 871 -237 0 feedthrough
rlabel pdiffusion 878 -237 878 -237 0 feedthrough
rlabel pdiffusion 885 -237 885 -237 0 feedthrough
rlabel pdiffusion 892 -237 892 -237 0 feedthrough
rlabel pdiffusion 899 -237 899 -237 0 feedthrough
rlabel pdiffusion 906 -237 906 -237 0 feedthrough
rlabel pdiffusion 913 -237 913 -237 0 feedthrough
rlabel pdiffusion 920 -237 920 -237 0 feedthrough
rlabel pdiffusion 927 -237 927 -237 0 feedthrough
rlabel pdiffusion 934 -237 934 -237 0 feedthrough
rlabel pdiffusion 941 -237 941 -237 0 feedthrough
rlabel pdiffusion 948 -237 948 -237 0 feedthrough
rlabel pdiffusion 955 -237 955 -237 0 feedthrough
rlabel pdiffusion 962 -237 962 -237 0 feedthrough
rlabel pdiffusion 969 -237 969 -237 0 feedthrough
rlabel pdiffusion 976 -237 976 -237 0 feedthrough
rlabel pdiffusion 983 -237 983 -237 0 feedthrough
rlabel pdiffusion 990 -237 990 -237 0 feedthrough
rlabel pdiffusion 997 -237 997 -237 0 feedthrough
rlabel pdiffusion 1004 -237 1004 -237 0 feedthrough
rlabel pdiffusion 1011 -237 1011 -237 0 feedthrough
rlabel pdiffusion 1018 -237 1018 -237 0 feedthrough
rlabel pdiffusion 1025 -237 1025 -237 0 feedthrough
rlabel pdiffusion 1039 -237 1039 -237 0 feedthrough
rlabel pdiffusion 1186 -237 1186 -237 0 feedthrough
rlabel pdiffusion 1326 -237 1326 -237 0 feedthrough
rlabel pdiffusion 3 -320 3 -320 0 cellNo=1013
rlabel pdiffusion 10 -320 10 -320 0 cellNo=1200
rlabel pdiffusion 17 -320 17 -320 0 cellNo=1048
rlabel pdiffusion 24 -320 24 -320 0 cellNo=1028
rlabel pdiffusion 31 -320 31 -320 0 cellNo=1198
rlabel pdiffusion 38 -320 38 -320 0 cellNo=1049
rlabel pdiffusion 45 -320 45 -320 0 cellNo=1063
rlabel pdiffusion 52 -320 52 -320 0 cellNo=1076
rlabel pdiffusion 59 -320 59 -320 0 cellNo=1095
rlabel pdiffusion 66 -320 66 -320 0 feedthrough
rlabel pdiffusion 73 -320 73 -320 0 cellNo=174
rlabel pdiffusion 80 -320 80 -320 0 feedthrough
rlabel pdiffusion 87 -320 87 -320 0 feedthrough
rlabel pdiffusion 94 -320 94 -320 0 feedthrough
rlabel pdiffusion 101 -320 101 -320 0 feedthrough
rlabel pdiffusion 108 -320 108 -320 0 feedthrough
rlabel pdiffusion 115 -320 115 -320 0 feedthrough
rlabel pdiffusion 122 -320 122 -320 0 feedthrough
rlabel pdiffusion 129 -320 129 -320 0 feedthrough
rlabel pdiffusion 136 -320 136 -320 0 cellNo=334
rlabel pdiffusion 143 -320 143 -320 0 cellNo=158
rlabel pdiffusion 150 -320 150 -320 0 feedthrough
rlabel pdiffusion 157 -320 157 -320 0 feedthrough
rlabel pdiffusion 164 -320 164 -320 0 feedthrough
rlabel pdiffusion 171 -320 171 -320 0 cellNo=46
rlabel pdiffusion 178 -320 178 -320 0 feedthrough
rlabel pdiffusion 185 -320 185 -320 0 cellNo=225
rlabel pdiffusion 192 -320 192 -320 0 feedthrough
rlabel pdiffusion 199 -320 199 -320 0 feedthrough
rlabel pdiffusion 206 -320 206 -320 0 cellNo=792
rlabel pdiffusion 213 -320 213 -320 0 feedthrough
rlabel pdiffusion 220 -320 220 -320 0 feedthrough
rlabel pdiffusion 227 -320 227 -320 0 feedthrough
rlabel pdiffusion 234 -320 234 -320 0 feedthrough
rlabel pdiffusion 241 -320 241 -320 0 feedthrough
rlabel pdiffusion 248 -320 248 -320 0 feedthrough
rlabel pdiffusion 255 -320 255 -320 0 feedthrough
rlabel pdiffusion 262 -320 262 -320 0 feedthrough
rlabel pdiffusion 269 -320 269 -320 0 feedthrough
rlabel pdiffusion 276 -320 276 -320 0 feedthrough
rlabel pdiffusion 283 -320 283 -320 0 feedthrough
rlabel pdiffusion 290 -320 290 -320 0 feedthrough
rlabel pdiffusion 297 -320 297 -320 0 feedthrough
rlabel pdiffusion 304 -320 304 -320 0 feedthrough
rlabel pdiffusion 311 -320 311 -320 0 cellNo=637
rlabel pdiffusion 318 -320 318 -320 0 feedthrough
rlabel pdiffusion 325 -320 325 -320 0 feedthrough
rlabel pdiffusion 332 -320 332 -320 0 feedthrough
rlabel pdiffusion 339 -320 339 -320 0 feedthrough
rlabel pdiffusion 346 -320 346 -320 0 feedthrough
rlabel pdiffusion 353 -320 353 -320 0 feedthrough
rlabel pdiffusion 360 -320 360 -320 0 feedthrough
rlabel pdiffusion 367 -320 367 -320 0 feedthrough
rlabel pdiffusion 374 -320 374 -320 0 cellNo=587
rlabel pdiffusion 381 -320 381 -320 0 cellNo=992
rlabel pdiffusion 388 -320 388 -320 0 cellNo=217
rlabel pdiffusion 395 -320 395 -320 0 feedthrough
rlabel pdiffusion 402 -320 402 -320 0 feedthrough
rlabel pdiffusion 409 -320 409 -320 0 feedthrough
rlabel pdiffusion 416 -320 416 -320 0 feedthrough
rlabel pdiffusion 423 -320 423 -320 0 feedthrough
rlabel pdiffusion 430 -320 430 -320 0 feedthrough
rlabel pdiffusion 437 -320 437 -320 0 feedthrough
rlabel pdiffusion 444 -320 444 -320 0 cellNo=170
rlabel pdiffusion 451 -320 451 -320 0 feedthrough
rlabel pdiffusion 458 -320 458 -320 0 feedthrough
rlabel pdiffusion 465 -320 465 -320 0 feedthrough
rlabel pdiffusion 472 -320 472 -320 0 feedthrough
rlabel pdiffusion 479 -320 479 -320 0 cellNo=326
rlabel pdiffusion 486 -320 486 -320 0 feedthrough
rlabel pdiffusion 493 -320 493 -320 0 feedthrough
rlabel pdiffusion 500 -320 500 -320 0 feedthrough
rlabel pdiffusion 507 -320 507 -320 0 feedthrough
rlabel pdiffusion 514 -320 514 -320 0 feedthrough
rlabel pdiffusion 521 -320 521 -320 0 feedthrough
rlabel pdiffusion 528 -320 528 -320 0 feedthrough
rlabel pdiffusion 535 -320 535 -320 0 cellNo=201
rlabel pdiffusion 542 -320 542 -320 0 feedthrough
rlabel pdiffusion 549 -320 549 -320 0 cellNo=509
rlabel pdiffusion 556 -320 556 -320 0 feedthrough
rlabel pdiffusion 563 -320 563 -320 0 feedthrough
rlabel pdiffusion 570 -320 570 -320 0 feedthrough
rlabel pdiffusion 577 -320 577 -320 0 feedthrough
rlabel pdiffusion 584 -320 584 -320 0 feedthrough
rlabel pdiffusion 591 -320 591 -320 0 cellNo=291
rlabel pdiffusion 598 -320 598 -320 0 cellNo=778
rlabel pdiffusion 605 -320 605 -320 0 cellNo=169
rlabel pdiffusion 612 -320 612 -320 0 feedthrough
rlabel pdiffusion 619 -320 619 -320 0 feedthrough
rlabel pdiffusion 626 -320 626 -320 0 cellNo=261
rlabel pdiffusion 633 -320 633 -320 0 feedthrough
rlabel pdiffusion 640 -320 640 -320 0 feedthrough
rlabel pdiffusion 647 -320 647 -320 0 cellNo=699
rlabel pdiffusion 654 -320 654 -320 0 feedthrough
rlabel pdiffusion 661 -320 661 -320 0 feedthrough
rlabel pdiffusion 668 -320 668 -320 0 cellNo=330
rlabel pdiffusion 675 -320 675 -320 0 feedthrough
rlabel pdiffusion 682 -320 682 -320 0 feedthrough
rlabel pdiffusion 689 -320 689 -320 0 feedthrough
rlabel pdiffusion 696 -320 696 -320 0 cellNo=978
rlabel pdiffusion 703 -320 703 -320 0 feedthrough
rlabel pdiffusion 710 -320 710 -320 0 feedthrough
rlabel pdiffusion 717 -320 717 -320 0 feedthrough
rlabel pdiffusion 724 -320 724 -320 0 feedthrough
rlabel pdiffusion 731 -320 731 -320 0 feedthrough
rlabel pdiffusion 738 -320 738 -320 0 feedthrough
rlabel pdiffusion 745 -320 745 -320 0 cellNo=219
rlabel pdiffusion 752 -320 752 -320 0 feedthrough
rlabel pdiffusion 759 -320 759 -320 0 feedthrough
rlabel pdiffusion 766 -320 766 -320 0 feedthrough
rlabel pdiffusion 773 -320 773 -320 0 feedthrough
rlabel pdiffusion 780 -320 780 -320 0 feedthrough
rlabel pdiffusion 787 -320 787 -320 0 feedthrough
rlabel pdiffusion 794 -320 794 -320 0 feedthrough
rlabel pdiffusion 801 -320 801 -320 0 feedthrough
rlabel pdiffusion 808 -320 808 -320 0 feedthrough
rlabel pdiffusion 815 -320 815 -320 0 feedthrough
rlabel pdiffusion 822 -320 822 -320 0 feedthrough
rlabel pdiffusion 829 -320 829 -320 0 feedthrough
rlabel pdiffusion 836 -320 836 -320 0 feedthrough
rlabel pdiffusion 843 -320 843 -320 0 feedthrough
rlabel pdiffusion 850 -320 850 -320 0 feedthrough
rlabel pdiffusion 857 -320 857 -320 0 feedthrough
rlabel pdiffusion 864 -320 864 -320 0 feedthrough
rlabel pdiffusion 871 -320 871 -320 0 feedthrough
rlabel pdiffusion 878 -320 878 -320 0 feedthrough
rlabel pdiffusion 885 -320 885 -320 0 feedthrough
rlabel pdiffusion 892 -320 892 -320 0 feedthrough
rlabel pdiffusion 899 -320 899 -320 0 feedthrough
rlabel pdiffusion 906 -320 906 -320 0 feedthrough
rlabel pdiffusion 913 -320 913 -320 0 feedthrough
rlabel pdiffusion 920 -320 920 -320 0 feedthrough
rlabel pdiffusion 927 -320 927 -320 0 feedthrough
rlabel pdiffusion 934 -320 934 -320 0 feedthrough
rlabel pdiffusion 941 -320 941 -320 0 feedthrough
rlabel pdiffusion 948 -320 948 -320 0 feedthrough
rlabel pdiffusion 955 -320 955 -320 0 feedthrough
rlabel pdiffusion 962 -320 962 -320 0 feedthrough
rlabel pdiffusion 969 -320 969 -320 0 feedthrough
rlabel pdiffusion 976 -320 976 -320 0 feedthrough
rlabel pdiffusion 983 -320 983 -320 0 feedthrough
rlabel pdiffusion 990 -320 990 -320 0 feedthrough
rlabel pdiffusion 997 -320 997 -320 0 feedthrough
rlabel pdiffusion 1004 -320 1004 -320 0 feedthrough
rlabel pdiffusion 1011 -320 1011 -320 0 feedthrough
rlabel pdiffusion 1018 -320 1018 -320 0 feedthrough
rlabel pdiffusion 1025 -320 1025 -320 0 feedthrough
rlabel pdiffusion 1032 -320 1032 -320 0 feedthrough
rlabel pdiffusion 1039 -320 1039 -320 0 feedthrough
rlabel pdiffusion 1046 -320 1046 -320 0 feedthrough
rlabel pdiffusion 1053 -320 1053 -320 0 feedthrough
rlabel pdiffusion 1060 -320 1060 -320 0 feedthrough
rlabel pdiffusion 1067 -320 1067 -320 0 feedthrough
rlabel pdiffusion 1074 -320 1074 -320 0 feedthrough
rlabel pdiffusion 1081 -320 1081 -320 0 feedthrough
rlabel pdiffusion 1088 -320 1088 -320 0 feedthrough
rlabel pdiffusion 1095 -320 1095 -320 0 feedthrough
rlabel pdiffusion 1102 -320 1102 -320 0 feedthrough
rlabel pdiffusion 1109 -320 1109 -320 0 feedthrough
rlabel pdiffusion 1116 -320 1116 -320 0 feedthrough
rlabel pdiffusion 1123 -320 1123 -320 0 feedthrough
rlabel pdiffusion 1207 -320 1207 -320 0 feedthrough
rlabel pdiffusion 1305 -320 1305 -320 0 cellNo=336
rlabel pdiffusion 1382 -320 1382 -320 0 feedthrough
rlabel pdiffusion 1459 -320 1459 -320 0 feedthrough
rlabel pdiffusion 3 -419 3 -419 0 cellNo=1011
rlabel pdiffusion 10 -419 10 -419 0 cellNo=1022
rlabel pdiffusion 17 -419 17 -419 0 cellNo=1100
rlabel pdiffusion 24 -419 24 -419 0 cellNo=1037
rlabel pdiffusion 31 -419 31 -419 0 cellNo=1047
rlabel pdiffusion 38 -419 38 -419 0 cellNo=1061
rlabel pdiffusion 45 -419 45 -419 0 cellNo=1074
rlabel pdiffusion 52 -419 52 -419 0 cellNo=1093
rlabel pdiffusion 59 -419 59 -419 0 cellNo=140
rlabel pdiffusion 66 -419 66 -419 0 cellNo=1156
rlabel pdiffusion 73 -419 73 -419 0 feedthrough
rlabel pdiffusion 80 -419 80 -419 0 feedthrough
rlabel pdiffusion 87 -419 87 -419 0 feedthrough
rlabel pdiffusion 94 -419 94 -419 0 feedthrough
rlabel pdiffusion 101 -419 101 -419 0 feedthrough
rlabel pdiffusion 108 -419 108 -419 0 feedthrough
rlabel pdiffusion 115 -419 115 -419 0 feedthrough
rlabel pdiffusion 122 -419 122 -419 0 feedthrough
rlabel pdiffusion 129 -419 129 -419 0 feedthrough
rlabel pdiffusion 136 -419 136 -419 0 feedthrough
rlabel pdiffusion 143 -419 143 -419 0 feedthrough
rlabel pdiffusion 150 -419 150 -419 0 cellNo=507
rlabel pdiffusion 157 -419 157 -419 0 feedthrough
rlabel pdiffusion 164 -419 164 -419 0 cellNo=167
rlabel pdiffusion 171 -419 171 -419 0 cellNo=407
rlabel pdiffusion 178 -419 178 -419 0 feedthrough
rlabel pdiffusion 185 -419 185 -419 0 cellNo=348
rlabel pdiffusion 192 -419 192 -419 0 cellNo=362
rlabel pdiffusion 199 -419 199 -419 0 feedthrough
rlabel pdiffusion 206 -419 206 -419 0 feedthrough
rlabel pdiffusion 213 -419 213 -419 0 feedthrough
rlabel pdiffusion 220 -419 220 -419 0 feedthrough
rlabel pdiffusion 227 -419 227 -419 0 feedthrough
rlabel pdiffusion 234 -419 234 -419 0 feedthrough
rlabel pdiffusion 241 -419 241 -419 0 feedthrough
rlabel pdiffusion 248 -419 248 -419 0 cellNo=277
rlabel pdiffusion 255 -419 255 -419 0 feedthrough
rlabel pdiffusion 262 -419 262 -419 0 feedthrough
rlabel pdiffusion 269 -419 269 -419 0 feedthrough
rlabel pdiffusion 276 -419 276 -419 0 feedthrough
rlabel pdiffusion 283 -419 283 -419 0 feedthrough
rlabel pdiffusion 290 -419 290 -419 0 feedthrough
rlabel pdiffusion 297 -419 297 -419 0 feedthrough
rlabel pdiffusion 304 -419 304 -419 0 feedthrough
rlabel pdiffusion 311 -419 311 -419 0 feedthrough
rlabel pdiffusion 318 -419 318 -419 0 feedthrough
rlabel pdiffusion 325 -419 325 -419 0 feedthrough
rlabel pdiffusion 332 -419 332 -419 0 feedthrough
rlabel pdiffusion 339 -419 339 -419 0 feedthrough
rlabel pdiffusion 346 -419 346 -419 0 feedthrough
rlabel pdiffusion 353 -419 353 -419 0 feedthrough
rlabel pdiffusion 360 -419 360 -419 0 cellNo=249
rlabel pdiffusion 367 -419 367 -419 0 cellNo=457
rlabel pdiffusion 374 -419 374 -419 0 feedthrough
rlabel pdiffusion 381 -419 381 -419 0 cellNo=69
rlabel pdiffusion 388 -419 388 -419 0 feedthrough
rlabel pdiffusion 395 -419 395 -419 0 feedthrough
rlabel pdiffusion 402 -419 402 -419 0 feedthrough
rlabel pdiffusion 409 -419 409 -419 0 feedthrough
rlabel pdiffusion 416 -419 416 -419 0 cellNo=71
rlabel pdiffusion 423 -419 423 -419 0 feedthrough
rlabel pdiffusion 430 -419 430 -419 0 feedthrough
rlabel pdiffusion 437 -419 437 -419 0 feedthrough
rlabel pdiffusion 444 -419 444 -419 0 feedthrough
rlabel pdiffusion 451 -419 451 -419 0 feedthrough
rlabel pdiffusion 458 -419 458 -419 0 feedthrough
rlabel pdiffusion 465 -419 465 -419 0 feedthrough
rlabel pdiffusion 472 -419 472 -419 0 feedthrough
rlabel pdiffusion 479 -419 479 -419 0 feedthrough
rlabel pdiffusion 486 -419 486 -419 0 feedthrough
rlabel pdiffusion 493 -419 493 -419 0 cellNo=322
rlabel pdiffusion 500 -419 500 -419 0 feedthrough
rlabel pdiffusion 507 -419 507 -419 0 feedthrough
rlabel pdiffusion 514 -419 514 -419 0 feedthrough
rlabel pdiffusion 521 -419 521 -419 0 feedthrough
rlabel pdiffusion 528 -419 528 -419 0 feedthrough
rlabel pdiffusion 535 -419 535 -419 0 feedthrough
rlabel pdiffusion 542 -419 542 -419 0 cellNo=931
rlabel pdiffusion 549 -419 549 -419 0 feedthrough
rlabel pdiffusion 556 -419 556 -419 0 feedthrough
rlabel pdiffusion 563 -419 563 -419 0 cellNo=22
rlabel pdiffusion 570 -419 570 -419 0 cellNo=741
rlabel pdiffusion 577 -419 577 -419 0 feedthrough
rlabel pdiffusion 584 -419 584 -419 0 cellNo=783
rlabel pdiffusion 591 -419 591 -419 0 feedthrough
rlabel pdiffusion 598 -419 598 -419 0 feedthrough
rlabel pdiffusion 605 -419 605 -419 0 feedthrough
rlabel pdiffusion 612 -419 612 -419 0 feedthrough
rlabel pdiffusion 619 -419 619 -419 0 feedthrough
rlabel pdiffusion 626 -419 626 -419 0 cellNo=677
rlabel pdiffusion 633 -419 633 -419 0 cellNo=952
rlabel pdiffusion 640 -419 640 -419 0 feedthrough
rlabel pdiffusion 647 -419 647 -419 0 feedthrough
rlabel pdiffusion 654 -419 654 -419 0 feedthrough
rlabel pdiffusion 661 -419 661 -419 0 feedthrough
rlabel pdiffusion 668 -419 668 -419 0 feedthrough
rlabel pdiffusion 675 -419 675 -419 0 feedthrough
rlabel pdiffusion 682 -419 682 -419 0 feedthrough
rlabel pdiffusion 689 -419 689 -419 0 cellNo=863
rlabel pdiffusion 696 -419 696 -419 0 feedthrough
rlabel pdiffusion 703 -419 703 -419 0 feedthrough
rlabel pdiffusion 710 -419 710 -419 0 feedthrough
rlabel pdiffusion 717 -419 717 -419 0 cellNo=789
rlabel pdiffusion 724 -419 724 -419 0 cellNo=835
rlabel pdiffusion 731 -419 731 -419 0 feedthrough
rlabel pdiffusion 738 -419 738 -419 0 feedthrough
rlabel pdiffusion 745 -419 745 -419 0 feedthrough
rlabel pdiffusion 752 -419 752 -419 0 feedthrough
rlabel pdiffusion 759 -419 759 -419 0 feedthrough
rlabel pdiffusion 766 -419 766 -419 0 feedthrough
rlabel pdiffusion 773 -419 773 -419 0 feedthrough
rlabel pdiffusion 780 -419 780 -419 0 feedthrough
rlabel pdiffusion 787 -419 787 -419 0 cellNo=817
rlabel pdiffusion 794 -419 794 -419 0 feedthrough
rlabel pdiffusion 801 -419 801 -419 0 feedthrough
rlabel pdiffusion 808 -419 808 -419 0 feedthrough
rlabel pdiffusion 815 -419 815 -419 0 feedthrough
rlabel pdiffusion 822 -419 822 -419 0 feedthrough
rlabel pdiffusion 829 -419 829 -419 0 feedthrough
rlabel pdiffusion 836 -419 836 -419 0 cellNo=458
rlabel pdiffusion 843 -419 843 -419 0 feedthrough
rlabel pdiffusion 850 -419 850 -419 0 feedthrough
rlabel pdiffusion 857 -419 857 -419 0 feedthrough
rlabel pdiffusion 864 -419 864 -419 0 feedthrough
rlabel pdiffusion 871 -419 871 -419 0 feedthrough
rlabel pdiffusion 878 -419 878 -419 0 feedthrough
rlabel pdiffusion 885 -419 885 -419 0 feedthrough
rlabel pdiffusion 892 -419 892 -419 0 feedthrough
rlabel pdiffusion 899 -419 899 -419 0 feedthrough
rlabel pdiffusion 906 -419 906 -419 0 feedthrough
rlabel pdiffusion 913 -419 913 -419 0 feedthrough
rlabel pdiffusion 920 -419 920 -419 0 feedthrough
rlabel pdiffusion 927 -419 927 -419 0 feedthrough
rlabel pdiffusion 934 -419 934 -419 0 feedthrough
rlabel pdiffusion 941 -419 941 -419 0 feedthrough
rlabel pdiffusion 948 -419 948 -419 0 feedthrough
rlabel pdiffusion 955 -419 955 -419 0 feedthrough
rlabel pdiffusion 962 -419 962 -419 0 feedthrough
rlabel pdiffusion 969 -419 969 -419 0 feedthrough
rlabel pdiffusion 976 -419 976 -419 0 feedthrough
rlabel pdiffusion 983 -419 983 -419 0 feedthrough
rlabel pdiffusion 990 -419 990 -419 0 feedthrough
rlabel pdiffusion 997 -419 997 -419 0 feedthrough
rlabel pdiffusion 1004 -419 1004 -419 0 feedthrough
rlabel pdiffusion 1011 -419 1011 -419 0 feedthrough
rlabel pdiffusion 1018 -419 1018 -419 0 feedthrough
rlabel pdiffusion 1025 -419 1025 -419 0 feedthrough
rlabel pdiffusion 1032 -419 1032 -419 0 feedthrough
rlabel pdiffusion 1039 -419 1039 -419 0 feedthrough
rlabel pdiffusion 1046 -419 1046 -419 0 feedthrough
rlabel pdiffusion 1053 -419 1053 -419 0 feedthrough
rlabel pdiffusion 1060 -419 1060 -419 0 feedthrough
rlabel pdiffusion 1067 -419 1067 -419 0 feedthrough
rlabel pdiffusion 1074 -419 1074 -419 0 feedthrough
rlabel pdiffusion 1081 -419 1081 -419 0 feedthrough
rlabel pdiffusion 1088 -419 1088 -419 0 feedthrough
rlabel pdiffusion 1095 -419 1095 -419 0 feedthrough
rlabel pdiffusion 1102 -419 1102 -419 0 feedthrough
rlabel pdiffusion 1109 -419 1109 -419 0 feedthrough
rlabel pdiffusion 1116 -419 1116 -419 0 feedthrough
rlabel pdiffusion 1123 -419 1123 -419 0 feedthrough
rlabel pdiffusion 1130 -419 1130 -419 0 feedthrough
rlabel pdiffusion 1137 -419 1137 -419 0 feedthrough
rlabel pdiffusion 1144 -419 1144 -419 0 feedthrough
rlabel pdiffusion 1151 -419 1151 -419 0 feedthrough
rlabel pdiffusion 1158 -419 1158 -419 0 feedthrough
rlabel pdiffusion 1165 -419 1165 -419 0 feedthrough
rlabel pdiffusion 1172 -419 1172 -419 0 feedthrough
rlabel pdiffusion 1179 -419 1179 -419 0 feedthrough
rlabel pdiffusion 1186 -419 1186 -419 0 feedthrough
rlabel pdiffusion 1193 -419 1193 -419 0 feedthrough
rlabel pdiffusion 1200 -419 1200 -419 0 feedthrough
rlabel pdiffusion 1207 -419 1207 -419 0 feedthrough
rlabel pdiffusion 1214 -419 1214 -419 0 feedthrough
rlabel pdiffusion 1221 -419 1221 -419 0 cellNo=215
rlabel pdiffusion 1389 -419 1389 -419 0 feedthrough
rlabel pdiffusion 1410 -419 1410 -419 0 feedthrough
rlabel pdiffusion 1522 -419 1522 -419 0 feedthrough
rlabel pdiffusion 3 -508 3 -508 0 cellNo=1021
rlabel pdiffusion 10 -508 10 -508 0 cellNo=1027
rlabel pdiffusion 17 -508 17 -508 0 cellNo=1035
rlabel pdiffusion 24 -508 24 -508 0 cellNo=1045
rlabel pdiffusion 31 -508 31 -508 0 cellNo=1060
rlabel pdiffusion 38 -508 38 -508 0 cellNo=1073
rlabel pdiffusion 45 -508 45 -508 0 cellNo=1092
rlabel pdiffusion 52 -508 52 -508 0 feedthrough
rlabel pdiffusion 59 -508 59 -508 0 feedthrough
rlabel pdiffusion 66 -508 66 -508 0 feedthrough
rlabel pdiffusion 73 -508 73 -508 0 feedthrough
rlabel pdiffusion 80 -508 80 -508 0 feedthrough
rlabel pdiffusion 87 -508 87 -508 0 feedthrough
rlabel pdiffusion 94 -508 94 -508 0 feedthrough
rlabel pdiffusion 101 -508 101 -508 0 feedthrough
rlabel pdiffusion 108 -508 108 -508 0 feedthrough
rlabel pdiffusion 115 -508 115 -508 0 feedthrough
rlabel pdiffusion 122 -508 122 -508 0 cellNo=493
rlabel pdiffusion 129 -508 129 -508 0 feedthrough
rlabel pdiffusion 136 -508 136 -508 0 cellNo=189
rlabel pdiffusion 143 -508 143 -508 0 cellNo=216
rlabel pdiffusion 150 -508 150 -508 0 feedthrough
rlabel pdiffusion 157 -508 157 -508 0 feedthrough
rlabel pdiffusion 164 -508 164 -508 0 cellNo=639
rlabel pdiffusion 171 -508 171 -508 0 feedthrough
rlabel pdiffusion 178 -508 178 -508 0 feedthrough
rlabel pdiffusion 185 -508 185 -508 0 feedthrough
rlabel pdiffusion 192 -508 192 -508 0 cellNo=208
rlabel pdiffusion 199 -508 199 -508 0 feedthrough
rlabel pdiffusion 206 -508 206 -508 0 feedthrough
rlabel pdiffusion 213 -508 213 -508 0 feedthrough
rlabel pdiffusion 220 -508 220 -508 0 feedthrough
rlabel pdiffusion 227 -508 227 -508 0 feedthrough
rlabel pdiffusion 234 -508 234 -508 0 cellNo=671
rlabel pdiffusion 241 -508 241 -508 0 feedthrough
rlabel pdiffusion 248 -508 248 -508 0 feedthrough
rlabel pdiffusion 255 -508 255 -508 0 cellNo=29
rlabel pdiffusion 262 -508 262 -508 0 feedthrough
rlabel pdiffusion 269 -508 269 -508 0 feedthrough
rlabel pdiffusion 276 -508 276 -508 0 feedthrough
rlabel pdiffusion 283 -508 283 -508 0 feedthrough
rlabel pdiffusion 290 -508 290 -508 0 feedthrough
rlabel pdiffusion 297 -508 297 -508 0 cellNo=750
rlabel pdiffusion 304 -508 304 -508 0 feedthrough
rlabel pdiffusion 311 -508 311 -508 0 feedthrough
rlabel pdiffusion 318 -508 318 -508 0 feedthrough
rlabel pdiffusion 325 -508 325 -508 0 feedthrough
rlabel pdiffusion 332 -508 332 -508 0 feedthrough
rlabel pdiffusion 339 -508 339 -508 0 feedthrough
rlabel pdiffusion 346 -508 346 -508 0 feedthrough
rlabel pdiffusion 353 -508 353 -508 0 feedthrough
rlabel pdiffusion 360 -508 360 -508 0 feedthrough
rlabel pdiffusion 367 -508 367 -508 0 feedthrough
rlabel pdiffusion 374 -508 374 -508 0 feedthrough
rlabel pdiffusion 381 -508 381 -508 0 feedthrough
rlabel pdiffusion 388 -508 388 -508 0 cellNo=560
rlabel pdiffusion 395 -508 395 -508 0 feedthrough
rlabel pdiffusion 402 -508 402 -508 0 cellNo=500
rlabel pdiffusion 409 -508 409 -508 0 feedthrough
rlabel pdiffusion 416 -508 416 -508 0 feedthrough
rlabel pdiffusion 423 -508 423 -508 0 cellNo=236
rlabel pdiffusion 430 -508 430 -508 0 feedthrough
rlabel pdiffusion 437 -508 437 -508 0 feedthrough
rlabel pdiffusion 444 -508 444 -508 0 feedthrough
rlabel pdiffusion 451 -508 451 -508 0 feedthrough
rlabel pdiffusion 458 -508 458 -508 0 feedthrough
rlabel pdiffusion 465 -508 465 -508 0 cellNo=657
rlabel pdiffusion 472 -508 472 -508 0 feedthrough
rlabel pdiffusion 479 -508 479 -508 0 feedthrough
rlabel pdiffusion 486 -508 486 -508 0 feedthrough
rlabel pdiffusion 493 -508 493 -508 0 feedthrough
rlabel pdiffusion 500 -508 500 -508 0 feedthrough
rlabel pdiffusion 507 -508 507 -508 0 feedthrough
rlabel pdiffusion 514 -508 514 -508 0 feedthrough
rlabel pdiffusion 521 -508 521 -508 0 feedthrough
rlabel pdiffusion 528 -508 528 -508 0 feedthrough
rlabel pdiffusion 535 -508 535 -508 0 feedthrough
rlabel pdiffusion 542 -508 542 -508 0 feedthrough
rlabel pdiffusion 549 -508 549 -508 0 cellNo=412
rlabel pdiffusion 556 -508 556 -508 0 cellNo=16
rlabel pdiffusion 563 -508 563 -508 0 feedthrough
rlabel pdiffusion 570 -508 570 -508 0 feedthrough
rlabel pdiffusion 577 -508 577 -508 0 feedthrough
rlabel pdiffusion 584 -508 584 -508 0 feedthrough
rlabel pdiffusion 591 -508 591 -508 0 cellNo=408
rlabel pdiffusion 598 -508 598 -508 0 feedthrough
rlabel pdiffusion 605 -508 605 -508 0 feedthrough
rlabel pdiffusion 612 -508 612 -508 0 feedthrough
rlabel pdiffusion 619 -508 619 -508 0 cellNo=205
rlabel pdiffusion 626 -508 626 -508 0 feedthrough
rlabel pdiffusion 633 -508 633 -508 0 feedthrough
rlabel pdiffusion 640 -508 640 -508 0 feedthrough
rlabel pdiffusion 647 -508 647 -508 0 cellNo=779
rlabel pdiffusion 654 -508 654 -508 0 cellNo=879
rlabel pdiffusion 661 -508 661 -508 0 cellNo=818
rlabel pdiffusion 668 -508 668 -508 0 feedthrough
rlabel pdiffusion 675 -508 675 -508 0 feedthrough
rlabel pdiffusion 682 -508 682 -508 0 cellNo=739
rlabel pdiffusion 689 -508 689 -508 0 feedthrough
rlabel pdiffusion 696 -508 696 -508 0 cellNo=802
rlabel pdiffusion 703 -508 703 -508 0 feedthrough
rlabel pdiffusion 710 -508 710 -508 0 feedthrough
rlabel pdiffusion 717 -508 717 -508 0 feedthrough
rlabel pdiffusion 724 -508 724 -508 0 feedthrough
rlabel pdiffusion 731 -508 731 -508 0 feedthrough
rlabel pdiffusion 738 -508 738 -508 0 feedthrough
rlabel pdiffusion 745 -508 745 -508 0 feedthrough
rlabel pdiffusion 752 -508 752 -508 0 cellNo=173
rlabel pdiffusion 759 -508 759 -508 0 feedthrough
rlabel pdiffusion 766 -508 766 -508 0 feedthrough
rlabel pdiffusion 773 -508 773 -508 0 feedthrough
rlabel pdiffusion 780 -508 780 -508 0 feedthrough
rlabel pdiffusion 787 -508 787 -508 0 feedthrough
rlabel pdiffusion 794 -508 794 -508 0 feedthrough
rlabel pdiffusion 801 -508 801 -508 0 feedthrough
rlabel pdiffusion 808 -508 808 -508 0 feedthrough
rlabel pdiffusion 815 -508 815 -508 0 feedthrough
rlabel pdiffusion 822 -508 822 -508 0 cellNo=283
rlabel pdiffusion 829 -508 829 -508 0 feedthrough
rlabel pdiffusion 836 -508 836 -508 0 feedthrough
rlabel pdiffusion 843 -508 843 -508 0 cellNo=428
rlabel pdiffusion 850 -508 850 -508 0 cellNo=360
rlabel pdiffusion 857 -508 857 -508 0 feedthrough
rlabel pdiffusion 864 -508 864 -508 0 feedthrough
rlabel pdiffusion 871 -508 871 -508 0 feedthrough
rlabel pdiffusion 878 -508 878 -508 0 feedthrough
rlabel pdiffusion 885 -508 885 -508 0 feedthrough
rlabel pdiffusion 892 -508 892 -508 0 feedthrough
rlabel pdiffusion 899 -508 899 -508 0 feedthrough
rlabel pdiffusion 906 -508 906 -508 0 feedthrough
rlabel pdiffusion 913 -508 913 -508 0 feedthrough
rlabel pdiffusion 920 -508 920 -508 0 feedthrough
rlabel pdiffusion 927 -508 927 -508 0 feedthrough
rlabel pdiffusion 934 -508 934 -508 0 feedthrough
rlabel pdiffusion 941 -508 941 -508 0 feedthrough
rlabel pdiffusion 948 -508 948 -508 0 feedthrough
rlabel pdiffusion 955 -508 955 -508 0 feedthrough
rlabel pdiffusion 962 -508 962 -508 0 feedthrough
rlabel pdiffusion 969 -508 969 -508 0 feedthrough
rlabel pdiffusion 976 -508 976 -508 0 feedthrough
rlabel pdiffusion 983 -508 983 -508 0 feedthrough
rlabel pdiffusion 990 -508 990 -508 0 feedthrough
rlabel pdiffusion 997 -508 997 -508 0 feedthrough
rlabel pdiffusion 1004 -508 1004 -508 0 feedthrough
rlabel pdiffusion 1011 -508 1011 -508 0 feedthrough
rlabel pdiffusion 1018 -508 1018 -508 0 feedthrough
rlabel pdiffusion 1025 -508 1025 -508 0 feedthrough
rlabel pdiffusion 1032 -508 1032 -508 0 feedthrough
rlabel pdiffusion 1039 -508 1039 -508 0 feedthrough
rlabel pdiffusion 1046 -508 1046 -508 0 feedthrough
rlabel pdiffusion 1053 -508 1053 -508 0 feedthrough
rlabel pdiffusion 1060 -508 1060 -508 0 feedthrough
rlabel pdiffusion 1067 -508 1067 -508 0 feedthrough
rlabel pdiffusion 1074 -508 1074 -508 0 feedthrough
rlabel pdiffusion 1081 -508 1081 -508 0 feedthrough
rlabel pdiffusion 1088 -508 1088 -508 0 feedthrough
rlabel pdiffusion 1095 -508 1095 -508 0 feedthrough
rlabel pdiffusion 1102 -508 1102 -508 0 feedthrough
rlabel pdiffusion 1109 -508 1109 -508 0 feedthrough
rlabel pdiffusion 1116 -508 1116 -508 0 feedthrough
rlabel pdiffusion 1123 -508 1123 -508 0 feedthrough
rlabel pdiffusion 1130 -508 1130 -508 0 feedthrough
rlabel pdiffusion 1137 -508 1137 -508 0 feedthrough
rlabel pdiffusion 1144 -508 1144 -508 0 feedthrough
rlabel pdiffusion 1151 -508 1151 -508 0 feedthrough
rlabel pdiffusion 1158 -508 1158 -508 0 feedthrough
rlabel pdiffusion 1165 -508 1165 -508 0 feedthrough
rlabel pdiffusion 1172 -508 1172 -508 0 feedthrough
rlabel pdiffusion 1179 -508 1179 -508 0 feedthrough
rlabel pdiffusion 1186 -508 1186 -508 0 feedthrough
rlabel pdiffusion 1193 -508 1193 -508 0 feedthrough
rlabel pdiffusion 1200 -508 1200 -508 0 feedthrough
rlabel pdiffusion 1207 -508 1207 -508 0 feedthrough
rlabel pdiffusion 1214 -508 1214 -508 0 feedthrough
rlabel pdiffusion 1221 -508 1221 -508 0 cellNo=465
rlabel pdiffusion 1228 -508 1228 -508 0 feedthrough
rlabel pdiffusion 1235 -508 1235 -508 0 feedthrough
rlabel pdiffusion 1242 -508 1242 -508 0 feedthrough
rlabel pdiffusion 1249 -508 1249 -508 0 cellNo=196
rlabel pdiffusion 1256 -508 1256 -508 0 feedthrough
rlabel pdiffusion 1431 -508 1431 -508 0 feedthrough
rlabel pdiffusion 1487 -508 1487 -508 0 feedthrough
rlabel pdiffusion 1543 -508 1543 -508 0 feedthrough
rlabel pdiffusion 3 -629 3 -629 0 cellNo=1034
rlabel pdiffusion 10 -629 10 -629 0 cellNo=1155
rlabel pdiffusion 17 -629 17 -629 0 cellNo=1044
rlabel pdiffusion 24 -629 24 -629 0 cellNo=1059
rlabel pdiffusion 31 -629 31 -629 0 cellNo=1072
rlabel pdiffusion 38 -629 38 -629 0 cellNo=1091
rlabel pdiffusion 45 -629 45 -629 0 feedthrough
rlabel pdiffusion 52 -629 52 -629 0 feedthrough
rlabel pdiffusion 59 -629 59 -629 0 feedthrough
rlabel pdiffusion 66 -629 66 -629 0 feedthrough
rlabel pdiffusion 73 -629 73 -629 0 feedthrough
rlabel pdiffusion 80 -629 80 -629 0 cellNo=266
rlabel pdiffusion 87 -629 87 -629 0 feedthrough
rlabel pdiffusion 94 -629 94 -629 0 feedthrough
rlabel pdiffusion 101 -629 101 -629 0 feedthrough
rlabel pdiffusion 108 -629 108 -629 0 cellNo=252
rlabel pdiffusion 115 -629 115 -629 0 feedthrough
rlabel pdiffusion 122 -629 122 -629 0 feedthrough
rlabel pdiffusion 129 -629 129 -629 0 feedthrough
rlabel pdiffusion 136 -629 136 -629 0 feedthrough
rlabel pdiffusion 143 -629 143 -629 0 feedthrough
rlabel pdiffusion 150 -629 150 -629 0 feedthrough
rlabel pdiffusion 157 -629 157 -629 0 feedthrough
rlabel pdiffusion 164 -629 164 -629 0 feedthrough
rlabel pdiffusion 171 -629 171 -629 0 feedthrough
rlabel pdiffusion 178 -629 178 -629 0 feedthrough
rlabel pdiffusion 185 -629 185 -629 0 feedthrough
rlabel pdiffusion 192 -629 192 -629 0 feedthrough
rlabel pdiffusion 199 -629 199 -629 0 cellNo=738
rlabel pdiffusion 206 -629 206 -629 0 feedthrough
rlabel pdiffusion 213 -629 213 -629 0 feedthrough
rlabel pdiffusion 220 -629 220 -629 0 feedthrough
rlabel pdiffusion 227 -629 227 -629 0 feedthrough
rlabel pdiffusion 234 -629 234 -629 0 cellNo=193
rlabel pdiffusion 241 -629 241 -629 0 cellNo=864
rlabel pdiffusion 248 -629 248 -629 0 feedthrough
rlabel pdiffusion 255 -629 255 -629 0 feedthrough
rlabel pdiffusion 262 -629 262 -629 0 cellNo=496
rlabel pdiffusion 269 -629 269 -629 0 feedthrough
rlabel pdiffusion 276 -629 276 -629 0 feedthrough
rlabel pdiffusion 283 -629 283 -629 0 feedthrough
rlabel pdiffusion 290 -629 290 -629 0 cellNo=826
rlabel pdiffusion 297 -629 297 -629 0 feedthrough
rlabel pdiffusion 304 -629 304 -629 0 feedthrough
rlabel pdiffusion 311 -629 311 -629 0 feedthrough
rlabel pdiffusion 318 -629 318 -629 0 feedthrough
rlabel pdiffusion 325 -629 325 -629 0 cellNo=882
rlabel pdiffusion 332 -629 332 -629 0 feedthrough
rlabel pdiffusion 339 -629 339 -629 0 feedthrough
rlabel pdiffusion 346 -629 346 -629 0 feedthrough
rlabel pdiffusion 353 -629 353 -629 0 cellNo=100
rlabel pdiffusion 360 -629 360 -629 0 feedthrough
rlabel pdiffusion 367 -629 367 -629 0 feedthrough
rlabel pdiffusion 374 -629 374 -629 0 feedthrough
rlabel pdiffusion 381 -629 381 -629 0 feedthrough
rlabel pdiffusion 388 -629 388 -629 0 cellNo=551
rlabel pdiffusion 395 -629 395 -629 0 feedthrough
rlabel pdiffusion 402 -629 402 -629 0 feedthrough
rlabel pdiffusion 409 -629 409 -629 0 feedthrough
rlabel pdiffusion 416 -629 416 -629 0 feedthrough
rlabel pdiffusion 423 -629 423 -629 0 cellNo=449
rlabel pdiffusion 430 -629 430 -629 0 feedthrough
rlabel pdiffusion 437 -629 437 -629 0 feedthrough
rlabel pdiffusion 444 -629 444 -629 0 feedthrough
rlabel pdiffusion 451 -629 451 -629 0 feedthrough
rlabel pdiffusion 458 -629 458 -629 0 cellNo=112
rlabel pdiffusion 465 -629 465 -629 0 feedthrough
rlabel pdiffusion 472 -629 472 -629 0 feedthrough
rlabel pdiffusion 479 -629 479 -629 0 cellNo=666
rlabel pdiffusion 486 -629 486 -629 0 feedthrough
rlabel pdiffusion 493 -629 493 -629 0 cellNo=293
rlabel pdiffusion 500 -629 500 -629 0 feedthrough
rlabel pdiffusion 507 -629 507 -629 0 feedthrough
rlabel pdiffusion 514 -629 514 -629 0 feedthrough
rlabel pdiffusion 521 -629 521 -629 0 feedthrough
rlabel pdiffusion 528 -629 528 -629 0 feedthrough
rlabel pdiffusion 535 -629 535 -629 0 feedthrough
rlabel pdiffusion 542 -629 542 -629 0 feedthrough
rlabel pdiffusion 549 -629 549 -629 0 feedthrough
rlabel pdiffusion 556 -629 556 -629 0 feedthrough
rlabel pdiffusion 563 -629 563 -629 0 feedthrough
rlabel pdiffusion 570 -629 570 -629 0 feedthrough
rlabel pdiffusion 577 -629 577 -629 0 feedthrough
rlabel pdiffusion 584 -629 584 -629 0 feedthrough
rlabel pdiffusion 591 -629 591 -629 0 feedthrough
rlabel pdiffusion 598 -629 598 -629 0 feedthrough
rlabel pdiffusion 605 -629 605 -629 0 cellNo=161
rlabel pdiffusion 612 -629 612 -629 0 feedthrough
rlabel pdiffusion 619 -629 619 -629 0 feedthrough
rlabel pdiffusion 626 -629 626 -629 0 feedthrough
rlabel pdiffusion 633 -629 633 -629 0 feedthrough
rlabel pdiffusion 640 -629 640 -629 0 cellNo=672
rlabel pdiffusion 647 -629 647 -629 0 cellNo=56
rlabel pdiffusion 654 -629 654 -629 0 feedthrough
rlabel pdiffusion 661 -629 661 -629 0 feedthrough
rlabel pdiffusion 668 -629 668 -629 0 feedthrough
rlabel pdiffusion 675 -629 675 -629 0 feedthrough
rlabel pdiffusion 682 -629 682 -629 0 cellNo=72
rlabel pdiffusion 689 -629 689 -629 0 feedthrough
rlabel pdiffusion 696 -629 696 -629 0 cellNo=141
rlabel pdiffusion 703 -629 703 -629 0 feedthrough
rlabel pdiffusion 710 -629 710 -629 0 feedthrough
rlabel pdiffusion 717 -629 717 -629 0 feedthrough
rlabel pdiffusion 724 -629 724 -629 0 feedthrough
rlabel pdiffusion 731 -629 731 -629 0 cellNo=109
rlabel pdiffusion 738 -629 738 -629 0 feedthrough
rlabel pdiffusion 745 -629 745 -629 0 cellNo=350
rlabel pdiffusion 752 -629 752 -629 0 feedthrough
rlabel pdiffusion 759 -629 759 -629 0 cellNo=297
rlabel pdiffusion 766 -629 766 -629 0 feedthrough
rlabel pdiffusion 773 -629 773 -629 0 feedthrough
rlabel pdiffusion 780 -629 780 -629 0 feedthrough
rlabel pdiffusion 787 -629 787 -629 0 cellNo=107
rlabel pdiffusion 794 -629 794 -629 0 feedthrough
rlabel pdiffusion 801 -629 801 -629 0 cellNo=113
rlabel pdiffusion 808 -629 808 -629 0 feedthrough
rlabel pdiffusion 815 -629 815 -629 0 feedthrough
rlabel pdiffusion 822 -629 822 -629 0 feedthrough
rlabel pdiffusion 829 -629 829 -629 0 feedthrough
rlabel pdiffusion 836 -629 836 -629 0 feedthrough
rlabel pdiffusion 843 -629 843 -629 0 cellNo=712
rlabel pdiffusion 850 -629 850 -629 0 feedthrough
rlabel pdiffusion 857 -629 857 -629 0 feedthrough
rlabel pdiffusion 864 -629 864 -629 0 feedthrough
rlabel pdiffusion 871 -629 871 -629 0 cellNo=763
rlabel pdiffusion 878 -629 878 -629 0 feedthrough
rlabel pdiffusion 885 -629 885 -629 0 feedthrough
rlabel pdiffusion 892 -629 892 -629 0 feedthrough
rlabel pdiffusion 899 -629 899 -629 0 feedthrough
rlabel pdiffusion 906 -629 906 -629 0 feedthrough
rlabel pdiffusion 913 -629 913 -629 0 feedthrough
rlabel pdiffusion 920 -629 920 -629 0 feedthrough
rlabel pdiffusion 927 -629 927 -629 0 feedthrough
rlabel pdiffusion 934 -629 934 -629 0 feedthrough
rlabel pdiffusion 941 -629 941 -629 0 feedthrough
rlabel pdiffusion 948 -629 948 -629 0 feedthrough
rlabel pdiffusion 955 -629 955 -629 0 feedthrough
rlabel pdiffusion 962 -629 962 -629 0 feedthrough
rlabel pdiffusion 969 -629 969 -629 0 feedthrough
rlabel pdiffusion 976 -629 976 -629 0 feedthrough
rlabel pdiffusion 983 -629 983 -629 0 feedthrough
rlabel pdiffusion 990 -629 990 -629 0 feedthrough
rlabel pdiffusion 997 -629 997 -629 0 feedthrough
rlabel pdiffusion 1004 -629 1004 -629 0 feedthrough
rlabel pdiffusion 1011 -629 1011 -629 0 feedthrough
rlabel pdiffusion 1018 -629 1018 -629 0 cellNo=242
rlabel pdiffusion 1025 -629 1025 -629 0 feedthrough
rlabel pdiffusion 1032 -629 1032 -629 0 cellNo=895
rlabel pdiffusion 1039 -629 1039 -629 0 feedthrough
rlabel pdiffusion 1046 -629 1046 -629 0 feedthrough
rlabel pdiffusion 1053 -629 1053 -629 0 feedthrough
rlabel pdiffusion 1060 -629 1060 -629 0 feedthrough
rlabel pdiffusion 1067 -629 1067 -629 0 feedthrough
rlabel pdiffusion 1074 -629 1074 -629 0 feedthrough
rlabel pdiffusion 1081 -629 1081 -629 0 feedthrough
rlabel pdiffusion 1088 -629 1088 -629 0 feedthrough
rlabel pdiffusion 1095 -629 1095 -629 0 feedthrough
rlabel pdiffusion 1102 -629 1102 -629 0 feedthrough
rlabel pdiffusion 1109 -629 1109 -629 0 feedthrough
rlabel pdiffusion 1116 -629 1116 -629 0 feedthrough
rlabel pdiffusion 1123 -629 1123 -629 0 feedthrough
rlabel pdiffusion 1130 -629 1130 -629 0 feedthrough
rlabel pdiffusion 1137 -629 1137 -629 0 feedthrough
rlabel pdiffusion 1144 -629 1144 -629 0 feedthrough
rlabel pdiffusion 1151 -629 1151 -629 0 feedthrough
rlabel pdiffusion 1158 -629 1158 -629 0 feedthrough
rlabel pdiffusion 1165 -629 1165 -629 0 feedthrough
rlabel pdiffusion 1172 -629 1172 -629 0 feedthrough
rlabel pdiffusion 1179 -629 1179 -629 0 feedthrough
rlabel pdiffusion 1186 -629 1186 -629 0 feedthrough
rlabel pdiffusion 1193 -629 1193 -629 0 feedthrough
rlabel pdiffusion 1200 -629 1200 -629 0 feedthrough
rlabel pdiffusion 1207 -629 1207 -629 0 feedthrough
rlabel pdiffusion 1214 -629 1214 -629 0 feedthrough
rlabel pdiffusion 1221 -629 1221 -629 0 feedthrough
rlabel pdiffusion 1228 -629 1228 -629 0 feedthrough
rlabel pdiffusion 1235 -629 1235 -629 0 feedthrough
rlabel pdiffusion 1242 -629 1242 -629 0 feedthrough
rlabel pdiffusion 1249 -629 1249 -629 0 feedthrough
rlabel pdiffusion 1256 -629 1256 -629 0 feedthrough
rlabel pdiffusion 1263 -629 1263 -629 0 feedthrough
rlabel pdiffusion 1270 -629 1270 -629 0 feedthrough
rlabel pdiffusion 1277 -629 1277 -629 0 feedthrough
rlabel pdiffusion 1284 -629 1284 -629 0 feedthrough
rlabel pdiffusion 1291 -629 1291 -629 0 feedthrough
rlabel pdiffusion 1298 -629 1298 -629 0 feedthrough
rlabel pdiffusion 1305 -629 1305 -629 0 feedthrough
rlabel pdiffusion 1312 -629 1312 -629 0 feedthrough
rlabel pdiffusion 1319 -629 1319 -629 0 feedthrough
rlabel pdiffusion 1326 -629 1326 -629 0 feedthrough
rlabel pdiffusion 1333 -629 1333 -629 0 feedthrough
rlabel pdiffusion 1340 -629 1340 -629 0 feedthrough
rlabel pdiffusion 1347 -629 1347 -629 0 feedthrough
rlabel pdiffusion 1354 -629 1354 -629 0 feedthrough
rlabel pdiffusion 1361 -629 1361 -629 0 feedthrough
rlabel pdiffusion 1368 -629 1368 -629 0 feedthrough
rlabel pdiffusion 1375 -629 1375 -629 0 feedthrough
rlabel pdiffusion 1382 -629 1382 -629 0 feedthrough
rlabel pdiffusion 1389 -629 1389 -629 0 feedthrough
rlabel pdiffusion 1396 -629 1396 -629 0 feedthrough
rlabel pdiffusion 1403 -629 1403 -629 0 feedthrough
rlabel pdiffusion 1410 -629 1410 -629 0 feedthrough
rlabel pdiffusion 1417 -629 1417 -629 0 cellNo=994
rlabel pdiffusion 1424 -629 1424 -629 0 feedthrough
rlabel pdiffusion 1431 -629 1431 -629 0 feedthrough
rlabel pdiffusion 1438 -629 1438 -629 0 feedthrough
rlabel pdiffusion 1445 -629 1445 -629 0 feedthrough
rlabel pdiffusion 1452 -629 1452 -629 0 feedthrough
rlabel pdiffusion 1459 -629 1459 -629 0 feedthrough
rlabel pdiffusion 1466 -629 1466 -629 0 feedthrough
rlabel pdiffusion 1529 -629 1529 -629 0 feedthrough
rlabel pdiffusion 1550 -629 1550 -629 0 feedthrough
rlabel pdiffusion 1620 -629 1620 -629 0 feedthrough
rlabel pdiffusion 3 -762 3 -762 0 cellNo=1033
rlabel pdiffusion 10 -762 10 -762 0 cellNo=1172
rlabel pdiffusion 17 -762 17 -762 0 cellNo=1126
rlabel pdiffusion 24 -762 24 -762 0 cellNo=1071
rlabel pdiffusion 31 -762 31 -762 0 cellNo=1090
rlabel pdiffusion 38 -762 38 -762 0 cellNo=1106
rlabel pdiffusion 45 -762 45 -762 0 feedthrough
rlabel pdiffusion 52 -762 52 -762 0 feedthrough
rlabel pdiffusion 59 -762 59 -762 0 cellNo=632
rlabel pdiffusion 66 -762 66 -762 0 cellNo=321
rlabel pdiffusion 73 -762 73 -762 0 feedthrough
rlabel pdiffusion 80 -762 80 -762 0 feedthrough
rlabel pdiffusion 87 -762 87 -762 0 feedthrough
rlabel pdiffusion 94 -762 94 -762 0 feedthrough
rlabel pdiffusion 101 -762 101 -762 0 feedthrough
rlabel pdiffusion 108 -762 108 -762 0 feedthrough
rlabel pdiffusion 115 -762 115 -762 0 cellNo=11
rlabel pdiffusion 122 -762 122 -762 0 feedthrough
rlabel pdiffusion 129 -762 129 -762 0 feedthrough
rlabel pdiffusion 136 -762 136 -762 0 feedthrough
rlabel pdiffusion 143 -762 143 -762 0 feedthrough
rlabel pdiffusion 150 -762 150 -762 0 feedthrough
rlabel pdiffusion 157 -762 157 -762 0 cellNo=146
rlabel pdiffusion 164 -762 164 -762 0 feedthrough
rlabel pdiffusion 171 -762 171 -762 0 feedthrough
rlabel pdiffusion 178 -762 178 -762 0 feedthrough
rlabel pdiffusion 185 -762 185 -762 0 feedthrough
rlabel pdiffusion 192 -762 192 -762 0 feedthrough
rlabel pdiffusion 199 -762 199 -762 0 feedthrough
rlabel pdiffusion 206 -762 206 -762 0 cellNo=357
rlabel pdiffusion 213 -762 213 -762 0 feedthrough
rlabel pdiffusion 220 -762 220 -762 0 cellNo=564
rlabel pdiffusion 227 -762 227 -762 0 feedthrough
rlabel pdiffusion 234 -762 234 -762 0 feedthrough
rlabel pdiffusion 241 -762 241 -762 0 feedthrough
rlabel pdiffusion 248 -762 248 -762 0 feedthrough
rlabel pdiffusion 255 -762 255 -762 0 cellNo=34
rlabel pdiffusion 262 -762 262 -762 0 feedthrough
rlabel pdiffusion 269 -762 269 -762 0 feedthrough
rlabel pdiffusion 276 -762 276 -762 0 feedthrough
rlabel pdiffusion 283 -762 283 -762 0 feedthrough
rlabel pdiffusion 290 -762 290 -762 0 feedthrough
rlabel pdiffusion 297 -762 297 -762 0 feedthrough
rlabel pdiffusion 304 -762 304 -762 0 feedthrough
rlabel pdiffusion 311 -762 311 -762 0 feedthrough
rlabel pdiffusion 318 -762 318 -762 0 feedthrough
rlabel pdiffusion 325 -762 325 -762 0 feedthrough
rlabel pdiffusion 332 -762 332 -762 0 cellNo=401
rlabel pdiffusion 339 -762 339 -762 0 feedthrough
rlabel pdiffusion 346 -762 346 -762 0 feedthrough
rlabel pdiffusion 353 -762 353 -762 0 feedthrough
rlabel pdiffusion 360 -762 360 -762 0 feedthrough
rlabel pdiffusion 367 -762 367 -762 0 feedthrough
rlabel pdiffusion 374 -762 374 -762 0 feedthrough
rlabel pdiffusion 381 -762 381 -762 0 feedthrough
rlabel pdiffusion 388 -762 388 -762 0 feedthrough
rlabel pdiffusion 395 -762 395 -762 0 feedthrough
rlabel pdiffusion 402 -762 402 -762 0 feedthrough
rlabel pdiffusion 409 -762 409 -762 0 feedthrough
rlabel pdiffusion 416 -762 416 -762 0 feedthrough
rlabel pdiffusion 423 -762 423 -762 0 feedthrough
rlabel pdiffusion 430 -762 430 -762 0 cellNo=181
rlabel pdiffusion 437 -762 437 -762 0 feedthrough
rlabel pdiffusion 444 -762 444 -762 0 feedthrough
rlabel pdiffusion 451 -762 451 -762 0 feedthrough
rlabel pdiffusion 458 -762 458 -762 0 feedthrough
rlabel pdiffusion 465 -762 465 -762 0 cellNo=409
rlabel pdiffusion 472 -762 472 -762 0 feedthrough
rlabel pdiffusion 479 -762 479 -762 0 feedthrough
rlabel pdiffusion 486 -762 486 -762 0 feedthrough
rlabel pdiffusion 493 -762 493 -762 0 cellNo=513
rlabel pdiffusion 500 -762 500 -762 0 feedthrough
rlabel pdiffusion 507 -762 507 -762 0 feedthrough
rlabel pdiffusion 514 -762 514 -762 0 feedthrough
rlabel pdiffusion 521 -762 521 -762 0 cellNo=413
rlabel pdiffusion 528 -762 528 -762 0 cellNo=269
rlabel pdiffusion 535 -762 535 -762 0 feedthrough
rlabel pdiffusion 542 -762 542 -762 0 feedthrough
rlabel pdiffusion 549 -762 549 -762 0 feedthrough
rlabel pdiffusion 556 -762 556 -762 0 cellNo=874
rlabel pdiffusion 563 -762 563 -762 0 feedthrough
rlabel pdiffusion 570 -762 570 -762 0 cellNo=143
rlabel pdiffusion 577 -762 577 -762 0 feedthrough
rlabel pdiffusion 584 -762 584 -762 0 feedthrough
rlabel pdiffusion 591 -762 591 -762 0 feedthrough
rlabel pdiffusion 598 -762 598 -762 0 feedthrough
rlabel pdiffusion 605 -762 605 -762 0 cellNo=372
rlabel pdiffusion 612 -762 612 -762 0 feedthrough
rlabel pdiffusion 619 -762 619 -762 0 feedthrough
rlabel pdiffusion 626 -762 626 -762 0 feedthrough
rlabel pdiffusion 633 -762 633 -762 0 cellNo=27
rlabel pdiffusion 640 -762 640 -762 0 feedthrough
rlabel pdiffusion 647 -762 647 -762 0 cellNo=786
rlabel pdiffusion 654 -762 654 -762 0 feedthrough
rlabel pdiffusion 661 -762 661 -762 0 feedthrough
rlabel pdiffusion 668 -762 668 -762 0 feedthrough
rlabel pdiffusion 675 -762 675 -762 0 cellNo=329
rlabel pdiffusion 682 -762 682 -762 0 feedthrough
rlabel pdiffusion 689 -762 689 -762 0 cellNo=280
rlabel pdiffusion 696 -762 696 -762 0 feedthrough
rlabel pdiffusion 703 -762 703 -762 0 feedthrough
rlabel pdiffusion 710 -762 710 -762 0 feedthrough
rlabel pdiffusion 717 -762 717 -762 0 cellNo=265
rlabel pdiffusion 724 -762 724 -762 0 feedthrough
rlabel pdiffusion 731 -762 731 -762 0 cellNo=689
rlabel pdiffusion 738 -762 738 -762 0 feedthrough
rlabel pdiffusion 745 -762 745 -762 0 feedthrough
rlabel pdiffusion 752 -762 752 -762 0 feedthrough
rlabel pdiffusion 759 -762 759 -762 0 feedthrough
rlabel pdiffusion 766 -762 766 -762 0 feedthrough
rlabel pdiffusion 773 -762 773 -762 0 feedthrough
rlabel pdiffusion 780 -762 780 -762 0 feedthrough
rlabel pdiffusion 787 -762 787 -762 0 feedthrough
rlabel pdiffusion 794 -762 794 -762 0 cellNo=492
rlabel pdiffusion 801 -762 801 -762 0 cellNo=947
rlabel pdiffusion 808 -762 808 -762 0 feedthrough
rlabel pdiffusion 815 -762 815 -762 0 feedthrough
rlabel pdiffusion 822 -762 822 -762 0 feedthrough
rlabel pdiffusion 829 -762 829 -762 0 cellNo=51
rlabel pdiffusion 836 -762 836 -762 0 cellNo=718
rlabel pdiffusion 843 -762 843 -762 0 feedthrough
rlabel pdiffusion 850 -762 850 -762 0 feedthrough
rlabel pdiffusion 857 -762 857 -762 0 feedthrough
rlabel pdiffusion 864 -762 864 -762 0 feedthrough
rlabel pdiffusion 871 -762 871 -762 0 cellNo=599
rlabel pdiffusion 878 -762 878 -762 0 feedthrough
rlabel pdiffusion 885 -762 885 -762 0 feedthrough
rlabel pdiffusion 892 -762 892 -762 0 feedthrough
rlabel pdiffusion 899 -762 899 -762 0 feedthrough
rlabel pdiffusion 906 -762 906 -762 0 cellNo=852
rlabel pdiffusion 913 -762 913 -762 0 feedthrough
rlabel pdiffusion 920 -762 920 -762 0 feedthrough
rlabel pdiffusion 927 -762 927 -762 0 cellNo=257
rlabel pdiffusion 934 -762 934 -762 0 feedthrough
rlabel pdiffusion 941 -762 941 -762 0 feedthrough
rlabel pdiffusion 948 -762 948 -762 0 feedthrough
rlabel pdiffusion 955 -762 955 -762 0 feedthrough
rlabel pdiffusion 962 -762 962 -762 0 feedthrough
rlabel pdiffusion 969 -762 969 -762 0 feedthrough
rlabel pdiffusion 976 -762 976 -762 0 feedthrough
rlabel pdiffusion 983 -762 983 -762 0 feedthrough
rlabel pdiffusion 990 -762 990 -762 0 feedthrough
rlabel pdiffusion 997 -762 997 -762 0 feedthrough
rlabel pdiffusion 1004 -762 1004 -762 0 feedthrough
rlabel pdiffusion 1011 -762 1011 -762 0 feedthrough
rlabel pdiffusion 1018 -762 1018 -762 0 feedthrough
rlabel pdiffusion 1025 -762 1025 -762 0 cellNo=965
rlabel pdiffusion 1032 -762 1032 -762 0 feedthrough
rlabel pdiffusion 1039 -762 1039 -762 0 feedthrough
rlabel pdiffusion 1046 -762 1046 -762 0 feedthrough
rlabel pdiffusion 1053 -762 1053 -762 0 feedthrough
rlabel pdiffusion 1060 -762 1060 -762 0 feedthrough
rlabel pdiffusion 1067 -762 1067 -762 0 feedthrough
rlabel pdiffusion 1074 -762 1074 -762 0 feedthrough
rlabel pdiffusion 1081 -762 1081 -762 0 feedthrough
rlabel pdiffusion 1088 -762 1088 -762 0 feedthrough
rlabel pdiffusion 1095 -762 1095 -762 0 feedthrough
rlabel pdiffusion 1102 -762 1102 -762 0 feedthrough
rlabel pdiffusion 1109 -762 1109 -762 0 feedthrough
rlabel pdiffusion 1116 -762 1116 -762 0 feedthrough
rlabel pdiffusion 1123 -762 1123 -762 0 feedthrough
rlabel pdiffusion 1130 -762 1130 -762 0 feedthrough
rlabel pdiffusion 1137 -762 1137 -762 0 feedthrough
rlabel pdiffusion 1144 -762 1144 -762 0 feedthrough
rlabel pdiffusion 1151 -762 1151 -762 0 feedthrough
rlabel pdiffusion 1158 -762 1158 -762 0 feedthrough
rlabel pdiffusion 1165 -762 1165 -762 0 feedthrough
rlabel pdiffusion 1172 -762 1172 -762 0 feedthrough
rlabel pdiffusion 1179 -762 1179 -762 0 feedthrough
rlabel pdiffusion 1186 -762 1186 -762 0 feedthrough
rlabel pdiffusion 1193 -762 1193 -762 0 feedthrough
rlabel pdiffusion 1200 -762 1200 -762 0 feedthrough
rlabel pdiffusion 1207 -762 1207 -762 0 feedthrough
rlabel pdiffusion 1214 -762 1214 -762 0 feedthrough
rlabel pdiffusion 1221 -762 1221 -762 0 feedthrough
rlabel pdiffusion 1228 -762 1228 -762 0 feedthrough
rlabel pdiffusion 1235 -762 1235 -762 0 feedthrough
rlabel pdiffusion 1242 -762 1242 -762 0 feedthrough
rlabel pdiffusion 1249 -762 1249 -762 0 feedthrough
rlabel pdiffusion 1256 -762 1256 -762 0 feedthrough
rlabel pdiffusion 1263 -762 1263 -762 0 feedthrough
rlabel pdiffusion 1270 -762 1270 -762 0 feedthrough
rlabel pdiffusion 1277 -762 1277 -762 0 feedthrough
rlabel pdiffusion 1284 -762 1284 -762 0 feedthrough
rlabel pdiffusion 1291 -762 1291 -762 0 feedthrough
rlabel pdiffusion 1298 -762 1298 -762 0 feedthrough
rlabel pdiffusion 1305 -762 1305 -762 0 feedthrough
rlabel pdiffusion 1312 -762 1312 -762 0 feedthrough
rlabel pdiffusion 1319 -762 1319 -762 0 feedthrough
rlabel pdiffusion 1326 -762 1326 -762 0 feedthrough
rlabel pdiffusion 1333 -762 1333 -762 0 feedthrough
rlabel pdiffusion 1340 -762 1340 -762 0 feedthrough
rlabel pdiffusion 1347 -762 1347 -762 0 feedthrough
rlabel pdiffusion 1354 -762 1354 -762 0 feedthrough
rlabel pdiffusion 1361 -762 1361 -762 0 feedthrough
rlabel pdiffusion 1368 -762 1368 -762 0 feedthrough
rlabel pdiffusion 1375 -762 1375 -762 0 feedthrough
rlabel pdiffusion 1382 -762 1382 -762 0 feedthrough
rlabel pdiffusion 1389 -762 1389 -762 0 feedthrough
rlabel pdiffusion 1396 -762 1396 -762 0 feedthrough
rlabel pdiffusion 1403 -762 1403 -762 0 feedthrough
rlabel pdiffusion 1410 -762 1410 -762 0 feedthrough
rlabel pdiffusion 1417 -762 1417 -762 0 feedthrough
rlabel pdiffusion 1424 -762 1424 -762 0 feedthrough
rlabel pdiffusion 1431 -762 1431 -762 0 feedthrough
rlabel pdiffusion 1438 -762 1438 -762 0 feedthrough
rlabel pdiffusion 1445 -762 1445 -762 0 feedthrough
rlabel pdiffusion 1452 -762 1452 -762 0 feedthrough
rlabel pdiffusion 1459 -762 1459 -762 0 feedthrough
rlabel pdiffusion 1466 -762 1466 -762 0 feedthrough
rlabel pdiffusion 1473 -762 1473 -762 0 feedthrough
rlabel pdiffusion 1480 -762 1480 -762 0 feedthrough
rlabel pdiffusion 1487 -762 1487 -762 0 feedthrough
rlabel pdiffusion 1529 -762 1529 -762 0 feedthrough
rlabel pdiffusion 1550 -762 1550 -762 0 feedthrough
rlabel pdiffusion 1557 -762 1557 -762 0 feedthrough
rlabel pdiffusion 1697 -762 1697 -762 0 feedthrough
rlabel pdiffusion 3 -875 3 -875 0 cellNo=1043
rlabel pdiffusion 10 -875 10 -875 0 cellNo=1058
rlabel pdiffusion 17 -875 17 -875 0 cellNo=1149
rlabel pdiffusion 24 -875 24 -875 0 cellNo=1089
rlabel pdiffusion 31 -875 31 -875 0 cellNo=1105
rlabel pdiffusion 38 -875 38 -875 0 feedthrough
rlabel pdiffusion 45 -875 45 -875 0 feedthrough
rlabel pdiffusion 52 -875 52 -875 0 feedthrough
rlabel pdiffusion 59 -875 59 -875 0 feedthrough
rlabel pdiffusion 66 -875 66 -875 0 feedthrough
rlabel pdiffusion 73 -875 73 -875 0 feedthrough
rlabel pdiffusion 80 -875 80 -875 0 feedthrough
rlabel pdiffusion 87 -875 87 -875 0 feedthrough
rlabel pdiffusion 94 -875 94 -875 0 feedthrough
rlabel pdiffusion 101 -875 101 -875 0 feedthrough
rlabel pdiffusion 108 -875 108 -875 0 cellNo=157
rlabel pdiffusion 115 -875 115 -875 0 feedthrough
rlabel pdiffusion 122 -875 122 -875 0 cellNo=767
rlabel pdiffusion 129 -875 129 -875 0 feedthrough
rlabel pdiffusion 136 -875 136 -875 0 feedthrough
rlabel pdiffusion 143 -875 143 -875 0 feedthrough
rlabel pdiffusion 150 -875 150 -875 0 cellNo=803
rlabel pdiffusion 157 -875 157 -875 0 feedthrough
rlabel pdiffusion 164 -875 164 -875 0 cellNo=349
rlabel pdiffusion 171 -875 171 -875 0 feedthrough
rlabel pdiffusion 178 -875 178 -875 0 feedthrough
rlabel pdiffusion 185 -875 185 -875 0 cellNo=197
rlabel pdiffusion 192 -875 192 -875 0 feedthrough
rlabel pdiffusion 199 -875 199 -875 0 feedthrough
rlabel pdiffusion 206 -875 206 -875 0 cellNo=384
rlabel pdiffusion 213 -875 213 -875 0 feedthrough
rlabel pdiffusion 220 -875 220 -875 0 cellNo=339
rlabel pdiffusion 227 -875 227 -875 0 feedthrough
rlabel pdiffusion 234 -875 234 -875 0 feedthrough
rlabel pdiffusion 241 -875 241 -875 0 feedthrough
rlabel pdiffusion 248 -875 248 -875 0 feedthrough
rlabel pdiffusion 255 -875 255 -875 0 cellNo=48
rlabel pdiffusion 262 -875 262 -875 0 feedthrough
rlabel pdiffusion 269 -875 269 -875 0 feedthrough
rlabel pdiffusion 276 -875 276 -875 0 feedthrough
rlabel pdiffusion 283 -875 283 -875 0 feedthrough
rlabel pdiffusion 290 -875 290 -875 0 feedthrough
rlabel pdiffusion 297 -875 297 -875 0 feedthrough
rlabel pdiffusion 304 -875 304 -875 0 feedthrough
rlabel pdiffusion 311 -875 311 -875 0 feedthrough
rlabel pdiffusion 318 -875 318 -875 0 feedthrough
rlabel pdiffusion 325 -875 325 -875 0 feedthrough
rlabel pdiffusion 332 -875 332 -875 0 feedthrough
rlabel pdiffusion 339 -875 339 -875 0 feedthrough
rlabel pdiffusion 346 -875 346 -875 0 feedthrough
rlabel pdiffusion 353 -875 353 -875 0 feedthrough
rlabel pdiffusion 360 -875 360 -875 0 feedthrough
rlabel pdiffusion 367 -875 367 -875 0 feedthrough
rlabel pdiffusion 374 -875 374 -875 0 feedthrough
rlabel pdiffusion 381 -875 381 -875 0 feedthrough
rlabel pdiffusion 388 -875 388 -875 0 feedthrough
rlabel pdiffusion 395 -875 395 -875 0 feedthrough
rlabel pdiffusion 402 -875 402 -875 0 feedthrough
rlabel pdiffusion 409 -875 409 -875 0 cellNo=341
rlabel pdiffusion 416 -875 416 -875 0 feedthrough
rlabel pdiffusion 423 -875 423 -875 0 feedthrough
rlabel pdiffusion 430 -875 430 -875 0 feedthrough
rlabel pdiffusion 437 -875 437 -875 0 feedthrough
rlabel pdiffusion 444 -875 444 -875 0 feedthrough
rlabel pdiffusion 451 -875 451 -875 0 feedthrough
rlabel pdiffusion 458 -875 458 -875 0 feedthrough
rlabel pdiffusion 465 -875 465 -875 0 feedthrough
rlabel pdiffusion 472 -875 472 -875 0 feedthrough
rlabel pdiffusion 479 -875 479 -875 0 feedthrough
rlabel pdiffusion 486 -875 486 -875 0 feedthrough
rlabel pdiffusion 493 -875 493 -875 0 feedthrough
rlabel pdiffusion 500 -875 500 -875 0 cellNo=307
rlabel pdiffusion 507 -875 507 -875 0 cellNo=471
rlabel pdiffusion 514 -875 514 -875 0 feedthrough
rlabel pdiffusion 521 -875 521 -875 0 cellNo=860
rlabel pdiffusion 528 -875 528 -875 0 cellNo=331
rlabel pdiffusion 535 -875 535 -875 0 cellNo=902
rlabel pdiffusion 542 -875 542 -875 0 feedthrough
rlabel pdiffusion 549 -875 549 -875 0 cellNo=191
rlabel pdiffusion 556 -875 556 -875 0 feedthrough
rlabel pdiffusion 563 -875 563 -875 0 feedthrough
rlabel pdiffusion 570 -875 570 -875 0 feedthrough
rlabel pdiffusion 577 -875 577 -875 0 feedthrough
rlabel pdiffusion 584 -875 584 -875 0 feedthrough
rlabel pdiffusion 591 -875 591 -875 0 feedthrough
rlabel pdiffusion 598 -875 598 -875 0 feedthrough
rlabel pdiffusion 605 -875 605 -875 0 feedthrough
rlabel pdiffusion 612 -875 612 -875 0 feedthrough
rlabel pdiffusion 619 -875 619 -875 0 feedthrough
rlabel pdiffusion 626 -875 626 -875 0 cellNo=499
rlabel pdiffusion 633 -875 633 -875 0 feedthrough
rlabel pdiffusion 640 -875 640 -875 0 feedthrough
rlabel pdiffusion 647 -875 647 -875 0 cellNo=160
rlabel pdiffusion 654 -875 654 -875 0 feedthrough
rlabel pdiffusion 661 -875 661 -875 0 feedthrough
rlabel pdiffusion 668 -875 668 -875 0 cellNo=33
rlabel pdiffusion 675 -875 675 -875 0 cellNo=235
rlabel pdiffusion 682 -875 682 -875 0 cellNo=586
rlabel pdiffusion 689 -875 689 -875 0 feedthrough
rlabel pdiffusion 696 -875 696 -875 0 feedthrough
rlabel pdiffusion 703 -875 703 -875 0 feedthrough
rlabel pdiffusion 710 -875 710 -875 0 feedthrough
rlabel pdiffusion 717 -875 717 -875 0 feedthrough
rlabel pdiffusion 724 -875 724 -875 0 feedthrough
rlabel pdiffusion 731 -875 731 -875 0 feedthrough
rlabel pdiffusion 738 -875 738 -875 0 feedthrough
rlabel pdiffusion 745 -875 745 -875 0 feedthrough
rlabel pdiffusion 752 -875 752 -875 0 feedthrough
rlabel pdiffusion 759 -875 759 -875 0 feedthrough
rlabel pdiffusion 766 -875 766 -875 0 feedthrough
rlabel pdiffusion 773 -875 773 -875 0 feedthrough
rlabel pdiffusion 780 -875 780 -875 0 cellNo=378
rlabel pdiffusion 787 -875 787 -875 0 feedthrough
rlabel pdiffusion 794 -875 794 -875 0 feedthrough
rlabel pdiffusion 801 -875 801 -875 0 feedthrough
rlabel pdiffusion 808 -875 808 -875 0 feedthrough
rlabel pdiffusion 815 -875 815 -875 0 cellNo=468
rlabel pdiffusion 822 -875 822 -875 0 feedthrough
rlabel pdiffusion 829 -875 829 -875 0 cellNo=845
rlabel pdiffusion 836 -875 836 -875 0 cellNo=990
rlabel pdiffusion 843 -875 843 -875 0 feedthrough
rlabel pdiffusion 850 -875 850 -875 0 feedthrough
rlabel pdiffusion 857 -875 857 -875 0 feedthrough
rlabel pdiffusion 864 -875 864 -875 0 feedthrough
rlabel pdiffusion 871 -875 871 -875 0 cellNo=28
rlabel pdiffusion 878 -875 878 -875 0 cellNo=663
rlabel pdiffusion 885 -875 885 -875 0 feedthrough
rlabel pdiffusion 892 -875 892 -875 0 feedthrough
rlabel pdiffusion 899 -875 899 -875 0 feedthrough
rlabel pdiffusion 906 -875 906 -875 0 feedthrough
rlabel pdiffusion 913 -875 913 -875 0 feedthrough
rlabel pdiffusion 920 -875 920 -875 0 cellNo=463
rlabel pdiffusion 927 -875 927 -875 0 feedthrough
rlabel pdiffusion 934 -875 934 -875 0 feedthrough
rlabel pdiffusion 941 -875 941 -875 0 feedthrough
rlabel pdiffusion 948 -875 948 -875 0 feedthrough
rlabel pdiffusion 955 -875 955 -875 0 feedthrough
rlabel pdiffusion 962 -875 962 -875 0 cellNo=675
rlabel pdiffusion 969 -875 969 -875 0 feedthrough
rlabel pdiffusion 976 -875 976 -875 0 feedthrough
rlabel pdiffusion 983 -875 983 -875 0 feedthrough
rlabel pdiffusion 990 -875 990 -875 0 feedthrough
rlabel pdiffusion 997 -875 997 -875 0 feedthrough
rlabel pdiffusion 1004 -875 1004 -875 0 feedthrough
rlabel pdiffusion 1011 -875 1011 -875 0 feedthrough
rlabel pdiffusion 1018 -875 1018 -875 0 feedthrough
rlabel pdiffusion 1025 -875 1025 -875 0 feedthrough
rlabel pdiffusion 1032 -875 1032 -875 0 feedthrough
rlabel pdiffusion 1039 -875 1039 -875 0 feedthrough
rlabel pdiffusion 1046 -875 1046 -875 0 feedthrough
rlabel pdiffusion 1053 -875 1053 -875 0 feedthrough
rlabel pdiffusion 1060 -875 1060 -875 0 feedthrough
rlabel pdiffusion 1067 -875 1067 -875 0 cellNo=967
rlabel pdiffusion 1074 -875 1074 -875 0 feedthrough
rlabel pdiffusion 1081 -875 1081 -875 0 feedthrough
rlabel pdiffusion 1088 -875 1088 -875 0 feedthrough
rlabel pdiffusion 1095 -875 1095 -875 0 feedthrough
rlabel pdiffusion 1102 -875 1102 -875 0 feedthrough
rlabel pdiffusion 1109 -875 1109 -875 0 feedthrough
rlabel pdiffusion 1116 -875 1116 -875 0 feedthrough
rlabel pdiffusion 1123 -875 1123 -875 0 feedthrough
rlabel pdiffusion 1130 -875 1130 -875 0 feedthrough
rlabel pdiffusion 1137 -875 1137 -875 0 feedthrough
rlabel pdiffusion 1144 -875 1144 -875 0 feedthrough
rlabel pdiffusion 1151 -875 1151 -875 0 feedthrough
rlabel pdiffusion 1158 -875 1158 -875 0 feedthrough
rlabel pdiffusion 1165 -875 1165 -875 0 feedthrough
rlabel pdiffusion 1172 -875 1172 -875 0 feedthrough
rlabel pdiffusion 1179 -875 1179 -875 0 feedthrough
rlabel pdiffusion 1186 -875 1186 -875 0 feedthrough
rlabel pdiffusion 1193 -875 1193 -875 0 feedthrough
rlabel pdiffusion 1200 -875 1200 -875 0 feedthrough
rlabel pdiffusion 1207 -875 1207 -875 0 feedthrough
rlabel pdiffusion 1214 -875 1214 -875 0 feedthrough
rlabel pdiffusion 1221 -875 1221 -875 0 feedthrough
rlabel pdiffusion 1228 -875 1228 -875 0 feedthrough
rlabel pdiffusion 1235 -875 1235 -875 0 feedthrough
rlabel pdiffusion 1242 -875 1242 -875 0 feedthrough
rlabel pdiffusion 1249 -875 1249 -875 0 feedthrough
rlabel pdiffusion 1256 -875 1256 -875 0 feedthrough
rlabel pdiffusion 1263 -875 1263 -875 0 feedthrough
rlabel pdiffusion 1270 -875 1270 -875 0 feedthrough
rlabel pdiffusion 1277 -875 1277 -875 0 feedthrough
rlabel pdiffusion 1284 -875 1284 -875 0 feedthrough
rlabel pdiffusion 1291 -875 1291 -875 0 feedthrough
rlabel pdiffusion 1298 -875 1298 -875 0 feedthrough
rlabel pdiffusion 1305 -875 1305 -875 0 feedthrough
rlabel pdiffusion 1312 -875 1312 -875 0 feedthrough
rlabel pdiffusion 1319 -875 1319 -875 0 feedthrough
rlabel pdiffusion 1326 -875 1326 -875 0 feedthrough
rlabel pdiffusion 1333 -875 1333 -875 0 feedthrough
rlabel pdiffusion 1340 -875 1340 -875 0 feedthrough
rlabel pdiffusion 1347 -875 1347 -875 0 feedthrough
rlabel pdiffusion 1354 -875 1354 -875 0 feedthrough
rlabel pdiffusion 1361 -875 1361 -875 0 feedthrough
rlabel pdiffusion 1368 -875 1368 -875 0 feedthrough
rlabel pdiffusion 1375 -875 1375 -875 0 feedthrough
rlabel pdiffusion 1382 -875 1382 -875 0 feedthrough
rlabel pdiffusion 1389 -875 1389 -875 0 feedthrough
rlabel pdiffusion 1396 -875 1396 -875 0 feedthrough
rlabel pdiffusion 1403 -875 1403 -875 0 feedthrough
rlabel pdiffusion 1410 -875 1410 -875 0 feedthrough
rlabel pdiffusion 1417 -875 1417 -875 0 feedthrough
rlabel pdiffusion 1424 -875 1424 -875 0 feedthrough
rlabel pdiffusion 1431 -875 1431 -875 0 feedthrough
rlabel pdiffusion 1438 -875 1438 -875 0 feedthrough
rlabel pdiffusion 1445 -875 1445 -875 0 feedthrough
rlabel pdiffusion 1452 -875 1452 -875 0 feedthrough
rlabel pdiffusion 1459 -875 1459 -875 0 feedthrough
rlabel pdiffusion 1466 -875 1466 -875 0 feedthrough
rlabel pdiffusion 1473 -875 1473 -875 0 feedthrough
rlabel pdiffusion 1480 -875 1480 -875 0 feedthrough
rlabel pdiffusion 1487 -875 1487 -875 0 feedthrough
rlabel pdiffusion 1494 -875 1494 -875 0 feedthrough
rlabel pdiffusion 1501 -875 1501 -875 0 feedthrough
rlabel pdiffusion 1508 -875 1508 -875 0 feedthrough
rlabel pdiffusion 1515 -875 1515 -875 0 feedthrough
rlabel pdiffusion 1522 -875 1522 -875 0 feedthrough
rlabel pdiffusion 1529 -875 1529 -875 0 feedthrough
rlabel pdiffusion 1536 -875 1536 -875 0 feedthrough
rlabel pdiffusion 1543 -875 1543 -875 0 feedthrough
rlabel pdiffusion 1550 -875 1550 -875 0 feedthrough
rlabel pdiffusion 1557 -875 1557 -875 0 cellNo=647
rlabel pdiffusion 1564 -875 1564 -875 0 cellNo=164
rlabel pdiffusion 1571 -875 1571 -875 0 feedthrough
rlabel pdiffusion 1578 -875 1578 -875 0 feedthrough
rlabel pdiffusion 1585 -875 1585 -875 0 feedthrough
rlabel pdiffusion 1725 -875 1725 -875 0 feedthrough
rlabel pdiffusion 3 -1002 3 -1002 0 cellNo=1057
rlabel pdiffusion 10 -1002 10 -1002 0 cellNo=1070
rlabel pdiffusion 17 -1002 17 -1002 0 cellNo=1088
rlabel pdiffusion 24 -1002 24 -1002 0 cellNo=1104
rlabel pdiffusion 31 -1002 31 -1002 0 feedthrough
rlabel pdiffusion 38 -1002 38 -1002 0 feedthrough
rlabel pdiffusion 45 -1002 45 -1002 0 feedthrough
rlabel pdiffusion 52 -1002 52 -1002 0 feedthrough
rlabel pdiffusion 59 -1002 59 -1002 0 feedthrough
rlabel pdiffusion 66 -1002 66 -1002 0 feedthrough
rlabel pdiffusion 73 -1002 73 -1002 0 feedthrough
rlabel pdiffusion 80 -1002 80 -1002 0 cellNo=410
rlabel pdiffusion 87 -1002 87 -1002 0 feedthrough
rlabel pdiffusion 94 -1002 94 -1002 0 feedthrough
rlabel pdiffusion 101 -1002 101 -1002 0 feedthrough
rlabel pdiffusion 108 -1002 108 -1002 0 feedthrough
rlabel pdiffusion 115 -1002 115 -1002 0 feedthrough
rlabel pdiffusion 122 -1002 122 -1002 0 feedthrough
rlabel pdiffusion 129 -1002 129 -1002 0 cellNo=21
rlabel pdiffusion 136 -1002 136 -1002 0 cellNo=958
rlabel pdiffusion 143 -1002 143 -1002 0 feedthrough
rlabel pdiffusion 150 -1002 150 -1002 0 cellNo=271
rlabel pdiffusion 157 -1002 157 -1002 0 feedthrough
rlabel pdiffusion 164 -1002 164 -1002 0 feedthrough
rlabel pdiffusion 171 -1002 171 -1002 0 feedthrough
rlabel pdiffusion 178 -1002 178 -1002 0 feedthrough
rlabel pdiffusion 185 -1002 185 -1002 0 feedthrough
rlabel pdiffusion 192 -1002 192 -1002 0 feedthrough
rlabel pdiffusion 199 -1002 199 -1002 0 feedthrough
rlabel pdiffusion 206 -1002 206 -1002 0 feedthrough
rlabel pdiffusion 213 -1002 213 -1002 0 feedthrough
rlabel pdiffusion 220 -1002 220 -1002 0 feedthrough
rlabel pdiffusion 227 -1002 227 -1002 0 feedthrough
rlabel pdiffusion 234 -1002 234 -1002 0 feedthrough
rlabel pdiffusion 241 -1002 241 -1002 0 feedthrough
rlabel pdiffusion 248 -1002 248 -1002 0 cellNo=274
rlabel pdiffusion 255 -1002 255 -1002 0 feedthrough
rlabel pdiffusion 262 -1002 262 -1002 0 feedthrough
rlabel pdiffusion 269 -1002 269 -1002 0 feedthrough
rlabel pdiffusion 276 -1002 276 -1002 0 feedthrough
rlabel pdiffusion 283 -1002 283 -1002 0 feedthrough
rlabel pdiffusion 290 -1002 290 -1002 0 feedthrough
rlabel pdiffusion 297 -1002 297 -1002 0 feedthrough
rlabel pdiffusion 304 -1002 304 -1002 0 feedthrough
rlabel pdiffusion 311 -1002 311 -1002 0 feedthrough
rlabel pdiffusion 318 -1002 318 -1002 0 feedthrough
rlabel pdiffusion 325 -1002 325 -1002 0 feedthrough
rlabel pdiffusion 332 -1002 332 -1002 0 feedthrough
rlabel pdiffusion 339 -1002 339 -1002 0 feedthrough
rlabel pdiffusion 346 -1002 346 -1002 0 feedthrough
rlabel pdiffusion 353 -1002 353 -1002 0 feedthrough
rlabel pdiffusion 360 -1002 360 -1002 0 feedthrough
rlabel pdiffusion 367 -1002 367 -1002 0 feedthrough
rlabel pdiffusion 374 -1002 374 -1002 0 feedthrough
rlabel pdiffusion 381 -1002 381 -1002 0 feedthrough
rlabel pdiffusion 388 -1002 388 -1002 0 feedthrough
rlabel pdiffusion 395 -1002 395 -1002 0 feedthrough
rlabel pdiffusion 402 -1002 402 -1002 0 feedthrough
rlabel pdiffusion 409 -1002 409 -1002 0 feedthrough
rlabel pdiffusion 416 -1002 416 -1002 0 feedthrough
rlabel pdiffusion 423 -1002 423 -1002 0 cellNo=188
rlabel pdiffusion 430 -1002 430 -1002 0 feedthrough
rlabel pdiffusion 437 -1002 437 -1002 0 feedthrough
rlabel pdiffusion 444 -1002 444 -1002 0 cellNo=697
rlabel pdiffusion 451 -1002 451 -1002 0 feedthrough
rlabel pdiffusion 458 -1002 458 -1002 0 feedthrough
rlabel pdiffusion 465 -1002 465 -1002 0 feedthrough
rlabel pdiffusion 472 -1002 472 -1002 0 feedthrough
rlabel pdiffusion 479 -1002 479 -1002 0 feedthrough
rlabel pdiffusion 486 -1002 486 -1002 0 feedthrough
rlabel pdiffusion 493 -1002 493 -1002 0 feedthrough
rlabel pdiffusion 500 -1002 500 -1002 0 cellNo=980
rlabel pdiffusion 507 -1002 507 -1002 0 cellNo=977
rlabel pdiffusion 514 -1002 514 -1002 0 feedthrough
rlabel pdiffusion 521 -1002 521 -1002 0 feedthrough
rlabel pdiffusion 528 -1002 528 -1002 0 feedthrough
rlabel pdiffusion 535 -1002 535 -1002 0 feedthrough
rlabel pdiffusion 542 -1002 542 -1002 0 feedthrough
rlabel pdiffusion 549 -1002 549 -1002 0 feedthrough
rlabel pdiffusion 556 -1002 556 -1002 0 feedthrough
rlabel pdiffusion 563 -1002 563 -1002 0 feedthrough
rlabel pdiffusion 570 -1002 570 -1002 0 feedthrough
rlabel pdiffusion 577 -1002 577 -1002 0 feedthrough
rlabel pdiffusion 584 -1002 584 -1002 0 cellNo=692
rlabel pdiffusion 591 -1002 591 -1002 0 feedthrough
rlabel pdiffusion 598 -1002 598 -1002 0 feedthrough
rlabel pdiffusion 605 -1002 605 -1002 0 feedthrough
rlabel pdiffusion 612 -1002 612 -1002 0 feedthrough
rlabel pdiffusion 619 -1002 619 -1002 0 cellNo=728
rlabel pdiffusion 626 -1002 626 -1002 0 feedthrough
rlabel pdiffusion 633 -1002 633 -1002 0 feedthrough
rlabel pdiffusion 640 -1002 640 -1002 0 cellNo=600
rlabel pdiffusion 647 -1002 647 -1002 0 cellNo=54
rlabel pdiffusion 654 -1002 654 -1002 0 cellNo=110
rlabel pdiffusion 661 -1002 661 -1002 0 feedthrough
rlabel pdiffusion 668 -1002 668 -1002 0 feedthrough
rlabel pdiffusion 675 -1002 675 -1002 0 feedthrough
rlabel pdiffusion 682 -1002 682 -1002 0 cellNo=646
rlabel pdiffusion 689 -1002 689 -1002 0 cellNo=645
rlabel pdiffusion 696 -1002 696 -1002 0 cellNo=434
rlabel pdiffusion 703 -1002 703 -1002 0 feedthrough
rlabel pdiffusion 710 -1002 710 -1002 0 feedthrough
rlabel pdiffusion 717 -1002 717 -1002 0 feedthrough
rlabel pdiffusion 724 -1002 724 -1002 0 feedthrough
rlabel pdiffusion 731 -1002 731 -1002 0 cellNo=416
rlabel pdiffusion 738 -1002 738 -1002 0 feedthrough
rlabel pdiffusion 745 -1002 745 -1002 0 feedthrough
rlabel pdiffusion 752 -1002 752 -1002 0 feedthrough
rlabel pdiffusion 759 -1002 759 -1002 0 feedthrough
rlabel pdiffusion 766 -1002 766 -1002 0 cellNo=706
rlabel pdiffusion 773 -1002 773 -1002 0 cellNo=452
rlabel pdiffusion 780 -1002 780 -1002 0 feedthrough
rlabel pdiffusion 787 -1002 787 -1002 0 feedthrough
rlabel pdiffusion 794 -1002 794 -1002 0 feedthrough
rlabel pdiffusion 801 -1002 801 -1002 0 feedthrough
rlabel pdiffusion 808 -1002 808 -1002 0 feedthrough
rlabel pdiffusion 815 -1002 815 -1002 0 feedthrough
rlabel pdiffusion 822 -1002 822 -1002 0 feedthrough
rlabel pdiffusion 829 -1002 829 -1002 0 feedthrough
rlabel pdiffusion 836 -1002 836 -1002 0 feedthrough
rlabel pdiffusion 843 -1002 843 -1002 0 cellNo=245
rlabel pdiffusion 850 -1002 850 -1002 0 feedthrough
rlabel pdiffusion 857 -1002 857 -1002 0 feedthrough
rlabel pdiffusion 864 -1002 864 -1002 0 feedthrough
rlabel pdiffusion 871 -1002 871 -1002 0 feedthrough
rlabel pdiffusion 878 -1002 878 -1002 0 feedthrough
rlabel pdiffusion 885 -1002 885 -1002 0 cellNo=766
rlabel pdiffusion 892 -1002 892 -1002 0 feedthrough
rlabel pdiffusion 899 -1002 899 -1002 0 cellNo=831
rlabel pdiffusion 906 -1002 906 -1002 0 feedthrough
rlabel pdiffusion 913 -1002 913 -1002 0 feedthrough
rlabel pdiffusion 920 -1002 920 -1002 0 feedthrough
rlabel pdiffusion 927 -1002 927 -1002 0 feedthrough
rlabel pdiffusion 934 -1002 934 -1002 0 feedthrough
rlabel pdiffusion 941 -1002 941 -1002 0 feedthrough
rlabel pdiffusion 948 -1002 948 -1002 0 feedthrough
rlabel pdiffusion 955 -1002 955 -1002 0 feedthrough
rlabel pdiffusion 962 -1002 962 -1002 0 cellNo=368
rlabel pdiffusion 969 -1002 969 -1002 0 feedthrough
rlabel pdiffusion 976 -1002 976 -1002 0 cellNo=584
rlabel pdiffusion 983 -1002 983 -1002 0 cellNo=390
rlabel pdiffusion 990 -1002 990 -1002 0 cellNo=798
rlabel pdiffusion 997 -1002 997 -1002 0 cellNo=371
rlabel pdiffusion 1004 -1002 1004 -1002 0 feedthrough
rlabel pdiffusion 1011 -1002 1011 -1002 0 cellNo=784
rlabel pdiffusion 1018 -1002 1018 -1002 0 feedthrough
rlabel pdiffusion 1025 -1002 1025 -1002 0 feedthrough
rlabel pdiffusion 1032 -1002 1032 -1002 0 feedthrough
rlabel pdiffusion 1039 -1002 1039 -1002 0 feedthrough
rlabel pdiffusion 1046 -1002 1046 -1002 0 feedthrough
rlabel pdiffusion 1053 -1002 1053 -1002 0 feedthrough
rlabel pdiffusion 1060 -1002 1060 -1002 0 feedthrough
rlabel pdiffusion 1067 -1002 1067 -1002 0 feedthrough
rlabel pdiffusion 1074 -1002 1074 -1002 0 feedthrough
rlabel pdiffusion 1081 -1002 1081 -1002 0 feedthrough
rlabel pdiffusion 1088 -1002 1088 -1002 0 feedthrough
rlabel pdiffusion 1095 -1002 1095 -1002 0 feedthrough
rlabel pdiffusion 1102 -1002 1102 -1002 0 feedthrough
rlabel pdiffusion 1109 -1002 1109 -1002 0 cellNo=65
rlabel pdiffusion 1116 -1002 1116 -1002 0 feedthrough
rlabel pdiffusion 1123 -1002 1123 -1002 0 feedthrough
rlabel pdiffusion 1130 -1002 1130 -1002 0 feedthrough
rlabel pdiffusion 1137 -1002 1137 -1002 0 feedthrough
rlabel pdiffusion 1144 -1002 1144 -1002 0 feedthrough
rlabel pdiffusion 1151 -1002 1151 -1002 0 feedthrough
rlabel pdiffusion 1158 -1002 1158 -1002 0 feedthrough
rlabel pdiffusion 1165 -1002 1165 -1002 0 feedthrough
rlabel pdiffusion 1172 -1002 1172 -1002 0 feedthrough
rlabel pdiffusion 1179 -1002 1179 -1002 0 feedthrough
rlabel pdiffusion 1186 -1002 1186 -1002 0 feedthrough
rlabel pdiffusion 1193 -1002 1193 -1002 0 feedthrough
rlabel pdiffusion 1200 -1002 1200 -1002 0 feedthrough
rlabel pdiffusion 1207 -1002 1207 -1002 0 feedthrough
rlabel pdiffusion 1214 -1002 1214 -1002 0 feedthrough
rlabel pdiffusion 1221 -1002 1221 -1002 0 feedthrough
rlabel pdiffusion 1228 -1002 1228 -1002 0 feedthrough
rlabel pdiffusion 1235 -1002 1235 -1002 0 feedthrough
rlabel pdiffusion 1242 -1002 1242 -1002 0 feedthrough
rlabel pdiffusion 1249 -1002 1249 -1002 0 feedthrough
rlabel pdiffusion 1256 -1002 1256 -1002 0 feedthrough
rlabel pdiffusion 1263 -1002 1263 -1002 0 feedthrough
rlabel pdiffusion 1270 -1002 1270 -1002 0 feedthrough
rlabel pdiffusion 1277 -1002 1277 -1002 0 feedthrough
rlabel pdiffusion 1284 -1002 1284 -1002 0 feedthrough
rlabel pdiffusion 1291 -1002 1291 -1002 0 feedthrough
rlabel pdiffusion 1298 -1002 1298 -1002 0 feedthrough
rlabel pdiffusion 1305 -1002 1305 -1002 0 feedthrough
rlabel pdiffusion 1312 -1002 1312 -1002 0 feedthrough
rlabel pdiffusion 1319 -1002 1319 -1002 0 feedthrough
rlabel pdiffusion 1326 -1002 1326 -1002 0 feedthrough
rlabel pdiffusion 1333 -1002 1333 -1002 0 feedthrough
rlabel pdiffusion 1340 -1002 1340 -1002 0 feedthrough
rlabel pdiffusion 1347 -1002 1347 -1002 0 feedthrough
rlabel pdiffusion 1354 -1002 1354 -1002 0 feedthrough
rlabel pdiffusion 1361 -1002 1361 -1002 0 feedthrough
rlabel pdiffusion 1368 -1002 1368 -1002 0 feedthrough
rlabel pdiffusion 1375 -1002 1375 -1002 0 feedthrough
rlabel pdiffusion 1382 -1002 1382 -1002 0 feedthrough
rlabel pdiffusion 1389 -1002 1389 -1002 0 feedthrough
rlabel pdiffusion 1396 -1002 1396 -1002 0 feedthrough
rlabel pdiffusion 1403 -1002 1403 -1002 0 feedthrough
rlabel pdiffusion 1410 -1002 1410 -1002 0 feedthrough
rlabel pdiffusion 1417 -1002 1417 -1002 0 feedthrough
rlabel pdiffusion 1424 -1002 1424 -1002 0 feedthrough
rlabel pdiffusion 1431 -1002 1431 -1002 0 feedthrough
rlabel pdiffusion 1438 -1002 1438 -1002 0 feedthrough
rlabel pdiffusion 1445 -1002 1445 -1002 0 feedthrough
rlabel pdiffusion 1452 -1002 1452 -1002 0 feedthrough
rlabel pdiffusion 1459 -1002 1459 -1002 0 feedthrough
rlabel pdiffusion 1466 -1002 1466 -1002 0 feedthrough
rlabel pdiffusion 1473 -1002 1473 -1002 0 feedthrough
rlabel pdiffusion 1480 -1002 1480 -1002 0 feedthrough
rlabel pdiffusion 1487 -1002 1487 -1002 0 feedthrough
rlabel pdiffusion 1494 -1002 1494 -1002 0 feedthrough
rlabel pdiffusion 1501 -1002 1501 -1002 0 feedthrough
rlabel pdiffusion 1508 -1002 1508 -1002 0 feedthrough
rlabel pdiffusion 1515 -1002 1515 -1002 0 feedthrough
rlabel pdiffusion 1522 -1002 1522 -1002 0 feedthrough
rlabel pdiffusion 1529 -1002 1529 -1002 0 feedthrough
rlabel pdiffusion 1536 -1002 1536 -1002 0 feedthrough
rlabel pdiffusion 1543 -1002 1543 -1002 0 feedthrough
rlabel pdiffusion 1550 -1002 1550 -1002 0 cellNo=694
rlabel pdiffusion 1557 -1002 1557 -1002 0 feedthrough
rlabel pdiffusion 1564 -1002 1564 -1002 0 cellNo=836
rlabel pdiffusion 1571 -1002 1571 -1002 0 cellNo=837
rlabel pdiffusion 1578 -1002 1578 -1002 0 feedthrough
rlabel pdiffusion 1585 -1002 1585 -1002 0 feedthrough
rlabel pdiffusion 1592 -1002 1592 -1002 0 feedthrough
rlabel pdiffusion 1599 -1002 1599 -1002 0 feedthrough
rlabel pdiffusion 1606 -1002 1606 -1002 0 feedthrough
rlabel pdiffusion 1613 -1002 1613 -1002 0 feedthrough
rlabel pdiffusion 1620 -1002 1620 -1002 0 feedthrough
rlabel pdiffusion 1627 -1002 1627 -1002 0 feedthrough
rlabel pdiffusion 1634 -1002 1634 -1002 0 feedthrough
rlabel pdiffusion 1739 -1002 1739 -1002 0 feedthrough
rlabel pdiffusion 3 -1103 3 -1103 0 cellNo=1069
rlabel pdiffusion 10 -1103 10 -1103 0 cellNo=1086
rlabel pdiffusion 17 -1103 17 -1103 0 cellNo=1103
rlabel pdiffusion 24 -1103 24 -1103 0 feedthrough
rlabel pdiffusion 31 -1103 31 -1103 0 feedthrough
rlabel pdiffusion 38 -1103 38 -1103 0 cellNo=1134
rlabel pdiffusion 45 -1103 45 -1103 0 feedthrough
rlabel pdiffusion 52 -1103 52 -1103 0 feedthrough
rlabel pdiffusion 59 -1103 59 -1103 0 feedthrough
rlabel pdiffusion 66 -1103 66 -1103 0 feedthrough
rlabel pdiffusion 73 -1103 73 -1103 0 cellNo=519
rlabel pdiffusion 80 -1103 80 -1103 0 feedthrough
rlabel pdiffusion 87 -1103 87 -1103 0 cellNo=583
rlabel pdiffusion 94 -1103 94 -1103 0 feedthrough
rlabel pdiffusion 101 -1103 101 -1103 0 feedthrough
rlabel pdiffusion 108 -1103 108 -1103 0 feedthrough
rlabel pdiffusion 115 -1103 115 -1103 0 feedthrough
rlabel pdiffusion 122 -1103 122 -1103 0 feedthrough
rlabel pdiffusion 129 -1103 129 -1103 0 feedthrough
rlabel pdiffusion 136 -1103 136 -1103 0 cellNo=998
rlabel pdiffusion 143 -1103 143 -1103 0 feedthrough
rlabel pdiffusion 150 -1103 150 -1103 0 feedthrough
rlabel pdiffusion 157 -1103 157 -1103 0 feedthrough
rlabel pdiffusion 164 -1103 164 -1103 0 feedthrough
rlabel pdiffusion 171 -1103 171 -1103 0 feedthrough
rlabel pdiffusion 178 -1103 178 -1103 0 feedthrough
rlabel pdiffusion 185 -1103 185 -1103 0 feedthrough
rlabel pdiffusion 192 -1103 192 -1103 0 feedthrough
rlabel pdiffusion 199 -1103 199 -1103 0 feedthrough
rlabel pdiffusion 206 -1103 206 -1103 0 feedthrough
rlabel pdiffusion 213 -1103 213 -1103 0 cellNo=185
rlabel pdiffusion 220 -1103 220 -1103 0 feedthrough
rlabel pdiffusion 227 -1103 227 -1103 0 feedthrough
rlabel pdiffusion 234 -1103 234 -1103 0 cellNo=281
rlabel pdiffusion 241 -1103 241 -1103 0 feedthrough
rlabel pdiffusion 248 -1103 248 -1103 0 cellNo=451
rlabel pdiffusion 255 -1103 255 -1103 0 feedthrough
rlabel pdiffusion 262 -1103 262 -1103 0 cellNo=431
rlabel pdiffusion 269 -1103 269 -1103 0 feedthrough
rlabel pdiffusion 276 -1103 276 -1103 0 feedthrough
rlabel pdiffusion 283 -1103 283 -1103 0 feedthrough
rlabel pdiffusion 290 -1103 290 -1103 0 feedthrough
rlabel pdiffusion 297 -1103 297 -1103 0 feedthrough
rlabel pdiffusion 304 -1103 304 -1103 0 feedthrough
rlabel pdiffusion 311 -1103 311 -1103 0 feedthrough
rlabel pdiffusion 318 -1103 318 -1103 0 feedthrough
rlabel pdiffusion 325 -1103 325 -1103 0 feedthrough
rlabel pdiffusion 332 -1103 332 -1103 0 feedthrough
rlabel pdiffusion 339 -1103 339 -1103 0 cellNo=594
rlabel pdiffusion 346 -1103 346 -1103 0 feedthrough
rlabel pdiffusion 353 -1103 353 -1103 0 feedthrough
rlabel pdiffusion 360 -1103 360 -1103 0 feedthrough
rlabel pdiffusion 367 -1103 367 -1103 0 feedthrough
rlabel pdiffusion 374 -1103 374 -1103 0 feedthrough
rlabel pdiffusion 381 -1103 381 -1103 0 feedthrough
rlabel pdiffusion 388 -1103 388 -1103 0 feedthrough
rlabel pdiffusion 395 -1103 395 -1103 0 cellNo=55
rlabel pdiffusion 402 -1103 402 -1103 0 feedthrough
rlabel pdiffusion 409 -1103 409 -1103 0 feedthrough
rlabel pdiffusion 416 -1103 416 -1103 0 feedthrough
rlabel pdiffusion 423 -1103 423 -1103 0 cellNo=397
rlabel pdiffusion 430 -1103 430 -1103 0 feedthrough
rlabel pdiffusion 437 -1103 437 -1103 0 feedthrough
rlabel pdiffusion 444 -1103 444 -1103 0 feedthrough
rlabel pdiffusion 451 -1103 451 -1103 0 feedthrough
rlabel pdiffusion 458 -1103 458 -1103 0 feedthrough
rlabel pdiffusion 465 -1103 465 -1103 0 feedthrough
rlabel pdiffusion 472 -1103 472 -1103 0 cellNo=285
rlabel pdiffusion 479 -1103 479 -1103 0 cellNo=106
rlabel pdiffusion 486 -1103 486 -1103 0 feedthrough
rlabel pdiffusion 493 -1103 493 -1103 0 feedthrough
rlabel pdiffusion 500 -1103 500 -1103 0 feedthrough
rlabel pdiffusion 507 -1103 507 -1103 0 feedthrough
rlabel pdiffusion 514 -1103 514 -1103 0 cellNo=490
rlabel pdiffusion 521 -1103 521 -1103 0 feedthrough
rlabel pdiffusion 528 -1103 528 -1103 0 feedthrough
rlabel pdiffusion 535 -1103 535 -1103 0 feedthrough
rlabel pdiffusion 542 -1103 542 -1103 0 feedthrough
rlabel pdiffusion 549 -1103 549 -1103 0 feedthrough
rlabel pdiffusion 556 -1103 556 -1103 0 feedthrough
rlabel pdiffusion 563 -1103 563 -1103 0 feedthrough
rlabel pdiffusion 570 -1103 570 -1103 0 feedthrough
rlabel pdiffusion 577 -1103 577 -1103 0 feedthrough
rlabel pdiffusion 584 -1103 584 -1103 0 feedthrough
rlabel pdiffusion 591 -1103 591 -1103 0 feedthrough
rlabel pdiffusion 598 -1103 598 -1103 0 feedthrough
rlabel pdiffusion 605 -1103 605 -1103 0 feedthrough
rlabel pdiffusion 612 -1103 612 -1103 0 feedthrough
rlabel pdiffusion 619 -1103 619 -1103 0 feedthrough
rlabel pdiffusion 626 -1103 626 -1103 0 cellNo=478
rlabel pdiffusion 633 -1103 633 -1103 0 feedthrough
rlabel pdiffusion 640 -1103 640 -1103 0 cellNo=690
rlabel pdiffusion 647 -1103 647 -1103 0 cellNo=133
rlabel pdiffusion 654 -1103 654 -1103 0 feedthrough
rlabel pdiffusion 661 -1103 661 -1103 0 feedthrough
rlabel pdiffusion 668 -1103 668 -1103 0 feedthrough
rlabel pdiffusion 675 -1103 675 -1103 0 cellNo=736
rlabel pdiffusion 682 -1103 682 -1103 0 feedthrough
rlabel pdiffusion 689 -1103 689 -1103 0 cellNo=121
rlabel pdiffusion 696 -1103 696 -1103 0 cellNo=820
rlabel pdiffusion 703 -1103 703 -1103 0 feedthrough
rlabel pdiffusion 710 -1103 710 -1103 0 feedthrough
rlabel pdiffusion 717 -1103 717 -1103 0 feedthrough
rlabel pdiffusion 724 -1103 724 -1103 0 feedthrough
rlabel pdiffusion 731 -1103 731 -1103 0 cellNo=572
rlabel pdiffusion 738 -1103 738 -1103 0 feedthrough
rlabel pdiffusion 745 -1103 745 -1103 0 feedthrough
rlabel pdiffusion 752 -1103 752 -1103 0 feedthrough
rlabel pdiffusion 759 -1103 759 -1103 0 feedthrough
rlabel pdiffusion 766 -1103 766 -1103 0 feedthrough
rlabel pdiffusion 773 -1103 773 -1103 0 feedthrough
rlabel pdiffusion 780 -1103 780 -1103 0 feedthrough
rlabel pdiffusion 787 -1103 787 -1103 0 feedthrough
rlabel pdiffusion 794 -1103 794 -1103 0 feedthrough
rlabel pdiffusion 801 -1103 801 -1103 0 cellNo=345
rlabel pdiffusion 808 -1103 808 -1103 0 feedthrough
rlabel pdiffusion 815 -1103 815 -1103 0 feedthrough
rlabel pdiffusion 822 -1103 822 -1103 0 feedthrough
rlabel pdiffusion 829 -1103 829 -1103 0 feedthrough
rlabel pdiffusion 836 -1103 836 -1103 0 feedthrough
rlabel pdiffusion 843 -1103 843 -1103 0 feedthrough
rlabel pdiffusion 850 -1103 850 -1103 0 feedthrough
rlabel pdiffusion 857 -1103 857 -1103 0 feedthrough
rlabel pdiffusion 864 -1103 864 -1103 0 cellNo=576
rlabel pdiffusion 871 -1103 871 -1103 0 feedthrough
rlabel pdiffusion 878 -1103 878 -1103 0 cellNo=550
rlabel pdiffusion 885 -1103 885 -1103 0 cellNo=361
rlabel pdiffusion 892 -1103 892 -1103 0 cellNo=365
rlabel pdiffusion 899 -1103 899 -1103 0 feedthrough
rlabel pdiffusion 906 -1103 906 -1103 0 feedthrough
rlabel pdiffusion 913 -1103 913 -1103 0 feedthrough
rlabel pdiffusion 920 -1103 920 -1103 0 feedthrough
rlabel pdiffusion 927 -1103 927 -1103 0 feedthrough
rlabel pdiffusion 934 -1103 934 -1103 0 feedthrough
rlabel pdiffusion 941 -1103 941 -1103 0 feedthrough
rlabel pdiffusion 948 -1103 948 -1103 0 feedthrough
rlabel pdiffusion 955 -1103 955 -1103 0 feedthrough
rlabel pdiffusion 962 -1103 962 -1103 0 feedthrough
rlabel pdiffusion 969 -1103 969 -1103 0 feedthrough
rlabel pdiffusion 976 -1103 976 -1103 0 feedthrough
rlabel pdiffusion 983 -1103 983 -1103 0 feedthrough
rlabel pdiffusion 990 -1103 990 -1103 0 feedthrough
rlabel pdiffusion 997 -1103 997 -1103 0 feedthrough
rlabel pdiffusion 1004 -1103 1004 -1103 0 cellNo=436
rlabel pdiffusion 1011 -1103 1011 -1103 0 feedthrough
rlabel pdiffusion 1018 -1103 1018 -1103 0 feedthrough
rlabel pdiffusion 1025 -1103 1025 -1103 0 feedthrough
rlabel pdiffusion 1032 -1103 1032 -1103 0 feedthrough
rlabel pdiffusion 1039 -1103 1039 -1103 0 feedthrough
rlabel pdiffusion 1046 -1103 1046 -1103 0 cellNo=47
rlabel pdiffusion 1053 -1103 1053 -1103 0 cellNo=497
rlabel pdiffusion 1060 -1103 1060 -1103 0 feedthrough
rlabel pdiffusion 1067 -1103 1067 -1103 0 feedthrough
rlabel pdiffusion 1074 -1103 1074 -1103 0 feedthrough
rlabel pdiffusion 1081 -1103 1081 -1103 0 feedthrough
rlabel pdiffusion 1088 -1103 1088 -1103 0 cellNo=212
rlabel pdiffusion 1095 -1103 1095 -1103 0 feedthrough
rlabel pdiffusion 1102 -1103 1102 -1103 0 feedthrough
rlabel pdiffusion 1109 -1103 1109 -1103 0 feedthrough
rlabel pdiffusion 1116 -1103 1116 -1103 0 feedthrough
rlabel pdiffusion 1123 -1103 1123 -1103 0 feedthrough
rlabel pdiffusion 1130 -1103 1130 -1103 0 feedthrough
rlabel pdiffusion 1137 -1103 1137 -1103 0 feedthrough
rlabel pdiffusion 1144 -1103 1144 -1103 0 feedthrough
rlabel pdiffusion 1151 -1103 1151 -1103 0 feedthrough
rlabel pdiffusion 1158 -1103 1158 -1103 0 feedthrough
rlabel pdiffusion 1165 -1103 1165 -1103 0 feedthrough
rlabel pdiffusion 1172 -1103 1172 -1103 0 feedthrough
rlabel pdiffusion 1179 -1103 1179 -1103 0 feedthrough
rlabel pdiffusion 1186 -1103 1186 -1103 0 feedthrough
rlabel pdiffusion 1193 -1103 1193 -1103 0 feedthrough
rlabel pdiffusion 1200 -1103 1200 -1103 0 feedthrough
rlabel pdiffusion 1207 -1103 1207 -1103 0 feedthrough
rlabel pdiffusion 1214 -1103 1214 -1103 0 feedthrough
rlabel pdiffusion 1221 -1103 1221 -1103 0 cellNo=729
rlabel pdiffusion 1228 -1103 1228 -1103 0 feedthrough
rlabel pdiffusion 1235 -1103 1235 -1103 0 feedthrough
rlabel pdiffusion 1242 -1103 1242 -1103 0 feedthrough
rlabel pdiffusion 1249 -1103 1249 -1103 0 feedthrough
rlabel pdiffusion 1256 -1103 1256 -1103 0 feedthrough
rlabel pdiffusion 1263 -1103 1263 -1103 0 feedthrough
rlabel pdiffusion 1270 -1103 1270 -1103 0 feedthrough
rlabel pdiffusion 1277 -1103 1277 -1103 0 feedthrough
rlabel pdiffusion 1284 -1103 1284 -1103 0 feedthrough
rlabel pdiffusion 1291 -1103 1291 -1103 0 feedthrough
rlabel pdiffusion 1298 -1103 1298 -1103 0 feedthrough
rlabel pdiffusion 1305 -1103 1305 -1103 0 feedthrough
rlabel pdiffusion 1312 -1103 1312 -1103 0 feedthrough
rlabel pdiffusion 1319 -1103 1319 -1103 0 feedthrough
rlabel pdiffusion 1326 -1103 1326 -1103 0 feedthrough
rlabel pdiffusion 1333 -1103 1333 -1103 0 feedthrough
rlabel pdiffusion 1340 -1103 1340 -1103 0 feedthrough
rlabel pdiffusion 1347 -1103 1347 -1103 0 feedthrough
rlabel pdiffusion 1354 -1103 1354 -1103 0 feedthrough
rlabel pdiffusion 1361 -1103 1361 -1103 0 feedthrough
rlabel pdiffusion 1368 -1103 1368 -1103 0 feedthrough
rlabel pdiffusion 1375 -1103 1375 -1103 0 feedthrough
rlabel pdiffusion 1382 -1103 1382 -1103 0 cellNo=824
rlabel pdiffusion 1389 -1103 1389 -1103 0 feedthrough
rlabel pdiffusion 1396 -1103 1396 -1103 0 feedthrough
rlabel pdiffusion 1403 -1103 1403 -1103 0 feedthrough
rlabel pdiffusion 1410 -1103 1410 -1103 0 feedthrough
rlabel pdiffusion 1417 -1103 1417 -1103 0 feedthrough
rlabel pdiffusion 1424 -1103 1424 -1103 0 feedthrough
rlabel pdiffusion 1431 -1103 1431 -1103 0 feedthrough
rlabel pdiffusion 1438 -1103 1438 -1103 0 feedthrough
rlabel pdiffusion 1445 -1103 1445 -1103 0 feedthrough
rlabel pdiffusion 1452 -1103 1452 -1103 0 cellNo=32
rlabel pdiffusion 1459 -1103 1459 -1103 0 feedthrough
rlabel pdiffusion 1466 -1103 1466 -1103 0 feedthrough
rlabel pdiffusion 1473 -1103 1473 -1103 0 cellNo=286
rlabel pdiffusion 1480 -1103 1480 -1103 0 feedthrough
rlabel pdiffusion 1487 -1103 1487 -1103 0 feedthrough
rlabel pdiffusion 1494 -1103 1494 -1103 0 cellNo=45
rlabel pdiffusion 1501 -1103 1501 -1103 0 feedthrough
rlabel pdiffusion 1508 -1103 1508 -1103 0 feedthrough
rlabel pdiffusion 1515 -1103 1515 -1103 0 feedthrough
rlabel pdiffusion 1522 -1103 1522 -1103 0 feedthrough
rlabel pdiffusion 1529 -1103 1529 -1103 0 feedthrough
rlabel pdiffusion 1536 -1103 1536 -1103 0 feedthrough
rlabel pdiffusion 1543 -1103 1543 -1103 0 feedthrough
rlabel pdiffusion 1550 -1103 1550 -1103 0 feedthrough
rlabel pdiffusion 1557 -1103 1557 -1103 0 feedthrough
rlabel pdiffusion 1564 -1103 1564 -1103 0 feedthrough
rlabel pdiffusion 1571 -1103 1571 -1103 0 feedthrough
rlabel pdiffusion 1578 -1103 1578 -1103 0 feedthrough
rlabel pdiffusion 1585 -1103 1585 -1103 0 feedthrough
rlabel pdiffusion 1592 -1103 1592 -1103 0 feedthrough
rlabel pdiffusion 1599 -1103 1599 -1103 0 feedthrough
rlabel pdiffusion 1606 -1103 1606 -1103 0 feedthrough
rlabel pdiffusion 1613 -1103 1613 -1103 0 feedthrough
rlabel pdiffusion 1620 -1103 1620 -1103 0 feedthrough
rlabel pdiffusion 1627 -1103 1627 -1103 0 feedthrough
rlabel pdiffusion 1634 -1103 1634 -1103 0 feedthrough
rlabel pdiffusion 1641 -1103 1641 -1103 0 feedthrough
rlabel pdiffusion 1648 -1103 1648 -1103 0 feedthrough
rlabel pdiffusion 1655 -1103 1655 -1103 0 feedthrough
rlabel pdiffusion 1676 -1103 1676 -1103 0 feedthrough
rlabel pdiffusion 1683 -1103 1683 -1103 0 feedthrough
rlabel pdiffusion 1746 -1103 1746 -1103 0 feedthrough
rlabel pdiffusion 3 -1222 3 -1222 0 cellNo=1084
rlabel pdiffusion 10 -1222 10 -1222 0 cellNo=1102
rlabel pdiffusion 17 -1222 17 -1222 0 cellNo=1110
rlabel pdiffusion 24 -1222 24 -1222 0 feedthrough
rlabel pdiffusion 31 -1222 31 -1222 0 feedthrough
rlabel pdiffusion 38 -1222 38 -1222 0 feedthrough
rlabel pdiffusion 45 -1222 45 -1222 0 feedthrough
rlabel pdiffusion 52 -1222 52 -1222 0 feedthrough
rlabel pdiffusion 59 -1222 59 -1222 0 feedthrough
rlabel pdiffusion 66 -1222 66 -1222 0 cellNo=968
rlabel pdiffusion 73 -1222 73 -1222 0 feedthrough
rlabel pdiffusion 80 -1222 80 -1222 0 feedthrough
rlabel pdiffusion 87 -1222 87 -1222 0 cellNo=423
rlabel pdiffusion 94 -1222 94 -1222 0 feedthrough
rlabel pdiffusion 101 -1222 101 -1222 0 feedthrough
rlabel pdiffusion 108 -1222 108 -1222 0 cellNo=574
rlabel pdiffusion 115 -1222 115 -1222 0 feedthrough
rlabel pdiffusion 122 -1222 122 -1222 0 cellNo=6
rlabel pdiffusion 129 -1222 129 -1222 0 feedthrough
rlabel pdiffusion 136 -1222 136 -1222 0 feedthrough
rlabel pdiffusion 143 -1222 143 -1222 0 cellNo=722
rlabel pdiffusion 150 -1222 150 -1222 0 feedthrough
rlabel pdiffusion 157 -1222 157 -1222 0 feedthrough
rlabel pdiffusion 164 -1222 164 -1222 0 feedthrough
rlabel pdiffusion 171 -1222 171 -1222 0 cellNo=223
rlabel pdiffusion 178 -1222 178 -1222 0 cellNo=737
rlabel pdiffusion 185 -1222 185 -1222 0 feedthrough
rlabel pdiffusion 192 -1222 192 -1222 0 feedthrough
rlabel pdiffusion 199 -1222 199 -1222 0 feedthrough
rlabel pdiffusion 206 -1222 206 -1222 0 feedthrough
rlabel pdiffusion 213 -1222 213 -1222 0 feedthrough
rlabel pdiffusion 220 -1222 220 -1222 0 feedthrough
rlabel pdiffusion 227 -1222 227 -1222 0 cellNo=31
rlabel pdiffusion 234 -1222 234 -1222 0 feedthrough
rlabel pdiffusion 241 -1222 241 -1222 0 cellNo=777
rlabel pdiffusion 248 -1222 248 -1222 0 feedthrough
rlabel pdiffusion 255 -1222 255 -1222 0 feedthrough
rlabel pdiffusion 262 -1222 262 -1222 0 cellNo=411
rlabel pdiffusion 269 -1222 269 -1222 0 feedthrough
rlabel pdiffusion 276 -1222 276 -1222 0 feedthrough
rlabel pdiffusion 283 -1222 283 -1222 0 feedthrough
rlabel pdiffusion 290 -1222 290 -1222 0 feedthrough
rlabel pdiffusion 297 -1222 297 -1222 0 feedthrough
rlabel pdiffusion 304 -1222 304 -1222 0 feedthrough
rlabel pdiffusion 311 -1222 311 -1222 0 feedthrough
rlabel pdiffusion 318 -1222 318 -1222 0 feedthrough
rlabel pdiffusion 325 -1222 325 -1222 0 feedthrough
rlabel pdiffusion 332 -1222 332 -1222 0 feedthrough
rlabel pdiffusion 339 -1222 339 -1222 0 feedthrough
rlabel pdiffusion 346 -1222 346 -1222 0 feedthrough
rlabel pdiffusion 353 -1222 353 -1222 0 feedthrough
rlabel pdiffusion 360 -1222 360 -1222 0 feedthrough
rlabel pdiffusion 367 -1222 367 -1222 0 feedthrough
rlabel pdiffusion 374 -1222 374 -1222 0 feedthrough
rlabel pdiffusion 381 -1222 381 -1222 0 feedthrough
rlabel pdiffusion 388 -1222 388 -1222 0 feedthrough
rlabel pdiffusion 395 -1222 395 -1222 0 feedthrough
rlabel pdiffusion 402 -1222 402 -1222 0 feedthrough
rlabel pdiffusion 409 -1222 409 -1222 0 feedthrough
rlabel pdiffusion 416 -1222 416 -1222 0 feedthrough
rlabel pdiffusion 423 -1222 423 -1222 0 feedthrough
rlabel pdiffusion 430 -1222 430 -1222 0 feedthrough
rlabel pdiffusion 437 -1222 437 -1222 0 cellNo=90
rlabel pdiffusion 444 -1222 444 -1222 0 feedthrough
rlabel pdiffusion 451 -1222 451 -1222 0 feedthrough
rlabel pdiffusion 458 -1222 458 -1222 0 feedthrough
rlabel pdiffusion 465 -1222 465 -1222 0 feedthrough
rlabel pdiffusion 472 -1222 472 -1222 0 feedthrough
rlabel pdiffusion 479 -1222 479 -1222 0 feedthrough
rlabel pdiffusion 486 -1222 486 -1222 0 feedthrough
rlabel pdiffusion 493 -1222 493 -1222 0 feedthrough
rlabel pdiffusion 500 -1222 500 -1222 0 feedthrough
rlabel pdiffusion 507 -1222 507 -1222 0 cellNo=900
rlabel pdiffusion 514 -1222 514 -1222 0 feedthrough
rlabel pdiffusion 521 -1222 521 -1222 0 feedthrough
rlabel pdiffusion 528 -1222 528 -1222 0 feedthrough
rlabel pdiffusion 535 -1222 535 -1222 0 feedthrough
rlabel pdiffusion 542 -1222 542 -1222 0 cellNo=617
rlabel pdiffusion 549 -1222 549 -1222 0 feedthrough
rlabel pdiffusion 556 -1222 556 -1222 0 feedthrough
rlabel pdiffusion 563 -1222 563 -1222 0 cellNo=389
rlabel pdiffusion 570 -1222 570 -1222 0 feedthrough
rlabel pdiffusion 577 -1222 577 -1222 0 feedthrough
rlabel pdiffusion 584 -1222 584 -1222 0 feedthrough
rlabel pdiffusion 591 -1222 591 -1222 0 feedthrough
rlabel pdiffusion 598 -1222 598 -1222 0 cellNo=63
rlabel pdiffusion 605 -1222 605 -1222 0 cellNo=314
rlabel pdiffusion 612 -1222 612 -1222 0 feedthrough
rlabel pdiffusion 619 -1222 619 -1222 0 feedthrough
rlabel pdiffusion 626 -1222 626 -1222 0 feedthrough
rlabel pdiffusion 633 -1222 633 -1222 0 cellNo=77
rlabel pdiffusion 640 -1222 640 -1222 0 feedthrough
rlabel pdiffusion 647 -1222 647 -1222 0 cellNo=237
rlabel pdiffusion 654 -1222 654 -1222 0 cellNo=923
rlabel pdiffusion 661 -1222 661 -1222 0 feedthrough
rlabel pdiffusion 668 -1222 668 -1222 0 feedthrough
rlabel pdiffusion 675 -1222 675 -1222 0 feedthrough
rlabel pdiffusion 682 -1222 682 -1222 0 feedthrough
rlabel pdiffusion 689 -1222 689 -1222 0 feedthrough
rlabel pdiffusion 696 -1222 696 -1222 0 cellNo=529
rlabel pdiffusion 703 -1222 703 -1222 0 cellNo=206
rlabel pdiffusion 710 -1222 710 -1222 0 feedthrough
rlabel pdiffusion 717 -1222 717 -1222 0 feedthrough
rlabel pdiffusion 724 -1222 724 -1222 0 feedthrough
rlabel pdiffusion 731 -1222 731 -1222 0 feedthrough
rlabel pdiffusion 738 -1222 738 -1222 0 cellNo=433
rlabel pdiffusion 745 -1222 745 -1222 0 feedthrough
rlabel pdiffusion 752 -1222 752 -1222 0 feedthrough
rlabel pdiffusion 759 -1222 759 -1222 0 feedthrough
rlabel pdiffusion 766 -1222 766 -1222 0 cellNo=19
rlabel pdiffusion 773 -1222 773 -1222 0 feedthrough
rlabel pdiffusion 780 -1222 780 -1222 0 feedthrough
rlabel pdiffusion 787 -1222 787 -1222 0 feedthrough
rlabel pdiffusion 794 -1222 794 -1222 0 cellNo=240
rlabel pdiffusion 801 -1222 801 -1222 0 feedthrough
rlabel pdiffusion 808 -1222 808 -1222 0 feedthrough
rlabel pdiffusion 815 -1222 815 -1222 0 cellNo=546
rlabel pdiffusion 822 -1222 822 -1222 0 cellNo=524
rlabel pdiffusion 829 -1222 829 -1222 0 cellNo=642
rlabel pdiffusion 836 -1222 836 -1222 0 feedthrough
rlabel pdiffusion 843 -1222 843 -1222 0 feedthrough
rlabel pdiffusion 850 -1222 850 -1222 0 feedthrough
rlabel pdiffusion 857 -1222 857 -1222 0 cellNo=183
rlabel pdiffusion 864 -1222 864 -1222 0 feedthrough
rlabel pdiffusion 871 -1222 871 -1222 0 feedthrough
rlabel pdiffusion 878 -1222 878 -1222 0 feedthrough
rlabel pdiffusion 885 -1222 885 -1222 0 feedthrough
rlabel pdiffusion 892 -1222 892 -1222 0 cellNo=503
rlabel pdiffusion 899 -1222 899 -1222 0 feedthrough
rlabel pdiffusion 906 -1222 906 -1222 0 feedthrough
rlabel pdiffusion 913 -1222 913 -1222 0 feedthrough
rlabel pdiffusion 920 -1222 920 -1222 0 feedthrough
rlabel pdiffusion 927 -1222 927 -1222 0 cellNo=604
rlabel pdiffusion 934 -1222 934 -1222 0 feedthrough
rlabel pdiffusion 941 -1222 941 -1222 0 feedthrough
rlabel pdiffusion 948 -1222 948 -1222 0 cellNo=448
rlabel pdiffusion 955 -1222 955 -1222 0 feedthrough
rlabel pdiffusion 962 -1222 962 -1222 0 feedthrough
rlabel pdiffusion 969 -1222 969 -1222 0 feedthrough
rlabel pdiffusion 976 -1222 976 -1222 0 feedthrough
rlabel pdiffusion 983 -1222 983 -1222 0 feedthrough
rlabel pdiffusion 990 -1222 990 -1222 0 feedthrough
rlabel pdiffusion 997 -1222 997 -1222 0 feedthrough
rlabel pdiffusion 1004 -1222 1004 -1222 0 feedthrough
rlabel pdiffusion 1011 -1222 1011 -1222 0 feedthrough
rlabel pdiffusion 1018 -1222 1018 -1222 0 feedthrough
rlabel pdiffusion 1025 -1222 1025 -1222 0 feedthrough
rlabel pdiffusion 1032 -1222 1032 -1222 0 feedthrough
rlabel pdiffusion 1039 -1222 1039 -1222 0 feedthrough
rlabel pdiffusion 1046 -1222 1046 -1222 0 feedthrough
rlabel pdiffusion 1053 -1222 1053 -1222 0 cellNo=538
rlabel pdiffusion 1060 -1222 1060 -1222 0 feedthrough
rlabel pdiffusion 1067 -1222 1067 -1222 0 feedthrough
rlabel pdiffusion 1074 -1222 1074 -1222 0 feedthrough
rlabel pdiffusion 1081 -1222 1081 -1222 0 feedthrough
rlabel pdiffusion 1088 -1222 1088 -1222 0 feedthrough
rlabel pdiffusion 1095 -1222 1095 -1222 0 feedthrough
rlabel pdiffusion 1102 -1222 1102 -1222 0 feedthrough
rlabel pdiffusion 1109 -1222 1109 -1222 0 feedthrough
rlabel pdiffusion 1116 -1222 1116 -1222 0 feedthrough
rlabel pdiffusion 1123 -1222 1123 -1222 0 feedthrough
rlabel pdiffusion 1130 -1222 1130 -1222 0 feedthrough
rlabel pdiffusion 1137 -1222 1137 -1222 0 feedthrough
rlabel pdiffusion 1144 -1222 1144 -1222 0 feedthrough
rlabel pdiffusion 1151 -1222 1151 -1222 0 feedthrough
rlabel pdiffusion 1158 -1222 1158 -1222 0 feedthrough
rlabel pdiffusion 1165 -1222 1165 -1222 0 feedthrough
rlabel pdiffusion 1172 -1222 1172 -1222 0 feedthrough
rlabel pdiffusion 1179 -1222 1179 -1222 0 feedthrough
rlabel pdiffusion 1186 -1222 1186 -1222 0 feedthrough
rlabel pdiffusion 1193 -1222 1193 -1222 0 feedthrough
rlabel pdiffusion 1200 -1222 1200 -1222 0 feedthrough
rlabel pdiffusion 1207 -1222 1207 -1222 0 feedthrough
rlabel pdiffusion 1214 -1222 1214 -1222 0 feedthrough
rlabel pdiffusion 1221 -1222 1221 -1222 0 feedthrough
rlabel pdiffusion 1228 -1222 1228 -1222 0 feedthrough
rlabel pdiffusion 1235 -1222 1235 -1222 0 feedthrough
rlabel pdiffusion 1242 -1222 1242 -1222 0 feedthrough
rlabel pdiffusion 1249 -1222 1249 -1222 0 feedthrough
rlabel pdiffusion 1256 -1222 1256 -1222 0 feedthrough
rlabel pdiffusion 1263 -1222 1263 -1222 0 feedthrough
rlabel pdiffusion 1270 -1222 1270 -1222 0 feedthrough
rlabel pdiffusion 1277 -1222 1277 -1222 0 feedthrough
rlabel pdiffusion 1284 -1222 1284 -1222 0 feedthrough
rlabel pdiffusion 1291 -1222 1291 -1222 0 feedthrough
rlabel pdiffusion 1298 -1222 1298 -1222 0 feedthrough
rlabel pdiffusion 1305 -1222 1305 -1222 0 feedthrough
rlabel pdiffusion 1312 -1222 1312 -1222 0 feedthrough
rlabel pdiffusion 1319 -1222 1319 -1222 0 feedthrough
rlabel pdiffusion 1326 -1222 1326 -1222 0 feedthrough
rlabel pdiffusion 1333 -1222 1333 -1222 0 feedthrough
rlabel pdiffusion 1340 -1222 1340 -1222 0 feedthrough
rlabel pdiffusion 1347 -1222 1347 -1222 0 feedthrough
rlabel pdiffusion 1354 -1222 1354 -1222 0 feedthrough
rlabel pdiffusion 1361 -1222 1361 -1222 0 feedthrough
rlabel pdiffusion 1368 -1222 1368 -1222 0 feedthrough
rlabel pdiffusion 1375 -1222 1375 -1222 0 feedthrough
rlabel pdiffusion 1382 -1222 1382 -1222 0 feedthrough
rlabel pdiffusion 1389 -1222 1389 -1222 0 feedthrough
rlabel pdiffusion 1396 -1222 1396 -1222 0 feedthrough
rlabel pdiffusion 1403 -1222 1403 -1222 0 feedthrough
rlabel pdiffusion 1410 -1222 1410 -1222 0 feedthrough
rlabel pdiffusion 1417 -1222 1417 -1222 0 feedthrough
rlabel pdiffusion 1424 -1222 1424 -1222 0 feedthrough
rlabel pdiffusion 1431 -1222 1431 -1222 0 feedthrough
rlabel pdiffusion 1438 -1222 1438 -1222 0 feedthrough
rlabel pdiffusion 1445 -1222 1445 -1222 0 feedthrough
rlabel pdiffusion 1452 -1222 1452 -1222 0 feedthrough
rlabel pdiffusion 1459 -1222 1459 -1222 0 feedthrough
rlabel pdiffusion 1466 -1222 1466 -1222 0 feedthrough
rlabel pdiffusion 1473 -1222 1473 -1222 0 feedthrough
rlabel pdiffusion 1480 -1222 1480 -1222 0 feedthrough
rlabel pdiffusion 1487 -1222 1487 -1222 0 feedthrough
rlabel pdiffusion 1494 -1222 1494 -1222 0 feedthrough
rlabel pdiffusion 1501 -1222 1501 -1222 0 feedthrough
rlabel pdiffusion 1508 -1222 1508 -1222 0 feedthrough
rlabel pdiffusion 1515 -1222 1515 -1222 0 feedthrough
rlabel pdiffusion 1522 -1222 1522 -1222 0 feedthrough
rlabel pdiffusion 1529 -1222 1529 -1222 0 feedthrough
rlabel pdiffusion 1536 -1222 1536 -1222 0 feedthrough
rlabel pdiffusion 1543 -1222 1543 -1222 0 feedthrough
rlabel pdiffusion 1550 -1222 1550 -1222 0 feedthrough
rlabel pdiffusion 1557 -1222 1557 -1222 0 feedthrough
rlabel pdiffusion 1564 -1222 1564 -1222 0 feedthrough
rlabel pdiffusion 1571 -1222 1571 -1222 0 feedthrough
rlabel pdiffusion 1578 -1222 1578 -1222 0 feedthrough
rlabel pdiffusion 1585 -1222 1585 -1222 0 feedthrough
rlabel pdiffusion 1592 -1222 1592 -1222 0 feedthrough
rlabel pdiffusion 1599 -1222 1599 -1222 0 feedthrough
rlabel pdiffusion 1606 -1222 1606 -1222 0 feedthrough
rlabel pdiffusion 1613 -1222 1613 -1222 0 feedthrough
rlabel pdiffusion 1620 -1222 1620 -1222 0 feedthrough
rlabel pdiffusion 1627 -1222 1627 -1222 0 feedthrough
rlabel pdiffusion 1634 -1222 1634 -1222 0 feedthrough
rlabel pdiffusion 1641 -1222 1641 -1222 0 feedthrough
rlabel pdiffusion 1648 -1222 1648 -1222 0 feedthrough
rlabel pdiffusion 1655 -1222 1655 -1222 0 feedthrough
rlabel pdiffusion 1662 -1222 1662 -1222 0 feedthrough
rlabel pdiffusion 1669 -1222 1669 -1222 0 feedthrough
rlabel pdiffusion 1676 -1222 1676 -1222 0 feedthrough
rlabel pdiffusion 1683 -1222 1683 -1222 0 feedthrough
rlabel pdiffusion 1690 -1222 1690 -1222 0 feedthrough
rlabel pdiffusion 1697 -1222 1697 -1222 0 feedthrough
rlabel pdiffusion 1704 -1222 1704 -1222 0 feedthrough
rlabel pdiffusion 1711 -1222 1711 -1222 0 feedthrough
rlabel pdiffusion 1718 -1222 1718 -1222 0 feedthrough
rlabel pdiffusion 1725 -1222 1725 -1222 0 feedthrough
rlabel pdiffusion 1732 -1222 1732 -1222 0 feedthrough
rlabel pdiffusion 1739 -1222 1739 -1222 0 feedthrough
rlabel pdiffusion 1746 -1222 1746 -1222 0 cellNo=395
rlabel pdiffusion 1753 -1222 1753 -1222 0 feedthrough
rlabel pdiffusion 1760 -1222 1760 -1222 0 feedthrough
rlabel pdiffusion 1767 -1222 1767 -1222 0 cellNo=279
rlabel pdiffusion 1774 -1222 1774 -1222 0 cellNo=340
rlabel pdiffusion 1781 -1222 1781 -1222 0 feedthrough
rlabel pdiffusion 1788 -1222 1788 -1222 0 feedthrough
rlabel pdiffusion 3 -1365 3 -1365 0 cellNo=1101
rlabel pdiffusion 10 -1365 10 -1365 0 cellNo=1109
rlabel pdiffusion 17 -1365 17 -1365 0 feedthrough
rlabel pdiffusion 24 -1365 24 -1365 0 feedthrough
rlabel pdiffusion 31 -1365 31 -1365 0 feedthrough
rlabel pdiffusion 38 -1365 38 -1365 0 cellNo=1123
rlabel pdiffusion 45 -1365 45 -1365 0 feedthrough
rlabel pdiffusion 52 -1365 52 -1365 0 cellNo=966
rlabel pdiffusion 59 -1365 59 -1365 0 cellNo=607
rlabel pdiffusion 66 -1365 66 -1365 0 feedthrough
rlabel pdiffusion 73 -1365 73 -1365 0 feedthrough
rlabel pdiffusion 80 -1365 80 -1365 0 cellNo=36
rlabel pdiffusion 87 -1365 87 -1365 0 feedthrough
rlabel pdiffusion 94 -1365 94 -1365 0 feedthrough
rlabel pdiffusion 101 -1365 101 -1365 0 cellNo=889
rlabel pdiffusion 108 -1365 108 -1365 0 cellNo=17
rlabel pdiffusion 115 -1365 115 -1365 0 feedthrough
rlabel pdiffusion 122 -1365 122 -1365 0 feedthrough
rlabel pdiffusion 129 -1365 129 -1365 0 cellNo=488
rlabel pdiffusion 136 -1365 136 -1365 0 feedthrough
rlabel pdiffusion 143 -1365 143 -1365 0 feedthrough
rlabel pdiffusion 150 -1365 150 -1365 0 feedthrough
rlabel pdiffusion 157 -1365 157 -1365 0 feedthrough
rlabel pdiffusion 164 -1365 164 -1365 0 feedthrough
rlabel pdiffusion 171 -1365 171 -1365 0 feedthrough
rlabel pdiffusion 178 -1365 178 -1365 0 feedthrough
rlabel pdiffusion 185 -1365 185 -1365 0 cellNo=76
rlabel pdiffusion 192 -1365 192 -1365 0 feedthrough
rlabel pdiffusion 199 -1365 199 -1365 0 cellNo=177
rlabel pdiffusion 206 -1365 206 -1365 0 cellNo=224
rlabel pdiffusion 213 -1365 213 -1365 0 feedthrough
rlabel pdiffusion 220 -1365 220 -1365 0 cellNo=405
rlabel pdiffusion 227 -1365 227 -1365 0 feedthrough
rlabel pdiffusion 234 -1365 234 -1365 0 feedthrough
rlabel pdiffusion 241 -1365 241 -1365 0 feedthrough
rlabel pdiffusion 248 -1365 248 -1365 0 feedthrough
rlabel pdiffusion 255 -1365 255 -1365 0 feedthrough
rlabel pdiffusion 262 -1365 262 -1365 0 feedthrough
rlabel pdiffusion 269 -1365 269 -1365 0 feedthrough
rlabel pdiffusion 276 -1365 276 -1365 0 feedthrough
rlabel pdiffusion 283 -1365 283 -1365 0 feedthrough
rlabel pdiffusion 290 -1365 290 -1365 0 cellNo=3
rlabel pdiffusion 297 -1365 297 -1365 0 feedthrough
rlabel pdiffusion 304 -1365 304 -1365 0 feedthrough
rlabel pdiffusion 311 -1365 311 -1365 0 feedthrough
rlabel pdiffusion 318 -1365 318 -1365 0 feedthrough
rlabel pdiffusion 325 -1365 325 -1365 0 feedthrough
rlabel pdiffusion 332 -1365 332 -1365 0 feedthrough
rlabel pdiffusion 339 -1365 339 -1365 0 feedthrough
rlabel pdiffusion 346 -1365 346 -1365 0 feedthrough
rlabel pdiffusion 353 -1365 353 -1365 0 feedthrough
rlabel pdiffusion 360 -1365 360 -1365 0 feedthrough
rlabel pdiffusion 367 -1365 367 -1365 0 feedthrough
rlabel pdiffusion 374 -1365 374 -1365 0 feedthrough
rlabel pdiffusion 381 -1365 381 -1365 0 feedthrough
rlabel pdiffusion 388 -1365 388 -1365 0 feedthrough
rlabel pdiffusion 395 -1365 395 -1365 0 feedthrough
rlabel pdiffusion 402 -1365 402 -1365 0 feedthrough
rlabel pdiffusion 409 -1365 409 -1365 0 feedthrough
rlabel pdiffusion 416 -1365 416 -1365 0 feedthrough
rlabel pdiffusion 423 -1365 423 -1365 0 feedthrough
rlabel pdiffusion 430 -1365 430 -1365 0 feedthrough
rlabel pdiffusion 437 -1365 437 -1365 0 feedthrough
rlabel pdiffusion 444 -1365 444 -1365 0 cellNo=866
rlabel pdiffusion 451 -1365 451 -1365 0 cellNo=811
rlabel pdiffusion 458 -1365 458 -1365 0 feedthrough
rlabel pdiffusion 465 -1365 465 -1365 0 feedthrough
rlabel pdiffusion 472 -1365 472 -1365 0 feedthrough
rlabel pdiffusion 479 -1365 479 -1365 0 feedthrough
rlabel pdiffusion 486 -1365 486 -1365 0 feedthrough
rlabel pdiffusion 493 -1365 493 -1365 0 feedthrough
rlabel pdiffusion 500 -1365 500 -1365 0 feedthrough
rlabel pdiffusion 507 -1365 507 -1365 0 feedthrough
rlabel pdiffusion 514 -1365 514 -1365 0 feedthrough
rlabel pdiffusion 521 -1365 521 -1365 0 feedthrough
rlabel pdiffusion 528 -1365 528 -1365 0 feedthrough
rlabel pdiffusion 535 -1365 535 -1365 0 feedthrough
rlabel pdiffusion 542 -1365 542 -1365 0 feedthrough
rlabel pdiffusion 549 -1365 549 -1365 0 cellNo=704
rlabel pdiffusion 556 -1365 556 -1365 0 cellNo=800
rlabel pdiffusion 563 -1365 563 -1365 0 cellNo=516
rlabel pdiffusion 570 -1365 570 -1365 0 cellNo=988
rlabel pdiffusion 577 -1365 577 -1365 0 feedthrough
rlabel pdiffusion 584 -1365 584 -1365 0 feedthrough
rlabel pdiffusion 591 -1365 591 -1365 0 feedthrough
rlabel pdiffusion 598 -1365 598 -1365 0 cellNo=466
rlabel pdiffusion 605 -1365 605 -1365 0 feedthrough
rlabel pdiffusion 612 -1365 612 -1365 0 feedthrough
rlabel pdiffusion 619 -1365 619 -1365 0 feedthrough
rlabel pdiffusion 626 -1365 626 -1365 0 feedthrough
rlabel pdiffusion 633 -1365 633 -1365 0 feedthrough
rlabel pdiffusion 640 -1365 640 -1365 0 feedthrough
rlabel pdiffusion 647 -1365 647 -1365 0 feedthrough
rlabel pdiffusion 654 -1365 654 -1365 0 feedthrough
rlabel pdiffusion 661 -1365 661 -1365 0 feedthrough
rlabel pdiffusion 668 -1365 668 -1365 0 feedthrough
rlabel pdiffusion 675 -1365 675 -1365 0 feedthrough
rlabel pdiffusion 682 -1365 682 -1365 0 feedthrough
rlabel pdiffusion 689 -1365 689 -1365 0 feedthrough
rlabel pdiffusion 696 -1365 696 -1365 0 feedthrough
rlabel pdiffusion 703 -1365 703 -1365 0 feedthrough
rlabel pdiffusion 710 -1365 710 -1365 0 feedthrough
rlabel pdiffusion 717 -1365 717 -1365 0 feedthrough
rlabel pdiffusion 724 -1365 724 -1365 0 feedthrough
rlabel pdiffusion 731 -1365 731 -1365 0 feedthrough
rlabel pdiffusion 738 -1365 738 -1365 0 cellNo=239
rlabel pdiffusion 745 -1365 745 -1365 0 feedthrough
rlabel pdiffusion 752 -1365 752 -1365 0 cellNo=187
rlabel pdiffusion 759 -1365 759 -1365 0 feedthrough
rlabel pdiffusion 766 -1365 766 -1365 0 feedthrough
rlabel pdiffusion 773 -1365 773 -1365 0 feedthrough
rlabel pdiffusion 780 -1365 780 -1365 0 feedthrough
rlabel pdiffusion 787 -1365 787 -1365 0 cellNo=873
rlabel pdiffusion 794 -1365 794 -1365 0 feedthrough
rlabel pdiffusion 801 -1365 801 -1365 0 feedthrough
rlabel pdiffusion 808 -1365 808 -1365 0 feedthrough
rlabel pdiffusion 815 -1365 815 -1365 0 cellNo=251
rlabel pdiffusion 822 -1365 822 -1365 0 cellNo=512
rlabel pdiffusion 829 -1365 829 -1365 0 cellNo=312
rlabel pdiffusion 836 -1365 836 -1365 0 feedthrough
rlabel pdiffusion 843 -1365 843 -1365 0 feedthrough
rlabel pdiffusion 850 -1365 850 -1365 0 cellNo=364
rlabel pdiffusion 857 -1365 857 -1365 0 feedthrough
rlabel pdiffusion 864 -1365 864 -1365 0 feedthrough
rlabel pdiffusion 871 -1365 871 -1365 0 feedthrough
rlabel pdiffusion 878 -1365 878 -1365 0 feedthrough
rlabel pdiffusion 885 -1365 885 -1365 0 feedthrough
rlabel pdiffusion 892 -1365 892 -1365 0 feedthrough
rlabel pdiffusion 899 -1365 899 -1365 0 feedthrough
rlabel pdiffusion 906 -1365 906 -1365 0 feedthrough
rlabel pdiffusion 913 -1365 913 -1365 0 feedthrough
rlabel pdiffusion 920 -1365 920 -1365 0 cellNo=721
rlabel pdiffusion 927 -1365 927 -1365 0 feedthrough
rlabel pdiffusion 934 -1365 934 -1365 0 cellNo=823
rlabel pdiffusion 941 -1365 941 -1365 0 feedthrough
rlabel pdiffusion 948 -1365 948 -1365 0 cellNo=391
rlabel pdiffusion 955 -1365 955 -1365 0 feedthrough
rlabel pdiffusion 962 -1365 962 -1365 0 feedthrough
rlabel pdiffusion 969 -1365 969 -1365 0 feedthrough
rlabel pdiffusion 976 -1365 976 -1365 0 feedthrough
rlabel pdiffusion 983 -1365 983 -1365 0 cellNo=669
rlabel pdiffusion 990 -1365 990 -1365 0 feedthrough
rlabel pdiffusion 997 -1365 997 -1365 0 feedthrough
rlabel pdiffusion 1004 -1365 1004 -1365 0 cellNo=42
rlabel pdiffusion 1011 -1365 1011 -1365 0 feedthrough
rlabel pdiffusion 1018 -1365 1018 -1365 0 cellNo=14
rlabel pdiffusion 1025 -1365 1025 -1365 0 feedthrough
rlabel pdiffusion 1032 -1365 1032 -1365 0 feedthrough
rlabel pdiffusion 1039 -1365 1039 -1365 0 feedthrough
rlabel pdiffusion 1046 -1365 1046 -1365 0 feedthrough
rlabel pdiffusion 1053 -1365 1053 -1365 0 feedthrough
rlabel pdiffusion 1060 -1365 1060 -1365 0 feedthrough
rlabel pdiffusion 1067 -1365 1067 -1365 0 feedthrough
rlabel pdiffusion 1074 -1365 1074 -1365 0 feedthrough
rlabel pdiffusion 1081 -1365 1081 -1365 0 feedthrough
rlabel pdiffusion 1088 -1365 1088 -1365 0 feedthrough
rlabel pdiffusion 1095 -1365 1095 -1365 0 feedthrough
rlabel pdiffusion 1102 -1365 1102 -1365 0 cellNo=830
rlabel pdiffusion 1109 -1365 1109 -1365 0 feedthrough
rlabel pdiffusion 1116 -1365 1116 -1365 0 feedthrough
rlabel pdiffusion 1123 -1365 1123 -1365 0 feedthrough
rlabel pdiffusion 1130 -1365 1130 -1365 0 feedthrough
rlabel pdiffusion 1137 -1365 1137 -1365 0 feedthrough
rlabel pdiffusion 1144 -1365 1144 -1365 0 cellNo=764
rlabel pdiffusion 1151 -1365 1151 -1365 0 feedthrough
rlabel pdiffusion 1158 -1365 1158 -1365 0 feedthrough
rlabel pdiffusion 1165 -1365 1165 -1365 0 feedthrough
rlabel pdiffusion 1172 -1365 1172 -1365 0 feedthrough
rlabel pdiffusion 1179 -1365 1179 -1365 0 feedthrough
rlabel pdiffusion 1186 -1365 1186 -1365 0 feedthrough
rlabel pdiffusion 1193 -1365 1193 -1365 0 feedthrough
rlabel pdiffusion 1200 -1365 1200 -1365 0 cellNo=256
rlabel pdiffusion 1207 -1365 1207 -1365 0 feedthrough
rlabel pdiffusion 1214 -1365 1214 -1365 0 cellNo=794
rlabel pdiffusion 1221 -1365 1221 -1365 0 feedthrough
rlabel pdiffusion 1228 -1365 1228 -1365 0 feedthrough
rlabel pdiffusion 1235 -1365 1235 -1365 0 feedthrough
rlabel pdiffusion 1242 -1365 1242 -1365 0 feedthrough
rlabel pdiffusion 1249 -1365 1249 -1365 0 feedthrough
rlabel pdiffusion 1256 -1365 1256 -1365 0 feedthrough
rlabel pdiffusion 1263 -1365 1263 -1365 0 feedthrough
rlabel pdiffusion 1270 -1365 1270 -1365 0 feedthrough
rlabel pdiffusion 1277 -1365 1277 -1365 0 feedthrough
rlabel pdiffusion 1284 -1365 1284 -1365 0 feedthrough
rlabel pdiffusion 1291 -1365 1291 -1365 0 feedthrough
rlabel pdiffusion 1298 -1365 1298 -1365 0 feedthrough
rlabel pdiffusion 1305 -1365 1305 -1365 0 feedthrough
rlabel pdiffusion 1312 -1365 1312 -1365 0 feedthrough
rlabel pdiffusion 1319 -1365 1319 -1365 0 feedthrough
rlabel pdiffusion 1326 -1365 1326 -1365 0 feedthrough
rlabel pdiffusion 1333 -1365 1333 -1365 0 feedthrough
rlabel pdiffusion 1340 -1365 1340 -1365 0 feedthrough
rlabel pdiffusion 1347 -1365 1347 -1365 0 feedthrough
rlabel pdiffusion 1354 -1365 1354 -1365 0 feedthrough
rlabel pdiffusion 1361 -1365 1361 -1365 0 feedthrough
rlabel pdiffusion 1368 -1365 1368 -1365 0 feedthrough
rlabel pdiffusion 1375 -1365 1375 -1365 0 feedthrough
rlabel pdiffusion 1382 -1365 1382 -1365 0 feedthrough
rlabel pdiffusion 1389 -1365 1389 -1365 0 feedthrough
rlabel pdiffusion 1396 -1365 1396 -1365 0 feedthrough
rlabel pdiffusion 1403 -1365 1403 -1365 0 feedthrough
rlabel pdiffusion 1410 -1365 1410 -1365 0 feedthrough
rlabel pdiffusion 1417 -1365 1417 -1365 0 feedthrough
rlabel pdiffusion 1424 -1365 1424 -1365 0 feedthrough
rlabel pdiffusion 1431 -1365 1431 -1365 0 feedthrough
rlabel pdiffusion 1438 -1365 1438 -1365 0 feedthrough
rlabel pdiffusion 1445 -1365 1445 -1365 0 feedthrough
rlabel pdiffusion 1452 -1365 1452 -1365 0 feedthrough
rlabel pdiffusion 1459 -1365 1459 -1365 0 feedthrough
rlabel pdiffusion 1466 -1365 1466 -1365 0 feedthrough
rlabel pdiffusion 1473 -1365 1473 -1365 0 feedthrough
rlabel pdiffusion 1480 -1365 1480 -1365 0 feedthrough
rlabel pdiffusion 1487 -1365 1487 -1365 0 feedthrough
rlabel pdiffusion 1494 -1365 1494 -1365 0 feedthrough
rlabel pdiffusion 1501 -1365 1501 -1365 0 feedthrough
rlabel pdiffusion 1508 -1365 1508 -1365 0 feedthrough
rlabel pdiffusion 1515 -1365 1515 -1365 0 feedthrough
rlabel pdiffusion 1522 -1365 1522 -1365 0 feedthrough
rlabel pdiffusion 1529 -1365 1529 -1365 0 feedthrough
rlabel pdiffusion 1536 -1365 1536 -1365 0 feedthrough
rlabel pdiffusion 1543 -1365 1543 -1365 0 feedthrough
rlabel pdiffusion 1550 -1365 1550 -1365 0 feedthrough
rlabel pdiffusion 1557 -1365 1557 -1365 0 feedthrough
rlabel pdiffusion 1564 -1365 1564 -1365 0 feedthrough
rlabel pdiffusion 1571 -1365 1571 -1365 0 feedthrough
rlabel pdiffusion 1578 -1365 1578 -1365 0 feedthrough
rlabel pdiffusion 1585 -1365 1585 -1365 0 feedthrough
rlabel pdiffusion 1592 -1365 1592 -1365 0 feedthrough
rlabel pdiffusion 1599 -1365 1599 -1365 0 feedthrough
rlabel pdiffusion 1606 -1365 1606 -1365 0 feedthrough
rlabel pdiffusion 1613 -1365 1613 -1365 0 feedthrough
rlabel pdiffusion 1620 -1365 1620 -1365 0 feedthrough
rlabel pdiffusion 1627 -1365 1627 -1365 0 feedthrough
rlabel pdiffusion 1634 -1365 1634 -1365 0 feedthrough
rlabel pdiffusion 1641 -1365 1641 -1365 0 feedthrough
rlabel pdiffusion 1648 -1365 1648 -1365 0 feedthrough
rlabel pdiffusion 1655 -1365 1655 -1365 0 feedthrough
rlabel pdiffusion 1662 -1365 1662 -1365 0 feedthrough
rlabel pdiffusion 1669 -1365 1669 -1365 0 feedthrough
rlabel pdiffusion 1676 -1365 1676 -1365 0 feedthrough
rlabel pdiffusion 1683 -1365 1683 -1365 0 feedthrough
rlabel pdiffusion 1690 -1365 1690 -1365 0 feedthrough
rlabel pdiffusion 1697 -1365 1697 -1365 0 feedthrough
rlabel pdiffusion 1704 -1365 1704 -1365 0 feedthrough
rlabel pdiffusion 1711 -1365 1711 -1365 0 feedthrough
rlabel pdiffusion 1718 -1365 1718 -1365 0 feedthrough
rlabel pdiffusion 1725 -1365 1725 -1365 0 feedthrough
rlabel pdiffusion 1732 -1365 1732 -1365 0 feedthrough
rlabel pdiffusion 1739 -1365 1739 -1365 0 feedthrough
rlabel pdiffusion 1746 -1365 1746 -1365 0 feedthrough
rlabel pdiffusion 1753 -1365 1753 -1365 0 feedthrough
rlabel pdiffusion 3 -1506 3 -1506 0 cellNo=1108
rlabel pdiffusion 10 -1506 10 -1506 0 cellNo=1113
rlabel pdiffusion 17 -1506 17 -1506 0 cellNo=1116
rlabel pdiffusion 24 -1506 24 -1506 0 feedthrough
rlabel pdiffusion 31 -1506 31 -1506 0 feedthrough
rlabel pdiffusion 38 -1506 38 -1506 0 feedthrough
rlabel pdiffusion 45 -1506 45 -1506 0 feedthrough
rlabel pdiffusion 52 -1506 52 -1506 0 feedthrough
rlabel pdiffusion 59 -1506 59 -1506 0 feedthrough
rlabel pdiffusion 66 -1506 66 -1506 0 cellNo=305
rlabel pdiffusion 73 -1506 73 -1506 0 feedthrough
rlabel pdiffusion 80 -1506 80 -1506 0 feedthrough
rlabel pdiffusion 87 -1506 87 -1506 0 feedthrough
rlabel pdiffusion 94 -1506 94 -1506 0 feedthrough
rlabel pdiffusion 101 -1506 101 -1506 0 feedthrough
rlabel pdiffusion 108 -1506 108 -1506 0 feedthrough
rlabel pdiffusion 115 -1506 115 -1506 0 feedthrough
rlabel pdiffusion 122 -1506 122 -1506 0 cellNo=13
rlabel pdiffusion 129 -1506 129 -1506 0 cellNo=74
rlabel pdiffusion 136 -1506 136 -1506 0 feedthrough
rlabel pdiffusion 143 -1506 143 -1506 0 feedthrough
rlabel pdiffusion 150 -1506 150 -1506 0 feedthrough
rlabel pdiffusion 157 -1506 157 -1506 0 cellNo=148
rlabel pdiffusion 164 -1506 164 -1506 0 feedthrough
rlabel pdiffusion 171 -1506 171 -1506 0 feedthrough
rlabel pdiffusion 178 -1506 178 -1506 0 feedthrough
rlabel pdiffusion 185 -1506 185 -1506 0 cellNo=230
rlabel pdiffusion 192 -1506 192 -1506 0 cellNo=179
rlabel pdiffusion 199 -1506 199 -1506 0 feedthrough
rlabel pdiffusion 206 -1506 206 -1506 0 feedthrough
rlabel pdiffusion 213 -1506 213 -1506 0 cellNo=549
rlabel pdiffusion 220 -1506 220 -1506 0 feedthrough
rlabel pdiffusion 227 -1506 227 -1506 0 cellNo=536
rlabel pdiffusion 234 -1506 234 -1506 0 feedthrough
rlabel pdiffusion 241 -1506 241 -1506 0 feedthrough
rlabel pdiffusion 248 -1506 248 -1506 0 feedthrough
rlabel pdiffusion 255 -1506 255 -1506 0 cellNo=983
rlabel pdiffusion 262 -1506 262 -1506 0 feedthrough
rlabel pdiffusion 269 -1506 269 -1506 0 feedthrough
rlabel pdiffusion 276 -1506 276 -1506 0 feedthrough
rlabel pdiffusion 283 -1506 283 -1506 0 feedthrough
rlabel pdiffusion 290 -1506 290 -1506 0 feedthrough
rlabel pdiffusion 297 -1506 297 -1506 0 feedthrough
rlabel pdiffusion 304 -1506 304 -1506 0 feedthrough
rlabel pdiffusion 311 -1506 311 -1506 0 feedthrough
rlabel pdiffusion 318 -1506 318 -1506 0 cellNo=501
rlabel pdiffusion 325 -1506 325 -1506 0 feedthrough
rlabel pdiffusion 332 -1506 332 -1506 0 feedthrough
rlabel pdiffusion 339 -1506 339 -1506 0 feedthrough
rlabel pdiffusion 346 -1506 346 -1506 0 feedthrough
rlabel pdiffusion 353 -1506 353 -1506 0 feedthrough
rlabel pdiffusion 360 -1506 360 -1506 0 feedthrough
rlabel pdiffusion 367 -1506 367 -1506 0 feedthrough
rlabel pdiffusion 374 -1506 374 -1506 0 feedthrough
rlabel pdiffusion 381 -1506 381 -1506 0 feedthrough
rlabel pdiffusion 388 -1506 388 -1506 0 feedthrough
rlabel pdiffusion 395 -1506 395 -1506 0 feedthrough
rlabel pdiffusion 402 -1506 402 -1506 0 feedthrough
rlabel pdiffusion 409 -1506 409 -1506 0 feedthrough
rlabel pdiffusion 416 -1506 416 -1506 0 cellNo=932
rlabel pdiffusion 423 -1506 423 -1506 0 feedthrough
rlabel pdiffusion 430 -1506 430 -1506 0 feedthrough
rlabel pdiffusion 437 -1506 437 -1506 0 feedthrough
rlabel pdiffusion 444 -1506 444 -1506 0 feedthrough
rlabel pdiffusion 451 -1506 451 -1506 0 feedthrough
rlabel pdiffusion 458 -1506 458 -1506 0 cellNo=103
rlabel pdiffusion 465 -1506 465 -1506 0 feedthrough
rlabel pdiffusion 472 -1506 472 -1506 0 feedthrough
rlabel pdiffusion 479 -1506 479 -1506 0 cellNo=278
rlabel pdiffusion 486 -1506 486 -1506 0 feedthrough
rlabel pdiffusion 493 -1506 493 -1506 0 feedthrough
rlabel pdiffusion 500 -1506 500 -1506 0 feedthrough
rlabel pdiffusion 507 -1506 507 -1506 0 feedthrough
rlabel pdiffusion 514 -1506 514 -1506 0 cellNo=142
rlabel pdiffusion 521 -1506 521 -1506 0 feedthrough
rlabel pdiffusion 528 -1506 528 -1506 0 feedthrough
rlabel pdiffusion 535 -1506 535 -1506 0 feedthrough
rlabel pdiffusion 542 -1506 542 -1506 0 feedthrough
rlabel pdiffusion 549 -1506 549 -1506 0 feedthrough
rlabel pdiffusion 556 -1506 556 -1506 0 feedthrough
rlabel pdiffusion 563 -1506 563 -1506 0 feedthrough
rlabel pdiffusion 570 -1506 570 -1506 0 feedthrough
rlabel pdiffusion 577 -1506 577 -1506 0 feedthrough
rlabel pdiffusion 584 -1506 584 -1506 0 feedthrough
rlabel pdiffusion 591 -1506 591 -1506 0 feedthrough
rlabel pdiffusion 598 -1506 598 -1506 0 feedthrough
rlabel pdiffusion 605 -1506 605 -1506 0 feedthrough
rlabel pdiffusion 612 -1506 612 -1506 0 feedthrough
rlabel pdiffusion 619 -1506 619 -1506 0 feedthrough
rlabel pdiffusion 626 -1506 626 -1506 0 cellNo=580
rlabel pdiffusion 633 -1506 633 -1506 0 feedthrough
rlabel pdiffusion 640 -1506 640 -1506 0 feedthrough
rlabel pdiffusion 647 -1506 647 -1506 0 feedthrough
rlabel pdiffusion 654 -1506 654 -1506 0 cellNo=30
rlabel pdiffusion 661 -1506 661 -1506 0 feedthrough
rlabel pdiffusion 668 -1506 668 -1506 0 cellNo=108
rlabel pdiffusion 675 -1506 675 -1506 0 feedthrough
rlabel pdiffusion 682 -1506 682 -1506 0 feedthrough
rlabel pdiffusion 689 -1506 689 -1506 0 feedthrough
rlabel pdiffusion 696 -1506 696 -1506 0 feedthrough
rlabel pdiffusion 703 -1506 703 -1506 0 feedthrough
rlabel pdiffusion 710 -1506 710 -1506 0 feedthrough
rlabel pdiffusion 717 -1506 717 -1506 0 cellNo=134
rlabel pdiffusion 724 -1506 724 -1506 0 cellNo=539
rlabel pdiffusion 731 -1506 731 -1506 0 feedthrough
rlabel pdiffusion 738 -1506 738 -1506 0 cellNo=470
rlabel pdiffusion 745 -1506 745 -1506 0 feedthrough
rlabel pdiffusion 752 -1506 752 -1506 0 feedthrough
rlabel pdiffusion 759 -1506 759 -1506 0 cellNo=222
rlabel pdiffusion 766 -1506 766 -1506 0 feedthrough
rlabel pdiffusion 773 -1506 773 -1506 0 feedthrough
rlabel pdiffusion 780 -1506 780 -1506 0 feedthrough
rlabel pdiffusion 787 -1506 787 -1506 0 cellNo=762
rlabel pdiffusion 794 -1506 794 -1506 0 feedthrough
rlabel pdiffusion 801 -1506 801 -1506 0 feedthrough
rlabel pdiffusion 808 -1506 808 -1506 0 feedthrough
rlabel pdiffusion 815 -1506 815 -1506 0 feedthrough
rlabel pdiffusion 822 -1506 822 -1506 0 cellNo=375
rlabel pdiffusion 829 -1506 829 -1506 0 cellNo=716
rlabel pdiffusion 836 -1506 836 -1506 0 feedthrough
rlabel pdiffusion 843 -1506 843 -1506 0 feedthrough
rlabel pdiffusion 850 -1506 850 -1506 0 feedthrough
rlabel pdiffusion 857 -1506 857 -1506 0 feedthrough
rlabel pdiffusion 864 -1506 864 -1506 0 cellNo=887
rlabel pdiffusion 871 -1506 871 -1506 0 feedthrough
rlabel pdiffusion 878 -1506 878 -1506 0 feedthrough
rlabel pdiffusion 885 -1506 885 -1506 0 feedthrough
rlabel pdiffusion 892 -1506 892 -1506 0 feedthrough
rlabel pdiffusion 899 -1506 899 -1506 0 feedthrough
rlabel pdiffusion 906 -1506 906 -1506 0 feedthrough
rlabel pdiffusion 913 -1506 913 -1506 0 feedthrough
rlabel pdiffusion 920 -1506 920 -1506 0 feedthrough
rlabel pdiffusion 927 -1506 927 -1506 0 feedthrough
rlabel pdiffusion 934 -1506 934 -1506 0 cellNo=356
rlabel pdiffusion 941 -1506 941 -1506 0 feedthrough
rlabel pdiffusion 948 -1506 948 -1506 0 cellNo=913
rlabel pdiffusion 955 -1506 955 -1506 0 feedthrough
rlabel pdiffusion 962 -1506 962 -1506 0 feedthrough
rlabel pdiffusion 969 -1506 969 -1506 0 feedthrough
rlabel pdiffusion 976 -1506 976 -1506 0 cellNo=659
rlabel pdiffusion 983 -1506 983 -1506 0 feedthrough
rlabel pdiffusion 990 -1506 990 -1506 0 feedthrough
rlabel pdiffusion 997 -1506 997 -1506 0 feedthrough
rlabel pdiffusion 1004 -1506 1004 -1506 0 feedthrough
rlabel pdiffusion 1011 -1506 1011 -1506 0 feedthrough
rlabel pdiffusion 1018 -1506 1018 -1506 0 feedthrough
rlabel pdiffusion 1025 -1506 1025 -1506 0 feedthrough
rlabel pdiffusion 1032 -1506 1032 -1506 0 cellNo=610
rlabel pdiffusion 1039 -1506 1039 -1506 0 feedthrough
rlabel pdiffusion 1046 -1506 1046 -1506 0 cellNo=300
rlabel pdiffusion 1053 -1506 1053 -1506 0 feedthrough
rlabel pdiffusion 1060 -1506 1060 -1506 0 feedthrough
rlabel pdiffusion 1067 -1506 1067 -1506 0 feedthrough
rlabel pdiffusion 1074 -1506 1074 -1506 0 feedthrough
rlabel pdiffusion 1081 -1506 1081 -1506 0 feedthrough
rlabel pdiffusion 1088 -1506 1088 -1506 0 feedthrough
rlabel pdiffusion 1095 -1506 1095 -1506 0 feedthrough
rlabel pdiffusion 1102 -1506 1102 -1506 0 feedthrough
rlabel pdiffusion 1109 -1506 1109 -1506 0 feedthrough
rlabel pdiffusion 1116 -1506 1116 -1506 0 feedthrough
rlabel pdiffusion 1123 -1506 1123 -1506 0 feedthrough
rlabel pdiffusion 1130 -1506 1130 -1506 0 feedthrough
rlabel pdiffusion 1137 -1506 1137 -1506 0 feedthrough
rlabel pdiffusion 1144 -1506 1144 -1506 0 feedthrough
rlabel pdiffusion 1151 -1506 1151 -1506 0 feedthrough
rlabel pdiffusion 1158 -1506 1158 -1506 0 feedthrough
rlabel pdiffusion 1165 -1506 1165 -1506 0 feedthrough
rlabel pdiffusion 1172 -1506 1172 -1506 0 feedthrough
rlabel pdiffusion 1179 -1506 1179 -1506 0 feedthrough
rlabel pdiffusion 1186 -1506 1186 -1506 0 feedthrough
rlabel pdiffusion 1193 -1506 1193 -1506 0 feedthrough
rlabel pdiffusion 1200 -1506 1200 -1506 0 feedthrough
rlabel pdiffusion 1207 -1506 1207 -1506 0 feedthrough
rlabel pdiffusion 1214 -1506 1214 -1506 0 feedthrough
rlabel pdiffusion 1221 -1506 1221 -1506 0 feedthrough
rlabel pdiffusion 1228 -1506 1228 -1506 0 feedthrough
rlabel pdiffusion 1235 -1506 1235 -1506 0 feedthrough
rlabel pdiffusion 1242 -1506 1242 -1506 0 feedthrough
rlabel pdiffusion 1249 -1506 1249 -1506 0 feedthrough
rlabel pdiffusion 1256 -1506 1256 -1506 0 feedthrough
rlabel pdiffusion 1263 -1506 1263 -1506 0 feedthrough
rlabel pdiffusion 1270 -1506 1270 -1506 0 feedthrough
rlabel pdiffusion 1277 -1506 1277 -1506 0 feedthrough
rlabel pdiffusion 1284 -1506 1284 -1506 0 feedthrough
rlabel pdiffusion 1291 -1506 1291 -1506 0 feedthrough
rlabel pdiffusion 1298 -1506 1298 -1506 0 feedthrough
rlabel pdiffusion 1305 -1506 1305 -1506 0 feedthrough
rlabel pdiffusion 1312 -1506 1312 -1506 0 feedthrough
rlabel pdiffusion 1319 -1506 1319 -1506 0 feedthrough
rlabel pdiffusion 1326 -1506 1326 -1506 0 feedthrough
rlabel pdiffusion 1333 -1506 1333 -1506 0 feedthrough
rlabel pdiffusion 1340 -1506 1340 -1506 0 feedthrough
rlabel pdiffusion 1347 -1506 1347 -1506 0 feedthrough
rlabel pdiffusion 1354 -1506 1354 -1506 0 feedthrough
rlabel pdiffusion 1361 -1506 1361 -1506 0 feedthrough
rlabel pdiffusion 1368 -1506 1368 -1506 0 feedthrough
rlabel pdiffusion 1375 -1506 1375 -1506 0 feedthrough
rlabel pdiffusion 1382 -1506 1382 -1506 0 feedthrough
rlabel pdiffusion 1389 -1506 1389 -1506 0 feedthrough
rlabel pdiffusion 1396 -1506 1396 -1506 0 feedthrough
rlabel pdiffusion 1403 -1506 1403 -1506 0 feedthrough
rlabel pdiffusion 1410 -1506 1410 -1506 0 feedthrough
rlabel pdiffusion 1417 -1506 1417 -1506 0 feedthrough
rlabel pdiffusion 1424 -1506 1424 -1506 0 feedthrough
rlabel pdiffusion 1431 -1506 1431 -1506 0 feedthrough
rlabel pdiffusion 1438 -1506 1438 -1506 0 feedthrough
rlabel pdiffusion 1445 -1506 1445 -1506 0 feedthrough
rlabel pdiffusion 1452 -1506 1452 -1506 0 feedthrough
rlabel pdiffusion 1459 -1506 1459 -1506 0 feedthrough
rlabel pdiffusion 1466 -1506 1466 -1506 0 feedthrough
rlabel pdiffusion 1473 -1506 1473 -1506 0 feedthrough
rlabel pdiffusion 1480 -1506 1480 -1506 0 feedthrough
rlabel pdiffusion 1487 -1506 1487 -1506 0 feedthrough
rlabel pdiffusion 1494 -1506 1494 -1506 0 feedthrough
rlabel pdiffusion 1501 -1506 1501 -1506 0 feedthrough
rlabel pdiffusion 1508 -1506 1508 -1506 0 feedthrough
rlabel pdiffusion 1515 -1506 1515 -1506 0 feedthrough
rlabel pdiffusion 1522 -1506 1522 -1506 0 feedthrough
rlabel pdiffusion 1529 -1506 1529 -1506 0 feedthrough
rlabel pdiffusion 1536 -1506 1536 -1506 0 cellNo=254
rlabel pdiffusion 1543 -1506 1543 -1506 0 feedthrough
rlabel pdiffusion 1550 -1506 1550 -1506 0 cellNo=859
rlabel pdiffusion 1557 -1506 1557 -1506 0 feedthrough
rlabel pdiffusion 1564 -1506 1564 -1506 0 feedthrough
rlabel pdiffusion 1571 -1506 1571 -1506 0 feedthrough
rlabel pdiffusion 1578 -1506 1578 -1506 0 feedthrough
rlabel pdiffusion 1585 -1506 1585 -1506 0 cellNo=43
rlabel pdiffusion 1592 -1506 1592 -1506 0 feedthrough
rlabel pdiffusion 1599 -1506 1599 -1506 0 feedthrough
rlabel pdiffusion 1606 -1506 1606 -1506 0 cellNo=559
rlabel pdiffusion 1613 -1506 1613 -1506 0 feedthrough
rlabel pdiffusion 1620 -1506 1620 -1506 0 feedthrough
rlabel pdiffusion 1627 -1506 1627 -1506 0 feedthrough
rlabel pdiffusion 1634 -1506 1634 -1506 0 feedthrough
rlabel pdiffusion 1641 -1506 1641 -1506 0 cellNo=685
rlabel pdiffusion 1648 -1506 1648 -1506 0 feedthrough
rlabel pdiffusion 1655 -1506 1655 -1506 0 feedthrough
rlabel pdiffusion 1662 -1506 1662 -1506 0 feedthrough
rlabel pdiffusion 1669 -1506 1669 -1506 0 feedthrough
rlabel pdiffusion 1676 -1506 1676 -1506 0 feedthrough
rlabel pdiffusion 1683 -1506 1683 -1506 0 feedthrough
rlabel pdiffusion 1690 -1506 1690 -1506 0 feedthrough
rlabel pdiffusion 1697 -1506 1697 -1506 0 feedthrough
rlabel pdiffusion 1704 -1506 1704 -1506 0 feedthrough
rlabel pdiffusion 1711 -1506 1711 -1506 0 feedthrough
rlabel pdiffusion 1718 -1506 1718 -1506 0 feedthrough
rlabel pdiffusion 1725 -1506 1725 -1506 0 feedthrough
rlabel pdiffusion 1732 -1506 1732 -1506 0 feedthrough
rlabel pdiffusion 1802 -1506 1802 -1506 0 feedthrough
rlabel pdiffusion 3 -1641 3 -1641 0 cellNo=1112
rlabel pdiffusion 10 -1641 10 -1641 0 cellNo=1115
rlabel pdiffusion 17 -1641 17 -1641 0 cellNo=1119
rlabel pdiffusion 24 -1641 24 -1641 0 feedthrough
rlabel pdiffusion 31 -1641 31 -1641 0 feedthrough
rlabel pdiffusion 38 -1641 38 -1641 0 feedthrough
rlabel pdiffusion 45 -1641 45 -1641 0 feedthrough
rlabel pdiffusion 52 -1641 52 -1641 0 feedthrough
rlabel pdiffusion 59 -1641 59 -1641 0 cellNo=486
rlabel pdiffusion 66 -1641 66 -1641 0 feedthrough
rlabel pdiffusion 73 -1641 73 -1641 0 feedthrough
rlabel pdiffusion 80 -1641 80 -1641 0 feedthrough
rlabel pdiffusion 87 -1641 87 -1641 0 feedthrough
rlabel pdiffusion 94 -1641 94 -1641 0 feedthrough
rlabel pdiffusion 101 -1641 101 -1641 0 feedthrough
rlabel pdiffusion 108 -1641 108 -1641 0 feedthrough
rlabel pdiffusion 115 -1641 115 -1641 0 feedthrough
rlabel pdiffusion 122 -1641 122 -1641 0 cellNo=595
rlabel pdiffusion 129 -1641 129 -1641 0 feedthrough
rlabel pdiffusion 136 -1641 136 -1641 0 feedthrough
rlabel pdiffusion 143 -1641 143 -1641 0 feedthrough
rlabel pdiffusion 150 -1641 150 -1641 0 feedthrough
rlabel pdiffusion 157 -1641 157 -1641 0 feedthrough
rlabel pdiffusion 164 -1641 164 -1641 0 cellNo=268
rlabel pdiffusion 171 -1641 171 -1641 0 feedthrough
rlabel pdiffusion 178 -1641 178 -1641 0 feedthrough
rlabel pdiffusion 185 -1641 185 -1641 0 cellNo=899
rlabel pdiffusion 192 -1641 192 -1641 0 feedthrough
rlabel pdiffusion 199 -1641 199 -1641 0 feedthrough
rlabel pdiffusion 206 -1641 206 -1641 0 feedthrough
rlabel pdiffusion 213 -1641 213 -1641 0 feedthrough
rlabel pdiffusion 220 -1641 220 -1641 0 cellNo=453
rlabel pdiffusion 227 -1641 227 -1641 0 feedthrough
rlabel pdiffusion 234 -1641 234 -1641 0 feedthrough
rlabel pdiffusion 241 -1641 241 -1641 0 feedthrough
rlabel pdiffusion 248 -1641 248 -1641 0 feedthrough
rlabel pdiffusion 255 -1641 255 -1641 0 feedthrough
rlabel pdiffusion 262 -1641 262 -1641 0 cellNo=713
rlabel pdiffusion 269 -1641 269 -1641 0 feedthrough
rlabel pdiffusion 276 -1641 276 -1641 0 feedthrough
rlabel pdiffusion 283 -1641 283 -1641 0 feedthrough
rlabel pdiffusion 290 -1641 290 -1641 0 feedthrough
rlabel pdiffusion 297 -1641 297 -1641 0 feedthrough
rlabel pdiffusion 304 -1641 304 -1641 0 feedthrough
rlabel pdiffusion 311 -1641 311 -1641 0 cellNo=462
rlabel pdiffusion 318 -1641 318 -1641 0 feedthrough
rlabel pdiffusion 325 -1641 325 -1641 0 feedthrough
rlabel pdiffusion 332 -1641 332 -1641 0 feedthrough
rlabel pdiffusion 339 -1641 339 -1641 0 feedthrough
rlabel pdiffusion 346 -1641 346 -1641 0 feedthrough
rlabel pdiffusion 353 -1641 353 -1641 0 feedthrough
rlabel pdiffusion 360 -1641 360 -1641 0 feedthrough
rlabel pdiffusion 367 -1641 367 -1641 0 feedthrough
rlabel pdiffusion 374 -1641 374 -1641 0 feedthrough
rlabel pdiffusion 381 -1641 381 -1641 0 feedthrough
rlabel pdiffusion 388 -1641 388 -1641 0 feedthrough
rlabel pdiffusion 395 -1641 395 -1641 0 feedthrough
rlabel pdiffusion 402 -1641 402 -1641 0 feedthrough
rlabel pdiffusion 409 -1641 409 -1641 0 feedthrough
rlabel pdiffusion 416 -1641 416 -1641 0 feedthrough
rlabel pdiffusion 423 -1641 423 -1641 0 feedthrough
rlabel pdiffusion 430 -1641 430 -1641 0 feedthrough
rlabel pdiffusion 437 -1641 437 -1641 0 feedthrough
rlabel pdiffusion 444 -1641 444 -1641 0 cellNo=445
rlabel pdiffusion 451 -1641 451 -1641 0 cellNo=370
rlabel pdiffusion 458 -1641 458 -1641 0 feedthrough
rlabel pdiffusion 465 -1641 465 -1641 0 feedthrough
rlabel pdiffusion 472 -1641 472 -1641 0 feedthrough
rlabel pdiffusion 479 -1641 479 -1641 0 feedthrough
rlabel pdiffusion 486 -1641 486 -1641 0 feedthrough
rlabel pdiffusion 493 -1641 493 -1641 0 feedthrough
rlabel pdiffusion 500 -1641 500 -1641 0 feedthrough
rlabel pdiffusion 507 -1641 507 -1641 0 feedthrough
rlabel pdiffusion 514 -1641 514 -1641 0 feedthrough
rlabel pdiffusion 521 -1641 521 -1641 0 feedthrough
rlabel pdiffusion 528 -1641 528 -1641 0 feedthrough
rlabel pdiffusion 535 -1641 535 -1641 0 feedthrough
rlabel pdiffusion 542 -1641 542 -1641 0 cellNo=898
rlabel pdiffusion 549 -1641 549 -1641 0 cellNo=426
rlabel pdiffusion 556 -1641 556 -1641 0 feedthrough
rlabel pdiffusion 563 -1641 563 -1641 0 feedthrough
rlabel pdiffusion 570 -1641 570 -1641 0 feedthrough
rlabel pdiffusion 577 -1641 577 -1641 0 feedthrough
rlabel pdiffusion 584 -1641 584 -1641 0 feedthrough
rlabel pdiffusion 591 -1641 591 -1641 0 feedthrough
rlabel pdiffusion 598 -1641 598 -1641 0 feedthrough
rlabel pdiffusion 605 -1641 605 -1641 0 cellNo=319
rlabel pdiffusion 612 -1641 612 -1641 0 feedthrough
rlabel pdiffusion 619 -1641 619 -1641 0 feedthrough
rlabel pdiffusion 626 -1641 626 -1641 0 feedthrough
rlabel pdiffusion 633 -1641 633 -1641 0 feedthrough
rlabel pdiffusion 640 -1641 640 -1641 0 feedthrough
rlabel pdiffusion 647 -1641 647 -1641 0 feedthrough
rlabel pdiffusion 654 -1641 654 -1641 0 feedthrough
rlabel pdiffusion 661 -1641 661 -1641 0 feedthrough
rlabel pdiffusion 668 -1641 668 -1641 0 feedthrough
rlabel pdiffusion 675 -1641 675 -1641 0 feedthrough
rlabel pdiffusion 682 -1641 682 -1641 0 feedthrough
rlabel pdiffusion 689 -1641 689 -1641 0 feedthrough
rlabel pdiffusion 696 -1641 696 -1641 0 feedthrough
rlabel pdiffusion 703 -1641 703 -1641 0 feedthrough
rlabel pdiffusion 710 -1641 710 -1641 0 feedthrough
rlabel pdiffusion 717 -1641 717 -1641 0 feedthrough
rlabel pdiffusion 724 -1641 724 -1641 0 cellNo=50
rlabel pdiffusion 731 -1641 731 -1641 0 cellNo=37
rlabel pdiffusion 738 -1641 738 -1641 0 feedthrough
rlabel pdiffusion 745 -1641 745 -1641 0 cellNo=680
rlabel pdiffusion 752 -1641 752 -1641 0 cellNo=195
rlabel pdiffusion 759 -1641 759 -1641 0 feedthrough
rlabel pdiffusion 766 -1641 766 -1641 0 feedthrough
rlabel pdiffusion 773 -1641 773 -1641 0 feedthrough
rlabel pdiffusion 780 -1641 780 -1641 0 feedthrough
rlabel pdiffusion 787 -1641 787 -1641 0 feedthrough
rlabel pdiffusion 794 -1641 794 -1641 0 feedthrough
rlabel pdiffusion 801 -1641 801 -1641 0 feedthrough
rlabel pdiffusion 808 -1641 808 -1641 0 feedthrough
rlabel pdiffusion 815 -1641 815 -1641 0 cellNo=89
rlabel pdiffusion 822 -1641 822 -1641 0 cellNo=318
rlabel pdiffusion 829 -1641 829 -1641 0 feedthrough
rlabel pdiffusion 836 -1641 836 -1641 0 feedthrough
rlabel pdiffusion 843 -1641 843 -1641 0 feedthrough
rlabel pdiffusion 850 -1641 850 -1641 0 feedthrough
rlabel pdiffusion 857 -1641 857 -1641 0 cellNo=862
rlabel pdiffusion 864 -1641 864 -1641 0 cellNo=869
rlabel pdiffusion 871 -1641 871 -1641 0 feedthrough
rlabel pdiffusion 878 -1641 878 -1641 0 cellNo=970
rlabel pdiffusion 885 -1641 885 -1641 0 feedthrough
rlabel pdiffusion 892 -1641 892 -1641 0 cellNo=964
rlabel pdiffusion 899 -1641 899 -1641 0 feedthrough
rlabel pdiffusion 906 -1641 906 -1641 0 feedthrough
rlabel pdiffusion 913 -1641 913 -1641 0 feedthrough
rlabel pdiffusion 920 -1641 920 -1641 0 feedthrough
rlabel pdiffusion 927 -1641 927 -1641 0 feedthrough
rlabel pdiffusion 934 -1641 934 -1641 0 feedthrough
rlabel pdiffusion 941 -1641 941 -1641 0 feedthrough
rlabel pdiffusion 948 -1641 948 -1641 0 feedthrough
rlabel pdiffusion 955 -1641 955 -1641 0 cellNo=244
rlabel pdiffusion 962 -1641 962 -1641 0 feedthrough
rlabel pdiffusion 969 -1641 969 -1641 0 feedthrough
rlabel pdiffusion 976 -1641 976 -1641 0 feedthrough
rlabel pdiffusion 983 -1641 983 -1641 0 feedthrough
rlabel pdiffusion 990 -1641 990 -1641 0 feedthrough
rlabel pdiffusion 997 -1641 997 -1641 0 feedthrough
rlabel pdiffusion 1004 -1641 1004 -1641 0 cellNo=437
rlabel pdiffusion 1011 -1641 1011 -1641 0 feedthrough
rlabel pdiffusion 1018 -1641 1018 -1641 0 cellNo=963
rlabel pdiffusion 1025 -1641 1025 -1641 0 feedthrough
rlabel pdiffusion 1032 -1641 1032 -1641 0 feedthrough
rlabel pdiffusion 1039 -1641 1039 -1641 0 feedthrough
rlabel pdiffusion 1046 -1641 1046 -1641 0 feedthrough
rlabel pdiffusion 1053 -1641 1053 -1641 0 feedthrough
rlabel pdiffusion 1060 -1641 1060 -1641 0 cellNo=567
rlabel pdiffusion 1067 -1641 1067 -1641 0 feedthrough
rlabel pdiffusion 1074 -1641 1074 -1641 0 feedthrough
rlabel pdiffusion 1081 -1641 1081 -1641 0 cellNo=57
rlabel pdiffusion 1088 -1641 1088 -1641 0 feedthrough
rlabel pdiffusion 1095 -1641 1095 -1641 0 feedthrough
rlabel pdiffusion 1102 -1641 1102 -1641 0 feedthrough
rlabel pdiffusion 1109 -1641 1109 -1641 0 cellNo=535
rlabel pdiffusion 1116 -1641 1116 -1641 0 feedthrough
rlabel pdiffusion 1123 -1641 1123 -1641 0 cellNo=592
rlabel pdiffusion 1130 -1641 1130 -1641 0 feedthrough
rlabel pdiffusion 1137 -1641 1137 -1641 0 feedthrough
rlabel pdiffusion 1144 -1641 1144 -1641 0 feedthrough
rlabel pdiffusion 1151 -1641 1151 -1641 0 feedthrough
rlabel pdiffusion 1158 -1641 1158 -1641 0 feedthrough
rlabel pdiffusion 1165 -1641 1165 -1641 0 feedthrough
rlabel pdiffusion 1172 -1641 1172 -1641 0 feedthrough
rlabel pdiffusion 1179 -1641 1179 -1641 0 feedthrough
rlabel pdiffusion 1186 -1641 1186 -1641 0 cellNo=829
rlabel pdiffusion 1193 -1641 1193 -1641 0 feedthrough
rlabel pdiffusion 1200 -1641 1200 -1641 0 feedthrough
rlabel pdiffusion 1207 -1641 1207 -1641 0 cellNo=414
rlabel pdiffusion 1214 -1641 1214 -1641 0 feedthrough
rlabel pdiffusion 1221 -1641 1221 -1641 0 feedthrough
rlabel pdiffusion 1228 -1641 1228 -1641 0 feedthrough
rlabel pdiffusion 1235 -1641 1235 -1641 0 feedthrough
rlabel pdiffusion 1242 -1641 1242 -1641 0 feedthrough
rlabel pdiffusion 1249 -1641 1249 -1641 0 feedthrough
rlabel pdiffusion 1256 -1641 1256 -1641 0 feedthrough
rlabel pdiffusion 1263 -1641 1263 -1641 0 feedthrough
rlabel pdiffusion 1270 -1641 1270 -1641 0 feedthrough
rlabel pdiffusion 1277 -1641 1277 -1641 0 feedthrough
rlabel pdiffusion 1284 -1641 1284 -1641 0 feedthrough
rlabel pdiffusion 1291 -1641 1291 -1641 0 feedthrough
rlabel pdiffusion 1298 -1641 1298 -1641 0 cellNo=427
rlabel pdiffusion 1305 -1641 1305 -1641 0 feedthrough
rlabel pdiffusion 1312 -1641 1312 -1641 0 feedthrough
rlabel pdiffusion 1319 -1641 1319 -1641 0 feedthrough
rlabel pdiffusion 1326 -1641 1326 -1641 0 feedthrough
rlabel pdiffusion 1333 -1641 1333 -1641 0 feedthrough
rlabel pdiffusion 1340 -1641 1340 -1641 0 feedthrough
rlabel pdiffusion 1347 -1641 1347 -1641 0 feedthrough
rlabel pdiffusion 1354 -1641 1354 -1641 0 feedthrough
rlabel pdiffusion 1361 -1641 1361 -1641 0 feedthrough
rlabel pdiffusion 1368 -1641 1368 -1641 0 feedthrough
rlabel pdiffusion 1375 -1641 1375 -1641 0 feedthrough
rlabel pdiffusion 1382 -1641 1382 -1641 0 feedthrough
rlabel pdiffusion 1389 -1641 1389 -1641 0 feedthrough
rlabel pdiffusion 1396 -1641 1396 -1641 0 feedthrough
rlabel pdiffusion 1403 -1641 1403 -1641 0 feedthrough
rlabel pdiffusion 1410 -1641 1410 -1641 0 feedthrough
rlabel pdiffusion 1417 -1641 1417 -1641 0 feedthrough
rlabel pdiffusion 1424 -1641 1424 -1641 0 feedthrough
rlabel pdiffusion 1431 -1641 1431 -1641 0 feedthrough
rlabel pdiffusion 1438 -1641 1438 -1641 0 feedthrough
rlabel pdiffusion 1445 -1641 1445 -1641 0 feedthrough
rlabel pdiffusion 1452 -1641 1452 -1641 0 feedthrough
rlabel pdiffusion 1459 -1641 1459 -1641 0 feedthrough
rlabel pdiffusion 1466 -1641 1466 -1641 0 feedthrough
rlabel pdiffusion 1473 -1641 1473 -1641 0 feedthrough
rlabel pdiffusion 1480 -1641 1480 -1641 0 feedthrough
rlabel pdiffusion 1487 -1641 1487 -1641 0 feedthrough
rlabel pdiffusion 1494 -1641 1494 -1641 0 feedthrough
rlabel pdiffusion 1501 -1641 1501 -1641 0 feedthrough
rlabel pdiffusion 1508 -1641 1508 -1641 0 feedthrough
rlabel pdiffusion 1515 -1641 1515 -1641 0 feedthrough
rlabel pdiffusion 1522 -1641 1522 -1641 0 feedthrough
rlabel pdiffusion 1529 -1641 1529 -1641 0 feedthrough
rlabel pdiffusion 1536 -1641 1536 -1641 0 feedthrough
rlabel pdiffusion 1543 -1641 1543 -1641 0 feedthrough
rlabel pdiffusion 1550 -1641 1550 -1641 0 feedthrough
rlabel pdiffusion 1557 -1641 1557 -1641 0 feedthrough
rlabel pdiffusion 1564 -1641 1564 -1641 0 feedthrough
rlabel pdiffusion 1571 -1641 1571 -1641 0 feedthrough
rlabel pdiffusion 1578 -1641 1578 -1641 0 feedthrough
rlabel pdiffusion 1585 -1641 1585 -1641 0 feedthrough
rlabel pdiffusion 1592 -1641 1592 -1641 0 feedthrough
rlabel pdiffusion 1599 -1641 1599 -1641 0 feedthrough
rlabel pdiffusion 1606 -1641 1606 -1641 0 feedthrough
rlabel pdiffusion 1613 -1641 1613 -1641 0 feedthrough
rlabel pdiffusion 1620 -1641 1620 -1641 0 feedthrough
rlabel pdiffusion 1627 -1641 1627 -1641 0 feedthrough
rlabel pdiffusion 1634 -1641 1634 -1641 0 feedthrough
rlabel pdiffusion 1641 -1641 1641 -1641 0 feedthrough
rlabel pdiffusion 1648 -1641 1648 -1641 0 cellNo=60
rlabel pdiffusion 1655 -1641 1655 -1641 0 feedthrough
rlabel pdiffusion 1662 -1641 1662 -1641 0 feedthrough
rlabel pdiffusion 1669 -1641 1669 -1641 0 feedthrough
rlabel pdiffusion 1676 -1641 1676 -1641 0 feedthrough
rlabel pdiffusion 1683 -1641 1683 -1641 0 cellNo=172
rlabel pdiffusion 1690 -1641 1690 -1641 0 feedthrough
rlabel pdiffusion 1697 -1641 1697 -1641 0 feedthrough
rlabel pdiffusion 1704 -1641 1704 -1641 0 cellNo=769
rlabel pdiffusion 1711 -1641 1711 -1641 0 feedthrough
rlabel pdiffusion 1718 -1641 1718 -1641 0 feedthrough
rlabel pdiffusion 1725 -1641 1725 -1641 0 feedthrough
rlabel pdiffusion 1823 -1641 1823 -1641 0 feedthrough
rlabel pdiffusion 3 -1788 3 -1788 0 cellNo=1114
rlabel pdiffusion 10 -1788 10 -1788 0 cellNo=1118
rlabel pdiffusion 17 -1788 17 -1788 0 cellNo=1122
rlabel pdiffusion 24 -1788 24 -1788 0 feedthrough
rlabel pdiffusion 31 -1788 31 -1788 0 feedthrough
rlabel pdiffusion 38 -1788 38 -1788 0 feedthrough
rlabel pdiffusion 45 -1788 45 -1788 0 feedthrough
rlabel pdiffusion 52 -1788 52 -1788 0 feedthrough
rlabel pdiffusion 59 -1788 59 -1788 0 feedthrough
rlabel pdiffusion 66 -1788 66 -1788 0 feedthrough
rlabel pdiffusion 73 -1788 73 -1788 0 cellNo=270
rlabel pdiffusion 80 -1788 80 -1788 0 feedthrough
rlabel pdiffusion 87 -1788 87 -1788 0 cellNo=839
rlabel pdiffusion 94 -1788 94 -1788 0 feedthrough
rlabel pdiffusion 101 -1788 101 -1788 0 feedthrough
rlabel pdiffusion 108 -1788 108 -1788 0 feedthrough
rlabel pdiffusion 115 -1788 115 -1788 0 cellNo=102
rlabel pdiffusion 122 -1788 122 -1788 0 feedthrough
rlabel pdiffusion 129 -1788 129 -1788 0 feedthrough
rlabel pdiffusion 136 -1788 136 -1788 0 feedthrough
rlabel pdiffusion 143 -1788 143 -1788 0 cellNo=24
rlabel pdiffusion 150 -1788 150 -1788 0 feedthrough
rlabel pdiffusion 157 -1788 157 -1788 0 cellNo=749
rlabel pdiffusion 164 -1788 164 -1788 0 feedthrough
rlabel pdiffusion 171 -1788 171 -1788 0 feedthrough
rlabel pdiffusion 178 -1788 178 -1788 0 feedthrough
rlabel pdiffusion 185 -1788 185 -1788 0 feedthrough
rlabel pdiffusion 192 -1788 192 -1788 0 feedthrough
rlabel pdiffusion 199 -1788 199 -1788 0 feedthrough
rlabel pdiffusion 206 -1788 206 -1788 0 feedthrough
rlabel pdiffusion 213 -1788 213 -1788 0 feedthrough
rlabel pdiffusion 220 -1788 220 -1788 0 cellNo=776
rlabel pdiffusion 227 -1788 227 -1788 0 feedthrough
rlabel pdiffusion 234 -1788 234 -1788 0 cellNo=788
rlabel pdiffusion 241 -1788 241 -1788 0 feedthrough
rlabel pdiffusion 248 -1788 248 -1788 0 feedthrough
rlabel pdiffusion 255 -1788 255 -1788 0 feedthrough
rlabel pdiffusion 262 -1788 262 -1788 0 cellNo=620
rlabel pdiffusion 269 -1788 269 -1788 0 feedthrough
rlabel pdiffusion 276 -1788 276 -1788 0 feedthrough
rlabel pdiffusion 283 -1788 283 -1788 0 feedthrough
rlabel pdiffusion 290 -1788 290 -1788 0 feedthrough
rlabel pdiffusion 297 -1788 297 -1788 0 feedthrough
rlabel pdiffusion 304 -1788 304 -1788 0 feedthrough
rlabel pdiffusion 311 -1788 311 -1788 0 feedthrough
rlabel pdiffusion 318 -1788 318 -1788 0 feedthrough
rlabel pdiffusion 325 -1788 325 -1788 0 feedthrough
rlabel pdiffusion 332 -1788 332 -1788 0 feedthrough
rlabel pdiffusion 339 -1788 339 -1788 0 feedthrough
rlabel pdiffusion 346 -1788 346 -1788 0 feedthrough
rlabel pdiffusion 353 -1788 353 -1788 0 feedthrough
rlabel pdiffusion 360 -1788 360 -1788 0 cellNo=99
rlabel pdiffusion 367 -1788 367 -1788 0 feedthrough
rlabel pdiffusion 374 -1788 374 -1788 0 feedthrough
rlabel pdiffusion 381 -1788 381 -1788 0 cellNo=555
rlabel pdiffusion 388 -1788 388 -1788 0 feedthrough
rlabel pdiffusion 395 -1788 395 -1788 0 feedthrough
rlabel pdiffusion 402 -1788 402 -1788 0 feedthrough
rlabel pdiffusion 409 -1788 409 -1788 0 feedthrough
rlabel pdiffusion 416 -1788 416 -1788 0 feedthrough
rlabel pdiffusion 423 -1788 423 -1788 0 feedthrough
rlabel pdiffusion 430 -1788 430 -1788 0 feedthrough
rlabel pdiffusion 437 -1788 437 -1788 0 feedthrough
rlabel pdiffusion 444 -1788 444 -1788 0 feedthrough
rlabel pdiffusion 451 -1788 451 -1788 0 feedthrough
rlabel pdiffusion 458 -1788 458 -1788 0 feedthrough
rlabel pdiffusion 465 -1788 465 -1788 0 feedthrough
rlabel pdiffusion 472 -1788 472 -1788 0 feedthrough
rlabel pdiffusion 479 -1788 479 -1788 0 feedthrough
rlabel pdiffusion 486 -1788 486 -1788 0 feedthrough
rlabel pdiffusion 493 -1788 493 -1788 0 feedthrough
rlabel pdiffusion 500 -1788 500 -1788 0 cellNo=993
rlabel pdiffusion 507 -1788 507 -1788 0 feedthrough
rlabel pdiffusion 514 -1788 514 -1788 0 feedthrough
rlabel pdiffusion 521 -1788 521 -1788 0 feedthrough
rlabel pdiffusion 528 -1788 528 -1788 0 feedthrough
rlabel pdiffusion 535 -1788 535 -1788 0 cellNo=385
rlabel pdiffusion 542 -1788 542 -1788 0 cellNo=18
rlabel pdiffusion 549 -1788 549 -1788 0 cellNo=987
rlabel pdiffusion 556 -1788 556 -1788 0 feedthrough
rlabel pdiffusion 563 -1788 563 -1788 0 feedthrough
rlabel pdiffusion 570 -1788 570 -1788 0 feedthrough
rlabel pdiffusion 577 -1788 577 -1788 0 cellNo=673
rlabel pdiffusion 584 -1788 584 -1788 0 cellNo=7
rlabel pdiffusion 591 -1788 591 -1788 0 cellNo=376
rlabel pdiffusion 598 -1788 598 -1788 0 feedthrough
rlabel pdiffusion 605 -1788 605 -1788 0 feedthrough
rlabel pdiffusion 612 -1788 612 -1788 0 feedthrough
rlabel pdiffusion 619 -1788 619 -1788 0 feedthrough
rlabel pdiffusion 626 -1788 626 -1788 0 feedthrough
rlabel pdiffusion 633 -1788 633 -1788 0 cellNo=358
rlabel pdiffusion 640 -1788 640 -1788 0 feedthrough
rlabel pdiffusion 647 -1788 647 -1788 0 feedthrough
rlabel pdiffusion 654 -1788 654 -1788 0 feedthrough
rlabel pdiffusion 661 -1788 661 -1788 0 feedthrough
rlabel pdiffusion 668 -1788 668 -1788 0 feedthrough
rlabel pdiffusion 675 -1788 675 -1788 0 cellNo=96
rlabel pdiffusion 682 -1788 682 -1788 0 feedthrough
rlabel pdiffusion 689 -1788 689 -1788 0 feedthrough
rlabel pdiffusion 696 -1788 696 -1788 0 feedthrough
rlabel pdiffusion 703 -1788 703 -1788 0 cellNo=204
rlabel pdiffusion 710 -1788 710 -1788 0 feedthrough
rlabel pdiffusion 717 -1788 717 -1788 0 cellNo=482
rlabel pdiffusion 724 -1788 724 -1788 0 cellNo=303
rlabel pdiffusion 731 -1788 731 -1788 0 cellNo=344
rlabel pdiffusion 738 -1788 738 -1788 0 feedthrough
rlabel pdiffusion 745 -1788 745 -1788 0 feedthrough
rlabel pdiffusion 752 -1788 752 -1788 0 feedthrough
rlabel pdiffusion 759 -1788 759 -1788 0 feedthrough
rlabel pdiffusion 766 -1788 766 -1788 0 feedthrough
rlabel pdiffusion 773 -1788 773 -1788 0 feedthrough
rlabel pdiffusion 780 -1788 780 -1788 0 cellNo=114
rlabel pdiffusion 787 -1788 787 -1788 0 cellNo=421
rlabel pdiffusion 794 -1788 794 -1788 0 feedthrough
rlabel pdiffusion 801 -1788 801 -1788 0 feedthrough
rlabel pdiffusion 808 -1788 808 -1788 0 feedthrough
rlabel pdiffusion 815 -1788 815 -1788 0 feedthrough
rlabel pdiffusion 822 -1788 822 -1788 0 cellNo=916
rlabel pdiffusion 829 -1788 829 -1788 0 feedthrough
rlabel pdiffusion 836 -1788 836 -1788 0 feedthrough
rlabel pdiffusion 843 -1788 843 -1788 0 feedthrough
rlabel pdiffusion 850 -1788 850 -1788 0 feedthrough
rlabel pdiffusion 857 -1788 857 -1788 0 feedthrough
rlabel pdiffusion 864 -1788 864 -1788 0 feedthrough
rlabel pdiffusion 871 -1788 871 -1788 0 feedthrough
rlabel pdiffusion 878 -1788 878 -1788 0 feedthrough
rlabel pdiffusion 885 -1788 885 -1788 0 cellNo=806
rlabel pdiffusion 892 -1788 892 -1788 0 feedthrough
rlabel pdiffusion 899 -1788 899 -1788 0 cellNo=117
rlabel pdiffusion 906 -1788 906 -1788 0 feedthrough
rlabel pdiffusion 913 -1788 913 -1788 0 feedthrough
rlabel pdiffusion 920 -1788 920 -1788 0 feedthrough
rlabel pdiffusion 927 -1788 927 -1788 0 feedthrough
rlabel pdiffusion 934 -1788 934 -1788 0 feedthrough
rlabel pdiffusion 941 -1788 941 -1788 0 feedthrough
rlabel pdiffusion 948 -1788 948 -1788 0 cellNo=597
rlabel pdiffusion 955 -1788 955 -1788 0 feedthrough
rlabel pdiffusion 962 -1788 962 -1788 0 feedthrough
rlabel pdiffusion 969 -1788 969 -1788 0 feedthrough
rlabel pdiffusion 976 -1788 976 -1788 0 cellNo=234
rlabel pdiffusion 983 -1788 983 -1788 0 feedthrough
rlabel pdiffusion 990 -1788 990 -1788 0 feedthrough
rlabel pdiffusion 997 -1788 997 -1788 0 feedthrough
rlabel pdiffusion 1004 -1788 1004 -1788 0 feedthrough
rlabel pdiffusion 1011 -1788 1011 -1788 0 feedthrough
rlabel pdiffusion 1018 -1788 1018 -1788 0 feedthrough
rlabel pdiffusion 1025 -1788 1025 -1788 0 cellNo=939
rlabel pdiffusion 1032 -1788 1032 -1788 0 feedthrough
rlabel pdiffusion 1039 -1788 1039 -1788 0 feedthrough
rlabel pdiffusion 1046 -1788 1046 -1788 0 feedthrough
rlabel pdiffusion 1053 -1788 1053 -1788 0 cellNo=796
rlabel pdiffusion 1060 -1788 1060 -1788 0 feedthrough
rlabel pdiffusion 1067 -1788 1067 -1788 0 feedthrough
rlabel pdiffusion 1074 -1788 1074 -1788 0 feedthrough
rlabel pdiffusion 1081 -1788 1081 -1788 0 feedthrough
rlabel pdiffusion 1088 -1788 1088 -1788 0 feedthrough
rlabel pdiffusion 1095 -1788 1095 -1788 0 feedthrough
rlabel pdiffusion 1102 -1788 1102 -1788 0 feedthrough
rlabel pdiffusion 1109 -1788 1109 -1788 0 feedthrough
rlabel pdiffusion 1116 -1788 1116 -1788 0 feedthrough
rlabel pdiffusion 1123 -1788 1123 -1788 0 feedthrough
rlabel pdiffusion 1130 -1788 1130 -1788 0 feedthrough
rlabel pdiffusion 1137 -1788 1137 -1788 0 feedthrough
rlabel pdiffusion 1144 -1788 1144 -1788 0 cellNo=455
rlabel pdiffusion 1151 -1788 1151 -1788 0 feedthrough
rlabel pdiffusion 1158 -1788 1158 -1788 0 feedthrough
rlabel pdiffusion 1165 -1788 1165 -1788 0 feedthrough
rlabel pdiffusion 1172 -1788 1172 -1788 0 feedthrough
rlabel pdiffusion 1179 -1788 1179 -1788 0 feedthrough
rlabel pdiffusion 1186 -1788 1186 -1788 0 feedthrough
rlabel pdiffusion 1193 -1788 1193 -1788 0 feedthrough
rlabel pdiffusion 1200 -1788 1200 -1788 0 feedthrough
rlabel pdiffusion 1207 -1788 1207 -1788 0 feedthrough
rlabel pdiffusion 1214 -1788 1214 -1788 0 feedthrough
rlabel pdiffusion 1221 -1788 1221 -1788 0 feedthrough
rlabel pdiffusion 1228 -1788 1228 -1788 0 feedthrough
rlabel pdiffusion 1235 -1788 1235 -1788 0 feedthrough
rlabel pdiffusion 1242 -1788 1242 -1788 0 feedthrough
rlabel pdiffusion 1249 -1788 1249 -1788 0 feedthrough
rlabel pdiffusion 1256 -1788 1256 -1788 0 feedthrough
rlabel pdiffusion 1263 -1788 1263 -1788 0 feedthrough
rlabel pdiffusion 1270 -1788 1270 -1788 0 feedthrough
rlabel pdiffusion 1277 -1788 1277 -1788 0 feedthrough
rlabel pdiffusion 1284 -1788 1284 -1788 0 feedthrough
rlabel pdiffusion 1291 -1788 1291 -1788 0 cellNo=511
rlabel pdiffusion 1298 -1788 1298 -1788 0 feedthrough
rlabel pdiffusion 1305 -1788 1305 -1788 0 feedthrough
rlabel pdiffusion 1312 -1788 1312 -1788 0 feedthrough
rlabel pdiffusion 1319 -1788 1319 -1788 0 feedthrough
rlabel pdiffusion 1326 -1788 1326 -1788 0 feedthrough
rlabel pdiffusion 1333 -1788 1333 -1788 0 feedthrough
rlabel pdiffusion 1340 -1788 1340 -1788 0 feedthrough
rlabel pdiffusion 1347 -1788 1347 -1788 0 feedthrough
rlabel pdiffusion 1354 -1788 1354 -1788 0 feedthrough
rlabel pdiffusion 1361 -1788 1361 -1788 0 feedthrough
rlabel pdiffusion 1368 -1788 1368 -1788 0 feedthrough
rlabel pdiffusion 1375 -1788 1375 -1788 0 feedthrough
rlabel pdiffusion 1382 -1788 1382 -1788 0 feedthrough
rlabel pdiffusion 1389 -1788 1389 -1788 0 feedthrough
rlabel pdiffusion 1396 -1788 1396 -1788 0 feedthrough
rlabel pdiffusion 1403 -1788 1403 -1788 0 feedthrough
rlabel pdiffusion 1410 -1788 1410 -1788 0 feedthrough
rlabel pdiffusion 1417 -1788 1417 -1788 0 feedthrough
rlabel pdiffusion 1424 -1788 1424 -1788 0 feedthrough
rlabel pdiffusion 1431 -1788 1431 -1788 0 feedthrough
rlabel pdiffusion 1438 -1788 1438 -1788 0 feedthrough
rlabel pdiffusion 1445 -1788 1445 -1788 0 feedthrough
rlabel pdiffusion 1452 -1788 1452 -1788 0 feedthrough
rlabel pdiffusion 1459 -1788 1459 -1788 0 feedthrough
rlabel pdiffusion 1466 -1788 1466 -1788 0 feedthrough
rlabel pdiffusion 1473 -1788 1473 -1788 0 feedthrough
rlabel pdiffusion 1480 -1788 1480 -1788 0 feedthrough
rlabel pdiffusion 1487 -1788 1487 -1788 0 feedthrough
rlabel pdiffusion 1494 -1788 1494 -1788 0 feedthrough
rlabel pdiffusion 1501 -1788 1501 -1788 0 feedthrough
rlabel pdiffusion 1508 -1788 1508 -1788 0 feedthrough
rlabel pdiffusion 1515 -1788 1515 -1788 0 feedthrough
rlabel pdiffusion 1522 -1788 1522 -1788 0 feedthrough
rlabel pdiffusion 1529 -1788 1529 -1788 0 feedthrough
rlabel pdiffusion 1536 -1788 1536 -1788 0 feedthrough
rlabel pdiffusion 1543 -1788 1543 -1788 0 feedthrough
rlabel pdiffusion 1550 -1788 1550 -1788 0 feedthrough
rlabel pdiffusion 1557 -1788 1557 -1788 0 feedthrough
rlabel pdiffusion 1564 -1788 1564 -1788 0 feedthrough
rlabel pdiffusion 1571 -1788 1571 -1788 0 feedthrough
rlabel pdiffusion 1578 -1788 1578 -1788 0 feedthrough
rlabel pdiffusion 1585 -1788 1585 -1788 0 feedthrough
rlabel pdiffusion 1592 -1788 1592 -1788 0 feedthrough
rlabel pdiffusion 1599 -1788 1599 -1788 0 feedthrough
rlabel pdiffusion 1606 -1788 1606 -1788 0 feedthrough
rlabel pdiffusion 1613 -1788 1613 -1788 0 feedthrough
rlabel pdiffusion 1620 -1788 1620 -1788 0 feedthrough
rlabel pdiffusion 1627 -1788 1627 -1788 0 feedthrough
rlabel pdiffusion 1634 -1788 1634 -1788 0 feedthrough
rlabel pdiffusion 1641 -1788 1641 -1788 0 feedthrough
rlabel pdiffusion 1648 -1788 1648 -1788 0 feedthrough
rlabel pdiffusion 1655 -1788 1655 -1788 0 feedthrough
rlabel pdiffusion 1662 -1788 1662 -1788 0 feedthrough
rlabel pdiffusion 1669 -1788 1669 -1788 0 feedthrough
rlabel pdiffusion 1676 -1788 1676 -1788 0 feedthrough
rlabel pdiffusion 1683 -1788 1683 -1788 0 feedthrough
rlabel pdiffusion 1690 -1788 1690 -1788 0 feedthrough
rlabel pdiffusion 1697 -1788 1697 -1788 0 feedthrough
rlabel pdiffusion 1704 -1788 1704 -1788 0 feedthrough
rlabel pdiffusion 1711 -1788 1711 -1788 0 feedthrough
rlabel pdiffusion 1718 -1788 1718 -1788 0 feedthrough
rlabel pdiffusion 1725 -1788 1725 -1788 0 feedthrough
rlabel pdiffusion 1732 -1788 1732 -1788 0 feedthrough
rlabel pdiffusion 1739 -1788 1739 -1788 0 feedthrough
rlabel pdiffusion 1746 -1788 1746 -1788 0 feedthrough
rlabel pdiffusion 1753 -1788 1753 -1788 0 feedthrough
rlabel pdiffusion 1760 -1788 1760 -1788 0 feedthrough
rlabel pdiffusion 1767 -1788 1767 -1788 0 feedthrough
rlabel pdiffusion 1774 -1788 1774 -1788 0 feedthrough
rlabel pdiffusion 1781 -1788 1781 -1788 0 feedthrough
rlabel pdiffusion 1788 -1788 1788 -1788 0 feedthrough
rlabel pdiffusion 1795 -1788 1795 -1788 0 feedthrough
rlabel pdiffusion 1802 -1788 1802 -1788 0 feedthrough
rlabel pdiffusion 1809 -1788 1809 -1788 0 feedthrough
rlabel pdiffusion 1816 -1788 1816 -1788 0 feedthrough
rlabel pdiffusion 1823 -1788 1823 -1788 0 feedthrough
rlabel pdiffusion 1830 -1788 1830 -1788 0 feedthrough
rlabel pdiffusion 1837 -1788 1837 -1788 0 cellNo=367
rlabel pdiffusion 3 -1927 3 -1927 0 cellNo=1117
rlabel pdiffusion 10 -1927 10 -1927 0 cellNo=1121
rlabel pdiffusion 17 -1927 17 -1927 0 cellNo=1127
rlabel pdiffusion 24 -1927 24 -1927 0 cellNo=1133
rlabel pdiffusion 31 -1927 31 -1927 0 feedthrough
rlabel pdiffusion 38 -1927 38 -1927 0 feedthrough
rlabel pdiffusion 45 -1927 45 -1927 0 feedthrough
rlabel pdiffusion 52 -1927 52 -1927 0 feedthrough
rlabel pdiffusion 59 -1927 59 -1927 0 cellNo=943
rlabel pdiffusion 66 -1927 66 -1927 0 cellNo=891
rlabel pdiffusion 73 -1927 73 -1927 0 feedthrough
rlabel pdiffusion 80 -1927 80 -1927 0 feedthrough
rlabel pdiffusion 87 -1927 87 -1927 0 feedthrough
rlabel pdiffusion 94 -1927 94 -1927 0 feedthrough
rlabel pdiffusion 101 -1927 101 -1927 0 feedthrough
rlabel pdiffusion 108 -1927 108 -1927 0 cellNo=137
rlabel pdiffusion 115 -1927 115 -1927 0 feedthrough
rlabel pdiffusion 122 -1927 122 -1927 0 feedthrough
rlabel pdiffusion 129 -1927 129 -1927 0 feedthrough
rlabel pdiffusion 136 -1927 136 -1927 0 feedthrough
rlabel pdiffusion 143 -1927 143 -1927 0 feedthrough
rlabel pdiffusion 150 -1927 150 -1927 0 feedthrough
rlabel pdiffusion 157 -1927 157 -1927 0 feedthrough
rlabel pdiffusion 164 -1927 164 -1927 0 feedthrough
rlabel pdiffusion 171 -1927 171 -1927 0 cellNo=258
rlabel pdiffusion 178 -1927 178 -1927 0 feedthrough
rlabel pdiffusion 185 -1927 185 -1927 0 feedthrough
rlabel pdiffusion 192 -1927 192 -1927 0 feedthrough
rlabel pdiffusion 199 -1927 199 -1927 0 feedthrough
rlabel pdiffusion 206 -1927 206 -1927 0 feedthrough
rlabel pdiffusion 213 -1927 213 -1927 0 feedthrough
rlabel pdiffusion 220 -1927 220 -1927 0 cellNo=678
rlabel pdiffusion 227 -1927 227 -1927 0 cellNo=726
rlabel pdiffusion 234 -1927 234 -1927 0 feedthrough
rlabel pdiffusion 241 -1927 241 -1927 0 cellNo=770
rlabel pdiffusion 248 -1927 248 -1927 0 cellNo=962
rlabel pdiffusion 255 -1927 255 -1927 0 feedthrough
rlabel pdiffusion 262 -1927 262 -1927 0 feedthrough
rlabel pdiffusion 269 -1927 269 -1927 0 feedthrough
rlabel pdiffusion 276 -1927 276 -1927 0 feedthrough
rlabel pdiffusion 283 -1927 283 -1927 0 feedthrough
rlabel pdiffusion 290 -1927 290 -1927 0 feedthrough
rlabel pdiffusion 297 -1927 297 -1927 0 feedthrough
rlabel pdiffusion 304 -1927 304 -1927 0 feedthrough
rlabel pdiffusion 311 -1927 311 -1927 0 feedthrough
rlabel pdiffusion 318 -1927 318 -1927 0 feedthrough
rlabel pdiffusion 325 -1927 325 -1927 0 feedthrough
rlabel pdiffusion 332 -1927 332 -1927 0 feedthrough
rlabel pdiffusion 339 -1927 339 -1927 0 cellNo=664
rlabel pdiffusion 346 -1927 346 -1927 0 feedthrough
rlabel pdiffusion 353 -1927 353 -1927 0 feedthrough
rlabel pdiffusion 360 -1927 360 -1927 0 feedthrough
rlabel pdiffusion 367 -1927 367 -1927 0 feedthrough
rlabel pdiffusion 374 -1927 374 -1927 0 feedthrough
rlabel pdiffusion 381 -1927 381 -1927 0 feedthrough
rlabel pdiffusion 388 -1927 388 -1927 0 feedthrough
rlabel pdiffusion 395 -1927 395 -1927 0 feedthrough
rlabel pdiffusion 402 -1927 402 -1927 0 cellNo=210
rlabel pdiffusion 409 -1927 409 -1927 0 feedthrough
rlabel pdiffusion 416 -1927 416 -1927 0 feedthrough
rlabel pdiffusion 423 -1927 423 -1927 0 feedthrough
rlabel pdiffusion 430 -1927 430 -1927 0 cellNo=366
rlabel pdiffusion 437 -1927 437 -1927 0 feedthrough
rlabel pdiffusion 444 -1927 444 -1927 0 feedthrough
rlabel pdiffusion 451 -1927 451 -1927 0 feedthrough
rlabel pdiffusion 458 -1927 458 -1927 0 feedthrough
rlabel pdiffusion 465 -1927 465 -1927 0 feedthrough
rlabel pdiffusion 472 -1927 472 -1927 0 feedthrough
rlabel pdiffusion 479 -1927 479 -1927 0 feedthrough
rlabel pdiffusion 486 -1927 486 -1927 0 feedthrough
rlabel pdiffusion 493 -1927 493 -1927 0 feedthrough
rlabel pdiffusion 500 -1927 500 -1927 0 feedthrough
rlabel pdiffusion 507 -1927 507 -1927 0 feedthrough
rlabel pdiffusion 514 -1927 514 -1927 0 feedthrough
rlabel pdiffusion 521 -1927 521 -1927 0 feedthrough
rlabel pdiffusion 528 -1927 528 -1927 0 cellNo=472
rlabel pdiffusion 535 -1927 535 -1927 0 feedthrough
rlabel pdiffusion 542 -1927 542 -1927 0 feedthrough
rlabel pdiffusion 549 -1927 549 -1927 0 feedthrough
rlabel pdiffusion 556 -1927 556 -1927 0 feedthrough
rlabel pdiffusion 563 -1927 563 -1927 0 feedthrough
rlabel pdiffusion 570 -1927 570 -1927 0 feedthrough
rlabel pdiffusion 577 -1927 577 -1927 0 feedthrough
rlabel pdiffusion 584 -1927 584 -1927 0 feedthrough
rlabel pdiffusion 591 -1927 591 -1927 0 cellNo=558
rlabel pdiffusion 598 -1927 598 -1927 0 feedthrough
rlabel pdiffusion 605 -1927 605 -1927 0 feedthrough
rlabel pdiffusion 612 -1927 612 -1927 0 feedthrough
rlabel pdiffusion 619 -1927 619 -1927 0 cellNo=446
rlabel pdiffusion 626 -1927 626 -1927 0 feedthrough
rlabel pdiffusion 633 -1927 633 -1927 0 feedthrough
rlabel pdiffusion 640 -1927 640 -1927 0 feedthrough
rlabel pdiffusion 647 -1927 647 -1927 0 feedthrough
rlabel pdiffusion 654 -1927 654 -1927 0 cellNo=773
rlabel pdiffusion 661 -1927 661 -1927 0 feedthrough
rlabel pdiffusion 668 -1927 668 -1927 0 cellNo=808
rlabel pdiffusion 675 -1927 675 -1927 0 feedthrough
rlabel pdiffusion 682 -1927 682 -1927 0 cellNo=961
rlabel pdiffusion 689 -1927 689 -1927 0 feedthrough
rlabel pdiffusion 696 -1927 696 -1927 0 feedthrough
rlabel pdiffusion 703 -1927 703 -1927 0 feedthrough
rlabel pdiffusion 710 -1927 710 -1927 0 feedthrough
rlabel pdiffusion 717 -1927 717 -1927 0 feedthrough
rlabel pdiffusion 724 -1927 724 -1927 0 cellNo=648
rlabel pdiffusion 731 -1927 731 -1927 0 feedthrough
rlabel pdiffusion 738 -1927 738 -1927 0 feedthrough
rlabel pdiffusion 745 -1927 745 -1927 0 feedthrough
rlabel pdiffusion 752 -1927 752 -1927 0 feedthrough
rlabel pdiffusion 759 -1927 759 -1927 0 feedthrough
rlabel pdiffusion 766 -1927 766 -1927 0 feedthrough
rlabel pdiffusion 773 -1927 773 -1927 0 cellNo=531
rlabel pdiffusion 780 -1927 780 -1927 0 feedthrough
rlabel pdiffusion 787 -1927 787 -1927 0 cellNo=243
rlabel pdiffusion 794 -1927 794 -1927 0 feedthrough
rlabel pdiffusion 801 -1927 801 -1927 0 feedthrough
rlabel pdiffusion 808 -1927 808 -1927 0 cellNo=658
rlabel pdiffusion 815 -1927 815 -1927 0 feedthrough
rlabel pdiffusion 822 -1927 822 -1927 0 feedthrough
rlabel pdiffusion 829 -1927 829 -1927 0 cellNo=144
rlabel pdiffusion 836 -1927 836 -1927 0 feedthrough
rlabel pdiffusion 843 -1927 843 -1927 0 feedthrough
rlabel pdiffusion 850 -1927 850 -1927 0 cellNo=430
rlabel pdiffusion 857 -1927 857 -1927 0 feedthrough
rlabel pdiffusion 864 -1927 864 -1927 0 feedthrough
rlabel pdiffusion 871 -1927 871 -1927 0 cellNo=556
rlabel pdiffusion 878 -1927 878 -1927 0 feedthrough
rlabel pdiffusion 885 -1927 885 -1927 0 feedthrough
rlabel pdiffusion 892 -1927 892 -1927 0 feedthrough
rlabel pdiffusion 899 -1927 899 -1927 0 feedthrough
rlabel pdiffusion 906 -1927 906 -1927 0 feedthrough
rlabel pdiffusion 913 -1927 913 -1927 0 cellNo=392
rlabel pdiffusion 920 -1927 920 -1927 0 feedthrough
rlabel pdiffusion 927 -1927 927 -1927 0 feedthrough
rlabel pdiffusion 934 -1927 934 -1927 0 feedthrough
rlabel pdiffusion 941 -1927 941 -1927 0 feedthrough
rlabel pdiffusion 948 -1927 948 -1927 0 feedthrough
rlabel pdiffusion 955 -1927 955 -1927 0 feedthrough
rlabel pdiffusion 962 -1927 962 -1927 0 feedthrough
rlabel pdiffusion 969 -1927 969 -1927 0 feedthrough
rlabel pdiffusion 976 -1927 976 -1927 0 feedthrough
rlabel pdiffusion 983 -1927 983 -1927 0 cellNo=636
rlabel pdiffusion 990 -1927 990 -1927 0 cellNo=982
rlabel pdiffusion 997 -1927 997 -1927 0 feedthrough
rlabel pdiffusion 1004 -1927 1004 -1927 0 feedthrough
rlabel pdiffusion 1011 -1927 1011 -1927 0 feedthrough
rlabel pdiffusion 1018 -1927 1018 -1927 0 feedthrough
rlabel pdiffusion 1025 -1927 1025 -1927 0 feedthrough
rlabel pdiffusion 1032 -1927 1032 -1927 0 feedthrough
rlabel pdiffusion 1039 -1927 1039 -1927 0 feedthrough
rlabel pdiffusion 1046 -1927 1046 -1927 0 feedthrough
rlabel pdiffusion 1053 -1927 1053 -1927 0 feedthrough
rlabel pdiffusion 1060 -1927 1060 -1927 0 feedthrough
rlabel pdiffusion 1067 -1927 1067 -1927 0 feedthrough
rlabel pdiffusion 1074 -1927 1074 -1927 0 feedthrough
rlabel pdiffusion 1081 -1927 1081 -1927 0 feedthrough
rlabel pdiffusion 1088 -1927 1088 -1927 0 feedthrough
rlabel pdiffusion 1095 -1927 1095 -1927 0 cellNo=479
rlabel pdiffusion 1102 -1927 1102 -1927 0 feedthrough
rlabel pdiffusion 1109 -1927 1109 -1927 0 feedthrough
rlabel pdiffusion 1116 -1927 1116 -1927 0 feedthrough
rlabel pdiffusion 1123 -1927 1123 -1927 0 cellNo=165
rlabel pdiffusion 1130 -1927 1130 -1927 0 feedthrough
rlabel pdiffusion 1137 -1927 1137 -1927 0 feedthrough
rlabel pdiffusion 1144 -1927 1144 -1927 0 feedthrough
rlabel pdiffusion 1151 -1927 1151 -1927 0 feedthrough
rlabel pdiffusion 1158 -1927 1158 -1927 0 cellNo=653
rlabel pdiffusion 1165 -1927 1165 -1927 0 cellNo=903
rlabel pdiffusion 1172 -1927 1172 -1927 0 feedthrough
rlabel pdiffusion 1179 -1927 1179 -1927 0 feedthrough
rlabel pdiffusion 1186 -1927 1186 -1927 0 feedthrough
rlabel pdiffusion 1193 -1927 1193 -1927 0 feedthrough
rlabel pdiffusion 1200 -1927 1200 -1927 0 feedthrough
rlabel pdiffusion 1207 -1927 1207 -1927 0 feedthrough
rlabel pdiffusion 1214 -1927 1214 -1927 0 feedthrough
rlabel pdiffusion 1221 -1927 1221 -1927 0 feedthrough
rlabel pdiffusion 1228 -1927 1228 -1927 0 cellNo=163
rlabel pdiffusion 1235 -1927 1235 -1927 0 feedthrough
rlabel pdiffusion 1242 -1927 1242 -1927 0 feedthrough
rlabel pdiffusion 1249 -1927 1249 -1927 0 feedthrough
rlabel pdiffusion 1256 -1927 1256 -1927 0 feedthrough
rlabel pdiffusion 1263 -1927 1263 -1927 0 feedthrough
rlabel pdiffusion 1270 -1927 1270 -1927 0 feedthrough
rlabel pdiffusion 1277 -1927 1277 -1927 0 feedthrough
rlabel pdiffusion 1284 -1927 1284 -1927 0 feedthrough
rlabel pdiffusion 1291 -1927 1291 -1927 0 feedthrough
rlabel pdiffusion 1298 -1927 1298 -1927 0 feedthrough
rlabel pdiffusion 1305 -1927 1305 -1927 0 feedthrough
rlabel pdiffusion 1312 -1927 1312 -1927 0 feedthrough
rlabel pdiffusion 1319 -1927 1319 -1927 0 feedthrough
rlabel pdiffusion 1326 -1927 1326 -1927 0 feedthrough
rlabel pdiffusion 1333 -1927 1333 -1927 0 feedthrough
rlabel pdiffusion 1340 -1927 1340 -1927 0 feedthrough
rlabel pdiffusion 1347 -1927 1347 -1927 0 feedthrough
rlabel pdiffusion 1354 -1927 1354 -1927 0 feedthrough
rlabel pdiffusion 1361 -1927 1361 -1927 0 feedthrough
rlabel pdiffusion 1368 -1927 1368 -1927 0 feedthrough
rlabel pdiffusion 1375 -1927 1375 -1927 0 feedthrough
rlabel pdiffusion 1382 -1927 1382 -1927 0 cellNo=480
rlabel pdiffusion 1389 -1927 1389 -1927 0 feedthrough
rlabel pdiffusion 1396 -1927 1396 -1927 0 feedthrough
rlabel pdiffusion 1403 -1927 1403 -1927 0 feedthrough
rlabel pdiffusion 1410 -1927 1410 -1927 0 feedthrough
rlabel pdiffusion 1417 -1927 1417 -1927 0 feedthrough
rlabel pdiffusion 1424 -1927 1424 -1927 0 feedthrough
rlabel pdiffusion 1431 -1927 1431 -1927 0 feedthrough
rlabel pdiffusion 1438 -1927 1438 -1927 0 feedthrough
rlabel pdiffusion 1445 -1927 1445 -1927 0 feedthrough
rlabel pdiffusion 1452 -1927 1452 -1927 0 feedthrough
rlabel pdiffusion 1459 -1927 1459 -1927 0 feedthrough
rlabel pdiffusion 1466 -1927 1466 -1927 0 feedthrough
rlabel pdiffusion 1473 -1927 1473 -1927 0 feedthrough
rlabel pdiffusion 1480 -1927 1480 -1927 0 feedthrough
rlabel pdiffusion 1487 -1927 1487 -1927 0 feedthrough
rlabel pdiffusion 1494 -1927 1494 -1927 0 feedthrough
rlabel pdiffusion 1501 -1927 1501 -1927 0 feedthrough
rlabel pdiffusion 1508 -1927 1508 -1927 0 feedthrough
rlabel pdiffusion 1515 -1927 1515 -1927 0 feedthrough
rlabel pdiffusion 1522 -1927 1522 -1927 0 feedthrough
rlabel pdiffusion 1529 -1927 1529 -1927 0 feedthrough
rlabel pdiffusion 1536 -1927 1536 -1927 0 feedthrough
rlabel pdiffusion 1543 -1927 1543 -1927 0 feedthrough
rlabel pdiffusion 1550 -1927 1550 -1927 0 feedthrough
rlabel pdiffusion 1557 -1927 1557 -1927 0 feedthrough
rlabel pdiffusion 1564 -1927 1564 -1927 0 feedthrough
rlabel pdiffusion 1571 -1927 1571 -1927 0 feedthrough
rlabel pdiffusion 1578 -1927 1578 -1927 0 feedthrough
rlabel pdiffusion 1585 -1927 1585 -1927 0 feedthrough
rlabel pdiffusion 1592 -1927 1592 -1927 0 feedthrough
rlabel pdiffusion 1599 -1927 1599 -1927 0 feedthrough
rlabel pdiffusion 1606 -1927 1606 -1927 0 feedthrough
rlabel pdiffusion 1613 -1927 1613 -1927 0 feedthrough
rlabel pdiffusion 1620 -1927 1620 -1927 0 feedthrough
rlabel pdiffusion 1627 -1927 1627 -1927 0 feedthrough
rlabel pdiffusion 1634 -1927 1634 -1927 0 feedthrough
rlabel pdiffusion 1641 -1927 1641 -1927 0 feedthrough
rlabel pdiffusion 1648 -1927 1648 -1927 0 feedthrough
rlabel pdiffusion 1655 -1927 1655 -1927 0 feedthrough
rlabel pdiffusion 1662 -1927 1662 -1927 0 feedthrough
rlabel pdiffusion 1669 -1927 1669 -1927 0 feedthrough
rlabel pdiffusion 1676 -1927 1676 -1927 0 feedthrough
rlabel pdiffusion 1683 -1927 1683 -1927 0 feedthrough
rlabel pdiffusion 1690 -1927 1690 -1927 0 feedthrough
rlabel pdiffusion 1697 -1927 1697 -1927 0 feedthrough
rlabel pdiffusion 1704 -1927 1704 -1927 0 feedthrough
rlabel pdiffusion 1711 -1927 1711 -1927 0 feedthrough
rlabel pdiffusion 1718 -1927 1718 -1927 0 feedthrough
rlabel pdiffusion 1725 -1927 1725 -1927 0 feedthrough
rlabel pdiffusion 1732 -1927 1732 -1927 0 feedthrough
rlabel pdiffusion 1739 -1927 1739 -1927 0 feedthrough
rlabel pdiffusion 1746 -1927 1746 -1927 0 feedthrough
rlabel pdiffusion 1753 -1927 1753 -1927 0 cellNo=880
rlabel pdiffusion 1760 -1927 1760 -1927 0 feedthrough
rlabel pdiffusion 1767 -1927 1767 -1927 0 feedthrough
rlabel pdiffusion 1795 -1927 1795 -1927 0 feedthrough
rlabel pdiffusion 3 -2054 3 -2054 0 cellNo=1120
rlabel pdiffusion 10 -2054 10 -2054 0 cellNo=1125
rlabel pdiffusion 17 -2054 17 -2054 0 cellNo=1131
rlabel pdiffusion 24 -2054 24 -2054 0 feedthrough
rlabel pdiffusion 31 -2054 31 -2054 0 cellNo=1142
rlabel pdiffusion 38 -2054 38 -2054 0 feedthrough
rlabel pdiffusion 45 -2054 45 -2054 0 feedthrough
rlabel pdiffusion 52 -2054 52 -2054 0 feedthrough
rlabel pdiffusion 59 -2054 59 -2054 0 feedthrough
rlabel pdiffusion 66 -2054 66 -2054 0 feedthrough
rlabel pdiffusion 73 -2054 73 -2054 0 feedthrough
rlabel pdiffusion 80 -2054 80 -2054 0 feedthrough
rlabel pdiffusion 87 -2054 87 -2054 0 feedthrough
rlabel pdiffusion 94 -2054 94 -2054 0 feedthrough
rlabel pdiffusion 101 -2054 101 -2054 0 feedthrough
rlabel pdiffusion 108 -2054 108 -2054 0 cellNo=79
rlabel pdiffusion 115 -2054 115 -2054 0 cellNo=832
rlabel pdiffusion 122 -2054 122 -2054 0 feedthrough
rlabel pdiffusion 129 -2054 129 -2054 0 cellNo=951
rlabel pdiffusion 136 -2054 136 -2054 0 cellNo=369
rlabel pdiffusion 143 -2054 143 -2054 0 feedthrough
rlabel pdiffusion 150 -2054 150 -2054 0 feedthrough
rlabel pdiffusion 157 -2054 157 -2054 0 cellNo=827
rlabel pdiffusion 164 -2054 164 -2054 0 cellNo=969
rlabel pdiffusion 171 -2054 171 -2054 0 feedthrough
rlabel pdiffusion 178 -2054 178 -2054 0 feedthrough
rlabel pdiffusion 185 -2054 185 -2054 0 feedthrough
rlabel pdiffusion 192 -2054 192 -2054 0 feedthrough
rlabel pdiffusion 199 -2054 199 -2054 0 feedthrough
rlabel pdiffusion 206 -2054 206 -2054 0 cellNo=182
rlabel pdiffusion 213 -2054 213 -2054 0 feedthrough
rlabel pdiffusion 220 -2054 220 -2054 0 feedthrough
rlabel pdiffusion 227 -2054 227 -2054 0 feedthrough
rlabel pdiffusion 234 -2054 234 -2054 0 feedthrough
rlabel pdiffusion 241 -2054 241 -2054 0 feedthrough
rlabel pdiffusion 248 -2054 248 -2054 0 feedthrough
rlabel pdiffusion 255 -2054 255 -2054 0 feedthrough
rlabel pdiffusion 262 -2054 262 -2054 0 feedthrough
rlabel pdiffusion 269 -2054 269 -2054 0 feedthrough
rlabel pdiffusion 276 -2054 276 -2054 0 feedthrough
rlabel pdiffusion 283 -2054 283 -2054 0 feedthrough
rlabel pdiffusion 290 -2054 290 -2054 0 feedthrough
rlabel pdiffusion 297 -2054 297 -2054 0 feedthrough
rlabel pdiffusion 304 -2054 304 -2054 0 feedthrough
rlabel pdiffusion 311 -2054 311 -2054 0 feedthrough
rlabel pdiffusion 318 -2054 318 -2054 0 feedthrough
rlabel pdiffusion 325 -2054 325 -2054 0 feedthrough
rlabel pdiffusion 332 -2054 332 -2054 0 feedthrough
rlabel pdiffusion 339 -2054 339 -2054 0 feedthrough
rlabel pdiffusion 346 -2054 346 -2054 0 feedthrough
rlabel pdiffusion 353 -2054 353 -2054 0 feedthrough
rlabel pdiffusion 360 -2054 360 -2054 0 feedthrough
rlabel pdiffusion 367 -2054 367 -2054 0 cellNo=147
rlabel pdiffusion 374 -2054 374 -2054 0 feedthrough
rlabel pdiffusion 381 -2054 381 -2054 0 feedthrough
rlabel pdiffusion 388 -2054 388 -2054 0 feedthrough
rlabel pdiffusion 395 -2054 395 -2054 0 feedthrough
rlabel pdiffusion 402 -2054 402 -2054 0 feedthrough
rlabel pdiffusion 409 -2054 409 -2054 0 feedthrough
rlabel pdiffusion 416 -2054 416 -2054 0 feedthrough
rlabel pdiffusion 423 -2054 423 -2054 0 feedthrough
rlabel pdiffusion 430 -2054 430 -2054 0 feedthrough
rlabel pdiffusion 437 -2054 437 -2054 0 feedthrough
rlabel pdiffusion 444 -2054 444 -2054 0 feedthrough
rlabel pdiffusion 451 -2054 451 -2054 0 feedthrough
rlabel pdiffusion 458 -2054 458 -2054 0 feedthrough
rlabel pdiffusion 465 -2054 465 -2054 0 feedthrough
rlabel pdiffusion 472 -2054 472 -2054 0 feedthrough
rlabel pdiffusion 479 -2054 479 -2054 0 feedthrough
rlabel pdiffusion 486 -2054 486 -2054 0 feedthrough
rlabel pdiffusion 493 -2054 493 -2054 0 feedthrough
rlabel pdiffusion 500 -2054 500 -2054 0 feedthrough
rlabel pdiffusion 507 -2054 507 -2054 0 feedthrough
rlabel pdiffusion 514 -2054 514 -2054 0 feedthrough
rlabel pdiffusion 521 -2054 521 -2054 0 feedthrough
rlabel pdiffusion 528 -2054 528 -2054 0 cellNo=667
rlabel pdiffusion 535 -2054 535 -2054 0 feedthrough
rlabel pdiffusion 542 -2054 542 -2054 0 feedthrough
rlabel pdiffusion 549 -2054 549 -2054 0 feedthrough
rlabel pdiffusion 556 -2054 556 -2054 0 feedthrough
rlabel pdiffusion 563 -2054 563 -2054 0 feedthrough
rlabel pdiffusion 570 -2054 570 -2054 0 feedthrough
rlabel pdiffusion 577 -2054 577 -2054 0 feedthrough
rlabel pdiffusion 584 -2054 584 -2054 0 feedthrough
rlabel pdiffusion 591 -2054 591 -2054 0 cellNo=797
rlabel pdiffusion 598 -2054 598 -2054 0 cellNo=485
rlabel pdiffusion 605 -2054 605 -2054 0 cellNo=220
rlabel pdiffusion 612 -2054 612 -2054 0 feedthrough
rlabel pdiffusion 619 -2054 619 -2054 0 cellNo=53
rlabel pdiffusion 626 -2054 626 -2054 0 feedthrough
rlabel pdiffusion 633 -2054 633 -2054 0 cellNo=398
rlabel pdiffusion 640 -2054 640 -2054 0 feedthrough
rlabel pdiffusion 647 -2054 647 -2054 0 feedthrough
rlabel pdiffusion 654 -2054 654 -2054 0 feedthrough
rlabel pdiffusion 661 -2054 661 -2054 0 cellNo=734
rlabel pdiffusion 668 -2054 668 -2054 0 cellNo=681
rlabel pdiffusion 675 -2054 675 -2054 0 feedthrough
rlabel pdiffusion 682 -2054 682 -2054 0 feedthrough
rlabel pdiffusion 689 -2054 689 -2054 0 cellNo=627
rlabel pdiffusion 696 -2054 696 -2054 0 feedthrough
rlabel pdiffusion 703 -2054 703 -2054 0 feedthrough
rlabel pdiffusion 710 -2054 710 -2054 0 feedthrough
rlabel pdiffusion 717 -2054 717 -2054 0 feedthrough
rlabel pdiffusion 724 -2054 724 -2054 0 feedthrough
rlabel pdiffusion 731 -2054 731 -2054 0 feedthrough
rlabel pdiffusion 738 -2054 738 -2054 0 feedthrough
rlabel pdiffusion 745 -2054 745 -2054 0 feedthrough
rlabel pdiffusion 752 -2054 752 -2054 0 cellNo=41
rlabel pdiffusion 759 -2054 759 -2054 0 feedthrough
rlabel pdiffusion 766 -2054 766 -2054 0 cellNo=273
rlabel pdiffusion 773 -2054 773 -2054 0 feedthrough
rlabel pdiffusion 780 -2054 780 -2054 0 cellNo=159
rlabel pdiffusion 787 -2054 787 -2054 0 feedthrough
rlabel pdiffusion 794 -2054 794 -2054 0 feedthrough
rlabel pdiffusion 801 -2054 801 -2054 0 cellNo=198
rlabel pdiffusion 808 -2054 808 -2054 0 feedthrough
rlabel pdiffusion 815 -2054 815 -2054 0 cellNo=787
rlabel pdiffusion 822 -2054 822 -2054 0 feedthrough
rlabel pdiffusion 829 -2054 829 -2054 0 feedthrough
rlabel pdiffusion 836 -2054 836 -2054 0 feedthrough
rlabel pdiffusion 843 -2054 843 -2054 0 feedthrough
rlabel pdiffusion 850 -2054 850 -2054 0 feedthrough
rlabel pdiffusion 857 -2054 857 -2054 0 feedthrough
rlabel pdiffusion 864 -2054 864 -2054 0 feedthrough
rlabel pdiffusion 871 -2054 871 -2054 0 feedthrough
rlabel pdiffusion 878 -2054 878 -2054 0 feedthrough
rlabel pdiffusion 885 -2054 885 -2054 0 feedthrough
rlabel pdiffusion 892 -2054 892 -2054 0 feedthrough
rlabel pdiffusion 899 -2054 899 -2054 0 feedthrough
rlabel pdiffusion 906 -2054 906 -2054 0 cellNo=338
rlabel pdiffusion 913 -2054 913 -2054 0 feedthrough
rlabel pdiffusion 920 -2054 920 -2054 0 feedthrough
rlabel pdiffusion 927 -2054 927 -2054 0 cellNo=851
rlabel pdiffusion 934 -2054 934 -2054 0 cellNo=460
rlabel pdiffusion 941 -2054 941 -2054 0 feedthrough
rlabel pdiffusion 948 -2054 948 -2054 0 cellNo=744
rlabel pdiffusion 955 -2054 955 -2054 0 feedthrough
rlabel pdiffusion 962 -2054 962 -2054 0 feedthrough
rlabel pdiffusion 969 -2054 969 -2054 0 feedthrough
rlabel pdiffusion 976 -2054 976 -2054 0 feedthrough
rlabel pdiffusion 983 -2054 983 -2054 0 cellNo=403
rlabel pdiffusion 990 -2054 990 -2054 0 feedthrough
rlabel pdiffusion 997 -2054 997 -2054 0 feedthrough
rlabel pdiffusion 1004 -2054 1004 -2054 0 feedthrough
rlabel pdiffusion 1011 -2054 1011 -2054 0 feedthrough
rlabel pdiffusion 1018 -2054 1018 -2054 0 cellNo=75
rlabel pdiffusion 1025 -2054 1025 -2054 0 feedthrough
rlabel pdiffusion 1032 -2054 1032 -2054 0 feedthrough
rlabel pdiffusion 1039 -2054 1039 -2054 0 feedthrough
rlabel pdiffusion 1046 -2054 1046 -2054 0 feedthrough
rlabel pdiffusion 1053 -2054 1053 -2054 0 feedthrough
rlabel pdiffusion 1060 -2054 1060 -2054 0 feedthrough
rlabel pdiffusion 1067 -2054 1067 -2054 0 feedthrough
rlabel pdiffusion 1074 -2054 1074 -2054 0 feedthrough
rlabel pdiffusion 1081 -2054 1081 -2054 0 feedthrough
rlabel pdiffusion 1088 -2054 1088 -2054 0 cellNo=719
rlabel pdiffusion 1095 -2054 1095 -2054 0 feedthrough
rlabel pdiffusion 1102 -2054 1102 -2054 0 feedthrough
rlabel pdiffusion 1109 -2054 1109 -2054 0 feedthrough
rlabel pdiffusion 1116 -2054 1116 -2054 0 feedthrough
rlabel pdiffusion 1123 -2054 1123 -2054 0 feedthrough
rlabel pdiffusion 1130 -2054 1130 -2054 0 feedthrough
rlabel pdiffusion 1137 -2054 1137 -2054 0 feedthrough
rlabel pdiffusion 1144 -2054 1144 -2054 0 feedthrough
rlabel pdiffusion 1151 -2054 1151 -2054 0 feedthrough
rlabel pdiffusion 1158 -2054 1158 -2054 0 feedthrough
rlabel pdiffusion 1165 -2054 1165 -2054 0 feedthrough
rlabel pdiffusion 1172 -2054 1172 -2054 0 feedthrough
rlabel pdiffusion 1179 -2054 1179 -2054 0 feedthrough
rlabel pdiffusion 1186 -2054 1186 -2054 0 feedthrough
rlabel pdiffusion 1193 -2054 1193 -2054 0 feedthrough
rlabel pdiffusion 1200 -2054 1200 -2054 0 feedthrough
rlabel pdiffusion 1207 -2054 1207 -2054 0 feedthrough
rlabel pdiffusion 1214 -2054 1214 -2054 0 feedthrough
rlabel pdiffusion 1221 -2054 1221 -2054 0 feedthrough
rlabel pdiffusion 1228 -2054 1228 -2054 0 feedthrough
rlabel pdiffusion 1235 -2054 1235 -2054 0 feedthrough
rlabel pdiffusion 1242 -2054 1242 -2054 0 feedthrough
rlabel pdiffusion 1249 -2054 1249 -2054 0 feedthrough
rlabel pdiffusion 1256 -2054 1256 -2054 0 cellNo=354
rlabel pdiffusion 1263 -2054 1263 -2054 0 feedthrough
rlabel pdiffusion 1270 -2054 1270 -2054 0 feedthrough
rlabel pdiffusion 1277 -2054 1277 -2054 0 feedthrough
rlabel pdiffusion 1284 -2054 1284 -2054 0 feedthrough
rlabel pdiffusion 1291 -2054 1291 -2054 0 feedthrough
rlabel pdiffusion 1298 -2054 1298 -2054 0 feedthrough
rlabel pdiffusion 1305 -2054 1305 -2054 0 feedthrough
rlabel pdiffusion 1312 -2054 1312 -2054 0 feedthrough
rlabel pdiffusion 1319 -2054 1319 -2054 0 feedthrough
rlabel pdiffusion 1326 -2054 1326 -2054 0 feedthrough
rlabel pdiffusion 1333 -2054 1333 -2054 0 feedthrough
rlabel pdiffusion 1340 -2054 1340 -2054 0 feedthrough
rlabel pdiffusion 1347 -2054 1347 -2054 0 feedthrough
rlabel pdiffusion 1354 -2054 1354 -2054 0 feedthrough
rlabel pdiffusion 1361 -2054 1361 -2054 0 feedthrough
rlabel pdiffusion 1368 -2054 1368 -2054 0 feedthrough
rlabel pdiffusion 1375 -2054 1375 -2054 0 feedthrough
rlabel pdiffusion 1382 -2054 1382 -2054 0 feedthrough
rlabel pdiffusion 1389 -2054 1389 -2054 0 feedthrough
rlabel pdiffusion 1396 -2054 1396 -2054 0 feedthrough
rlabel pdiffusion 1403 -2054 1403 -2054 0 feedthrough
rlabel pdiffusion 1410 -2054 1410 -2054 0 feedthrough
rlabel pdiffusion 1417 -2054 1417 -2054 0 feedthrough
rlabel pdiffusion 1424 -2054 1424 -2054 0 feedthrough
rlabel pdiffusion 1431 -2054 1431 -2054 0 feedthrough
rlabel pdiffusion 1438 -2054 1438 -2054 0 feedthrough
rlabel pdiffusion 1445 -2054 1445 -2054 0 feedthrough
rlabel pdiffusion 1452 -2054 1452 -2054 0 cellNo=260
rlabel pdiffusion 1459 -2054 1459 -2054 0 feedthrough
rlabel pdiffusion 1466 -2054 1466 -2054 0 feedthrough
rlabel pdiffusion 1473 -2054 1473 -2054 0 feedthrough
rlabel pdiffusion 1480 -2054 1480 -2054 0 feedthrough
rlabel pdiffusion 1487 -2054 1487 -2054 0 feedthrough
rlabel pdiffusion 1494 -2054 1494 -2054 0 feedthrough
rlabel pdiffusion 1501 -2054 1501 -2054 0 feedthrough
rlabel pdiffusion 1508 -2054 1508 -2054 0 feedthrough
rlabel pdiffusion 1515 -2054 1515 -2054 0 feedthrough
rlabel pdiffusion 1522 -2054 1522 -2054 0 feedthrough
rlabel pdiffusion 1529 -2054 1529 -2054 0 feedthrough
rlabel pdiffusion 1536 -2054 1536 -2054 0 feedthrough
rlabel pdiffusion 1543 -2054 1543 -2054 0 feedthrough
rlabel pdiffusion 1550 -2054 1550 -2054 0 feedthrough
rlabel pdiffusion 1557 -2054 1557 -2054 0 feedthrough
rlabel pdiffusion 1564 -2054 1564 -2054 0 feedthrough
rlabel pdiffusion 1571 -2054 1571 -2054 0 feedthrough
rlabel pdiffusion 1578 -2054 1578 -2054 0 feedthrough
rlabel pdiffusion 1585 -2054 1585 -2054 0 feedthrough
rlabel pdiffusion 1592 -2054 1592 -2054 0 feedthrough
rlabel pdiffusion 1599 -2054 1599 -2054 0 feedthrough
rlabel pdiffusion 1606 -2054 1606 -2054 0 feedthrough
rlabel pdiffusion 1613 -2054 1613 -2054 0 feedthrough
rlabel pdiffusion 1620 -2054 1620 -2054 0 feedthrough
rlabel pdiffusion 1627 -2054 1627 -2054 0 feedthrough
rlabel pdiffusion 1634 -2054 1634 -2054 0 feedthrough
rlabel pdiffusion 1641 -2054 1641 -2054 0 feedthrough
rlabel pdiffusion 1648 -2054 1648 -2054 0 feedthrough
rlabel pdiffusion 1655 -2054 1655 -2054 0 feedthrough
rlabel pdiffusion 1662 -2054 1662 -2054 0 feedthrough
rlabel pdiffusion 1669 -2054 1669 -2054 0 feedthrough
rlabel pdiffusion 1676 -2054 1676 -2054 0 feedthrough
rlabel pdiffusion 1683 -2054 1683 -2054 0 feedthrough
rlabel pdiffusion 1690 -2054 1690 -2054 0 feedthrough
rlabel pdiffusion 1697 -2054 1697 -2054 0 feedthrough
rlabel pdiffusion 1704 -2054 1704 -2054 0 feedthrough
rlabel pdiffusion 1711 -2054 1711 -2054 0 feedthrough
rlabel pdiffusion 1718 -2054 1718 -2054 0 feedthrough
rlabel pdiffusion 1725 -2054 1725 -2054 0 feedthrough
rlabel pdiffusion 1732 -2054 1732 -2054 0 feedthrough
rlabel pdiffusion 1739 -2054 1739 -2054 0 feedthrough
rlabel pdiffusion 1746 -2054 1746 -2054 0 cellNo=533
rlabel pdiffusion 1753 -2054 1753 -2054 0 cellNo=127
rlabel pdiffusion 1760 -2054 1760 -2054 0 cellNo=710
rlabel pdiffusion 1767 -2054 1767 -2054 0 feedthrough
rlabel pdiffusion 1774 -2054 1774 -2054 0 feedthrough
rlabel pdiffusion 3 -2193 3 -2193 0 cellNo=1124
rlabel pdiffusion 10 -2193 10 -2193 0 cellNo=1129
rlabel pdiffusion 17 -2193 17 -2193 0 cellNo=1137
rlabel pdiffusion 24 -2193 24 -2193 0 cellNo=1141
rlabel pdiffusion 31 -2193 31 -2193 0 feedthrough
rlabel pdiffusion 38 -2193 38 -2193 0 cellNo=674
rlabel pdiffusion 45 -2193 45 -2193 0 cellNo=571
rlabel pdiffusion 52 -2193 52 -2193 0 cellNo=542
rlabel pdiffusion 59 -2193 59 -2193 0 feedthrough
rlabel pdiffusion 66 -2193 66 -2193 0 cellNo=9
rlabel pdiffusion 73 -2193 73 -2193 0 feedthrough
rlabel pdiffusion 80 -2193 80 -2193 0 feedthrough
rlabel pdiffusion 87 -2193 87 -2193 0 cellNo=406
rlabel pdiffusion 94 -2193 94 -2193 0 cellNo=194
rlabel pdiffusion 101 -2193 101 -2193 0 feedthrough
rlabel pdiffusion 108 -2193 108 -2193 0 feedthrough
rlabel pdiffusion 115 -2193 115 -2193 0 feedthrough
rlabel pdiffusion 122 -2193 122 -2193 0 feedthrough
rlabel pdiffusion 129 -2193 129 -2193 0 cellNo=650
rlabel pdiffusion 136 -2193 136 -2193 0 feedthrough
rlabel pdiffusion 143 -2193 143 -2193 0 feedthrough
rlabel pdiffusion 150 -2193 150 -2193 0 cellNo=481
rlabel pdiffusion 157 -2193 157 -2193 0 feedthrough
rlabel pdiffusion 164 -2193 164 -2193 0 feedthrough
rlabel pdiffusion 171 -2193 171 -2193 0 cellNo=129
rlabel pdiffusion 178 -2193 178 -2193 0 feedthrough
rlabel pdiffusion 185 -2193 185 -2193 0 feedthrough
rlabel pdiffusion 192 -2193 192 -2193 0 feedthrough
rlabel pdiffusion 199 -2193 199 -2193 0 feedthrough
rlabel pdiffusion 206 -2193 206 -2193 0 feedthrough
rlabel pdiffusion 213 -2193 213 -2193 0 feedthrough
rlabel pdiffusion 220 -2193 220 -2193 0 feedthrough
rlabel pdiffusion 227 -2193 227 -2193 0 cellNo=598
rlabel pdiffusion 234 -2193 234 -2193 0 feedthrough
rlabel pdiffusion 241 -2193 241 -2193 0 feedthrough
rlabel pdiffusion 248 -2193 248 -2193 0 feedthrough
rlabel pdiffusion 255 -2193 255 -2193 0 feedthrough
rlabel pdiffusion 262 -2193 262 -2193 0 feedthrough
rlabel pdiffusion 269 -2193 269 -2193 0 cellNo=547
rlabel pdiffusion 276 -2193 276 -2193 0 feedthrough
rlabel pdiffusion 283 -2193 283 -2193 0 feedthrough
rlabel pdiffusion 290 -2193 290 -2193 0 feedthrough
rlabel pdiffusion 297 -2193 297 -2193 0 feedthrough
rlabel pdiffusion 304 -2193 304 -2193 0 feedthrough
rlabel pdiffusion 311 -2193 311 -2193 0 feedthrough
rlabel pdiffusion 318 -2193 318 -2193 0 feedthrough
rlabel pdiffusion 325 -2193 325 -2193 0 feedthrough
rlabel pdiffusion 332 -2193 332 -2193 0 feedthrough
rlabel pdiffusion 339 -2193 339 -2193 0 feedthrough
rlabel pdiffusion 346 -2193 346 -2193 0 feedthrough
rlabel pdiffusion 353 -2193 353 -2193 0 feedthrough
rlabel pdiffusion 360 -2193 360 -2193 0 cellNo=337
rlabel pdiffusion 367 -2193 367 -2193 0 feedthrough
rlabel pdiffusion 374 -2193 374 -2193 0 feedthrough
rlabel pdiffusion 381 -2193 381 -2193 0 feedthrough
rlabel pdiffusion 388 -2193 388 -2193 0 feedthrough
rlabel pdiffusion 395 -2193 395 -2193 0 feedthrough
rlabel pdiffusion 402 -2193 402 -2193 0 feedthrough
rlabel pdiffusion 409 -2193 409 -2193 0 cellNo=662
rlabel pdiffusion 416 -2193 416 -2193 0 feedthrough
rlabel pdiffusion 423 -2193 423 -2193 0 feedthrough
rlabel pdiffusion 430 -2193 430 -2193 0 feedthrough
rlabel pdiffusion 437 -2193 437 -2193 0 feedthrough
rlabel pdiffusion 444 -2193 444 -2193 0 feedthrough
rlabel pdiffusion 451 -2193 451 -2193 0 cellNo=10
rlabel pdiffusion 458 -2193 458 -2193 0 feedthrough
rlabel pdiffusion 465 -2193 465 -2193 0 feedthrough
rlabel pdiffusion 472 -2193 472 -2193 0 feedthrough
rlabel pdiffusion 479 -2193 479 -2193 0 feedthrough
rlabel pdiffusion 486 -2193 486 -2193 0 feedthrough
rlabel pdiffusion 493 -2193 493 -2193 0 feedthrough
rlabel pdiffusion 500 -2193 500 -2193 0 feedthrough
rlabel pdiffusion 507 -2193 507 -2193 0 feedthrough
rlabel pdiffusion 514 -2193 514 -2193 0 feedthrough
rlabel pdiffusion 521 -2193 521 -2193 0 cellNo=655
rlabel pdiffusion 528 -2193 528 -2193 0 feedthrough
rlabel pdiffusion 535 -2193 535 -2193 0 feedthrough
rlabel pdiffusion 542 -2193 542 -2193 0 feedthrough
rlabel pdiffusion 549 -2193 549 -2193 0 feedthrough
rlabel pdiffusion 556 -2193 556 -2193 0 feedthrough
rlabel pdiffusion 563 -2193 563 -2193 0 feedthrough
rlabel pdiffusion 570 -2193 570 -2193 0 feedthrough
rlabel pdiffusion 577 -2193 577 -2193 0 feedthrough
rlabel pdiffusion 584 -2193 584 -2193 0 feedthrough
rlabel pdiffusion 591 -2193 591 -2193 0 feedthrough
rlabel pdiffusion 598 -2193 598 -2193 0 feedthrough
rlabel pdiffusion 605 -2193 605 -2193 0 cellNo=15
rlabel pdiffusion 612 -2193 612 -2193 0 feedthrough
rlabel pdiffusion 619 -2193 619 -2193 0 cellNo=184
rlabel pdiffusion 626 -2193 626 -2193 0 feedthrough
rlabel pdiffusion 633 -2193 633 -2193 0 feedthrough
rlabel pdiffusion 640 -2193 640 -2193 0 feedthrough
rlabel pdiffusion 647 -2193 647 -2193 0 feedthrough
rlabel pdiffusion 654 -2193 654 -2193 0 feedthrough
rlabel pdiffusion 661 -2193 661 -2193 0 feedthrough
rlabel pdiffusion 668 -2193 668 -2193 0 feedthrough
rlabel pdiffusion 675 -2193 675 -2193 0 feedthrough
rlabel pdiffusion 682 -2193 682 -2193 0 feedthrough
rlabel pdiffusion 689 -2193 689 -2193 0 feedthrough
rlabel pdiffusion 696 -2193 696 -2193 0 feedthrough
rlabel pdiffusion 703 -2193 703 -2193 0 cellNo=799
rlabel pdiffusion 710 -2193 710 -2193 0 feedthrough
rlabel pdiffusion 717 -2193 717 -2193 0 feedthrough
rlabel pdiffusion 724 -2193 724 -2193 0 cellNo=622
rlabel pdiffusion 731 -2193 731 -2193 0 cellNo=554
rlabel pdiffusion 738 -2193 738 -2193 0 feedthrough
rlabel pdiffusion 745 -2193 745 -2193 0 cellNo=171
rlabel pdiffusion 752 -2193 752 -2193 0 feedthrough
rlabel pdiffusion 759 -2193 759 -2193 0 cellNo=540
rlabel pdiffusion 766 -2193 766 -2193 0 feedthrough
rlabel pdiffusion 773 -2193 773 -2193 0 cellNo=857
rlabel pdiffusion 780 -2193 780 -2193 0 feedthrough
rlabel pdiffusion 787 -2193 787 -2193 0 feedthrough
rlabel pdiffusion 794 -2193 794 -2193 0 cellNo=211
rlabel pdiffusion 801 -2193 801 -2193 0 feedthrough
rlabel pdiffusion 808 -2193 808 -2193 0 feedthrough
rlabel pdiffusion 815 -2193 815 -2193 0 cellNo=888
rlabel pdiffusion 822 -2193 822 -2193 0 feedthrough
rlabel pdiffusion 829 -2193 829 -2193 0 cellNo=579
rlabel pdiffusion 836 -2193 836 -2193 0 feedthrough
rlabel pdiffusion 843 -2193 843 -2193 0 feedthrough
rlabel pdiffusion 850 -2193 850 -2193 0 feedthrough
rlabel pdiffusion 857 -2193 857 -2193 0 feedthrough
rlabel pdiffusion 864 -2193 864 -2193 0 feedthrough
rlabel pdiffusion 871 -2193 871 -2193 0 cellNo=61
rlabel pdiffusion 878 -2193 878 -2193 0 feedthrough
rlabel pdiffusion 885 -2193 885 -2193 0 feedthrough
rlabel pdiffusion 892 -2193 892 -2193 0 feedthrough
rlabel pdiffusion 899 -2193 899 -2193 0 feedthrough
rlabel pdiffusion 906 -2193 906 -2193 0 feedthrough
rlabel pdiffusion 913 -2193 913 -2193 0 feedthrough
rlabel pdiffusion 920 -2193 920 -2193 0 feedthrough
rlabel pdiffusion 927 -2193 927 -2193 0 feedthrough
rlabel pdiffusion 934 -2193 934 -2193 0 cellNo=955
rlabel pdiffusion 941 -2193 941 -2193 0 feedthrough
rlabel pdiffusion 948 -2193 948 -2193 0 feedthrough
rlabel pdiffusion 955 -2193 955 -2193 0 feedthrough
rlabel pdiffusion 962 -2193 962 -2193 0 feedthrough
rlabel pdiffusion 969 -2193 969 -2193 0 feedthrough
rlabel pdiffusion 976 -2193 976 -2193 0 cellNo=707
rlabel pdiffusion 983 -2193 983 -2193 0 feedthrough
rlabel pdiffusion 990 -2193 990 -2193 0 feedthrough
rlabel pdiffusion 997 -2193 997 -2193 0 cellNo=473
rlabel pdiffusion 1004 -2193 1004 -2193 0 feedthrough
rlabel pdiffusion 1011 -2193 1011 -2193 0 cellNo=815
rlabel pdiffusion 1018 -2193 1018 -2193 0 feedthrough
rlabel pdiffusion 1025 -2193 1025 -2193 0 feedthrough
rlabel pdiffusion 1032 -2193 1032 -2193 0 feedthrough
rlabel pdiffusion 1039 -2193 1039 -2193 0 feedthrough
rlabel pdiffusion 1046 -2193 1046 -2193 0 feedthrough
rlabel pdiffusion 1053 -2193 1053 -2193 0 feedthrough
rlabel pdiffusion 1060 -2193 1060 -2193 0 feedthrough
rlabel pdiffusion 1067 -2193 1067 -2193 0 feedthrough
rlabel pdiffusion 1074 -2193 1074 -2193 0 feedthrough
rlabel pdiffusion 1081 -2193 1081 -2193 0 feedthrough
rlabel pdiffusion 1088 -2193 1088 -2193 0 feedthrough
rlabel pdiffusion 1095 -2193 1095 -2193 0 feedthrough
rlabel pdiffusion 1102 -2193 1102 -2193 0 cellNo=125
rlabel pdiffusion 1109 -2193 1109 -2193 0 feedthrough
rlabel pdiffusion 1116 -2193 1116 -2193 0 cellNo=404
rlabel pdiffusion 1123 -2193 1123 -2193 0 feedthrough
rlabel pdiffusion 1130 -2193 1130 -2193 0 feedthrough
rlabel pdiffusion 1137 -2193 1137 -2193 0 feedthrough
rlabel pdiffusion 1144 -2193 1144 -2193 0 feedthrough
rlabel pdiffusion 1151 -2193 1151 -2193 0 feedthrough
rlabel pdiffusion 1158 -2193 1158 -2193 0 feedthrough
rlabel pdiffusion 1165 -2193 1165 -2193 0 feedthrough
rlabel pdiffusion 1172 -2193 1172 -2193 0 feedthrough
rlabel pdiffusion 1179 -2193 1179 -2193 0 feedthrough
rlabel pdiffusion 1186 -2193 1186 -2193 0 feedthrough
rlabel pdiffusion 1193 -2193 1193 -2193 0 feedthrough
rlabel pdiffusion 1200 -2193 1200 -2193 0 feedthrough
rlabel pdiffusion 1207 -2193 1207 -2193 0 feedthrough
rlabel pdiffusion 1214 -2193 1214 -2193 0 feedthrough
rlabel pdiffusion 1221 -2193 1221 -2193 0 feedthrough
rlabel pdiffusion 1228 -2193 1228 -2193 0 feedthrough
rlabel pdiffusion 1235 -2193 1235 -2193 0 feedthrough
rlabel pdiffusion 1242 -2193 1242 -2193 0 feedthrough
rlabel pdiffusion 1249 -2193 1249 -2193 0 feedthrough
rlabel pdiffusion 1256 -2193 1256 -2193 0 feedthrough
rlabel pdiffusion 1263 -2193 1263 -2193 0 feedthrough
rlabel pdiffusion 1270 -2193 1270 -2193 0 feedthrough
rlabel pdiffusion 1277 -2193 1277 -2193 0 feedthrough
rlabel pdiffusion 1284 -2193 1284 -2193 0 feedthrough
rlabel pdiffusion 1291 -2193 1291 -2193 0 feedthrough
rlabel pdiffusion 1298 -2193 1298 -2193 0 feedthrough
rlabel pdiffusion 1305 -2193 1305 -2193 0 feedthrough
rlabel pdiffusion 1312 -2193 1312 -2193 0 feedthrough
rlabel pdiffusion 1319 -2193 1319 -2193 0 feedthrough
rlabel pdiffusion 1326 -2193 1326 -2193 0 feedthrough
rlabel pdiffusion 1333 -2193 1333 -2193 0 feedthrough
rlabel pdiffusion 1340 -2193 1340 -2193 0 feedthrough
rlabel pdiffusion 1347 -2193 1347 -2193 0 feedthrough
rlabel pdiffusion 1354 -2193 1354 -2193 0 feedthrough
rlabel pdiffusion 1361 -2193 1361 -2193 0 feedthrough
rlabel pdiffusion 1368 -2193 1368 -2193 0 feedthrough
rlabel pdiffusion 1375 -2193 1375 -2193 0 feedthrough
rlabel pdiffusion 1382 -2193 1382 -2193 0 feedthrough
rlabel pdiffusion 1389 -2193 1389 -2193 0 feedthrough
rlabel pdiffusion 1396 -2193 1396 -2193 0 feedthrough
rlabel pdiffusion 1403 -2193 1403 -2193 0 feedthrough
rlabel pdiffusion 1410 -2193 1410 -2193 0 feedthrough
rlabel pdiffusion 1417 -2193 1417 -2193 0 feedthrough
rlabel pdiffusion 1424 -2193 1424 -2193 0 feedthrough
rlabel pdiffusion 1431 -2193 1431 -2193 0 feedthrough
rlabel pdiffusion 1438 -2193 1438 -2193 0 feedthrough
rlabel pdiffusion 1445 -2193 1445 -2193 0 feedthrough
rlabel pdiffusion 1452 -2193 1452 -2193 0 feedthrough
rlabel pdiffusion 1459 -2193 1459 -2193 0 feedthrough
rlabel pdiffusion 1466 -2193 1466 -2193 0 feedthrough
rlabel pdiffusion 1473 -2193 1473 -2193 0 feedthrough
rlabel pdiffusion 1480 -2193 1480 -2193 0 feedthrough
rlabel pdiffusion 1487 -2193 1487 -2193 0 feedthrough
rlabel pdiffusion 1494 -2193 1494 -2193 0 feedthrough
rlabel pdiffusion 1501 -2193 1501 -2193 0 feedthrough
rlabel pdiffusion 1508 -2193 1508 -2193 0 feedthrough
rlabel pdiffusion 1515 -2193 1515 -2193 0 feedthrough
rlabel pdiffusion 1522 -2193 1522 -2193 0 feedthrough
rlabel pdiffusion 1529 -2193 1529 -2193 0 feedthrough
rlabel pdiffusion 1536 -2193 1536 -2193 0 feedthrough
rlabel pdiffusion 1543 -2193 1543 -2193 0 feedthrough
rlabel pdiffusion 1550 -2193 1550 -2193 0 feedthrough
rlabel pdiffusion 1557 -2193 1557 -2193 0 feedthrough
rlabel pdiffusion 1564 -2193 1564 -2193 0 feedthrough
rlabel pdiffusion 1571 -2193 1571 -2193 0 feedthrough
rlabel pdiffusion 1578 -2193 1578 -2193 0 feedthrough
rlabel pdiffusion 1585 -2193 1585 -2193 0 feedthrough
rlabel pdiffusion 1592 -2193 1592 -2193 0 feedthrough
rlabel pdiffusion 1599 -2193 1599 -2193 0 feedthrough
rlabel pdiffusion 1606 -2193 1606 -2193 0 feedthrough
rlabel pdiffusion 1613 -2193 1613 -2193 0 feedthrough
rlabel pdiffusion 1620 -2193 1620 -2193 0 feedthrough
rlabel pdiffusion 1627 -2193 1627 -2193 0 feedthrough
rlabel pdiffusion 1634 -2193 1634 -2193 0 feedthrough
rlabel pdiffusion 1641 -2193 1641 -2193 0 feedthrough
rlabel pdiffusion 1648 -2193 1648 -2193 0 feedthrough
rlabel pdiffusion 1655 -2193 1655 -2193 0 feedthrough
rlabel pdiffusion 1662 -2193 1662 -2193 0 feedthrough
rlabel pdiffusion 1669 -2193 1669 -2193 0 feedthrough
rlabel pdiffusion 1676 -2193 1676 -2193 0 feedthrough
rlabel pdiffusion 1683 -2193 1683 -2193 0 feedthrough
rlabel pdiffusion 1690 -2193 1690 -2193 0 feedthrough
rlabel pdiffusion 1697 -2193 1697 -2193 0 feedthrough
rlabel pdiffusion 1704 -2193 1704 -2193 0 feedthrough
rlabel pdiffusion 1711 -2193 1711 -2193 0 feedthrough
rlabel pdiffusion 1718 -2193 1718 -2193 0 feedthrough
rlabel pdiffusion 1725 -2193 1725 -2193 0 feedthrough
rlabel pdiffusion 1732 -2193 1732 -2193 0 feedthrough
rlabel pdiffusion 1739 -2193 1739 -2193 0 feedthrough
rlabel pdiffusion 1746 -2193 1746 -2193 0 feedthrough
rlabel pdiffusion 1753 -2193 1753 -2193 0 cellNo=705
rlabel pdiffusion 1760 -2193 1760 -2193 0 feedthrough
rlabel pdiffusion 1767 -2193 1767 -2193 0 feedthrough
rlabel pdiffusion 3 -2328 3 -2328 0 cellNo=1128
rlabel pdiffusion 10 -2328 10 -2328 0 cellNo=1136
rlabel pdiffusion 17 -2328 17 -2328 0 cellNo=1140
rlabel pdiffusion 24 -2328 24 -2328 0 cellNo=1147
rlabel pdiffusion 31 -2328 31 -2328 0 cellNo=1175
rlabel pdiffusion 38 -2328 38 -2328 0 cellNo=1167
rlabel pdiffusion 45 -2328 45 -2328 0 feedthrough
rlabel pdiffusion 52 -2328 52 -2328 0 feedthrough
rlabel pdiffusion 59 -2328 59 -2328 0 feedthrough
rlabel pdiffusion 66 -2328 66 -2328 0 feedthrough
rlabel pdiffusion 73 -2328 73 -2328 0 feedthrough
rlabel pdiffusion 80 -2328 80 -2328 0 feedthrough
rlabel pdiffusion 87 -2328 87 -2328 0 cellNo=62
rlabel pdiffusion 94 -2328 94 -2328 0 cellNo=229
rlabel pdiffusion 101 -2328 101 -2328 0 feedthrough
rlabel pdiffusion 108 -2328 108 -2328 0 feedthrough
rlabel pdiffusion 115 -2328 115 -2328 0 cellNo=494
rlabel pdiffusion 122 -2328 122 -2328 0 feedthrough
rlabel pdiffusion 129 -2328 129 -2328 0 feedthrough
rlabel pdiffusion 136 -2328 136 -2328 0 cellNo=166
rlabel pdiffusion 143 -2328 143 -2328 0 feedthrough
rlabel pdiffusion 150 -2328 150 -2328 0 feedthrough
rlabel pdiffusion 157 -2328 157 -2328 0 feedthrough
rlabel pdiffusion 164 -2328 164 -2328 0 feedthrough
rlabel pdiffusion 171 -2328 171 -2328 0 cellNo=111
rlabel pdiffusion 178 -2328 178 -2328 0 feedthrough
rlabel pdiffusion 185 -2328 185 -2328 0 feedthrough
rlabel pdiffusion 192 -2328 192 -2328 0 feedthrough
rlabel pdiffusion 199 -2328 199 -2328 0 feedthrough
rlabel pdiffusion 206 -2328 206 -2328 0 feedthrough
rlabel pdiffusion 213 -2328 213 -2328 0 cellNo=386
rlabel pdiffusion 220 -2328 220 -2328 0 feedthrough
rlabel pdiffusion 227 -2328 227 -2328 0 feedthrough
rlabel pdiffusion 234 -2328 234 -2328 0 cellNo=629
rlabel pdiffusion 241 -2328 241 -2328 0 feedthrough
rlabel pdiffusion 248 -2328 248 -2328 0 feedthrough
rlabel pdiffusion 255 -2328 255 -2328 0 feedthrough
rlabel pdiffusion 262 -2328 262 -2328 0 feedthrough
rlabel pdiffusion 269 -2328 269 -2328 0 feedthrough
rlabel pdiffusion 276 -2328 276 -2328 0 feedthrough
rlabel pdiffusion 283 -2328 283 -2328 0 feedthrough
rlabel pdiffusion 290 -2328 290 -2328 0 feedthrough
rlabel pdiffusion 297 -2328 297 -2328 0 feedthrough
rlabel pdiffusion 304 -2328 304 -2328 0 feedthrough
rlabel pdiffusion 311 -2328 311 -2328 0 feedthrough
rlabel pdiffusion 318 -2328 318 -2328 0 feedthrough
rlabel pdiffusion 325 -2328 325 -2328 0 feedthrough
rlabel pdiffusion 332 -2328 332 -2328 0 feedthrough
rlabel pdiffusion 339 -2328 339 -2328 0 feedthrough
rlabel pdiffusion 346 -2328 346 -2328 0 feedthrough
rlabel pdiffusion 353 -2328 353 -2328 0 feedthrough
rlabel pdiffusion 360 -2328 360 -2328 0 feedthrough
rlabel pdiffusion 367 -2328 367 -2328 0 feedthrough
rlabel pdiffusion 374 -2328 374 -2328 0 feedthrough
rlabel pdiffusion 381 -2328 381 -2328 0 feedthrough
rlabel pdiffusion 388 -2328 388 -2328 0 feedthrough
rlabel pdiffusion 395 -2328 395 -2328 0 feedthrough
rlabel pdiffusion 402 -2328 402 -2328 0 feedthrough
rlabel pdiffusion 409 -2328 409 -2328 0 feedthrough
rlabel pdiffusion 416 -2328 416 -2328 0 feedthrough
rlabel pdiffusion 423 -2328 423 -2328 0 feedthrough
rlabel pdiffusion 430 -2328 430 -2328 0 feedthrough
rlabel pdiffusion 437 -2328 437 -2328 0 feedthrough
rlabel pdiffusion 444 -2328 444 -2328 0 feedthrough
rlabel pdiffusion 451 -2328 451 -2328 0 feedthrough
rlabel pdiffusion 458 -2328 458 -2328 0 feedthrough
rlabel pdiffusion 465 -2328 465 -2328 0 feedthrough
rlabel pdiffusion 472 -2328 472 -2328 0 feedthrough
rlabel pdiffusion 479 -2328 479 -2328 0 feedthrough
rlabel pdiffusion 486 -2328 486 -2328 0 feedthrough
rlabel pdiffusion 493 -2328 493 -2328 0 feedthrough
rlabel pdiffusion 500 -2328 500 -2328 0 feedthrough
rlabel pdiffusion 507 -2328 507 -2328 0 feedthrough
rlabel pdiffusion 514 -2328 514 -2328 0 feedthrough
rlabel pdiffusion 521 -2328 521 -2328 0 feedthrough
rlabel pdiffusion 528 -2328 528 -2328 0 feedthrough
rlabel pdiffusion 535 -2328 535 -2328 0 cellNo=38
rlabel pdiffusion 542 -2328 542 -2328 0 feedthrough
rlabel pdiffusion 549 -2328 549 -2328 0 feedthrough
rlabel pdiffusion 556 -2328 556 -2328 0 feedthrough
rlabel pdiffusion 563 -2328 563 -2328 0 feedthrough
rlabel pdiffusion 570 -2328 570 -2328 0 feedthrough
rlabel pdiffusion 577 -2328 577 -2328 0 feedthrough
rlabel pdiffusion 584 -2328 584 -2328 0 cellNo=854
rlabel pdiffusion 591 -2328 591 -2328 0 feedthrough
rlabel pdiffusion 598 -2328 598 -2328 0 feedthrough
rlabel pdiffusion 605 -2328 605 -2328 0 feedthrough
rlabel pdiffusion 612 -2328 612 -2328 0 feedthrough
rlabel pdiffusion 619 -2328 619 -2328 0 feedthrough
rlabel pdiffusion 626 -2328 626 -2328 0 feedthrough
rlabel pdiffusion 633 -2328 633 -2328 0 feedthrough
rlabel pdiffusion 640 -2328 640 -2328 0 cellNo=847
rlabel pdiffusion 647 -2328 647 -2328 0 feedthrough
rlabel pdiffusion 654 -2328 654 -2328 0 cellNo=577
rlabel pdiffusion 661 -2328 661 -2328 0 feedthrough
rlabel pdiffusion 668 -2328 668 -2328 0 feedthrough
rlabel pdiffusion 675 -2328 675 -2328 0 feedthrough
rlabel pdiffusion 682 -2328 682 -2328 0 feedthrough
rlabel pdiffusion 689 -2328 689 -2328 0 cellNo=454
rlabel pdiffusion 696 -2328 696 -2328 0 feedthrough
rlabel pdiffusion 703 -2328 703 -2328 0 cellNo=299
rlabel pdiffusion 710 -2328 710 -2328 0 feedthrough
rlabel pdiffusion 717 -2328 717 -2328 0 feedthrough
rlabel pdiffusion 724 -2328 724 -2328 0 feedthrough
rlabel pdiffusion 731 -2328 731 -2328 0 cellNo=589
rlabel pdiffusion 738 -2328 738 -2328 0 feedthrough
rlabel pdiffusion 745 -2328 745 -2328 0 cellNo=975
rlabel pdiffusion 752 -2328 752 -2328 0 feedthrough
rlabel pdiffusion 759 -2328 759 -2328 0 feedthrough
rlabel pdiffusion 766 -2328 766 -2328 0 feedthrough
rlabel pdiffusion 773 -2328 773 -2328 0 cellNo=487
rlabel pdiffusion 780 -2328 780 -2328 0 feedthrough
rlabel pdiffusion 787 -2328 787 -2328 0 feedthrough
rlabel pdiffusion 794 -2328 794 -2328 0 feedthrough
rlabel pdiffusion 801 -2328 801 -2328 0 feedthrough
rlabel pdiffusion 808 -2328 808 -2328 0 feedthrough
rlabel pdiffusion 815 -2328 815 -2328 0 feedthrough
rlabel pdiffusion 822 -2328 822 -2328 0 feedthrough
rlabel pdiffusion 829 -2328 829 -2328 0 feedthrough
rlabel pdiffusion 836 -2328 836 -2328 0 feedthrough
rlabel pdiffusion 843 -2328 843 -2328 0 feedthrough
rlabel pdiffusion 850 -2328 850 -2328 0 cellNo=262
rlabel pdiffusion 857 -2328 857 -2328 0 feedthrough
rlabel pdiffusion 864 -2328 864 -2328 0 feedthrough
rlabel pdiffusion 871 -2328 871 -2328 0 cellNo=997
rlabel pdiffusion 878 -2328 878 -2328 0 feedthrough
rlabel pdiffusion 885 -2328 885 -2328 0 feedthrough
rlabel pdiffusion 892 -2328 892 -2328 0 feedthrough
rlabel pdiffusion 899 -2328 899 -2328 0 cellNo=924
rlabel pdiffusion 906 -2328 906 -2328 0 feedthrough
rlabel pdiffusion 913 -2328 913 -2328 0 feedthrough
rlabel pdiffusion 920 -2328 920 -2328 0 feedthrough
rlabel pdiffusion 927 -2328 927 -2328 0 feedthrough
rlabel pdiffusion 934 -2328 934 -2328 0 feedthrough
rlabel pdiffusion 941 -2328 941 -2328 0 feedthrough
rlabel pdiffusion 948 -2328 948 -2328 0 feedthrough
rlabel pdiffusion 955 -2328 955 -2328 0 cellNo=981
rlabel pdiffusion 962 -2328 962 -2328 0 feedthrough
rlabel pdiffusion 969 -2328 969 -2328 0 cellNo=232
rlabel pdiffusion 976 -2328 976 -2328 0 feedthrough
rlabel pdiffusion 983 -2328 983 -2328 0 feedthrough
rlabel pdiffusion 990 -2328 990 -2328 0 feedthrough
rlabel pdiffusion 997 -2328 997 -2328 0 cellNo=937
rlabel pdiffusion 1004 -2328 1004 -2328 0 feedthrough
rlabel pdiffusion 1011 -2328 1011 -2328 0 feedthrough
rlabel pdiffusion 1018 -2328 1018 -2328 0 feedthrough
rlabel pdiffusion 1025 -2328 1025 -2328 0 feedthrough
rlabel pdiffusion 1032 -2328 1032 -2328 0 feedthrough
rlabel pdiffusion 1039 -2328 1039 -2328 0 feedthrough
rlabel pdiffusion 1046 -2328 1046 -2328 0 feedthrough
rlabel pdiffusion 1053 -2328 1053 -2328 0 feedthrough
rlabel pdiffusion 1060 -2328 1060 -2328 0 feedthrough
rlabel pdiffusion 1067 -2328 1067 -2328 0 feedthrough
rlabel pdiffusion 1074 -2328 1074 -2328 0 feedthrough
rlabel pdiffusion 1081 -2328 1081 -2328 0 cellNo=918
rlabel pdiffusion 1088 -2328 1088 -2328 0 feedthrough
rlabel pdiffusion 1095 -2328 1095 -2328 0 cellNo=917
rlabel pdiffusion 1102 -2328 1102 -2328 0 feedthrough
rlabel pdiffusion 1109 -2328 1109 -2328 0 feedthrough
rlabel pdiffusion 1116 -2328 1116 -2328 0 feedthrough
rlabel pdiffusion 1123 -2328 1123 -2328 0 cellNo=302
rlabel pdiffusion 1130 -2328 1130 -2328 0 feedthrough
rlabel pdiffusion 1137 -2328 1137 -2328 0 feedthrough
rlabel pdiffusion 1144 -2328 1144 -2328 0 cellNo=138
rlabel pdiffusion 1151 -2328 1151 -2328 0 feedthrough
rlabel pdiffusion 1158 -2328 1158 -2328 0 feedthrough
rlabel pdiffusion 1165 -2328 1165 -2328 0 feedthrough
rlabel pdiffusion 1172 -2328 1172 -2328 0 cellNo=288
rlabel pdiffusion 1179 -2328 1179 -2328 0 feedthrough
rlabel pdiffusion 1186 -2328 1186 -2328 0 feedthrough
rlabel pdiffusion 1193 -2328 1193 -2328 0 feedthrough
rlabel pdiffusion 1200 -2328 1200 -2328 0 feedthrough
rlabel pdiffusion 1207 -2328 1207 -2328 0 feedthrough
rlabel pdiffusion 1214 -2328 1214 -2328 0 feedthrough
rlabel pdiffusion 1221 -2328 1221 -2328 0 feedthrough
rlabel pdiffusion 1228 -2328 1228 -2328 0 feedthrough
rlabel pdiffusion 1235 -2328 1235 -2328 0 cellNo=209
rlabel pdiffusion 1242 -2328 1242 -2328 0 feedthrough
rlabel pdiffusion 1249 -2328 1249 -2328 0 feedthrough
rlabel pdiffusion 1256 -2328 1256 -2328 0 feedthrough
rlabel pdiffusion 1263 -2328 1263 -2328 0 feedthrough
rlabel pdiffusion 1270 -2328 1270 -2328 0 feedthrough
rlabel pdiffusion 1277 -2328 1277 -2328 0 feedthrough
rlabel pdiffusion 1284 -2328 1284 -2328 0 feedthrough
rlabel pdiffusion 1291 -2328 1291 -2328 0 feedthrough
rlabel pdiffusion 1298 -2328 1298 -2328 0 feedthrough
rlabel pdiffusion 1305 -2328 1305 -2328 0 cellNo=130
rlabel pdiffusion 1312 -2328 1312 -2328 0 feedthrough
rlabel pdiffusion 1319 -2328 1319 -2328 0 feedthrough
rlabel pdiffusion 1326 -2328 1326 -2328 0 feedthrough
rlabel pdiffusion 1333 -2328 1333 -2328 0 cellNo=382
rlabel pdiffusion 1340 -2328 1340 -2328 0 feedthrough
rlabel pdiffusion 1347 -2328 1347 -2328 0 feedthrough
rlabel pdiffusion 1354 -2328 1354 -2328 0 feedthrough
rlabel pdiffusion 1361 -2328 1361 -2328 0 feedthrough
rlabel pdiffusion 1368 -2328 1368 -2328 0 feedthrough
rlabel pdiffusion 1375 -2328 1375 -2328 0 feedthrough
rlabel pdiffusion 1382 -2328 1382 -2328 0 feedthrough
rlabel pdiffusion 1389 -2328 1389 -2328 0 feedthrough
rlabel pdiffusion 1396 -2328 1396 -2328 0 feedthrough
rlabel pdiffusion 1403 -2328 1403 -2328 0 feedthrough
rlabel pdiffusion 1410 -2328 1410 -2328 0 feedthrough
rlabel pdiffusion 1417 -2328 1417 -2328 0 feedthrough
rlabel pdiffusion 1424 -2328 1424 -2328 0 feedthrough
rlabel pdiffusion 1431 -2328 1431 -2328 0 feedthrough
rlabel pdiffusion 1438 -2328 1438 -2328 0 feedthrough
rlabel pdiffusion 1445 -2328 1445 -2328 0 feedthrough
rlabel pdiffusion 1452 -2328 1452 -2328 0 feedthrough
rlabel pdiffusion 1459 -2328 1459 -2328 0 feedthrough
rlabel pdiffusion 1466 -2328 1466 -2328 0 feedthrough
rlabel pdiffusion 1473 -2328 1473 -2328 0 feedthrough
rlabel pdiffusion 1480 -2328 1480 -2328 0 feedthrough
rlabel pdiffusion 1487 -2328 1487 -2328 0 feedthrough
rlabel pdiffusion 1494 -2328 1494 -2328 0 feedthrough
rlabel pdiffusion 1501 -2328 1501 -2328 0 feedthrough
rlabel pdiffusion 1508 -2328 1508 -2328 0 feedthrough
rlabel pdiffusion 1515 -2328 1515 -2328 0 feedthrough
rlabel pdiffusion 1522 -2328 1522 -2328 0 feedthrough
rlabel pdiffusion 1529 -2328 1529 -2328 0 feedthrough
rlabel pdiffusion 1536 -2328 1536 -2328 0 feedthrough
rlabel pdiffusion 1543 -2328 1543 -2328 0 feedthrough
rlabel pdiffusion 1550 -2328 1550 -2328 0 feedthrough
rlabel pdiffusion 1557 -2328 1557 -2328 0 feedthrough
rlabel pdiffusion 1564 -2328 1564 -2328 0 feedthrough
rlabel pdiffusion 1571 -2328 1571 -2328 0 feedthrough
rlabel pdiffusion 1578 -2328 1578 -2328 0 feedthrough
rlabel pdiffusion 1585 -2328 1585 -2328 0 feedthrough
rlabel pdiffusion 1592 -2328 1592 -2328 0 feedthrough
rlabel pdiffusion 1599 -2328 1599 -2328 0 feedthrough
rlabel pdiffusion 1606 -2328 1606 -2328 0 feedthrough
rlabel pdiffusion 1613 -2328 1613 -2328 0 feedthrough
rlabel pdiffusion 1620 -2328 1620 -2328 0 feedthrough
rlabel pdiffusion 1627 -2328 1627 -2328 0 feedthrough
rlabel pdiffusion 1634 -2328 1634 -2328 0 feedthrough
rlabel pdiffusion 1641 -2328 1641 -2328 0 feedthrough
rlabel pdiffusion 1648 -2328 1648 -2328 0 feedthrough
rlabel pdiffusion 1655 -2328 1655 -2328 0 feedthrough
rlabel pdiffusion 1662 -2328 1662 -2328 0 feedthrough
rlabel pdiffusion 1669 -2328 1669 -2328 0 feedthrough
rlabel pdiffusion 1676 -2328 1676 -2328 0 feedthrough
rlabel pdiffusion 1683 -2328 1683 -2328 0 feedthrough
rlabel pdiffusion 1690 -2328 1690 -2328 0 feedthrough
rlabel pdiffusion 1697 -2328 1697 -2328 0 feedthrough
rlabel pdiffusion 1704 -2328 1704 -2328 0 cellNo=640
rlabel pdiffusion 1711 -2328 1711 -2328 0 cellNo=644
rlabel pdiffusion 1718 -2328 1718 -2328 0 feedthrough
rlabel pdiffusion 1725 -2328 1725 -2328 0 feedthrough
rlabel pdiffusion 1732 -2328 1732 -2328 0 feedthrough
rlabel pdiffusion 1739 -2328 1739 -2328 0 feedthrough
rlabel pdiffusion 3 -2443 3 -2443 0 cellNo=1135
rlabel pdiffusion 10 -2443 10 -2443 0 cellNo=1139
rlabel pdiffusion 17 -2443 17 -2443 0 cellNo=1146
rlabel pdiffusion 24 -2443 24 -2443 0 cellNo=1153
rlabel pdiffusion 31 -2443 31 -2443 0 cellNo=1165
rlabel pdiffusion 52 -2443 52 -2443 0 feedthrough
rlabel pdiffusion 59 -2443 59 -2443 0 feedthrough
rlabel pdiffusion 66 -2443 66 -2443 0 feedthrough
rlabel pdiffusion 73 -2443 73 -2443 0 feedthrough
rlabel pdiffusion 80 -2443 80 -2443 0 feedthrough
rlabel pdiffusion 87 -2443 87 -2443 0 feedthrough
rlabel pdiffusion 94 -2443 94 -2443 0 feedthrough
rlabel pdiffusion 101 -2443 101 -2443 0 feedthrough
rlabel pdiffusion 108 -2443 108 -2443 0 feedthrough
rlabel pdiffusion 115 -2443 115 -2443 0 feedthrough
rlabel pdiffusion 122 -2443 122 -2443 0 feedthrough
rlabel pdiffusion 129 -2443 129 -2443 0 feedthrough
rlabel pdiffusion 136 -2443 136 -2443 0 feedthrough
rlabel pdiffusion 143 -2443 143 -2443 0 feedthrough
rlabel pdiffusion 150 -2443 150 -2443 0 feedthrough
rlabel pdiffusion 157 -2443 157 -2443 0 feedthrough
rlabel pdiffusion 164 -2443 164 -2443 0 feedthrough
rlabel pdiffusion 171 -2443 171 -2443 0 feedthrough
rlabel pdiffusion 178 -2443 178 -2443 0 cellNo=292
rlabel pdiffusion 185 -2443 185 -2443 0 feedthrough
rlabel pdiffusion 192 -2443 192 -2443 0 feedthrough
rlabel pdiffusion 199 -2443 199 -2443 0 feedthrough
rlabel pdiffusion 206 -2443 206 -2443 0 feedthrough
rlabel pdiffusion 213 -2443 213 -2443 0 cellNo=570
rlabel pdiffusion 220 -2443 220 -2443 0 feedthrough
rlabel pdiffusion 227 -2443 227 -2443 0 feedthrough
rlabel pdiffusion 234 -2443 234 -2443 0 feedthrough
rlabel pdiffusion 241 -2443 241 -2443 0 feedthrough
rlabel pdiffusion 248 -2443 248 -2443 0 feedthrough
rlabel pdiffusion 255 -2443 255 -2443 0 cellNo=945
rlabel pdiffusion 262 -2443 262 -2443 0 feedthrough
rlabel pdiffusion 269 -2443 269 -2443 0 feedthrough
rlabel pdiffusion 276 -2443 276 -2443 0 feedthrough
rlabel pdiffusion 283 -2443 283 -2443 0 feedthrough
rlabel pdiffusion 290 -2443 290 -2443 0 feedthrough
rlabel pdiffusion 297 -2443 297 -2443 0 feedthrough
rlabel pdiffusion 304 -2443 304 -2443 0 feedthrough
rlabel pdiffusion 311 -2443 311 -2443 0 cellNo=154
rlabel pdiffusion 318 -2443 318 -2443 0 feedthrough
rlabel pdiffusion 325 -2443 325 -2443 0 feedthrough
rlabel pdiffusion 332 -2443 332 -2443 0 feedthrough
rlabel pdiffusion 339 -2443 339 -2443 0 feedthrough
rlabel pdiffusion 346 -2443 346 -2443 0 feedthrough
rlabel pdiffusion 353 -2443 353 -2443 0 feedthrough
rlabel pdiffusion 360 -2443 360 -2443 0 feedthrough
rlabel pdiffusion 367 -2443 367 -2443 0 feedthrough
rlabel pdiffusion 374 -2443 374 -2443 0 feedthrough
rlabel pdiffusion 381 -2443 381 -2443 0 feedthrough
rlabel pdiffusion 388 -2443 388 -2443 0 feedthrough
rlabel pdiffusion 395 -2443 395 -2443 0 feedthrough
rlabel pdiffusion 402 -2443 402 -2443 0 feedthrough
rlabel pdiffusion 409 -2443 409 -2443 0 feedthrough
rlabel pdiffusion 416 -2443 416 -2443 0 feedthrough
rlabel pdiffusion 423 -2443 423 -2443 0 feedthrough
rlabel pdiffusion 430 -2443 430 -2443 0 cellNo=907
rlabel pdiffusion 437 -2443 437 -2443 0 feedthrough
rlabel pdiffusion 444 -2443 444 -2443 0 feedthrough
rlabel pdiffusion 451 -2443 451 -2443 0 feedthrough
rlabel pdiffusion 458 -2443 458 -2443 0 feedthrough
rlabel pdiffusion 465 -2443 465 -2443 0 feedthrough
rlabel pdiffusion 472 -2443 472 -2443 0 cellNo=925
rlabel pdiffusion 479 -2443 479 -2443 0 feedthrough
rlabel pdiffusion 486 -2443 486 -2443 0 feedthrough
rlabel pdiffusion 493 -2443 493 -2443 0 feedthrough
rlabel pdiffusion 500 -2443 500 -2443 0 cellNo=308
rlabel pdiffusion 507 -2443 507 -2443 0 feedthrough
rlabel pdiffusion 514 -2443 514 -2443 0 feedthrough
rlabel pdiffusion 521 -2443 521 -2443 0 feedthrough
rlabel pdiffusion 528 -2443 528 -2443 0 cellNo=941
rlabel pdiffusion 535 -2443 535 -2443 0 feedthrough
rlabel pdiffusion 542 -2443 542 -2443 0 cellNo=2
rlabel pdiffusion 549 -2443 549 -2443 0 feedthrough
rlabel pdiffusion 556 -2443 556 -2443 0 feedthrough
rlabel pdiffusion 563 -2443 563 -2443 0 feedthrough
rlabel pdiffusion 570 -2443 570 -2443 0 feedthrough
rlabel pdiffusion 577 -2443 577 -2443 0 feedthrough
rlabel pdiffusion 584 -2443 584 -2443 0 feedthrough
rlabel pdiffusion 591 -2443 591 -2443 0 feedthrough
rlabel pdiffusion 598 -2443 598 -2443 0 feedthrough
rlabel pdiffusion 605 -2443 605 -2443 0 feedthrough
rlabel pdiffusion 612 -2443 612 -2443 0 cellNo=686
rlabel pdiffusion 619 -2443 619 -2443 0 feedthrough
rlabel pdiffusion 626 -2443 626 -2443 0 feedthrough
rlabel pdiffusion 633 -2443 633 -2443 0 feedthrough
rlabel pdiffusion 640 -2443 640 -2443 0 cellNo=150
rlabel pdiffusion 647 -2443 647 -2443 0 feedthrough
rlabel pdiffusion 654 -2443 654 -2443 0 feedthrough
rlabel pdiffusion 661 -2443 661 -2443 0 feedthrough
rlabel pdiffusion 668 -2443 668 -2443 0 feedthrough
rlabel pdiffusion 675 -2443 675 -2443 0 cellNo=464
rlabel pdiffusion 682 -2443 682 -2443 0 cellNo=95
rlabel pdiffusion 689 -2443 689 -2443 0 feedthrough
rlabel pdiffusion 696 -2443 696 -2443 0 feedthrough
rlabel pdiffusion 703 -2443 703 -2443 0 cellNo=276
rlabel pdiffusion 710 -2443 710 -2443 0 feedthrough
rlabel pdiffusion 717 -2443 717 -2443 0 feedthrough
rlabel pdiffusion 724 -2443 724 -2443 0 feedthrough
rlabel pdiffusion 731 -2443 731 -2443 0 cellNo=1
rlabel pdiffusion 738 -2443 738 -2443 0 feedthrough
rlabel pdiffusion 745 -2443 745 -2443 0 cellNo=343
rlabel pdiffusion 752 -2443 752 -2443 0 feedthrough
rlabel pdiffusion 759 -2443 759 -2443 0 feedthrough
rlabel pdiffusion 766 -2443 766 -2443 0 feedthrough
rlabel pdiffusion 773 -2443 773 -2443 0 feedthrough
rlabel pdiffusion 780 -2443 780 -2443 0 feedthrough
rlabel pdiffusion 787 -2443 787 -2443 0 feedthrough
rlabel pdiffusion 794 -2443 794 -2443 0 feedthrough
rlabel pdiffusion 801 -2443 801 -2443 0 feedthrough
rlabel pdiffusion 808 -2443 808 -2443 0 cellNo=552
rlabel pdiffusion 815 -2443 815 -2443 0 feedthrough
rlabel pdiffusion 822 -2443 822 -2443 0 cellNo=724
rlabel pdiffusion 829 -2443 829 -2443 0 feedthrough
rlabel pdiffusion 836 -2443 836 -2443 0 feedthrough
rlabel pdiffusion 843 -2443 843 -2443 0 cellNo=606
rlabel pdiffusion 850 -2443 850 -2443 0 cellNo=202
rlabel pdiffusion 857 -2443 857 -2443 0 cellNo=119
rlabel pdiffusion 864 -2443 864 -2443 0 feedthrough
rlabel pdiffusion 871 -2443 871 -2443 0 feedthrough
rlabel pdiffusion 878 -2443 878 -2443 0 feedthrough
rlabel pdiffusion 885 -2443 885 -2443 0 feedthrough
rlabel pdiffusion 892 -2443 892 -2443 0 cellNo=264
rlabel pdiffusion 899 -2443 899 -2443 0 cellNo=809
rlabel pdiffusion 906 -2443 906 -2443 0 feedthrough
rlabel pdiffusion 913 -2443 913 -2443 0 feedthrough
rlabel pdiffusion 920 -2443 920 -2443 0 feedthrough
rlabel pdiffusion 927 -2443 927 -2443 0 feedthrough
rlabel pdiffusion 934 -2443 934 -2443 0 feedthrough
rlabel pdiffusion 941 -2443 941 -2443 0 feedthrough
rlabel pdiffusion 948 -2443 948 -2443 0 feedthrough
rlabel pdiffusion 955 -2443 955 -2443 0 feedthrough
rlabel pdiffusion 962 -2443 962 -2443 0 feedthrough
rlabel pdiffusion 969 -2443 969 -2443 0 cellNo=20
rlabel pdiffusion 976 -2443 976 -2443 0 feedthrough
rlabel pdiffusion 983 -2443 983 -2443 0 feedthrough
rlabel pdiffusion 990 -2443 990 -2443 0 feedthrough
rlabel pdiffusion 997 -2443 997 -2443 0 feedthrough
rlabel pdiffusion 1004 -2443 1004 -2443 0 feedthrough
rlabel pdiffusion 1011 -2443 1011 -2443 0 feedthrough
rlabel pdiffusion 1018 -2443 1018 -2443 0 feedthrough
rlabel pdiffusion 1025 -2443 1025 -2443 0 feedthrough
rlabel pdiffusion 1032 -2443 1032 -2443 0 feedthrough
rlabel pdiffusion 1039 -2443 1039 -2443 0 feedthrough
rlabel pdiffusion 1046 -2443 1046 -2443 0 feedthrough
rlabel pdiffusion 1053 -2443 1053 -2443 0 feedthrough
rlabel pdiffusion 1060 -2443 1060 -2443 0 feedthrough
rlabel pdiffusion 1067 -2443 1067 -2443 0 feedthrough
rlabel pdiffusion 1074 -2443 1074 -2443 0 cellNo=175
rlabel pdiffusion 1081 -2443 1081 -2443 0 feedthrough
rlabel pdiffusion 1088 -2443 1088 -2443 0 feedthrough
rlabel pdiffusion 1095 -2443 1095 -2443 0 feedthrough
rlabel pdiffusion 1102 -2443 1102 -2443 0 feedthrough
rlabel pdiffusion 1109 -2443 1109 -2443 0 feedthrough
rlabel pdiffusion 1116 -2443 1116 -2443 0 feedthrough
rlabel pdiffusion 1123 -2443 1123 -2443 0 feedthrough
rlabel pdiffusion 1130 -2443 1130 -2443 0 feedthrough
rlabel pdiffusion 1137 -2443 1137 -2443 0 feedthrough
rlabel pdiffusion 1144 -2443 1144 -2443 0 feedthrough
rlabel pdiffusion 1151 -2443 1151 -2443 0 feedthrough
rlabel pdiffusion 1158 -2443 1158 -2443 0 feedthrough
rlabel pdiffusion 1165 -2443 1165 -2443 0 feedthrough
rlabel pdiffusion 1172 -2443 1172 -2443 0 feedthrough
rlabel pdiffusion 1179 -2443 1179 -2443 0 feedthrough
rlabel pdiffusion 1186 -2443 1186 -2443 0 feedthrough
rlabel pdiffusion 1193 -2443 1193 -2443 0 cellNo=115
rlabel pdiffusion 1200 -2443 1200 -2443 0 feedthrough
rlabel pdiffusion 1207 -2443 1207 -2443 0 cellNo=561
rlabel pdiffusion 1214 -2443 1214 -2443 0 feedthrough
rlabel pdiffusion 1221 -2443 1221 -2443 0 feedthrough
rlabel pdiffusion 1228 -2443 1228 -2443 0 feedthrough
rlabel pdiffusion 1235 -2443 1235 -2443 0 feedthrough
rlabel pdiffusion 1242 -2443 1242 -2443 0 cellNo=979
rlabel pdiffusion 1249 -2443 1249 -2443 0 feedthrough
rlabel pdiffusion 1256 -2443 1256 -2443 0 feedthrough
rlabel pdiffusion 1263 -2443 1263 -2443 0 feedthrough
rlabel pdiffusion 1270 -2443 1270 -2443 0 feedthrough
rlabel pdiffusion 1277 -2443 1277 -2443 0 feedthrough
rlabel pdiffusion 1284 -2443 1284 -2443 0 feedthrough
rlabel pdiffusion 1291 -2443 1291 -2443 0 feedthrough
rlabel pdiffusion 1298 -2443 1298 -2443 0 cellNo=609
rlabel pdiffusion 1305 -2443 1305 -2443 0 feedthrough
rlabel pdiffusion 1312 -2443 1312 -2443 0 cellNo=373
rlabel pdiffusion 1319 -2443 1319 -2443 0 feedthrough
rlabel pdiffusion 1326 -2443 1326 -2443 0 feedthrough
rlabel pdiffusion 1333 -2443 1333 -2443 0 feedthrough
rlabel pdiffusion 1340 -2443 1340 -2443 0 feedthrough
rlabel pdiffusion 1347 -2443 1347 -2443 0 feedthrough
rlabel pdiffusion 1354 -2443 1354 -2443 0 feedthrough
rlabel pdiffusion 1361 -2443 1361 -2443 0 feedthrough
rlabel pdiffusion 1368 -2443 1368 -2443 0 feedthrough
rlabel pdiffusion 1375 -2443 1375 -2443 0 feedthrough
rlabel pdiffusion 1382 -2443 1382 -2443 0 cellNo=933
rlabel pdiffusion 1389 -2443 1389 -2443 0 feedthrough
rlabel pdiffusion 1396 -2443 1396 -2443 0 feedthrough
rlabel pdiffusion 1403 -2443 1403 -2443 0 feedthrough
rlabel pdiffusion 1410 -2443 1410 -2443 0 feedthrough
rlabel pdiffusion 1417 -2443 1417 -2443 0 feedthrough
rlabel pdiffusion 1424 -2443 1424 -2443 0 feedthrough
rlabel pdiffusion 1431 -2443 1431 -2443 0 feedthrough
rlabel pdiffusion 1438 -2443 1438 -2443 0 feedthrough
rlabel pdiffusion 1445 -2443 1445 -2443 0 feedthrough
rlabel pdiffusion 1452 -2443 1452 -2443 0 feedthrough
rlabel pdiffusion 1459 -2443 1459 -2443 0 feedthrough
rlabel pdiffusion 1466 -2443 1466 -2443 0 feedthrough
rlabel pdiffusion 1473 -2443 1473 -2443 0 feedthrough
rlabel pdiffusion 1480 -2443 1480 -2443 0 feedthrough
rlabel pdiffusion 1487 -2443 1487 -2443 0 feedthrough
rlabel pdiffusion 1494 -2443 1494 -2443 0 feedthrough
rlabel pdiffusion 1501 -2443 1501 -2443 0 feedthrough
rlabel pdiffusion 1508 -2443 1508 -2443 0 feedthrough
rlabel pdiffusion 1515 -2443 1515 -2443 0 feedthrough
rlabel pdiffusion 1522 -2443 1522 -2443 0 feedthrough
rlabel pdiffusion 1529 -2443 1529 -2443 0 feedthrough
rlabel pdiffusion 1536 -2443 1536 -2443 0 cellNo=80
rlabel pdiffusion 1543 -2443 1543 -2443 0 feedthrough
rlabel pdiffusion 1550 -2443 1550 -2443 0 feedthrough
rlabel pdiffusion 1557 -2443 1557 -2443 0 feedthrough
rlabel pdiffusion 1564 -2443 1564 -2443 0 feedthrough
rlabel pdiffusion 1571 -2443 1571 -2443 0 feedthrough
rlabel pdiffusion 1578 -2443 1578 -2443 0 cellNo=527
rlabel pdiffusion 1585 -2443 1585 -2443 0 feedthrough
rlabel pdiffusion 1592 -2443 1592 -2443 0 feedthrough
rlabel pdiffusion 1599 -2443 1599 -2443 0 feedthrough
rlabel pdiffusion 1606 -2443 1606 -2443 0 feedthrough
rlabel pdiffusion 1676 -2443 1676 -2443 0 feedthrough
rlabel pdiffusion 3 -2560 3 -2560 0 cellNo=1138
rlabel pdiffusion 10 -2560 10 -2560 0 cellNo=1145
rlabel pdiffusion 17 -2560 17 -2560 0 cellNo=1152
rlabel pdiffusion 24 -2560 24 -2560 0 cellNo=1163
rlabel pdiffusion 31 -2560 31 -2560 0 cellNo=1177
rlabel pdiffusion 38 -2560 38 -2560 0 cellNo=1186
rlabel pdiffusion 45 -2560 45 -2560 0 feedthrough
rlabel pdiffusion 52 -2560 52 -2560 0 feedthrough
rlabel pdiffusion 59 -2560 59 -2560 0 feedthrough
rlabel pdiffusion 66 -2560 66 -2560 0 cellNo=317
rlabel pdiffusion 73 -2560 73 -2560 0 cellNo=921
rlabel pdiffusion 80 -2560 80 -2560 0 feedthrough
rlabel pdiffusion 87 -2560 87 -2560 0 feedthrough
rlabel pdiffusion 94 -2560 94 -2560 0 feedthrough
rlabel pdiffusion 101 -2560 101 -2560 0 cellNo=190
rlabel pdiffusion 108 -2560 108 -2560 0 feedthrough
rlabel pdiffusion 115 -2560 115 -2560 0 feedthrough
rlabel pdiffusion 122 -2560 122 -2560 0 feedthrough
rlabel pdiffusion 129 -2560 129 -2560 0 feedthrough
rlabel pdiffusion 136 -2560 136 -2560 0 feedthrough
rlabel pdiffusion 143 -2560 143 -2560 0 feedthrough
rlabel pdiffusion 150 -2560 150 -2560 0 cellNo=226
rlabel pdiffusion 157 -2560 157 -2560 0 feedthrough
rlabel pdiffusion 164 -2560 164 -2560 0 cellNo=927
rlabel pdiffusion 171 -2560 171 -2560 0 cellNo=214
rlabel pdiffusion 178 -2560 178 -2560 0 feedthrough
rlabel pdiffusion 185 -2560 185 -2560 0 feedthrough
rlabel pdiffusion 192 -2560 192 -2560 0 feedthrough
rlabel pdiffusion 199 -2560 199 -2560 0 feedthrough
rlabel pdiffusion 206 -2560 206 -2560 0 feedthrough
rlabel pdiffusion 213 -2560 213 -2560 0 feedthrough
rlabel pdiffusion 220 -2560 220 -2560 0 feedthrough
rlabel pdiffusion 227 -2560 227 -2560 0 feedthrough
rlabel pdiffusion 234 -2560 234 -2560 0 feedthrough
rlabel pdiffusion 241 -2560 241 -2560 0 feedthrough
rlabel pdiffusion 248 -2560 248 -2560 0 feedthrough
rlabel pdiffusion 255 -2560 255 -2560 0 cellNo=904
rlabel pdiffusion 262 -2560 262 -2560 0 feedthrough
rlabel pdiffusion 269 -2560 269 -2560 0 feedthrough
rlabel pdiffusion 276 -2560 276 -2560 0 feedthrough
rlabel pdiffusion 283 -2560 283 -2560 0 feedthrough
rlabel pdiffusion 290 -2560 290 -2560 0 feedthrough
rlabel pdiffusion 297 -2560 297 -2560 0 feedthrough
rlabel pdiffusion 304 -2560 304 -2560 0 feedthrough
rlabel pdiffusion 311 -2560 311 -2560 0 feedthrough
rlabel pdiffusion 318 -2560 318 -2560 0 feedthrough
rlabel pdiffusion 325 -2560 325 -2560 0 feedthrough
rlabel pdiffusion 332 -2560 332 -2560 0 feedthrough
rlabel pdiffusion 339 -2560 339 -2560 0 feedthrough
rlabel pdiffusion 346 -2560 346 -2560 0 feedthrough
rlabel pdiffusion 353 -2560 353 -2560 0 feedthrough
rlabel pdiffusion 360 -2560 360 -2560 0 feedthrough
rlabel pdiffusion 367 -2560 367 -2560 0 feedthrough
rlabel pdiffusion 374 -2560 374 -2560 0 feedthrough
rlabel pdiffusion 381 -2560 381 -2560 0 feedthrough
rlabel pdiffusion 388 -2560 388 -2560 0 feedthrough
rlabel pdiffusion 395 -2560 395 -2560 0 feedthrough
rlabel pdiffusion 402 -2560 402 -2560 0 feedthrough
rlabel pdiffusion 409 -2560 409 -2560 0 cellNo=631
rlabel pdiffusion 416 -2560 416 -2560 0 feedthrough
rlabel pdiffusion 423 -2560 423 -2560 0 feedthrough
rlabel pdiffusion 430 -2560 430 -2560 0 cellNo=687
rlabel pdiffusion 437 -2560 437 -2560 0 feedthrough
rlabel pdiffusion 444 -2560 444 -2560 0 cellNo=740
rlabel pdiffusion 451 -2560 451 -2560 0 feedthrough
rlabel pdiffusion 458 -2560 458 -2560 0 feedthrough
rlabel pdiffusion 465 -2560 465 -2560 0 feedthrough
rlabel pdiffusion 472 -2560 472 -2560 0 feedthrough
rlabel pdiffusion 479 -2560 479 -2560 0 feedthrough
rlabel pdiffusion 486 -2560 486 -2560 0 feedthrough
rlabel pdiffusion 493 -2560 493 -2560 0 feedthrough
rlabel pdiffusion 500 -2560 500 -2560 0 feedthrough
rlabel pdiffusion 507 -2560 507 -2560 0 feedthrough
rlabel pdiffusion 514 -2560 514 -2560 0 feedthrough
rlabel pdiffusion 521 -2560 521 -2560 0 feedthrough
rlabel pdiffusion 528 -2560 528 -2560 0 feedthrough
rlabel pdiffusion 535 -2560 535 -2560 0 feedthrough
rlabel pdiffusion 542 -2560 542 -2560 0 feedthrough
rlabel pdiffusion 549 -2560 549 -2560 0 cellNo=323
rlabel pdiffusion 556 -2560 556 -2560 0 feedthrough
rlabel pdiffusion 563 -2560 563 -2560 0 feedthrough
rlabel pdiffusion 570 -2560 570 -2560 0 feedthrough
rlabel pdiffusion 577 -2560 577 -2560 0 feedthrough
rlabel pdiffusion 584 -2560 584 -2560 0 feedthrough
rlabel pdiffusion 591 -2560 591 -2560 0 cellNo=936
rlabel pdiffusion 598 -2560 598 -2560 0 feedthrough
rlabel pdiffusion 605 -2560 605 -2560 0 feedthrough
rlabel pdiffusion 612 -2560 612 -2560 0 feedthrough
rlabel pdiffusion 619 -2560 619 -2560 0 feedthrough
rlabel pdiffusion 626 -2560 626 -2560 0 cellNo=168
rlabel pdiffusion 633 -2560 633 -2560 0 feedthrough
rlabel pdiffusion 640 -2560 640 -2560 0 feedthrough
rlabel pdiffusion 647 -2560 647 -2560 0 cellNo=227
rlabel pdiffusion 654 -2560 654 -2560 0 feedthrough
rlabel pdiffusion 661 -2560 661 -2560 0 cellNo=67
rlabel pdiffusion 668 -2560 668 -2560 0 feedthrough
rlabel pdiffusion 675 -2560 675 -2560 0 feedthrough
rlabel pdiffusion 682 -2560 682 -2560 0 feedthrough
rlabel pdiffusion 689 -2560 689 -2560 0 feedthrough
rlabel pdiffusion 696 -2560 696 -2560 0 feedthrough
rlabel pdiffusion 703 -2560 703 -2560 0 feedthrough
rlabel pdiffusion 710 -2560 710 -2560 0 feedthrough
rlabel pdiffusion 717 -2560 717 -2560 0 feedthrough
rlabel pdiffusion 724 -2560 724 -2560 0 feedthrough
rlabel pdiffusion 731 -2560 731 -2560 0 cellNo=450
rlabel pdiffusion 738 -2560 738 -2560 0 cellNo=298
rlabel pdiffusion 745 -2560 745 -2560 0 cellNo=435
rlabel pdiffusion 752 -2560 752 -2560 0 cellNo=335
rlabel pdiffusion 759 -2560 759 -2560 0 feedthrough
rlabel pdiffusion 766 -2560 766 -2560 0 feedthrough
rlabel pdiffusion 773 -2560 773 -2560 0 feedthrough
rlabel pdiffusion 780 -2560 780 -2560 0 feedthrough
rlabel pdiffusion 787 -2560 787 -2560 0 cellNo=304
rlabel pdiffusion 794 -2560 794 -2560 0 feedthrough
rlabel pdiffusion 801 -2560 801 -2560 0 feedthrough
rlabel pdiffusion 808 -2560 808 -2560 0 feedthrough
rlabel pdiffusion 815 -2560 815 -2560 0 feedthrough
rlabel pdiffusion 822 -2560 822 -2560 0 cellNo=444
rlabel pdiffusion 829 -2560 829 -2560 0 feedthrough
rlabel pdiffusion 836 -2560 836 -2560 0 feedthrough
rlabel pdiffusion 843 -2560 843 -2560 0 feedthrough
rlabel pdiffusion 850 -2560 850 -2560 0 feedthrough
rlabel pdiffusion 857 -2560 857 -2560 0 feedthrough
rlabel pdiffusion 864 -2560 864 -2560 0 feedthrough
rlabel pdiffusion 871 -2560 871 -2560 0 cellNo=267
rlabel pdiffusion 878 -2560 878 -2560 0 feedthrough
rlabel pdiffusion 885 -2560 885 -2560 0 feedthrough
rlabel pdiffusion 892 -2560 892 -2560 0 feedthrough
rlabel pdiffusion 899 -2560 899 -2560 0 feedthrough
rlabel pdiffusion 906 -2560 906 -2560 0 feedthrough
rlabel pdiffusion 913 -2560 913 -2560 0 feedthrough
rlabel pdiffusion 920 -2560 920 -2560 0 feedthrough
rlabel pdiffusion 927 -2560 927 -2560 0 cellNo=83
rlabel pdiffusion 934 -2560 934 -2560 0 feedthrough
rlabel pdiffusion 941 -2560 941 -2560 0 feedthrough
rlabel pdiffusion 948 -2560 948 -2560 0 feedthrough
rlabel pdiffusion 955 -2560 955 -2560 0 cellNo=241
rlabel pdiffusion 962 -2560 962 -2560 0 feedthrough
rlabel pdiffusion 969 -2560 969 -2560 0 feedthrough
rlabel pdiffusion 976 -2560 976 -2560 0 feedthrough
rlabel pdiffusion 983 -2560 983 -2560 0 feedthrough
rlabel pdiffusion 990 -2560 990 -2560 0 feedthrough
rlabel pdiffusion 997 -2560 997 -2560 0 feedthrough
rlabel pdiffusion 1004 -2560 1004 -2560 0 feedthrough
rlabel pdiffusion 1011 -2560 1011 -2560 0 feedthrough
rlabel pdiffusion 1018 -2560 1018 -2560 0 feedthrough
rlabel pdiffusion 1025 -2560 1025 -2560 0 feedthrough
rlabel pdiffusion 1032 -2560 1032 -2560 0 feedthrough
rlabel pdiffusion 1039 -2560 1039 -2560 0 feedthrough
rlabel pdiffusion 1046 -2560 1046 -2560 0 feedthrough
rlabel pdiffusion 1053 -2560 1053 -2560 0 feedthrough
rlabel pdiffusion 1060 -2560 1060 -2560 0 cellNo=12
rlabel pdiffusion 1067 -2560 1067 -2560 0 feedthrough
rlabel pdiffusion 1074 -2560 1074 -2560 0 feedthrough
rlabel pdiffusion 1081 -2560 1081 -2560 0 cellNo=821
rlabel pdiffusion 1088 -2560 1088 -2560 0 cellNo=960
rlabel pdiffusion 1095 -2560 1095 -2560 0 feedthrough
rlabel pdiffusion 1102 -2560 1102 -2560 0 feedthrough
rlabel pdiffusion 1109 -2560 1109 -2560 0 feedthrough
rlabel pdiffusion 1116 -2560 1116 -2560 0 feedthrough
rlabel pdiffusion 1123 -2560 1123 -2560 0 feedthrough
rlabel pdiffusion 1130 -2560 1130 -2560 0 feedthrough
rlabel pdiffusion 1137 -2560 1137 -2560 0 feedthrough
rlabel pdiffusion 1144 -2560 1144 -2560 0 feedthrough
rlabel pdiffusion 1151 -2560 1151 -2560 0 feedthrough
rlabel pdiffusion 1158 -2560 1158 -2560 0 feedthrough
rlabel pdiffusion 1165 -2560 1165 -2560 0 cellNo=702
rlabel pdiffusion 1172 -2560 1172 -2560 0 feedthrough
rlabel pdiffusion 1179 -2560 1179 -2560 0 feedthrough
rlabel pdiffusion 1186 -2560 1186 -2560 0 cellNo=795
rlabel pdiffusion 1193 -2560 1193 -2560 0 feedthrough
rlabel pdiffusion 1200 -2560 1200 -2560 0 feedthrough
rlabel pdiffusion 1207 -2560 1207 -2560 0 feedthrough
rlabel pdiffusion 1214 -2560 1214 -2560 0 feedthrough
rlabel pdiffusion 1221 -2560 1221 -2560 0 feedthrough
rlabel pdiffusion 1228 -2560 1228 -2560 0 feedthrough
rlabel pdiffusion 1235 -2560 1235 -2560 0 feedthrough
rlabel pdiffusion 1242 -2560 1242 -2560 0 feedthrough
rlabel pdiffusion 1249 -2560 1249 -2560 0 feedthrough
rlabel pdiffusion 1256 -2560 1256 -2560 0 feedthrough
rlabel pdiffusion 1263 -2560 1263 -2560 0 feedthrough
rlabel pdiffusion 1270 -2560 1270 -2560 0 feedthrough
rlabel pdiffusion 1277 -2560 1277 -2560 0 feedthrough
rlabel pdiffusion 1284 -2560 1284 -2560 0 feedthrough
rlabel pdiffusion 1291 -2560 1291 -2560 0 feedthrough
rlabel pdiffusion 1298 -2560 1298 -2560 0 feedthrough
rlabel pdiffusion 1305 -2560 1305 -2560 0 feedthrough
rlabel pdiffusion 1312 -2560 1312 -2560 0 feedthrough
rlabel pdiffusion 1319 -2560 1319 -2560 0 feedthrough
rlabel pdiffusion 1326 -2560 1326 -2560 0 feedthrough
rlabel pdiffusion 1333 -2560 1333 -2560 0 feedthrough
rlabel pdiffusion 1340 -2560 1340 -2560 0 feedthrough
rlabel pdiffusion 1347 -2560 1347 -2560 0 feedthrough
rlabel pdiffusion 1354 -2560 1354 -2560 0 feedthrough
rlabel pdiffusion 1361 -2560 1361 -2560 0 feedthrough
rlabel pdiffusion 1368 -2560 1368 -2560 0 feedthrough
rlabel pdiffusion 1375 -2560 1375 -2560 0 feedthrough
rlabel pdiffusion 1382 -2560 1382 -2560 0 feedthrough
rlabel pdiffusion 1389 -2560 1389 -2560 0 feedthrough
rlabel pdiffusion 1396 -2560 1396 -2560 0 feedthrough
rlabel pdiffusion 1403 -2560 1403 -2560 0 feedthrough
rlabel pdiffusion 1410 -2560 1410 -2560 0 feedthrough
rlabel pdiffusion 1417 -2560 1417 -2560 0 feedthrough
rlabel pdiffusion 1424 -2560 1424 -2560 0 feedthrough
rlabel pdiffusion 1431 -2560 1431 -2560 0 feedthrough
rlabel pdiffusion 1438 -2560 1438 -2560 0 feedthrough
rlabel pdiffusion 1445 -2560 1445 -2560 0 feedthrough
rlabel pdiffusion 1452 -2560 1452 -2560 0 feedthrough
rlabel pdiffusion 1459 -2560 1459 -2560 0 feedthrough
rlabel pdiffusion 1466 -2560 1466 -2560 0 feedthrough
rlabel pdiffusion 1473 -2560 1473 -2560 0 feedthrough
rlabel pdiffusion 1480 -2560 1480 -2560 0 feedthrough
rlabel pdiffusion 1487 -2560 1487 -2560 0 feedthrough
rlabel pdiffusion 1494 -2560 1494 -2560 0 feedthrough
rlabel pdiffusion 1501 -2560 1501 -2560 0 feedthrough
rlabel pdiffusion 1508 -2560 1508 -2560 0 feedthrough
rlabel pdiffusion 1515 -2560 1515 -2560 0 feedthrough
rlabel pdiffusion 1522 -2560 1522 -2560 0 feedthrough
rlabel pdiffusion 1529 -2560 1529 -2560 0 feedthrough
rlabel pdiffusion 1536 -2560 1536 -2560 0 feedthrough
rlabel pdiffusion 1543 -2560 1543 -2560 0 feedthrough
rlabel pdiffusion 1550 -2560 1550 -2560 0 feedthrough
rlabel pdiffusion 1557 -2560 1557 -2560 0 feedthrough
rlabel pdiffusion 1564 -2560 1564 -2560 0 feedthrough
rlabel pdiffusion 1571 -2560 1571 -2560 0 feedthrough
rlabel pdiffusion 1578 -2560 1578 -2560 0 feedthrough
rlabel pdiffusion 1585 -2560 1585 -2560 0 feedthrough
rlabel pdiffusion 1592 -2560 1592 -2560 0 feedthrough
rlabel pdiffusion 1599 -2560 1599 -2560 0 feedthrough
rlabel pdiffusion 1606 -2560 1606 -2560 0 feedthrough
rlabel pdiffusion 1613 -2560 1613 -2560 0 feedthrough
rlabel pdiffusion 1620 -2560 1620 -2560 0 feedthrough
rlabel pdiffusion 1627 -2560 1627 -2560 0 feedthrough
rlabel pdiffusion 1634 -2560 1634 -2560 0 feedthrough
rlabel pdiffusion 1641 -2560 1641 -2560 0 feedthrough
rlabel pdiffusion 1648 -2560 1648 -2560 0 feedthrough
rlabel pdiffusion 1655 -2560 1655 -2560 0 feedthrough
rlabel pdiffusion 1662 -2560 1662 -2560 0 feedthrough
rlabel pdiffusion 1669 -2560 1669 -2560 0 feedthrough
rlabel pdiffusion 1676 -2560 1676 -2560 0 cellNo=363
rlabel pdiffusion 1683 -2560 1683 -2560 0 feedthrough
rlabel pdiffusion 1690 -2560 1690 -2560 0 feedthrough
rlabel pdiffusion 1697 -2560 1697 -2560 0 feedthrough
rlabel pdiffusion 1704 -2560 1704 -2560 0 cellNo=771
rlabel pdiffusion 1711 -2560 1711 -2560 0 feedthrough
rlabel pdiffusion 1718 -2560 1718 -2560 0 feedthrough
rlabel pdiffusion 1725 -2560 1725 -2560 0 feedthrough
rlabel pdiffusion 1732 -2560 1732 -2560 0 feedthrough
rlabel pdiffusion 1739 -2560 1739 -2560 0 feedthrough
rlabel pdiffusion 3 -2689 3 -2689 0 cellNo=1144
rlabel pdiffusion 10 -2689 10 -2689 0 cellNo=1151
rlabel pdiffusion 17 -2689 17 -2689 0 cellNo=1162
rlabel pdiffusion 24 -2689 24 -2689 0 cellNo=1176
rlabel pdiffusion 31 -2689 31 -2689 0 cellNo=1185
rlabel pdiffusion 38 -2689 38 -2689 0 cellNo=1196
rlabel pdiffusion 45 -2689 45 -2689 0 feedthrough
rlabel pdiffusion 52 -2689 52 -2689 0 feedthrough
rlabel pdiffusion 59 -2689 59 -2689 0 feedthrough
rlabel pdiffusion 66 -2689 66 -2689 0 cellNo=944
rlabel pdiffusion 73 -2689 73 -2689 0 feedthrough
rlabel pdiffusion 80 -2689 80 -2689 0 cellNo=422
rlabel pdiffusion 87 -2689 87 -2689 0 cellNo=248
rlabel pdiffusion 94 -2689 94 -2689 0 feedthrough
rlabel pdiffusion 101 -2689 101 -2689 0 feedthrough
rlabel pdiffusion 108 -2689 108 -2689 0 feedthrough
rlabel pdiffusion 115 -2689 115 -2689 0 cellNo=328
rlabel pdiffusion 122 -2689 122 -2689 0 feedthrough
rlabel pdiffusion 129 -2689 129 -2689 0 feedthrough
rlabel pdiffusion 136 -2689 136 -2689 0 feedthrough
rlabel pdiffusion 143 -2689 143 -2689 0 feedthrough
rlabel pdiffusion 150 -2689 150 -2689 0 feedthrough
rlabel pdiffusion 157 -2689 157 -2689 0 feedthrough
rlabel pdiffusion 164 -2689 164 -2689 0 cellNo=957
rlabel pdiffusion 171 -2689 171 -2689 0 feedthrough
rlabel pdiffusion 178 -2689 178 -2689 0 feedthrough
rlabel pdiffusion 185 -2689 185 -2689 0 feedthrough
rlabel pdiffusion 192 -2689 192 -2689 0 feedthrough
rlabel pdiffusion 199 -2689 199 -2689 0 cellNo=861
rlabel pdiffusion 206 -2689 206 -2689 0 feedthrough
rlabel pdiffusion 213 -2689 213 -2689 0 feedthrough
rlabel pdiffusion 220 -2689 220 -2689 0 feedthrough
rlabel pdiffusion 227 -2689 227 -2689 0 feedthrough
rlabel pdiffusion 234 -2689 234 -2689 0 feedthrough
rlabel pdiffusion 241 -2689 241 -2689 0 feedthrough
rlabel pdiffusion 248 -2689 248 -2689 0 cellNo=91
rlabel pdiffusion 255 -2689 255 -2689 0 feedthrough
rlabel pdiffusion 262 -2689 262 -2689 0 feedthrough
rlabel pdiffusion 269 -2689 269 -2689 0 feedthrough
rlabel pdiffusion 276 -2689 276 -2689 0 feedthrough
rlabel pdiffusion 283 -2689 283 -2689 0 feedthrough
rlabel pdiffusion 290 -2689 290 -2689 0 feedthrough
rlabel pdiffusion 297 -2689 297 -2689 0 feedthrough
rlabel pdiffusion 304 -2689 304 -2689 0 feedthrough
rlabel pdiffusion 311 -2689 311 -2689 0 feedthrough
rlabel pdiffusion 318 -2689 318 -2689 0 feedthrough
rlabel pdiffusion 325 -2689 325 -2689 0 feedthrough
rlabel pdiffusion 332 -2689 332 -2689 0 feedthrough
rlabel pdiffusion 339 -2689 339 -2689 0 feedthrough
rlabel pdiffusion 346 -2689 346 -2689 0 feedthrough
rlabel pdiffusion 353 -2689 353 -2689 0 feedthrough
rlabel pdiffusion 360 -2689 360 -2689 0 feedthrough
rlabel pdiffusion 367 -2689 367 -2689 0 feedthrough
rlabel pdiffusion 374 -2689 374 -2689 0 feedthrough
rlabel pdiffusion 381 -2689 381 -2689 0 feedthrough
rlabel pdiffusion 388 -2689 388 -2689 0 feedthrough
rlabel pdiffusion 395 -2689 395 -2689 0 feedthrough
rlabel pdiffusion 402 -2689 402 -2689 0 feedthrough
rlabel pdiffusion 409 -2689 409 -2689 0 cellNo=86
rlabel pdiffusion 416 -2689 416 -2689 0 cellNo=26
rlabel pdiffusion 423 -2689 423 -2689 0 feedthrough
rlabel pdiffusion 430 -2689 430 -2689 0 feedthrough
rlabel pdiffusion 437 -2689 437 -2689 0 feedthrough
rlabel pdiffusion 444 -2689 444 -2689 0 feedthrough
rlabel pdiffusion 451 -2689 451 -2689 0 cellNo=287
rlabel pdiffusion 458 -2689 458 -2689 0 cellNo=731
rlabel pdiffusion 465 -2689 465 -2689 0 cellNo=615
rlabel pdiffusion 472 -2689 472 -2689 0 feedthrough
rlabel pdiffusion 479 -2689 479 -2689 0 cellNo=327
rlabel pdiffusion 486 -2689 486 -2689 0 feedthrough
rlabel pdiffusion 493 -2689 493 -2689 0 feedthrough
rlabel pdiffusion 500 -2689 500 -2689 0 feedthrough
rlabel pdiffusion 507 -2689 507 -2689 0 feedthrough
rlabel pdiffusion 514 -2689 514 -2689 0 feedthrough
rlabel pdiffusion 521 -2689 521 -2689 0 feedthrough
rlabel pdiffusion 528 -2689 528 -2689 0 feedthrough
rlabel pdiffusion 535 -2689 535 -2689 0 feedthrough
rlabel pdiffusion 542 -2689 542 -2689 0 feedthrough
rlabel pdiffusion 549 -2689 549 -2689 0 feedthrough
rlabel pdiffusion 556 -2689 556 -2689 0 feedthrough
rlabel pdiffusion 563 -2689 563 -2689 0 feedthrough
rlabel pdiffusion 570 -2689 570 -2689 0 feedthrough
rlabel pdiffusion 577 -2689 577 -2689 0 cellNo=875
rlabel pdiffusion 584 -2689 584 -2689 0 feedthrough
rlabel pdiffusion 591 -2689 591 -2689 0 feedthrough
rlabel pdiffusion 598 -2689 598 -2689 0 cellNo=456
rlabel pdiffusion 605 -2689 605 -2689 0 feedthrough
rlabel pdiffusion 612 -2689 612 -2689 0 feedthrough
rlabel pdiffusion 619 -2689 619 -2689 0 feedthrough
rlabel pdiffusion 626 -2689 626 -2689 0 cellNo=139
rlabel pdiffusion 633 -2689 633 -2689 0 feedthrough
rlabel pdiffusion 640 -2689 640 -2689 0 feedthrough
rlabel pdiffusion 647 -2689 647 -2689 0 feedthrough
rlabel pdiffusion 654 -2689 654 -2689 0 feedthrough
rlabel pdiffusion 661 -2689 661 -2689 0 feedthrough
rlabel pdiffusion 668 -2689 668 -2689 0 cellNo=566
rlabel pdiffusion 675 -2689 675 -2689 0 cellNo=59
rlabel pdiffusion 682 -2689 682 -2689 0 feedthrough
rlabel pdiffusion 689 -2689 689 -2689 0 cellNo=621
rlabel pdiffusion 696 -2689 696 -2689 0 feedthrough
rlabel pdiffusion 703 -2689 703 -2689 0 feedthrough
rlabel pdiffusion 710 -2689 710 -2689 0 feedthrough
rlabel pdiffusion 717 -2689 717 -2689 0 feedthrough
rlabel pdiffusion 724 -2689 724 -2689 0 feedthrough
rlabel pdiffusion 731 -2689 731 -2689 0 cellNo=429
rlabel pdiffusion 738 -2689 738 -2689 0 feedthrough
rlabel pdiffusion 745 -2689 745 -2689 0 feedthrough
rlabel pdiffusion 752 -2689 752 -2689 0 cellNo=325
rlabel pdiffusion 759 -2689 759 -2689 0 feedthrough
rlabel pdiffusion 766 -2689 766 -2689 0 cellNo=735
rlabel pdiffusion 773 -2689 773 -2689 0 feedthrough
rlabel pdiffusion 780 -2689 780 -2689 0 feedthrough
rlabel pdiffusion 787 -2689 787 -2689 0 feedthrough
rlabel pdiffusion 794 -2689 794 -2689 0 feedthrough
rlabel pdiffusion 801 -2689 801 -2689 0 cellNo=954
rlabel pdiffusion 808 -2689 808 -2689 0 feedthrough
rlabel pdiffusion 815 -2689 815 -2689 0 feedthrough
rlabel pdiffusion 822 -2689 822 -2689 0 feedthrough
rlabel pdiffusion 829 -2689 829 -2689 0 feedthrough
rlabel pdiffusion 836 -2689 836 -2689 0 cellNo=120
rlabel pdiffusion 843 -2689 843 -2689 0 cellNo=865
rlabel pdiffusion 850 -2689 850 -2689 0 feedthrough
rlabel pdiffusion 857 -2689 857 -2689 0 feedthrough
rlabel pdiffusion 864 -2689 864 -2689 0 feedthrough
rlabel pdiffusion 871 -2689 871 -2689 0 cellNo=730
rlabel pdiffusion 878 -2689 878 -2689 0 feedthrough
rlabel pdiffusion 885 -2689 885 -2689 0 feedthrough
rlabel pdiffusion 892 -2689 892 -2689 0 cellNo=250
rlabel pdiffusion 899 -2689 899 -2689 0 feedthrough
rlabel pdiffusion 906 -2689 906 -2689 0 feedthrough
rlabel pdiffusion 913 -2689 913 -2689 0 feedthrough
rlabel pdiffusion 920 -2689 920 -2689 0 feedthrough
rlabel pdiffusion 927 -2689 927 -2689 0 feedthrough
rlabel pdiffusion 934 -2689 934 -2689 0 feedthrough
rlabel pdiffusion 941 -2689 941 -2689 0 feedthrough
rlabel pdiffusion 948 -2689 948 -2689 0 feedthrough
rlabel pdiffusion 955 -2689 955 -2689 0 cellNo=346
rlabel pdiffusion 962 -2689 962 -2689 0 feedthrough
rlabel pdiffusion 969 -2689 969 -2689 0 feedthrough
rlabel pdiffusion 976 -2689 976 -2689 0 feedthrough
rlabel pdiffusion 983 -2689 983 -2689 0 feedthrough
rlabel pdiffusion 990 -2689 990 -2689 0 cellNo=709
rlabel pdiffusion 997 -2689 997 -2689 0 feedthrough
rlabel pdiffusion 1004 -2689 1004 -2689 0 feedthrough
rlabel pdiffusion 1011 -2689 1011 -2689 0 feedthrough
rlabel pdiffusion 1018 -2689 1018 -2689 0 feedthrough
rlabel pdiffusion 1025 -2689 1025 -2689 0 feedthrough
rlabel pdiffusion 1032 -2689 1032 -2689 0 cellNo=218
rlabel pdiffusion 1039 -2689 1039 -2689 0 feedthrough
rlabel pdiffusion 1046 -2689 1046 -2689 0 feedthrough
rlabel pdiffusion 1053 -2689 1053 -2689 0 feedthrough
rlabel pdiffusion 1060 -2689 1060 -2689 0 feedthrough
rlabel pdiffusion 1067 -2689 1067 -2689 0 feedthrough
rlabel pdiffusion 1074 -2689 1074 -2689 0 feedthrough
rlabel pdiffusion 1081 -2689 1081 -2689 0 feedthrough
rlabel pdiffusion 1088 -2689 1088 -2689 0 feedthrough
rlabel pdiffusion 1095 -2689 1095 -2689 0 cellNo=698
rlabel pdiffusion 1102 -2689 1102 -2689 0 feedthrough
rlabel pdiffusion 1109 -2689 1109 -2689 0 feedthrough
rlabel pdiffusion 1116 -2689 1116 -2689 0 feedthrough
rlabel pdiffusion 1123 -2689 1123 -2689 0 feedthrough
rlabel pdiffusion 1130 -2689 1130 -2689 0 feedthrough
rlabel pdiffusion 1137 -2689 1137 -2689 0 feedthrough
rlabel pdiffusion 1144 -2689 1144 -2689 0 feedthrough
rlabel pdiffusion 1151 -2689 1151 -2689 0 feedthrough
rlabel pdiffusion 1158 -2689 1158 -2689 0 feedthrough
rlabel pdiffusion 1165 -2689 1165 -2689 0 feedthrough
rlabel pdiffusion 1172 -2689 1172 -2689 0 feedthrough
rlabel pdiffusion 1179 -2689 1179 -2689 0 feedthrough
rlabel pdiffusion 1186 -2689 1186 -2689 0 feedthrough
rlabel pdiffusion 1193 -2689 1193 -2689 0 feedthrough
rlabel pdiffusion 1200 -2689 1200 -2689 0 feedthrough
rlabel pdiffusion 1207 -2689 1207 -2689 0 feedthrough
rlabel pdiffusion 1214 -2689 1214 -2689 0 feedthrough
rlabel pdiffusion 1221 -2689 1221 -2689 0 feedthrough
rlabel pdiffusion 1228 -2689 1228 -2689 0 feedthrough
rlabel pdiffusion 1235 -2689 1235 -2689 0 feedthrough
rlabel pdiffusion 1242 -2689 1242 -2689 0 feedthrough
rlabel pdiffusion 1249 -2689 1249 -2689 0 feedthrough
rlabel pdiffusion 1256 -2689 1256 -2689 0 feedthrough
rlabel pdiffusion 1263 -2689 1263 -2689 0 feedthrough
rlabel pdiffusion 1270 -2689 1270 -2689 0 feedthrough
rlabel pdiffusion 1277 -2689 1277 -2689 0 feedthrough
rlabel pdiffusion 1284 -2689 1284 -2689 0 feedthrough
rlabel pdiffusion 1291 -2689 1291 -2689 0 feedthrough
rlabel pdiffusion 1298 -2689 1298 -2689 0 feedthrough
rlabel pdiffusion 1305 -2689 1305 -2689 0 feedthrough
rlabel pdiffusion 1312 -2689 1312 -2689 0 feedthrough
rlabel pdiffusion 1319 -2689 1319 -2689 0 feedthrough
rlabel pdiffusion 1326 -2689 1326 -2689 0 feedthrough
rlabel pdiffusion 1333 -2689 1333 -2689 0 feedthrough
rlabel pdiffusion 1340 -2689 1340 -2689 0 feedthrough
rlabel pdiffusion 1347 -2689 1347 -2689 0 feedthrough
rlabel pdiffusion 1354 -2689 1354 -2689 0 feedthrough
rlabel pdiffusion 1361 -2689 1361 -2689 0 feedthrough
rlabel pdiffusion 1368 -2689 1368 -2689 0 feedthrough
rlabel pdiffusion 1375 -2689 1375 -2689 0 feedthrough
rlabel pdiffusion 1382 -2689 1382 -2689 0 feedthrough
rlabel pdiffusion 1389 -2689 1389 -2689 0 feedthrough
rlabel pdiffusion 1396 -2689 1396 -2689 0 feedthrough
rlabel pdiffusion 1403 -2689 1403 -2689 0 feedthrough
rlabel pdiffusion 1410 -2689 1410 -2689 0 feedthrough
rlabel pdiffusion 1417 -2689 1417 -2689 0 feedthrough
rlabel pdiffusion 1424 -2689 1424 -2689 0 feedthrough
rlabel pdiffusion 1431 -2689 1431 -2689 0 feedthrough
rlabel pdiffusion 1438 -2689 1438 -2689 0 feedthrough
rlabel pdiffusion 1445 -2689 1445 -2689 0 feedthrough
rlabel pdiffusion 1452 -2689 1452 -2689 0 feedthrough
rlabel pdiffusion 1459 -2689 1459 -2689 0 feedthrough
rlabel pdiffusion 1466 -2689 1466 -2689 0 feedthrough
rlabel pdiffusion 1473 -2689 1473 -2689 0 feedthrough
rlabel pdiffusion 1480 -2689 1480 -2689 0 feedthrough
rlabel pdiffusion 1487 -2689 1487 -2689 0 feedthrough
rlabel pdiffusion 1494 -2689 1494 -2689 0 feedthrough
rlabel pdiffusion 1501 -2689 1501 -2689 0 feedthrough
rlabel pdiffusion 1508 -2689 1508 -2689 0 feedthrough
rlabel pdiffusion 1515 -2689 1515 -2689 0 feedthrough
rlabel pdiffusion 1522 -2689 1522 -2689 0 feedthrough
rlabel pdiffusion 1529 -2689 1529 -2689 0 feedthrough
rlabel pdiffusion 1536 -2689 1536 -2689 0 feedthrough
rlabel pdiffusion 1543 -2689 1543 -2689 0 feedthrough
rlabel pdiffusion 1550 -2689 1550 -2689 0 feedthrough
rlabel pdiffusion 1557 -2689 1557 -2689 0 feedthrough
rlabel pdiffusion 1564 -2689 1564 -2689 0 feedthrough
rlabel pdiffusion 1571 -2689 1571 -2689 0 feedthrough
rlabel pdiffusion 1578 -2689 1578 -2689 0 feedthrough
rlabel pdiffusion 1585 -2689 1585 -2689 0 feedthrough
rlabel pdiffusion 1592 -2689 1592 -2689 0 feedthrough
rlabel pdiffusion 1599 -2689 1599 -2689 0 feedthrough
rlabel pdiffusion 1606 -2689 1606 -2689 0 feedthrough
rlabel pdiffusion 1613 -2689 1613 -2689 0 feedthrough
rlabel pdiffusion 1620 -2689 1620 -2689 0 feedthrough
rlabel pdiffusion 1627 -2689 1627 -2689 0 feedthrough
rlabel pdiffusion 1634 -2689 1634 -2689 0 feedthrough
rlabel pdiffusion 1641 -2689 1641 -2689 0 feedthrough
rlabel pdiffusion 1648 -2689 1648 -2689 0 feedthrough
rlabel pdiffusion 1655 -2689 1655 -2689 0 feedthrough
rlabel pdiffusion 1662 -2689 1662 -2689 0 feedthrough
rlabel pdiffusion 1669 -2689 1669 -2689 0 feedthrough
rlabel pdiffusion 1676 -2689 1676 -2689 0 feedthrough
rlabel pdiffusion 1683 -2689 1683 -2689 0 feedthrough
rlabel pdiffusion 1690 -2689 1690 -2689 0 feedthrough
rlabel pdiffusion 1697 -2689 1697 -2689 0 feedthrough
rlabel pdiffusion 1704 -2689 1704 -2689 0 feedthrough
rlabel pdiffusion 3 -2838 3 -2838 0 cellNo=1150
rlabel pdiffusion 10 -2838 10 -2838 0 cellNo=1160
rlabel pdiffusion 17 -2838 17 -2838 0 cellNo=1174
rlabel pdiffusion 24 -2838 24 -2838 0 cellNo=1184
rlabel pdiffusion 31 -2838 31 -2838 0 cellNo=1195
rlabel pdiffusion 38 -2838 38 -2838 0 feedthrough
rlabel pdiffusion 45 -2838 45 -2838 0 feedthrough
rlabel pdiffusion 52 -2838 52 -2838 0 feedthrough
rlabel pdiffusion 59 -2838 59 -2838 0 feedthrough
rlabel pdiffusion 66 -2838 66 -2838 0 feedthrough
rlabel pdiffusion 73 -2838 73 -2838 0 feedthrough
rlabel pdiffusion 80 -2838 80 -2838 0 feedthrough
rlabel pdiffusion 87 -2838 87 -2838 0 cellNo=581
rlabel pdiffusion 94 -2838 94 -2838 0 cellNo=98
rlabel pdiffusion 101 -2838 101 -2838 0 feedthrough
rlabel pdiffusion 108 -2838 108 -2838 0 cellNo=420
rlabel pdiffusion 115 -2838 115 -2838 0 feedthrough
rlabel pdiffusion 122 -2838 122 -2838 0 feedthrough
rlabel pdiffusion 129 -2838 129 -2838 0 cellNo=868
rlabel pdiffusion 136 -2838 136 -2838 0 feedthrough
rlabel pdiffusion 143 -2838 143 -2838 0 feedthrough
rlabel pdiffusion 150 -2838 150 -2838 0 feedthrough
rlabel pdiffusion 157 -2838 157 -2838 0 feedthrough
rlabel pdiffusion 164 -2838 164 -2838 0 cellNo=88
rlabel pdiffusion 171 -2838 171 -2838 0 feedthrough
rlabel pdiffusion 178 -2838 178 -2838 0 cellNo=178
rlabel pdiffusion 185 -2838 185 -2838 0 feedthrough
rlabel pdiffusion 192 -2838 192 -2838 0 feedthrough
rlabel pdiffusion 199 -2838 199 -2838 0 feedthrough
rlabel pdiffusion 206 -2838 206 -2838 0 feedthrough
rlabel pdiffusion 213 -2838 213 -2838 0 feedthrough
rlabel pdiffusion 220 -2838 220 -2838 0 feedthrough
rlabel pdiffusion 227 -2838 227 -2838 0 cellNo=930
rlabel pdiffusion 234 -2838 234 -2838 0 feedthrough
rlabel pdiffusion 241 -2838 241 -2838 0 feedthrough
rlabel pdiffusion 248 -2838 248 -2838 0 cellNo=934
rlabel pdiffusion 255 -2838 255 -2838 0 feedthrough
rlabel pdiffusion 262 -2838 262 -2838 0 feedthrough
rlabel pdiffusion 269 -2838 269 -2838 0 feedthrough
rlabel pdiffusion 276 -2838 276 -2838 0 feedthrough
rlabel pdiffusion 283 -2838 283 -2838 0 feedthrough
rlabel pdiffusion 290 -2838 290 -2838 0 feedthrough
rlabel pdiffusion 297 -2838 297 -2838 0 feedthrough
rlabel pdiffusion 304 -2838 304 -2838 0 feedthrough
rlabel pdiffusion 311 -2838 311 -2838 0 feedthrough
rlabel pdiffusion 318 -2838 318 -2838 0 feedthrough
rlabel pdiffusion 325 -2838 325 -2838 0 feedthrough
rlabel pdiffusion 332 -2838 332 -2838 0 feedthrough
rlabel pdiffusion 339 -2838 339 -2838 0 feedthrough
rlabel pdiffusion 346 -2838 346 -2838 0 feedthrough
rlabel pdiffusion 353 -2838 353 -2838 0 feedthrough
rlabel pdiffusion 360 -2838 360 -2838 0 feedthrough
rlabel pdiffusion 367 -2838 367 -2838 0 feedthrough
rlabel pdiffusion 374 -2838 374 -2838 0 feedthrough
rlabel pdiffusion 381 -2838 381 -2838 0 cellNo=162
rlabel pdiffusion 388 -2838 388 -2838 0 feedthrough
rlabel pdiffusion 395 -2838 395 -2838 0 feedthrough
rlabel pdiffusion 402 -2838 402 -2838 0 feedthrough
rlabel pdiffusion 409 -2838 409 -2838 0 feedthrough
rlabel pdiffusion 416 -2838 416 -2838 0 feedthrough
rlabel pdiffusion 423 -2838 423 -2838 0 feedthrough
rlabel pdiffusion 430 -2838 430 -2838 0 feedthrough
rlabel pdiffusion 437 -2838 437 -2838 0 feedthrough
rlabel pdiffusion 444 -2838 444 -2838 0 feedthrough
rlabel pdiffusion 451 -2838 451 -2838 0 cellNo=603
rlabel pdiffusion 458 -2838 458 -2838 0 feedthrough
rlabel pdiffusion 465 -2838 465 -2838 0 feedthrough
rlabel pdiffusion 472 -2838 472 -2838 0 feedthrough
rlabel pdiffusion 479 -2838 479 -2838 0 feedthrough
rlabel pdiffusion 486 -2838 486 -2838 0 feedthrough
rlabel pdiffusion 493 -2838 493 -2838 0 feedthrough
rlabel pdiffusion 500 -2838 500 -2838 0 feedthrough
rlabel pdiffusion 507 -2838 507 -2838 0 feedthrough
rlabel pdiffusion 514 -2838 514 -2838 0 feedthrough
rlabel pdiffusion 521 -2838 521 -2838 0 cellNo=284
rlabel pdiffusion 528 -2838 528 -2838 0 feedthrough
rlabel pdiffusion 535 -2838 535 -2838 0 feedthrough
rlabel pdiffusion 542 -2838 542 -2838 0 feedthrough
rlabel pdiffusion 549 -2838 549 -2838 0 feedthrough
rlabel pdiffusion 556 -2838 556 -2838 0 feedthrough
rlabel pdiffusion 563 -2838 563 -2838 0 feedthrough
rlabel pdiffusion 570 -2838 570 -2838 0 feedthrough
rlabel pdiffusion 577 -2838 577 -2838 0 feedthrough
rlabel pdiffusion 584 -2838 584 -2838 0 feedthrough
rlabel pdiffusion 591 -2838 591 -2838 0 cellNo=522
rlabel pdiffusion 598 -2838 598 -2838 0 feedthrough
rlabel pdiffusion 605 -2838 605 -2838 0 feedthrough
rlabel pdiffusion 612 -2838 612 -2838 0 feedthrough
rlabel pdiffusion 619 -2838 619 -2838 0 feedthrough
rlabel pdiffusion 626 -2838 626 -2838 0 feedthrough
rlabel pdiffusion 633 -2838 633 -2838 0 feedthrough
rlabel pdiffusion 640 -2838 640 -2838 0 feedthrough
rlabel pdiffusion 647 -2838 647 -2838 0 cellNo=484
rlabel pdiffusion 654 -2838 654 -2838 0 cellNo=517
rlabel pdiffusion 661 -2838 661 -2838 0 feedthrough
rlabel pdiffusion 668 -2838 668 -2838 0 feedthrough
rlabel pdiffusion 675 -2838 675 -2838 0 feedthrough
rlabel pdiffusion 682 -2838 682 -2838 0 cellNo=309
rlabel pdiffusion 689 -2838 689 -2838 0 feedthrough
rlabel pdiffusion 696 -2838 696 -2838 0 feedthrough
rlabel pdiffusion 703 -2838 703 -2838 0 feedthrough
rlabel pdiffusion 710 -2838 710 -2838 0 feedthrough
rlabel pdiffusion 717 -2838 717 -2838 0 feedthrough
rlabel pdiffusion 724 -2838 724 -2838 0 feedthrough
rlabel pdiffusion 731 -2838 731 -2838 0 feedthrough
rlabel pdiffusion 738 -2838 738 -2838 0 feedthrough
rlabel pdiffusion 745 -2838 745 -2838 0 feedthrough
rlabel pdiffusion 752 -2838 752 -2838 0 feedthrough
rlabel pdiffusion 759 -2838 759 -2838 0 cellNo=315
rlabel pdiffusion 766 -2838 766 -2838 0 cellNo=402
rlabel pdiffusion 773 -2838 773 -2838 0 cellNo=828
rlabel pdiffusion 780 -2838 780 -2838 0 feedthrough
rlabel pdiffusion 787 -2838 787 -2838 0 feedthrough
rlabel pdiffusion 794 -2838 794 -2838 0 feedthrough
rlabel pdiffusion 801 -2838 801 -2838 0 cellNo=101
rlabel pdiffusion 808 -2838 808 -2838 0 feedthrough
rlabel pdiffusion 815 -2838 815 -2838 0 feedthrough
rlabel pdiffusion 822 -2838 822 -2838 0 feedthrough
rlabel pdiffusion 829 -2838 829 -2838 0 feedthrough
rlabel pdiffusion 836 -2838 836 -2838 0 feedthrough
rlabel pdiffusion 843 -2838 843 -2838 0 feedthrough
rlabel pdiffusion 850 -2838 850 -2838 0 feedthrough
rlabel pdiffusion 857 -2838 857 -2838 0 feedthrough
rlabel pdiffusion 864 -2838 864 -2838 0 feedthrough
rlabel pdiffusion 871 -2838 871 -2838 0 feedthrough
rlabel pdiffusion 878 -2838 878 -2838 0 feedthrough
rlabel pdiffusion 885 -2838 885 -2838 0 cellNo=66
rlabel pdiffusion 892 -2838 892 -2838 0 cellNo=105
rlabel pdiffusion 899 -2838 899 -2838 0 cellNo=619
rlabel pdiffusion 906 -2838 906 -2838 0 feedthrough
rlabel pdiffusion 913 -2838 913 -2838 0 feedthrough
rlabel pdiffusion 920 -2838 920 -2838 0 feedthrough
rlabel pdiffusion 927 -2838 927 -2838 0 feedthrough
rlabel pdiffusion 934 -2838 934 -2838 0 feedthrough
rlabel pdiffusion 941 -2838 941 -2838 0 feedthrough
rlabel pdiffusion 948 -2838 948 -2838 0 feedthrough
rlabel pdiffusion 955 -2838 955 -2838 0 feedthrough
rlabel pdiffusion 962 -2838 962 -2838 0 feedthrough
rlabel pdiffusion 969 -2838 969 -2838 0 feedthrough
rlabel pdiffusion 976 -2838 976 -2838 0 feedthrough
rlabel pdiffusion 983 -2838 983 -2838 0 cellNo=417
rlabel pdiffusion 990 -2838 990 -2838 0 feedthrough
rlabel pdiffusion 997 -2838 997 -2838 0 cellNo=126
rlabel pdiffusion 1004 -2838 1004 -2838 0 feedthrough
rlabel pdiffusion 1011 -2838 1011 -2838 0 feedthrough
rlabel pdiffusion 1018 -2838 1018 -2838 0 feedthrough
rlabel pdiffusion 1025 -2838 1025 -2838 0 feedthrough
rlabel pdiffusion 1032 -2838 1032 -2838 0 feedthrough
rlabel pdiffusion 1039 -2838 1039 -2838 0 feedthrough
rlabel pdiffusion 1046 -2838 1046 -2838 0 cellNo=654
rlabel pdiffusion 1053 -2838 1053 -2838 0 feedthrough
rlabel pdiffusion 1060 -2838 1060 -2838 0 feedthrough
rlabel pdiffusion 1067 -2838 1067 -2838 0 feedthrough
rlabel pdiffusion 1074 -2838 1074 -2838 0 feedthrough
rlabel pdiffusion 1081 -2838 1081 -2838 0 feedthrough
rlabel pdiffusion 1088 -2838 1088 -2838 0 feedthrough
rlabel pdiffusion 1095 -2838 1095 -2838 0 cellNo=841
rlabel pdiffusion 1102 -2838 1102 -2838 0 feedthrough
rlabel pdiffusion 1109 -2838 1109 -2838 0 feedthrough
rlabel pdiffusion 1116 -2838 1116 -2838 0 cellNo=49
rlabel pdiffusion 1123 -2838 1123 -2838 0 feedthrough
rlabel pdiffusion 1130 -2838 1130 -2838 0 feedthrough
rlabel pdiffusion 1137 -2838 1137 -2838 0 feedthrough
rlabel pdiffusion 1144 -2838 1144 -2838 0 feedthrough
rlabel pdiffusion 1151 -2838 1151 -2838 0 feedthrough
rlabel pdiffusion 1158 -2838 1158 -2838 0 feedthrough
rlabel pdiffusion 1165 -2838 1165 -2838 0 feedthrough
rlabel pdiffusion 1172 -2838 1172 -2838 0 feedthrough
rlabel pdiffusion 1179 -2838 1179 -2838 0 feedthrough
rlabel pdiffusion 1186 -2838 1186 -2838 0 cellNo=553
rlabel pdiffusion 1193 -2838 1193 -2838 0 feedthrough
rlabel pdiffusion 1200 -2838 1200 -2838 0 feedthrough
rlabel pdiffusion 1207 -2838 1207 -2838 0 feedthrough
rlabel pdiffusion 1214 -2838 1214 -2838 0 feedthrough
rlabel pdiffusion 1221 -2838 1221 -2838 0 feedthrough
rlabel pdiffusion 1228 -2838 1228 -2838 0 feedthrough
rlabel pdiffusion 1235 -2838 1235 -2838 0 feedthrough
rlabel pdiffusion 1242 -2838 1242 -2838 0 feedthrough
rlabel pdiffusion 1249 -2838 1249 -2838 0 feedthrough
rlabel pdiffusion 1256 -2838 1256 -2838 0 feedthrough
rlabel pdiffusion 1263 -2838 1263 -2838 0 feedthrough
rlabel pdiffusion 1270 -2838 1270 -2838 0 feedthrough
rlabel pdiffusion 1277 -2838 1277 -2838 0 cellNo=755
rlabel pdiffusion 1284 -2838 1284 -2838 0 feedthrough
rlabel pdiffusion 1291 -2838 1291 -2838 0 feedthrough
rlabel pdiffusion 1298 -2838 1298 -2838 0 feedthrough
rlabel pdiffusion 1305 -2838 1305 -2838 0 feedthrough
rlabel pdiffusion 1312 -2838 1312 -2838 0 feedthrough
rlabel pdiffusion 1319 -2838 1319 -2838 0 feedthrough
rlabel pdiffusion 1326 -2838 1326 -2838 0 feedthrough
rlabel pdiffusion 1333 -2838 1333 -2838 0 feedthrough
rlabel pdiffusion 1340 -2838 1340 -2838 0 feedthrough
rlabel pdiffusion 1347 -2838 1347 -2838 0 feedthrough
rlabel pdiffusion 1354 -2838 1354 -2838 0 feedthrough
rlabel pdiffusion 1361 -2838 1361 -2838 0 feedthrough
rlabel pdiffusion 1368 -2838 1368 -2838 0 feedthrough
rlabel pdiffusion 1375 -2838 1375 -2838 0 feedthrough
rlabel pdiffusion 1382 -2838 1382 -2838 0 feedthrough
rlabel pdiffusion 1389 -2838 1389 -2838 0 feedthrough
rlabel pdiffusion 1396 -2838 1396 -2838 0 feedthrough
rlabel pdiffusion 1403 -2838 1403 -2838 0 feedthrough
rlabel pdiffusion 1410 -2838 1410 -2838 0 feedthrough
rlabel pdiffusion 1417 -2838 1417 -2838 0 feedthrough
rlabel pdiffusion 1424 -2838 1424 -2838 0 feedthrough
rlabel pdiffusion 1431 -2838 1431 -2838 0 feedthrough
rlabel pdiffusion 1438 -2838 1438 -2838 0 feedthrough
rlabel pdiffusion 1445 -2838 1445 -2838 0 feedthrough
rlabel pdiffusion 1452 -2838 1452 -2838 0 feedthrough
rlabel pdiffusion 1459 -2838 1459 -2838 0 feedthrough
rlabel pdiffusion 1466 -2838 1466 -2838 0 feedthrough
rlabel pdiffusion 1473 -2838 1473 -2838 0 feedthrough
rlabel pdiffusion 1480 -2838 1480 -2838 0 feedthrough
rlabel pdiffusion 1487 -2838 1487 -2838 0 feedthrough
rlabel pdiffusion 1494 -2838 1494 -2838 0 feedthrough
rlabel pdiffusion 1501 -2838 1501 -2838 0 feedthrough
rlabel pdiffusion 1508 -2838 1508 -2838 0 cellNo=419
rlabel pdiffusion 1515 -2838 1515 -2838 0 cellNo=635
rlabel pdiffusion 1522 -2838 1522 -2838 0 feedthrough
rlabel pdiffusion 1529 -2838 1529 -2838 0 feedthrough
rlabel pdiffusion 1536 -2838 1536 -2838 0 feedthrough
rlabel pdiffusion 1543 -2838 1543 -2838 0 feedthrough
rlabel pdiffusion 1550 -2838 1550 -2838 0 feedthrough
rlabel pdiffusion 1557 -2838 1557 -2838 0 feedthrough
rlabel pdiffusion 3 -2949 3 -2949 0 cellNo=1159
rlabel pdiffusion 10 -2949 10 -2949 0 cellNo=1173
rlabel pdiffusion 17 -2949 17 -2949 0 cellNo=1183
rlabel pdiffusion 24 -2949 24 -2949 0 cellNo=1194
rlabel pdiffusion 31 -2949 31 -2949 0 feedthrough
rlabel pdiffusion 38 -2949 38 -2949 0 feedthrough
rlabel pdiffusion 45 -2949 45 -2949 0 feedthrough
rlabel pdiffusion 52 -2949 52 -2949 0 feedthrough
rlabel pdiffusion 59 -2949 59 -2949 0 feedthrough
rlabel pdiffusion 66 -2949 66 -2949 0 feedthrough
rlabel pdiffusion 73 -2949 73 -2949 0 cellNo=135
rlabel pdiffusion 80 -2949 80 -2949 0 feedthrough
rlabel pdiffusion 87 -2949 87 -2949 0 feedthrough
rlabel pdiffusion 94 -2949 94 -2949 0 feedthrough
rlabel pdiffusion 101 -2949 101 -2949 0 feedthrough
rlabel pdiffusion 108 -2949 108 -2949 0 feedthrough
rlabel pdiffusion 115 -2949 115 -2949 0 cellNo=701
rlabel pdiffusion 122 -2949 122 -2949 0 feedthrough
rlabel pdiffusion 129 -2949 129 -2949 0 feedthrough
rlabel pdiffusion 136 -2949 136 -2949 0 feedthrough
rlabel pdiffusion 143 -2949 143 -2949 0 feedthrough
rlabel pdiffusion 150 -2949 150 -2949 0 feedthrough
rlabel pdiffusion 157 -2949 157 -2949 0 cellNo=801
rlabel pdiffusion 164 -2949 164 -2949 0 feedthrough
rlabel pdiffusion 171 -2949 171 -2949 0 feedthrough
rlabel pdiffusion 178 -2949 178 -2949 0 cellNo=491
rlabel pdiffusion 185 -2949 185 -2949 0 feedthrough
rlabel pdiffusion 192 -2949 192 -2949 0 feedthrough
rlabel pdiffusion 199 -2949 199 -2949 0 feedthrough
rlabel pdiffusion 206 -2949 206 -2949 0 feedthrough
rlabel pdiffusion 213 -2949 213 -2949 0 feedthrough
rlabel pdiffusion 220 -2949 220 -2949 0 feedthrough
rlabel pdiffusion 227 -2949 227 -2949 0 feedthrough
rlabel pdiffusion 234 -2949 234 -2949 0 feedthrough
rlabel pdiffusion 241 -2949 241 -2949 0 feedthrough
rlabel pdiffusion 248 -2949 248 -2949 0 cellNo=905
rlabel pdiffusion 255 -2949 255 -2949 0 cellNo=333
rlabel pdiffusion 262 -2949 262 -2949 0 cellNo=526
rlabel pdiffusion 269 -2949 269 -2949 0 feedthrough
rlabel pdiffusion 276 -2949 276 -2949 0 feedthrough
rlabel pdiffusion 283 -2949 283 -2949 0 feedthrough
rlabel pdiffusion 290 -2949 290 -2949 0 feedthrough
rlabel pdiffusion 297 -2949 297 -2949 0 feedthrough
rlabel pdiffusion 304 -2949 304 -2949 0 feedthrough
rlabel pdiffusion 311 -2949 311 -2949 0 feedthrough
rlabel pdiffusion 318 -2949 318 -2949 0 feedthrough
rlabel pdiffusion 325 -2949 325 -2949 0 feedthrough
rlabel pdiffusion 332 -2949 332 -2949 0 feedthrough
rlabel pdiffusion 339 -2949 339 -2949 0 feedthrough
rlabel pdiffusion 346 -2949 346 -2949 0 feedthrough
rlabel pdiffusion 353 -2949 353 -2949 0 feedthrough
rlabel pdiffusion 360 -2949 360 -2949 0 feedthrough
rlabel pdiffusion 367 -2949 367 -2949 0 feedthrough
rlabel pdiffusion 374 -2949 374 -2949 0 cellNo=510
rlabel pdiffusion 381 -2949 381 -2949 0 feedthrough
rlabel pdiffusion 388 -2949 388 -2949 0 feedthrough
rlabel pdiffusion 395 -2949 395 -2949 0 feedthrough
rlabel pdiffusion 402 -2949 402 -2949 0 cellNo=885
rlabel pdiffusion 409 -2949 409 -2949 0 cellNo=203
rlabel pdiffusion 416 -2949 416 -2949 0 feedthrough
rlabel pdiffusion 423 -2949 423 -2949 0 feedthrough
rlabel pdiffusion 430 -2949 430 -2949 0 feedthrough
rlabel pdiffusion 437 -2949 437 -2949 0 feedthrough
rlabel pdiffusion 444 -2949 444 -2949 0 feedthrough
rlabel pdiffusion 451 -2949 451 -2949 0 feedthrough
rlabel pdiffusion 458 -2949 458 -2949 0 feedthrough
rlabel pdiffusion 465 -2949 465 -2949 0 feedthrough
rlabel pdiffusion 472 -2949 472 -2949 0 cellNo=469
rlabel pdiffusion 479 -2949 479 -2949 0 cellNo=914
rlabel pdiffusion 486 -2949 486 -2949 0 feedthrough
rlabel pdiffusion 493 -2949 493 -2949 0 feedthrough
rlabel pdiffusion 500 -2949 500 -2949 0 cellNo=374
rlabel pdiffusion 507 -2949 507 -2949 0 feedthrough
rlabel pdiffusion 514 -2949 514 -2949 0 feedthrough
rlabel pdiffusion 521 -2949 521 -2949 0 feedthrough
rlabel pdiffusion 528 -2949 528 -2949 0 feedthrough
rlabel pdiffusion 535 -2949 535 -2949 0 feedthrough
rlabel pdiffusion 542 -2949 542 -2949 0 feedthrough
rlabel pdiffusion 549 -2949 549 -2949 0 feedthrough
rlabel pdiffusion 556 -2949 556 -2949 0 feedthrough
rlabel pdiffusion 563 -2949 563 -2949 0 cellNo=541
rlabel pdiffusion 570 -2949 570 -2949 0 feedthrough
rlabel pdiffusion 577 -2949 577 -2949 0 feedthrough
rlabel pdiffusion 584 -2949 584 -2949 0 feedthrough
rlabel pdiffusion 591 -2949 591 -2949 0 feedthrough
rlabel pdiffusion 598 -2949 598 -2949 0 feedthrough
rlabel pdiffusion 605 -2949 605 -2949 0 cellNo=459
rlabel pdiffusion 612 -2949 612 -2949 0 feedthrough
rlabel pdiffusion 619 -2949 619 -2949 0 feedthrough
rlabel pdiffusion 626 -2949 626 -2949 0 feedthrough
rlabel pdiffusion 633 -2949 633 -2949 0 cellNo=753
rlabel pdiffusion 640 -2949 640 -2949 0 feedthrough
rlabel pdiffusion 647 -2949 647 -2949 0 feedthrough
rlabel pdiffusion 654 -2949 654 -2949 0 feedthrough
rlabel pdiffusion 661 -2949 661 -2949 0 feedthrough
rlabel pdiffusion 668 -2949 668 -2949 0 cellNo=723
rlabel pdiffusion 675 -2949 675 -2949 0 feedthrough
rlabel pdiffusion 682 -2949 682 -2949 0 feedthrough
rlabel pdiffusion 689 -2949 689 -2949 0 cellNo=986
rlabel pdiffusion 696 -2949 696 -2949 0 feedthrough
rlabel pdiffusion 703 -2949 703 -2949 0 cellNo=543
rlabel pdiffusion 710 -2949 710 -2949 0 feedthrough
rlabel pdiffusion 717 -2949 717 -2949 0 feedthrough
rlabel pdiffusion 724 -2949 724 -2949 0 feedthrough
rlabel pdiffusion 731 -2949 731 -2949 0 cellNo=582
rlabel pdiffusion 738 -2949 738 -2949 0 feedthrough
rlabel pdiffusion 745 -2949 745 -2949 0 feedthrough
rlabel pdiffusion 752 -2949 752 -2949 0 feedthrough
rlabel pdiffusion 759 -2949 759 -2949 0 cellNo=757
rlabel pdiffusion 766 -2949 766 -2949 0 feedthrough
rlabel pdiffusion 773 -2949 773 -2949 0 feedthrough
rlabel pdiffusion 780 -2949 780 -2949 0 feedthrough
rlabel pdiffusion 787 -2949 787 -2949 0 feedthrough
rlabel pdiffusion 794 -2949 794 -2949 0 feedthrough
rlabel pdiffusion 801 -2949 801 -2949 0 feedthrough
rlabel pdiffusion 808 -2949 808 -2949 0 feedthrough
rlabel pdiffusion 815 -2949 815 -2949 0 feedthrough
rlabel pdiffusion 822 -2949 822 -2949 0 feedthrough
rlabel pdiffusion 829 -2949 829 -2949 0 feedthrough
rlabel pdiffusion 836 -2949 836 -2949 0 feedthrough
rlabel pdiffusion 843 -2949 843 -2949 0 feedthrough
rlabel pdiffusion 850 -2949 850 -2949 0 feedthrough
rlabel pdiffusion 857 -2949 857 -2949 0 feedthrough
rlabel pdiffusion 864 -2949 864 -2949 0 cellNo=946
rlabel pdiffusion 871 -2949 871 -2949 0 feedthrough
rlabel pdiffusion 878 -2949 878 -2949 0 feedthrough
rlabel pdiffusion 885 -2949 885 -2949 0 feedthrough
rlabel pdiffusion 892 -2949 892 -2949 0 feedthrough
rlabel pdiffusion 899 -2949 899 -2949 0 feedthrough
rlabel pdiffusion 906 -2949 906 -2949 0 feedthrough
rlabel pdiffusion 913 -2949 913 -2949 0 cellNo=5
rlabel pdiffusion 920 -2949 920 -2949 0 feedthrough
rlabel pdiffusion 927 -2949 927 -2949 0 cellNo=4
rlabel pdiffusion 934 -2949 934 -2949 0 cellNo=641
rlabel pdiffusion 941 -2949 941 -2949 0 feedthrough
rlabel pdiffusion 948 -2949 948 -2949 0 feedthrough
rlabel pdiffusion 955 -2949 955 -2949 0 feedthrough
rlabel pdiffusion 962 -2949 962 -2949 0 feedthrough
rlabel pdiffusion 969 -2949 969 -2949 0 feedthrough
rlabel pdiffusion 976 -2949 976 -2949 0 feedthrough
rlabel pdiffusion 983 -2949 983 -2949 0 feedthrough
rlabel pdiffusion 990 -2949 990 -2949 0 feedthrough
rlabel pdiffusion 997 -2949 997 -2949 0 cellNo=521
rlabel pdiffusion 1004 -2949 1004 -2949 0 feedthrough
rlabel pdiffusion 1011 -2949 1011 -2949 0 feedthrough
rlabel pdiffusion 1018 -2949 1018 -2949 0 cellNo=929
rlabel pdiffusion 1025 -2949 1025 -2949 0 cellNo=876
rlabel pdiffusion 1032 -2949 1032 -2949 0 feedthrough
rlabel pdiffusion 1039 -2949 1039 -2949 0 feedthrough
rlabel pdiffusion 1046 -2949 1046 -2949 0 feedthrough
rlabel pdiffusion 1053 -2949 1053 -2949 0 feedthrough
rlabel pdiffusion 1060 -2949 1060 -2949 0 feedthrough
rlabel pdiffusion 1067 -2949 1067 -2949 0 feedthrough
rlabel pdiffusion 1074 -2949 1074 -2949 0 feedthrough
rlabel pdiffusion 1081 -2949 1081 -2949 0 feedthrough
rlabel pdiffusion 1088 -2949 1088 -2949 0 feedthrough
rlabel pdiffusion 1095 -2949 1095 -2949 0 feedthrough
rlabel pdiffusion 1102 -2949 1102 -2949 0 feedthrough
rlabel pdiffusion 1109 -2949 1109 -2949 0 feedthrough
rlabel pdiffusion 1116 -2949 1116 -2949 0 feedthrough
rlabel pdiffusion 1123 -2949 1123 -2949 0 feedthrough
rlabel pdiffusion 1130 -2949 1130 -2949 0 feedthrough
rlabel pdiffusion 1137 -2949 1137 -2949 0 feedthrough
rlabel pdiffusion 1144 -2949 1144 -2949 0 feedthrough
rlabel pdiffusion 1151 -2949 1151 -2949 0 feedthrough
rlabel pdiffusion 1158 -2949 1158 -2949 0 feedthrough
rlabel pdiffusion 1165 -2949 1165 -2949 0 feedthrough
rlabel pdiffusion 1172 -2949 1172 -2949 0 feedthrough
rlabel pdiffusion 1179 -2949 1179 -2949 0 feedthrough
rlabel pdiffusion 1186 -2949 1186 -2949 0 feedthrough
rlabel pdiffusion 1193 -2949 1193 -2949 0 feedthrough
rlabel pdiffusion 1200 -2949 1200 -2949 0 cellNo=919
rlabel pdiffusion 1207 -2949 1207 -2949 0 feedthrough
rlabel pdiffusion 1214 -2949 1214 -2949 0 feedthrough
rlabel pdiffusion 1221 -2949 1221 -2949 0 feedthrough
rlabel pdiffusion 1228 -2949 1228 -2949 0 feedthrough
rlabel pdiffusion 1235 -2949 1235 -2949 0 feedthrough
rlabel pdiffusion 1242 -2949 1242 -2949 0 feedthrough
rlabel pdiffusion 1249 -2949 1249 -2949 0 feedthrough
rlabel pdiffusion 1256 -2949 1256 -2949 0 feedthrough
rlabel pdiffusion 1263 -2949 1263 -2949 0 feedthrough
rlabel pdiffusion 1270 -2949 1270 -2949 0 feedthrough
rlabel pdiffusion 1277 -2949 1277 -2949 0 feedthrough
rlabel pdiffusion 1284 -2949 1284 -2949 0 feedthrough
rlabel pdiffusion 1291 -2949 1291 -2949 0 feedthrough
rlabel pdiffusion 1298 -2949 1298 -2949 0 feedthrough
rlabel pdiffusion 1305 -2949 1305 -2949 0 feedthrough
rlabel pdiffusion 1312 -2949 1312 -2949 0 feedthrough
rlabel pdiffusion 1319 -2949 1319 -2949 0 feedthrough
rlabel pdiffusion 1326 -2949 1326 -2949 0 feedthrough
rlabel pdiffusion 1333 -2949 1333 -2949 0 feedthrough
rlabel pdiffusion 1340 -2949 1340 -2949 0 feedthrough
rlabel pdiffusion 1347 -2949 1347 -2949 0 feedthrough
rlabel pdiffusion 1354 -2949 1354 -2949 0 feedthrough
rlabel pdiffusion 1361 -2949 1361 -2949 0 feedthrough
rlabel pdiffusion 1368 -2949 1368 -2949 0 feedthrough
rlabel pdiffusion 1375 -2949 1375 -2949 0 feedthrough
rlabel pdiffusion 1382 -2949 1382 -2949 0 feedthrough
rlabel pdiffusion 1389 -2949 1389 -2949 0 feedthrough
rlabel pdiffusion 1396 -2949 1396 -2949 0 feedthrough
rlabel pdiffusion 1403 -2949 1403 -2949 0 feedthrough
rlabel pdiffusion 1410 -2949 1410 -2949 0 feedthrough
rlabel pdiffusion 1417 -2949 1417 -2949 0 feedthrough
rlabel pdiffusion 1424 -2949 1424 -2949 0 feedthrough
rlabel pdiffusion 1431 -2949 1431 -2949 0 feedthrough
rlabel pdiffusion 1438 -2949 1438 -2949 0 feedthrough
rlabel pdiffusion 1445 -2949 1445 -2949 0 cellNo=684
rlabel pdiffusion 1452 -2949 1452 -2949 0 feedthrough
rlabel pdiffusion 1459 -2949 1459 -2949 0 feedthrough
rlabel pdiffusion 1466 -2949 1466 -2949 0 feedthrough
rlabel pdiffusion 1480 -2949 1480 -2949 0 feedthrough
rlabel pdiffusion 1487 -2949 1487 -2949 0 feedthrough
rlabel pdiffusion 1494 -2949 1494 -2949 0 feedthrough
rlabel pdiffusion 1501 -2949 1501 -2949 0 feedthrough
rlabel pdiffusion 3 -3068 3 -3068 0 cellNo=1171
rlabel pdiffusion 10 -3068 10 -3068 0 cellNo=1182
rlabel pdiffusion 17 -3068 17 -3068 0 cellNo=1192
rlabel pdiffusion 38 -3068 38 -3068 0 feedthrough
rlabel pdiffusion 45 -3068 45 -3068 0 feedthrough
rlabel pdiffusion 52 -3068 52 -3068 0 feedthrough
rlabel pdiffusion 59 -3068 59 -3068 0 feedthrough
rlabel pdiffusion 66 -3068 66 -3068 0 feedthrough
rlabel pdiffusion 73 -3068 73 -3068 0 feedthrough
rlabel pdiffusion 80 -3068 80 -3068 0 feedthrough
rlabel pdiffusion 87 -3068 87 -3068 0 feedthrough
rlabel pdiffusion 94 -3068 94 -3068 0 cellNo=691
rlabel pdiffusion 101 -3068 101 -3068 0 feedthrough
rlabel pdiffusion 108 -3068 108 -3068 0 feedthrough
rlabel pdiffusion 115 -3068 115 -3068 0 feedthrough
rlabel pdiffusion 122 -3068 122 -3068 0 cellNo=124
rlabel pdiffusion 129 -3068 129 -3068 0 feedthrough
rlabel pdiffusion 136 -3068 136 -3068 0 feedthrough
rlabel pdiffusion 143 -3068 143 -3068 0 feedthrough
rlabel pdiffusion 150 -3068 150 -3068 0 feedthrough
rlabel pdiffusion 157 -3068 157 -3068 0 feedthrough
rlabel pdiffusion 164 -3068 164 -3068 0 feedthrough
rlabel pdiffusion 171 -3068 171 -3068 0 feedthrough
rlabel pdiffusion 178 -3068 178 -3068 0 cellNo=259
rlabel pdiffusion 185 -3068 185 -3068 0 feedthrough
rlabel pdiffusion 192 -3068 192 -3068 0 feedthrough
rlabel pdiffusion 199 -3068 199 -3068 0 cellNo=525
rlabel pdiffusion 206 -3068 206 -3068 0 feedthrough
rlabel pdiffusion 213 -3068 213 -3068 0 feedthrough
rlabel pdiffusion 220 -3068 220 -3068 0 cellNo=906
rlabel pdiffusion 227 -3068 227 -3068 0 feedthrough
rlabel pdiffusion 234 -3068 234 -3068 0 feedthrough
rlabel pdiffusion 241 -3068 241 -3068 0 cellNo=971
rlabel pdiffusion 248 -3068 248 -3068 0 cellNo=355
rlabel pdiffusion 255 -3068 255 -3068 0 feedthrough
rlabel pdiffusion 262 -3068 262 -3068 0 cellNo=856
rlabel pdiffusion 269 -3068 269 -3068 0 feedthrough
rlabel pdiffusion 276 -3068 276 -3068 0 feedthrough
rlabel pdiffusion 283 -3068 283 -3068 0 feedthrough
rlabel pdiffusion 290 -3068 290 -3068 0 feedthrough
rlabel pdiffusion 297 -3068 297 -3068 0 cellNo=39
rlabel pdiffusion 304 -3068 304 -3068 0 feedthrough
rlabel pdiffusion 311 -3068 311 -3068 0 feedthrough
rlabel pdiffusion 318 -3068 318 -3068 0 feedthrough
rlabel pdiffusion 325 -3068 325 -3068 0 feedthrough
rlabel pdiffusion 332 -3068 332 -3068 0 feedthrough
rlabel pdiffusion 339 -3068 339 -3068 0 feedthrough
rlabel pdiffusion 346 -3068 346 -3068 0 feedthrough
rlabel pdiffusion 353 -3068 353 -3068 0 cellNo=745
rlabel pdiffusion 360 -3068 360 -3068 0 feedthrough
rlabel pdiffusion 367 -3068 367 -3068 0 feedthrough
rlabel pdiffusion 374 -3068 374 -3068 0 feedthrough
rlabel pdiffusion 381 -3068 381 -3068 0 feedthrough
rlabel pdiffusion 388 -3068 388 -3068 0 feedthrough
rlabel pdiffusion 395 -3068 395 -3068 0 feedthrough
rlabel pdiffusion 402 -3068 402 -3068 0 feedthrough
rlabel pdiffusion 409 -3068 409 -3068 0 cellNo=122
rlabel pdiffusion 416 -3068 416 -3068 0 feedthrough
rlabel pdiffusion 423 -3068 423 -3068 0 feedthrough
rlabel pdiffusion 430 -3068 430 -3068 0 feedthrough
rlabel pdiffusion 437 -3068 437 -3068 0 feedthrough
rlabel pdiffusion 444 -3068 444 -3068 0 feedthrough
rlabel pdiffusion 451 -3068 451 -3068 0 feedthrough
rlabel pdiffusion 458 -3068 458 -3068 0 feedthrough
rlabel pdiffusion 465 -3068 465 -3068 0 feedthrough
rlabel pdiffusion 472 -3068 472 -3068 0 feedthrough
rlabel pdiffusion 479 -3068 479 -3068 0 feedthrough
rlabel pdiffusion 486 -3068 486 -3068 0 feedthrough
rlabel pdiffusion 493 -3068 493 -3068 0 feedthrough
rlabel pdiffusion 500 -3068 500 -3068 0 feedthrough
rlabel pdiffusion 507 -3068 507 -3068 0 feedthrough
rlabel pdiffusion 514 -3068 514 -3068 0 feedthrough
rlabel pdiffusion 521 -3068 521 -3068 0 cellNo=352
rlabel pdiffusion 528 -3068 528 -3068 0 feedthrough
rlabel pdiffusion 535 -3068 535 -3068 0 feedthrough
rlabel pdiffusion 542 -3068 542 -3068 0 feedthrough
rlabel pdiffusion 549 -3068 549 -3068 0 feedthrough
rlabel pdiffusion 556 -3068 556 -3068 0 feedthrough
rlabel pdiffusion 563 -3068 563 -3068 0 feedthrough
rlabel pdiffusion 570 -3068 570 -3068 0 feedthrough
rlabel pdiffusion 577 -3068 577 -3068 0 feedthrough
rlabel pdiffusion 584 -3068 584 -3068 0 feedthrough
rlabel pdiffusion 591 -3068 591 -3068 0 feedthrough
rlabel pdiffusion 598 -3068 598 -3068 0 feedthrough
rlabel pdiffusion 605 -3068 605 -3068 0 cellNo=310
rlabel pdiffusion 612 -3068 612 -3068 0 feedthrough
rlabel pdiffusion 619 -3068 619 -3068 0 cellNo=848
rlabel pdiffusion 626 -3068 626 -3068 0 feedthrough
rlabel pdiffusion 633 -3068 633 -3068 0 feedthrough
rlabel pdiffusion 640 -3068 640 -3068 0 cellNo=760
rlabel pdiffusion 647 -3068 647 -3068 0 feedthrough
rlabel pdiffusion 654 -3068 654 -3068 0 feedthrough
rlabel pdiffusion 661 -3068 661 -3068 0 feedthrough
rlabel pdiffusion 668 -3068 668 -3068 0 feedthrough
rlabel pdiffusion 675 -3068 675 -3068 0 feedthrough
rlabel pdiffusion 682 -3068 682 -3068 0 cellNo=825
rlabel pdiffusion 689 -3068 689 -3068 0 feedthrough
rlabel pdiffusion 696 -3068 696 -3068 0 feedthrough
rlabel pdiffusion 703 -3068 703 -3068 0 cellNo=565
rlabel pdiffusion 710 -3068 710 -3068 0 feedthrough
rlabel pdiffusion 717 -3068 717 -3068 0 feedthrough
rlabel pdiffusion 724 -3068 724 -3068 0 feedthrough
rlabel pdiffusion 731 -3068 731 -3068 0 feedthrough
rlabel pdiffusion 738 -3068 738 -3068 0 cellNo=104
rlabel pdiffusion 745 -3068 745 -3068 0 feedthrough
rlabel pdiffusion 752 -3068 752 -3068 0 feedthrough
rlabel pdiffusion 759 -3068 759 -3068 0 feedthrough
rlabel pdiffusion 766 -3068 766 -3068 0 feedthrough
rlabel pdiffusion 773 -3068 773 -3068 0 feedthrough
rlabel pdiffusion 780 -3068 780 -3068 0 feedthrough
rlabel pdiffusion 787 -3068 787 -3068 0 feedthrough
rlabel pdiffusion 794 -3068 794 -3068 0 cellNo=537
rlabel pdiffusion 801 -3068 801 -3068 0 feedthrough
rlabel pdiffusion 808 -3068 808 -3068 0 feedthrough
rlabel pdiffusion 815 -3068 815 -3068 0 feedthrough
rlabel pdiffusion 822 -3068 822 -3068 0 feedthrough
rlabel pdiffusion 829 -3068 829 -3068 0 feedthrough
rlabel pdiffusion 836 -3068 836 -3068 0 feedthrough
rlabel pdiffusion 843 -3068 843 -3068 0 feedthrough
rlabel pdiffusion 850 -3068 850 -3068 0 cellNo=231
rlabel pdiffusion 857 -3068 857 -3068 0 feedthrough
rlabel pdiffusion 864 -3068 864 -3068 0 feedthrough
rlabel pdiffusion 871 -3068 871 -3068 0 cellNo=819
rlabel pdiffusion 878 -3068 878 -3068 0 feedthrough
rlabel pdiffusion 885 -3068 885 -3068 0 feedthrough
rlabel pdiffusion 892 -3068 892 -3068 0 feedthrough
rlabel pdiffusion 899 -3068 899 -3068 0 feedthrough
rlabel pdiffusion 906 -3068 906 -3068 0 feedthrough
rlabel pdiffusion 913 -3068 913 -3068 0 feedthrough
rlabel pdiffusion 920 -3068 920 -3068 0 cellNo=909
rlabel pdiffusion 927 -3068 927 -3068 0 cellNo=881
rlabel pdiffusion 934 -3068 934 -3068 0 feedthrough
rlabel pdiffusion 941 -3068 941 -3068 0 feedthrough
rlabel pdiffusion 948 -3068 948 -3068 0 feedthrough
rlabel pdiffusion 955 -3068 955 -3068 0 feedthrough
rlabel pdiffusion 962 -3068 962 -3068 0 cellNo=351
rlabel pdiffusion 969 -3068 969 -3068 0 feedthrough
rlabel pdiffusion 976 -3068 976 -3068 0 feedthrough
rlabel pdiffusion 983 -3068 983 -3068 0 feedthrough
rlabel pdiffusion 990 -3068 990 -3068 0 feedthrough
rlabel pdiffusion 997 -3068 997 -3068 0 cellNo=935
rlabel pdiffusion 1004 -3068 1004 -3068 0 feedthrough
rlabel pdiffusion 1011 -3068 1011 -3068 0 feedthrough
rlabel pdiffusion 1018 -3068 1018 -3068 0 feedthrough
rlabel pdiffusion 1025 -3068 1025 -3068 0 feedthrough
rlabel pdiffusion 1032 -3068 1032 -3068 0 feedthrough
rlabel pdiffusion 1039 -3068 1039 -3068 0 feedthrough
rlabel pdiffusion 1046 -3068 1046 -3068 0 feedthrough
rlabel pdiffusion 1053 -3068 1053 -3068 0 feedthrough
rlabel pdiffusion 1060 -3068 1060 -3068 0 cellNo=949
rlabel pdiffusion 1067 -3068 1067 -3068 0 feedthrough
rlabel pdiffusion 1074 -3068 1074 -3068 0 feedthrough
rlabel pdiffusion 1081 -3068 1081 -3068 0 feedthrough
rlabel pdiffusion 1088 -3068 1088 -3068 0 cellNo=593
rlabel pdiffusion 1095 -3068 1095 -3068 0 feedthrough
rlabel pdiffusion 1102 -3068 1102 -3068 0 feedthrough
rlabel pdiffusion 1109 -3068 1109 -3068 0 feedthrough
rlabel pdiffusion 1116 -3068 1116 -3068 0 feedthrough
rlabel pdiffusion 1123 -3068 1123 -3068 0 feedthrough
rlabel pdiffusion 1130 -3068 1130 -3068 0 feedthrough
rlabel pdiffusion 1137 -3068 1137 -3068 0 feedthrough
rlabel pdiffusion 1144 -3068 1144 -3068 0 feedthrough
rlabel pdiffusion 1151 -3068 1151 -3068 0 feedthrough
rlabel pdiffusion 1158 -3068 1158 -3068 0 feedthrough
rlabel pdiffusion 1165 -3068 1165 -3068 0 feedthrough
rlabel pdiffusion 1172 -3068 1172 -3068 0 feedthrough
rlabel pdiffusion 1179 -3068 1179 -3068 0 feedthrough
rlabel pdiffusion 1186 -3068 1186 -3068 0 feedthrough
rlabel pdiffusion 1193 -3068 1193 -3068 0 feedthrough
rlabel pdiffusion 1200 -3068 1200 -3068 0 feedthrough
rlabel pdiffusion 1207 -3068 1207 -3068 0 feedthrough
rlabel pdiffusion 1214 -3068 1214 -3068 0 feedthrough
rlabel pdiffusion 1221 -3068 1221 -3068 0 cellNo=768
rlabel pdiffusion 1228 -3068 1228 -3068 0 feedthrough
rlabel pdiffusion 1235 -3068 1235 -3068 0 feedthrough
rlabel pdiffusion 1242 -3068 1242 -3068 0 feedthrough
rlabel pdiffusion 1249 -3068 1249 -3068 0 feedthrough
rlabel pdiffusion 1256 -3068 1256 -3068 0 feedthrough
rlabel pdiffusion 1263 -3068 1263 -3068 0 feedthrough
rlabel pdiffusion 1270 -3068 1270 -3068 0 feedthrough
rlabel pdiffusion 1277 -3068 1277 -3068 0 feedthrough
rlabel pdiffusion 1284 -3068 1284 -3068 0 cellNo=996
rlabel pdiffusion 1291 -3068 1291 -3068 0 feedthrough
rlabel pdiffusion 1298 -3068 1298 -3068 0 feedthrough
rlabel pdiffusion 1305 -3068 1305 -3068 0 feedthrough
rlabel pdiffusion 1312 -3068 1312 -3068 0 feedthrough
rlabel pdiffusion 1319 -3068 1319 -3068 0 feedthrough
rlabel pdiffusion 1326 -3068 1326 -3068 0 feedthrough
rlabel pdiffusion 1333 -3068 1333 -3068 0 feedthrough
rlabel pdiffusion 1340 -3068 1340 -3068 0 feedthrough
rlabel pdiffusion 1347 -3068 1347 -3068 0 feedthrough
rlabel pdiffusion 1375 -3068 1375 -3068 0 feedthrough
rlabel pdiffusion 1382 -3068 1382 -3068 0 feedthrough
rlabel pdiffusion 1417 -3068 1417 -3068 0 feedthrough
rlabel pdiffusion 1459 -3068 1459 -3068 0 feedthrough
rlabel pdiffusion 1466 -3068 1466 -3068 0 feedthrough
rlabel pdiffusion 1473 -3068 1473 -3068 0 feedthrough
rlabel pdiffusion 3 -3157 3 -3157 0 cellNo=1181
rlabel pdiffusion 10 -3157 10 -3157 0 cellNo=1191
rlabel pdiffusion 80 -3157 80 -3157 0 feedthrough
rlabel pdiffusion 87 -3157 87 -3157 0 feedthrough
rlabel pdiffusion 94 -3157 94 -3157 0 feedthrough
rlabel pdiffusion 101 -3157 101 -3157 0 feedthrough
rlabel pdiffusion 108 -3157 108 -3157 0 feedthrough
rlabel pdiffusion 115 -3157 115 -3157 0 feedthrough
rlabel pdiffusion 122 -3157 122 -3157 0 feedthrough
rlabel pdiffusion 129 -3157 129 -3157 0 feedthrough
rlabel pdiffusion 136 -3157 136 -3157 0 feedthrough
rlabel pdiffusion 143 -3157 143 -3157 0 feedthrough
rlabel pdiffusion 150 -3157 150 -3157 0 feedthrough
rlabel pdiffusion 157 -3157 157 -3157 0 feedthrough
rlabel pdiffusion 164 -3157 164 -3157 0 feedthrough
rlabel pdiffusion 171 -3157 171 -3157 0 feedthrough
rlabel pdiffusion 178 -3157 178 -3157 0 feedthrough
rlabel pdiffusion 185 -3157 185 -3157 0 cellNo=207
rlabel pdiffusion 192 -3157 192 -3157 0 feedthrough
rlabel pdiffusion 199 -3157 199 -3157 0 feedthrough
rlabel pdiffusion 206 -3157 206 -3157 0 feedthrough
rlabel pdiffusion 213 -3157 213 -3157 0 cellNo=871
rlabel pdiffusion 220 -3157 220 -3157 0 cellNo=192
rlabel pdiffusion 227 -3157 227 -3157 0 feedthrough
rlabel pdiffusion 234 -3157 234 -3157 0 feedthrough
rlabel pdiffusion 241 -3157 241 -3157 0 feedthrough
rlabel pdiffusion 248 -3157 248 -3157 0 feedthrough
rlabel pdiffusion 255 -3157 255 -3157 0 feedthrough
rlabel pdiffusion 262 -3157 262 -3157 0 feedthrough
rlabel pdiffusion 269 -3157 269 -3157 0 feedthrough
rlabel pdiffusion 276 -3157 276 -3157 0 feedthrough
rlabel pdiffusion 283 -3157 283 -3157 0 feedthrough
rlabel pdiffusion 290 -3157 290 -3157 0 feedthrough
rlabel pdiffusion 297 -3157 297 -3157 0 feedthrough
rlabel pdiffusion 304 -3157 304 -3157 0 cellNo=186
rlabel pdiffusion 311 -3157 311 -3157 0 feedthrough
rlabel pdiffusion 318 -3157 318 -3157 0 feedthrough
rlabel pdiffusion 325 -3157 325 -3157 0 feedthrough
rlabel pdiffusion 332 -3157 332 -3157 0 feedthrough
rlabel pdiffusion 339 -3157 339 -3157 0 feedthrough
rlabel pdiffusion 346 -3157 346 -3157 0 feedthrough
rlabel pdiffusion 353 -3157 353 -3157 0 feedthrough
rlabel pdiffusion 360 -3157 360 -3157 0 cellNo=44
rlabel pdiffusion 367 -3157 367 -3157 0 feedthrough
rlabel pdiffusion 374 -3157 374 -3157 0 feedthrough
rlabel pdiffusion 381 -3157 381 -3157 0 feedthrough
rlabel pdiffusion 388 -3157 388 -3157 0 feedthrough
rlabel pdiffusion 395 -3157 395 -3157 0 feedthrough
rlabel pdiffusion 402 -3157 402 -3157 0 feedthrough
rlabel pdiffusion 409 -3157 409 -3157 0 feedthrough
rlabel pdiffusion 416 -3157 416 -3157 0 feedthrough
rlabel pdiffusion 423 -3157 423 -3157 0 feedthrough
rlabel pdiffusion 430 -3157 430 -3157 0 cellNo=920
rlabel pdiffusion 437 -3157 437 -3157 0 feedthrough
rlabel pdiffusion 444 -3157 444 -3157 0 feedthrough
rlabel pdiffusion 451 -3157 451 -3157 0 feedthrough
rlabel pdiffusion 458 -3157 458 -3157 0 feedthrough
rlabel pdiffusion 465 -3157 465 -3157 0 feedthrough
rlabel pdiffusion 472 -3157 472 -3157 0 feedthrough
rlabel pdiffusion 479 -3157 479 -3157 0 feedthrough
rlabel pdiffusion 486 -3157 486 -3157 0 feedthrough
rlabel pdiffusion 493 -3157 493 -3157 0 feedthrough
rlabel pdiffusion 500 -3157 500 -3157 0 feedthrough
rlabel pdiffusion 507 -3157 507 -3157 0 feedthrough
rlabel pdiffusion 514 -3157 514 -3157 0 feedthrough
rlabel pdiffusion 521 -3157 521 -3157 0 feedthrough
rlabel pdiffusion 528 -3157 528 -3157 0 feedthrough
rlabel pdiffusion 535 -3157 535 -3157 0 feedthrough
rlabel pdiffusion 542 -3157 542 -3157 0 feedthrough
rlabel pdiffusion 549 -3157 549 -3157 0 feedthrough
rlabel pdiffusion 556 -3157 556 -3157 0 feedthrough
rlabel pdiffusion 563 -3157 563 -3157 0 feedthrough
rlabel pdiffusion 570 -3157 570 -3157 0 feedthrough
rlabel pdiffusion 577 -3157 577 -3157 0 cellNo=748
rlabel pdiffusion 584 -3157 584 -3157 0 feedthrough
rlabel pdiffusion 591 -3157 591 -3157 0 feedthrough
rlabel pdiffusion 598 -3157 598 -3157 0 feedthrough
rlabel pdiffusion 605 -3157 605 -3157 0 cellNo=759
rlabel pdiffusion 612 -3157 612 -3157 0 feedthrough
rlabel pdiffusion 619 -3157 619 -3157 0 cellNo=320
rlabel pdiffusion 626 -3157 626 -3157 0 feedthrough
rlabel pdiffusion 633 -3157 633 -3157 0 cellNo=92
rlabel pdiffusion 640 -3157 640 -3157 0 feedthrough
rlabel pdiffusion 647 -3157 647 -3157 0 feedthrough
rlabel pdiffusion 654 -3157 654 -3157 0 cellNo=761
rlabel pdiffusion 661 -3157 661 -3157 0 cellNo=377
rlabel pdiffusion 668 -3157 668 -3157 0 feedthrough
rlabel pdiffusion 675 -3157 675 -3157 0 feedthrough
rlabel pdiffusion 682 -3157 682 -3157 0 feedthrough
rlabel pdiffusion 689 -3157 689 -3157 0 cellNo=474
rlabel pdiffusion 696 -3157 696 -3157 0 feedthrough
rlabel pdiffusion 703 -3157 703 -3157 0 cellNo=858
rlabel pdiffusion 710 -3157 710 -3157 0 feedthrough
rlabel pdiffusion 717 -3157 717 -3157 0 feedthrough
rlabel pdiffusion 724 -3157 724 -3157 0 feedthrough
rlabel pdiffusion 731 -3157 731 -3157 0 cellNo=275
rlabel pdiffusion 738 -3157 738 -3157 0 feedthrough
rlabel pdiffusion 745 -3157 745 -3157 0 feedthrough
rlabel pdiffusion 752 -3157 752 -3157 0 feedthrough
rlabel pdiffusion 759 -3157 759 -3157 0 feedthrough
rlabel pdiffusion 766 -3157 766 -3157 0 feedthrough
rlabel pdiffusion 773 -3157 773 -3157 0 cellNo=199
rlabel pdiffusion 780 -3157 780 -3157 0 cellNo=152
rlabel pdiffusion 787 -3157 787 -3157 0 feedthrough
rlabel pdiffusion 794 -3157 794 -3157 0 feedthrough
rlabel pdiffusion 801 -3157 801 -3157 0 feedthrough
rlabel pdiffusion 808 -3157 808 -3157 0 feedthrough
rlabel pdiffusion 815 -3157 815 -3157 0 feedthrough
rlabel pdiffusion 822 -3157 822 -3157 0 feedthrough
rlabel pdiffusion 829 -3157 829 -3157 0 feedthrough
rlabel pdiffusion 836 -3157 836 -3157 0 feedthrough
rlabel pdiffusion 843 -3157 843 -3157 0 cellNo=393
rlabel pdiffusion 850 -3157 850 -3157 0 feedthrough
rlabel pdiffusion 857 -3157 857 -3157 0 cellNo=568
rlabel pdiffusion 864 -3157 864 -3157 0 feedthrough
rlabel pdiffusion 871 -3157 871 -3157 0 feedthrough
rlabel pdiffusion 878 -3157 878 -3157 0 cellNo=447
rlabel pdiffusion 885 -3157 885 -3157 0 feedthrough
rlabel pdiffusion 892 -3157 892 -3157 0 feedthrough
rlabel pdiffusion 899 -3157 899 -3157 0 feedthrough
rlabel pdiffusion 906 -3157 906 -3157 0 feedthrough
rlabel pdiffusion 913 -3157 913 -3157 0 feedthrough
rlabel pdiffusion 920 -3157 920 -3157 0 feedthrough
rlabel pdiffusion 927 -3157 927 -3157 0 feedthrough
rlabel pdiffusion 934 -3157 934 -3157 0 feedthrough
rlabel pdiffusion 941 -3157 941 -3157 0 feedthrough
rlabel pdiffusion 948 -3157 948 -3157 0 feedthrough
rlabel pdiffusion 955 -3157 955 -3157 0 feedthrough
rlabel pdiffusion 962 -3157 962 -3157 0 cellNo=676
rlabel pdiffusion 969 -3157 969 -3157 0 feedthrough
rlabel pdiffusion 976 -3157 976 -3157 0 feedthrough
rlabel pdiffusion 983 -3157 983 -3157 0 feedthrough
rlabel pdiffusion 990 -3157 990 -3157 0 feedthrough
rlabel pdiffusion 997 -3157 997 -3157 0 cellNo=467
rlabel pdiffusion 1004 -3157 1004 -3157 0 feedthrough
rlabel pdiffusion 1011 -3157 1011 -3157 0 feedthrough
rlabel pdiffusion 1018 -3157 1018 -3157 0 feedthrough
rlabel pdiffusion 1025 -3157 1025 -3157 0 feedthrough
rlabel pdiffusion 1032 -3157 1032 -3157 0 feedthrough
rlabel pdiffusion 1039 -3157 1039 -3157 0 feedthrough
rlabel pdiffusion 1046 -3157 1046 -3157 0 feedthrough
rlabel pdiffusion 1053 -3157 1053 -3157 0 feedthrough
rlabel pdiffusion 1060 -3157 1060 -3157 0 feedthrough
rlabel pdiffusion 1067 -3157 1067 -3157 0 feedthrough
rlabel pdiffusion 1074 -3157 1074 -3157 0 feedthrough
rlabel pdiffusion 1081 -3157 1081 -3157 0 feedthrough
rlabel pdiffusion 1088 -3157 1088 -3157 0 cellNo=733
rlabel pdiffusion 1095 -3157 1095 -3157 0 feedthrough
rlabel pdiffusion 1102 -3157 1102 -3157 0 feedthrough
rlabel pdiffusion 1109 -3157 1109 -3157 0 feedthrough
rlabel pdiffusion 1116 -3157 1116 -3157 0 feedthrough
rlabel pdiffusion 1123 -3157 1123 -3157 0 feedthrough
rlabel pdiffusion 1130 -3157 1130 -3157 0 feedthrough
rlabel pdiffusion 1137 -3157 1137 -3157 0 feedthrough
rlabel pdiffusion 1144 -3157 1144 -3157 0 feedthrough
rlabel pdiffusion 1151 -3157 1151 -3157 0 feedthrough
rlabel pdiffusion 1158 -3157 1158 -3157 0 feedthrough
rlabel pdiffusion 1165 -3157 1165 -3157 0 feedthrough
rlabel pdiffusion 1172 -3157 1172 -3157 0 feedthrough
rlabel pdiffusion 1179 -3157 1179 -3157 0 feedthrough
rlabel pdiffusion 1186 -3157 1186 -3157 0 cellNo=530
rlabel pdiffusion 1193 -3157 1193 -3157 0 feedthrough
rlabel pdiffusion 1200 -3157 1200 -3157 0 feedthrough
rlabel pdiffusion 1207 -3157 1207 -3157 0 feedthrough
rlabel pdiffusion 1214 -3157 1214 -3157 0 feedthrough
rlabel pdiffusion 1221 -3157 1221 -3157 0 feedthrough
rlabel pdiffusion 1228 -3157 1228 -3157 0 cellNo=253
rlabel pdiffusion 1235 -3157 1235 -3157 0 cellNo=812
rlabel pdiffusion 1242 -3157 1242 -3157 0 cellNo=665
rlabel pdiffusion 1263 -3157 1263 -3157 0 feedthrough
rlabel pdiffusion 1277 -3157 1277 -3157 0 feedthrough
rlabel pdiffusion 1291 -3157 1291 -3157 0 cellNo=754
rlabel pdiffusion 1347 -3157 1347 -3157 0 feedthrough
rlabel pdiffusion 1354 -3157 1354 -3157 0 feedthrough
rlabel pdiffusion 1368 -3157 1368 -3157 0 feedthrough
rlabel pdiffusion 1410 -3157 1410 -3157 0 feedthrough
rlabel pdiffusion 1452 -3157 1452 -3157 0 feedthrough
rlabel pdiffusion 1459 -3157 1459 -3157 0 feedthrough
rlabel pdiffusion 1466 -3157 1466 -3157 0 feedthrough
rlabel pdiffusion 3 -3218 3 -3218 0 cellNo=1190
rlabel pdiffusion 59 -3218 59 -3218 0 feedthrough
rlabel pdiffusion 66 -3218 66 -3218 0 feedthrough
rlabel pdiffusion 73 -3218 73 -3218 0 feedthrough
rlabel pdiffusion 80 -3218 80 -3218 0 feedthrough
rlabel pdiffusion 87 -3218 87 -3218 0 feedthrough
rlabel pdiffusion 94 -3218 94 -3218 0 feedthrough
rlabel pdiffusion 101 -3218 101 -3218 0 feedthrough
rlabel pdiffusion 108 -3218 108 -3218 0 feedthrough
rlabel pdiffusion 115 -3218 115 -3218 0 cellNo=557
rlabel pdiffusion 122 -3218 122 -3218 0 feedthrough
rlabel pdiffusion 129 -3218 129 -3218 0 cellNo=596
rlabel pdiffusion 136 -3218 136 -3218 0 feedthrough
rlabel pdiffusion 143 -3218 143 -3218 0 cellNo=534
rlabel pdiffusion 150 -3218 150 -3218 0 cellNo=379
rlabel pdiffusion 157 -3218 157 -3218 0 feedthrough
rlabel pdiffusion 164 -3218 164 -3218 0 feedthrough
rlabel pdiffusion 171 -3218 171 -3218 0 cellNo=628
rlabel pdiffusion 178 -3218 178 -3218 0 cellNo=282
rlabel pdiffusion 185 -3218 185 -3218 0 feedthrough
rlabel pdiffusion 192 -3218 192 -3218 0 cellNo=506
rlabel pdiffusion 199 -3218 199 -3218 0 cellNo=714
rlabel pdiffusion 206 -3218 206 -3218 0 cellNo=752
rlabel pdiffusion 213 -3218 213 -3218 0 feedthrough
rlabel pdiffusion 220 -3218 220 -3218 0 feedthrough
rlabel pdiffusion 227 -3218 227 -3218 0 feedthrough
rlabel pdiffusion 234 -3218 234 -3218 0 feedthrough
rlabel pdiffusion 241 -3218 241 -3218 0 feedthrough
rlabel pdiffusion 248 -3218 248 -3218 0 cellNo=94
rlabel pdiffusion 255 -3218 255 -3218 0 feedthrough
rlabel pdiffusion 262 -3218 262 -3218 0 cellNo=85
rlabel pdiffusion 269 -3218 269 -3218 0 feedthrough
rlabel pdiffusion 276 -3218 276 -3218 0 feedthrough
rlabel pdiffusion 283 -3218 283 -3218 0 feedthrough
rlabel pdiffusion 290 -3218 290 -3218 0 feedthrough
rlabel pdiffusion 297 -3218 297 -3218 0 feedthrough
rlabel pdiffusion 304 -3218 304 -3218 0 feedthrough
rlabel pdiffusion 311 -3218 311 -3218 0 feedthrough
rlabel pdiffusion 318 -3218 318 -3218 0 feedthrough
rlabel pdiffusion 325 -3218 325 -3218 0 cellNo=656
rlabel pdiffusion 332 -3218 332 -3218 0 feedthrough
rlabel pdiffusion 339 -3218 339 -3218 0 feedthrough
rlabel pdiffusion 346 -3218 346 -3218 0 feedthrough
rlabel pdiffusion 353 -3218 353 -3218 0 feedthrough
rlabel pdiffusion 360 -3218 360 -3218 0 feedthrough
rlabel pdiffusion 367 -3218 367 -3218 0 feedthrough
rlabel pdiffusion 374 -3218 374 -3218 0 feedthrough
rlabel pdiffusion 381 -3218 381 -3218 0 feedthrough
rlabel pdiffusion 388 -3218 388 -3218 0 feedthrough
rlabel pdiffusion 395 -3218 395 -3218 0 feedthrough
rlabel pdiffusion 402 -3218 402 -3218 0 feedthrough
rlabel pdiffusion 409 -3218 409 -3218 0 feedthrough
rlabel pdiffusion 416 -3218 416 -3218 0 feedthrough
rlabel pdiffusion 423 -3218 423 -3218 0 feedthrough
rlabel pdiffusion 430 -3218 430 -3218 0 feedthrough
rlabel pdiffusion 437 -3218 437 -3218 0 feedthrough
rlabel pdiffusion 444 -3218 444 -3218 0 feedthrough
rlabel pdiffusion 451 -3218 451 -3218 0 feedthrough
rlabel pdiffusion 458 -3218 458 -3218 0 feedthrough
rlabel pdiffusion 465 -3218 465 -3218 0 feedthrough
rlabel pdiffusion 472 -3218 472 -3218 0 feedthrough
rlabel pdiffusion 479 -3218 479 -3218 0 feedthrough
rlabel pdiffusion 486 -3218 486 -3218 0 feedthrough
rlabel pdiffusion 493 -3218 493 -3218 0 feedthrough
rlabel pdiffusion 500 -3218 500 -3218 0 feedthrough
rlabel pdiffusion 507 -3218 507 -3218 0 feedthrough
rlabel pdiffusion 514 -3218 514 -3218 0 feedthrough
rlabel pdiffusion 521 -3218 521 -3218 0 feedthrough
rlabel pdiffusion 528 -3218 528 -3218 0 feedthrough
rlabel pdiffusion 535 -3218 535 -3218 0 feedthrough
rlabel pdiffusion 542 -3218 542 -3218 0 feedthrough
rlabel pdiffusion 549 -3218 549 -3218 0 feedthrough
rlabel pdiffusion 556 -3218 556 -3218 0 cellNo=892
rlabel pdiffusion 563 -3218 563 -3218 0 feedthrough
rlabel pdiffusion 570 -3218 570 -3218 0 feedthrough
rlabel pdiffusion 577 -3218 577 -3218 0 cellNo=942
rlabel pdiffusion 584 -3218 584 -3218 0 feedthrough
rlabel pdiffusion 591 -3218 591 -3218 0 feedthrough
rlabel pdiffusion 598 -3218 598 -3218 0 feedthrough
rlabel pdiffusion 605 -3218 605 -3218 0 cellNo=263
rlabel pdiffusion 612 -3218 612 -3218 0 feedthrough
rlabel pdiffusion 619 -3218 619 -3218 0 feedthrough
rlabel pdiffusion 626 -3218 626 -3218 0 cellNo=247
rlabel pdiffusion 633 -3218 633 -3218 0 cellNo=246
rlabel pdiffusion 640 -3218 640 -3218 0 feedthrough
rlabel pdiffusion 647 -3218 647 -3218 0 feedthrough
rlabel pdiffusion 654 -3218 654 -3218 0 feedthrough
rlabel pdiffusion 661 -3218 661 -3218 0 cellNo=791
rlabel pdiffusion 668 -3218 668 -3218 0 feedthrough
rlabel pdiffusion 675 -3218 675 -3218 0 feedthrough
rlabel pdiffusion 682 -3218 682 -3218 0 feedthrough
rlabel pdiffusion 689 -3218 689 -3218 0 feedthrough
rlabel pdiffusion 696 -3218 696 -3218 0 feedthrough
rlabel pdiffusion 703 -3218 703 -3218 0 feedthrough
rlabel pdiffusion 710 -3218 710 -3218 0 feedthrough
rlabel pdiffusion 717 -3218 717 -3218 0 feedthrough
rlabel pdiffusion 724 -3218 724 -3218 0 feedthrough
rlabel pdiffusion 731 -3218 731 -3218 0 feedthrough
rlabel pdiffusion 738 -3218 738 -3218 0 feedthrough
rlabel pdiffusion 745 -3218 745 -3218 0 feedthrough
rlabel pdiffusion 752 -3218 752 -3218 0 feedthrough
rlabel pdiffusion 759 -3218 759 -3218 0 cellNo=922
rlabel pdiffusion 766 -3218 766 -3218 0 feedthrough
rlabel pdiffusion 773 -3218 773 -3218 0 feedthrough
rlabel pdiffusion 780 -3218 780 -3218 0 feedthrough
rlabel pdiffusion 787 -3218 787 -3218 0 feedthrough
rlabel pdiffusion 794 -3218 794 -3218 0 feedthrough
rlabel pdiffusion 801 -3218 801 -3218 0 feedthrough
rlabel pdiffusion 808 -3218 808 -3218 0 feedthrough
rlabel pdiffusion 815 -3218 815 -3218 0 feedthrough
rlabel pdiffusion 822 -3218 822 -3218 0 feedthrough
rlabel pdiffusion 829 -3218 829 -3218 0 feedthrough
rlabel pdiffusion 836 -3218 836 -3218 0 feedthrough
rlabel pdiffusion 843 -3218 843 -3218 0 feedthrough
rlabel pdiffusion 850 -3218 850 -3218 0 feedthrough
rlabel pdiffusion 857 -3218 857 -3218 0 feedthrough
rlabel pdiffusion 864 -3218 864 -3218 0 cellNo=128
rlabel pdiffusion 871 -3218 871 -3218 0 feedthrough
rlabel pdiffusion 878 -3218 878 -3218 0 feedthrough
rlabel pdiffusion 885 -3218 885 -3218 0 feedthrough
rlabel pdiffusion 892 -3218 892 -3218 0 feedthrough
rlabel pdiffusion 899 -3218 899 -3218 0 feedthrough
rlabel pdiffusion 906 -3218 906 -3218 0 feedthrough
rlabel pdiffusion 913 -3218 913 -3218 0 feedthrough
rlabel pdiffusion 920 -3218 920 -3218 0 feedthrough
rlabel pdiffusion 927 -3218 927 -3218 0 feedthrough
rlabel pdiffusion 934 -3218 934 -3218 0 feedthrough
rlabel pdiffusion 941 -3218 941 -3218 0 feedthrough
rlabel pdiffusion 948 -3218 948 -3218 0 feedthrough
rlabel pdiffusion 955 -3218 955 -3218 0 feedthrough
rlabel pdiffusion 962 -3218 962 -3218 0 feedthrough
rlabel pdiffusion 969 -3218 969 -3218 0 feedthrough
rlabel pdiffusion 976 -3218 976 -3218 0 feedthrough
rlabel pdiffusion 983 -3218 983 -3218 0 cellNo=780
rlabel pdiffusion 990 -3218 990 -3218 0 feedthrough
rlabel pdiffusion 997 -3218 997 -3218 0 feedthrough
rlabel pdiffusion 1004 -3218 1004 -3218 0 cellNo=838
rlabel pdiffusion 1011 -3218 1011 -3218 0 feedthrough
rlabel pdiffusion 1018 -3218 1018 -3218 0 feedthrough
rlabel pdiffusion 1025 -3218 1025 -3218 0 feedthrough
rlabel pdiffusion 1032 -3218 1032 -3218 0 feedthrough
rlabel pdiffusion 1039 -3218 1039 -3218 0 feedthrough
rlabel pdiffusion 1046 -3218 1046 -3218 0 feedthrough
rlabel pdiffusion 1053 -3218 1053 -3218 0 feedthrough
rlabel pdiffusion 1060 -3218 1060 -3218 0 cellNo=532
rlabel pdiffusion 1074 -3218 1074 -3218 0 feedthrough
rlabel pdiffusion 1081 -3218 1081 -3218 0 feedthrough
rlabel pdiffusion 1088 -3218 1088 -3218 0 feedthrough
rlabel pdiffusion 1095 -3218 1095 -3218 0 feedthrough
rlabel pdiffusion 1102 -3218 1102 -3218 0 feedthrough
rlabel pdiffusion 1109 -3218 1109 -3218 0 cellNo=742
rlabel pdiffusion 1116 -3218 1116 -3218 0 feedthrough
rlabel pdiffusion 1123 -3218 1123 -3218 0 feedthrough
rlabel pdiffusion 1130 -3218 1130 -3218 0 feedthrough
rlabel pdiffusion 1137 -3218 1137 -3218 0 feedthrough
rlabel pdiffusion 1144 -3218 1144 -3218 0 feedthrough
rlabel pdiffusion 1151 -3218 1151 -3218 0 feedthrough
rlabel pdiffusion 1158 -3218 1158 -3218 0 cellNo=255
rlabel pdiffusion 1165 -3218 1165 -3218 0 cellNo=688
rlabel pdiffusion 1172 -3218 1172 -3218 0 feedthrough
rlabel pdiffusion 1186 -3218 1186 -3218 0 feedthrough
rlabel pdiffusion 1193 -3218 1193 -3218 0 feedthrough
rlabel pdiffusion 1200 -3218 1200 -3218 0 feedthrough
rlabel pdiffusion 1207 -3218 1207 -3218 0 feedthrough
rlabel pdiffusion 1214 -3218 1214 -3218 0 feedthrough
rlabel pdiffusion 1235 -3218 1235 -3218 0 feedthrough
rlabel pdiffusion 1333 -3218 1333 -3218 0 feedthrough
rlabel pdiffusion 1361 -3218 1361 -3218 0 feedthrough
rlabel pdiffusion 1368 -3218 1368 -3218 0 feedthrough
rlabel pdiffusion 1410 -3218 1410 -3218 0 feedthrough
rlabel pdiffusion 1452 -3218 1452 -3218 0 feedthrough
rlabel pdiffusion 1459 -3218 1459 -3218 0 feedthrough
rlabel pdiffusion 1466 -3218 1466 -3218 0 feedthrough
rlabel pdiffusion 157 -3273 157 -3273 0 feedthrough
rlabel pdiffusion 164 -3273 164 -3273 0 feedthrough
rlabel pdiffusion 171 -3273 171 -3273 0 feedthrough
rlabel pdiffusion 178 -3273 178 -3273 0 feedthrough
rlabel pdiffusion 185 -3273 185 -3273 0 cellNo=573
rlabel pdiffusion 192 -3273 192 -3273 0 feedthrough
rlabel pdiffusion 199 -3273 199 -3273 0 feedthrough
rlabel pdiffusion 206 -3273 206 -3273 0 cellNo=995
rlabel pdiffusion 213 -3273 213 -3273 0 feedthrough
rlabel pdiffusion 220 -3273 220 -3273 0 feedthrough
rlabel pdiffusion 227 -3273 227 -3273 0 feedthrough
rlabel pdiffusion 234 -3273 234 -3273 0 feedthrough
rlabel pdiffusion 241 -3273 241 -3273 0 cellNo=884
rlabel pdiffusion 248 -3273 248 -3273 0 cellNo=301
rlabel pdiffusion 255 -3273 255 -3273 0 feedthrough
rlabel pdiffusion 262 -3273 262 -3273 0 cellNo=136
rlabel pdiffusion 269 -3273 269 -3273 0 feedthrough
rlabel pdiffusion 276 -3273 276 -3273 0 feedthrough
rlabel pdiffusion 283 -3273 283 -3273 0 feedthrough
rlabel pdiffusion 290 -3273 290 -3273 0 feedthrough
rlabel pdiffusion 297 -3273 297 -3273 0 feedthrough
rlabel pdiffusion 304 -3273 304 -3273 0 feedthrough
rlabel pdiffusion 311 -3273 311 -3273 0 feedthrough
rlabel pdiffusion 318 -3273 318 -3273 0 feedthrough
rlabel pdiffusion 325 -3273 325 -3273 0 feedthrough
rlabel pdiffusion 332 -3273 332 -3273 0 feedthrough
rlabel pdiffusion 339 -3273 339 -3273 0 feedthrough
rlabel pdiffusion 346 -3273 346 -3273 0 feedthrough
rlabel pdiffusion 353 -3273 353 -3273 0 feedthrough
rlabel pdiffusion 360 -3273 360 -3273 0 feedthrough
rlabel pdiffusion 367 -3273 367 -3273 0 feedthrough
rlabel pdiffusion 374 -3273 374 -3273 0 feedthrough
rlabel pdiffusion 381 -3273 381 -3273 0 feedthrough
rlabel pdiffusion 388 -3273 388 -3273 0 feedthrough
rlabel pdiffusion 395 -3273 395 -3273 0 cellNo=715
rlabel pdiffusion 402 -3273 402 -3273 0 cellNo=813
rlabel pdiffusion 409 -3273 409 -3273 0 feedthrough
rlabel pdiffusion 416 -3273 416 -3273 0 feedthrough
rlabel pdiffusion 423 -3273 423 -3273 0 feedthrough
rlabel pdiffusion 430 -3273 430 -3273 0 feedthrough
rlabel pdiffusion 437 -3273 437 -3273 0 feedthrough
rlabel pdiffusion 444 -3273 444 -3273 0 feedthrough
rlabel pdiffusion 451 -3273 451 -3273 0 feedthrough
rlabel pdiffusion 458 -3273 458 -3273 0 feedthrough
rlabel pdiffusion 465 -3273 465 -3273 0 feedthrough
rlabel pdiffusion 472 -3273 472 -3273 0 cellNo=633
rlabel pdiffusion 479 -3273 479 -3273 0 feedthrough
rlabel pdiffusion 486 -3273 486 -3273 0 cellNo=40
rlabel pdiffusion 493 -3273 493 -3273 0 feedthrough
rlabel pdiffusion 500 -3273 500 -3273 0 feedthrough
rlabel pdiffusion 507 -3273 507 -3273 0 feedthrough
rlabel pdiffusion 514 -3273 514 -3273 0 feedthrough
rlabel pdiffusion 521 -3273 521 -3273 0 feedthrough
rlabel pdiffusion 528 -3273 528 -3273 0 feedthrough
rlabel pdiffusion 535 -3273 535 -3273 0 feedthrough
rlabel pdiffusion 542 -3273 542 -3273 0 feedthrough
rlabel pdiffusion 549 -3273 549 -3273 0 feedthrough
rlabel pdiffusion 556 -3273 556 -3273 0 feedthrough
rlabel pdiffusion 563 -3273 563 -3273 0 feedthrough
rlabel pdiffusion 570 -3273 570 -3273 0 feedthrough
rlabel pdiffusion 577 -3273 577 -3273 0 feedthrough
rlabel pdiffusion 584 -3273 584 -3273 0 feedthrough
rlabel pdiffusion 591 -3273 591 -3273 0 cellNo=984
rlabel pdiffusion 598 -3273 598 -3273 0 feedthrough
rlabel pdiffusion 605 -3273 605 -3273 0 feedthrough
rlabel pdiffusion 612 -3273 612 -3273 0 feedthrough
rlabel pdiffusion 619 -3273 619 -3273 0 feedthrough
rlabel pdiffusion 626 -3273 626 -3273 0 feedthrough
rlabel pdiffusion 633 -3273 633 -3273 0 cellNo=974
rlabel pdiffusion 640 -3273 640 -3273 0 feedthrough
rlabel pdiffusion 647 -3273 647 -3273 0 feedthrough
rlabel pdiffusion 654 -3273 654 -3273 0 feedthrough
rlabel pdiffusion 661 -3273 661 -3273 0 feedthrough
rlabel pdiffusion 668 -3273 668 -3273 0 feedthrough
rlabel pdiffusion 675 -3273 675 -3273 0 feedthrough
rlabel pdiffusion 682 -3273 682 -3273 0 feedthrough
rlabel pdiffusion 689 -3273 689 -3273 0 feedthrough
rlabel pdiffusion 696 -3273 696 -3273 0 feedthrough
rlabel pdiffusion 703 -3273 703 -3273 0 feedthrough
rlabel pdiffusion 710 -3273 710 -3273 0 feedthrough
rlabel pdiffusion 717 -3273 717 -3273 0 feedthrough
rlabel pdiffusion 724 -3273 724 -3273 0 cellNo=461
rlabel pdiffusion 731 -3273 731 -3273 0 cellNo=295
rlabel pdiffusion 738 -3273 738 -3273 0 feedthrough
rlabel pdiffusion 745 -3273 745 -3273 0 feedthrough
rlabel pdiffusion 752 -3273 752 -3273 0 feedthrough
rlabel pdiffusion 759 -3273 759 -3273 0 feedthrough
rlabel pdiffusion 766 -3273 766 -3273 0 feedthrough
rlabel pdiffusion 773 -3273 773 -3273 0 feedthrough
rlabel pdiffusion 780 -3273 780 -3273 0 cellNo=720
rlabel pdiffusion 787 -3273 787 -3273 0 feedthrough
rlabel pdiffusion 794 -3273 794 -3273 0 feedthrough
rlabel pdiffusion 801 -3273 801 -3273 0 feedthrough
rlabel pdiffusion 808 -3273 808 -3273 0 feedthrough
rlabel pdiffusion 815 -3273 815 -3273 0 feedthrough
rlabel pdiffusion 822 -3273 822 -3273 0 feedthrough
rlabel pdiffusion 829 -3273 829 -3273 0 feedthrough
rlabel pdiffusion 843 -3273 843 -3273 0 feedthrough
rlabel pdiffusion 871 -3273 871 -3273 0 feedthrough
rlabel pdiffusion 878 -3273 878 -3273 0 cellNo=601
rlabel pdiffusion 885 -3273 885 -3273 0 feedthrough
rlabel pdiffusion 892 -3273 892 -3273 0 feedthrough
rlabel pdiffusion 899 -3273 899 -3273 0 feedthrough
rlabel pdiffusion 906 -3273 906 -3273 0 feedthrough
rlabel pdiffusion 913 -3273 913 -3273 0 feedthrough
rlabel pdiffusion 920 -3273 920 -3273 0 feedthrough
rlabel pdiffusion 927 -3273 927 -3273 0 feedthrough
rlabel pdiffusion 934 -3273 934 -3273 0 feedthrough
rlabel pdiffusion 941 -3273 941 -3273 0 feedthrough
rlabel pdiffusion 948 -3273 948 -3273 0 feedthrough
rlabel pdiffusion 955 -3273 955 -3273 0 feedthrough
rlabel pdiffusion 962 -3273 962 -3273 0 feedthrough
rlabel pdiffusion 983 -3273 983 -3273 0 feedthrough
rlabel pdiffusion 990 -3273 990 -3273 0 cellNo=238
rlabel pdiffusion 997 -3273 997 -3273 0 feedthrough
rlabel pdiffusion 1004 -3273 1004 -3273 0 feedthrough
rlabel pdiffusion 1067 -3273 1067 -3273 0 feedthrough
rlabel pdiffusion 1074 -3273 1074 -3273 0 feedthrough
rlabel pdiffusion 1081 -3273 1081 -3273 0 feedthrough
rlabel pdiffusion 1095 -3273 1095 -3273 0 feedthrough
rlabel pdiffusion 1102 -3273 1102 -3273 0 feedthrough
rlabel pdiffusion 1109 -3273 1109 -3273 0 feedthrough
rlabel pdiffusion 1123 -3273 1123 -3273 0 cellNo=78
rlabel pdiffusion 1130 -3273 1130 -3273 0 feedthrough
rlabel pdiffusion 1137 -3273 1137 -3273 0 feedthrough
rlabel pdiffusion 1144 -3273 1144 -3273 0 feedthrough
rlabel pdiffusion 1151 -3273 1151 -3273 0 feedthrough
rlabel pdiffusion 1158 -3273 1158 -3273 0 cellNo=670
rlabel pdiffusion 1165 -3273 1165 -3273 0 feedthrough
rlabel pdiffusion 1172 -3273 1172 -3273 0 feedthrough
rlabel pdiffusion 1186 -3273 1186 -3273 0 cellNo=910
rlabel pdiffusion 1207 -3273 1207 -3273 0 feedthrough
rlabel pdiffusion 1214 -3273 1214 -3273 0 cellNo=585
rlabel pdiffusion 1221 -3273 1221 -3273 0 feedthrough
rlabel pdiffusion 1235 -3273 1235 -3273 0 cellNo=233
rlabel pdiffusion 1249 -3273 1249 -3273 0 cellNo=625
rlabel pdiffusion 1291 -3273 1291 -3273 0 feedthrough
rlabel pdiffusion 1326 -3273 1326 -3273 0 cellNo=717
rlabel pdiffusion 1361 -3273 1361 -3273 0 feedthrough
rlabel pdiffusion 1368 -3273 1368 -3273 0 feedthrough
rlabel pdiffusion 1410 -3273 1410 -3273 0 feedthrough
rlabel pdiffusion 1452 -3273 1452 -3273 0 feedthrough
rlabel pdiffusion 1459 -3273 1459 -3273 0 cellNo=489
rlabel pdiffusion 1466 -3273 1466 -3273 0 feedthrough
rlabel pdiffusion 178 -3336 178 -3336 0 feedthrough
rlabel pdiffusion 185 -3336 185 -3336 0 feedthrough
rlabel pdiffusion 192 -3336 192 -3336 0 feedthrough
rlabel pdiffusion 199 -3336 199 -3336 0 feedthrough
rlabel pdiffusion 206 -3336 206 -3336 0 feedthrough
rlabel pdiffusion 213 -3336 213 -3336 0 feedthrough
rlabel pdiffusion 220 -3336 220 -3336 0 feedthrough
rlabel pdiffusion 227 -3336 227 -3336 0 cellNo=483
rlabel pdiffusion 234 -3336 234 -3336 0 feedthrough
rlabel pdiffusion 241 -3336 241 -3336 0 feedthrough
rlabel pdiffusion 248 -3336 248 -3336 0 feedthrough
rlabel pdiffusion 255 -3336 255 -3336 0 feedthrough
rlabel pdiffusion 262 -3336 262 -3336 0 cellNo=822
rlabel pdiffusion 269 -3336 269 -3336 0 feedthrough
rlabel pdiffusion 276 -3336 276 -3336 0 feedthrough
rlabel pdiffusion 283 -3336 283 -3336 0 feedthrough
rlabel pdiffusion 290 -3336 290 -3336 0 feedthrough
rlabel pdiffusion 297 -3336 297 -3336 0 feedthrough
rlabel pdiffusion 304 -3336 304 -3336 0 feedthrough
rlabel pdiffusion 311 -3336 311 -3336 0 feedthrough
rlabel pdiffusion 318 -3336 318 -3336 0 feedthrough
rlabel pdiffusion 325 -3336 325 -3336 0 feedthrough
rlabel pdiffusion 332 -3336 332 -3336 0 feedthrough
rlabel pdiffusion 339 -3336 339 -3336 0 feedthrough
rlabel pdiffusion 346 -3336 346 -3336 0 feedthrough
rlabel pdiffusion 353 -3336 353 -3336 0 feedthrough
rlabel pdiffusion 360 -3336 360 -3336 0 feedthrough
rlabel pdiffusion 367 -3336 367 -3336 0 feedthrough
rlabel pdiffusion 374 -3336 374 -3336 0 feedthrough
rlabel pdiffusion 381 -3336 381 -3336 0 cellNo=807
rlabel pdiffusion 388 -3336 388 -3336 0 feedthrough
rlabel pdiffusion 395 -3336 395 -3336 0 feedthrough
rlabel pdiffusion 402 -3336 402 -3336 0 feedthrough
rlabel pdiffusion 409 -3336 409 -3336 0 cellNo=853
rlabel pdiffusion 416 -3336 416 -3336 0 feedthrough
rlabel pdiffusion 423 -3336 423 -3336 0 feedthrough
rlabel pdiffusion 430 -3336 430 -3336 0 feedthrough
rlabel pdiffusion 437 -3336 437 -3336 0 feedthrough
rlabel pdiffusion 444 -3336 444 -3336 0 cellNo=911
rlabel pdiffusion 451 -3336 451 -3336 0 feedthrough
rlabel pdiffusion 458 -3336 458 -3336 0 feedthrough
rlabel pdiffusion 465 -3336 465 -3336 0 cellNo=894
rlabel pdiffusion 472 -3336 472 -3336 0 feedthrough
rlabel pdiffusion 479 -3336 479 -3336 0 feedthrough
rlabel pdiffusion 486 -3336 486 -3336 0 feedthrough
rlabel pdiffusion 493 -3336 493 -3336 0 feedthrough
rlabel pdiffusion 500 -3336 500 -3336 0 feedthrough
rlabel pdiffusion 507 -3336 507 -3336 0 feedthrough
rlabel pdiffusion 514 -3336 514 -3336 0 feedthrough
rlabel pdiffusion 521 -3336 521 -3336 0 feedthrough
rlabel pdiffusion 528 -3336 528 -3336 0 feedthrough
rlabel pdiffusion 535 -3336 535 -3336 0 feedthrough
rlabel pdiffusion 542 -3336 542 -3336 0 cellNo=514
rlabel pdiffusion 549 -3336 549 -3336 0 feedthrough
rlabel pdiffusion 556 -3336 556 -3336 0 feedthrough
rlabel pdiffusion 563 -3336 563 -3336 0 feedthrough
rlabel pdiffusion 570 -3336 570 -3336 0 cellNo=432
rlabel pdiffusion 577 -3336 577 -3336 0 feedthrough
rlabel pdiffusion 584 -3336 584 -3336 0 feedthrough
rlabel pdiffusion 591 -3336 591 -3336 0 cellNo=652
rlabel pdiffusion 598 -3336 598 -3336 0 feedthrough
rlabel pdiffusion 605 -3336 605 -3336 0 feedthrough
rlabel pdiffusion 612 -3336 612 -3336 0 feedthrough
rlabel pdiffusion 619 -3336 619 -3336 0 cellNo=926
rlabel pdiffusion 626 -3336 626 -3336 0 feedthrough
rlabel pdiffusion 633 -3336 633 -3336 0 feedthrough
rlabel pdiffusion 640 -3336 640 -3336 0 feedthrough
rlabel pdiffusion 647 -3336 647 -3336 0 feedthrough
rlabel pdiffusion 654 -3336 654 -3336 0 feedthrough
rlabel pdiffusion 661 -3336 661 -3336 0 feedthrough
rlabel pdiffusion 668 -3336 668 -3336 0 cellNo=743
rlabel pdiffusion 675 -3336 675 -3336 0 feedthrough
rlabel pdiffusion 682 -3336 682 -3336 0 cellNo=793
rlabel pdiffusion 689 -3336 689 -3336 0 feedthrough
rlabel pdiffusion 696 -3336 696 -3336 0 feedthrough
rlabel pdiffusion 703 -3336 703 -3336 0 feedthrough
rlabel pdiffusion 710 -3336 710 -3336 0 cellNo=872
rlabel pdiffusion 717 -3336 717 -3336 0 feedthrough
rlabel pdiffusion 724 -3336 724 -3336 0 feedthrough
rlabel pdiffusion 731 -3336 731 -3336 0 feedthrough
rlabel pdiffusion 738 -3336 738 -3336 0 cellNo=805
rlabel pdiffusion 745 -3336 745 -3336 0 feedthrough
rlabel pdiffusion 752 -3336 752 -3336 0 feedthrough
rlabel pdiffusion 759 -3336 759 -3336 0 feedthrough
rlabel pdiffusion 766 -3336 766 -3336 0 feedthrough
rlabel pdiffusion 773 -3336 773 -3336 0 feedthrough
rlabel pdiffusion 780 -3336 780 -3336 0 feedthrough
rlabel pdiffusion 787 -3336 787 -3336 0 feedthrough
rlabel pdiffusion 794 -3336 794 -3336 0 feedthrough
rlabel pdiffusion 801 -3336 801 -3336 0 feedthrough
rlabel pdiffusion 808 -3336 808 -3336 0 feedthrough
rlabel pdiffusion 815 -3336 815 -3336 0 feedthrough
rlabel pdiffusion 822 -3336 822 -3336 0 feedthrough
rlabel pdiffusion 829 -3336 829 -3336 0 feedthrough
rlabel pdiffusion 836 -3336 836 -3336 0 cellNo=415
rlabel pdiffusion 843 -3336 843 -3336 0 cellNo=758
rlabel pdiffusion 850 -3336 850 -3336 0 feedthrough
rlabel pdiffusion 857 -3336 857 -3336 0 feedthrough
rlabel pdiffusion 864 -3336 864 -3336 0 feedthrough
rlabel pdiffusion 871 -3336 871 -3336 0 feedthrough
rlabel pdiffusion 878 -3336 878 -3336 0 feedthrough
rlabel pdiffusion 885 -3336 885 -3336 0 feedthrough
rlabel pdiffusion 892 -3336 892 -3336 0 feedthrough
rlabel pdiffusion 899 -3336 899 -3336 0 feedthrough
rlabel pdiffusion 906 -3336 906 -3336 0 feedthrough
rlabel pdiffusion 913 -3336 913 -3336 0 feedthrough
rlabel pdiffusion 920 -3336 920 -3336 0 feedthrough
rlabel pdiffusion 927 -3336 927 -3336 0 feedthrough
rlabel pdiffusion 934 -3336 934 -3336 0 cellNo=213
rlabel pdiffusion 941 -3336 941 -3336 0 feedthrough
rlabel pdiffusion 948 -3336 948 -3336 0 cellNo=97
rlabel pdiffusion 955 -3336 955 -3336 0 feedthrough
rlabel pdiffusion 962 -3336 962 -3336 0 feedthrough
rlabel pdiffusion 976 -3336 976 -3336 0 feedthrough
rlabel pdiffusion 990 -3336 990 -3336 0 feedthrough
rlabel pdiffusion 1060 -3336 1060 -3336 0 cellNo=940
rlabel pdiffusion 1067 -3336 1067 -3336 0 feedthrough
rlabel pdiffusion 1074 -3336 1074 -3336 0 feedthrough
rlabel pdiffusion 1081 -3336 1081 -3336 0 feedthrough
rlabel pdiffusion 1095 -3336 1095 -3336 0 cellNo=523
rlabel pdiffusion 1109 -3336 1109 -3336 0 feedthrough
rlabel pdiffusion 1116 -3336 1116 -3336 0 feedthrough
rlabel pdiffusion 1137 -3336 1137 -3336 0 cellNo=562
rlabel pdiffusion 1144 -3336 1144 -3336 0 feedthrough
rlabel pdiffusion 1214 -3336 1214 -3336 0 feedthrough
rlabel pdiffusion 1291 -3336 1291 -3336 0 feedthrough
rlabel pdiffusion 1361 -3336 1361 -3336 0 feedthrough
rlabel pdiffusion 1368 -3336 1368 -3336 0 feedthrough
rlabel pdiffusion 1410 -3336 1410 -3336 0 feedthrough
rlabel pdiffusion 178 -3401 178 -3401 0 feedthrough
rlabel pdiffusion 185 -3401 185 -3401 0 feedthrough
rlabel pdiffusion 192 -3401 192 -3401 0 feedthrough
rlabel pdiffusion 199 -3401 199 -3401 0 feedthrough
rlabel pdiffusion 206 -3401 206 -3401 0 feedthrough
rlabel pdiffusion 213 -3401 213 -3401 0 feedthrough
rlabel pdiffusion 220 -3401 220 -3401 0 feedthrough
rlabel pdiffusion 227 -3401 227 -3401 0 cellNo=73
rlabel pdiffusion 234 -3401 234 -3401 0 feedthrough
rlabel pdiffusion 241 -3401 241 -3401 0 feedthrough
rlabel pdiffusion 248 -3401 248 -3401 0 feedthrough
rlabel pdiffusion 255 -3401 255 -3401 0 feedthrough
rlabel pdiffusion 262 -3401 262 -3401 0 feedthrough
rlabel pdiffusion 269 -3401 269 -3401 0 feedthrough
rlabel pdiffusion 276 -3401 276 -3401 0 feedthrough
rlabel pdiffusion 283 -3401 283 -3401 0 feedthrough
rlabel pdiffusion 290 -3401 290 -3401 0 feedthrough
rlabel pdiffusion 297 -3401 297 -3401 0 feedthrough
rlabel pdiffusion 304 -3401 304 -3401 0 feedthrough
rlabel pdiffusion 311 -3401 311 -3401 0 feedthrough
rlabel pdiffusion 318 -3401 318 -3401 0 feedthrough
rlabel pdiffusion 325 -3401 325 -3401 0 feedthrough
rlabel pdiffusion 332 -3401 332 -3401 0 feedthrough
rlabel pdiffusion 339 -3401 339 -3401 0 cellNo=915
rlabel pdiffusion 346 -3401 346 -3401 0 feedthrough
rlabel pdiffusion 353 -3401 353 -3401 0 cellNo=890
rlabel pdiffusion 360 -3401 360 -3401 0 feedthrough
rlabel pdiffusion 367 -3401 367 -3401 0 feedthrough
rlabel pdiffusion 374 -3401 374 -3401 0 feedthrough
rlabel pdiffusion 381 -3401 381 -3401 0 cellNo=708
rlabel pdiffusion 388 -3401 388 -3401 0 feedthrough
rlabel pdiffusion 395 -3401 395 -3401 0 cellNo=772
rlabel pdiffusion 402 -3401 402 -3401 0 feedthrough
rlabel pdiffusion 409 -3401 409 -3401 0 feedthrough
rlabel pdiffusion 416 -3401 416 -3401 0 feedthrough
rlabel pdiffusion 423 -3401 423 -3401 0 feedthrough
rlabel pdiffusion 430 -3401 430 -3401 0 feedthrough
rlabel pdiffusion 437 -3401 437 -3401 0 feedthrough
rlabel pdiffusion 444 -3401 444 -3401 0 feedthrough
rlabel pdiffusion 451 -3401 451 -3401 0 feedthrough
rlabel pdiffusion 458 -3401 458 -3401 0 feedthrough
rlabel pdiffusion 465 -3401 465 -3401 0 cellNo=498
rlabel pdiffusion 472 -3401 472 -3401 0 feedthrough
rlabel pdiffusion 479 -3401 479 -3401 0 feedthrough
rlabel pdiffusion 486 -3401 486 -3401 0 cellNo=725
rlabel pdiffusion 493 -3401 493 -3401 0 cellNo=35
rlabel pdiffusion 500 -3401 500 -3401 0 feedthrough
rlabel pdiffusion 507 -3401 507 -3401 0 cellNo=180
rlabel pdiffusion 514 -3401 514 -3401 0 feedthrough
rlabel pdiffusion 521 -3401 521 -3401 0 feedthrough
rlabel pdiffusion 528 -3401 528 -3401 0 feedthrough
rlabel pdiffusion 535 -3401 535 -3401 0 cellNo=683
rlabel pdiffusion 542 -3401 542 -3401 0 cellNo=388
rlabel pdiffusion 549 -3401 549 -3401 0 feedthrough
rlabel pdiffusion 556 -3401 556 -3401 0 cellNo=611
rlabel pdiffusion 563 -3401 563 -3401 0 feedthrough
rlabel pdiffusion 570 -3401 570 -3401 0 feedthrough
rlabel pdiffusion 577 -3401 577 -3401 0 cellNo=495
rlabel pdiffusion 584 -3401 584 -3401 0 feedthrough
rlabel pdiffusion 591 -3401 591 -3401 0 feedthrough
rlabel pdiffusion 598 -3401 598 -3401 0 feedthrough
rlabel pdiffusion 605 -3401 605 -3401 0 feedthrough
rlabel pdiffusion 612 -3401 612 -3401 0 feedthrough
rlabel pdiffusion 619 -3401 619 -3401 0 feedthrough
rlabel pdiffusion 626 -3401 626 -3401 0 feedthrough
rlabel pdiffusion 633 -3401 633 -3401 0 feedthrough
rlabel pdiffusion 640 -3401 640 -3401 0 feedthrough
rlabel pdiffusion 647 -3401 647 -3401 0 feedthrough
rlabel pdiffusion 654 -3401 654 -3401 0 feedthrough
rlabel pdiffusion 661 -3401 661 -3401 0 feedthrough
rlabel pdiffusion 668 -3401 668 -3401 0 feedthrough
rlabel pdiffusion 675 -3401 675 -3401 0 feedthrough
rlabel pdiffusion 682 -3401 682 -3401 0 feedthrough
rlabel pdiffusion 689 -3401 689 -3401 0 feedthrough
rlabel pdiffusion 696 -3401 696 -3401 0 feedthrough
rlabel pdiffusion 703 -3401 703 -3401 0 cellNo=842
rlabel pdiffusion 710 -3401 710 -3401 0 feedthrough
rlabel pdiffusion 717 -3401 717 -3401 0 feedthrough
rlabel pdiffusion 724 -3401 724 -3401 0 feedthrough
rlabel pdiffusion 731 -3401 731 -3401 0 feedthrough
rlabel pdiffusion 738 -3401 738 -3401 0 feedthrough
rlabel pdiffusion 745 -3401 745 -3401 0 feedthrough
rlabel pdiffusion 752 -3401 752 -3401 0 feedthrough
rlabel pdiffusion 759 -3401 759 -3401 0 feedthrough
rlabel pdiffusion 766 -3401 766 -3401 0 feedthrough
rlabel pdiffusion 773 -3401 773 -3401 0 cellNo=901
rlabel pdiffusion 780 -3401 780 -3401 0 feedthrough
rlabel pdiffusion 815 -3401 815 -3401 0 feedthrough
rlabel pdiffusion 822 -3401 822 -3401 0 feedthrough
rlabel pdiffusion 829 -3401 829 -3401 0 cellNo=311
rlabel pdiffusion 836 -3401 836 -3401 0 feedthrough
rlabel pdiffusion 843 -3401 843 -3401 0 cellNo=81
rlabel pdiffusion 850 -3401 850 -3401 0 feedthrough
rlabel pdiffusion 857 -3401 857 -3401 0 feedthrough
rlabel pdiffusion 864 -3401 864 -3401 0 cellNo=575
rlabel pdiffusion 871 -3401 871 -3401 0 feedthrough
rlabel pdiffusion 878 -3401 878 -3401 0 feedthrough
rlabel pdiffusion 885 -3401 885 -3401 0 feedthrough
rlabel pdiffusion 892 -3401 892 -3401 0 cellNo=775
rlabel pdiffusion 906 -3401 906 -3401 0 feedthrough
rlabel pdiffusion 913 -3401 913 -3401 0 feedthrough
rlabel pdiffusion 920 -3401 920 -3401 0 feedthrough
rlabel pdiffusion 927 -3401 927 -3401 0 feedthrough
rlabel pdiffusion 941 -3401 941 -3401 0 feedthrough
rlabel pdiffusion 990 -3401 990 -3401 0 feedthrough
rlabel pdiffusion 997 -3401 997 -3401 0 feedthrough
rlabel pdiffusion 1074 -3401 1074 -3401 0 feedthrough
rlabel pdiffusion 1116 -3401 1116 -3401 0 feedthrough
rlabel pdiffusion 1123 -3401 1123 -3401 0 feedthrough
rlabel pdiffusion 1214 -3401 1214 -3401 0 feedthrough
rlabel pdiffusion 1354 -3401 1354 -3401 0 feedthrough
rlabel pdiffusion 1361 -3401 1361 -3401 0 feedthrough
rlabel pdiffusion 1368 -3401 1368 -3401 0 feedthrough
rlabel pdiffusion 1410 -3401 1410 -3401 0 feedthrough
rlabel pdiffusion 220 -3444 220 -3444 0 cellNo=912
rlabel pdiffusion 241 -3444 241 -3444 0 feedthrough
rlabel pdiffusion 255 -3444 255 -3444 0 feedthrough
rlabel pdiffusion 262 -3444 262 -3444 0 cellNo=87
rlabel pdiffusion 269 -3444 269 -3444 0 feedthrough
rlabel pdiffusion 276 -3444 276 -3444 0 feedthrough
rlabel pdiffusion 283 -3444 283 -3444 0 feedthrough
rlabel pdiffusion 290 -3444 290 -3444 0 cellNo=387
rlabel pdiffusion 297 -3444 297 -3444 0 feedthrough
rlabel pdiffusion 304 -3444 304 -3444 0 cellNo=418
rlabel pdiffusion 311 -3444 311 -3444 0 feedthrough
rlabel pdiffusion 318 -3444 318 -3444 0 feedthrough
rlabel pdiffusion 325 -3444 325 -3444 0 cellNo=508
rlabel pdiffusion 339 -3444 339 -3444 0 cellNo=588
rlabel pdiffusion 346 -3444 346 -3444 0 feedthrough
rlabel pdiffusion 353 -3444 353 -3444 0 feedthrough
rlabel pdiffusion 360 -3444 360 -3444 0 feedthrough
rlabel pdiffusion 374 -3444 374 -3444 0 feedthrough
rlabel pdiffusion 388 -3444 388 -3444 0 feedthrough
rlabel pdiffusion 395 -3444 395 -3444 0 feedthrough
rlabel pdiffusion 402 -3444 402 -3444 0 feedthrough
rlabel pdiffusion 409 -3444 409 -3444 0 feedthrough
rlabel pdiffusion 423 -3444 423 -3444 0 feedthrough
rlabel pdiffusion 430 -3444 430 -3444 0 feedthrough
rlabel pdiffusion 437 -3444 437 -3444 0 feedthrough
rlabel pdiffusion 444 -3444 444 -3444 0 feedthrough
rlabel pdiffusion 451 -3444 451 -3444 0 feedthrough
rlabel pdiffusion 472 -3444 472 -3444 0 feedthrough
rlabel pdiffusion 486 -3444 486 -3444 0 feedthrough
rlabel pdiffusion 493 -3444 493 -3444 0 feedthrough
rlabel pdiffusion 500 -3444 500 -3444 0 cellNo=438
rlabel pdiffusion 535 -3444 535 -3444 0 feedthrough
rlabel pdiffusion 542 -3444 542 -3444 0 feedthrough
rlabel pdiffusion 549 -3444 549 -3444 0 feedthrough
rlabel pdiffusion 556 -3444 556 -3444 0 feedthrough
rlabel pdiffusion 563 -3444 563 -3444 0 feedthrough
rlabel pdiffusion 570 -3444 570 -3444 0 cellNo=727
rlabel pdiffusion 577 -3444 577 -3444 0 feedthrough
rlabel pdiffusion 584 -3444 584 -3444 0 feedthrough
rlabel pdiffusion 598 -3444 598 -3444 0 feedthrough
rlabel pdiffusion 626 -3444 626 -3444 0 feedthrough
rlabel pdiffusion 633 -3444 633 -3444 0 feedthrough
rlabel pdiffusion 640 -3444 640 -3444 0 cellNo=272
rlabel pdiffusion 647 -3444 647 -3444 0 feedthrough
rlabel pdiffusion 654 -3444 654 -3444 0 feedthrough
rlabel pdiffusion 661 -3444 661 -3444 0 feedthrough
rlabel pdiffusion 668 -3444 668 -3444 0 feedthrough
rlabel pdiffusion 675 -3444 675 -3444 0 feedthrough
rlabel pdiffusion 682 -3444 682 -3444 0 feedthrough
rlabel pdiffusion 689 -3444 689 -3444 0 feedthrough
rlabel pdiffusion 696 -3444 696 -3444 0 feedthrough
rlabel pdiffusion 703 -3444 703 -3444 0 feedthrough
rlabel pdiffusion 710 -3444 710 -3444 0 feedthrough
rlabel pdiffusion 717 -3444 717 -3444 0 cellNo=844
rlabel pdiffusion 724 -3444 724 -3444 0 cellNo=476
rlabel pdiffusion 731 -3444 731 -3444 0 feedthrough
rlabel pdiffusion 738 -3444 738 -3444 0 cellNo=441
rlabel pdiffusion 745 -3444 745 -3444 0 feedthrough
rlabel pdiffusion 752 -3444 752 -3444 0 feedthrough
rlabel pdiffusion 759 -3444 759 -3444 0 feedthrough
rlabel pdiffusion 766 -3444 766 -3444 0 feedthrough
rlabel pdiffusion 773 -3444 773 -3444 0 cellNo=751
rlabel pdiffusion 780 -3444 780 -3444 0 cellNo=504
rlabel pdiffusion 822 -3444 822 -3444 0 feedthrough
rlabel pdiffusion 829 -3444 829 -3444 0 cellNo=999
rlabel pdiffusion 836 -3444 836 -3444 0 feedthrough
rlabel pdiffusion 843 -3444 843 -3444 0 feedthrough
rlabel pdiffusion 850 -3444 850 -3444 0 feedthrough
rlabel pdiffusion 857 -3444 857 -3444 0 feedthrough
rlabel pdiffusion 864 -3444 864 -3444 0 feedthrough
rlabel pdiffusion 871 -3444 871 -3444 0 feedthrough
rlabel pdiffusion 885 -3444 885 -3444 0 feedthrough
rlabel pdiffusion 913 -3444 913 -3444 0 feedthrough
rlabel pdiffusion 920 -3444 920 -3444 0 feedthrough
rlabel pdiffusion 927 -3444 927 -3444 0 feedthrough
rlabel pdiffusion 941 -3444 941 -3444 0 feedthrough
rlabel pdiffusion 948 -3444 948 -3444 0 feedthrough
rlabel pdiffusion 955 -3444 955 -3444 0 cellNo=991
rlabel pdiffusion 962 -3444 962 -3444 0 cellNo=643
rlabel pdiffusion 969 -3444 969 -3444 0 feedthrough
rlabel pdiffusion 976 -3444 976 -3444 0 cellNo=93
rlabel pdiffusion 983 -3444 983 -3444 0 feedthrough
rlabel pdiffusion 990 -3444 990 -3444 0 feedthrough
rlabel pdiffusion 997 -3444 997 -3444 0 feedthrough
rlabel pdiffusion 1011 -3444 1011 -3444 0 feedthrough
rlabel pdiffusion 1074 -3444 1074 -3444 0 feedthrough
rlabel pdiffusion 1095 -3444 1095 -3444 0 feedthrough
rlabel pdiffusion 1116 -3444 1116 -3444 0 feedthrough
rlabel pdiffusion 1123 -3444 1123 -3444 0 feedthrough
rlabel pdiffusion 1214 -3444 1214 -3444 0 feedthrough
rlabel pdiffusion 1354 -3444 1354 -3444 0 feedthrough
rlabel pdiffusion 1361 -3444 1361 -3444 0 feedthrough
rlabel pdiffusion 1396 -3444 1396 -3444 0 feedthrough
rlabel pdiffusion 1410 -3444 1410 -3444 0 feedthrough
rlabel pdiffusion 255 -3471 255 -3471 0 feedthrough
rlabel pdiffusion 262 -3471 262 -3471 0 feedthrough
rlabel pdiffusion 304 -3471 304 -3471 0 feedthrough
rlabel pdiffusion 318 -3471 318 -3471 0 feedthrough
rlabel pdiffusion 325 -3471 325 -3471 0 cellNo=638
rlabel pdiffusion 332 -3471 332 -3471 0 feedthrough
rlabel pdiffusion 339 -3471 339 -3471 0 feedthrough
rlabel pdiffusion 353 -3471 353 -3471 0 feedthrough
rlabel pdiffusion 360 -3471 360 -3471 0 feedthrough
rlabel pdiffusion 381 -3471 381 -3471 0 feedthrough
rlabel pdiffusion 395 -3471 395 -3471 0 feedthrough
rlabel pdiffusion 402 -3471 402 -3471 0 feedthrough
rlabel pdiffusion 409 -3471 409 -3471 0 cellNo=563
rlabel pdiffusion 416 -3471 416 -3471 0 feedthrough
rlabel pdiffusion 423 -3471 423 -3471 0 cellNo=394
rlabel pdiffusion 430 -3471 430 -3471 0 feedthrough
rlabel pdiffusion 437 -3471 437 -3471 0 cellNo=959
rlabel pdiffusion 444 -3471 444 -3471 0 feedthrough
rlabel pdiffusion 458 -3471 458 -3471 0 cellNo=989
rlabel pdiffusion 465 -3471 465 -3471 0 cellNo=850
rlabel pdiffusion 472 -3471 472 -3471 0 cellNo=950
rlabel pdiffusion 479 -3471 479 -3471 0 feedthrough
rlabel pdiffusion 486 -3471 486 -3471 0 feedthrough
rlabel pdiffusion 493 -3471 493 -3471 0 feedthrough
rlabel pdiffusion 500 -3471 500 -3471 0 cellNo=630
rlabel pdiffusion 507 -3471 507 -3471 0 feedthrough
rlabel pdiffusion 514 -3471 514 -3471 0 cellNo=855
rlabel pdiffusion 521 -3471 521 -3471 0 feedthrough
rlabel pdiffusion 542 -3471 542 -3471 0 feedthrough
rlabel pdiffusion 549 -3471 549 -3471 0 feedthrough
rlabel pdiffusion 556 -3471 556 -3471 0 feedthrough
rlabel pdiffusion 563 -3471 563 -3471 0 feedthrough
rlabel pdiffusion 570 -3471 570 -3471 0 feedthrough
rlabel pdiffusion 577 -3471 577 -3471 0 feedthrough
rlabel pdiffusion 584 -3471 584 -3471 0 feedthrough
rlabel pdiffusion 605 -3471 605 -3471 0 feedthrough
rlabel pdiffusion 612 -3471 612 -3471 0 cellNo=578
rlabel pdiffusion 619 -3471 619 -3471 0 cellNo=985
rlabel pdiffusion 626 -3471 626 -3471 0 feedthrough
rlabel pdiffusion 647 -3471 647 -3471 0 feedthrough
rlabel pdiffusion 654 -3471 654 -3471 0 feedthrough
rlabel pdiffusion 661 -3471 661 -3471 0 feedthrough
rlabel pdiffusion 675 -3471 675 -3471 0 feedthrough
rlabel pdiffusion 682 -3471 682 -3471 0 feedthrough
rlabel pdiffusion 689 -3471 689 -3471 0 cellNo=679
rlabel pdiffusion 696 -3471 696 -3471 0 cellNo=313
rlabel pdiffusion 710 -3471 710 -3471 0 feedthrough
rlabel pdiffusion 738 -3471 738 -3471 0 feedthrough
rlabel pdiffusion 759 -3471 759 -3471 0 feedthrough
rlabel pdiffusion 822 -3471 822 -3471 0 cellNo=353
rlabel pdiffusion 836 -3471 836 -3471 0 feedthrough
rlabel pdiffusion 843 -3471 843 -3471 0 feedthrough
rlabel pdiffusion 850 -3471 850 -3471 0 cellNo=668
rlabel pdiffusion 857 -3471 857 -3471 0 feedthrough
rlabel pdiffusion 871 -3471 871 -3471 0 feedthrough
rlabel pdiffusion 885 -3471 885 -3471 0 feedthrough
rlabel pdiffusion 892 -3471 892 -3471 0 feedthrough
rlabel pdiffusion 913 -3471 913 -3471 0 feedthrough
rlabel pdiffusion 920 -3471 920 -3471 0 feedthrough
rlabel pdiffusion 927 -3471 927 -3471 0 feedthrough
rlabel pdiffusion 934 -3471 934 -3471 0 feedthrough
rlabel pdiffusion 941 -3471 941 -3471 0 feedthrough
rlabel pdiffusion 990 -3471 990 -3471 0 feedthrough
rlabel pdiffusion 997 -3471 997 -3471 0 feedthrough
rlabel pdiffusion 1067 -3471 1067 -3471 0 feedthrough
rlabel pdiffusion 1074 -3471 1074 -3471 0 cellNo=502
rlabel pdiffusion 1116 -3471 1116 -3471 0 feedthrough
rlabel pdiffusion 1123 -3471 1123 -3471 0 feedthrough
rlabel pdiffusion 1214 -3471 1214 -3471 0 feedthrough
rlabel pdiffusion 1221 -3471 1221 -3471 0 cellNo=515
rlabel pdiffusion 1228 -3471 1228 -3471 0 feedthrough
rlabel pdiffusion 1354 -3471 1354 -3471 0 feedthrough
rlabel pdiffusion 1361 -3471 1361 -3471 0 feedthrough
rlabel pdiffusion 1410 -3471 1410 -3471 0 feedthrough
rlabel pdiffusion 1417 -3471 1417 -3471 0 feedthrough
rlabel pdiffusion 262 -3494 262 -3494 0 feedthrough
rlabel pdiffusion 269 -3494 269 -3494 0 feedthrough
rlabel pdiffusion 311 -3494 311 -3494 0 feedthrough
rlabel pdiffusion 332 -3494 332 -3494 0 feedthrough
rlabel pdiffusion 339 -3494 339 -3494 0 feedthrough
rlabel pdiffusion 346 -3494 346 -3494 0 cellNo=608
rlabel pdiffusion 353 -3494 353 -3494 0 feedthrough
rlabel pdiffusion 409 -3494 409 -3494 0 feedthrough
rlabel pdiffusion 416 -3494 416 -3494 0 cellNo=616
rlabel pdiffusion 430 -3494 430 -3494 0 cellNo=746
rlabel pdiffusion 437 -3494 437 -3494 0 feedthrough
rlabel pdiffusion 479 -3494 479 -3494 0 feedthrough
rlabel pdiffusion 542 -3494 542 -3494 0 feedthrough
rlabel pdiffusion 549 -3494 549 -3494 0 feedthrough
rlabel pdiffusion 556 -3494 556 -3494 0 feedthrough
rlabel pdiffusion 570 -3494 570 -3494 0 feedthrough
rlabel pdiffusion 577 -3494 577 -3494 0 feedthrough
rlabel pdiffusion 584 -3494 584 -3494 0 feedthrough
rlabel pdiffusion 591 -3494 591 -3494 0 feedthrough
rlabel pdiffusion 598 -3494 598 -3494 0 cellNo=878
rlabel pdiffusion 647 -3494 647 -3494 0 cellNo=626
rlabel pdiffusion 654 -3494 654 -3494 0 feedthrough
rlabel pdiffusion 661 -3494 661 -3494 0 feedthrough
rlabel pdiffusion 682 -3494 682 -3494 0 feedthrough
rlabel pdiffusion 689 -3494 689 -3494 0 feedthrough
rlabel pdiffusion 717 -3494 717 -3494 0 feedthrough
rlabel pdiffusion 724 -3494 724 -3494 0 cellNo=614
rlabel pdiffusion 829 -3494 829 -3494 0 feedthrough
rlabel pdiffusion 836 -3494 836 -3494 0 feedthrough
rlabel pdiffusion 843 -3494 843 -3494 0 cellNo=425
rlabel pdiffusion 850 -3494 850 -3494 0 feedthrough
rlabel pdiffusion 878 -3494 878 -3494 0 feedthrough
rlabel pdiffusion 885 -3494 885 -3494 0 cellNo=123
rlabel pdiffusion 899 -3494 899 -3494 0 cellNo=695
rlabel pdiffusion 906 -3494 906 -3494 0 feedthrough
rlabel pdiffusion 913 -3494 913 -3494 0 feedthrough
rlabel pdiffusion 920 -3494 920 -3494 0 feedthrough
rlabel pdiffusion 927 -3494 927 -3494 0 feedthrough
rlabel pdiffusion 941 -3494 941 -3494 0 feedthrough
rlabel pdiffusion 948 -3494 948 -3494 0 cellNo=908
rlabel pdiffusion 990 -3494 990 -3494 0 cellNo=956
rlabel pdiffusion 997 -3494 997 -3494 0 feedthrough
rlabel pdiffusion 1095 -3494 1095 -3494 0 feedthrough
rlabel pdiffusion 1116 -3494 1116 -3494 0 cellNo=893
rlabel pdiffusion 1123 -3494 1123 -3494 0 feedthrough
rlabel pdiffusion 1221 -3494 1221 -3494 0 cellNo=332
rlabel pdiffusion 1354 -3494 1354 -3494 0 feedthrough
rlabel pdiffusion 1361 -3494 1361 -3494 0 feedthrough
rlabel pdiffusion 1410 -3494 1410 -3494 0 cellNo=660
rlabel pdiffusion 1417 -3494 1417 -3494 0 feedthrough
rlabel pdiffusion 269 -3509 269 -3509 0 cellNo=765
rlabel pdiffusion 276 -3509 276 -3509 0 feedthrough
rlabel pdiffusion 325 -3509 325 -3509 0 cellNo=52
rlabel pdiffusion 332 -3509 332 -3509 0 feedthrough
rlabel pdiffusion 353 -3509 353 -3509 0 cellNo=810
rlabel pdiffusion 360 -3509 360 -3509 0 feedthrough
rlabel pdiffusion 542 -3509 542 -3509 0 feedthrough
rlabel pdiffusion 549 -3509 549 -3509 0 cellNo=399
rlabel pdiffusion 556 -3509 556 -3509 0 cellNo=528
rlabel pdiffusion 563 -3509 563 -3509 0 cellNo=877
rlabel pdiffusion 570 -3509 570 -3509 0 feedthrough
rlabel pdiffusion 577 -3509 577 -3509 0 cellNo=294
rlabel pdiffusion 584 -3509 584 -3509 0 feedthrough
rlabel pdiffusion 661 -3509 661 -3509 0 cellNo=347
rlabel pdiffusion 668 -3509 668 -3509 0 feedthrough
rlabel pdiffusion 689 -3509 689 -3509 0 cellNo=693
rlabel pdiffusion 857 -3509 857 -3509 0 cellNo=953
rlabel pdiffusion 871 -3509 871 -3509 0 feedthrough
rlabel pdiffusion 878 -3509 878 -3509 0 feedthrough
rlabel pdiffusion 913 -3509 913 -3509 0 cellNo=545
rlabel pdiffusion 920 -3509 920 -3509 0 cellNo=700
rlabel pdiffusion 1354 -3509 1354 -3509 0 feedthrough
rlabel pdiffusion 1361 -3509 1361 -3509 0 cellNo=938
rlabel pdiffusion 1368 -3509 1368 -3509 0 feedthrough
rlabel polysilicon 282 -6 282 -6 0 1
rlabel polysilicon 285 -12 285 -12 0 4
rlabel polysilicon 317 -6 317 -6 0 1
rlabel polysilicon 317 -12 317 -12 0 3
rlabel polysilicon 345 -6 345 -6 0 1
rlabel polysilicon 345 -12 345 -12 0 3
rlabel polysilicon 352 -6 352 -6 0 1
rlabel polysilicon 352 -12 352 -12 0 3
rlabel polysilicon 425 -6 425 -6 0 2
rlabel polysilicon 425 -12 425 -12 0 4
rlabel polysilicon 436 -6 436 -6 0 1
rlabel polysilicon 436 -12 436 -12 0 3
rlabel polysilicon 443 -6 443 -6 0 1
rlabel polysilicon 443 -12 443 -12 0 3
rlabel polysilicon 450 -6 450 -6 0 1
rlabel polysilicon 450 -12 450 -12 0 3
rlabel polysilicon 457 -6 457 -6 0 1
rlabel polysilicon 460 -12 460 -12 0 4
rlabel polysilicon 464 -6 464 -6 0 1
rlabel polysilicon 464 -12 464 -12 0 3
rlabel polysilicon 478 -6 478 -6 0 1
rlabel polysilicon 478 -12 478 -12 0 3
rlabel polysilicon 506 -12 506 -12 0 3
rlabel polysilicon 509 -12 509 -12 0 4
rlabel polysilicon 513 -6 513 -6 0 1
rlabel polysilicon 513 -12 513 -12 0 3
rlabel polysilicon 905 -6 905 -6 0 1
rlabel polysilicon 905 -12 905 -12 0 3
rlabel polysilicon 947 -6 947 -6 0 1
rlabel polysilicon 950 -6 950 -6 0 2
rlabel polysilicon 989 -6 989 -6 0 1
rlabel polysilicon 989 -12 989 -12 0 3
rlabel polysilicon 226 -25 226 -25 0 1
rlabel polysilicon 226 -31 226 -31 0 3
rlabel polysilicon 289 -25 289 -25 0 1
rlabel polysilicon 289 -31 289 -31 0 3
rlabel polysilicon 303 -25 303 -25 0 1
rlabel polysilicon 303 -31 303 -31 0 3
rlabel polysilicon 338 -25 338 -25 0 1
rlabel polysilicon 338 -31 338 -31 0 3
rlabel polysilicon 345 -25 345 -25 0 1
rlabel polysilicon 348 -25 348 -25 0 2
rlabel polysilicon 352 -25 352 -25 0 1
rlabel polysilicon 352 -31 352 -31 0 3
rlabel polysilicon 359 -25 359 -25 0 1
rlabel polysilicon 362 -25 362 -25 0 2
rlabel polysilicon 366 -25 366 -25 0 1
rlabel polysilicon 366 -31 366 -31 0 3
rlabel polysilicon 373 -25 373 -25 0 1
rlabel polysilicon 373 -31 373 -31 0 3
rlabel polysilicon 380 -25 380 -25 0 1
rlabel polysilicon 380 -31 380 -31 0 3
rlabel polysilicon 387 -25 387 -25 0 1
rlabel polysilicon 387 -31 387 -31 0 3
rlabel polysilicon 394 -25 394 -25 0 1
rlabel polysilicon 394 -31 394 -31 0 3
rlabel polysilicon 408 -25 408 -25 0 1
rlabel polysilicon 408 -31 408 -31 0 3
rlabel polysilicon 418 -25 418 -25 0 2
rlabel polysilicon 418 -31 418 -31 0 4
rlabel polysilicon 422 -25 422 -25 0 1
rlabel polysilicon 422 -31 422 -31 0 3
rlabel polysilicon 436 -25 436 -25 0 1
rlabel polysilicon 436 -31 436 -31 0 3
rlabel polysilicon 450 -25 450 -25 0 1
rlabel polysilicon 450 -31 450 -31 0 3
rlabel polysilicon 457 -25 457 -25 0 1
rlabel polysilicon 457 -31 457 -31 0 3
rlabel polysilicon 464 -25 464 -25 0 1
rlabel polysilicon 464 -31 464 -31 0 3
rlabel polysilicon 499 -25 499 -25 0 1
rlabel polysilicon 499 -31 499 -31 0 3
rlabel polysilicon 509 -25 509 -25 0 2
rlabel polysilicon 506 -31 506 -31 0 3
rlabel polysilicon 513 -25 513 -25 0 1
rlabel polysilicon 513 -31 513 -31 0 3
rlabel polysilicon 520 -31 520 -31 0 3
rlabel polysilicon 523 -31 523 -31 0 4
rlabel polysilicon 527 -25 527 -25 0 1
rlabel polysilicon 527 -31 527 -31 0 3
rlabel polysilicon 537 -25 537 -25 0 2
rlabel polysilicon 537 -31 537 -31 0 4
rlabel polysilicon 541 -25 541 -25 0 1
rlabel polysilicon 541 -31 541 -31 0 3
rlabel polysilicon 548 -25 548 -25 0 1
rlabel polysilicon 548 -31 548 -31 0 3
rlabel polysilicon 579 -25 579 -25 0 2
rlabel polysilicon 583 -25 583 -25 0 1
rlabel polysilicon 590 -25 590 -25 0 1
rlabel polysilicon 590 -31 590 -31 0 3
rlabel polysilicon 597 -25 597 -25 0 1
rlabel polysilicon 597 -31 597 -31 0 3
rlabel polysilicon 604 -25 604 -25 0 1
rlabel polysilicon 604 -31 604 -31 0 3
rlabel polysilicon 611 -25 611 -25 0 1
rlabel polysilicon 611 -31 611 -31 0 3
rlabel polysilicon 618 -25 618 -25 0 1
rlabel polysilicon 625 -25 625 -25 0 1
rlabel polysilicon 625 -31 625 -31 0 3
rlabel polysilicon 635 -31 635 -31 0 4
rlabel polysilicon 639 -25 639 -25 0 1
rlabel polysilicon 639 -31 639 -31 0 3
rlabel polysilicon 674 -25 674 -25 0 1
rlabel polysilicon 674 -31 674 -31 0 3
rlabel polysilicon 891 -25 891 -25 0 1
rlabel polysilicon 891 -31 891 -31 0 3
rlabel polysilicon 1003 -25 1003 -25 0 1
rlabel polysilicon 1003 -31 1003 -31 0 3
rlabel polysilicon 219 -48 219 -48 0 1
rlabel polysilicon 219 -54 219 -54 0 3
rlabel polysilicon 275 -48 275 -48 0 1
rlabel polysilicon 275 -54 275 -54 0 3
rlabel polysilicon 282 -48 282 -48 0 1
rlabel polysilicon 282 -54 282 -54 0 3
rlabel polysilicon 296 -48 296 -48 0 1
rlabel polysilicon 299 -54 299 -54 0 4
rlabel polysilicon 303 -48 303 -48 0 1
rlabel polysilicon 303 -54 303 -54 0 3
rlabel polysilicon 320 -54 320 -54 0 4
rlabel polysilicon 324 -48 324 -48 0 1
rlabel polysilicon 324 -54 324 -54 0 3
rlabel polysilicon 331 -48 331 -48 0 1
rlabel polysilicon 331 -54 331 -54 0 3
rlabel polysilicon 338 -48 338 -48 0 1
rlabel polysilicon 341 -48 341 -48 0 2
rlabel polysilicon 338 -54 338 -54 0 3
rlabel polysilicon 341 -54 341 -54 0 4
rlabel polysilicon 345 -48 345 -48 0 1
rlabel polysilicon 345 -54 345 -54 0 3
rlabel polysilicon 352 -48 352 -48 0 1
rlabel polysilicon 352 -54 352 -54 0 3
rlabel polysilicon 359 -48 359 -48 0 1
rlabel polysilicon 359 -54 359 -54 0 3
rlabel polysilicon 366 -48 366 -48 0 1
rlabel polysilicon 366 -54 366 -54 0 3
rlabel polysilicon 373 -48 373 -48 0 1
rlabel polysilicon 373 -54 373 -54 0 3
rlabel polysilicon 380 -48 380 -48 0 1
rlabel polysilicon 380 -54 380 -54 0 3
rlabel polysilicon 387 -48 387 -48 0 1
rlabel polysilicon 390 -54 390 -54 0 4
rlabel polysilicon 394 -48 394 -48 0 1
rlabel polysilicon 394 -54 394 -54 0 3
rlabel polysilicon 401 -48 401 -48 0 1
rlabel polysilicon 401 -54 401 -54 0 3
rlabel polysilicon 408 -48 408 -48 0 1
rlabel polysilicon 408 -54 408 -54 0 3
rlabel polysilicon 415 -48 415 -48 0 1
rlabel polysilicon 415 -54 415 -54 0 3
rlabel polysilicon 422 -48 422 -48 0 1
rlabel polysilicon 422 -54 422 -54 0 3
rlabel polysilicon 429 -48 429 -48 0 1
rlabel polysilicon 432 -48 432 -48 0 2
rlabel polysilicon 429 -54 429 -54 0 3
rlabel polysilicon 436 -48 436 -48 0 1
rlabel polysilicon 436 -54 436 -54 0 3
rlabel polysilicon 443 -48 443 -48 0 1
rlabel polysilicon 443 -54 443 -54 0 3
rlabel polysilicon 450 -48 450 -48 0 1
rlabel polysilicon 450 -54 450 -54 0 3
rlabel polysilicon 457 -48 457 -48 0 1
rlabel polysilicon 457 -54 457 -54 0 3
rlabel polysilicon 464 -48 464 -48 0 1
rlabel polysilicon 464 -54 464 -54 0 3
rlabel polysilicon 471 -48 471 -48 0 1
rlabel polysilicon 471 -54 471 -54 0 3
rlabel polysilicon 485 -48 485 -48 0 1
rlabel polysilicon 485 -54 485 -54 0 3
rlabel polysilicon 492 -48 492 -48 0 1
rlabel polysilicon 492 -54 492 -54 0 3
rlabel polysilicon 499 -48 499 -48 0 1
rlabel polysilicon 499 -54 499 -54 0 3
rlabel polysilicon 506 -48 506 -48 0 1
rlabel polysilicon 506 -54 506 -54 0 3
rlabel polysilicon 520 -48 520 -48 0 1
rlabel polysilicon 520 -54 520 -54 0 3
rlabel polysilicon 541 -48 541 -48 0 1
rlabel polysilicon 541 -54 541 -54 0 3
rlabel polysilicon 551 -48 551 -48 0 2
rlabel polysilicon 548 -54 548 -54 0 3
rlabel polysilicon 555 -48 555 -48 0 1
rlabel polysilicon 555 -54 555 -54 0 3
rlabel polysilicon 565 -48 565 -48 0 2
rlabel polysilicon 562 -54 562 -54 0 3
rlabel polysilicon 569 -54 569 -54 0 3
rlabel polysilicon 572 -54 572 -54 0 4
rlabel polysilicon 576 -48 576 -48 0 1
rlabel polysilicon 576 -54 576 -54 0 3
rlabel polysilicon 583 -48 583 -48 0 1
rlabel polysilicon 583 -54 583 -54 0 3
rlabel polysilicon 590 -48 590 -48 0 1
rlabel polysilicon 590 -54 590 -54 0 3
rlabel polysilicon 597 -48 597 -48 0 1
rlabel polysilicon 597 -54 597 -54 0 3
rlabel polysilicon 604 -48 604 -48 0 1
rlabel polysilicon 604 -54 604 -54 0 3
rlabel polysilicon 611 -54 611 -54 0 3
rlabel polysilicon 614 -54 614 -54 0 4
rlabel polysilicon 621 -48 621 -48 0 2
rlabel polysilicon 621 -54 621 -54 0 4
rlabel polysilicon 625 -48 625 -48 0 1
rlabel polysilicon 625 -54 625 -54 0 3
rlabel polysilicon 632 -48 632 -48 0 1
rlabel polysilicon 632 -54 632 -54 0 3
rlabel polysilicon 639 -48 639 -48 0 1
rlabel polysilicon 639 -54 639 -54 0 3
rlabel polysilicon 653 -48 653 -48 0 1
rlabel polysilicon 653 -54 653 -54 0 3
rlabel polysilicon 674 -48 674 -48 0 1
rlabel polysilicon 674 -54 674 -54 0 3
rlabel polysilicon 681 -48 681 -48 0 1
rlabel polysilicon 681 -54 681 -54 0 3
rlabel polysilicon 723 -48 723 -48 0 1
rlabel polysilicon 723 -54 723 -54 0 3
rlabel polysilicon 730 -48 730 -48 0 1
rlabel polysilicon 730 -54 730 -54 0 3
rlabel polysilicon 758 -48 758 -48 0 1
rlabel polysilicon 758 -54 758 -54 0 3
rlabel polysilicon 828 -48 828 -48 0 1
rlabel polysilicon 828 -54 828 -54 0 3
rlabel polysilicon 884 -48 884 -48 0 1
rlabel polysilicon 884 -54 884 -54 0 3
rlabel polysilicon 1010 -48 1010 -48 0 1
rlabel polysilicon 1010 -54 1010 -54 0 3
rlabel polysilicon 191 -99 191 -99 0 1
rlabel polysilicon 191 -105 191 -105 0 3
rlabel polysilicon 205 -99 205 -99 0 1
rlabel polysilicon 205 -105 205 -105 0 3
rlabel polysilicon 219 -99 219 -99 0 1
rlabel polysilicon 219 -105 219 -105 0 3
rlabel polysilicon 233 -99 233 -99 0 1
rlabel polysilicon 233 -105 233 -105 0 3
rlabel polysilicon 240 -99 240 -99 0 1
rlabel polysilicon 243 -99 243 -99 0 2
rlabel polysilicon 247 -99 247 -99 0 1
rlabel polysilicon 247 -105 247 -105 0 3
rlabel polysilicon 254 -99 254 -99 0 1
rlabel polysilicon 254 -105 254 -105 0 3
rlabel polysilicon 257 -105 257 -105 0 4
rlabel polysilicon 261 -99 261 -99 0 1
rlabel polysilicon 261 -105 261 -105 0 3
rlabel polysilicon 271 -105 271 -105 0 4
rlabel polysilicon 275 -99 275 -99 0 1
rlabel polysilicon 278 -99 278 -99 0 2
rlabel polysilicon 275 -105 275 -105 0 3
rlabel polysilicon 282 -99 282 -99 0 1
rlabel polysilicon 282 -105 282 -105 0 3
rlabel polysilicon 289 -99 289 -99 0 1
rlabel polysilicon 289 -105 289 -105 0 3
rlabel polysilicon 296 -99 296 -99 0 1
rlabel polysilicon 299 -99 299 -99 0 2
rlabel polysilicon 299 -105 299 -105 0 4
rlabel polysilicon 303 -99 303 -99 0 1
rlabel polysilicon 303 -105 303 -105 0 3
rlabel polysilicon 310 -99 310 -99 0 1
rlabel polysilicon 310 -105 310 -105 0 3
rlabel polysilicon 317 -99 317 -99 0 1
rlabel polysilicon 317 -105 317 -105 0 3
rlabel polysilicon 324 -99 324 -99 0 1
rlabel polysilicon 324 -105 324 -105 0 3
rlabel polysilicon 331 -99 331 -99 0 1
rlabel polysilicon 331 -105 331 -105 0 3
rlabel polysilicon 338 -99 338 -99 0 1
rlabel polysilicon 338 -105 338 -105 0 3
rlabel polysilicon 345 -99 345 -99 0 1
rlabel polysilicon 345 -105 345 -105 0 3
rlabel polysilicon 352 -99 352 -99 0 1
rlabel polysilicon 352 -105 352 -105 0 3
rlabel polysilicon 359 -99 359 -99 0 1
rlabel polysilicon 359 -105 359 -105 0 3
rlabel polysilicon 366 -99 366 -99 0 1
rlabel polysilicon 366 -105 366 -105 0 3
rlabel polysilicon 373 -99 373 -99 0 1
rlabel polysilicon 373 -105 373 -105 0 3
rlabel polysilicon 380 -99 380 -99 0 1
rlabel polysilicon 383 -99 383 -99 0 2
rlabel polysilicon 383 -105 383 -105 0 4
rlabel polysilicon 390 -99 390 -99 0 2
rlabel polysilicon 387 -105 387 -105 0 3
rlabel polysilicon 390 -105 390 -105 0 4
rlabel polysilicon 394 -99 394 -99 0 1
rlabel polysilicon 394 -105 394 -105 0 3
rlabel polysilicon 401 -99 401 -99 0 1
rlabel polysilicon 401 -105 401 -105 0 3
rlabel polysilicon 408 -99 408 -99 0 1
rlabel polysilicon 408 -105 408 -105 0 3
rlabel polysilicon 415 -99 415 -99 0 1
rlabel polysilicon 415 -105 415 -105 0 3
rlabel polysilicon 422 -99 422 -99 0 1
rlabel polysilicon 422 -105 422 -105 0 3
rlabel polysilicon 429 -99 429 -99 0 1
rlabel polysilicon 429 -105 429 -105 0 3
rlabel polysilicon 436 -99 436 -99 0 1
rlabel polysilicon 436 -105 436 -105 0 3
rlabel polysilicon 443 -99 443 -99 0 1
rlabel polysilicon 443 -105 443 -105 0 3
rlabel polysilicon 450 -99 450 -99 0 1
rlabel polysilicon 450 -105 450 -105 0 3
rlabel polysilicon 457 -99 457 -99 0 1
rlabel polysilicon 457 -105 457 -105 0 3
rlabel polysilicon 464 -99 464 -99 0 1
rlabel polysilicon 464 -105 464 -105 0 3
rlabel polysilicon 471 -99 471 -99 0 1
rlabel polysilicon 471 -105 471 -105 0 3
rlabel polysilicon 478 -99 478 -99 0 1
rlabel polysilicon 478 -105 478 -105 0 3
rlabel polysilicon 485 -99 485 -99 0 1
rlabel polysilicon 485 -105 485 -105 0 3
rlabel polysilicon 492 -99 492 -99 0 1
rlabel polysilicon 492 -105 492 -105 0 3
rlabel polysilicon 499 -99 499 -99 0 1
rlabel polysilicon 499 -105 499 -105 0 3
rlabel polysilicon 509 -99 509 -99 0 2
rlabel polysilicon 506 -105 506 -105 0 3
rlabel polysilicon 509 -105 509 -105 0 4
rlabel polysilicon 513 -99 513 -99 0 1
rlabel polysilicon 516 -99 516 -99 0 2
rlabel polysilicon 513 -105 513 -105 0 3
rlabel polysilicon 516 -105 516 -105 0 4
rlabel polysilicon 520 -99 520 -99 0 1
rlabel polysilicon 523 -99 523 -99 0 2
rlabel polysilicon 520 -105 520 -105 0 3
rlabel polysilicon 527 -99 527 -99 0 1
rlabel polysilicon 527 -105 527 -105 0 3
rlabel polysilicon 534 -99 534 -99 0 1
rlabel polysilicon 537 -105 537 -105 0 4
rlabel polysilicon 541 -105 541 -105 0 3
rlabel polysilicon 548 -99 548 -99 0 1
rlabel polysilicon 548 -105 548 -105 0 3
rlabel polysilicon 555 -99 555 -99 0 1
rlabel polysilicon 555 -105 555 -105 0 3
rlabel polysilicon 562 -105 562 -105 0 3
rlabel polysilicon 565 -105 565 -105 0 4
rlabel polysilicon 569 -99 569 -99 0 1
rlabel polysilicon 569 -105 569 -105 0 3
rlabel polysilicon 576 -99 576 -99 0 1
rlabel polysilicon 576 -105 576 -105 0 3
rlabel polysilicon 586 -99 586 -99 0 2
rlabel polysilicon 583 -105 583 -105 0 3
rlabel polysilicon 586 -105 586 -105 0 4
rlabel polysilicon 590 -99 590 -99 0 1
rlabel polysilicon 590 -105 590 -105 0 3
rlabel polysilicon 597 -99 597 -99 0 1
rlabel polysilicon 597 -105 597 -105 0 3
rlabel polysilicon 604 -99 604 -99 0 1
rlabel polysilicon 604 -105 604 -105 0 3
rlabel polysilicon 611 -99 611 -99 0 1
rlabel polysilicon 611 -105 611 -105 0 3
rlabel polysilicon 618 -99 618 -99 0 1
rlabel polysilicon 618 -105 618 -105 0 3
rlabel polysilicon 628 -99 628 -99 0 2
rlabel polysilicon 625 -105 625 -105 0 3
rlabel polysilicon 628 -105 628 -105 0 4
rlabel polysilicon 632 -99 632 -99 0 1
rlabel polysilicon 632 -105 632 -105 0 3
rlabel polysilicon 639 -99 639 -99 0 1
rlabel polysilicon 639 -105 639 -105 0 3
rlabel polysilicon 646 -99 646 -99 0 1
rlabel polysilicon 646 -105 646 -105 0 3
rlabel polysilicon 653 -99 653 -99 0 1
rlabel polysilicon 653 -105 653 -105 0 3
rlabel polysilicon 660 -99 660 -99 0 1
rlabel polysilicon 660 -105 660 -105 0 3
rlabel polysilicon 667 -99 667 -99 0 1
rlabel polysilicon 667 -105 667 -105 0 3
rlabel polysilicon 681 -99 681 -99 0 1
rlabel polysilicon 681 -105 681 -105 0 3
rlabel polysilicon 688 -99 688 -99 0 1
rlabel polysilicon 688 -105 688 -105 0 3
rlabel polysilicon 702 -99 702 -99 0 1
rlabel polysilicon 702 -105 702 -105 0 3
rlabel polysilicon 709 -99 709 -99 0 1
rlabel polysilicon 709 -105 709 -105 0 3
rlabel polysilicon 723 -99 723 -99 0 1
rlabel polysilicon 723 -105 723 -105 0 3
rlabel polysilicon 730 -99 730 -99 0 1
rlabel polysilicon 730 -105 730 -105 0 3
rlabel polysilicon 737 -99 737 -99 0 1
rlabel polysilicon 737 -105 737 -105 0 3
rlabel polysilicon 779 -99 779 -99 0 1
rlabel polysilicon 782 -99 782 -99 0 2
rlabel polysilicon 782 -105 782 -105 0 4
rlabel polysilicon 789 -99 789 -99 0 2
rlabel polysilicon 786 -105 786 -105 0 3
rlabel polysilicon 793 -99 793 -99 0 1
rlabel polysilicon 793 -105 793 -105 0 3
rlabel polysilicon 800 -99 800 -99 0 1
rlabel polysilicon 800 -105 800 -105 0 3
rlabel polysilicon 807 -99 807 -99 0 1
rlabel polysilicon 807 -105 807 -105 0 3
rlabel polysilicon 863 -99 863 -99 0 1
rlabel polysilicon 863 -105 863 -105 0 3
rlabel polysilicon 891 -99 891 -99 0 1
rlabel polysilicon 891 -105 891 -105 0 3
rlabel polysilicon 898 -99 898 -99 0 1
rlabel polysilicon 898 -105 898 -105 0 3
rlabel polysilicon 1017 -99 1017 -99 0 1
rlabel polysilicon 1017 -105 1017 -105 0 3
rlabel polysilicon 114 -166 114 -166 0 1
rlabel polysilicon 114 -172 114 -172 0 3
rlabel polysilicon 121 -166 121 -166 0 1
rlabel polysilicon 121 -172 121 -172 0 3
rlabel polysilicon 128 -166 128 -166 0 1
rlabel polysilicon 128 -172 128 -172 0 3
rlabel polysilicon 135 -166 135 -166 0 1
rlabel polysilicon 135 -172 135 -172 0 3
rlabel polysilicon 142 -166 142 -166 0 1
rlabel polysilicon 142 -172 142 -172 0 3
rlabel polysilicon 149 -166 149 -166 0 1
rlabel polysilicon 149 -172 149 -172 0 3
rlabel polysilicon 156 -166 156 -166 0 1
rlabel polysilicon 156 -172 156 -172 0 3
rlabel polysilicon 163 -166 163 -166 0 1
rlabel polysilicon 163 -172 163 -172 0 3
rlabel polysilicon 170 -166 170 -166 0 1
rlabel polysilicon 170 -172 170 -172 0 3
rlabel polysilicon 177 -166 177 -166 0 1
rlabel polysilicon 177 -172 177 -172 0 3
rlabel polysilicon 184 -166 184 -166 0 1
rlabel polysilicon 184 -172 184 -172 0 3
rlabel polysilicon 191 -166 191 -166 0 1
rlabel polysilicon 191 -172 191 -172 0 3
rlabel polysilicon 198 -166 198 -166 0 1
rlabel polysilicon 198 -172 198 -172 0 3
rlabel polysilicon 205 -166 205 -166 0 1
rlabel polysilicon 205 -172 205 -172 0 3
rlabel polysilicon 212 -166 212 -166 0 1
rlabel polysilicon 212 -172 212 -172 0 3
rlabel polysilicon 219 -166 219 -166 0 1
rlabel polysilicon 219 -172 219 -172 0 3
rlabel polysilicon 226 -166 226 -166 0 1
rlabel polysilicon 229 -166 229 -166 0 2
rlabel polysilicon 226 -172 226 -172 0 3
rlabel polysilicon 233 -166 233 -166 0 1
rlabel polysilicon 233 -172 233 -172 0 3
rlabel polysilicon 240 -166 240 -166 0 1
rlabel polysilicon 240 -172 240 -172 0 3
rlabel polysilicon 247 -166 247 -166 0 1
rlabel polysilicon 247 -172 247 -172 0 3
rlabel polysilicon 254 -166 254 -166 0 1
rlabel polysilicon 254 -172 254 -172 0 3
rlabel polysilicon 261 -166 261 -166 0 1
rlabel polysilicon 261 -172 261 -172 0 3
rlabel polysilicon 268 -166 268 -166 0 1
rlabel polysilicon 268 -172 268 -172 0 3
rlabel polysilicon 275 -166 275 -166 0 1
rlabel polysilicon 275 -172 275 -172 0 3
rlabel polysilicon 282 -166 282 -166 0 1
rlabel polysilicon 282 -172 282 -172 0 3
rlabel polysilicon 289 -166 289 -166 0 1
rlabel polysilicon 289 -172 289 -172 0 3
rlabel polysilicon 296 -166 296 -166 0 1
rlabel polysilicon 299 -166 299 -166 0 2
rlabel polysilicon 296 -172 296 -172 0 3
rlabel polysilicon 303 -166 303 -166 0 1
rlabel polysilicon 303 -172 303 -172 0 3
rlabel polysilicon 310 -166 310 -166 0 1
rlabel polysilicon 310 -172 310 -172 0 3
rlabel polysilicon 317 -166 317 -166 0 1
rlabel polysilicon 317 -172 317 -172 0 3
rlabel polysilicon 324 -166 324 -166 0 1
rlabel polysilicon 324 -172 324 -172 0 3
rlabel polysilicon 331 -166 331 -166 0 1
rlabel polysilicon 334 -166 334 -166 0 2
rlabel polysilicon 331 -172 331 -172 0 3
rlabel polysilicon 334 -172 334 -172 0 4
rlabel polysilicon 338 -166 338 -166 0 1
rlabel polysilicon 338 -172 338 -172 0 3
rlabel polysilicon 345 -166 345 -166 0 1
rlabel polysilicon 345 -172 345 -172 0 3
rlabel polysilicon 352 -166 352 -166 0 1
rlabel polysilicon 352 -172 352 -172 0 3
rlabel polysilicon 359 -166 359 -166 0 1
rlabel polysilicon 359 -172 359 -172 0 3
rlabel polysilicon 366 -166 366 -166 0 1
rlabel polysilicon 369 -166 369 -166 0 2
rlabel polysilicon 369 -172 369 -172 0 4
rlabel polysilicon 373 -166 373 -166 0 1
rlabel polysilicon 373 -172 373 -172 0 3
rlabel polysilicon 380 -166 380 -166 0 1
rlabel polysilicon 380 -172 380 -172 0 3
rlabel polysilicon 390 -166 390 -166 0 2
rlabel polysilicon 387 -172 387 -172 0 3
rlabel polysilicon 390 -172 390 -172 0 4
rlabel polysilicon 394 -166 394 -166 0 1
rlabel polysilicon 394 -172 394 -172 0 3
rlabel polysilicon 401 -166 401 -166 0 1
rlabel polysilicon 401 -172 401 -172 0 3
rlabel polysilicon 404 -172 404 -172 0 4
rlabel polysilicon 408 -166 408 -166 0 1
rlabel polysilicon 408 -172 408 -172 0 3
rlabel polysilicon 415 -166 415 -166 0 1
rlabel polysilicon 415 -172 415 -172 0 3
rlabel polysilicon 422 -166 422 -166 0 1
rlabel polysilicon 422 -172 422 -172 0 3
rlabel polysilicon 429 -166 429 -166 0 1
rlabel polysilicon 429 -172 429 -172 0 3
rlabel polysilicon 436 -166 436 -166 0 1
rlabel polysilicon 436 -172 436 -172 0 3
rlabel polysilicon 443 -166 443 -166 0 1
rlabel polysilicon 443 -172 443 -172 0 3
rlabel polysilicon 450 -166 450 -166 0 1
rlabel polysilicon 453 -166 453 -166 0 2
rlabel polysilicon 450 -172 450 -172 0 3
rlabel polysilicon 457 -166 457 -166 0 1
rlabel polysilicon 457 -172 457 -172 0 3
rlabel polysilicon 464 -166 464 -166 0 1
rlabel polysilicon 464 -172 464 -172 0 3
rlabel polysilicon 471 -166 471 -166 0 1
rlabel polysilicon 471 -172 471 -172 0 3
rlabel polysilicon 478 -166 478 -166 0 1
rlabel polysilicon 478 -172 478 -172 0 3
rlabel polysilicon 485 -166 485 -166 0 1
rlabel polysilicon 485 -172 485 -172 0 3
rlabel polysilicon 492 -166 492 -166 0 1
rlabel polysilicon 492 -172 492 -172 0 3
rlabel polysilicon 499 -166 499 -166 0 1
rlabel polysilicon 502 -166 502 -166 0 2
rlabel polysilicon 499 -172 499 -172 0 3
rlabel polysilicon 506 -166 506 -166 0 1
rlabel polysilicon 506 -172 506 -172 0 3
rlabel polysilicon 513 -166 513 -166 0 1
rlabel polysilicon 516 -166 516 -166 0 2
rlabel polysilicon 513 -172 513 -172 0 3
rlabel polysilicon 523 -166 523 -166 0 2
rlabel polysilicon 520 -172 520 -172 0 3
rlabel polysilicon 523 -172 523 -172 0 4
rlabel polysilicon 527 -166 527 -166 0 1
rlabel polysilicon 530 -166 530 -166 0 2
rlabel polysilicon 530 -172 530 -172 0 4
rlabel polysilicon 534 -166 534 -166 0 1
rlabel polysilicon 534 -172 534 -172 0 3
rlabel polysilicon 541 -166 541 -166 0 1
rlabel polysilicon 541 -172 541 -172 0 3
rlabel polysilicon 548 -166 548 -166 0 1
rlabel polysilicon 548 -172 548 -172 0 3
rlabel polysilicon 555 -166 555 -166 0 1
rlabel polysilicon 558 -166 558 -166 0 2
rlabel polysilicon 558 -172 558 -172 0 4
rlabel polysilicon 562 -166 562 -166 0 1
rlabel polysilicon 562 -172 562 -172 0 3
rlabel polysilicon 569 -166 569 -166 0 1
rlabel polysilicon 572 -166 572 -166 0 2
rlabel polysilicon 569 -172 569 -172 0 3
rlabel polysilicon 576 -166 576 -166 0 1
rlabel polysilicon 576 -172 576 -172 0 3
rlabel polysilicon 583 -166 583 -166 0 1
rlabel polysilicon 583 -172 583 -172 0 3
rlabel polysilicon 593 -166 593 -166 0 2
rlabel polysilicon 593 -172 593 -172 0 4
rlabel polysilicon 597 -166 597 -166 0 1
rlabel polysilicon 597 -172 597 -172 0 3
rlabel polysilicon 604 -166 604 -166 0 1
rlabel polysilicon 607 -172 607 -172 0 4
rlabel polysilicon 611 -166 611 -166 0 1
rlabel polysilicon 614 -166 614 -166 0 2
rlabel polysilicon 611 -172 611 -172 0 3
rlabel polysilicon 618 -166 618 -166 0 1
rlabel polysilicon 618 -172 618 -172 0 3
rlabel polysilicon 625 -166 625 -166 0 1
rlabel polysilicon 625 -172 625 -172 0 3
rlabel polysilicon 632 -166 632 -166 0 1
rlabel polysilicon 632 -172 632 -172 0 3
rlabel polysilicon 639 -166 639 -166 0 1
rlabel polysilicon 639 -172 639 -172 0 3
rlabel polysilicon 646 -166 646 -166 0 1
rlabel polysilicon 646 -172 646 -172 0 3
rlabel polysilicon 653 -166 653 -166 0 1
rlabel polysilicon 656 -166 656 -166 0 2
rlabel polysilicon 656 -172 656 -172 0 4
rlabel polysilicon 660 -166 660 -166 0 1
rlabel polysilicon 660 -172 660 -172 0 3
rlabel polysilicon 667 -166 667 -166 0 1
rlabel polysilicon 667 -172 667 -172 0 3
rlabel polysilicon 674 -166 674 -166 0 1
rlabel polysilicon 674 -172 674 -172 0 3
rlabel polysilicon 681 -166 681 -166 0 1
rlabel polysilicon 681 -172 681 -172 0 3
rlabel polysilicon 688 -166 688 -166 0 1
rlabel polysilicon 688 -172 688 -172 0 3
rlabel polysilicon 695 -166 695 -166 0 1
rlabel polysilicon 695 -172 695 -172 0 3
rlabel polysilicon 702 -166 702 -166 0 1
rlabel polysilicon 702 -172 702 -172 0 3
rlabel polysilicon 709 -166 709 -166 0 1
rlabel polysilicon 709 -172 709 -172 0 3
rlabel polysilicon 716 -166 716 -166 0 1
rlabel polysilicon 716 -172 716 -172 0 3
rlabel polysilicon 723 -166 723 -166 0 1
rlabel polysilicon 723 -172 723 -172 0 3
rlabel polysilicon 730 -166 730 -166 0 1
rlabel polysilicon 737 -166 737 -166 0 1
rlabel polysilicon 737 -172 737 -172 0 3
rlabel polysilicon 744 -166 744 -166 0 1
rlabel polysilicon 744 -172 744 -172 0 3
rlabel polysilicon 751 -166 751 -166 0 1
rlabel polysilicon 751 -172 751 -172 0 3
rlabel polysilicon 758 -166 758 -166 0 1
rlabel polysilicon 758 -172 758 -172 0 3
rlabel polysilicon 765 -166 765 -166 0 1
rlabel polysilicon 765 -172 765 -172 0 3
rlabel polysilicon 772 -166 772 -166 0 1
rlabel polysilicon 772 -172 772 -172 0 3
rlabel polysilicon 779 -166 779 -166 0 1
rlabel polysilicon 779 -172 779 -172 0 3
rlabel polysilicon 786 -166 786 -166 0 1
rlabel polysilicon 786 -172 786 -172 0 3
rlabel polysilicon 793 -166 793 -166 0 1
rlabel polysilicon 793 -172 793 -172 0 3
rlabel polysilicon 800 -166 800 -166 0 1
rlabel polysilicon 800 -172 800 -172 0 3
rlabel polysilicon 807 -166 807 -166 0 1
rlabel polysilicon 807 -172 807 -172 0 3
rlabel polysilicon 814 -166 814 -166 0 1
rlabel polysilicon 814 -172 814 -172 0 3
rlabel polysilicon 821 -166 821 -166 0 1
rlabel polysilicon 821 -172 821 -172 0 3
rlabel polysilicon 828 -166 828 -166 0 1
rlabel polysilicon 828 -172 828 -172 0 3
rlabel polysilicon 835 -166 835 -166 0 1
rlabel polysilicon 835 -172 835 -172 0 3
rlabel polysilicon 842 -166 842 -166 0 1
rlabel polysilicon 842 -172 842 -172 0 3
rlabel polysilicon 849 -166 849 -166 0 1
rlabel polysilicon 849 -172 849 -172 0 3
rlabel polysilicon 856 -166 856 -166 0 1
rlabel polysilicon 856 -172 856 -172 0 3
rlabel polysilicon 863 -166 863 -166 0 1
rlabel polysilicon 863 -172 863 -172 0 3
rlabel polysilicon 870 -166 870 -166 0 1
rlabel polysilicon 870 -172 870 -172 0 3
rlabel polysilicon 877 -166 877 -166 0 1
rlabel polysilicon 877 -172 877 -172 0 3
rlabel polysilicon 898 -166 898 -166 0 1
rlabel polysilicon 898 -172 898 -172 0 3
rlabel polysilicon 919 -166 919 -166 0 1
rlabel polysilicon 919 -172 919 -172 0 3
rlabel polysilicon 940 -166 940 -166 0 1
rlabel polysilicon 940 -172 940 -172 0 3
rlabel polysilicon 1010 -166 1010 -166 0 1
rlabel polysilicon 1013 -166 1013 -166 0 2
rlabel polysilicon 1024 -166 1024 -166 0 1
rlabel polysilicon 1024 -172 1024 -172 0 3
rlabel polysilicon 1136 -166 1136 -166 0 1
rlabel polysilicon 1136 -172 1136 -172 0 3
rlabel polysilicon 1171 -166 1171 -166 0 1
rlabel polysilicon 1171 -172 1171 -172 0 3
rlabel polysilicon 72 -233 72 -233 0 1
rlabel polysilicon 72 -239 72 -239 0 3
rlabel polysilicon 79 -233 79 -233 0 1
rlabel polysilicon 79 -239 79 -239 0 3
rlabel polysilicon 86 -233 86 -233 0 1
rlabel polysilicon 86 -239 86 -239 0 3
rlabel polysilicon 93 -233 93 -233 0 1
rlabel polysilicon 93 -239 93 -239 0 3
rlabel polysilicon 100 -233 100 -233 0 1
rlabel polysilicon 100 -239 100 -239 0 3
rlabel polysilicon 107 -233 107 -233 0 1
rlabel polysilicon 107 -239 107 -239 0 3
rlabel polysilicon 114 -233 114 -233 0 1
rlabel polysilicon 114 -239 114 -239 0 3
rlabel polysilicon 121 -233 121 -233 0 1
rlabel polysilicon 121 -239 121 -239 0 3
rlabel polysilicon 128 -233 128 -233 0 1
rlabel polysilicon 128 -239 128 -239 0 3
rlabel polysilicon 135 -233 135 -233 0 1
rlabel polysilicon 135 -239 135 -239 0 3
rlabel polysilicon 142 -233 142 -233 0 1
rlabel polysilicon 142 -239 142 -239 0 3
rlabel polysilicon 149 -233 149 -233 0 1
rlabel polysilicon 149 -239 149 -239 0 3
rlabel polysilicon 156 -239 156 -239 0 3
rlabel polysilicon 159 -239 159 -239 0 4
rlabel polysilicon 163 -233 163 -233 0 1
rlabel polysilicon 163 -239 163 -239 0 3
rlabel polysilicon 170 -233 170 -233 0 1
rlabel polysilicon 170 -239 170 -239 0 3
rlabel polysilicon 177 -233 177 -233 0 1
rlabel polysilicon 177 -239 177 -239 0 3
rlabel polysilicon 184 -233 184 -233 0 1
rlabel polysilicon 184 -239 184 -239 0 3
rlabel polysilicon 191 -233 191 -233 0 1
rlabel polysilicon 191 -239 191 -239 0 3
rlabel polysilicon 198 -233 198 -233 0 1
rlabel polysilicon 198 -239 198 -239 0 3
rlabel polysilicon 205 -233 205 -233 0 1
rlabel polysilicon 208 -233 208 -233 0 2
rlabel polysilicon 205 -239 205 -239 0 3
rlabel polysilicon 208 -239 208 -239 0 4
rlabel polysilicon 212 -233 212 -233 0 1
rlabel polysilicon 212 -239 212 -239 0 3
rlabel polysilicon 219 -233 219 -233 0 1
rlabel polysilicon 222 -233 222 -233 0 2
rlabel polysilicon 219 -239 219 -239 0 3
rlabel polysilicon 229 -233 229 -233 0 2
rlabel polysilicon 226 -239 226 -239 0 3
rlabel polysilicon 233 -233 233 -233 0 1
rlabel polysilicon 236 -233 236 -233 0 2
rlabel polysilicon 236 -239 236 -239 0 4
rlabel polysilicon 243 -233 243 -233 0 2
rlabel polysilicon 243 -239 243 -239 0 4
rlabel polysilicon 247 -233 247 -233 0 1
rlabel polysilicon 247 -239 247 -239 0 3
rlabel polysilicon 254 -233 254 -233 0 1
rlabel polysilicon 254 -239 254 -239 0 3
rlabel polysilicon 257 -239 257 -239 0 4
rlabel polysilicon 261 -233 261 -233 0 1
rlabel polysilicon 261 -239 261 -239 0 3
rlabel polysilicon 268 -233 268 -233 0 1
rlabel polysilicon 268 -239 268 -239 0 3
rlabel polysilicon 275 -233 275 -233 0 1
rlabel polysilicon 275 -239 275 -239 0 3
rlabel polysilicon 282 -233 282 -233 0 1
rlabel polysilicon 282 -239 282 -239 0 3
rlabel polysilicon 289 -233 289 -233 0 1
rlabel polysilicon 289 -239 289 -239 0 3
rlabel polysilicon 296 -233 296 -233 0 1
rlabel polysilicon 296 -239 296 -239 0 3
rlabel polysilicon 303 -233 303 -233 0 1
rlabel polysilicon 303 -239 303 -239 0 3
rlabel polysilicon 310 -233 310 -233 0 1
rlabel polysilicon 310 -239 310 -239 0 3
rlabel polysilicon 317 -233 317 -233 0 1
rlabel polysilicon 317 -239 317 -239 0 3
rlabel polysilicon 324 -233 324 -233 0 1
rlabel polysilicon 324 -239 324 -239 0 3
rlabel polysilicon 331 -233 331 -233 0 1
rlabel polysilicon 331 -239 331 -239 0 3
rlabel polysilicon 338 -233 338 -233 0 1
rlabel polysilicon 338 -239 338 -239 0 3
rlabel polysilicon 345 -233 345 -233 0 1
rlabel polysilicon 345 -239 345 -239 0 3
rlabel polysilicon 352 -233 352 -233 0 1
rlabel polysilicon 352 -239 352 -239 0 3
rlabel polysilicon 359 -233 359 -233 0 1
rlabel polysilicon 359 -239 359 -239 0 3
rlabel polysilicon 366 -233 366 -233 0 1
rlabel polysilicon 366 -239 366 -239 0 3
rlabel polysilicon 369 -239 369 -239 0 4
rlabel polysilicon 373 -233 373 -233 0 1
rlabel polysilicon 373 -239 373 -239 0 3
rlabel polysilicon 380 -233 380 -233 0 1
rlabel polysilicon 380 -239 380 -239 0 3
rlabel polysilicon 387 -233 387 -233 0 1
rlabel polysilicon 387 -239 387 -239 0 3
rlabel polysilicon 394 -233 394 -233 0 1
rlabel polysilicon 394 -239 394 -239 0 3
rlabel polysilicon 401 -233 401 -233 0 1
rlabel polysilicon 401 -239 401 -239 0 3
rlabel polysilicon 408 -233 408 -233 0 1
rlabel polysilicon 411 -239 411 -239 0 4
rlabel polysilicon 415 -233 415 -233 0 1
rlabel polysilicon 415 -239 415 -239 0 3
rlabel polysilicon 422 -233 422 -233 0 1
rlabel polysilicon 422 -239 422 -239 0 3
rlabel polysilicon 429 -233 429 -233 0 1
rlabel polysilicon 432 -233 432 -233 0 2
rlabel polysilicon 429 -239 429 -239 0 3
rlabel polysilicon 436 -233 436 -233 0 1
rlabel polysilicon 436 -239 436 -239 0 3
rlabel polysilicon 443 -233 443 -233 0 1
rlabel polysilicon 446 -233 446 -233 0 2
rlabel polysilicon 446 -239 446 -239 0 4
rlabel polysilicon 450 -233 450 -233 0 1
rlabel polysilicon 453 -233 453 -233 0 2
rlabel polysilicon 450 -239 450 -239 0 3
rlabel polysilicon 453 -239 453 -239 0 4
rlabel polysilicon 457 -233 457 -233 0 1
rlabel polysilicon 457 -239 457 -239 0 3
rlabel polysilicon 464 -233 464 -233 0 1
rlabel polysilicon 464 -239 464 -239 0 3
rlabel polysilicon 471 -233 471 -233 0 1
rlabel polysilicon 471 -239 471 -239 0 3
rlabel polysilicon 478 -233 478 -233 0 1
rlabel polysilicon 478 -239 478 -239 0 3
rlabel polysilicon 481 -239 481 -239 0 4
rlabel polysilicon 485 -233 485 -233 0 1
rlabel polysilicon 485 -239 485 -239 0 3
rlabel polysilicon 488 -239 488 -239 0 4
rlabel polysilicon 492 -233 492 -233 0 1
rlabel polysilicon 492 -239 492 -239 0 3
rlabel polysilicon 499 -233 499 -233 0 1
rlabel polysilicon 499 -239 499 -239 0 3
rlabel polysilicon 502 -239 502 -239 0 4
rlabel polysilicon 506 -233 506 -233 0 1
rlabel polysilicon 506 -239 506 -239 0 3
rlabel polysilicon 513 -233 513 -233 0 1
rlabel polysilicon 513 -239 513 -239 0 3
rlabel polysilicon 520 -233 520 -233 0 1
rlabel polysilicon 520 -239 520 -239 0 3
rlabel polysilicon 527 -233 527 -233 0 1
rlabel polysilicon 527 -239 527 -239 0 3
rlabel polysilicon 534 -233 534 -233 0 1
rlabel polysilicon 534 -239 534 -239 0 3
rlabel polysilicon 541 -233 541 -233 0 1
rlabel polysilicon 541 -239 541 -239 0 3
rlabel polysilicon 551 -233 551 -233 0 2
rlabel polysilicon 551 -239 551 -239 0 4
rlabel polysilicon 555 -233 555 -233 0 1
rlabel polysilicon 555 -239 555 -239 0 3
rlabel polysilicon 562 -233 562 -233 0 1
rlabel polysilicon 562 -239 562 -239 0 3
rlabel polysilicon 569 -233 569 -233 0 1
rlabel polysilicon 569 -239 569 -239 0 3
rlabel polysilicon 576 -233 576 -233 0 1
rlabel polysilicon 576 -239 576 -239 0 3
rlabel polysilicon 583 -233 583 -233 0 1
rlabel polysilicon 583 -239 583 -239 0 3
rlabel polysilicon 590 -233 590 -233 0 1
rlabel polysilicon 590 -239 590 -239 0 3
rlabel polysilicon 597 -233 597 -233 0 1
rlabel polysilicon 597 -239 597 -239 0 3
rlabel polysilicon 604 -233 604 -233 0 1
rlabel polysilicon 604 -239 604 -239 0 3
rlabel polysilicon 611 -233 611 -233 0 1
rlabel polysilicon 614 -233 614 -233 0 2
rlabel polysilicon 611 -239 611 -239 0 3
rlabel polysilicon 618 -233 618 -233 0 1
rlabel polysilicon 618 -239 618 -239 0 3
rlabel polysilicon 625 -233 625 -233 0 1
rlabel polysilicon 628 -233 628 -233 0 2
rlabel polysilicon 628 -239 628 -239 0 4
rlabel polysilicon 632 -233 632 -233 0 1
rlabel polysilicon 632 -239 632 -239 0 3
rlabel polysilicon 639 -233 639 -233 0 1
rlabel polysilicon 639 -239 639 -239 0 3
rlabel polysilicon 646 -233 646 -233 0 1
rlabel polysilicon 646 -239 646 -239 0 3
rlabel polysilicon 653 -233 653 -233 0 1
rlabel polysilicon 653 -239 653 -239 0 3
rlabel polysilicon 660 -233 660 -233 0 1
rlabel polysilicon 660 -239 660 -239 0 3
rlabel polysilicon 667 -233 667 -233 0 1
rlabel polysilicon 667 -239 667 -239 0 3
rlabel polysilicon 674 -233 674 -233 0 1
rlabel polysilicon 674 -239 674 -239 0 3
rlabel polysilicon 681 -233 681 -233 0 1
rlabel polysilicon 681 -239 681 -239 0 3
rlabel polysilicon 688 -233 688 -233 0 1
rlabel polysilicon 688 -239 688 -239 0 3
rlabel polysilicon 695 -233 695 -233 0 1
rlabel polysilicon 695 -239 695 -239 0 3
rlabel polysilicon 702 -233 702 -233 0 1
rlabel polysilicon 702 -239 702 -239 0 3
rlabel polysilicon 709 -233 709 -233 0 1
rlabel polysilicon 709 -239 709 -239 0 3
rlabel polysilicon 716 -233 716 -233 0 1
rlabel polysilicon 716 -239 716 -239 0 3
rlabel polysilicon 723 -233 723 -233 0 1
rlabel polysilicon 723 -239 723 -239 0 3
rlabel polysilicon 730 -233 730 -233 0 1
rlabel polysilicon 730 -239 730 -239 0 3
rlabel polysilicon 737 -233 737 -233 0 1
rlabel polysilicon 737 -239 737 -239 0 3
rlabel polysilicon 744 -233 744 -233 0 1
rlabel polysilicon 744 -239 744 -239 0 3
rlabel polysilicon 751 -233 751 -233 0 1
rlabel polysilicon 754 -239 754 -239 0 4
rlabel polysilicon 758 -233 758 -233 0 1
rlabel polysilicon 758 -239 758 -239 0 3
rlabel polysilicon 765 -233 765 -233 0 1
rlabel polysilicon 765 -239 765 -239 0 3
rlabel polysilicon 772 -233 772 -233 0 1
rlabel polysilicon 772 -239 772 -239 0 3
rlabel polysilicon 779 -233 779 -233 0 1
rlabel polysilicon 779 -239 779 -239 0 3
rlabel polysilicon 786 -233 786 -233 0 1
rlabel polysilicon 786 -239 786 -239 0 3
rlabel polysilicon 793 -233 793 -233 0 1
rlabel polysilicon 793 -239 793 -239 0 3
rlabel polysilicon 800 -233 800 -233 0 1
rlabel polysilicon 800 -239 800 -239 0 3
rlabel polysilicon 807 -233 807 -233 0 1
rlabel polysilicon 807 -239 807 -239 0 3
rlabel polysilicon 814 -233 814 -233 0 1
rlabel polysilicon 814 -239 814 -239 0 3
rlabel polysilicon 821 -233 821 -233 0 1
rlabel polysilicon 821 -239 821 -239 0 3
rlabel polysilicon 831 -233 831 -233 0 2
rlabel polysilicon 828 -239 828 -239 0 3
rlabel polysilicon 835 -233 835 -233 0 1
rlabel polysilicon 835 -239 835 -239 0 3
rlabel polysilicon 842 -233 842 -233 0 1
rlabel polysilicon 842 -239 842 -239 0 3
rlabel polysilicon 849 -233 849 -233 0 1
rlabel polysilicon 849 -239 849 -239 0 3
rlabel polysilicon 856 -233 856 -233 0 1
rlabel polysilicon 856 -239 856 -239 0 3
rlabel polysilicon 863 -233 863 -233 0 1
rlabel polysilicon 863 -239 863 -239 0 3
rlabel polysilicon 870 -233 870 -233 0 1
rlabel polysilicon 870 -239 870 -239 0 3
rlabel polysilicon 877 -233 877 -233 0 1
rlabel polysilicon 877 -239 877 -239 0 3
rlabel polysilicon 884 -233 884 -233 0 1
rlabel polysilicon 884 -239 884 -239 0 3
rlabel polysilicon 891 -233 891 -233 0 1
rlabel polysilicon 891 -239 891 -239 0 3
rlabel polysilicon 898 -233 898 -233 0 1
rlabel polysilicon 898 -239 898 -239 0 3
rlabel polysilicon 905 -233 905 -233 0 1
rlabel polysilicon 905 -239 905 -239 0 3
rlabel polysilicon 912 -233 912 -233 0 1
rlabel polysilicon 912 -239 912 -239 0 3
rlabel polysilicon 919 -233 919 -233 0 1
rlabel polysilicon 919 -239 919 -239 0 3
rlabel polysilicon 926 -233 926 -233 0 1
rlabel polysilicon 926 -239 926 -239 0 3
rlabel polysilicon 933 -233 933 -233 0 1
rlabel polysilicon 933 -239 933 -239 0 3
rlabel polysilicon 940 -233 940 -233 0 1
rlabel polysilicon 940 -239 940 -239 0 3
rlabel polysilicon 947 -233 947 -233 0 1
rlabel polysilicon 947 -239 947 -239 0 3
rlabel polysilicon 954 -233 954 -233 0 1
rlabel polysilicon 954 -239 954 -239 0 3
rlabel polysilicon 961 -233 961 -233 0 1
rlabel polysilicon 961 -239 961 -239 0 3
rlabel polysilicon 968 -233 968 -233 0 1
rlabel polysilicon 968 -239 968 -239 0 3
rlabel polysilicon 975 -233 975 -233 0 1
rlabel polysilicon 975 -239 975 -239 0 3
rlabel polysilicon 982 -233 982 -233 0 1
rlabel polysilicon 982 -239 982 -239 0 3
rlabel polysilicon 989 -233 989 -233 0 1
rlabel polysilicon 989 -239 989 -239 0 3
rlabel polysilicon 996 -233 996 -233 0 1
rlabel polysilicon 996 -239 996 -239 0 3
rlabel polysilicon 1003 -233 1003 -233 0 1
rlabel polysilicon 1003 -239 1003 -239 0 3
rlabel polysilicon 1010 -233 1010 -233 0 1
rlabel polysilicon 1010 -239 1010 -239 0 3
rlabel polysilicon 1017 -233 1017 -233 0 1
rlabel polysilicon 1017 -239 1017 -239 0 3
rlabel polysilicon 1024 -233 1024 -233 0 1
rlabel polysilicon 1024 -239 1024 -239 0 3
rlabel polysilicon 1038 -233 1038 -233 0 1
rlabel polysilicon 1038 -239 1038 -239 0 3
rlabel polysilicon 1185 -233 1185 -233 0 1
rlabel polysilicon 1185 -239 1185 -239 0 3
rlabel polysilicon 1325 -233 1325 -233 0 1
rlabel polysilicon 1325 -239 1325 -239 0 3
rlabel polysilicon 65 -316 65 -316 0 1
rlabel polysilicon 65 -322 65 -322 0 3
rlabel polysilicon 72 -316 72 -316 0 1
rlabel polysilicon 72 -322 72 -322 0 3
rlabel polysilicon 79 -316 79 -316 0 1
rlabel polysilicon 79 -322 79 -322 0 3
rlabel polysilicon 86 -316 86 -316 0 1
rlabel polysilicon 86 -322 86 -322 0 3
rlabel polysilicon 93 -316 93 -316 0 1
rlabel polysilicon 93 -322 93 -322 0 3
rlabel polysilicon 100 -316 100 -316 0 1
rlabel polysilicon 100 -322 100 -322 0 3
rlabel polysilicon 107 -316 107 -316 0 1
rlabel polysilicon 107 -322 107 -322 0 3
rlabel polysilicon 114 -316 114 -316 0 1
rlabel polysilicon 114 -322 114 -322 0 3
rlabel polysilicon 121 -316 121 -316 0 1
rlabel polysilicon 121 -322 121 -322 0 3
rlabel polysilicon 128 -316 128 -316 0 1
rlabel polysilicon 128 -322 128 -322 0 3
rlabel polysilicon 138 -316 138 -316 0 2
rlabel polysilicon 138 -322 138 -322 0 4
rlabel polysilicon 142 -316 142 -316 0 1
rlabel polysilicon 145 -316 145 -316 0 2
rlabel polysilicon 142 -322 142 -322 0 3
rlabel polysilicon 149 -316 149 -316 0 1
rlabel polysilicon 149 -322 149 -322 0 3
rlabel polysilicon 156 -316 156 -316 0 1
rlabel polysilicon 156 -322 156 -322 0 3
rlabel polysilicon 163 -316 163 -316 0 1
rlabel polysilicon 163 -322 163 -322 0 3
rlabel polysilicon 170 -316 170 -316 0 1
rlabel polysilicon 173 -316 173 -316 0 2
rlabel polysilicon 170 -322 170 -322 0 3
rlabel polysilicon 173 -322 173 -322 0 4
rlabel polysilicon 177 -316 177 -316 0 1
rlabel polysilicon 177 -322 177 -322 0 3
rlabel polysilicon 184 -316 184 -316 0 1
rlabel polysilicon 187 -316 187 -316 0 2
rlabel polysilicon 184 -322 184 -322 0 3
rlabel polysilicon 187 -322 187 -322 0 4
rlabel polysilicon 191 -316 191 -316 0 1
rlabel polysilicon 191 -322 191 -322 0 3
rlabel polysilicon 198 -316 198 -316 0 1
rlabel polysilicon 198 -322 198 -322 0 3
rlabel polysilicon 208 -316 208 -316 0 2
rlabel polysilicon 205 -322 205 -322 0 3
rlabel polysilicon 208 -322 208 -322 0 4
rlabel polysilicon 212 -316 212 -316 0 1
rlabel polysilicon 212 -322 212 -322 0 3
rlabel polysilicon 219 -316 219 -316 0 1
rlabel polysilicon 219 -322 219 -322 0 3
rlabel polysilicon 226 -316 226 -316 0 1
rlabel polysilicon 226 -322 226 -322 0 3
rlabel polysilicon 233 -316 233 -316 0 1
rlabel polysilicon 233 -322 233 -322 0 3
rlabel polysilicon 240 -316 240 -316 0 1
rlabel polysilicon 240 -322 240 -322 0 3
rlabel polysilicon 247 -316 247 -316 0 1
rlabel polysilicon 247 -322 247 -322 0 3
rlabel polysilicon 254 -316 254 -316 0 1
rlabel polysilicon 254 -322 254 -322 0 3
rlabel polysilicon 261 -316 261 -316 0 1
rlabel polysilicon 261 -322 261 -322 0 3
rlabel polysilicon 268 -316 268 -316 0 1
rlabel polysilicon 268 -322 268 -322 0 3
rlabel polysilicon 275 -316 275 -316 0 1
rlabel polysilicon 275 -322 275 -322 0 3
rlabel polysilicon 282 -316 282 -316 0 1
rlabel polysilicon 282 -322 282 -322 0 3
rlabel polysilicon 289 -316 289 -316 0 1
rlabel polysilicon 289 -322 289 -322 0 3
rlabel polysilicon 296 -316 296 -316 0 1
rlabel polysilicon 296 -322 296 -322 0 3
rlabel polysilicon 303 -316 303 -316 0 1
rlabel polysilicon 303 -322 303 -322 0 3
rlabel polysilicon 310 -316 310 -316 0 1
rlabel polysilicon 310 -322 310 -322 0 3
rlabel polysilicon 313 -322 313 -322 0 4
rlabel polysilicon 317 -316 317 -316 0 1
rlabel polysilicon 317 -322 317 -322 0 3
rlabel polysilicon 324 -316 324 -316 0 1
rlabel polysilicon 324 -322 324 -322 0 3
rlabel polysilicon 331 -316 331 -316 0 1
rlabel polysilicon 331 -322 331 -322 0 3
rlabel polysilicon 338 -316 338 -316 0 1
rlabel polysilicon 338 -322 338 -322 0 3
rlabel polysilicon 345 -316 345 -316 0 1
rlabel polysilicon 345 -322 345 -322 0 3
rlabel polysilicon 352 -316 352 -316 0 1
rlabel polysilicon 352 -322 352 -322 0 3
rlabel polysilicon 359 -316 359 -316 0 1
rlabel polysilicon 359 -322 359 -322 0 3
rlabel polysilicon 366 -316 366 -316 0 1
rlabel polysilicon 366 -322 366 -322 0 3
rlabel polysilicon 373 -316 373 -316 0 1
rlabel polysilicon 376 -316 376 -316 0 2
rlabel polysilicon 376 -322 376 -322 0 4
rlabel polysilicon 380 -316 380 -316 0 1
rlabel polysilicon 383 -316 383 -316 0 2
rlabel polysilicon 383 -322 383 -322 0 4
rlabel polysilicon 387 -316 387 -316 0 1
rlabel polysilicon 390 -316 390 -316 0 2
rlabel polysilicon 387 -322 387 -322 0 3
rlabel polysilicon 390 -322 390 -322 0 4
rlabel polysilicon 394 -316 394 -316 0 1
rlabel polysilicon 394 -322 394 -322 0 3
rlabel polysilicon 401 -316 401 -316 0 1
rlabel polysilicon 401 -322 401 -322 0 3
rlabel polysilicon 408 -316 408 -316 0 1
rlabel polysilicon 408 -322 408 -322 0 3
rlabel polysilicon 415 -316 415 -316 0 1
rlabel polysilicon 415 -322 415 -322 0 3
rlabel polysilicon 422 -316 422 -316 0 1
rlabel polysilicon 422 -322 422 -322 0 3
rlabel polysilicon 429 -316 429 -316 0 1
rlabel polysilicon 429 -322 429 -322 0 3
rlabel polysilicon 436 -316 436 -316 0 1
rlabel polysilicon 436 -322 436 -322 0 3
rlabel polysilicon 443 -316 443 -316 0 1
rlabel polysilicon 446 -316 446 -316 0 2
rlabel polysilicon 443 -322 443 -322 0 3
rlabel polysilicon 446 -322 446 -322 0 4
rlabel polysilicon 450 -316 450 -316 0 1
rlabel polysilicon 450 -322 450 -322 0 3
rlabel polysilicon 457 -316 457 -316 0 1
rlabel polysilicon 457 -322 457 -322 0 3
rlabel polysilicon 464 -316 464 -316 0 1
rlabel polysilicon 464 -322 464 -322 0 3
rlabel polysilicon 471 -316 471 -316 0 1
rlabel polysilicon 471 -322 471 -322 0 3
rlabel polysilicon 478 -316 478 -316 0 1
rlabel polysilicon 481 -322 481 -322 0 4
rlabel polysilicon 485 -316 485 -316 0 1
rlabel polysilicon 485 -322 485 -322 0 3
rlabel polysilicon 492 -316 492 -316 0 1
rlabel polysilicon 492 -322 492 -322 0 3
rlabel polysilicon 499 -316 499 -316 0 1
rlabel polysilicon 499 -322 499 -322 0 3
rlabel polysilicon 506 -316 506 -316 0 1
rlabel polysilicon 506 -322 506 -322 0 3
rlabel polysilicon 513 -316 513 -316 0 1
rlabel polysilicon 513 -322 513 -322 0 3
rlabel polysilicon 520 -316 520 -316 0 1
rlabel polysilicon 520 -322 520 -322 0 3
rlabel polysilicon 527 -316 527 -316 0 1
rlabel polysilicon 527 -322 527 -322 0 3
rlabel polysilicon 534 -316 534 -316 0 1
rlabel polysilicon 537 -316 537 -316 0 2
rlabel polysilicon 534 -322 534 -322 0 3
rlabel polysilicon 537 -322 537 -322 0 4
rlabel polysilicon 541 -316 541 -316 0 1
rlabel polysilicon 541 -322 541 -322 0 3
rlabel polysilicon 548 -316 548 -316 0 1
rlabel polysilicon 551 -316 551 -316 0 2
rlabel polysilicon 548 -322 548 -322 0 3
rlabel polysilicon 551 -322 551 -322 0 4
rlabel polysilicon 555 -316 555 -316 0 1
rlabel polysilicon 555 -322 555 -322 0 3
rlabel polysilicon 562 -316 562 -316 0 1
rlabel polysilicon 562 -322 562 -322 0 3
rlabel polysilicon 569 -316 569 -316 0 1
rlabel polysilicon 569 -322 569 -322 0 3
rlabel polysilicon 576 -316 576 -316 0 1
rlabel polysilicon 576 -322 576 -322 0 3
rlabel polysilicon 583 -316 583 -316 0 1
rlabel polysilicon 583 -322 583 -322 0 3
rlabel polysilicon 590 -316 590 -316 0 1
rlabel polysilicon 590 -322 590 -322 0 3
rlabel polysilicon 593 -322 593 -322 0 4
rlabel polysilicon 597 -316 597 -316 0 1
rlabel polysilicon 600 -316 600 -316 0 2
rlabel polysilicon 597 -322 597 -322 0 3
rlabel polysilicon 600 -322 600 -322 0 4
rlabel polysilicon 604 -316 604 -316 0 1
rlabel polysilicon 607 -316 607 -316 0 2
rlabel polysilicon 604 -322 604 -322 0 3
rlabel polysilicon 611 -316 611 -316 0 1
rlabel polysilicon 611 -322 611 -322 0 3
rlabel polysilicon 618 -316 618 -316 0 1
rlabel polysilicon 618 -322 618 -322 0 3
rlabel polysilicon 625 -316 625 -316 0 1
rlabel polysilicon 628 -316 628 -316 0 2
rlabel polysilicon 625 -322 625 -322 0 3
rlabel polysilicon 628 -322 628 -322 0 4
rlabel polysilicon 632 -316 632 -316 0 1
rlabel polysilicon 632 -322 632 -322 0 3
rlabel polysilicon 639 -316 639 -316 0 1
rlabel polysilicon 639 -322 639 -322 0 3
rlabel polysilicon 646 -316 646 -316 0 1
rlabel polysilicon 649 -322 649 -322 0 4
rlabel polysilicon 653 -316 653 -316 0 1
rlabel polysilicon 653 -322 653 -322 0 3
rlabel polysilicon 660 -316 660 -316 0 1
rlabel polysilicon 660 -322 660 -322 0 3
rlabel polysilicon 667 -316 667 -316 0 1
rlabel polysilicon 670 -316 670 -316 0 2
rlabel polysilicon 670 -322 670 -322 0 4
rlabel polysilicon 674 -316 674 -316 0 1
rlabel polysilicon 674 -322 674 -322 0 3
rlabel polysilicon 681 -316 681 -316 0 1
rlabel polysilicon 681 -322 681 -322 0 3
rlabel polysilicon 688 -316 688 -316 0 1
rlabel polysilicon 688 -322 688 -322 0 3
rlabel polysilicon 695 -316 695 -316 0 1
rlabel polysilicon 695 -322 695 -322 0 3
rlabel polysilicon 702 -316 702 -316 0 1
rlabel polysilicon 702 -322 702 -322 0 3
rlabel polysilicon 709 -316 709 -316 0 1
rlabel polysilicon 709 -322 709 -322 0 3
rlabel polysilicon 716 -316 716 -316 0 1
rlabel polysilicon 716 -322 716 -322 0 3
rlabel polysilicon 723 -316 723 -316 0 1
rlabel polysilicon 723 -322 723 -322 0 3
rlabel polysilicon 730 -316 730 -316 0 1
rlabel polysilicon 730 -322 730 -322 0 3
rlabel polysilicon 737 -316 737 -316 0 1
rlabel polysilicon 737 -322 737 -322 0 3
rlabel polysilicon 744 -316 744 -316 0 1
rlabel polysilicon 747 -316 747 -316 0 2
rlabel polysilicon 747 -322 747 -322 0 4
rlabel polysilicon 751 -316 751 -316 0 1
rlabel polysilicon 751 -322 751 -322 0 3
rlabel polysilicon 758 -316 758 -316 0 1
rlabel polysilicon 758 -322 758 -322 0 3
rlabel polysilicon 765 -316 765 -316 0 1
rlabel polysilicon 765 -322 765 -322 0 3
rlabel polysilicon 772 -316 772 -316 0 1
rlabel polysilicon 772 -322 772 -322 0 3
rlabel polysilicon 779 -316 779 -316 0 1
rlabel polysilicon 779 -322 779 -322 0 3
rlabel polysilicon 786 -316 786 -316 0 1
rlabel polysilicon 786 -322 786 -322 0 3
rlabel polysilicon 793 -316 793 -316 0 1
rlabel polysilicon 793 -322 793 -322 0 3
rlabel polysilicon 800 -316 800 -316 0 1
rlabel polysilicon 800 -322 800 -322 0 3
rlabel polysilicon 807 -316 807 -316 0 1
rlabel polysilicon 807 -322 807 -322 0 3
rlabel polysilicon 814 -316 814 -316 0 1
rlabel polysilicon 814 -322 814 -322 0 3
rlabel polysilicon 821 -316 821 -316 0 1
rlabel polysilicon 821 -322 821 -322 0 3
rlabel polysilicon 828 -316 828 -316 0 1
rlabel polysilicon 828 -322 828 -322 0 3
rlabel polysilicon 835 -316 835 -316 0 1
rlabel polysilicon 835 -322 835 -322 0 3
rlabel polysilicon 842 -316 842 -316 0 1
rlabel polysilicon 842 -322 842 -322 0 3
rlabel polysilicon 849 -316 849 -316 0 1
rlabel polysilicon 849 -322 849 -322 0 3
rlabel polysilicon 856 -316 856 -316 0 1
rlabel polysilicon 856 -322 856 -322 0 3
rlabel polysilicon 863 -316 863 -316 0 1
rlabel polysilicon 863 -322 863 -322 0 3
rlabel polysilicon 870 -316 870 -316 0 1
rlabel polysilicon 870 -322 870 -322 0 3
rlabel polysilicon 877 -316 877 -316 0 1
rlabel polysilicon 877 -322 877 -322 0 3
rlabel polysilicon 884 -316 884 -316 0 1
rlabel polysilicon 884 -322 884 -322 0 3
rlabel polysilicon 891 -316 891 -316 0 1
rlabel polysilicon 891 -322 891 -322 0 3
rlabel polysilicon 898 -316 898 -316 0 1
rlabel polysilicon 898 -322 898 -322 0 3
rlabel polysilicon 905 -316 905 -316 0 1
rlabel polysilicon 905 -322 905 -322 0 3
rlabel polysilicon 912 -316 912 -316 0 1
rlabel polysilicon 912 -322 912 -322 0 3
rlabel polysilicon 919 -316 919 -316 0 1
rlabel polysilicon 919 -322 919 -322 0 3
rlabel polysilicon 926 -316 926 -316 0 1
rlabel polysilicon 926 -322 926 -322 0 3
rlabel polysilicon 933 -316 933 -316 0 1
rlabel polysilicon 933 -322 933 -322 0 3
rlabel polysilicon 940 -316 940 -316 0 1
rlabel polysilicon 940 -322 940 -322 0 3
rlabel polysilicon 947 -316 947 -316 0 1
rlabel polysilicon 947 -322 947 -322 0 3
rlabel polysilicon 954 -316 954 -316 0 1
rlabel polysilicon 954 -322 954 -322 0 3
rlabel polysilicon 961 -316 961 -316 0 1
rlabel polysilicon 961 -322 961 -322 0 3
rlabel polysilicon 968 -316 968 -316 0 1
rlabel polysilicon 968 -322 968 -322 0 3
rlabel polysilicon 975 -316 975 -316 0 1
rlabel polysilicon 975 -322 975 -322 0 3
rlabel polysilicon 982 -316 982 -316 0 1
rlabel polysilicon 982 -322 982 -322 0 3
rlabel polysilicon 989 -316 989 -316 0 1
rlabel polysilicon 989 -322 989 -322 0 3
rlabel polysilicon 996 -316 996 -316 0 1
rlabel polysilicon 996 -322 996 -322 0 3
rlabel polysilicon 1003 -316 1003 -316 0 1
rlabel polysilicon 1003 -322 1003 -322 0 3
rlabel polysilicon 1010 -316 1010 -316 0 1
rlabel polysilicon 1010 -322 1010 -322 0 3
rlabel polysilicon 1017 -316 1017 -316 0 1
rlabel polysilicon 1017 -322 1017 -322 0 3
rlabel polysilicon 1024 -316 1024 -316 0 1
rlabel polysilicon 1024 -322 1024 -322 0 3
rlabel polysilicon 1031 -316 1031 -316 0 1
rlabel polysilicon 1031 -322 1031 -322 0 3
rlabel polysilicon 1038 -316 1038 -316 0 1
rlabel polysilicon 1038 -322 1038 -322 0 3
rlabel polysilicon 1045 -316 1045 -316 0 1
rlabel polysilicon 1045 -322 1045 -322 0 3
rlabel polysilicon 1052 -316 1052 -316 0 1
rlabel polysilicon 1052 -322 1052 -322 0 3
rlabel polysilicon 1059 -316 1059 -316 0 1
rlabel polysilicon 1059 -322 1059 -322 0 3
rlabel polysilicon 1066 -316 1066 -316 0 1
rlabel polysilicon 1066 -322 1066 -322 0 3
rlabel polysilicon 1073 -316 1073 -316 0 1
rlabel polysilicon 1073 -322 1073 -322 0 3
rlabel polysilicon 1080 -316 1080 -316 0 1
rlabel polysilicon 1080 -322 1080 -322 0 3
rlabel polysilicon 1087 -316 1087 -316 0 1
rlabel polysilicon 1087 -322 1087 -322 0 3
rlabel polysilicon 1094 -316 1094 -316 0 1
rlabel polysilicon 1094 -322 1094 -322 0 3
rlabel polysilicon 1101 -316 1101 -316 0 1
rlabel polysilicon 1101 -322 1101 -322 0 3
rlabel polysilicon 1108 -316 1108 -316 0 1
rlabel polysilicon 1108 -322 1108 -322 0 3
rlabel polysilicon 1115 -316 1115 -316 0 1
rlabel polysilicon 1115 -322 1115 -322 0 3
rlabel polysilicon 1122 -316 1122 -316 0 1
rlabel polysilicon 1122 -322 1122 -322 0 3
rlabel polysilicon 1206 -316 1206 -316 0 1
rlabel polysilicon 1206 -322 1206 -322 0 3
rlabel polysilicon 1307 -316 1307 -316 0 2
rlabel polysilicon 1307 -322 1307 -322 0 4
rlabel polysilicon 1381 -316 1381 -316 0 1
rlabel polysilicon 1381 -322 1381 -322 0 3
rlabel polysilicon 1458 -316 1458 -316 0 1
rlabel polysilicon 1458 -322 1458 -322 0 3
rlabel polysilicon 58 -415 58 -415 0 1
rlabel polysilicon 72 -415 72 -415 0 1
rlabel polysilicon 72 -421 72 -421 0 3
rlabel polysilicon 79 -415 79 -415 0 1
rlabel polysilicon 79 -421 79 -421 0 3
rlabel polysilicon 86 -415 86 -415 0 1
rlabel polysilicon 86 -421 86 -421 0 3
rlabel polysilicon 93 -415 93 -415 0 1
rlabel polysilicon 93 -421 93 -421 0 3
rlabel polysilicon 100 -415 100 -415 0 1
rlabel polysilicon 100 -421 100 -421 0 3
rlabel polysilicon 107 -415 107 -415 0 1
rlabel polysilicon 107 -421 107 -421 0 3
rlabel polysilicon 114 -415 114 -415 0 1
rlabel polysilicon 114 -421 114 -421 0 3
rlabel polysilicon 121 -415 121 -415 0 1
rlabel polysilicon 121 -421 121 -421 0 3
rlabel polysilicon 128 -415 128 -415 0 1
rlabel polysilicon 128 -421 128 -421 0 3
rlabel polysilicon 135 -415 135 -415 0 1
rlabel polysilicon 135 -421 135 -421 0 3
rlabel polysilicon 142 -415 142 -415 0 1
rlabel polysilicon 142 -421 142 -421 0 3
rlabel polysilicon 149 -415 149 -415 0 1
rlabel polysilicon 149 -421 149 -421 0 3
rlabel polysilicon 152 -421 152 -421 0 4
rlabel polysilicon 156 -415 156 -415 0 1
rlabel polysilicon 156 -421 156 -421 0 3
rlabel polysilicon 166 -415 166 -415 0 2
rlabel polysilicon 163 -421 163 -421 0 3
rlabel polysilicon 166 -421 166 -421 0 4
rlabel polysilicon 173 -415 173 -415 0 2
rlabel polysilicon 173 -421 173 -421 0 4
rlabel polysilicon 177 -415 177 -415 0 1
rlabel polysilicon 177 -421 177 -421 0 3
rlabel polysilicon 184 -415 184 -415 0 1
rlabel polysilicon 187 -415 187 -415 0 2
rlabel polysilicon 187 -421 187 -421 0 4
rlabel polysilicon 194 -415 194 -415 0 2
rlabel polysilicon 191 -421 191 -421 0 3
rlabel polysilicon 194 -421 194 -421 0 4
rlabel polysilicon 198 -415 198 -415 0 1
rlabel polysilicon 198 -421 198 -421 0 3
rlabel polysilicon 205 -415 205 -415 0 1
rlabel polysilicon 205 -421 205 -421 0 3
rlabel polysilicon 212 -415 212 -415 0 1
rlabel polysilicon 212 -421 212 -421 0 3
rlabel polysilicon 219 -415 219 -415 0 1
rlabel polysilicon 219 -421 219 -421 0 3
rlabel polysilicon 226 -415 226 -415 0 1
rlabel polysilicon 226 -421 226 -421 0 3
rlabel polysilicon 233 -415 233 -415 0 1
rlabel polysilicon 233 -421 233 -421 0 3
rlabel polysilicon 240 -415 240 -415 0 1
rlabel polysilicon 240 -421 240 -421 0 3
rlabel polysilicon 247 -415 247 -415 0 1
rlabel polysilicon 250 -415 250 -415 0 2
rlabel polysilicon 247 -421 247 -421 0 3
rlabel polysilicon 250 -421 250 -421 0 4
rlabel polysilicon 254 -415 254 -415 0 1
rlabel polysilicon 254 -421 254 -421 0 3
rlabel polysilicon 261 -415 261 -415 0 1
rlabel polysilicon 261 -421 261 -421 0 3
rlabel polysilicon 268 -415 268 -415 0 1
rlabel polysilicon 268 -421 268 -421 0 3
rlabel polysilicon 275 -415 275 -415 0 1
rlabel polysilicon 275 -421 275 -421 0 3
rlabel polysilicon 282 -415 282 -415 0 1
rlabel polysilicon 282 -421 282 -421 0 3
rlabel polysilicon 289 -415 289 -415 0 1
rlabel polysilicon 289 -421 289 -421 0 3
rlabel polysilicon 296 -415 296 -415 0 1
rlabel polysilicon 296 -421 296 -421 0 3
rlabel polysilicon 303 -415 303 -415 0 1
rlabel polysilicon 303 -421 303 -421 0 3
rlabel polysilicon 310 -415 310 -415 0 1
rlabel polysilicon 310 -421 310 -421 0 3
rlabel polysilicon 317 -415 317 -415 0 1
rlabel polysilicon 317 -421 317 -421 0 3
rlabel polysilicon 324 -415 324 -415 0 1
rlabel polysilicon 324 -421 324 -421 0 3
rlabel polysilicon 331 -415 331 -415 0 1
rlabel polysilicon 331 -421 331 -421 0 3
rlabel polysilicon 338 -415 338 -415 0 1
rlabel polysilicon 338 -421 338 -421 0 3
rlabel polysilicon 345 -415 345 -415 0 1
rlabel polysilicon 345 -421 345 -421 0 3
rlabel polysilicon 352 -415 352 -415 0 1
rlabel polysilicon 352 -421 352 -421 0 3
rlabel polysilicon 362 -415 362 -415 0 2
rlabel polysilicon 359 -421 359 -421 0 3
rlabel polysilicon 362 -421 362 -421 0 4
rlabel polysilicon 369 -415 369 -415 0 2
rlabel polysilicon 366 -421 366 -421 0 3
rlabel polysilicon 369 -421 369 -421 0 4
rlabel polysilicon 373 -415 373 -415 0 1
rlabel polysilicon 373 -421 373 -421 0 3
rlabel polysilicon 380 -415 380 -415 0 1
rlabel polysilicon 383 -415 383 -415 0 2
rlabel polysilicon 380 -421 380 -421 0 3
rlabel polysilicon 383 -421 383 -421 0 4
rlabel polysilicon 387 -415 387 -415 0 1
rlabel polysilicon 387 -421 387 -421 0 3
rlabel polysilicon 394 -415 394 -415 0 1
rlabel polysilicon 394 -421 394 -421 0 3
rlabel polysilicon 401 -415 401 -415 0 1
rlabel polysilicon 401 -421 401 -421 0 3
rlabel polysilicon 408 -415 408 -415 0 1
rlabel polysilicon 408 -421 408 -421 0 3
rlabel polysilicon 415 -415 415 -415 0 1
rlabel polysilicon 418 -415 418 -415 0 2
rlabel polysilicon 415 -421 415 -421 0 3
rlabel polysilicon 418 -421 418 -421 0 4
rlabel polysilicon 422 -415 422 -415 0 1
rlabel polysilicon 422 -421 422 -421 0 3
rlabel polysilicon 429 -415 429 -415 0 1
rlabel polysilicon 429 -421 429 -421 0 3
rlabel polysilicon 436 -415 436 -415 0 1
rlabel polysilicon 436 -421 436 -421 0 3
rlabel polysilicon 443 -415 443 -415 0 1
rlabel polysilicon 443 -421 443 -421 0 3
rlabel polysilicon 450 -415 450 -415 0 1
rlabel polysilicon 450 -421 450 -421 0 3
rlabel polysilicon 457 -415 457 -415 0 1
rlabel polysilicon 457 -421 457 -421 0 3
rlabel polysilicon 464 -415 464 -415 0 1
rlabel polysilicon 464 -421 464 -421 0 3
rlabel polysilicon 471 -415 471 -415 0 1
rlabel polysilicon 471 -421 471 -421 0 3
rlabel polysilicon 478 -415 478 -415 0 1
rlabel polysilicon 478 -421 478 -421 0 3
rlabel polysilicon 485 -415 485 -415 0 1
rlabel polysilicon 485 -421 485 -421 0 3
rlabel polysilicon 492 -415 492 -415 0 1
rlabel polysilicon 495 -415 495 -415 0 2
rlabel polysilicon 495 -421 495 -421 0 4
rlabel polysilicon 499 -415 499 -415 0 1
rlabel polysilicon 499 -421 499 -421 0 3
rlabel polysilicon 506 -415 506 -415 0 1
rlabel polysilicon 506 -421 506 -421 0 3
rlabel polysilicon 513 -415 513 -415 0 1
rlabel polysilicon 513 -421 513 -421 0 3
rlabel polysilicon 520 -415 520 -415 0 1
rlabel polysilicon 520 -421 520 -421 0 3
rlabel polysilicon 527 -415 527 -415 0 1
rlabel polysilicon 527 -421 527 -421 0 3
rlabel polysilicon 534 -415 534 -415 0 1
rlabel polysilicon 534 -421 534 -421 0 3
rlabel polysilicon 541 -415 541 -415 0 1
rlabel polysilicon 541 -421 541 -421 0 3
rlabel polysilicon 544 -421 544 -421 0 4
rlabel polysilicon 548 -415 548 -415 0 1
rlabel polysilicon 548 -421 548 -421 0 3
rlabel polysilicon 555 -415 555 -415 0 1
rlabel polysilicon 555 -421 555 -421 0 3
rlabel polysilicon 565 -415 565 -415 0 2
rlabel polysilicon 562 -421 562 -421 0 3
rlabel polysilicon 569 -415 569 -415 0 1
rlabel polysilicon 572 -415 572 -415 0 2
rlabel polysilicon 569 -421 569 -421 0 3
rlabel polysilicon 572 -421 572 -421 0 4
rlabel polysilicon 576 -415 576 -415 0 1
rlabel polysilicon 576 -421 576 -421 0 3
rlabel polysilicon 583 -415 583 -415 0 1
rlabel polysilicon 586 -415 586 -415 0 2
rlabel polysilicon 583 -421 583 -421 0 3
rlabel polysilicon 586 -421 586 -421 0 4
rlabel polysilicon 590 -415 590 -415 0 1
rlabel polysilicon 590 -421 590 -421 0 3
rlabel polysilicon 597 -415 597 -415 0 1
rlabel polysilicon 597 -421 597 -421 0 3
rlabel polysilicon 604 -415 604 -415 0 1
rlabel polysilicon 604 -421 604 -421 0 3
rlabel polysilicon 611 -415 611 -415 0 1
rlabel polysilicon 611 -421 611 -421 0 3
rlabel polysilicon 618 -415 618 -415 0 1
rlabel polysilicon 618 -421 618 -421 0 3
rlabel polysilicon 625 -415 625 -415 0 1
rlabel polysilicon 625 -421 625 -421 0 3
rlabel polysilicon 628 -421 628 -421 0 4
rlabel polysilicon 632 -415 632 -415 0 1
rlabel polysilicon 635 -415 635 -415 0 2
rlabel polysilicon 632 -421 632 -421 0 3
rlabel polysilicon 639 -415 639 -415 0 1
rlabel polysilicon 639 -421 639 -421 0 3
rlabel polysilicon 646 -415 646 -415 0 1
rlabel polysilicon 646 -421 646 -421 0 3
rlabel polysilicon 653 -415 653 -415 0 1
rlabel polysilicon 653 -421 653 -421 0 3
rlabel polysilicon 660 -415 660 -415 0 1
rlabel polysilicon 660 -421 660 -421 0 3
rlabel polysilicon 667 -415 667 -415 0 1
rlabel polysilicon 667 -421 667 -421 0 3
rlabel polysilicon 674 -415 674 -415 0 1
rlabel polysilicon 674 -421 674 -421 0 3
rlabel polysilicon 681 -415 681 -415 0 1
rlabel polysilicon 681 -421 681 -421 0 3
rlabel polysilicon 688 -415 688 -415 0 1
rlabel polysilicon 691 -415 691 -415 0 2
rlabel polysilicon 688 -421 688 -421 0 3
rlabel polysilicon 691 -421 691 -421 0 4
rlabel polysilicon 695 -415 695 -415 0 1
rlabel polysilicon 695 -421 695 -421 0 3
rlabel polysilicon 702 -415 702 -415 0 1
rlabel polysilicon 702 -421 702 -421 0 3
rlabel polysilicon 709 -415 709 -415 0 1
rlabel polysilicon 709 -421 709 -421 0 3
rlabel polysilicon 716 -415 716 -415 0 1
rlabel polysilicon 719 -421 719 -421 0 4
rlabel polysilicon 723 -415 723 -415 0 1
rlabel polysilicon 723 -421 723 -421 0 3
rlabel polysilicon 726 -421 726 -421 0 4
rlabel polysilicon 730 -415 730 -415 0 1
rlabel polysilicon 730 -421 730 -421 0 3
rlabel polysilicon 737 -415 737 -415 0 1
rlabel polysilicon 737 -421 737 -421 0 3
rlabel polysilicon 744 -415 744 -415 0 1
rlabel polysilicon 744 -421 744 -421 0 3
rlabel polysilicon 751 -415 751 -415 0 1
rlabel polysilicon 751 -421 751 -421 0 3
rlabel polysilicon 758 -415 758 -415 0 1
rlabel polysilicon 758 -421 758 -421 0 3
rlabel polysilicon 765 -415 765 -415 0 1
rlabel polysilicon 765 -421 765 -421 0 3
rlabel polysilicon 772 -415 772 -415 0 1
rlabel polysilicon 772 -421 772 -421 0 3
rlabel polysilicon 779 -415 779 -415 0 1
rlabel polysilicon 779 -421 779 -421 0 3
rlabel polysilicon 786 -415 786 -415 0 1
rlabel polysilicon 789 -415 789 -415 0 2
rlabel polysilicon 789 -421 789 -421 0 4
rlabel polysilicon 793 -415 793 -415 0 1
rlabel polysilicon 793 -421 793 -421 0 3
rlabel polysilicon 800 -415 800 -415 0 1
rlabel polysilicon 800 -421 800 -421 0 3
rlabel polysilicon 807 -415 807 -415 0 1
rlabel polysilicon 807 -421 807 -421 0 3
rlabel polysilicon 814 -415 814 -415 0 1
rlabel polysilicon 814 -421 814 -421 0 3
rlabel polysilicon 821 -415 821 -415 0 1
rlabel polysilicon 821 -421 821 -421 0 3
rlabel polysilicon 828 -415 828 -415 0 1
rlabel polysilicon 828 -421 828 -421 0 3
rlabel polysilicon 835 -415 835 -415 0 1
rlabel polysilicon 835 -421 835 -421 0 3
rlabel polysilicon 838 -421 838 -421 0 4
rlabel polysilicon 842 -415 842 -415 0 1
rlabel polysilicon 842 -421 842 -421 0 3
rlabel polysilicon 849 -415 849 -415 0 1
rlabel polysilicon 849 -421 849 -421 0 3
rlabel polysilicon 856 -415 856 -415 0 1
rlabel polysilicon 856 -421 856 -421 0 3
rlabel polysilicon 863 -415 863 -415 0 1
rlabel polysilicon 863 -421 863 -421 0 3
rlabel polysilicon 870 -415 870 -415 0 1
rlabel polysilicon 870 -421 870 -421 0 3
rlabel polysilicon 877 -415 877 -415 0 1
rlabel polysilicon 877 -421 877 -421 0 3
rlabel polysilicon 884 -415 884 -415 0 1
rlabel polysilicon 884 -421 884 -421 0 3
rlabel polysilicon 891 -415 891 -415 0 1
rlabel polysilicon 891 -421 891 -421 0 3
rlabel polysilicon 898 -415 898 -415 0 1
rlabel polysilicon 898 -421 898 -421 0 3
rlabel polysilicon 905 -415 905 -415 0 1
rlabel polysilicon 905 -421 905 -421 0 3
rlabel polysilicon 912 -415 912 -415 0 1
rlabel polysilicon 912 -421 912 -421 0 3
rlabel polysilicon 919 -415 919 -415 0 1
rlabel polysilicon 919 -421 919 -421 0 3
rlabel polysilicon 926 -415 926 -415 0 1
rlabel polysilicon 926 -421 926 -421 0 3
rlabel polysilicon 933 -415 933 -415 0 1
rlabel polysilicon 933 -421 933 -421 0 3
rlabel polysilicon 940 -415 940 -415 0 1
rlabel polysilicon 940 -421 940 -421 0 3
rlabel polysilicon 947 -415 947 -415 0 1
rlabel polysilicon 947 -421 947 -421 0 3
rlabel polysilicon 954 -415 954 -415 0 1
rlabel polysilicon 954 -421 954 -421 0 3
rlabel polysilicon 961 -415 961 -415 0 1
rlabel polysilicon 961 -421 961 -421 0 3
rlabel polysilicon 968 -415 968 -415 0 1
rlabel polysilicon 968 -421 968 -421 0 3
rlabel polysilicon 975 -415 975 -415 0 1
rlabel polysilicon 975 -421 975 -421 0 3
rlabel polysilicon 982 -415 982 -415 0 1
rlabel polysilicon 982 -421 982 -421 0 3
rlabel polysilicon 989 -415 989 -415 0 1
rlabel polysilicon 989 -421 989 -421 0 3
rlabel polysilicon 996 -415 996 -415 0 1
rlabel polysilicon 996 -421 996 -421 0 3
rlabel polysilicon 1003 -415 1003 -415 0 1
rlabel polysilicon 1003 -421 1003 -421 0 3
rlabel polysilicon 1010 -415 1010 -415 0 1
rlabel polysilicon 1010 -421 1010 -421 0 3
rlabel polysilicon 1017 -415 1017 -415 0 1
rlabel polysilicon 1017 -421 1017 -421 0 3
rlabel polysilicon 1024 -415 1024 -415 0 1
rlabel polysilicon 1024 -421 1024 -421 0 3
rlabel polysilicon 1031 -415 1031 -415 0 1
rlabel polysilicon 1031 -421 1031 -421 0 3
rlabel polysilicon 1038 -415 1038 -415 0 1
rlabel polysilicon 1038 -421 1038 -421 0 3
rlabel polysilicon 1045 -415 1045 -415 0 1
rlabel polysilicon 1045 -421 1045 -421 0 3
rlabel polysilicon 1052 -415 1052 -415 0 1
rlabel polysilicon 1052 -421 1052 -421 0 3
rlabel polysilicon 1059 -415 1059 -415 0 1
rlabel polysilicon 1059 -421 1059 -421 0 3
rlabel polysilicon 1066 -415 1066 -415 0 1
rlabel polysilicon 1066 -421 1066 -421 0 3
rlabel polysilicon 1073 -415 1073 -415 0 1
rlabel polysilicon 1073 -421 1073 -421 0 3
rlabel polysilicon 1080 -415 1080 -415 0 1
rlabel polysilicon 1080 -421 1080 -421 0 3
rlabel polysilicon 1087 -415 1087 -415 0 1
rlabel polysilicon 1087 -421 1087 -421 0 3
rlabel polysilicon 1094 -415 1094 -415 0 1
rlabel polysilicon 1094 -421 1094 -421 0 3
rlabel polysilicon 1101 -415 1101 -415 0 1
rlabel polysilicon 1101 -421 1101 -421 0 3
rlabel polysilicon 1108 -415 1108 -415 0 1
rlabel polysilicon 1108 -421 1108 -421 0 3
rlabel polysilicon 1115 -415 1115 -415 0 1
rlabel polysilicon 1115 -421 1115 -421 0 3
rlabel polysilicon 1122 -415 1122 -415 0 1
rlabel polysilicon 1122 -421 1122 -421 0 3
rlabel polysilicon 1129 -415 1129 -415 0 1
rlabel polysilicon 1129 -421 1129 -421 0 3
rlabel polysilicon 1136 -415 1136 -415 0 1
rlabel polysilicon 1136 -421 1136 -421 0 3
rlabel polysilicon 1143 -415 1143 -415 0 1
rlabel polysilicon 1143 -421 1143 -421 0 3
rlabel polysilicon 1150 -415 1150 -415 0 1
rlabel polysilicon 1150 -421 1150 -421 0 3
rlabel polysilicon 1157 -415 1157 -415 0 1
rlabel polysilicon 1157 -421 1157 -421 0 3
rlabel polysilicon 1164 -415 1164 -415 0 1
rlabel polysilicon 1164 -421 1164 -421 0 3
rlabel polysilicon 1171 -415 1171 -415 0 1
rlabel polysilicon 1171 -421 1171 -421 0 3
rlabel polysilicon 1178 -415 1178 -415 0 1
rlabel polysilicon 1178 -421 1178 -421 0 3
rlabel polysilicon 1185 -415 1185 -415 0 1
rlabel polysilicon 1185 -421 1185 -421 0 3
rlabel polysilicon 1192 -415 1192 -415 0 1
rlabel polysilicon 1192 -421 1192 -421 0 3
rlabel polysilicon 1199 -415 1199 -415 0 1
rlabel polysilicon 1199 -421 1199 -421 0 3
rlabel polysilicon 1206 -415 1206 -415 0 1
rlabel polysilicon 1206 -421 1206 -421 0 3
rlabel polysilicon 1213 -415 1213 -415 0 1
rlabel polysilicon 1213 -421 1213 -421 0 3
rlabel polysilicon 1223 -415 1223 -415 0 2
rlabel polysilicon 1220 -421 1220 -421 0 3
rlabel polysilicon 1223 -421 1223 -421 0 4
rlabel polysilicon 1388 -415 1388 -415 0 1
rlabel polysilicon 1388 -421 1388 -421 0 3
rlabel polysilicon 1409 -415 1409 -415 0 1
rlabel polysilicon 1409 -421 1409 -421 0 3
rlabel polysilicon 1521 -415 1521 -415 0 1
rlabel polysilicon 1521 -421 1521 -421 0 3
rlabel polysilicon 51 -504 51 -504 0 1
rlabel polysilicon 51 -510 51 -510 0 3
rlabel polysilicon 58 -504 58 -504 0 1
rlabel polysilicon 58 -510 58 -510 0 3
rlabel polysilicon 65 -504 65 -504 0 1
rlabel polysilicon 65 -510 65 -510 0 3
rlabel polysilicon 72 -504 72 -504 0 1
rlabel polysilicon 72 -510 72 -510 0 3
rlabel polysilicon 79 -504 79 -504 0 1
rlabel polysilicon 79 -510 79 -510 0 3
rlabel polysilicon 86 -504 86 -504 0 1
rlabel polysilicon 86 -510 86 -510 0 3
rlabel polysilicon 93 -504 93 -504 0 1
rlabel polysilicon 93 -510 93 -510 0 3
rlabel polysilicon 100 -504 100 -504 0 1
rlabel polysilicon 100 -510 100 -510 0 3
rlabel polysilicon 107 -504 107 -504 0 1
rlabel polysilicon 107 -510 107 -510 0 3
rlabel polysilicon 114 -504 114 -504 0 1
rlabel polysilicon 114 -510 114 -510 0 3
rlabel polysilicon 121 -504 121 -504 0 1
rlabel polysilicon 124 -504 124 -504 0 2
rlabel polysilicon 124 -510 124 -510 0 4
rlabel polysilicon 128 -504 128 -504 0 1
rlabel polysilicon 128 -510 128 -510 0 3
rlabel polysilicon 135 -504 135 -504 0 1
rlabel polysilicon 138 -504 138 -504 0 2
rlabel polysilicon 142 -504 142 -504 0 1
rlabel polysilicon 145 -504 145 -504 0 2
rlabel polysilicon 142 -510 142 -510 0 3
rlabel polysilicon 145 -510 145 -510 0 4
rlabel polysilicon 149 -504 149 -504 0 1
rlabel polysilicon 149 -510 149 -510 0 3
rlabel polysilicon 156 -504 156 -504 0 1
rlabel polysilicon 156 -510 156 -510 0 3
rlabel polysilicon 163 -504 163 -504 0 1
rlabel polysilicon 166 -504 166 -504 0 2
rlabel polysilicon 163 -510 163 -510 0 3
rlabel polysilicon 166 -510 166 -510 0 4
rlabel polysilicon 170 -504 170 -504 0 1
rlabel polysilicon 170 -510 170 -510 0 3
rlabel polysilicon 177 -504 177 -504 0 1
rlabel polysilicon 177 -510 177 -510 0 3
rlabel polysilicon 184 -504 184 -504 0 1
rlabel polysilicon 184 -510 184 -510 0 3
rlabel polysilicon 191 -504 191 -504 0 1
rlabel polysilicon 194 -504 194 -504 0 2
rlabel polysilicon 191 -510 191 -510 0 3
rlabel polysilicon 194 -510 194 -510 0 4
rlabel polysilicon 198 -504 198 -504 0 1
rlabel polysilicon 198 -510 198 -510 0 3
rlabel polysilicon 205 -504 205 -504 0 1
rlabel polysilicon 205 -510 205 -510 0 3
rlabel polysilicon 212 -504 212 -504 0 1
rlabel polysilicon 212 -510 212 -510 0 3
rlabel polysilicon 219 -504 219 -504 0 1
rlabel polysilicon 219 -510 219 -510 0 3
rlabel polysilicon 226 -504 226 -504 0 1
rlabel polysilicon 226 -510 226 -510 0 3
rlabel polysilicon 233 -510 233 -510 0 3
rlabel polysilicon 240 -504 240 -504 0 1
rlabel polysilicon 240 -510 240 -510 0 3
rlabel polysilicon 247 -504 247 -504 0 1
rlabel polysilicon 247 -510 247 -510 0 3
rlabel polysilicon 254 -504 254 -504 0 1
rlabel polysilicon 257 -504 257 -504 0 2
rlabel polysilicon 261 -504 261 -504 0 1
rlabel polysilicon 261 -510 261 -510 0 3
rlabel polysilicon 268 -504 268 -504 0 1
rlabel polysilicon 268 -510 268 -510 0 3
rlabel polysilicon 275 -504 275 -504 0 1
rlabel polysilicon 275 -510 275 -510 0 3
rlabel polysilicon 282 -504 282 -504 0 1
rlabel polysilicon 282 -510 282 -510 0 3
rlabel polysilicon 289 -504 289 -504 0 1
rlabel polysilicon 289 -510 289 -510 0 3
rlabel polysilicon 296 -504 296 -504 0 1
rlabel polysilicon 299 -504 299 -504 0 2
rlabel polysilicon 296 -510 296 -510 0 3
rlabel polysilicon 299 -510 299 -510 0 4
rlabel polysilicon 303 -504 303 -504 0 1
rlabel polysilicon 303 -510 303 -510 0 3
rlabel polysilicon 310 -504 310 -504 0 1
rlabel polysilicon 310 -510 310 -510 0 3
rlabel polysilicon 317 -504 317 -504 0 1
rlabel polysilicon 317 -510 317 -510 0 3
rlabel polysilicon 324 -504 324 -504 0 1
rlabel polysilicon 324 -510 324 -510 0 3
rlabel polysilicon 331 -504 331 -504 0 1
rlabel polysilicon 331 -510 331 -510 0 3
rlabel polysilicon 338 -504 338 -504 0 1
rlabel polysilicon 338 -510 338 -510 0 3
rlabel polysilicon 345 -504 345 -504 0 1
rlabel polysilicon 345 -510 345 -510 0 3
rlabel polysilicon 352 -504 352 -504 0 1
rlabel polysilicon 352 -510 352 -510 0 3
rlabel polysilicon 359 -504 359 -504 0 1
rlabel polysilicon 359 -510 359 -510 0 3
rlabel polysilicon 366 -504 366 -504 0 1
rlabel polysilicon 366 -510 366 -510 0 3
rlabel polysilicon 373 -504 373 -504 0 1
rlabel polysilicon 373 -510 373 -510 0 3
rlabel polysilicon 380 -504 380 -504 0 1
rlabel polysilicon 380 -510 380 -510 0 3
rlabel polysilicon 387 -504 387 -504 0 1
rlabel polysilicon 390 -504 390 -504 0 2
rlabel polysilicon 387 -510 387 -510 0 3
rlabel polysilicon 390 -510 390 -510 0 4
rlabel polysilicon 394 -504 394 -504 0 1
rlabel polysilicon 394 -510 394 -510 0 3
rlabel polysilicon 404 -504 404 -504 0 2
rlabel polysilicon 404 -510 404 -510 0 4
rlabel polysilicon 408 -504 408 -504 0 1
rlabel polysilicon 408 -510 408 -510 0 3
rlabel polysilicon 415 -504 415 -504 0 1
rlabel polysilicon 415 -510 415 -510 0 3
rlabel polysilicon 422 -504 422 -504 0 1
rlabel polysilicon 425 -504 425 -504 0 2
rlabel polysilicon 422 -510 422 -510 0 3
rlabel polysilicon 425 -510 425 -510 0 4
rlabel polysilicon 429 -504 429 -504 0 1
rlabel polysilicon 429 -510 429 -510 0 3
rlabel polysilicon 436 -504 436 -504 0 1
rlabel polysilicon 436 -510 436 -510 0 3
rlabel polysilicon 443 -504 443 -504 0 1
rlabel polysilicon 443 -510 443 -510 0 3
rlabel polysilicon 450 -504 450 -504 0 1
rlabel polysilicon 450 -510 450 -510 0 3
rlabel polysilicon 457 -504 457 -504 0 1
rlabel polysilicon 457 -510 457 -510 0 3
rlabel polysilicon 464 -504 464 -504 0 1
rlabel polysilicon 467 -504 467 -504 0 2
rlabel polysilicon 464 -510 464 -510 0 3
rlabel polysilicon 467 -510 467 -510 0 4
rlabel polysilicon 471 -504 471 -504 0 1
rlabel polysilicon 471 -510 471 -510 0 3
rlabel polysilicon 478 -504 478 -504 0 1
rlabel polysilicon 478 -510 478 -510 0 3
rlabel polysilicon 485 -504 485 -504 0 1
rlabel polysilicon 485 -510 485 -510 0 3
rlabel polysilicon 492 -504 492 -504 0 1
rlabel polysilicon 492 -510 492 -510 0 3
rlabel polysilicon 499 -504 499 -504 0 1
rlabel polysilicon 499 -510 499 -510 0 3
rlabel polysilicon 506 -504 506 -504 0 1
rlabel polysilicon 506 -510 506 -510 0 3
rlabel polysilicon 513 -504 513 -504 0 1
rlabel polysilicon 513 -510 513 -510 0 3
rlabel polysilicon 520 -504 520 -504 0 1
rlabel polysilicon 520 -510 520 -510 0 3
rlabel polysilicon 527 -504 527 -504 0 1
rlabel polysilicon 527 -510 527 -510 0 3
rlabel polysilicon 534 -504 534 -504 0 1
rlabel polysilicon 534 -510 534 -510 0 3
rlabel polysilicon 541 -504 541 -504 0 1
rlabel polysilicon 541 -510 541 -510 0 3
rlabel polysilicon 548 -504 548 -504 0 1
rlabel polysilicon 551 -504 551 -504 0 2
rlabel polysilicon 555 -504 555 -504 0 1
rlabel polysilicon 558 -504 558 -504 0 2
rlabel polysilicon 555 -510 555 -510 0 3
rlabel polysilicon 562 -504 562 -504 0 1
rlabel polysilicon 562 -510 562 -510 0 3
rlabel polysilicon 569 -504 569 -504 0 1
rlabel polysilicon 569 -510 569 -510 0 3
rlabel polysilicon 576 -504 576 -504 0 1
rlabel polysilicon 576 -510 576 -510 0 3
rlabel polysilicon 583 -504 583 -504 0 1
rlabel polysilicon 583 -510 583 -510 0 3
rlabel polysilicon 590 -504 590 -504 0 1
rlabel polysilicon 593 -504 593 -504 0 2
rlabel polysilicon 590 -510 590 -510 0 3
rlabel polysilicon 593 -510 593 -510 0 4
rlabel polysilicon 597 -504 597 -504 0 1
rlabel polysilicon 597 -510 597 -510 0 3
rlabel polysilicon 604 -504 604 -504 0 1
rlabel polysilicon 604 -510 604 -510 0 3
rlabel polysilicon 611 -504 611 -504 0 1
rlabel polysilicon 611 -510 611 -510 0 3
rlabel polysilicon 618 -504 618 -504 0 1
rlabel polysilicon 621 -504 621 -504 0 2
rlabel polysilicon 618 -510 618 -510 0 3
rlabel polysilicon 621 -510 621 -510 0 4
rlabel polysilicon 625 -504 625 -504 0 1
rlabel polysilicon 625 -510 625 -510 0 3
rlabel polysilicon 632 -504 632 -504 0 1
rlabel polysilicon 632 -510 632 -510 0 3
rlabel polysilicon 639 -504 639 -504 0 1
rlabel polysilicon 639 -510 639 -510 0 3
rlabel polysilicon 649 -504 649 -504 0 2
rlabel polysilicon 646 -510 646 -510 0 3
rlabel polysilicon 649 -510 649 -510 0 4
rlabel polysilicon 653 -504 653 -504 0 1
rlabel polysilicon 656 -504 656 -504 0 2
rlabel polysilicon 653 -510 653 -510 0 3
rlabel polysilicon 656 -510 656 -510 0 4
rlabel polysilicon 663 -504 663 -504 0 2
rlabel polysilicon 660 -510 660 -510 0 3
rlabel polysilicon 663 -510 663 -510 0 4
rlabel polysilicon 667 -504 667 -504 0 1
rlabel polysilicon 667 -510 667 -510 0 3
rlabel polysilicon 674 -504 674 -504 0 1
rlabel polysilicon 674 -510 674 -510 0 3
rlabel polysilicon 681 -504 681 -504 0 1
rlabel polysilicon 684 -504 684 -504 0 2
rlabel polysilicon 684 -510 684 -510 0 4
rlabel polysilicon 688 -504 688 -504 0 1
rlabel polysilicon 688 -510 688 -510 0 3
rlabel polysilicon 698 -504 698 -504 0 2
rlabel polysilicon 695 -510 695 -510 0 3
rlabel polysilicon 698 -510 698 -510 0 4
rlabel polysilicon 702 -504 702 -504 0 1
rlabel polysilicon 702 -510 702 -510 0 3
rlabel polysilicon 709 -504 709 -504 0 1
rlabel polysilicon 709 -510 709 -510 0 3
rlabel polysilicon 716 -504 716 -504 0 1
rlabel polysilicon 716 -510 716 -510 0 3
rlabel polysilicon 723 -504 723 -504 0 1
rlabel polysilicon 723 -510 723 -510 0 3
rlabel polysilicon 730 -504 730 -504 0 1
rlabel polysilicon 730 -510 730 -510 0 3
rlabel polysilicon 737 -504 737 -504 0 1
rlabel polysilicon 737 -510 737 -510 0 3
rlabel polysilicon 744 -504 744 -504 0 1
rlabel polysilicon 744 -510 744 -510 0 3
rlabel polysilicon 751 -504 751 -504 0 1
rlabel polysilicon 754 -504 754 -504 0 2
rlabel polysilicon 751 -510 751 -510 0 3
rlabel polysilicon 754 -510 754 -510 0 4
rlabel polysilicon 758 -504 758 -504 0 1
rlabel polysilicon 758 -510 758 -510 0 3
rlabel polysilicon 765 -504 765 -504 0 1
rlabel polysilicon 765 -510 765 -510 0 3
rlabel polysilicon 772 -504 772 -504 0 1
rlabel polysilicon 772 -510 772 -510 0 3
rlabel polysilicon 779 -504 779 -504 0 1
rlabel polysilicon 779 -510 779 -510 0 3
rlabel polysilicon 786 -504 786 -504 0 1
rlabel polysilicon 786 -510 786 -510 0 3
rlabel polysilicon 793 -504 793 -504 0 1
rlabel polysilicon 793 -510 793 -510 0 3
rlabel polysilicon 800 -504 800 -504 0 1
rlabel polysilicon 800 -510 800 -510 0 3
rlabel polysilicon 807 -504 807 -504 0 1
rlabel polysilicon 807 -510 807 -510 0 3
rlabel polysilicon 814 -504 814 -504 0 1
rlabel polysilicon 814 -510 814 -510 0 3
rlabel polysilicon 821 -504 821 -504 0 1
rlabel polysilicon 824 -504 824 -504 0 2
rlabel polysilicon 821 -510 821 -510 0 3
rlabel polysilicon 824 -510 824 -510 0 4
rlabel polysilicon 828 -504 828 -504 0 1
rlabel polysilicon 828 -510 828 -510 0 3
rlabel polysilicon 835 -504 835 -504 0 1
rlabel polysilicon 835 -510 835 -510 0 3
rlabel polysilicon 845 -504 845 -504 0 2
rlabel polysilicon 842 -510 842 -510 0 3
rlabel polysilicon 845 -510 845 -510 0 4
rlabel polysilicon 852 -504 852 -504 0 2
rlabel polysilicon 852 -510 852 -510 0 4
rlabel polysilicon 856 -504 856 -504 0 1
rlabel polysilicon 856 -510 856 -510 0 3
rlabel polysilicon 863 -504 863 -504 0 1
rlabel polysilicon 863 -510 863 -510 0 3
rlabel polysilicon 870 -504 870 -504 0 1
rlabel polysilicon 870 -510 870 -510 0 3
rlabel polysilicon 877 -504 877 -504 0 1
rlabel polysilicon 877 -510 877 -510 0 3
rlabel polysilicon 884 -504 884 -504 0 1
rlabel polysilicon 884 -510 884 -510 0 3
rlabel polysilicon 891 -504 891 -504 0 1
rlabel polysilicon 891 -510 891 -510 0 3
rlabel polysilicon 898 -504 898 -504 0 1
rlabel polysilicon 898 -510 898 -510 0 3
rlabel polysilicon 905 -504 905 -504 0 1
rlabel polysilicon 905 -510 905 -510 0 3
rlabel polysilicon 912 -504 912 -504 0 1
rlabel polysilicon 912 -510 912 -510 0 3
rlabel polysilicon 919 -504 919 -504 0 1
rlabel polysilicon 919 -510 919 -510 0 3
rlabel polysilicon 926 -504 926 -504 0 1
rlabel polysilicon 926 -510 926 -510 0 3
rlabel polysilicon 933 -504 933 -504 0 1
rlabel polysilicon 933 -510 933 -510 0 3
rlabel polysilicon 940 -504 940 -504 0 1
rlabel polysilicon 940 -510 940 -510 0 3
rlabel polysilicon 947 -504 947 -504 0 1
rlabel polysilicon 947 -510 947 -510 0 3
rlabel polysilicon 954 -504 954 -504 0 1
rlabel polysilicon 954 -510 954 -510 0 3
rlabel polysilicon 961 -504 961 -504 0 1
rlabel polysilicon 961 -510 961 -510 0 3
rlabel polysilicon 968 -504 968 -504 0 1
rlabel polysilicon 968 -510 968 -510 0 3
rlabel polysilicon 975 -504 975 -504 0 1
rlabel polysilicon 975 -510 975 -510 0 3
rlabel polysilicon 982 -504 982 -504 0 1
rlabel polysilicon 982 -510 982 -510 0 3
rlabel polysilicon 989 -504 989 -504 0 1
rlabel polysilicon 989 -510 989 -510 0 3
rlabel polysilicon 996 -504 996 -504 0 1
rlabel polysilicon 996 -510 996 -510 0 3
rlabel polysilicon 1003 -504 1003 -504 0 1
rlabel polysilicon 1003 -510 1003 -510 0 3
rlabel polysilicon 1010 -504 1010 -504 0 1
rlabel polysilicon 1010 -510 1010 -510 0 3
rlabel polysilicon 1017 -504 1017 -504 0 1
rlabel polysilicon 1017 -510 1017 -510 0 3
rlabel polysilicon 1024 -504 1024 -504 0 1
rlabel polysilicon 1024 -510 1024 -510 0 3
rlabel polysilicon 1031 -504 1031 -504 0 1
rlabel polysilicon 1031 -510 1031 -510 0 3
rlabel polysilicon 1038 -504 1038 -504 0 1
rlabel polysilicon 1038 -510 1038 -510 0 3
rlabel polysilicon 1045 -504 1045 -504 0 1
rlabel polysilicon 1045 -510 1045 -510 0 3
rlabel polysilicon 1052 -504 1052 -504 0 1
rlabel polysilicon 1052 -510 1052 -510 0 3
rlabel polysilicon 1059 -504 1059 -504 0 1
rlabel polysilicon 1059 -510 1059 -510 0 3
rlabel polysilicon 1066 -504 1066 -504 0 1
rlabel polysilicon 1066 -510 1066 -510 0 3
rlabel polysilicon 1073 -504 1073 -504 0 1
rlabel polysilicon 1073 -510 1073 -510 0 3
rlabel polysilicon 1080 -504 1080 -504 0 1
rlabel polysilicon 1080 -510 1080 -510 0 3
rlabel polysilicon 1087 -504 1087 -504 0 1
rlabel polysilicon 1087 -510 1087 -510 0 3
rlabel polysilicon 1094 -504 1094 -504 0 1
rlabel polysilicon 1094 -510 1094 -510 0 3
rlabel polysilicon 1101 -504 1101 -504 0 1
rlabel polysilicon 1101 -510 1101 -510 0 3
rlabel polysilicon 1108 -504 1108 -504 0 1
rlabel polysilicon 1108 -510 1108 -510 0 3
rlabel polysilicon 1115 -504 1115 -504 0 1
rlabel polysilicon 1115 -510 1115 -510 0 3
rlabel polysilicon 1122 -504 1122 -504 0 1
rlabel polysilicon 1122 -510 1122 -510 0 3
rlabel polysilicon 1129 -504 1129 -504 0 1
rlabel polysilicon 1129 -510 1129 -510 0 3
rlabel polysilicon 1136 -504 1136 -504 0 1
rlabel polysilicon 1136 -510 1136 -510 0 3
rlabel polysilicon 1143 -504 1143 -504 0 1
rlabel polysilicon 1143 -510 1143 -510 0 3
rlabel polysilicon 1150 -504 1150 -504 0 1
rlabel polysilicon 1150 -510 1150 -510 0 3
rlabel polysilicon 1157 -504 1157 -504 0 1
rlabel polysilicon 1157 -510 1157 -510 0 3
rlabel polysilicon 1164 -504 1164 -504 0 1
rlabel polysilicon 1164 -510 1164 -510 0 3
rlabel polysilicon 1171 -504 1171 -504 0 1
rlabel polysilicon 1171 -510 1171 -510 0 3
rlabel polysilicon 1178 -504 1178 -504 0 1
rlabel polysilicon 1178 -510 1178 -510 0 3
rlabel polysilicon 1185 -504 1185 -504 0 1
rlabel polysilicon 1185 -510 1185 -510 0 3
rlabel polysilicon 1192 -504 1192 -504 0 1
rlabel polysilicon 1192 -510 1192 -510 0 3
rlabel polysilicon 1199 -504 1199 -504 0 1
rlabel polysilicon 1199 -510 1199 -510 0 3
rlabel polysilicon 1206 -504 1206 -504 0 1
rlabel polysilicon 1206 -510 1206 -510 0 3
rlabel polysilicon 1213 -504 1213 -504 0 1
rlabel polysilicon 1213 -510 1213 -510 0 3
rlabel polysilicon 1223 -510 1223 -510 0 4
rlabel polysilicon 1227 -504 1227 -504 0 1
rlabel polysilicon 1227 -510 1227 -510 0 3
rlabel polysilicon 1234 -504 1234 -504 0 1
rlabel polysilicon 1234 -510 1234 -510 0 3
rlabel polysilicon 1241 -504 1241 -504 0 1
rlabel polysilicon 1241 -510 1241 -510 0 3
rlabel polysilicon 1251 -504 1251 -504 0 2
rlabel polysilicon 1251 -510 1251 -510 0 4
rlabel polysilicon 1255 -504 1255 -504 0 1
rlabel polysilicon 1255 -510 1255 -510 0 3
rlabel polysilicon 1430 -504 1430 -504 0 1
rlabel polysilicon 1430 -510 1430 -510 0 3
rlabel polysilicon 1486 -504 1486 -504 0 1
rlabel polysilicon 1486 -510 1486 -510 0 3
rlabel polysilicon 1542 -504 1542 -504 0 1
rlabel polysilicon 1542 -510 1542 -510 0 3
rlabel polysilicon 44 -625 44 -625 0 1
rlabel polysilicon 44 -631 44 -631 0 3
rlabel polysilicon 51 -625 51 -625 0 1
rlabel polysilicon 51 -631 51 -631 0 3
rlabel polysilicon 58 -625 58 -625 0 1
rlabel polysilicon 58 -631 58 -631 0 3
rlabel polysilicon 65 -625 65 -625 0 1
rlabel polysilicon 65 -631 65 -631 0 3
rlabel polysilicon 72 -625 72 -625 0 1
rlabel polysilicon 72 -631 72 -631 0 3
rlabel polysilicon 79 -625 79 -625 0 1
rlabel polysilicon 79 -631 79 -631 0 3
rlabel polysilicon 86 -625 86 -625 0 1
rlabel polysilicon 86 -631 86 -631 0 3
rlabel polysilicon 93 -625 93 -625 0 1
rlabel polysilicon 93 -631 93 -631 0 3
rlabel polysilicon 100 -625 100 -625 0 1
rlabel polysilicon 100 -631 100 -631 0 3
rlabel polysilicon 107 -625 107 -625 0 1
rlabel polysilicon 110 -625 110 -625 0 2
rlabel polysilicon 107 -631 107 -631 0 3
rlabel polysilicon 114 -625 114 -625 0 1
rlabel polysilicon 114 -631 114 -631 0 3
rlabel polysilicon 121 -625 121 -625 0 1
rlabel polysilicon 121 -631 121 -631 0 3
rlabel polysilicon 128 -625 128 -625 0 1
rlabel polysilicon 128 -631 128 -631 0 3
rlabel polysilicon 135 -625 135 -625 0 1
rlabel polysilicon 135 -631 135 -631 0 3
rlabel polysilicon 142 -625 142 -625 0 1
rlabel polysilicon 142 -631 142 -631 0 3
rlabel polysilicon 149 -625 149 -625 0 1
rlabel polysilicon 149 -631 149 -631 0 3
rlabel polysilicon 156 -625 156 -625 0 1
rlabel polysilicon 156 -631 156 -631 0 3
rlabel polysilicon 163 -625 163 -625 0 1
rlabel polysilicon 163 -631 163 -631 0 3
rlabel polysilicon 170 -625 170 -625 0 1
rlabel polysilicon 170 -631 170 -631 0 3
rlabel polysilicon 177 -625 177 -625 0 1
rlabel polysilicon 177 -631 177 -631 0 3
rlabel polysilicon 184 -625 184 -625 0 1
rlabel polysilicon 184 -631 184 -631 0 3
rlabel polysilicon 191 -625 191 -625 0 1
rlabel polysilicon 191 -631 191 -631 0 3
rlabel polysilicon 198 -625 198 -625 0 1
rlabel polysilicon 198 -631 198 -631 0 3
rlabel polysilicon 201 -631 201 -631 0 4
rlabel polysilicon 205 -625 205 -625 0 1
rlabel polysilicon 205 -631 205 -631 0 3
rlabel polysilicon 212 -625 212 -625 0 1
rlabel polysilicon 212 -631 212 -631 0 3
rlabel polysilicon 219 -625 219 -625 0 1
rlabel polysilicon 219 -631 219 -631 0 3
rlabel polysilicon 226 -625 226 -625 0 1
rlabel polysilicon 226 -631 226 -631 0 3
rlabel polysilicon 233 -625 233 -625 0 1
rlabel polysilicon 236 -625 236 -625 0 2
rlabel polysilicon 233 -631 233 -631 0 3
rlabel polysilicon 240 -625 240 -625 0 1
rlabel polysilicon 240 -631 240 -631 0 3
rlabel polysilicon 243 -631 243 -631 0 4
rlabel polysilicon 247 -625 247 -625 0 1
rlabel polysilicon 247 -631 247 -631 0 3
rlabel polysilicon 254 -625 254 -625 0 1
rlabel polysilicon 254 -631 254 -631 0 3
rlabel polysilicon 261 -625 261 -625 0 1
rlabel polysilicon 264 -625 264 -625 0 2
rlabel polysilicon 261 -631 261 -631 0 3
rlabel polysilicon 264 -631 264 -631 0 4
rlabel polysilicon 268 -625 268 -625 0 1
rlabel polysilicon 268 -631 268 -631 0 3
rlabel polysilicon 275 -625 275 -625 0 1
rlabel polysilicon 275 -631 275 -631 0 3
rlabel polysilicon 282 -625 282 -625 0 1
rlabel polysilicon 282 -631 282 -631 0 3
rlabel polysilicon 289 -625 289 -625 0 1
rlabel polysilicon 292 -625 292 -625 0 2
rlabel polysilicon 289 -631 289 -631 0 3
rlabel polysilicon 296 -625 296 -625 0 1
rlabel polysilicon 296 -631 296 -631 0 3
rlabel polysilicon 303 -625 303 -625 0 1
rlabel polysilicon 303 -631 303 -631 0 3
rlabel polysilicon 310 -625 310 -625 0 1
rlabel polysilicon 310 -631 310 -631 0 3
rlabel polysilicon 317 -625 317 -625 0 1
rlabel polysilicon 317 -631 317 -631 0 3
rlabel polysilicon 324 -625 324 -625 0 1
rlabel polysilicon 327 -625 327 -625 0 2
rlabel polysilicon 324 -631 324 -631 0 3
rlabel polysilicon 327 -631 327 -631 0 4
rlabel polysilicon 331 -625 331 -625 0 1
rlabel polysilicon 331 -631 331 -631 0 3
rlabel polysilicon 338 -625 338 -625 0 1
rlabel polysilicon 338 -631 338 -631 0 3
rlabel polysilicon 345 -625 345 -625 0 1
rlabel polysilicon 345 -631 345 -631 0 3
rlabel polysilicon 352 -625 352 -625 0 1
rlabel polysilicon 355 -625 355 -625 0 2
rlabel polysilicon 352 -631 352 -631 0 3
rlabel polysilicon 355 -631 355 -631 0 4
rlabel polysilicon 359 -625 359 -625 0 1
rlabel polysilicon 359 -631 359 -631 0 3
rlabel polysilicon 366 -625 366 -625 0 1
rlabel polysilicon 366 -631 366 -631 0 3
rlabel polysilicon 373 -625 373 -625 0 1
rlabel polysilicon 373 -631 373 -631 0 3
rlabel polysilicon 380 -625 380 -625 0 1
rlabel polysilicon 380 -631 380 -631 0 3
rlabel polysilicon 387 -625 387 -625 0 1
rlabel polysilicon 390 -625 390 -625 0 2
rlabel polysilicon 387 -631 387 -631 0 3
rlabel polysilicon 394 -625 394 -625 0 1
rlabel polysilicon 394 -631 394 -631 0 3
rlabel polysilicon 401 -625 401 -625 0 1
rlabel polysilicon 401 -631 401 -631 0 3
rlabel polysilicon 408 -625 408 -625 0 1
rlabel polysilicon 408 -631 408 -631 0 3
rlabel polysilicon 415 -625 415 -625 0 1
rlabel polysilicon 415 -631 415 -631 0 3
rlabel polysilicon 422 -625 422 -625 0 1
rlabel polysilicon 425 -625 425 -625 0 2
rlabel polysilicon 422 -631 422 -631 0 3
rlabel polysilicon 425 -631 425 -631 0 4
rlabel polysilicon 429 -625 429 -625 0 1
rlabel polysilicon 429 -631 429 -631 0 3
rlabel polysilicon 436 -625 436 -625 0 1
rlabel polysilicon 436 -631 436 -631 0 3
rlabel polysilicon 443 -625 443 -625 0 1
rlabel polysilicon 443 -631 443 -631 0 3
rlabel polysilicon 450 -625 450 -625 0 1
rlabel polysilicon 450 -631 450 -631 0 3
rlabel polysilicon 457 -625 457 -625 0 1
rlabel polysilicon 460 -625 460 -625 0 2
rlabel polysilicon 457 -631 457 -631 0 3
rlabel polysilicon 460 -631 460 -631 0 4
rlabel polysilicon 464 -625 464 -625 0 1
rlabel polysilicon 464 -631 464 -631 0 3
rlabel polysilicon 471 -625 471 -625 0 1
rlabel polysilicon 471 -631 471 -631 0 3
rlabel polysilicon 478 -625 478 -625 0 1
rlabel polysilicon 481 -625 481 -625 0 2
rlabel polysilicon 478 -631 478 -631 0 3
rlabel polysilicon 481 -631 481 -631 0 4
rlabel polysilicon 485 -625 485 -625 0 1
rlabel polysilicon 485 -631 485 -631 0 3
rlabel polysilicon 492 -625 492 -625 0 1
rlabel polysilicon 495 -625 495 -625 0 2
rlabel polysilicon 492 -631 492 -631 0 3
rlabel polysilicon 499 -625 499 -625 0 1
rlabel polysilicon 499 -631 499 -631 0 3
rlabel polysilicon 506 -625 506 -625 0 1
rlabel polysilicon 506 -631 506 -631 0 3
rlabel polysilicon 513 -625 513 -625 0 1
rlabel polysilicon 513 -631 513 -631 0 3
rlabel polysilicon 520 -625 520 -625 0 1
rlabel polysilicon 520 -631 520 -631 0 3
rlabel polysilicon 527 -625 527 -625 0 1
rlabel polysilicon 527 -631 527 -631 0 3
rlabel polysilicon 534 -625 534 -625 0 1
rlabel polysilicon 534 -631 534 -631 0 3
rlabel polysilicon 541 -625 541 -625 0 1
rlabel polysilicon 541 -631 541 -631 0 3
rlabel polysilicon 548 -625 548 -625 0 1
rlabel polysilicon 548 -631 548 -631 0 3
rlabel polysilicon 555 -625 555 -625 0 1
rlabel polysilicon 555 -631 555 -631 0 3
rlabel polysilicon 562 -625 562 -625 0 1
rlabel polysilicon 562 -631 562 -631 0 3
rlabel polysilicon 569 -625 569 -625 0 1
rlabel polysilicon 569 -631 569 -631 0 3
rlabel polysilicon 576 -625 576 -625 0 1
rlabel polysilicon 576 -631 576 -631 0 3
rlabel polysilicon 583 -625 583 -625 0 1
rlabel polysilicon 583 -631 583 -631 0 3
rlabel polysilicon 590 -625 590 -625 0 1
rlabel polysilicon 590 -631 590 -631 0 3
rlabel polysilicon 597 -625 597 -625 0 1
rlabel polysilicon 597 -631 597 -631 0 3
rlabel polysilicon 604 -625 604 -625 0 1
rlabel polysilicon 607 -625 607 -625 0 2
rlabel polysilicon 604 -631 604 -631 0 3
rlabel polysilicon 607 -631 607 -631 0 4
rlabel polysilicon 611 -625 611 -625 0 1
rlabel polysilicon 611 -631 611 -631 0 3
rlabel polysilicon 618 -625 618 -625 0 1
rlabel polysilicon 618 -631 618 -631 0 3
rlabel polysilicon 625 -625 625 -625 0 1
rlabel polysilicon 625 -631 625 -631 0 3
rlabel polysilicon 632 -625 632 -625 0 1
rlabel polysilicon 632 -631 632 -631 0 3
rlabel polysilicon 639 -625 639 -625 0 1
rlabel polysilicon 642 -625 642 -625 0 2
rlabel polysilicon 642 -631 642 -631 0 4
rlabel polysilicon 646 -625 646 -625 0 1
rlabel polysilicon 649 -625 649 -625 0 2
rlabel polysilicon 653 -625 653 -625 0 1
rlabel polysilicon 653 -631 653 -631 0 3
rlabel polysilicon 660 -625 660 -625 0 1
rlabel polysilicon 660 -631 660 -631 0 3
rlabel polysilicon 667 -625 667 -625 0 1
rlabel polysilicon 667 -631 667 -631 0 3
rlabel polysilicon 674 -625 674 -625 0 1
rlabel polysilicon 674 -631 674 -631 0 3
rlabel polysilicon 681 -625 681 -625 0 1
rlabel polysilicon 684 -625 684 -625 0 2
rlabel polysilicon 681 -631 681 -631 0 3
rlabel polysilicon 684 -631 684 -631 0 4
rlabel polysilicon 688 -625 688 -625 0 1
rlabel polysilicon 688 -631 688 -631 0 3
rlabel polysilicon 695 -625 695 -625 0 1
rlabel polysilicon 698 -625 698 -625 0 2
rlabel polysilicon 698 -631 698 -631 0 4
rlabel polysilicon 702 -625 702 -625 0 1
rlabel polysilicon 702 -631 702 -631 0 3
rlabel polysilicon 709 -625 709 -625 0 1
rlabel polysilicon 709 -631 709 -631 0 3
rlabel polysilicon 716 -625 716 -625 0 1
rlabel polysilicon 716 -631 716 -631 0 3
rlabel polysilicon 723 -625 723 -625 0 1
rlabel polysilicon 723 -631 723 -631 0 3
rlabel polysilicon 730 -631 730 -631 0 3
rlabel polysilicon 733 -631 733 -631 0 4
rlabel polysilicon 737 -625 737 -625 0 1
rlabel polysilicon 737 -631 737 -631 0 3
rlabel polysilicon 744 -625 744 -625 0 1
rlabel polysilicon 747 -625 747 -625 0 2
rlabel polysilicon 744 -631 744 -631 0 3
rlabel polysilicon 751 -625 751 -625 0 1
rlabel polysilicon 751 -631 751 -631 0 3
rlabel polysilicon 758 -625 758 -625 0 1
rlabel polysilicon 761 -625 761 -625 0 2
rlabel polysilicon 758 -631 758 -631 0 3
rlabel polysilicon 761 -631 761 -631 0 4
rlabel polysilicon 765 -625 765 -625 0 1
rlabel polysilicon 765 -631 765 -631 0 3
rlabel polysilicon 772 -625 772 -625 0 1
rlabel polysilicon 772 -631 772 -631 0 3
rlabel polysilicon 779 -625 779 -625 0 1
rlabel polysilicon 779 -631 779 -631 0 3
rlabel polysilicon 789 -625 789 -625 0 2
rlabel polysilicon 786 -631 786 -631 0 3
rlabel polysilicon 789 -631 789 -631 0 4
rlabel polysilicon 793 -625 793 -625 0 1
rlabel polysilicon 793 -631 793 -631 0 3
rlabel polysilicon 803 -625 803 -625 0 2
rlabel polysilicon 800 -631 800 -631 0 3
rlabel polysilicon 807 -625 807 -625 0 1
rlabel polysilicon 807 -631 807 -631 0 3
rlabel polysilicon 814 -625 814 -625 0 1
rlabel polysilicon 814 -631 814 -631 0 3
rlabel polysilicon 821 -625 821 -625 0 1
rlabel polysilicon 821 -631 821 -631 0 3
rlabel polysilicon 828 -625 828 -625 0 1
rlabel polysilicon 828 -631 828 -631 0 3
rlabel polysilicon 835 -625 835 -625 0 1
rlabel polysilicon 835 -631 835 -631 0 3
rlabel polysilicon 845 -625 845 -625 0 2
rlabel polysilicon 842 -631 842 -631 0 3
rlabel polysilicon 845 -631 845 -631 0 4
rlabel polysilicon 849 -625 849 -625 0 1
rlabel polysilicon 849 -631 849 -631 0 3
rlabel polysilicon 856 -625 856 -625 0 1
rlabel polysilicon 856 -631 856 -631 0 3
rlabel polysilicon 863 -625 863 -625 0 1
rlabel polysilicon 863 -631 863 -631 0 3
rlabel polysilicon 870 -625 870 -625 0 1
rlabel polysilicon 873 -625 873 -625 0 2
rlabel polysilicon 873 -631 873 -631 0 4
rlabel polysilicon 877 -625 877 -625 0 1
rlabel polysilicon 877 -631 877 -631 0 3
rlabel polysilicon 884 -625 884 -625 0 1
rlabel polysilicon 884 -631 884 -631 0 3
rlabel polysilicon 891 -625 891 -625 0 1
rlabel polysilicon 891 -631 891 -631 0 3
rlabel polysilicon 898 -625 898 -625 0 1
rlabel polysilicon 898 -631 898 -631 0 3
rlabel polysilicon 905 -625 905 -625 0 1
rlabel polysilicon 905 -631 905 -631 0 3
rlabel polysilicon 912 -625 912 -625 0 1
rlabel polysilicon 912 -631 912 -631 0 3
rlabel polysilicon 919 -625 919 -625 0 1
rlabel polysilicon 919 -631 919 -631 0 3
rlabel polysilicon 926 -625 926 -625 0 1
rlabel polysilicon 926 -631 926 -631 0 3
rlabel polysilicon 933 -625 933 -625 0 1
rlabel polysilicon 933 -631 933 -631 0 3
rlabel polysilicon 940 -625 940 -625 0 1
rlabel polysilicon 940 -631 940 -631 0 3
rlabel polysilicon 947 -625 947 -625 0 1
rlabel polysilicon 947 -631 947 -631 0 3
rlabel polysilicon 954 -625 954 -625 0 1
rlabel polysilicon 954 -631 954 -631 0 3
rlabel polysilicon 961 -625 961 -625 0 1
rlabel polysilicon 961 -631 961 -631 0 3
rlabel polysilicon 968 -625 968 -625 0 1
rlabel polysilicon 968 -631 968 -631 0 3
rlabel polysilicon 975 -625 975 -625 0 1
rlabel polysilicon 975 -631 975 -631 0 3
rlabel polysilicon 982 -625 982 -625 0 1
rlabel polysilicon 982 -631 982 -631 0 3
rlabel polysilicon 989 -625 989 -625 0 1
rlabel polysilicon 989 -631 989 -631 0 3
rlabel polysilicon 996 -625 996 -625 0 1
rlabel polysilicon 996 -631 996 -631 0 3
rlabel polysilicon 1003 -625 1003 -625 0 1
rlabel polysilicon 1003 -631 1003 -631 0 3
rlabel polysilicon 1010 -625 1010 -625 0 1
rlabel polysilicon 1010 -631 1010 -631 0 3
rlabel polysilicon 1017 -625 1017 -625 0 1
rlabel polysilicon 1017 -631 1017 -631 0 3
rlabel polysilicon 1020 -631 1020 -631 0 4
rlabel polysilicon 1024 -625 1024 -625 0 1
rlabel polysilicon 1024 -631 1024 -631 0 3
rlabel polysilicon 1034 -625 1034 -625 0 2
rlabel polysilicon 1038 -625 1038 -625 0 1
rlabel polysilicon 1038 -631 1038 -631 0 3
rlabel polysilicon 1045 -625 1045 -625 0 1
rlabel polysilicon 1045 -631 1045 -631 0 3
rlabel polysilicon 1052 -625 1052 -625 0 1
rlabel polysilicon 1052 -631 1052 -631 0 3
rlabel polysilicon 1059 -625 1059 -625 0 1
rlabel polysilicon 1059 -631 1059 -631 0 3
rlabel polysilicon 1066 -625 1066 -625 0 1
rlabel polysilicon 1066 -631 1066 -631 0 3
rlabel polysilicon 1073 -625 1073 -625 0 1
rlabel polysilicon 1073 -631 1073 -631 0 3
rlabel polysilicon 1080 -625 1080 -625 0 1
rlabel polysilicon 1080 -631 1080 -631 0 3
rlabel polysilicon 1087 -625 1087 -625 0 1
rlabel polysilicon 1087 -631 1087 -631 0 3
rlabel polysilicon 1094 -625 1094 -625 0 1
rlabel polysilicon 1094 -631 1094 -631 0 3
rlabel polysilicon 1101 -625 1101 -625 0 1
rlabel polysilicon 1101 -631 1101 -631 0 3
rlabel polysilicon 1108 -625 1108 -625 0 1
rlabel polysilicon 1108 -631 1108 -631 0 3
rlabel polysilicon 1115 -625 1115 -625 0 1
rlabel polysilicon 1115 -631 1115 -631 0 3
rlabel polysilicon 1122 -625 1122 -625 0 1
rlabel polysilicon 1122 -631 1122 -631 0 3
rlabel polysilicon 1129 -625 1129 -625 0 1
rlabel polysilicon 1129 -631 1129 -631 0 3
rlabel polysilicon 1136 -625 1136 -625 0 1
rlabel polysilicon 1136 -631 1136 -631 0 3
rlabel polysilicon 1143 -625 1143 -625 0 1
rlabel polysilicon 1143 -631 1143 -631 0 3
rlabel polysilicon 1150 -625 1150 -625 0 1
rlabel polysilicon 1150 -631 1150 -631 0 3
rlabel polysilicon 1157 -625 1157 -625 0 1
rlabel polysilicon 1157 -631 1157 -631 0 3
rlabel polysilicon 1164 -625 1164 -625 0 1
rlabel polysilicon 1164 -631 1164 -631 0 3
rlabel polysilicon 1171 -625 1171 -625 0 1
rlabel polysilicon 1171 -631 1171 -631 0 3
rlabel polysilicon 1178 -625 1178 -625 0 1
rlabel polysilicon 1178 -631 1178 -631 0 3
rlabel polysilicon 1185 -625 1185 -625 0 1
rlabel polysilicon 1185 -631 1185 -631 0 3
rlabel polysilicon 1192 -625 1192 -625 0 1
rlabel polysilicon 1192 -631 1192 -631 0 3
rlabel polysilicon 1199 -625 1199 -625 0 1
rlabel polysilicon 1199 -631 1199 -631 0 3
rlabel polysilicon 1206 -625 1206 -625 0 1
rlabel polysilicon 1206 -631 1206 -631 0 3
rlabel polysilicon 1213 -625 1213 -625 0 1
rlabel polysilicon 1213 -631 1213 -631 0 3
rlabel polysilicon 1220 -625 1220 -625 0 1
rlabel polysilicon 1220 -631 1220 -631 0 3
rlabel polysilicon 1227 -625 1227 -625 0 1
rlabel polysilicon 1227 -631 1227 -631 0 3
rlabel polysilicon 1234 -625 1234 -625 0 1
rlabel polysilicon 1234 -631 1234 -631 0 3
rlabel polysilicon 1241 -625 1241 -625 0 1
rlabel polysilicon 1241 -631 1241 -631 0 3
rlabel polysilicon 1248 -625 1248 -625 0 1
rlabel polysilicon 1248 -631 1248 -631 0 3
rlabel polysilicon 1255 -625 1255 -625 0 1
rlabel polysilicon 1255 -631 1255 -631 0 3
rlabel polysilicon 1262 -625 1262 -625 0 1
rlabel polysilicon 1262 -631 1262 -631 0 3
rlabel polysilicon 1269 -625 1269 -625 0 1
rlabel polysilicon 1269 -631 1269 -631 0 3
rlabel polysilicon 1276 -625 1276 -625 0 1
rlabel polysilicon 1276 -631 1276 -631 0 3
rlabel polysilicon 1283 -625 1283 -625 0 1
rlabel polysilicon 1283 -631 1283 -631 0 3
rlabel polysilicon 1290 -625 1290 -625 0 1
rlabel polysilicon 1290 -631 1290 -631 0 3
rlabel polysilicon 1297 -625 1297 -625 0 1
rlabel polysilicon 1297 -631 1297 -631 0 3
rlabel polysilicon 1304 -625 1304 -625 0 1
rlabel polysilicon 1304 -631 1304 -631 0 3
rlabel polysilicon 1311 -625 1311 -625 0 1
rlabel polysilicon 1311 -631 1311 -631 0 3
rlabel polysilicon 1318 -625 1318 -625 0 1
rlabel polysilicon 1318 -631 1318 -631 0 3
rlabel polysilicon 1325 -625 1325 -625 0 1
rlabel polysilicon 1325 -631 1325 -631 0 3
rlabel polysilicon 1332 -625 1332 -625 0 1
rlabel polysilicon 1332 -631 1332 -631 0 3
rlabel polysilicon 1339 -625 1339 -625 0 1
rlabel polysilicon 1339 -631 1339 -631 0 3
rlabel polysilicon 1346 -625 1346 -625 0 1
rlabel polysilicon 1346 -631 1346 -631 0 3
rlabel polysilicon 1353 -625 1353 -625 0 1
rlabel polysilicon 1353 -631 1353 -631 0 3
rlabel polysilicon 1360 -625 1360 -625 0 1
rlabel polysilicon 1360 -631 1360 -631 0 3
rlabel polysilicon 1367 -625 1367 -625 0 1
rlabel polysilicon 1367 -631 1367 -631 0 3
rlabel polysilicon 1374 -625 1374 -625 0 1
rlabel polysilicon 1374 -631 1374 -631 0 3
rlabel polysilicon 1381 -625 1381 -625 0 1
rlabel polysilicon 1381 -631 1381 -631 0 3
rlabel polysilicon 1388 -625 1388 -625 0 1
rlabel polysilicon 1388 -631 1388 -631 0 3
rlabel polysilicon 1395 -625 1395 -625 0 1
rlabel polysilicon 1395 -631 1395 -631 0 3
rlabel polysilicon 1402 -625 1402 -625 0 1
rlabel polysilicon 1402 -631 1402 -631 0 3
rlabel polysilicon 1409 -625 1409 -625 0 1
rlabel polysilicon 1409 -631 1409 -631 0 3
rlabel polysilicon 1419 -625 1419 -625 0 2
rlabel polysilicon 1416 -631 1416 -631 0 3
rlabel polysilicon 1419 -631 1419 -631 0 4
rlabel polysilicon 1423 -625 1423 -625 0 1
rlabel polysilicon 1423 -631 1423 -631 0 3
rlabel polysilicon 1430 -625 1430 -625 0 1
rlabel polysilicon 1430 -631 1430 -631 0 3
rlabel polysilicon 1437 -625 1437 -625 0 1
rlabel polysilicon 1437 -631 1437 -631 0 3
rlabel polysilicon 1444 -625 1444 -625 0 1
rlabel polysilicon 1444 -631 1444 -631 0 3
rlabel polysilicon 1451 -625 1451 -625 0 1
rlabel polysilicon 1451 -631 1451 -631 0 3
rlabel polysilicon 1458 -625 1458 -625 0 1
rlabel polysilicon 1458 -631 1458 -631 0 3
rlabel polysilicon 1465 -625 1465 -625 0 1
rlabel polysilicon 1465 -631 1465 -631 0 3
rlabel polysilicon 1528 -625 1528 -625 0 1
rlabel polysilicon 1528 -631 1528 -631 0 3
rlabel polysilicon 1549 -625 1549 -625 0 1
rlabel polysilicon 1549 -631 1549 -631 0 3
rlabel polysilicon 1619 -625 1619 -625 0 1
rlabel polysilicon 1619 -631 1619 -631 0 3
rlabel polysilicon 44 -758 44 -758 0 1
rlabel polysilicon 44 -764 44 -764 0 3
rlabel polysilicon 51 -758 51 -758 0 1
rlabel polysilicon 51 -764 51 -764 0 3
rlabel polysilicon 58 -758 58 -758 0 1
rlabel polysilicon 61 -764 61 -764 0 4
rlabel polysilicon 68 -758 68 -758 0 2
rlabel polysilicon 65 -764 65 -764 0 3
rlabel polysilicon 72 -758 72 -758 0 1
rlabel polysilicon 72 -764 72 -764 0 3
rlabel polysilicon 79 -758 79 -758 0 1
rlabel polysilicon 79 -764 79 -764 0 3
rlabel polysilicon 86 -758 86 -758 0 1
rlabel polysilicon 86 -764 86 -764 0 3
rlabel polysilicon 93 -758 93 -758 0 1
rlabel polysilicon 93 -764 93 -764 0 3
rlabel polysilicon 100 -758 100 -758 0 1
rlabel polysilicon 100 -764 100 -764 0 3
rlabel polysilicon 107 -758 107 -758 0 1
rlabel polysilicon 107 -764 107 -764 0 3
rlabel polysilicon 114 -758 114 -758 0 1
rlabel polysilicon 117 -758 117 -758 0 2
rlabel polysilicon 117 -764 117 -764 0 4
rlabel polysilicon 121 -758 121 -758 0 1
rlabel polysilicon 121 -764 121 -764 0 3
rlabel polysilicon 128 -758 128 -758 0 1
rlabel polysilicon 128 -764 128 -764 0 3
rlabel polysilicon 135 -758 135 -758 0 1
rlabel polysilicon 135 -764 135 -764 0 3
rlabel polysilicon 142 -758 142 -758 0 1
rlabel polysilicon 142 -764 142 -764 0 3
rlabel polysilicon 149 -758 149 -758 0 1
rlabel polysilicon 149 -764 149 -764 0 3
rlabel polysilicon 156 -758 156 -758 0 1
rlabel polysilicon 159 -758 159 -758 0 2
rlabel polysilicon 156 -764 156 -764 0 3
rlabel polysilicon 159 -764 159 -764 0 4
rlabel polysilicon 163 -758 163 -758 0 1
rlabel polysilicon 163 -764 163 -764 0 3
rlabel polysilicon 170 -758 170 -758 0 1
rlabel polysilicon 170 -764 170 -764 0 3
rlabel polysilicon 177 -758 177 -758 0 1
rlabel polysilicon 177 -764 177 -764 0 3
rlabel polysilicon 184 -758 184 -758 0 1
rlabel polysilicon 184 -764 184 -764 0 3
rlabel polysilicon 191 -758 191 -758 0 1
rlabel polysilicon 191 -764 191 -764 0 3
rlabel polysilicon 198 -758 198 -758 0 1
rlabel polysilicon 198 -764 198 -764 0 3
rlabel polysilicon 205 -758 205 -758 0 1
rlabel polysilicon 205 -764 205 -764 0 3
rlabel polysilicon 208 -764 208 -764 0 4
rlabel polysilicon 212 -758 212 -758 0 1
rlabel polysilicon 212 -764 212 -764 0 3
rlabel polysilicon 219 -758 219 -758 0 1
rlabel polysilicon 222 -758 222 -758 0 2
rlabel polysilicon 226 -758 226 -758 0 1
rlabel polysilicon 226 -764 226 -764 0 3
rlabel polysilicon 233 -758 233 -758 0 1
rlabel polysilicon 233 -764 233 -764 0 3
rlabel polysilicon 240 -758 240 -758 0 1
rlabel polysilicon 240 -764 240 -764 0 3
rlabel polysilicon 247 -758 247 -758 0 1
rlabel polysilicon 247 -764 247 -764 0 3
rlabel polysilicon 254 -758 254 -758 0 1
rlabel polysilicon 257 -758 257 -758 0 2
rlabel polysilicon 261 -758 261 -758 0 1
rlabel polysilicon 261 -764 261 -764 0 3
rlabel polysilicon 268 -758 268 -758 0 1
rlabel polysilicon 268 -764 268 -764 0 3
rlabel polysilicon 275 -758 275 -758 0 1
rlabel polysilicon 275 -764 275 -764 0 3
rlabel polysilicon 282 -758 282 -758 0 1
rlabel polysilicon 282 -764 282 -764 0 3
rlabel polysilicon 289 -758 289 -758 0 1
rlabel polysilicon 289 -764 289 -764 0 3
rlabel polysilicon 296 -758 296 -758 0 1
rlabel polysilicon 296 -764 296 -764 0 3
rlabel polysilicon 303 -758 303 -758 0 1
rlabel polysilicon 303 -764 303 -764 0 3
rlabel polysilicon 310 -758 310 -758 0 1
rlabel polysilicon 310 -764 310 -764 0 3
rlabel polysilicon 317 -758 317 -758 0 1
rlabel polysilicon 317 -764 317 -764 0 3
rlabel polysilicon 324 -758 324 -758 0 1
rlabel polysilicon 324 -764 324 -764 0 3
rlabel polysilicon 331 -758 331 -758 0 1
rlabel polysilicon 334 -758 334 -758 0 2
rlabel polysilicon 331 -764 331 -764 0 3
rlabel polysilicon 338 -758 338 -758 0 1
rlabel polysilicon 338 -764 338 -764 0 3
rlabel polysilicon 345 -758 345 -758 0 1
rlabel polysilicon 345 -764 345 -764 0 3
rlabel polysilicon 352 -758 352 -758 0 1
rlabel polysilicon 352 -764 352 -764 0 3
rlabel polysilicon 359 -758 359 -758 0 1
rlabel polysilicon 359 -764 359 -764 0 3
rlabel polysilicon 366 -758 366 -758 0 1
rlabel polysilicon 366 -764 366 -764 0 3
rlabel polysilicon 373 -758 373 -758 0 1
rlabel polysilicon 373 -764 373 -764 0 3
rlabel polysilicon 380 -758 380 -758 0 1
rlabel polysilicon 380 -764 380 -764 0 3
rlabel polysilicon 387 -758 387 -758 0 1
rlabel polysilicon 387 -764 387 -764 0 3
rlabel polysilicon 394 -758 394 -758 0 1
rlabel polysilicon 394 -764 394 -764 0 3
rlabel polysilicon 401 -758 401 -758 0 1
rlabel polysilicon 401 -764 401 -764 0 3
rlabel polysilicon 408 -758 408 -758 0 1
rlabel polysilicon 408 -764 408 -764 0 3
rlabel polysilicon 415 -758 415 -758 0 1
rlabel polysilicon 415 -764 415 -764 0 3
rlabel polysilicon 422 -758 422 -758 0 1
rlabel polysilicon 422 -764 422 -764 0 3
rlabel polysilicon 429 -758 429 -758 0 1
rlabel polysilicon 432 -758 432 -758 0 2
rlabel polysilicon 429 -764 429 -764 0 3
rlabel polysilicon 432 -764 432 -764 0 4
rlabel polysilicon 436 -758 436 -758 0 1
rlabel polysilicon 436 -764 436 -764 0 3
rlabel polysilicon 443 -758 443 -758 0 1
rlabel polysilicon 443 -764 443 -764 0 3
rlabel polysilicon 450 -758 450 -758 0 1
rlabel polysilicon 450 -764 450 -764 0 3
rlabel polysilicon 457 -758 457 -758 0 1
rlabel polysilicon 457 -764 457 -764 0 3
rlabel polysilicon 464 -758 464 -758 0 1
rlabel polysilicon 467 -758 467 -758 0 2
rlabel polysilicon 464 -764 464 -764 0 3
rlabel polysilicon 471 -758 471 -758 0 1
rlabel polysilicon 471 -764 471 -764 0 3
rlabel polysilicon 478 -758 478 -758 0 1
rlabel polysilicon 478 -764 478 -764 0 3
rlabel polysilicon 485 -758 485 -758 0 1
rlabel polysilicon 485 -764 485 -764 0 3
rlabel polysilicon 492 -758 492 -758 0 1
rlabel polysilicon 495 -758 495 -758 0 2
rlabel polysilicon 492 -764 492 -764 0 3
rlabel polysilicon 499 -758 499 -758 0 1
rlabel polysilicon 499 -764 499 -764 0 3
rlabel polysilicon 506 -758 506 -758 0 1
rlabel polysilicon 506 -764 506 -764 0 3
rlabel polysilicon 513 -758 513 -758 0 1
rlabel polysilicon 513 -764 513 -764 0 3
rlabel polysilicon 523 -758 523 -758 0 2
rlabel polysilicon 520 -764 520 -764 0 3
rlabel polysilicon 523 -764 523 -764 0 4
rlabel polysilicon 527 -758 527 -758 0 1
rlabel polysilicon 530 -758 530 -758 0 2
rlabel polysilicon 527 -764 527 -764 0 3
rlabel polysilicon 530 -764 530 -764 0 4
rlabel polysilicon 534 -758 534 -758 0 1
rlabel polysilicon 534 -764 534 -764 0 3
rlabel polysilicon 541 -758 541 -758 0 1
rlabel polysilicon 541 -764 541 -764 0 3
rlabel polysilicon 548 -758 548 -758 0 1
rlabel polysilicon 548 -764 548 -764 0 3
rlabel polysilicon 555 -758 555 -758 0 1
rlabel polysilicon 558 -758 558 -758 0 2
rlabel polysilicon 555 -764 555 -764 0 3
rlabel polysilicon 558 -764 558 -764 0 4
rlabel polysilicon 562 -758 562 -758 0 1
rlabel polysilicon 562 -764 562 -764 0 3
rlabel polysilicon 569 -758 569 -758 0 1
rlabel polysilicon 572 -758 572 -758 0 2
rlabel polysilicon 572 -764 572 -764 0 4
rlabel polysilicon 576 -758 576 -758 0 1
rlabel polysilicon 576 -764 576 -764 0 3
rlabel polysilicon 583 -758 583 -758 0 1
rlabel polysilicon 583 -764 583 -764 0 3
rlabel polysilicon 590 -758 590 -758 0 1
rlabel polysilicon 590 -764 590 -764 0 3
rlabel polysilicon 597 -758 597 -758 0 1
rlabel polysilicon 597 -764 597 -764 0 3
rlabel polysilicon 604 -758 604 -758 0 1
rlabel polysilicon 607 -758 607 -758 0 2
rlabel polysilicon 604 -764 604 -764 0 3
rlabel polysilicon 607 -764 607 -764 0 4
rlabel polysilicon 611 -758 611 -758 0 1
rlabel polysilicon 611 -764 611 -764 0 3
rlabel polysilicon 618 -758 618 -758 0 1
rlabel polysilicon 618 -764 618 -764 0 3
rlabel polysilicon 625 -758 625 -758 0 1
rlabel polysilicon 625 -764 625 -764 0 3
rlabel polysilicon 632 -758 632 -758 0 1
rlabel polysilicon 635 -758 635 -758 0 2
rlabel polysilicon 635 -764 635 -764 0 4
rlabel polysilicon 639 -758 639 -758 0 1
rlabel polysilicon 639 -764 639 -764 0 3
rlabel polysilicon 646 -758 646 -758 0 1
rlabel polysilicon 649 -758 649 -758 0 2
rlabel polysilicon 646 -764 646 -764 0 3
rlabel polysilicon 649 -764 649 -764 0 4
rlabel polysilicon 653 -758 653 -758 0 1
rlabel polysilicon 653 -764 653 -764 0 3
rlabel polysilicon 660 -758 660 -758 0 1
rlabel polysilicon 660 -764 660 -764 0 3
rlabel polysilicon 667 -758 667 -758 0 1
rlabel polysilicon 667 -764 667 -764 0 3
rlabel polysilicon 674 -758 674 -758 0 1
rlabel polysilicon 677 -758 677 -758 0 2
rlabel polysilicon 674 -764 674 -764 0 3
rlabel polysilicon 677 -764 677 -764 0 4
rlabel polysilicon 681 -758 681 -758 0 1
rlabel polysilicon 681 -764 681 -764 0 3
rlabel polysilicon 691 -758 691 -758 0 2
rlabel polysilicon 688 -764 688 -764 0 3
rlabel polysilicon 691 -764 691 -764 0 4
rlabel polysilicon 695 -758 695 -758 0 1
rlabel polysilicon 695 -764 695 -764 0 3
rlabel polysilicon 702 -758 702 -758 0 1
rlabel polysilicon 702 -764 702 -764 0 3
rlabel polysilicon 709 -758 709 -758 0 1
rlabel polysilicon 709 -764 709 -764 0 3
rlabel polysilicon 716 -758 716 -758 0 1
rlabel polysilicon 719 -758 719 -758 0 2
rlabel polysilicon 716 -764 716 -764 0 3
rlabel polysilicon 719 -764 719 -764 0 4
rlabel polysilicon 723 -758 723 -758 0 1
rlabel polysilicon 723 -764 723 -764 0 3
rlabel polysilicon 733 -758 733 -758 0 2
rlabel polysilicon 730 -764 730 -764 0 3
rlabel polysilicon 737 -758 737 -758 0 1
rlabel polysilicon 737 -764 737 -764 0 3
rlabel polysilicon 744 -758 744 -758 0 1
rlabel polysilicon 744 -764 744 -764 0 3
rlabel polysilicon 751 -758 751 -758 0 1
rlabel polysilicon 751 -764 751 -764 0 3
rlabel polysilicon 758 -758 758 -758 0 1
rlabel polysilicon 758 -764 758 -764 0 3
rlabel polysilicon 765 -758 765 -758 0 1
rlabel polysilicon 765 -764 765 -764 0 3
rlabel polysilicon 772 -758 772 -758 0 1
rlabel polysilicon 772 -764 772 -764 0 3
rlabel polysilicon 779 -758 779 -758 0 1
rlabel polysilicon 779 -764 779 -764 0 3
rlabel polysilicon 786 -758 786 -758 0 1
rlabel polysilicon 786 -764 786 -764 0 3
rlabel polysilicon 796 -758 796 -758 0 2
rlabel polysilicon 793 -764 793 -764 0 3
rlabel polysilicon 796 -764 796 -764 0 4
rlabel polysilicon 800 -758 800 -758 0 1
rlabel polysilicon 803 -758 803 -758 0 2
rlabel polysilicon 800 -764 800 -764 0 3
rlabel polysilicon 807 -758 807 -758 0 1
rlabel polysilicon 807 -764 807 -764 0 3
rlabel polysilicon 814 -758 814 -758 0 1
rlabel polysilicon 814 -764 814 -764 0 3
rlabel polysilicon 821 -758 821 -758 0 1
rlabel polysilicon 821 -764 821 -764 0 3
rlabel polysilicon 828 -758 828 -758 0 1
rlabel polysilicon 831 -758 831 -758 0 2
rlabel polysilicon 828 -764 828 -764 0 3
rlabel polysilicon 831 -764 831 -764 0 4
rlabel polysilicon 835 -758 835 -758 0 1
rlabel polysilicon 838 -758 838 -758 0 2
rlabel polysilicon 835 -764 835 -764 0 3
rlabel polysilicon 838 -764 838 -764 0 4
rlabel polysilicon 842 -758 842 -758 0 1
rlabel polysilicon 842 -764 842 -764 0 3
rlabel polysilicon 849 -758 849 -758 0 1
rlabel polysilicon 849 -764 849 -764 0 3
rlabel polysilicon 856 -758 856 -758 0 1
rlabel polysilicon 856 -764 856 -764 0 3
rlabel polysilicon 863 -758 863 -758 0 1
rlabel polysilicon 863 -764 863 -764 0 3
rlabel polysilicon 870 -758 870 -758 0 1
rlabel polysilicon 870 -764 870 -764 0 3
rlabel polysilicon 873 -764 873 -764 0 4
rlabel polysilicon 877 -758 877 -758 0 1
rlabel polysilicon 877 -764 877 -764 0 3
rlabel polysilicon 884 -758 884 -758 0 1
rlabel polysilicon 884 -764 884 -764 0 3
rlabel polysilicon 891 -758 891 -758 0 1
rlabel polysilicon 891 -764 891 -764 0 3
rlabel polysilicon 898 -758 898 -758 0 1
rlabel polysilicon 898 -764 898 -764 0 3
rlabel polysilicon 905 -758 905 -758 0 1
rlabel polysilicon 908 -758 908 -758 0 2
rlabel polysilicon 905 -764 905 -764 0 3
rlabel polysilicon 908 -764 908 -764 0 4
rlabel polysilicon 912 -758 912 -758 0 1
rlabel polysilicon 912 -764 912 -764 0 3
rlabel polysilicon 919 -758 919 -758 0 1
rlabel polysilicon 919 -764 919 -764 0 3
rlabel polysilicon 929 -758 929 -758 0 2
rlabel polysilicon 926 -764 926 -764 0 3
rlabel polysilicon 929 -764 929 -764 0 4
rlabel polysilicon 933 -758 933 -758 0 1
rlabel polysilicon 933 -764 933 -764 0 3
rlabel polysilicon 940 -758 940 -758 0 1
rlabel polysilicon 940 -764 940 -764 0 3
rlabel polysilicon 947 -758 947 -758 0 1
rlabel polysilicon 947 -764 947 -764 0 3
rlabel polysilicon 954 -758 954 -758 0 1
rlabel polysilicon 954 -764 954 -764 0 3
rlabel polysilicon 961 -758 961 -758 0 1
rlabel polysilicon 961 -764 961 -764 0 3
rlabel polysilicon 968 -758 968 -758 0 1
rlabel polysilicon 968 -764 968 -764 0 3
rlabel polysilicon 975 -758 975 -758 0 1
rlabel polysilicon 975 -764 975 -764 0 3
rlabel polysilicon 982 -758 982 -758 0 1
rlabel polysilicon 982 -764 982 -764 0 3
rlabel polysilicon 989 -758 989 -758 0 1
rlabel polysilicon 989 -764 989 -764 0 3
rlabel polysilicon 996 -758 996 -758 0 1
rlabel polysilicon 996 -764 996 -764 0 3
rlabel polysilicon 1003 -758 1003 -758 0 1
rlabel polysilicon 1003 -764 1003 -764 0 3
rlabel polysilicon 1010 -758 1010 -758 0 1
rlabel polysilicon 1010 -764 1010 -764 0 3
rlabel polysilicon 1017 -758 1017 -758 0 1
rlabel polysilicon 1017 -764 1017 -764 0 3
rlabel polysilicon 1024 -758 1024 -758 0 1
rlabel polysilicon 1024 -764 1024 -764 0 3
rlabel polysilicon 1027 -764 1027 -764 0 4
rlabel polysilicon 1031 -758 1031 -758 0 1
rlabel polysilicon 1031 -764 1031 -764 0 3
rlabel polysilicon 1038 -758 1038 -758 0 1
rlabel polysilicon 1038 -764 1038 -764 0 3
rlabel polysilicon 1045 -758 1045 -758 0 1
rlabel polysilicon 1045 -764 1045 -764 0 3
rlabel polysilicon 1052 -758 1052 -758 0 1
rlabel polysilicon 1052 -764 1052 -764 0 3
rlabel polysilicon 1059 -758 1059 -758 0 1
rlabel polysilicon 1059 -764 1059 -764 0 3
rlabel polysilicon 1066 -758 1066 -758 0 1
rlabel polysilicon 1066 -764 1066 -764 0 3
rlabel polysilicon 1073 -758 1073 -758 0 1
rlabel polysilicon 1073 -764 1073 -764 0 3
rlabel polysilicon 1080 -758 1080 -758 0 1
rlabel polysilicon 1080 -764 1080 -764 0 3
rlabel polysilicon 1087 -758 1087 -758 0 1
rlabel polysilicon 1087 -764 1087 -764 0 3
rlabel polysilicon 1094 -758 1094 -758 0 1
rlabel polysilicon 1094 -764 1094 -764 0 3
rlabel polysilicon 1101 -758 1101 -758 0 1
rlabel polysilicon 1101 -764 1101 -764 0 3
rlabel polysilicon 1108 -758 1108 -758 0 1
rlabel polysilicon 1108 -764 1108 -764 0 3
rlabel polysilicon 1115 -758 1115 -758 0 1
rlabel polysilicon 1115 -764 1115 -764 0 3
rlabel polysilicon 1122 -758 1122 -758 0 1
rlabel polysilicon 1122 -764 1122 -764 0 3
rlabel polysilicon 1129 -758 1129 -758 0 1
rlabel polysilicon 1129 -764 1129 -764 0 3
rlabel polysilicon 1136 -758 1136 -758 0 1
rlabel polysilicon 1136 -764 1136 -764 0 3
rlabel polysilicon 1143 -758 1143 -758 0 1
rlabel polysilicon 1143 -764 1143 -764 0 3
rlabel polysilicon 1150 -758 1150 -758 0 1
rlabel polysilicon 1150 -764 1150 -764 0 3
rlabel polysilicon 1157 -758 1157 -758 0 1
rlabel polysilicon 1157 -764 1157 -764 0 3
rlabel polysilicon 1164 -758 1164 -758 0 1
rlabel polysilicon 1164 -764 1164 -764 0 3
rlabel polysilicon 1171 -758 1171 -758 0 1
rlabel polysilicon 1171 -764 1171 -764 0 3
rlabel polysilicon 1178 -758 1178 -758 0 1
rlabel polysilicon 1178 -764 1178 -764 0 3
rlabel polysilicon 1185 -758 1185 -758 0 1
rlabel polysilicon 1185 -764 1185 -764 0 3
rlabel polysilicon 1192 -758 1192 -758 0 1
rlabel polysilicon 1192 -764 1192 -764 0 3
rlabel polysilicon 1199 -758 1199 -758 0 1
rlabel polysilicon 1199 -764 1199 -764 0 3
rlabel polysilicon 1206 -758 1206 -758 0 1
rlabel polysilicon 1206 -764 1206 -764 0 3
rlabel polysilicon 1213 -758 1213 -758 0 1
rlabel polysilicon 1213 -764 1213 -764 0 3
rlabel polysilicon 1220 -758 1220 -758 0 1
rlabel polysilicon 1220 -764 1220 -764 0 3
rlabel polysilicon 1227 -758 1227 -758 0 1
rlabel polysilicon 1227 -764 1227 -764 0 3
rlabel polysilicon 1234 -758 1234 -758 0 1
rlabel polysilicon 1234 -764 1234 -764 0 3
rlabel polysilicon 1241 -758 1241 -758 0 1
rlabel polysilicon 1241 -764 1241 -764 0 3
rlabel polysilicon 1248 -758 1248 -758 0 1
rlabel polysilicon 1248 -764 1248 -764 0 3
rlabel polysilicon 1255 -758 1255 -758 0 1
rlabel polysilicon 1255 -764 1255 -764 0 3
rlabel polysilicon 1262 -758 1262 -758 0 1
rlabel polysilicon 1262 -764 1262 -764 0 3
rlabel polysilicon 1269 -758 1269 -758 0 1
rlabel polysilicon 1269 -764 1269 -764 0 3
rlabel polysilicon 1276 -758 1276 -758 0 1
rlabel polysilicon 1276 -764 1276 -764 0 3
rlabel polysilicon 1283 -758 1283 -758 0 1
rlabel polysilicon 1283 -764 1283 -764 0 3
rlabel polysilicon 1290 -758 1290 -758 0 1
rlabel polysilicon 1290 -764 1290 -764 0 3
rlabel polysilicon 1297 -758 1297 -758 0 1
rlabel polysilicon 1297 -764 1297 -764 0 3
rlabel polysilicon 1304 -758 1304 -758 0 1
rlabel polysilicon 1304 -764 1304 -764 0 3
rlabel polysilicon 1311 -758 1311 -758 0 1
rlabel polysilicon 1311 -764 1311 -764 0 3
rlabel polysilicon 1318 -758 1318 -758 0 1
rlabel polysilicon 1318 -764 1318 -764 0 3
rlabel polysilicon 1325 -758 1325 -758 0 1
rlabel polysilicon 1325 -764 1325 -764 0 3
rlabel polysilicon 1332 -758 1332 -758 0 1
rlabel polysilicon 1332 -764 1332 -764 0 3
rlabel polysilicon 1339 -758 1339 -758 0 1
rlabel polysilicon 1339 -764 1339 -764 0 3
rlabel polysilicon 1346 -758 1346 -758 0 1
rlabel polysilicon 1346 -764 1346 -764 0 3
rlabel polysilicon 1353 -758 1353 -758 0 1
rlabel polysilicon 1353 -764 1353 -764 0 3
rlabel polysilicon 1360 -758 1360 -758 0 1
rlabel polysilicon 1360 -764 1360 -764 0 3
rlabel polysilicon 1367 -758 1367 -758 0 1
rlabel polysilicon 1367 -764 1367 -764 0 3
rlabel polysilicon 1374 -758 1374 -758 0 1
rlabel polysilicon 1374 -764 1374 -764 0 3
rlabel polysilicon 1381 -758 1381 -758 0 1
rlabel polysilicon 1381 -764 1381 -764 0 3
rlabel polysilicon 1388 -758 1388 -758 0 1
rlabel polysilicon 1388 -764 1388 -764 0 3
rlabel polysilicon 1395 -758 1395 -758 0 1
rlabel polysilicon 1395 -764 1395 -764 0 3
rlabel polysilicon 1402 -758 1402 -758 0 1
rlabel polysilicon 1402 -764 1402 -764 0 3
rlabel polysilicon 1409 -758 1409 -758 0 1
rlabel polysilicon 1409 -764 1409 -764 0 3
rlabel polysilicon 1416 -758 1416 -758 0 1
rlabel polysilicon 1416 -764 1416 -764 0 3
rlabel polysilicon 1423 -758 1423 -758 0 1
rlabel polysilicon 1423 -764 1423 -764 0 3
rlabel polysilicon 1430 -758 1430 -758 0 1
rlabel polysilicon 1430 -764 1430 -764 0 3
rlabel polysilicon 1437 -758 1437 -758 0 1
rlabel polysilicon 1437 -764 1437 -764 0 3
rlabel polysilicon 1444 -758 1444 -758 0 1
rlabel polysilicon 1444 -764 1444 -764 0 3
rlabel polysilicon 1451 -758 1451 -758 0 1
rlabel polysilicon 1451 -764 1451 -764 0 3
rlabel polysilicon 1458 -758 1458 -758 0 1
rlabel polysilicon 1458 -764 1458 -764 0 3
rlabel polysilicon 1465 -758 1465 -758 0 1
rlabel polysilicon 1465 -764 1465 -764 0 3
rlabel polysilicon 1472 -758 1472 -758 0 1
rlabel polysilicon 1472 -764 1472 -764 0 3
rlabel polysilicon 1479 -758 1479 -758 0 1
rlabel polysilicon 1479 -764 1479 -764 0 3
rlabel polysilicon 1486 -758 1486 -758 0 1
rlabel polysilicon 1486 -764 1486 -764 0 3
rlabel polysilicon 1528 -758 1528 -758 0 1
rlabel polysilicon 1528 -764 1528 -764 0 3
rlabel polysilicon 1549 -758 1549 -758 0 1
rlabel polysilicon 1549 -764 1549 -764 0 3
rlabel polysilicon 1556 -758 1556 -758 0 1
rlabel polysilicon 1556 -764 1556 -764 0 3
rlabel polysilicon 1696 -758 1696 -758 0 1
rlabel polysilicon 1696 -764 1696 -764 0 3
rlabel polysilicon 37 -871 37 -871 0 1
rlabel polysilicon 37 -877 37 -877 0 3
rlabel polysilicon 44 -871 44 -871 0 1
rlabel polysilicon 44 -877 44 -877 0 3
rlabel polysilicon 51 -871 51 -871 0 1
rlabel polysilicon 51 -877 51 -877 0 3
rlabel polysilicon 58 -871 58 -871 0 1
rlabel polysilicon 58 -877 58 -877 0 3
rlabel polysilicon 65 -871 65 -871 0 1
rlabel polysilicon 65 -877 65 -877 0 3
rlabel polysilicon 72 -871 72 -871 0 1
rlabel polysilicon 72 -877 72 -877 0 3
rlabel polysilicon 79 -871 79 -871 0 1
rlabel polysilicon 79 -877 79 -877 0 3
rlabel polysilicon 86 -871 86 -871 0 1
rlabel polysilicon 86 -877 86 -877 0 3
rlabel polysilicon 93 -871 93 -871 0 1
rlabel polysilicon 93 -877 93 -877 0 3
rlabel polysilicon 100 -871 100 -871 0 1
rlabel polysilicon 100 -877 100 -877 0 3
rlabel polysilicon 107 -871 107 -871 0 1
rlabel polysilicon 107 -877 107 -877 0 3
rlabel polysilicon 110 -877 110 -877 0 4
rlabel polysilicon 114 -871 114 -871 0 1
rlabel polysilicon 114 -877 114 -877 0 3
rlabel polysilicon 121 -871 121 -871 0 1
rlabel polysilicon 124 -871 124 -871 0 2
rlabel polysilicon 121 -877 121 -877 0 3
rlabel polysilicon 124 -877 124 -877 0 4
rlabel polysilicon 128 -871 128 -871 0 1
rlabel polysilicon 128 -877 128 -877 0 3
rlabel polysilicon 135 -871 135 -871 0 1
rlabel polysilicon 135 -877 135 -877 0 3
rlabel polysilicon 142 -871 142 -871 0 1
rlabel polysilicon 142 -877 142 -877 0 3
rlabel polysilicon 149 -871 149 -871 0 1
rlabel polysilicon 152 -871 152 -871 0 2
rlabel polysilicon 149 -877 149 -877 0 3
rlabel polysilicon 156 -871 156 -871 0 1
rlabel polysilicon 156 -877 156 -877 0 3
rlabel polysilicon 163 -871 163 -871 0 1
rlabel polysilicon 166 -871 166 -871 0 2
rlabel polysilicon 163 -877 163 -877 0 3
rlabel polysilicon 166 -877 166 -877 0 4
rlabel polysilicon 170 -871 170 -871 0 1
rlabel polysilicon 170 -877 170 -877 0 3
rlabel polysilicon 177 -871 177 -871 0 1
rlabel polysilicon 177 -877 177 -877 0 3
rlabel polysilicon 184 -871 184 -871 0 1
rlabel polysilicon 187 -871 187 -871 0 2
rlabel polysilicon 184 -877 184 -877 0 3
rlabel polysilicon 191 -871 191 -871 0 1
rlabel polysilicon 191 -877 191 -877 0 3
rlabel polysilicon 198 -871 198 -871 0 1
rlabel polysilicon 198 -877 198 -877 0 3
rlabel polysilicon 205 -871 205 -871 0 1
rlabel polysilicon 208 -871 208 -871 0 2
rlabel polysilicon 205 -877 205 -877 0 3
rlabel polysilicon 208 -877 208 -877 0 4
rlabel polysilicon 212 -871 212 -871 0 1
rlabel polysilicon 212 -877 212 -877 0 3
rlabel polysilicon 222 -877 222 -877 0 4
rlabel polysilicon 226 -871 226 -871 0 1
rlabel polysilicon 226 -877 226 -877 0 3
rlabel polysilicon 233 -871 233 -871 0 1
rlabel polysilicon 233 -877 233 -877 0 3
rlabel polysilicon 240 -871 240 -871 0 1
rlabel polysilicon 240 -877 240 -877 0 3
rlabel polysilicon 247 -871 247 -871 0 1
rlabel polysilicon 247 -877 247 -877 0 3
rlabel polysilicon 254 -871 254 -871 0 1
rlabel polysilicon 254 -877 254 -877 0 3
rlabel polysilicon 257 -877 257 -877 0 4
rlabel polysilicon 261 -871 261 -871 0 1
rlabel polysilicon 261 -877 261 -877 0 3
rlabel polysilicon 268 -871 268 -871 0 1
rlabel polysilicon 268 -877 268 -877 0 3
rlabel polysilicon 275 -871 275 -871 0 1
rlabel polysilicon 275 -877 275 -877 0 3
rlabel polysilicon 282 -871 282 -871 0 1
rlabel polysilicon 282 -877 282 -877 0 3
rlabel polysilicon 289 -871 289 -871 0 1
rlabel polysilicon 289 -877 289 -877 0 3
rlabel polysilicon 296 -871 296 -871 0 1
rlabel polysilicon 296 -877 296 -877 0 3
rlabel polysilicon 303 -871 303 -871 0 1
rlabel polysilicon 303 -877 303 -877 0 3
rlabel polysilicon 310 -871 310 -871 0 1
rlabel polysilicon 310 -877 310 -877 0 3
rlabel polysilicon 317 -871 317 -871 0 1
rlabel polysilicon 317 -877 317 -877 0 3
rlabel polysilicon 324 -871 324 -871 0 1
rlabel polysilicon 331 -871 331 -871 0 1
rlabel polysilicon 331 -877 331 -877 0 3
rlabel polysilicon 338 -871 338 -871 0 1
rlabel polysilicon 338 -877 338 -877 0 3
rlabel polysilicon 345 -871 345 -871 0 1
rlabel polysilicon 345 -877 345 -877 0 3
rlabel polysilicon 352 -871 352 -871 0 1
rlabel polysilicon 352 -877 352 -877 0 3
rlabel polysilicon 359 -871 359 -871 0 1
rlabel polysilicon 359 -877 359 -877 0 3
rlabel polysilicon 366 -871 366 -871 0 1
rlabel polysilicon 366 -877 366 -877 0 3
rlabel polysilicon 373 -871 373 -871 0 1
rlabel polysilicon 373 -877 373 -877 0 3
rlabel polysilicon 380 -871 380 -871 0 1
rlabel polysilicon 380 -877 380 -877 0 3
rlabel polysilicon 387 -871 387 -871 0 1
rlabel polysilicon 387 -877 387 -877 0 3
rlabel polysilicon 394 -871 394 -871 0 1
rlabel polysilicon 394 -877 394 -877 0 3
rlabel polysilicon 401 -871 401 -871 0 1
rlabel polysilicon 401 -877 401 -877 0 3
rlabel polysilicon 411 -871 411 -871 0 2
rlabel polysilicon 408 -877 408 -877 0 3
rlabel polysilicon 411 -877 411 -877 0 4
rlabel polysilicon 415 -871 415 -871 0 1
rlabel polysilicon 415 -877 415 -877 0 3
rlabel polysilicon 422 -871 422 -871 0 1
rlabel polysilicon 422 -877 422 -877 0 3
rlabel polysilicon 429 -871 429 -871 0 1
rlabel polysilicon 429 -877 429 -877 0 3
rlabel polysilicon 436 -871 436 -871 0 1
rlabel polysilicon 436 -877 436 -877 0 3
rlabel polysilicon 443 -871 443 -871 0 1
rlabel polysilicon 443 -877 443 -877 0 3
rlabel polysilicon 450 -871 450 -871 0 1
rlabel polysilicon 450 -877 450 -877 0 3
rlabel polysilicon 457 -871 457 -871 0 1
rlabel polysilicon 457 -877 457 -877 0 3
rlabel polysilicon 464 -871 464 -871 0 1
rlabel polysilicon 464 -877 464 -877 0 3
rlabel polysilicon 471 -871 471 -871 0 1
rlabel polysilicon 471 -877 471 -877 0 3
rlabel polysilicon 478 -871 478 -871 0 1
rlabel polysilicon 478 -877 478 -877 0 3
rlabel polysilicon 485 -871 485 -871 0 1
rlabel polysilicon 485 -877 485 -877 0 3
rlabel polysilicon 492 -871 492 -871 0 1
rlabel polysilicon 492 -877 492 -877 0 3
rlabel polysilicon 499 -871 499 -871 0 1
rlabel polysilicon 499 -877 499 -877 0 3
rlabel polysilicon 502 -877 502 -877 0 4
rlabel polysilicon 506 -871 506 -871 0 1
rlabel polysilicon 509 -871 509 -871 0 2
rlabel polysilicon 506 -877 506 -877 0 3
rlabel polysilicon 509 -877 509 -877 0 4
rlabel polysilicon 513 -871 513 -871 0 1
rlabel polysilicon 513 -877 513 -877 0 3
rlabel polysilicon 520 -871 520 -871 0 1
rlabel polysilicon 523 -871 523 -871 0 2
rlabel polysilicon 520 -877 520 -877 0 3
rlabel polysilicon 523 -877 523 -877 0 4
rlabel polysilicon 527 -871 527 -871 0 1
rlabel polysilicon 530 -871 530 -871 0 2
rlabel polysilicon 527 -877 527 -877 0 3
rlabel polysilicon 530 -877 530 -877 0 4
rlabel polysilicon 534 -871 534 -871 0 1
rlabel polysilicon 534 -877 534 -877 0 3
rlabel polysilicon 537 -877 537 -877 0 4
rlabel polysilicon 541 -871 541 -871 0 1
rlabel polysilicon 541 -877 541 -877 0 3
rlabel polysilicon 548 -871 548 -871 0 1
rlabel polysilicon 551 -871 551 -871 0 2
rlabel polysilicon 548 -877 548 -877 0 3
rlabel polysilicon 551 -877 551 -877 0 4
rlabel polysilicon 555 -871 555 -871 0 1
rlabel polysilicon 555 -877 555 -877 0 3
rlabel polysilicon 562 -871 562 -871 0 1
rlabel polysilicon 562 -877 562 -877 0 3
rlabel polysilicon 569 -871 569 -871 0 1
rlabel polysilicon 569 -877 569 -877 0 3
rlabel polysilicon 576 -871 576 -871 0 1
rlabel polysilicon 576 -877 576 -877 0 3
rlabel polysilicon 583 -871 583 -871 0 1
rlabel polysilicon 583 -877 583 -877 0 3
rlabel polysilicon 590 -871 590 -871 0 1
rlabel polysilicon 590 -877 590 -877 0 3
rlabel polysilicon 597 -871 597 -871 0 1
rlabel polysilicon 597 -877 597 -877 0 3
rlabel polysilicon 604 -871 604 -871 0 1
rlabel polysilicon 604 -877 604 -877 0 3
rlabel polysilicon 611 -871 611 -871 0 1
rlabel polysilicon 611 -877 611 -877 0 3
rlabel polysilicon 618 -871 618 -871 0 1
rlabel polysilicon 618 -877 618 -877 0 3
rlabel polysilicon 625 -877 625 -877 0 3
rlabel polysilicon 628 -877 628 -877 0 4
rlabel polysilicon 632 -871 632 -871 0 1
rlabel polysilicon 632 -877 632 -877 0 3
rlabel polysilicon 639 -871 639 -871 0 1
rlabel polysilicon 639 -877 639 -877 0 3
rlabel polysilicon 646 -871 646 -871 0 1
rlabel polysilicon 649 -871 649 -871 0 2
rlabel polysilicon 646 -877 646 -877 0 3
rlabel polysilicon 649 -877 649 -877 0 4
rlabel polysilicon 653 -871 653 -871 0 1
rlabel polysilicon 653 -877 653 -877 0 3
rlabel polysilicon 660 -871 660 -871 0 1
rlabel polysilicon 660 -877 660 -877 0 3
rlabel polysilicon 667 -871 667 -871 0 1
rlabel polysilicon 667 -877 667 -877 0 3
rlabel polysilicon 670 -877 670 -877 0 4
rlabel polysilicon 674 -871 674 -871 0 1
rlabel polysilicon 674 -877 674 -877 0 3
rlabel polysilicon 677 -877 677 -877 0 4
rlabel polysilicon 681 -871 681 -871 0 1
rlabel polysilicon 684 -871 684 -871 0 2
rlabel polysilicon 681 -877 681 -877 0 3
rlabel polysilicon 684 -877 684 -877 0 4
rlabel polysilicon 688 -871 688 -871 0 1
rlabel polysilicon 688 -877 688 -877 0 3
rlabel polysilicon 695 -871 695 -871 0 1
rlabel polysilicon 695 -877 695 -877 0 3
rlabel polysilicon 702 -871 702 -871 0 1
rlabel polysilicon 702 -877 702 -877 0 3
rlabel polysilicon 709 -871 709 -871 0 1
rlabel polysilicon 709 -877 709 -877 0 3
rlabel polysilicon 716 -871 716 -871 0 1
rlabel polysilicon 716 -877 716 -877 0 3
rlabel polysilicon 723 -871 723 -871 0 1
rlabel polysilicon 723 -877 723 -877 0 3
rlabel polysilicon 730 -871 730 -871 0 1
rlabel polysilicon 730 -877 730 -877 0 3
rlabel polysilicon 737 -871 737 -871 0 1
rlabel polysilicon 737 -877 737 -877 0 3
rlabel polysilicon 744 -871 744 -871 0 1
rlabel polysilicon 744 -877 744 -877 0 3
rlabel polysilicon 751 -871 751 -871 0 1
rlabel polysilicon 751 -877 751 -877 0 3
rlabel polysilicon 758 -871 758 -871 0 1
rlabel polysilicon 758 -877 758 -877 0 3
rlabel polysilicon 765 -871 765 -871 0 1
rlabel polysilicon 765 -877 765 -877 0 3
rlabel polysilicon 772 -871 772 -871 0 1
rlabel polysilicon 772 -877 772 -877 0 3
rlabel polysilicon 779 -871 779 -871 0 1
rlabel polysilicon 782 -871 782 -871 0 2
rlabel polysilicon 782 -877 782 -877 0 4
rlabel polysilicon 786 -871 786 -871 0 1
rlabel polysilicon 786 -877 786 -877 0 3
rlabel polysilicon 793 -871 793 -871 0 1
rlabel polysilicon 793 -877 793 -877 0 3
rlabel polysilicon 800 -871 800 -871 0 1
rlabel polysilicon 800 -877 800 -877 0 3
rlabel polysilicon 807 -871 807 -871 0 1
rlabel polysilicon 807 -877 807 -877 0 3
rlabel polysilicon 814 -871 814 -871 0 1
rlabel polysilicon 814 -877 814 -877 0 3
rlabel polysilicon 821 -871 821 -871 0 1
rlabel polysilicon 821 -877 821 -877 0 3
rlabel polysilicon 828 -871 828 -871 0 1
rlabel polysilicon 831 -871 831 -871 0 2
rlabel polysilicon 828 -877 828 -877 0 3
rlabel polysilicon 831 -877 831 -877 0 4
rlabel polysilicon 835 -871 835 -871 0 1
rlabel polysilicon 838 -871 838 -871 0 2
rlabel polysilicon 835 -877 835 -877 0 3
rlabel polysilicon 838 -877 838 -877 0 4
rlabel polysilicon 842 -871 842 -871 0 1
rlabel polysilicon 842 -877 842 -877 0 3
rlabel polysilicon 849 -871 849 -871 0 1
rlabel polysilicon 849 -877 849 -877 0 3
rlabel polysilicon 856 -871 856 -871 0 1
rlabel polysilicon 856 -877 856 -877 0 3
rlabel polysilicon 863 -871 863 -871 0 1
rlabel polysilicon 863 -877 863 -877 0 3
rlabel polysilicon 870 -871 870 -871 0 1
rlabel polysilicon 873 -871 873 -871 0 2
rlabel polysilicon 870 -877 870 -877 0 3
rlabel polysilicon 873 -877 873 -877 0 4
rlabel polysilicon 877 -871 877 -871 0 1
rlabel polysilicon 880 -871 880 -871 0 2
rlabel polysilicon 877 -877 877 -877 0 3
rlabel polysilicon 880 -877 880 -877 0 4
rlabel polysilicon 884 -871 884 -871 0 1
rlabel polysilicon 884 -877 884 -877 0 3
rlabel polysilicon 891 -871 891 -871 0 1
rlabel polysilicon 891 -877 891 -877 0 3
rlabel polysilicon 898 -871 898 -871 0 1
rlabel polysilicon 898 -877 898 -877 0 3
rlabel polysilicon 905 -871 905 -871 0 1
rlabel polysilicon 905 -877 905 -877 0 3
rlabel polysilicon 912 -871 912 -871 0 1
rlabel polysilicon 912 -877 912 -877 0 3
rlabel polysilicon 919 -871 919 -871 0 1
rlabel polysilicon 922 -871 922 -871 0 2
rlabel polysilicon 919 -877 919 -877 0 3
rlabel polysilicon 922 -877 922 -877 0 4
rlabel polysilicon 926 -871 926 -871 0 1
rlabel polysilicon 926 -877 926 -877 0 3
rlabel polysilicon 929 -877 929 -877 0 4
rlabel polysilicon 933 -871 933 -871 0 1
rlabel polysilicon 933 -877 933 -877 0 3
rlabel polysilicon 940 -871 940 -871 0 1
rlabel polysilicon 940 -877 940 -877 0 3
rlabel polysilicon 947 -871 947 -871 0 1
rlabel polysilicon 947 -877 947 -877 0 3
rlabel polysilicon 954 -871 954 -871 0 1
rlabel polysilicon 954 -877 954 -877 0 3
rlabel polysilicon 961 -871 961 -871 0 1
rlabel polysilicon 964 -871 964 -871 0 2
rlabel polysilicon 964 -877 964 -877 0 4
rlabel polysilicon 968 -871 968 -871 0 1
rlabel polysilicon 968 -877 968 -877 0 3
rlabel polysilicon 975 -871 975 -871 0 1
rlabel polysilicon 975 -877 975 -877 0 3
rlabel polysilicon 982 -871 982 -871 0 1
rlabel polysilicon 982 -877 982 -877 0 3
rlabel polysilicon 989 -871 989 -871 0 1
rlabel polysilicon 989 -877 989 -877 0 3
rlabel polysilicon 996 -871 996 -871 0 1
rlabel polysilicon 996 -877 996 -877 0 3
rlabel polysilicon 1003 -871 1003 -871 0 1
rlabel polysilicon 1003 -877 1003 -877 0 3
rlabel polysilicon 1010 -871 1010 -871 0 1
rlabel polysilicon 1010 -877 1010 -877 0 3
rlabel polysilicon 1017 -871 1017 -871 0 1
rlabel polysilicon 1017 -877 1017 -877 0 3
rlabel polysilicon 1024 -871 1024 -871 0 1
rlabel polysilicon 1024 -877 1024 -877 0 3
rlabel polysilicon 1031 -871 1031 -871 0 1
rlabel polysilicon 1031 -877 1031 -877 0 3
rlabel polysilicon 1038 -871 1038 -871 0 1
rlabel polysilicon 1038 -877 1038 -877 0 3
rlabel polysilicon 1045 -871 1045 -871 0 1
rlabel polysilicon 1045 -877 1045 -877 0 3
rlabel polysilicon 1052 -871 1052 -871 0 1
rlabel polysilicon 1052 -877 1052 -877 0 3
rlabel polysilicon 1059 -871 1059 -871 0 1
rlabel polysilicon 1059 -877 1059 -877 0 3
rlabel polysilicon 1066 -871 1066 -871 0 1
rlabel polysilicon 1066 -877 1066 -877 0 3
rlabel polysilicon 1069 -877 1069 -877 0 4
rlabel polysilicon 1073 -871 1073 -871 0 1
rlabel polysilicon 1073 -877 1073 -877 0 3
rlabel polysilicon 1080 -871 1080 -871 0 1
rlabel polysilicon 1080 -877 1080 -877 0 3
rlabel polysilicon 1087 -871 1087 -871 0 1
rlabel polysilicon 1087 -877 1087 -877 0 3
rlabel polysilicon 1094 -871 1094 -871 0 1
rlabel polysilicon 1094 -877 1094 -877 0 3
rlabel polysilicon 1101 -871 1101 -871 0 1
rlabel polysilicon 1101 -877 1101 -877 0 3
rlabel polysilicon 1108 -871 1108 -871 0 1
rlabel polysilicon 1108 -877 1108 -877 0 3
rlabel polysilicon 1115 -871 1115 -871 0 1
rlabel polysilicon 1115 -877 1115 -877 0 3
rlabel polysilicon 1122 -871 1122 -871 0 1
rlabel polysilicon 1122 -877 1122 -877 0 3
rlabel polysilicon 1129 -871 1129 -871 0 1
rlabel polysilicon 1129 -877 1129 -877 0 3
rlabel polysilicon 1136 -871 1136 -871 0 1
rlabel polysilicon 1136 -877 1136 -877 0 3
rlabel polysilicon 1143 -871 1143 -871 0 1
rlabel polysilicon 1143 -877 1143 -877 0 3
rlabel polysilicon 1150 -871 1150 -871 0 1
rlabel polysilicon 1150 -877 1150 -877 0 3
rlabel polysilicon 1157 -871 1157 -871 0 1
rlabel polysilicon 1157 -877 1157 -877 0 3
rlabel polysilicon 1164 -871 1164 -871 0 1
rlabel polysilicon 1164 -877 1164 -877 0 3
rlabel polysilicon 1171 -871 1171 -871 0 1
rlabel polysilicon 1171 -877 1171 -877 0 3
rlabel polysilicon 1178 -871 1178 -871 0 1
rlabel polysilicon 1178 -877 1178 -877 0 3
rlabel polysilicon 1185 -871 1185 -871 0 1
rlabel polysilicon 1185 -877 1185 -877 0 3
rlabel polysilicon 1192 -871 1192 -871 0 1
rlabel polysilicon 1192 -877 1192 -877 0 3
rlabel polysilicon 1199 -871 1199 -871 0 1
rlabel polysilicon 1199 -877 1199 -877 0 3
rlabel polysilicon 1206 -871 1206 -871 0 1
rlabel polysilicon 1206 -877 1206 -877 0 3
rlabel polysilicon 1213 -871 1213 -871 0 1
rlabel polysilicon 1213 -877 1213 -877 0 3
rlabel polysilicon 1220 -871 1220 -871 0 1
rlabel polysilicon 1220 -877 1220 -877 0 3
rlabel polysilicon 1227 -871 1227 -871 0 1
rlabel polysilicon 1227 -877 1227 -877 0 3
rlabel polysilicon 1234 -871 1234 -871 0 1
rlabel polysilicon 1234 -877 1234 -877 0 3
rlabel polysilicon 1241 -871 1241 -871 0 1
rlabel polysilicon 1241 -877 1241 -877 0 3
rlabel polysilicon 1248 -871 1248 -871 0 1
rlabel polysilicon 1248 -877 1248 -877 0 3
rlabel polysilicon 1255 -871 1255 -871 0 1
rlabel polysilicon 1255 -877 1255 -877 0 3
rlabel polysilicon 1262 -871 1262 -871 0 1
rlabel polysilicon 1262 -877 1262 -877 0 3
rlabel polysilicon 1269 -871 1269 -871 0 1
rlabel polysilicon 1269 -877 1269 -877 0 3
rlabel polysilicon 1276 -871 1276 -871 0 1
rlabel polysilicon 1276 -877 1276 -877 0 3
rlabel polysilicon 1283 -871 1283 -871 0 1
rlabel polysilicon 1283 -877 1283 -877 0 3
rlabel polysilicon 1290 -871 1290 -871 0 1
rlabel polysilicon 1290 -877 1290 -877 0 3
rlabel polysilicon 1297 -871 1297 -871 0 1
rlabel polysilicon 1297 -877 1297 -877 0 3
rlabel polysilicon 1304 -871 1304 -871 0 1
rlabel polysilicon 1304 -877 1304 -877 0 3
rlabel polysilicon 1311 -871 1311 -871 0 1
rlabel polysilicon 1311 -877 1311 -877 0 3
rlabel polysilicon 1318 -871 1318 -871 0 1
rlabel polysilicon 1318 -877 1318 -877 0 3
rlabel polysilicon 1325 -871 1325 -871 0 1
rlabel polysilicon 1325 -877 1325 -877 0 3
rlabel polysilicon 1332 -871 1332 -871 0 1
rlabel polysilicon 1332 -877 1332 -877 0 3
rlabel polysilicon 1339 -871 1339 -871 0 1
rlabel polysilicon 1339 -877 1339 -877 0 3
rlabel polysilicon 1346 -871 1346 -871 0 1
rlabel polysilicon 1346 -877 1346 -877 0 3
rlabel polysilicon 1353 -871 1353 -871 0 1
rlabel polysilicon 1353 -877 1353 -877 0 3
rlabel polysilicon 1360 -871 1360 -871 0 1
rlabel polysilicon 1360 -877 1360 -877 0 3
rlabel polysilicon 1367 -871 1367 -871 0 1
rlabel polysilicon 1367 -877 1367 -877 0 3
rlabel polysilicon 1374 -871 1374 -871 0 1
rlabel polysilicon 1374 -877 1374 -877 0 3
rlabel polysilicon 1381 -871 1381 -871 0 1
rlabel polysilicon 1381 -877 1381 -877 0 3
rlabel polysilicon 1388 -871 1388 -871 0 1
rlabel polysilicon 1388 -877 1388 -877 0 3
rlabel polysilicon 1395 -871 1395 -871 0 1
rlabel polysilicon 1395 -877 1395 -877 0 3
rlabel polysilicon 1402 -871 1402 -871 0 1
rlabel polysilicon 1402 -877 1402 -877 0 3
rlabel polysilicon 1409 -871 1409 -871 0 1
rlabel polysilicon 1409 -877 1409 -877 0 3
rlabel polysilicon 1416 -871 1416 -871 0 1
rlabel polysilicon 1416 -877 1416 -877 0 3
rlabel polysilicon 1423 -871 1423 -871 0 1
rlabel polysilicon 1423 -877 1423 -877 0 3
rlabel polysilicon 1430 -871 1430 -871 0 1
rlabel polysilicon 1430 -877 1430 -877 0 3
rlabel polysilicon 1437 -871 1437 -871 0 1
rlabel polysilicon 1437 -877 1437 -877 0 3
rlabel polysilicon 1444 -871 1444 -871 0 1
rlabel polysilicon 1444 -877 1444 -877 0 3
rlabel polysilicon 1451 -871 1451 -871 0 1
rlabel polysilicon 1451 -877 1451 -877 0 3
rlabel polysilicon 1458 -871 1458 -871 0 1
rlabel polysilicon 1458 -877 1458 -877 0 3
rlabel polysilicon 1465 -871 1465 -871 0 1
rlabel polysilicon 1465 -877 1465 -877 0 3
rlabel polysilicon 1472 -871 1472 -871 0 1
rlabel polysilicon 1472 -877 1472 -877 0 3
rlabel polysilicon 1479 -871 1479 -871 0 1
rlabel polysilicon 1479 -877 1479 -877 0 3
rlabel polysilicon 1486 -871 1486 -871 0 1
rlabel polysilicon 1486 -877 1486 -877 0 3
rlabel polysilicon 1493 -871 1493 -871 0 1
rlabel polysilicon 1493 -877 1493 -877 0 3
rlabel polysilicon 1500 -871 1500 -871 0 1
rlabel polysilicon 1500 -877 1500 -877 0 3
rlabel polysilicon 1507 -871 1507 -871 0 1
rlabel polysilicon 1507 -877 1507 -877 0 3
rlabel polysilicon 1514 -871 1514 -871 0 1
rlabel polysilicon 1514 -877 1514 -877 0 3
rlabel polysilicon 1521 -871 1521 -871 0 1
rlabel polysilicon 1521 -877 1521 -877 0 3
rlabel polysilicon 1528 -871 1528 -871 0 1
rlabel polysilicon 1528 -877 1528 -877 0 3
rlabel polysilicon 1535 -871 1535 -871 0 1
rlabel polysilicon 1535 -877 1535 -877 0 3
rlabel polysilicon 1542 -871 1542 -871 0 1
rlabel polysilicon 1542 -877 1542 -877 0 3
rlabel polysilicon 1549 -871 1549 -871 0 1
rlabel polysilicon 1549 -877 1549 -877 0 3
rlabel polysilicon 1556 -871 1556 -871 0 1
rlabel polysilicon 1559 -871 1559 -871 0 2
rlabel polysilicon 1556 -877 1556 -877 0 3
rlabel polysilicon 1563 -877 1563 -877 0 3
rlabel polysilicon 1570 -871 1570 -871 0 1
rlabel polysilicon 1570 -877 1570 -877 0 3
rlabel polysilicon 1577 -871 1577 -871 0 1
rlabel polysilicon 1577 -877 1577 -877 0 3
rlabel polysilicon 1584 -871 1584 -871 0 1
rlabel polysilicon 1584 -877 1584 -877 0 3
rlabel polysilicon 1724 -871 1724 -871 0 1
rlabel polysilicon 1724 -877 1724 -877 0 3
rlabel polysilicon 30 -998 30 -998 0 1
rlabel polysilicon 30 -1004 30 -1004 0 3
rlabel polysilicon 37 -998 37 -998 0 1
rlabel polysilicon 37 -1004 37 -1004 0 3
rlabel polysilicon 44 -998 44 -998 0 1
rlabel polysilicon 44 -1004 44 -1004 0 3
rlabel polysilicon 51 -998 51 -998 0 1
rlabel polysilicon 51 -1004 51 -1004 0 3
rlabel polysilicon 58 -998 58 -998 0 1
rlabel polysilicon 58 -1004 58 -1004 0 3
rlabel polysilicon 65 -998 65 -998 0 1
rlabel polysilicon 72 -998 72 -998 0 1
rlabel polysilicon 72 -1004 72 -1004 0 3
rlabel polysilicon 79 -998 79 -998 0 1
rlabel polysilicon 82 -998 82 -998 0 2
rlabel polysilicon 79 -1004 79 -1004 0 3
rlabel polysilicon 82 -1004 82 -1004 0 4
rlabel polysilicon 86 -998 86 -998 0 1
rlabel polysilicon 86 -1004 86 -1004 0 3
rlabel polysilicon 93 -998 93 -998 0 1
rlabel polysilicon 93 -1004 93 -1004 0 3
rlabel polysilicon 100 -998 100 -998 0 1
rlabel polysilicon 100 -1004 100 -1004 0 3
rlabel polysilicon 107 -998 107 -998 0 1
rlabel polysilicon 107 -1004 107 -1004 0 3
rlabel polysilicon 114 -998 114 -998 0 1
rlabel polysilicon 114 -1004 114 -1004 0 3
rlabel polysilicon 121 -998 121 -998 0 1
rlabel polysilicon 121 -1004 121 -1004 0 3
rlabel polysilicon 128 -998 128 -998 0 1
rlabel polysilicon 128 -1004 128 -1004 0 3
rlabel polysilicon 131 -1004 131 -1004 0 4
rlabel polysilicon 135 -998 135 -998 0 1
rlabel polysilicon 138 -998 138 -998 0 2
rlabel polysilicon 138 -1004 138 -1004 0 4
rlabel polysilicon 142 -998 142 -998 0 1
rlabel polysilicon 142 -1004 142 -1004 0 3
rlabel polysilicon 149 -998 149 -998 0 1
rlabel polysilicon 152 -998 152 -998 0 2
rlabel polysilicon 156 -998 156 -998 0 1
rlabel polysilicon 156 -1004 156 -1004 0 3
rlabel polysilicon 163 -998 163 -998 0 1
rlabel polysilicon 163 -1004 163 -1004 0 3
rlabel polysilicon 170 -998 170 -998 0 1
rlabel polysilicon 170 -1004 170 -1004 0 3
rlabel polysilicon 177 -998 177 -998 0 1
rlabel polysilicon 177 -1004 177 -1004 0 3
rlabel polysilicon 184 -998 184 -998 0 1
rlabel polysilicon 184 -1004 184 -1004 0 3
rlabel polysilicon 191 -998 191 -998 0 1
rlabel polysilicon 191 -1004 191 -1004 0 3
rlabel polysilicon 198 -998 198 -998 0 1
rlabel polysilicon 198 -1004 198 -1004 0 3
rlabel polysilicon 205 -998 205 -998 0 1
rlabel polysilicon 205 -1004 205 -1004 0 3
rlabel polysilicon 212 -998 212 -998 0 1
rlabel polysilicon 212 -1004 212 -1004 0 3
rlabel polysilicon 219 -998 219 -998 0 1
rlabel polysilicon 219 -1004 219 -1004 0 3
rlabel polysilicon 226 -998 226 -998 0 1
rlabel polysilicon 226 -1004 226 -1004 0 3
rlabel polysilicon 233 -998 233 -998 0 1
rlabel polysilicon 233 -1004 233 -1004 0 3
rlabel polysilicon 240 -998 240 -998 0 1
rlabel polysilicon 250 -998 250 -998 0 2
rlabel polysilicon 250 -1004 250 -1004 0 4
rlabel polysilicon 254 -998 254 -998 0 1
rlabel polysilicon 254 -1004 254 -1004 0 3
rlabel polysilicon 261 -998 261 -998 0 1
rlabel polysilicon 261 -1004 261 -1004 0 3
rlabel polysilicon 268 -998 268 -998 0 1
rlabel polysilicon 268 -1004 268 -1004 0 3
rlabel polysilicon 275 -998 275 -998 0 1
rlabel polysilicon 275 -1004 275 -1004 0 3
rlabel polysilicon 282 -998 282 -998 0 1
rlabel polysilicon 282 -1004 282 -1004 0 3
rlabel polysilicon 289 -998 289 -998 0 1
rlabel polysilicon 289 -1004 289 -1004 0 3
rlabel polysilicon 296 -998 296 -998 0 1
rlabel polysilicon 296 -1004 296 -1004 0 3
rlabel polysilicon 303 -998 303 -998 0 1
rlabel polysilicon 303 -1004 303 -1004 0 3
rlabel polysilicon 310 -998 310 -998 0 1
rlabel polysilicon 310 -1004 310 -1004 0 3
rlabel polysilicon 317 -998 317 -998 0 1
rlabel polysilicon 317 -1004 317 -1004 0 3
rlabel polysilicon 324 -1004 324 -1004 0 3
rlabel polysilicon 331 -998 331 -998 0 1
rlabel polysilicon 331 -1004 331 -1004 0 3
rlabel polysilicon 338 -998 338 -998 0 1
rlabel polysilicon 338 -1004 338 -1004 0 3
rlabel polysilicon 345 -998 345 -998 0 1
rlabel polysilicon 345 -1004 345 -1004 0 3
rlabel polysilicon 352 -998 352 -998 0 1
rlabel polysilicon 352 -1004 352 -1004 0 3
rlabel polysilicon 359 -998 359 -998 0 1
rlabel polysilicon 359 -1004 359 -1004 0 3
rlabel polysilicon 366 -998 366 -998 0 1
rlabel polysilicon 366 -1004 366 -1004 0 3
rlabel polysilicon 373 -998 373 -998 0 1
rlabel polysilicon 373 -1004 373 -1004 0 3
rlabel polysilicon 380 -998 380 -998 0 1
rlabel polysilicon 380 -1004 380 -1004 0 3
rlabel polysilicon 387 -998 387 -998 0 1
rlabel polysilicon 387 -1004 387 -1004 0 3
rlabel polysilicon 394 -998 394 -998 0 1
rlabel polysilicon 394 -1004 394 -1004 0 3
rlabel polysilicon 401 -998 401 -998 0 1
rlabel polysilicon 401 -1004 401 -1004 0 3
rlabel polysilicon 408 -998 408 -998 0 1
rlabel polysilicon 408 -1004 408 -1004 0 3
rlabel polysilicon 415 -998 415 -998 0 1
rlabel polysilicon 415 -1004 415 -1004 0 3
rlabel polysilicon 422 -998 422 -998 0 1
rlabel polysilicon 425 -998 425 -998 0 2
rlabel polysilicon 422 -1004 422 -1004 0 3
rlabel polysilicon 425 -1004 425 -1004 0 4
rlabel polysilicon 429 -998 429 -998 0 1
rlabel polysilicon 429 -1004 429 -1004 0 3
rlabel polysilicon 436 -998 436 -998 0 1
rlabel polysilicon 436 -1004 436 -1004 0 3
rlabel polysilicon 443 -998 443 -998 0 1
rlabel polysilicon 446 -998 446 -998 0 2
rlabel polysilicon 443 -1004 443 -1004 0 3
rlabel polysilicon 446 -1004 446 -1004 0 4
rlabel polysilicon 450 -998 450 -998 0 1
rlabel polysilicon 450 -1004 450 -1004 0 3
rlabel polysilicon 457 -998 457 -998 0 1
rlabel polysilicon 457 -1004 457 -1004 0 3
rlabel polysilicon 464 -998 464 -998 0 1
rlabel polysilicon 464 -1004 464 -1004 0 3
rlabel polysilicon 471 -998 471 -998 0 1
rlabel polysilicon 471 -1004 471 -1004 0 3
rlabel polysilicon 478 -998 478 -998 0 1
rlabel polysilicon 478 -1004 478 -1004 0 3
rlabel polysilicon 485 -998 485 -998 0 1
rlabel polysilicon 485 -1004 485 -1004 0 3
rlabel polysilicon 492 -998 492 -998 0 1
rlabel polysilicon 492 -1004 492 -1004 0 3
rlabel polysilicon 499 -998 499 -998 0 1
rlabel polysilicon 502 -998 502 -998 0 2
rlabel polysilicon 499 -1004 499 -1004 0 3
rlabel polysilicon 502 -1004 502 -1004 0 4
rlabel polysilicon 506 -998 506 -998 0 1
rlabel polysilicon 509 -998 509 -998 0 2
rlabel polysilicon 506 -1004 506 -1004 0 3
rlabel polysilicon 509 -1004 509 -1004 0 4
rlabel polysilicon 513 -998 513 -998 0 1
rlabel polysilicon 513 -1004 513 -1004 0 3
rlabel polysilicon 520 -998 520 -998 0 1
rlabel polysilicon 520 -1004 520 -1004 0 3
rlabel polysilicon 527 -998 527 -998 0 1
rlabel polysilicon 527 -1004 527 -1004 0 3
rlabel polysilicon 534 -998 534 -998 0 1
rlabel polysilicon 534 -1004 534 -1004 0 3
rlabel polysilicon 541 -998 541 -998 0 1
rlabel polysilicon 541 -1004 541 -1004 0 3
rlabel polysilicon 548 -998 548 -998 0 1
rlabel polysilicon 548 -1004 548 -1004 0 3
rlabel polysilicon 555 -998 555 -998 0 1
rlabel polysilicon 555 -1004 555 -1004 0 3
rlabel polysilicon 562 -998 562 -998 0 1
rlabel polysilicon 562 -1004 562 -1004 0 3
rlabel polysilicon 569 -998 569 -998 0 1
rlabel polysilicon 569 -1004 569 -1004 0 3
rlabel polysilicon 576 -998 576 -998 0 1
rlabel polysilicon 576 -1004 576 -1004 0 3
rlabel polysilicon 583 -998 583 -998 0 1
rlabel polysilicon 586 -998 586 -998 0 2
rlabel polysilicon 583 -1004 583 -1004 0 3
rlabel polysilicon 586 -1004 586 -1004 0 4
rlabel polysilicon 590 -998 590 -998 0 1
rlabel polysilicon 590 -1004 590 -1004 0 3
rlabel polysilicon 597 -998 597 -998 0 1
rlabel polysilicon 597 -1004 597 -1004 0 3
rlabel polysilicon 604 -998 604 -998 0 1
rlabel polysilicon 604 -1004 604 -1004 0 3
rlabel polysilicon 611 -998 611 -998 0 1
rlabel polysilicon 611 -1004 611 -1004 0 3
rlabel polysilicon 618 -1004 618 -1004 0 3
rlabel polysilicon 621 -1004 621 -1004 0 4
rlabel polysilicon 625 -998 625 -998 0 1
rlabel polysilicon 625 -1004 625 -1004 0 3
rlabel polysilicon 632 -998 632 -998 0 1
rlabel polysilicon 632 -1004 632 -1004 0 3
rlabel polysilicon 639 -998 639 -998 0 1
rlabel polysilicon 642 -998 642 -998 0 2
rlabel polysilicon 639 -1004 639 -1004 0 3
rlabel polysilicon 646 -998 646 -998 0 1
rlabel polysilicon 649 -998 649 -998 0 2
rlabel polysilicon 646 -1004 646 -1004 0 3
rlabel polysilicon 649 -1004 649 -1004 0 4
rlabel polysilicon 653 -998 653 -998 0 1
rlabel polysilicon 656 -998 656 -998 0 2
rlabel polysilicon 653 -1004 653 -1004 0 3
rlabel polysilicon 656 -1004 656 -1004 0 4
rlabel polysilicon 660 -998 660 -998 0 1
rlabel polysilicon 660 -1004 660 -1004 0 3
rlabel polysilicon 667 -998 667 -998 0 1
rlabel polysilicon 667 -1004 667 -1004 0 3
rlabel polysilicon 674 -998 674 -998 0 1
rlabel polysilicon 674 -1004 674 -1004 0 3
rlabel polysilicon 681 -998 681 -998 0 1
rlabel polysilicon 684 -998 684 -998 0 2
rlabel polysilicon 681 -1004 681 -1004 0 3
rlabel polysilicon 684 -1004 684 -1004 0 4
rlabel polysilicon 688 -998 688 -998 0 1
rlabel polysilicon 691 -1004 691 -1004 0 4
rlabel polysilicon 695 -998 695 -998 0 1
rlabel polysilicon 698 -998 698 -998 0 2
rlabel polysilicon 695 -1004 695 -1004 0 3
rlabel polysilicon 698 -1004 698 -1004 0 4
rlabel polysilicon 702 -998 702 -998 0 1
rlabel polysilicon 702 -1004 702 -1004 0 3
rlabel polysilicon 709 -998 709 -998 0 1
rlabel polysilicon 709 -1004 709 -1004 0 3
rlabel polysilicon 716 -998 716 -998 0 1
rlabel polysilicon 716 -1004 716 -1004 0 3
rlabel polysilicon 723 -998 723 -998 0 1
rlabel polysilicon 723 -1004 723 -1004 0 3
rlabel polysilicon 730 -998 730 -998 0 1
rlabel polysilicon 733 -998 733 -998 0 2
rlabel polysilicon 730 -1004 730 -1004 0 3
rlabel polysilicon 733 -1004 733 -1004 0 4
rlabel polysilicon 737 -998 737 -998 0 1
rlabel polysilicon 737 -1004 737 -1004 0 3
rlabel polysilicon 744 -998 744 -998 0 1
rlabel polysilicon 744 -1004 744 -1004 0 3
rlabel polysilicon 751 -998 751 -998 0 1
rlabel polysilicon 751 -1004 751 -1004 0 3
rlabel polysilicon 758 -998 758 -998 0 1
rlabel polysilicon 758 -1004 758 -1004 0 3
rlabel polysilicon 765 -998 765 -998 0 1
rlabel polysilicon 768 -998 768 -998 0 2
rlabel polysilicon 765 -1004 765 -1004 0 3
rlabel polysilicon 768 -1004 768 -1004 0 4
rlabel polysilicon 772 -998 772 -998 0 1
rlabel polysilicon 775 -998 775 -998 0 2
rlabel polysilicon 775 -1004 775 -1004 0 4
rlabel polysilicon 779 -998 779 -998 0 1
rlabel polysilicon 779 -1004 779 -1004 0 3
rlabel polysilicon 786 -998 786 -998 0 1
rlabel polysilicon 786 -1004 786 -1004 0 3
rlabel polysilicon 793 -998 793 -998 0 1
rlabel polysilicon 793 -1004 793 -1004 0 3
rlabel polysilicon 800 -998 800 -998 0 1
rlabel polysilicon 800 -1004 800 -1004 0 3
rlabel polysilicon 807 -998 807 -998 0 1
rlabel polysilicon 807 -1004 807 -1004 0 3
rlabel polysilicon 814 -998 814 -998 0 1
rlabel polysilicon 814 -1004 814 -1004 0 3
rlabel polysilicon 821 -998 821 -998 0 1
rlabel polysilicon 821 -1004 821 -1004 0 3
rlabel polysilicon 828 -998 828 -998 0 1
rlabel polysilicon 828 -1004 828 -1004 0 3
rlabel polysilicon 835 -998 835 -998 0 1
rlabel polysilicon 835 -1004 835 -1004 0 3
rlabel polysilicon 842 -998 842 -998 0 1
rlabel polysilicon 845 -998 845 -998 0 2
rlabel polysilicon 842 -1004 842 -1004 0 3
rlabel polysilicon 845 -1004 845 -1004 0 4
rlabel polysilicon 849 -998 849 -998 0 1
rlabel polysilicon 849 -1004 849 -1004 0 3
rlabel polysilicon 856 -998 856 -998 0 1
rlabel polysilicon 856 -1004 856 -1004 0 3
rlabel polysilicon 863 -998 863 -998 0 1
rlabel polysilicon 863 -1004 863 -1004 0 3
rlabel polysilicon 870 -998 870 -998 0 1
rlabel polysilicon 870 -1004 870 -1004 0 3
rlabel polysilicon 877 -998 877 -998 0 1
rlabel polysilicon 877 -1004 877 -1004 0 3
rlabel polysilicon 884 -998 884 -998 0 1
rlabel polysilicon 887 -1004 887 -1004 0 4
rlabel polysilicon 891 -998 891 -998 0 1
rlabel polysilicon 891 -1004 891 -1004 0 3
rlabel polysilicon 898 -998 898 -998 0 1
rlabel polysilicon 901 -998 901 -998 0 2
rlabel polysilicon 898 -1004 898 -1004 0 3
rlabel polysilicon 901 -1004 901 -1004 0 4
rlabel polysilicon 905 -998 905 -998 0 1
rlabel polysilicon 905 -1004 905 -1004 0 3
rlabel polysilicon 912 -998 912 -998 0 1
rlabel polysilicon 912 -1004 912 -1004 0 3
rlabel polysilicon 919 -998 919 -998 0 1
rlabel polysilicon 919 -1004 919 -1004 0 3
rlabel polysilicon 926 -998 926 -998 0 1
rlabel polysilicon 929 -998 929 -998 0 2
rlabel polysilicon 926 -1004 926 -1004 0 3
rlabel polysilicon 933 -998 933 -998 0 1
rlabel polysilicon 933 -1004 933 -1004 0 3
rlabel polysilicon 940 -998 940 -998 0 1
rlabel polysilicon 940 -1004 940 -1004 0 3
rlabel polysilicon 947 -998 947 -998 0 1
rlabel polysilicon 947 -1004 947 -1004 0 3
rlabel polysilicon 954 -998 954 -998 0 1
rlabel polysilicon 954 -1004 954 -1004 0 3
rlabel polysilicon 961 -998 961 -998 0 1
rlabel polysilicon 964 -998 964 -998 0 2
rlabel polysilicon 961 -1004 961 -1004 0 3
rlabel polysilicon 968 -998 968 -998 0 1
rlabel polysilicon 968 -1004 968 -1004 0 3
rlabel polysilicon 975 -998 975 -998 0 1
rlabel polysilicon 978 -998 978 -998 0 2
rlabel polysilicon 978 -1004 978 -1004 0 4
rlabel polysilicon 982 -998 982 -998 0 1
rlabel polysilicon 985 -998 985 -998 0 2
rlabel polysilicon 982 -1004 982 -1004 0 3
rlabel polysilicon 985 -1004 985 -1004 0 4
rlabel polysilicon 992 -998 992 -998 0 2
rlabel polysilicon 989 -1004 989 -1004 0 3
rlabel polysilicon 992 -1004 992 -1004 0 4
rlabel polysilicon 996 -998 996 -998 0 1
rlabel polysilicon 999 -998 999 -998 0 2
rlabel polysilicon 996 -1004 996 -1004 0 3
rlabel polysilicon 999 -1004 999 -1004 0 4
rlabel polysilicon 1003 -998 1003 -998 0 1
rlabel polysilicon 1003 -1004 1003 -1004 0 3
rlabel polysilicon 1010 -998 1010 -998 0 1
rlabel polysilicon 1010 -1004 1010 -1004 0 3
rlabel polysilicon 1013 -1004 1013 -1004 0 4
rlabel polysilicon 1017 -998 1017 -998 0 1
rlabel polysilicon 1017 -1004 1017 -1004 0 3
rlabel polysilicon 1024 -998 1024 -998 0 1
rlabel polysilicon 1024 -1004 1024 -1004 0 3
rlabel polysilicon 1027 -1004 1027 -1004 0 4
rlabel polysilicon 1031 -998 1031 -998 0 1
rlabel polysilicon 1031 -1004 1031 -1004 0 3
rlabel polysilicon 1038 -998 1038 -998 0 1
rlabel polysilicon 1038 -1004 1038 -1004 0 3
rlabel polysilicon 1045 -998 1045 -998 0 1
rlabel polysilicon 1045 -1004 1045 -1004 0 3
rlabel polysilicon 1052 -998 1052 -998 0 1
rlabel polysilicon 1052 -1004 1052 -1004 0 3
rlabel polysilicon 1059 -998 1059 -998 0 1
rlabel polysilicon 1059 -1004 1059 -1004 0 3
rlabel polysilicon 1066 -998 1066 -998 0 1
rlabel polysilicon 1066 -1004 1066 -1004 0 3
rlabel polysilicon 1073 -998 1073 -998 0 1
rlabel polysilicon 1073 -1004 1073 -1004 0 3
rlabel polysilicon 1080 -998 1080 -998 0 1
rlabel polysilicon 1080 -1004 1080 -1004 0 3
rlabel polysilicon 1087 -998 1087 -998 0 1
rlabel polysilicon 1087 -1004 1087 -1004 0 3
rlabel polysilicon 1094 -998 1094 -998 0 1
rlabel polysilicon 1094 -1004 1094 -1004 0 3
rlabel polysilicon 1101 -998 1101 -998 0 1
rlabel polysilicon 1101 -1004 1101 -1004 0 3
rlabel polysilicon 1111 -998 1111 -998 0 2
rlabel polysilicon 1108 -1004 1108 -1004 0 3
rlabel polysilicon 1111 -1004 1111 -1004 0 4
rlabel polysilicon 1115 -998 1115 -998 0 1
rlabel polysilicon 1115 -1004 1115 -1004 0 3
rlabel polysilicon 1122 -998 1122 -998 0 1
rlabel polysilicon 1122 -1004 1122 -1004 0 3
rlabel polysilicon 1129 -998 1129 -998 0 1
rlabel polysilicon 1129 -1004 1129 -1004 0 3
rlabel polysilicon 1132 -1004 1132 -1004 0 4
rlabel polysilicon 1136 -998 1136 -998 0 1
rlabel polysilicon 1136 -1004 1136 -1004 0 3
rlabel polysilicon 1143 -998 1143 -998 0 1
rlabel polysilicon 1143 -1004 1143 -1004 0 3
rlabel polysilicon 1150 -998 1150 -998 0 1
rlabel polysilicon 1150 -1004 1150 -1004 0 3
rlabel polysilicon 1157 -998 1157 -998 0 1
rlabel polysilicon 1157 -1004 1157 -1004 0 3
rlabel polysilicon 1164 -998 1164 -998 0 1
rlabel polysilicon 1164 -1004 1164 -1004 0 3
rlabel polysilicon 1171 -998 1171 -998 0 1
rlabel polysilicon 1171 -1004 1171 -1004 0 3
rlabel polysilicon 1178 -998 1178 -998 0 1
rlabel polysilicon 1178 -1004 1178 -1004 0 3
rlabel polysilicon 1185 -998 1185 -998 0 1
rlabel polysilicon 1185 -1004 1185 -1004 0 3
rlabel polysilicon 1192 -998 1192 -998 0 1
rlabel polysilicon 1192 -1004 1192 -1004 0 3
rlabel polysilicon 1199 -998 1199 -998 0 1
rlabel polysilicon 1199 -1004 1199 -1004 0 3
rlabel polysilicon 1206 -998 1206 -998 0 1
rlabel polysilicon 1206 -1004 1206 -1004 0 3
rlabel polysilicon 1213 -998 1213 -998 0 1
rlabel polysilicon 1213 -1004 1213 -1004 0 3
rlabel polysilicon 1220 -998 1220 -998 0 1
rlabel polysilicon 1220 -1004 1220 -1004 0 3
rlabel polysilicon 1227 -998 1227 -998 0 1
rlabel polysilicon 1227 -1004 1227 -1004 0 3
rlabel polysilicon 1234 -998 1234 -998 0 1
rlabel polysilicon 1234 -1004 1234 -1004 0 3
rlabel polysilicon 1241 -998 1241 -998 0 1
rlabel polysilicon 1241 -1004 1241 -1004 0 3
rlabel polysilicon 1248 -998 1248 -998 0 1
rlabel polysilicon 1248 -1004 1248 -1004 0 3
rlabel polysilicon 1255 -998 1255 -998 0 1
rlabel polysilicon 1255 -1004 1255 -1004 0 3
rlabel polysilicon 1262 -998 1262 -998 0 1
rlabel polysilicon 1262 -1004 1262 -1004 0 3
rlabel polysilicon 1269 -998 1269 -998 0 1
rlabel polysilicon 1269 -1004 1269 -1004 0 3
rlabel polysilicon 1276 -998 1276 -998 0 1
rlabel polysilicon 1276 -1004 1276 -1004 0 3
rlabel polysilicon 1283 -998 1283 -998 0 1
rlabel polysilicon 1283 -1004 1283 -1004 0 3
rlabel polysilicon 1290 -998 1290 -998 0 1
rlabel polysilicon 1290 -1004 1290 -1004 0 3
rlabel polysilicon 1297 -998 1297 -998 0 1
rlabel polysilicon 1297 -1004 1297 -1004 0 3
rlabel polysilicon 1304 -998 1304 -998 0 1
rlabel polysilicon 1304 -1004 1304 -1004 0 3
rlabel polysilicon 1311 -998 1311 -998 0 1
rlabel polysilicon 1311 -1004 1311 -1004 0 3
rlabel polysilicon 1318 -998 1318 -998 0 1
rlabel polysilicon 1318 -1004 1318 -1004 0 3
rlabel polysilicon 1325 -998 1325 -998 0 1
rlabel polysilicon 1325 -1004 1325 -1004 0 3
rlabel polysilicon 1332 -998 1332 -998 0 1
rlabel polysilicon 1332 -1004 1332 -1004 0 3
rlabel polysilicon 1339 -998 1339 -998 0 1
rlabel polysilicon 1339 -1004 1339 -1004 0 3
rlabel polysilicon 1346 -998 1346 -998 0 1
rlabel polysilicon 1346 -1004 1346 -1004 0 3
rlabel polysilicon 1353 -998 1353 -998 0 1
rlabel polysilicon 1353 -1004 1353 -1004 0 3
rlabel polysilicon 1360 -998 1360 -998 0 1
rlabel polysilicon 1360 -1004 1360 -1004 0 3
rlabel polysilicon 1367 -998 1367 -998 0 1
rlabel polysilicon 1367 -1004 1367 -1004 0 3
rlabel polysilicon 1374 -998 1374 -998 0 1
rlabel polysilicon 1374 -1004 1374 -1004 0 3
rlabel polysilicon 1381 -998 1381 -998 0 1
rlabel polysilicon 1381 -1004 1381 -1004 0 3
rlabel polysilicon 1388 -998 1388 -998 0 1
rlabel polysilicon 1388 -1004 1388 -1004 0 3
rlabel polysilicon 1395 -998 1395 -998 0 1
rlabel polysilicon 1395 -1004 1395 -1004 0 3
rlabel polysilicon 1402 -998 1402 -998 0 1
rlabel polysilicon 1402 -1004 1402 -1004 0 3
rlabel polysilicon 1409 -998 1409 -998 0 1
rlabel polysilicon 1409 -1004 1409 -1004 0 3
rlabel polysilicon 1416 -998 1416 -998 0 1
rlabel polysilicon 1416 -1004 1416 -1004 0 3
rlabel polysilicon 1423 -998 1423 -998 0 1
rlabel polysilicon 1423 -1004 1423 -1004 0 3
rlabel polysilicon 1430 -998 1430 -998 0 1
rlabel polysilicon 1430 -1004 1430 -1004 0 3
rlabel polysilicon 1437 -998 1437 -998 0 1
rlabel polysilicon 1437 -1004 1437 -1004 0 3
rlabel polysilicon 1444 -998 1444 -998 0 1
rlabel polysilicon 1444 -1004 1444 -1004 0 3
rlabel polysilicon 1451 -998 1451 -998 0 1
rlabel polysilicon 1451 -1004 1451 -1004 0 3
rlabel polysilicon 1458 -998 1458 -998 0 1
rlabel polysilicon 1458 -1004 1458 -1004 0 3
rlabel polysilicon 1465 -998 1465 -998 0 1
rlabel polysilicon 1465 -1004 1465 -1004 0 3
rlabel polysilicon 1472 -998 1472 -998 0 1
rlabel polysilicon 1472 -1004 1472 -1004 0 3
rlabel polysilicon 1479 -998 1479 -998 0 1
rlabel polysilicon 1479 -1004 1479 -1004 0 3
rlabel polysilicon 1486 -998 1486 -998 0 1
rlabel polysilicon 1486 -1004 1486 -1004 0 3
rlabel polysilicon 1493 -998 1493 -998 0 1
rlabel polysilicon 1493 -1004 1493 -1004 0 3
rlabel polysilicon 1500 -998 1500 -998 0 1
rlabel polysilicon 1500 -1004 1500 -1004 0 3
rlabel polysilicon 1507 -998 1507 -998 0 1
rlabel polysilicon 1507 -1004 1507 -1004 0 3
rlabel polysilicon 1514 -998 1514 -998 0 1
rlabel polysilicon 1514 -1004 1514 -1004 0 3
rlabel polysilicon 1521 -998 1521 -998 0 1
rlabel polysilicon 1521 -1004 1521 -1004 0 3
rlabel polysilicon 1528 -998 1528 -998 0 1
rlabel polysilicon 1528 -1004 1528 -1004 0 3
rlabel polysilicon 1535 -998 1535 -998 0 1
rlabel polysilicon 1535 -1004 1535 -1004 0 3
rlabel polysilicon 1542 -998 1542 -998 0 1
rlabel polysilicon 1542 -1004 1542 -1004 0 3
rlabel polysilicon 1549 -998 1549 -998 0 1
rlabel polysilicon 1549 -1004 1549 -1004 0 3
rlabel polysilicon 1552 -1004 1552 -1004 0 4
rlabel polysilicon 1556 -998 1556 -998 0 1
rlabel polysilicon 1556 -1004 1556 -1004 0 3
rlabel polysilicon 1563 -998 1563 -998 0 1
rlabel polysilicon 1566 -998 1566 -998 0 2
rlabel polysilicon 1563 -1004 1563 -1004 0 3
rlabel polysilicon 1566 -1004 1566 -1004 0 4
rlabel polysilicon 1570 -998 1570 -998 0 1
rlabel polysilicon 1573 -998 1573 -998 0 2
rlabel polysilicon 1570 -1004 1570 -1004 0 3
rlabel polysilicon 1577 -998 1577 -998 0 1
rlabel polysilicon 1577 -1004 1577 -1004 0 3
rlabel polysilicon 1584 -998 1584 -998 0 1
rlabel polysilicon 1584 -1004 1584 -1004 0 3
rlabel polysilicon 1591 -998 1591 -998 0 1
rlabel polysilicon 1591 -1004 1591 -1004 0 3
rlabel polysilicon 1598 -998 1598 -998 0 1
rlabel polysilicon 1598 -1004 1598 -1004 0 3
rlabel polysilicon 1605 -998 1605 -998 0 1
rlabel polysilicon 1605 -1004 1605 -1004 0 3
rlabel polysilicon 1612 -998 1612 -998 0 1
rlabel polysilicon 1612 -1004 1612 -1004 0 3
rlabel polysilicon 1619 -998 1619 -998 0 1
rlabel polysilicon 1619 -1004 1619 -1004 0 3
rlabel polysilicon 1626 -998 1626 -998 0 1
rlabel polysilicon 1626 -1004 1626 -1004 0 3
rlabel polysilicon 1633 -998 1633 -998 0 1
rlabel polysilicon 1633 -1004 1633 -1004 0 3
rlabel polysilicon 1738 -998 1738 -998 0 1
rlabel polysilicon 1738 -1004 1738 -1004 0 3
rlabel polysilicon 23 -1099 23 -1099 0 1
rlabel polysilicon 23 -1105 23 -1105 0 3
rlabel polysilicon 30 -1099 30 -1099 0 1
rlabel polysilicon 30 -1105 30 -1105 0 3
rlabel polysilicon 44 -1099 44 -1099 0 1
rlabel polysilicon 44 -1105 44 -1105 0 3
rlabel polysilicon 51 -1099 51 -1099 0 1
rlabel polysilicon 51 -1105 51 -1105 0 3
rlabel polysilicon 58 -1099 58 -1099 0 1
rlabel polysilicon 58 -1105 58 -1105 0 3
rlabel polysilicon 65 -1105 65 -1105 0 3
rlabel polysilicon 72 -1099 72 -1099 0 1
rlabel polysilicon 75 -1099 75 -1099 0 2
rlabel polysilicon 75 -1105 75 -1105 0 4
rlabel polysilicon 79 -1099 79 -1099 0 1
rlabel polysilicon 79 -1105 79 -1105 0 3
rlabel polysilicon 86 -1099 86 -1099 0 1
rlabel polysilicon 89 -1099 89 -1099 0 2
rlabel polysilicon 86 -1105 86 -1105 0 3
rlabel polysilicon 89 -1105 89 -1105 0 4
rlabel polysilicon 93 -1099 93 -1099 0 1
rlabel polysilicon 93 -1105 93 -1105 0 3
rlabel polysilicon 100 -1099 100 -1099 0 1
rlabel polysilicon 100 -1105 100 -1105 0 3
rlabel polysilicon 107 -1099 107 -1099 0 1
rlabel polysilicon 107 -1105 107 -1105 0 3
rlabel polysilicon 114 -1099 114 -1099 0 1
rlabel polysilicon 114 -1105 114 -1105 0 3
rlabel polysilicon 121 -1099 121 -1099 0 1
rlabel polysilicon 121 -1105 121 -1105 0 3
rlabel polysilicon 128 -1099 128 -1099 0 1
rlabel polysilicon 128 -1105 128 -1105 0 3
rlabel polysilicon 135 -1099 135 -1099 0 1
rlabel polysilicon 138 -1099 138 -1099 0 2
rlabel polysilicon 138 -1105 138 -1105 0 4
rlabel polysilicon 142 -1099 142 -1099 0 1
rlabel polysilicon 142 -1105 142 -1105 0 3
rlabel polysilicon 149 -1099 149 -1099 0 1
rlabel polysilicon 149 -1105 149 -1105 0 3
rlabel polysilicon 156 -1099 156 -1099 0 1
rlabel polysilicon 156 -1105 156 -1105 0 3
rlabel polysilicon 163 -1099 163 -1099 0 1
rlabel polysilicon 163 -1105 163 -1105 0 3
rlabel polysilicon 170 -1099 170 -1099 0 1
rlabel polysilicon 170 -1105 170 -1105 0 3
rlabel polysilicon 177 -1099 177 -1099 0 1
rlabel polysilicon 177 -1105 177 -1105 0 3
rlabel polysilicon 184 -1099 184 -1099 0 1
rlabel polysilicon 184 -1105 184 -1105 0 3
rlabel polysilicon 191 -1099 191 -1099 0 1
rlabel polysilicon 191 -1105 191 -1105 0 3
rlabel polysilicon 198 -1099 198 -1099 0 1
rlabel polysilicon 198 -1105 198 -1105 0 3
rlabel polysilicon 205 -1099 205 -1099 0 1
rlabel polysilicon 205 -1105 205 -1105 0 3
rlabel polysilicon 212 -1099 212 -1099 0 1
rlabel polysilicon 215 -1099 215 -1099 0 2
rlabel polysilicon 212 -1105 212 -1105 0 3
rlabel polysilicon 219 -1099 219 -1099 0 1
rlabel polysilicon 219 -1105 219 -1105 0 3
rlabel polysilicon 226 -1099 226 -1099 0 1
rlabel polysilicon 226 -1105 226 -1105 0 3
rlabel polysilicon 236 -1099 236 -1099 0 2
rlabel polysilicon 233 -1105 233 -1105 0 3
rlabel polysilicon 236 -1105 236 -1105 0 4
rlabel polysilicon 240 -1105 240 -1105 0 3
rlabel polysilicon 250 -1099 250 -1099 0 2
rlabel polysilicon 247 -1105 247 -1105 0 3
rlabel polysilicon 250 -1105 250 -1105 0 4
rlabel polysilicon 254 -1099 254 -1099 0 1
rlabel polysilicon 254 -1105 254 -1105 0 3
rlabel polysilicon 261 -1105 261 -1105 0 3
rlabel polysilicon 268 -1099 268 -1099 0 1
rlabel polysilicon 268 -1105 268 -1105 0 3
rlabel polysilicon 275 -1099 275 -1099 0 1
rlabel polysilicon 275 -1105 275 -1105 0 3
rlabel polysilicon 282 -1099 282 -1099 0 1
rlabel polysilicon 282 -1105 282 -1105 0 3
rlabel polysilicon 289 -1099 289 -1099 0 1
rlabel polysilicon 289 -1105 289 -1105 0 3
rlabel polysilicon 296 -1099 296 -1099 0 1
rlabel polysilicon 296 -1105 296 -1105 0 3
rlabel polysilicon 303 -1099 303 -1099 0 1
rlabel polysilicon 303 -1105 303 -1105 0 3
rlabel polysilicon 310 -1099 310 -1099 0 1
rlabel polysilicon 310 -1105 310 -1105 0 3
rlabel polysilicon 317 -1099 317 -1099 0 1
rlabel polysilicon 317 -1105 317 -1105 0 3
rlabel polysilicon 324 -1099 324 -1099 0 1
rlabel polysilicon 324 -1105 324 -1105 0 3
rlabel polysilicon 331 -1099 331 -1099 0 1
rlabel polysilicon 331 -1105 331 -1105 0 3
rlabel polysilicon 338 -1099 338 -1099 0 1
rlabel polysilicon 338 -1105 338 -1105 0 3
rlabel polysilicon 341 -1105 341 -1105 0 4
rlabel polysilicon 345 -1099 345 -1099 0 1
rlabel polysilicon 345 -1105 345 -1105 0 3
rlabel polysilicon 352 -1099 352 -1099 0 1
rlabel polysilicon 352 -1105 352 -1105 0 3
rlabel polysilicon 359 -1099 359 -1099 0 1
rlabel polysilicon 359 -1105 359 -1105 0 3
rlabel polysilicon 366 -1099 366 -1099 0 1
rlabel polysilicon 366 -1105 366 -1105 0 3
rlabel polysilicon 373 -1099 373 -1099 0 1
rlabel polysilicon 373 -1105 373 -1105 0 3
rlabel polysilicon 380 -1099 380 -1099 0 1
rlabel polysilicon 380 -1105 380 -1105 0 3
rlabel polysilicon 387 -1099 387 -1099 0 1
rlabel polysilicon 387 -1105 387 -1105 0 3
rlabel polysilicon 394 -1099 394 -1099 0 1
rlabel polysilicon 397 -1099 397 -1099 0 2
rlabel polysilicon 394 -1105 394 -1105 0 3
rlabel polysilicon 397 -1105 397 -1105 0 4
rlabel polysilicon 401 -1099 401 -1099 0 1
rlabel polysilicon 401 -1105 401 -1105 0 3
rlabel polysilicon 408 -1099 408 -1099 0 1
rlabel polysilicon 408 -1105 408 -1105 0 3
rlabel polysilicon 415 -1099 415 -1099 0 1
rlabel polysilicon 415 -1105 415 -1105 0 3
rlabel polysilicon 425 -1105 425 -1105 0 4
rlabel polysilicon 429 -1099 429 -1099 0 1
rlabel polysilicon 429 -1105 429 -1105 0 3
rlabel polysilicon 436 -1099 436 -1099 0 1
rlabel polysilicon 436 -1105 436 -1105 0 3
rlabel polysilicon 443 -1099 443 -1099 0 1
rlabel polysilicon 443 -1105 443 -1105 0 3
rlabel polysilicon 450 -1099 450 -1099 0 1
rlabel polysilicon 450 -1105 450 -1105 0 3
rlabel polysilicon 457 -1099 457 -1099 0 1
rlabel polysilicon 457 -1105 457 -1105 0 3
rlabel polysilicon 464 -1099 464 -1099 0 1
rlabel polysilicon 464 -1105 464 -1105 0 3
rlabel polysilicon 471 -1099 471 -1099 0 1
rlabel polysilicon 471 -1105 471 -1105 0 3
rlabel polysilicon 481 -1099 481 -1099 0 2
rlabel polysilicon 481 -1105 481 -1105 0 4
rlabel polysilicon 485 -1099 485 -1099 0 1
rlabel polysilicon 485 -1105 485 -1105 0 3
rlabel polysilicon 492 -1099 492 -1099 0 1
rlabel polysilicon 492 -1105 492 -1105 0 3
rlabel polysilicon 499 -1099 499 -1099 0 1
rlabel polysilicon 499 -1105 499 -1105 0 3
rlabel polysilicon 506 -1099 506 -1099 0 1
rlabel polysilicon 506 -1105 506 -1105 0 3
rlabel polysilicon 513 -1099 513 -1099 0 1
rlabel polysilicon 516 -1099 516 -1099 0 2
rlabel polysilicon 516 -1105 516 -1105 0 4
rlabel polysilicon 520 -1099 520 -1099 0 1
rlabel polysilicon 520 -1105 520 -1105 0 3
rlabel polysilicon 527 -1099 527 -1099 0 1
rlabel polysilicon 527 -1105 527 -1105 0 3
rlabel polysilicon 534 -1099 534 -1099 0 1
rlabel polysilicon 534 -1105 534 -1105 0 3
rlabel polysilicon 541 -1099 541 -1099 0 1
rlabel polysilicon 541 -1105 541 -1105 0 3
rlabel polysilicon 548 -1099 548 -1099 0 1
rlabel polysilicon 548 -1105 548 -1105 0 3
rlabel polysilicon 555 -1099 555 -1099 0 1
rlabel polysilicon 555 -1105 555 -1105 0 3
rlabel polysilicon 562 -1099 562 -1099 0 1
rlabel polysilicon 562 -1105 562 -1105 0 3
rlabel polysilicon 569 -1099 569 -1099 0 1
rlabel polysilicon 569 -1105 569 -1105 0 3
rlabel polysilicon 576 -1099 576 -1099 0 1
rlabel polysilicon 576 -1105 576 -1105 0 3
rlabel polysilicon 583 -1099 583 -1099 0 1
rlabel polysilicon 583 -1105 583 -1105 0 3
rlabel polysilicon 590 -1099 590 -1099 0 1
rlabel polysilicon 590 -1105 590 -1105 0 3
rlabel polysilicon 597 -1099 597 -1099 0 1
rlabel polysilicon 597 -1105 597 -1105 0 3
rlabel polysilicon 604 -1099 604 -1099 0 1
rlabel polysilicon 604 -1105 604 -1105 0 3
rlabel polysilicon 611 -1099 611 -1099 0 1
rlabel polysilicon 611 -1105 611 -1105 0 3
rlabel polysilicon 618 -1099 618 -1099 0 1
rlabel polysilicon 618 -1105 618 -1105 0 3
rlabel polysilicon 625 -1099 625 -1099 0 1
rlabel polysilicon 628 -1099 628 -1099 0 2
rlabel polysilicon 625 -1105 625 -1105 0 3
rlabel polysilicon 632 -1099 632 -1099 0 1
rlabel polysilicon 632 -1105 632 -1105 0 3
rlabel polysilicon 639 -1099 639 -1099 0 1
rlabel polysilicon 642 -1099 642 -1099 0 2
rlabel polysilicon 639 -1105 639 -1105 0 3
rlabel polysilicon 646 -1099 646 -1099 0 1
rlabel polysilicon 649 -1099 649 -1099 0 2
rlabel polysilicon 649 -1105 649 -1105 0 4
rlabel polysilicon 653 -1099 653 -1099 0 1
rlabel polysilicon 653 -1105 653 -1105 0 3
rlabel polysilicon 660 -1099 660 -1099 0 1
rlabel polysilicon 660 -1105 660 -1105 0 3
rlabel polysilicon 667 -1099 667 -1099 0 1
rlabel polysilicon 667 -1105 667 -1105 0 3
rlabel polysilicon 674 -1099 674 -1099 0 1
rlabel polysilicon 677 -1099 677 -1099 0 2
rlabel polysilicon 674 -1105 674 -1105 0 3
rlabel polysilicon 677 -1105 677 -1105 0 4
rlabel polysilicon 681 -1099 681 -1099 0 1
rlabel polysilicon 681 -1105 681 -1105 0 3
rlabel polysilicon 688 -1099 688 -1099 0 1
rlabel polysilicon 688 -1105 688 -1105 0 3
rlabel polysilicon 691 -1105 691 -1105 0 4
rlabel polysilicon 695 -1099 695 -1099 0 1
rlabel polysilicon 698 -1099 698 -1099 0 2
rlabel polysilicon 695 -1105 695 -1105 0 3
rlabel polysilicon 698 -1105 698 -1105 0 4
rlabel polysilicon 702 -1099 702 -1099 0 1
rlabel polysilicon 702 -1105 702 -1105 0 3
rlabel polysilicon 709 -1099 709 -1099 0 1
rlabel polysilicon 709 -1105 709 -1105 0 3
rlabel polysilicon 716 -1099 716 -1099 0 1
rlabel polysilicon 716 -1105 716 -1105 0 3
rlabel polysilicon 723 -1099 723 -1099 0 1
rlabel polysilicon 723 -1105 723 -1105 0 3
rlabel polysilicon 730 -1099 730 -1099 0 1
rlabel polysilicon 733 -1099 733 -1099 0 2
rlabel polysilicon 730 -1105 730 -1105 0 3
rlabel polysilicon 733 -1105 733 -1105 0 4
rlabel polysilicon 737 -1099 737 -1099 0 1
rlabel polysilicon 737 -1105 737 -1105 0 3
rlabel polysilicon 744 -1099 744 -1099 0 1
rlabel polysilicon 744 -1105 744 -1105 0 3
rlabel polysilicon 751 -1099 751 -1099 0 1
rlabel polysilicon 751 -1105 751 -1105 0 3
rlabel polysilicon 758 -1099 758 -1099 0 1
rlabel polysilicon 758 -1105 758 -1105 0 3
rlabel polysilicon 765 -1099 765 -1099 0 1
rlabel polysilicon 765 -1105 765 -1105 0 3
rlabel polysilicon 772 -1099 772 -1099 0 1
rlabel polysilicon 772 -1105 772 -1105 0 3
rlabel polysilicon 779 -1099 779 -1099 0 1
rlabel polysilicon 779 -1105 779 -1105 0 3
rlabel polysilicon 786 -1099 786 -1099 0 1
rlabel polysilicon 786 -1105 786 -1105 0 3
rlabel polysilicon 793 -1099 793 -1099 0 1
rlabel polysilicon 793 -1105 793 -1105 0 3
rlabel polysilicon 800 -1099 800 -1099 0 1
rlabel polysilicon 803 -1099 803 -1099 0 2
rlabel polysilicon 803 -1105 803 -1105 0 4
rlabel polysilicon 807 -1099 807 -1099 0 1
rlabel polysilicon 807 -1105 807 -1105 0 3
rlabel polysilicon 814 -1099 814 -1099 0 1
rlabel polysilicon 814 -1105 814 -1105 0 3
rlabel polysilicon 821 -1099 821 -1099 0 1
rlabel polysilicon 821 -1105 821 -1105 0 3
rlabel polysilicon 828 -1099 828 -1099 0 1
rlabel polysilicon 828 -1105 828 -1105 0 3
rlabel polysilicon 835 -1099 835 -1099 0 1
rlabel polysilicon 835 -1105 835 -1105 0 3
rlabel polysilicon 842 -1099 842 -1099 0 1
rlabel polysilicon 842 -1105 842 -1105 0 3
rlabel polysilicon 849 -1099 849 -1099 0 1
rlabel polysilicon 849 -1105 849 -1105 0 3
rlabel polysilicon 856 -1099 856 -1099 0 1
rlabel polysilicon 856 -1105 856 -1105 0 3
rlabel polysilicon 863 -1099 863 -1099 0 1
rlabel polysilicon 866 -1099 866 -1099 0 2
rlabel polysilicon 863 -1105 863 -1105 0 3
rlabel polysilicon 866 -1105 866 -1105 0 4
rlabel polysilicon 870 -1099 870 -1099 0 1
rlabel polysilicon 870 -1105 870 -1105 0 3
rlabel polysilicon 877 -1099 877 -1099 0 1
rlabel polysilicon 880 -1099 880 -1099 0 2
rlabel polysilicon 877 -1105 877 -1105 0 3
rlabel polysilicon 880 -1105 880 -1105 0 4
rlabel polysilicon 884 -1099 884 -1099 0 1
rlabel polysilicon 887 -1099 887 -1099 0 2
rlabel polysilicon 887 -1105 887 -1105 0 4
rlabel polysilicon 891 -1099 891 -1099 0 1
rlabel polysilicon 894 -1099 894 -1099 0 2
rlabel polysilicon 891 -1105 891 -1105 0 3
rlabel polysilicon 894 -1105 894 -1105 0 4
rlabel polysilicon 898 -1099 898 -1099 0 1
rlabel polysilicon 898 -1105 898 -1105 0 3
rlabel polysilicon 905 -1099 905 -1099 0 1
rlabel polysilicon 905 -1105 905 -1105 0 3
rlabel polysilicon 912 -1099 912 -1099 0 1
rlabel polysilicon 912 -1105 912 -1105 0 3
rlabel polysilicon 919 -1099 919 -1099 0 1
rlabel polysilicon 919 -1105 919 -1105 0 3
rlabel polysilicon 926 -1099 926 -1099 0 1
rlabel polysilicon 926 -1105 926 -1105 0 3
rlabel polysilicon 933 -1099 933 -1099 0 1
rlabel polysilicon 933 -1105 933 -1105 0 3
rlabel polysilicon 940 -1099 940 -1099 0 1
rlabel polysilicon 940 -1105 940 -1105 0 3
rlabel polysilicon 947 -1099 947 -1099 0 1
rlabel polysilicon 947 -1105 947 -1105 0 3
rlabel polysilicon 954 -1099 954 -1099 0 1
rlabel polysilicon 954 -1105 954 -1105 0 3
rlabel polysilicon 961 -1099 961 -1099 0 1
rlabel polysilicon 961 -1105 961 -1105 0 3
rlabel polysilicon 968 -1099 968 -1099 0 1
rlabel polysilicon 968 -1105 968 -1105 0 3
rlabel polysilicon 975 -1099 975 -1099 0 1
rlabel polysilicon 975 -1105 975 -1105 0 3
rlabel polysilicon 982 -1099 982 -1099 0 1
rlabel polysilicon 982 -1105 982 -1105 0 3
rlabel polysilicon 989 -1099 989 -1099 0 1
rlabel polysilicon 989 -1105 989 -1105 0 3
rlabel polysilicon 996 -1099 996 -1099 0 1
rlabel polysilicon 996 -1105 996 -1105 0 3
rlabel polysilicon 1003 -1099 1003 -1099 0 1
rlabel polysilicon 1006 -1099 1006 -1099 0 2
rlabel polysilicon 1003 -1105 1003 -1105 0 3
rlabel polysilicon 1010 -1099 1010 -1099 0 1
rlabel polysilicon 1010 -1105 1010 -1105 0 3
rlabel polysilicon 1017 -1099 1017 -1099 0 1
rlabel polysilicon 1017 -1105 1017 -1105 0 3
rlabel polysilicon 1024 -1099 1024 -1099 0 1
rlabel polysilicon 1027 -1099 1027 -1099 0 2
rlabel polysilicon 1024 -1105 1024 -1105 0 3
rlabel polysilicon 1031 -1099 1031 -1099 0 1
rlabel polysilicon 1031 -1105 1031 -1105 0 3
rlabel polysilicon 1038 -1099 1038 -1099 0 1
rlabel polysilicon 1038 -1105 1038 -1105 0 3
rlabel polysilicon 1045 -1099 1045 -1099 0 1
rlabel polysilicon 1045 -1105 1045 -1105 0 3
rlabel polysilicon 1048 -1105 1048 -1105 0 4
rlabel polysilicon 1055 -1099 1055 -1099 0 2
rlabel polysilicon 1052 -1105 1052 -1105 0 3
rlabel polysilicon 1055 -1105 1055 -1105 0 4
rlabel polysilicon 1059 -1099 1059 -1099 0 1
rlabel polysilicon 1059 -1105 1059 -1105 0 3
rlabel polysilicon 1066 -1099 1066 -1099 0 1
rlabel polysilicon 1066 -1105 1066 -1105 0 3
rlabel polysilicon 1073 -1099 1073 -1099 0 1
rlabel polysilicon 1073 -1105 1073 -1105 0 3
rlabel polysilicon 1080 -1099 1080 -1099 0 1
rlabel polysilicon 1080 -1105 1080 -1105 0 3
rlabel polysilicon 1087 -1099 1087 -1099 0 1
rlabel polysilicon 1090 -1099 1090 -1099 0 2
rlabel polysilicon 1087 -1105 1087 -1105 0 3
rlabel polysilicon 1094 -1099 1094 -1099 0 1
rlabel polysilicon 1094 -1105 1094 -1105 0 3
rlabel polysilicon 1101 -1099 1101 -1099 0 1
rlabel polysilicon 1101 -1105 1101 -1105 0 3
rlabel polysilicon 1108 -1099 1108 -1099 0 1
rlabel polysilicon 1108 -1105 1108 -1105 0 3
rlabel polysilicon 1115 -1099 1115 -1099 0 1
rlabel polysilicon 1115 -1105 1115 -1105 0 3
rlabel polysilicon 1122 -1099 1122 -1099 0 1
rlabel polysilicon 1122 -1105 1122 -1105 0 3
rlabel polysilicon 1129 -1099 1129 -1099 0 1
rlabel polysilicon 1132 -1099 1132 -1099 0 2
rlabel polysilicon 1129 -1105 1129 -1105 0 3
rlabel polysilicon 1136 -1099 1136 -1099 0 1
rlabel polysilicon 1136 -1105 1136 -1105 0 3
rlabel polysilicon 1143 -1099 1143 -1099 0 1
rlabel polysilicon 1143 -1105 1143 -1105 0 3
rlabel polysilicon 1150 -1099 1150 -1099 0 1
rlabel polysilicon 1150 -1105 1150 -1105 0 3
rlabel polysilicon 1157 -1099 1157 -1099 0 1
rlabel polysilicon 1157 -1105 1157 -1105 0 3
rlabel polysilicon 1164 -1099 1164 -1099 0 1
rlabel polysilicon 1164 -1105 1164 -1105 0 3
rlabel polysilicon 1171 -1099 1171 -1099 0 1
rlabel polysilicon 1171 -1105 1171 -1105 0 3
rlabel polysilicon 1178 -1099 1178 -1099 0 1
rlabel polysilicon 1178 -1105 1178 -1105 0 3
rlabel polysilicon 1185 -1099 1185 -1099 0 1
rlabel polysilicon 1185 -1105 1185 -1105 0 3
rlabel polysilicon 1192 -1099 1192 -1099 0 1
rlabel polysilicon 1192 -1105 1192 -1105 0 3
rlabel polysilicon 1199 -1099 1199 -1099 0 1
rlabel polysilicon 1199 -1105 1199 -1105 0 3
rlabel polysilicon 1206 -1099 1206 -1099 0 1
rlabel polysilicon 1206 -1105 1206 -1105 0 3
rlabel polysilicon 1213 -1099 1213 -1099 0 1
rlabel polysilicon 1213 -1105 1213 -1105 0 3
rlabel polysilicon 1220 -1099 1220 -1099 0 1
rlabel polysilicon 1220 -1105 1220 -1105 0 3
rlabel polysilicon 1227 -1099 1227 -1099 0 1
rlabel polysilicon 1227 -1105 1227 -1105 0 3
rlabel polysilicon 1234 -1099 1234 -1099 0 1
rlabel polysilicon 1234 -1105 1234 -1105 0 3
rlabel polysilicon 1241 -1099 1241 -1099 0 1
rlabel polysilicon 1241 -1105 1241 -1105 0 3
rlabel polysilicon 1248 -1099 1248 -1099 0 1
rlabel polysilicon 1248 -1105 1248 -1105 0 3
rlabel polysilicon 1255 -1099 1255 -1099 0 1
rlabel polysilicon 1255 -1105 1255 -1105 0 3
rlabel polysilicon 1262 -1099 1262 -1099 0 1
rlabel polysilicon 1262 -1105 1262 -1105 0 3
rlabel polysilicon 1269 -1099 1269 -1099 0 1
rlabel polysilicon 1269 -1105 1269 -1105 0 3
rlabel polysilicon 1276 -1099 1276 -1099 0 1
rlabel polysilicon 1276 -1105 1276 -1105 0 3
rlabel polysilicon 1283 -1099 1283 -1099 0 1
rlabel polysilicon 1283 -1105 1283 -1105 0 3
rlabel polysilicon 1290 -1099 1290 -1099 0 1
rlabel polysilicon 1290 -1105 1290 -1105 0 3
rlabel polysilicon 1297 -1099 1297 -1099 0 1
rlabel polysilicon 1297 -1105 1297 -1105 0 3
rlabel polysilicon 1304 -1099 1304 -1099 0 1
rlabel polysilicon 1304 -1105 1304 -1105 0 3
rlabel polysilicon 1311 -1099 1311 -1099 0 1
rlabel polysilicon 1311 -1105 1311 -1105 0 3
rlabel polysilicon 1318 -1099 1318 -1099 0 1
rlabel polysilicon 1318 -1105 1318 -1105 0 3
rlabel polysilicon 1325 -1099 1325 -1099 0 1
rlabel polysilicon 1325 -1105 1325 -1105 0 3
rlabel polysilicon 1332 -1099 1332 -1099 0 1
rlabel polysilicon 1332 -1105 1332 -1105 0 3
rlabel polysilicon 1339 -1099 1339 -1099 0 1
rlabel polysilicon 1339 -1105 1339 -1105 0 3
rlabel polysilicon 1346 -1099 1346 -1099 0 1
rlabel polysilicon 1346 -1105 1346 -1105 0 3
rlabel polysilicon 1353 -1099 1353 -1099 0 1
rlabel polysilicon 1353 -1105 1353 -1105 0 3
rlabel polysilicon 1360 -1099 1360 -1099 0 1
rlabel polysilicon 1360 -1105 1360 -1105 0 3
rlabel polysilicon 1367 -1099 1367 -1099 0 1
rlabel polysilicon 1367 -1105 1367 -1105 0 3
rlabel polysilicon 1374 -1099 1374 -1099 0 1
rlabel polysilicon 1374 -1105 1374 -1105 0 3
rlabel polysilicon 1381 -1099 1381 -1099 0 1
rlabel polysilicon 1384 -1099 1384 -1099 0 2
rlabel polysilicon 1381 -1105 1381 -1105 0 3
rlabel polysilicon 1384 -1105 1384 -1105 0 4
rlabel polysilicon 1388 -1099 1388 -1099 0 1
rlabel polysilicon 1388 -1105 1388 -1105 0 3
rlabel polysilicon 1395 -1099 1395 -1099 0 1
rlabel polysilicon 1395 -1105 1395 -1105 0 3
rlabel polysilicon 1402 -1099 1402 -1099 0 1
rlabel polysilicon 1402 -1105 1402 -1105 0 3
rlabel polysilicon 1409 -1099 1409 -1099 0 1
rlabel polysilicon 1409 -1105 1409 -1105 0 3
rlabel polysilicon 1416 -1099 1416 -1099 0 1
rlabel polysilicon 1416 -1105 1416 -1105 0 3
rlabel polysilicon 1423 -1099 1423 -1099 0 1
rlabel polysilicon 1423 -1105 1423 -1105 0 3
rlabel polysilicon 1430 -1099 1430 -1099 0 1
rlabel polysilicon 1430 -1105 1430 -1105 0 3
rlabel polysilicon 1437 -1099 1437 -1099 0 1
rlabel polysilicon 1437 -1105 1437 -1105 0 3
rlabel polysilicon 1444 -1099 1444 -1099 0 1
rlabel polysilicon 1444 -1105 1444 -1105 0 3
rlabel polysilicon 1451 -1099 1451 -1099 0 1
rlabel polysilicon 1451 -1105 1451 -1105 0 3
rlabel polysilicon 1454 -1105 1454 -1105 0 4
rlabel polysilicon 1458 -1099 1458 -1099 0 1
rlabel polysilicon 1458 -1105 1458 -1105 0 3
rlabel polysilicon 1465 -1099 1465 -1099 0 1
rlabel polysilicon 1465 -1105 1465 -1105 0 3
rlabel polysilicon 1472 -1099 1472 -1099 0 1
rlabel polysilicon 1475 -1099 1475 -1099 0 2
rlabel polysilicon 1475 -1105 1475 -1105 0 4
rlabel polysilicon 1479 -1099 1479 -1099 0 1
rlabel polysilicon 1479 -1105 1479 -1105 0 3
rlabel polysilicon 1486 -1099 1486 -1099 0 1
rlabel polysilicon 1486 -1105 1486 -1105 0 3
rlabel polysilicon 1493 -1099 1493 -1099 0 1
rlabel polysilicon 1493 -1105 1493 -1105 0 3
rlabel polysilicon 1496 -1105 1496 -1105 0 4
rlabel polysilicon 1500 -1099 1500 -1099 0 1
rlabel polysilicon 1500 -1105 1500 -1105 0 3
rlabel polysilicon 1507 -1099 1507 -1099 0 1
rlabel polysilicon 1507 -1105 1507 -1105 0 3
rlabel polysilicon 1514 -1099 1514 -1099 0 1
rlabel polysilicon 1514 -1105 1514 -1105 0 3
rlabel polysilicon 1521 -1099 1521 -1099 0 1
rlabel polysilicon 1521 -1105 1521 -1105 0 3
rlabel polysilicon 1528 -1099 1528 -1099 0 1
rlabel polysilicon 1528 -1105 1528 -1105 0 3
rlabel polysilicon 1535 -1099 1535 -1099 0 1
rlabel polysilicon 1535 -1105 1535 -1105 0 3
rlabel polysilicon 1542 -1099 1542 -1099 0 1
rlabel polysilicon 1542 -1105 1542 -1105 0 3
rlabel polysilicon 1549 -1099 1549 -1099 0 1
rlabel polysilicon 1549 -1105 1549 -1105 0 3
rlabel polysilicon 1556 -1099 1556 -1099 0 1
rlabel polysilicon 1556 -1105 1556 -1105 0 3
rlabel polysilicon 1563 -1099 1563 -1099 0 1
rlabel polysilicon 1563 -1105 1563 -1105 0 3
rlabel polysilicon 1570 -1099 1570 -1099 0 1
rlabel polysilicon 1570 -1105 1570 -1105 0 3
rlabel polysilicon 1577 -1099 1577 -1099 0 1
rlabel polysilicon 1577 -1105 1577 -1105 0 3
rlabel polysilicon 1584 -1099 1584 -1099 0 1
rlabel polysilicon 1584 -1105 1584 -1105 0 3
rlabel polysilicon 1591 -1099 1591 -1099 0 1
rlabel polysilicon 1591 -1105 1591 -1105 0 3
rlabel polysilicon 1598 -1099 1598 -1099 0 1
rlabel polysilicon 1598 -1105 1598 -1105 0 3
rlabel polysilicon 1605 -1099 1605 -1099 0 1
rlabel polysilicon 1605 -1105 1605 -1105 0 3
rlabel polysilicon 1612 -1099 1612 -1099 0 1
rlabel polysilicon 1612 -1105 1612 -1105 0 3
rlabel polysilicon 1619 -1099 1619 -1099 0 1
rlabel polysilicon 1619 -1105 1619 -1105 0 3
rlabel polysilicon 1626 -1099 1626 -1099 0 1
rlabel polysilicon 1626 -1105 1626 -1105 0 3
rlabel polysilicon 1633 -1099 1633 -1099 0 1
rlabel polysilicon 1633 -1105 1633 -1105 0 3
rlabel polysilicon 1640 -1099 1640 -1099 0 1
rlabel polysilicon 1640 -1105 1640 -1105 0 3
rlabel polysilicon 1647 -1099 1647 -1099 0 1
rlabel polysilicon 1647 -1105 1647 -1105 0 3
rlabel polysilicon 1654 -1099 1654 -1099 0 1
rlabel polysilicon 1654 -1105 1654 -1105 0 3
rlabel polysilicon 1675 -1099 1675 -1099 0 1
rlabel polysilicon 1675 -1105 1675 -1105 0 3
rlabel polysilicon 1682 -1099 1682 -1099 0 1
rlabel polysilicon 1682 -1105 1682 -1105 0 3
rlabel polysilicon 1745 -1099 1745 -1099 0 1
rlabel polysilicon 1745 -1105 1745 -1105 0 3
rlabel polysilicon 23 -1218 23 -1218 0 1
rlabel polysilicon 23 -1224 23 -1224 0 3
rlabel polysilicon 30 -1218 30 -1218 0 1
rlabel polysilicon 30 -1224 30 -1224 0 3
rlabel polysilicon 37 -1218 37 -1218 0 1
rlabel polysilicon 37 -1224 37 -1224 0 3
rlabel polysilicon 44 -1218 44 -1218 0 1
rlabel polysilicon 44 -1224 44 -1224 0 3
rlabel polysilicon 51 -1218 51 -1218 0 1
rlabel polysilicon 51 -1224 51 -1224 0 3
rlabel polysilicon 58 -1218 58 -1218 0 1
rlabel polysilicon 58 -1224 58 -1224 0 3
rlabel polysilicon 65 -1218 65 -1218 0 1
rlabel polysilicon 68 -1218 68 -1218 0 2
rlabel polysilicon 65 -1224 65 -1224 0 3
rlabel polysilicon 68 -1224 68 -1224 0 4
rlabel polysilicon 72 -1218 72 -1218 0 1
rlabel polysilicon 72 -1224 72 -1224 0 3
rlabel polysilicon 79 -1218 79 -1218 0 1
rlabel polysilicon 79 -1224 79 -1224 0 3
rlabel polysilicon 86 -1218 86 -1218 0 1
rlabel polysilicon 89 -1218 89 -1218 0 2
rlabel polysilicon 86 -1224 86 -1224 0 3
rlabel polysilicon 89 -1224 89 -1224 0 4
rlabel polysilicon 93 -1218 93 -1218 0 1
rlabel polysilicon 93 -1224 93 -1224 0 3
rlabel polysilicon 100 -1218 100 -1218 0 1
rlabel polysilicon 100 -1224 100 -1224 0 3
rlabel polysilicon 110 -1218 110 -1218 0 2
rlabel polysilicon 107 -1224 107 -1224 0 3
rlabel polysilicon 110 -1224 110 -1224 0 4
rlabel polysilicon 114 -1218 114 -1218 0 1
rlabel polysilicon 114 -1224 114 -1224 0 3
rlabel polysilicon 121 -1218 121 -1218 0 1
rlabel polysilicon 124 -1218 124 -1218 0 2
rlabel polysilicon 121 -1224 121 -1224 0 3
rlabel polysilicon 124 -1224 124 -1224 0 4
rlabel polysilicon 128 -1218 128 -1218 0 1
rlabel polysilicon 128 -1224 128 -1224 0 3
rlabel polysilicon 135 -1218 135 -1218 0 1
rlabel polysilicon 135 -1224 135 -1224 0 3
rlabel polysilicon 142 -1218 142 -1218 0 1
rlabel polysilicon 145 -1218 145 -1218 0 2
rlabel polysilicon 142 -1224 142 -1224 0 3
rlabel polysilicon 145 -1224 145 -1224 0 4
rlabel polysilicon 149 -1218 149 -1218 0 1
rlabel polysilicon 149 -1224 149 -1224 0 3
rlabel polysilicon 156 -1218 156 -1218 0 1
rlabel polysilicon 156 -1224 156 -1224 0 3
rlabel polysilicon 163 -1218 163 -1218 0 1
rlabel polysilicon 163 -1224 163 -1224 0 3
rlabel polysilicon 170 -1218 170 -1218 0 1
rlabel polysilicon 173 -1218 173 -1218 0 2
rlabel polysilicon 170 -1224 170 -1224 0 3
rlabel polysilicon 173 -1224 173 -1224 0 4
rlabel polysilicon 177 -1218 177 -1218 0 1
rlabel polysilicon 180 -1218 180 -1218 0 2
rlabel polysilicon 177 -1224 177 -1224 0 3
rlabel polysilicon 180 -1224 180 -1224 0 4
rlabel polysilicon 184 -1218 184 -1218 0 1
rlabel polysilicon 184 -1224 184 -1224 0 3
rlabel polysilicon 191 -1218 191 -1218 0 1
rlabel polysilicon 191 -1224 191 -1224 0 3
rlabel polysilicon 198 -1218 198 -1218 0 1
rlabel polysilicon 198 -1224 198 -1224 0 3
rlabel polysilicon 205 -1218 205 -1218 0 1
rlabel polysilicon 205 -1224 205 -1224 0 3
rlabel polysilicon 212 -1218 212 -1218 0 1
rlabel polysilicon 212 -1224 212 -1224 0 3
rlabel polysilicon 219 -1218 219 -1218 0 1
rlabel polysilicon 219 -1224 219 -1224 0 3
rlabel polysilicon 226 -1218 226 -1218 0 1
rlabel polysilicon 229 -1218 229 -1218 0 2
rlabel polysilicon 226 -1224 226 -1224 0 3
rlabel polysilicon 233 -1218 233 -1218 0 1
rlabel polysilicon 233 -1224 233 -1224 0 3
rlabel polysilicon 240 -1218 240 -1218 0 1
rlabel polysilicon 243 -1218 243 -1218 0 2
rlabel polysilicon 243 -1224 243 -1224 0 4
rlabel polysilicon 247 -1218 247 -1218 0 1
rlabel polysilicon 247 -1224 247 -1224 0 3
rlabel polysilicon 254 -1218 254 -1218 0 1
rlabel polysilicon 254 -1224 254 -1224 0 3
rlabel polysilicon 264 -1218 264 -1218 0 2
rlabel polysilicon 264 -1224 264 -1224 0 4
rlabel polysilicon 268 -1218 268 -1218 0 1
rlabel polysilicon 268 -1224 268 -1224 0 3
rlabel polysilicon 275 -1218 275 -1218 0 1
rlabel polysilicon 275 -1224 275 -1224 0 3
rlabel polysilicon 282 -1218 282 -1218 0 1
rlabel polysilicon 282 -1224 282 -1224 0 3
rlabel polysilicon 289 -1218 289 -1218 0 1
rlabel polysilicon 289 -1224 289 -1224 0 3
rlabel polysilicon 296 -1218 296 -1218 0 1
rlabel polysilicon 296 -1224 296 -1224 0 3
rlabel polysilicon 303 -1218 303 -1218 0 1
rlabel polysilicon 303 -1224 303 -1224 0 3
rlabel polysilicon 310 -1218 310 -1218 0 1
rlabel polysilicon 310 -1224 310 -1224 0 3
rlabel polysilicon 317 -1218 317 -1218 0 1
rlabel polysilicon 317 -1224 317 -1224 0 3
rlabel polysilicon 324 -1218 324 -1218 0 1
rlabel polysilicon 324 -1224 324 -1224 0 3
rlabel polysilicon 331 -1218 331 -1218 0 1
rlabel polysilicon 331 -1224 331 -1224 0 3
rlabel polysilicon 338 -1218 338 -1218 0 1
rlabel polysilicon 338 -1224 338 -1224 0 3
rlabel polysilicon 345 -1218 345 -1218 0 1
rlabel polysilicon 345 -1224 345 -1224 0 3
rlabel polysilicon 352 -1218 352 -1218 0 1
rlabel polysilicon 352 -1224 352 -1224 0 3
rlabel polysilicon 359 -1218 359 -1218 0 1
rlabel polysilicon 359 -1224 359 -1224 0 3
rlabel polysilicon 366 -1218 366 -1218 0 1
rlabel polysilicon 366 -1224 366 -1224 0 3
rlabel polysilicon 373 -1218 373 -1218 0 1
rlabel polysilicon 373 -1224 373 -1224 0 3
rlabel polysilicon 380 -1218 380 -1218 0 1
rlabel polysilicon 380 -1224 380 -1224 0 3
rlabel polysilicon 387 -1218 387 -1218 0 1
rlabel polysilicon 387 -1224 387 -1224 0 3
rlabel polysilicon 394 -1218 394 -1218 0 1
rlabel polysilicon 394 -1224 394 -1224 0 3
rlabel polysilicon 401 -1218 401 -1218 0 1
rlabel polysilicon 401 -1224 401 -1224 0 3
rlabel polysilicon 408 -1218 408 -1218 0 1
rlabel polysilicon 408 -1224 408 -1224 0 3
rlabel polysilicon 415 -1218 415 -1218 0 1
rlabel polysilicon 415 -1224 415 -1224 0 3
rlabel polysilicon 422 -1218 422 -1218 0 1
rlabel polysilicon 422 -1224 422 -1224 0 3
rlabel polysilicon 429 -1218 429 -1218 0 1
rlabel polysilicon 429 -1224 429 -1224 0 3
rlabel polysilicon 436 -1218 436 -1218 0 1
rlabel polysilicon 439 -1218 439 -1218 0 2
rlabel polysilicon 436 -1224 436 -1224 0 3
rlabel polysilicon 443 -1218 443 -1218 0 1
rlabel polysilicon 443 -1224 443 -1224 0 3
rlabel polysilicon 450 -1218 450 -1218 0 1
rlabel polysilicon 450 -1224 450 -1224 0 3
rlabel polysilicon 457 -1218 457 -1218 0 1
rlabel polysilicon 457 -1224 457 -1224 0 3
rlabel polysilicon 464 -1218 464 -1218 0 1
rlabel polysilicon 464 -1224 464 -1224 0 3
rlabel polysilicon 471 -1218 471 -1218 0 1
rlabel polysilicon 471 -1224 471 -1224 0 3
rlabel polysilicon 478 -1218 478 -1218 0 1
rlabel polysilicon 478 -1224 478 -1224 0 3
rlabel polysilicon 485 -1218 485 -1218 0 1
rlabel polysilicon 485 -1224 485 -1224 0 3
rlabel polysilicon 492 -1218 492 -1218 0 1
rlabel polysilicon 492 -1224 492 -1224 0 3
rlabel polysilicon 499 -1218 499 -1218 0 1
rlabel polysilicon 499 -1224 499 -1224 0 3
rlabel polysilicon 506 -1224 506 -1224 0 3
rlabel polysilicon 509 -1224 509 -1224 0 4
rlabel polysilicon 513 -1218 513 -1218 0 1
rlabel polysilicon 513 -1224 513 -1224 0 3
rlabel polysilicon 520 -1218 520 -1218 0 1
rlabel polysilicon 520 -1224 520 -1224 0 3
rlabel polysilicon 527 -1218 527 -1218 0 1
rlabel polysilicon 527 -1224 527 -1224 0 3
rlabel polysilicon 534 -1218 534 -1218 0 1
rlabel polysilicon 534 -1224 534 -1224 0 3
rlabel polysilicon 541 -1218 541 -1218 0 1
rlabel polysilicon 544 -1218 544 -1218 0 2
rlabel polysilicon 541 -1224 541 -1224 0 3
rlabel polysilicon 548 -1218 548 -1218 0 1
rlabel polysilicon 548 -1224 548 -1224 0 3
rlabel polysilicon 555 -1218 555 -1218 0 1
rlabel polysilicon 555 -1224 555 -1224 0 3
rlabel polysilicon 562 -1218 562 -1218 0 1
rlabel polysilicon 562 -1224 562 -1224 0 3
rlabel polysilicon 565 -1224 565 -1224 0 4
rlabel polysilicon 569 -1218 569 -1218 0 1
rlabel polysilicon 569 -1224 569 -1224 0 3
rlabel polysilicon 576 -1218 576 -1218 0 1
rlabel polysilicon 576 -1224 576 -1224 0 3
rlabel polysilicon 583 -1218 583 -1218 0 1
rlabel polysilicon 583 -1224 583 -1224 0 3
rlabel polysilicon 590 -1218 590 -1218 0 1
rlabel polysilicon 590 -1224 590 -1224 0 3
rlabel polysilicon 597 -1218 597 -1218 0 1
rlabel polysilicon 597 -1224 597 -1224 0 3
rlabel polysilicon 604 -1218 604 -1218 0 1
rlabel polysilicon 604 -1224 604 -1224 0 3
rlabel polysilicon 607 -1224 607 -1224 0 4
rlabel polysilicon 611 -1218 611 -1218 0 1
rlabel polysilicon 611 -1224 611 -1224 0 3
rlabel polysilicon 618 -1218 618 -1218 0 1
rlabel polysilicon 618 -1224 618 -1224 0 3
rlabel polysilicon 625 -1218 625 -1218 0 1
rlabel polysilicon 625 -1224 625 -1224 0 3
rlabel polysilicon 635 -1218 635 -1218 0 2
rlabel polysilicon 632 -1224 632 -1224 0 3
rlabel polysilicon 635 -1224 635 -1224 0 4
rlabel polysilicon 639 -1218 639 -1218 0 1
rlabel polysilicon 639 -1224 639 -1224 0 3
rlabel polysilicon 646 -1218 646 -1218 0 1
rlabel polysilicon 649 -1218 649 -1218 0 2
rlabel polysilicon 656 -1218 656 -1218 0 2
rlabel polysilicon 656 -1224 656 -1224 0 4
rlabel polysilicon 660 -1218 660 -1218 0 1
rlabel polysilicon 660 -1224 660 -1224 0 3
rlabel polysilicon 667 -1218 667 -1218 0 1
rlabel polysilicon 667 -1224 667 -1224 0 3
rlabel polysilicon 674 -1218 674 -1218 0 1
rlabel polysilicon 674 -1224 674 -1224 0 3
rlabel polysilicon 681 -1218 681 -1218 0 1
rlabel polysilicon 681 -1224 681 -1224 0 3
rlabel polysilicon 688 -1218 688 -1218 0 1
rlabel polysilicon 688 -1224 688 -1224 0 3
rlabel polysilicon 695 -1218 695 -1218 0 1
rlabel polysilicon 698 -1218 698 -1218 0 2
rlabel polysilicon 695 -1224 695 -1224 0 3
rlabel polysilicon 698 -1224 698 -1224 0 4
rlabel polysilicon 702 -1218 702 -1218 0 1
rlabel polysilicon 702 -1224 702 -1224 0 3
rlabel polysilicon 705 -1224 705 -1224 0 4
rlabel polysilicon 709 -1218 709 -1218 0 1
rlabel polysilicon 709 -1224 709 -1224 0 3
rlabel polysilicon 716 -1218 716 -1218 0 1
rlabel polysilicon 716 -1224 716 -1224 0 3
rlabel polysilicon 723 -1218 723 -1218 0 1
rlabel polysilicon 723 -1224 723 -1224 0 3
rlabel polysilicon 730 -1218 730 -1218 0 1
rlabel polysilicon 730 -1224 730 -1224 0 3
rlabel polysilicon 737 -1218 737 -1218 0 1
rlabel polysilicon 740 -1218 740 -1218 0 2
rlabel polysilicon 737 -1224 737 -1224 0 3
rlabel polysilicon 740 -1224 740 -1224 0 4
rlabel polysilicon 744 -1218 744 -1218 0 1
rlabel polysilicon 744 -1224 744 -1224 0 3
rlabel polysilicon 751 -1218 751 -1218 0 1
rlabel polysilicon 751 -1224 751 -1224 0 3
rlabel polysilicon 758 -1218 758 -1218 0 1
rlabel polysilicon 758 -1224 758 -1224 0 3
rlabel polysilicon 765 -1218 765 -1218 0 1
rlabel polysilicon 768 -1218 768 -1218 0 2
rlabel polysilicon 768 -1224 768 -1224 0 4
rlabel polysilicon 772 -1218 772 -1218 0 1
rlabel polysilicon 772 -1224 772 -1224 0 3
rlabel polysilicon 779 -1218 779 -1218 0 1
rlabel polysilicon 779 -1224 779 -1224 0 3
rlabel polysilicon 786 -1218 786 -1218 0 1
rlabel polysilicon 786 -1224 786 -1224 0 3
rlabel polysilicon 793 -1218 793 -1218 0 1
rlabel polysilicon 796 -1218 796 -1218 0 2
rlabel polysilicon 793 -1224 793 -1224 0 3
rlabel polysilicon 796 -1224 796 -1224 0 4
rlabel polysilicon 800 -1218 800 -1218 0 1
rlabel polysilicon 800 -1224 800 -1224 0 3
rlabel polysilicon 807 -1218 807 -1218 0 1
rlabel polysilicon 807 -1224 807 -1224 0 3
rlabel polysilicon 814 -1218 814 -1218 0 1
rlabel polysilicon 817 -1218 817 -1218 0 2
rlabel polysilicon 814 -1224 814 -1224 0 3
rlabel polysilicon 817 -1224 817 -1224 0 4
rlabel polysilicon 821 -1218 821 -1218 0 1
rlabel polysilicon 824 -1218 824 -1218 0 2
rlabel polysilicon 821 -1224 821 -1224 0 3
rlabel polysilicon 828 -1218 828 -1218 0 1
rlabel polysilicon 831 -1218 831 -1218 0 2
rlabel polysilicon 828 -1224 828 -1224 0 3
rlabel polysilicon 831 -1224 831 -1224 0 4
rlabel polysilicon 835 -1218 835 -1218 0 1
rlabel polysilicon 835 -1224 835 -1224 0 3
rlabel polysilicon 842 -1218 842 -1218 0 1
rlabel polysilicon 842 -1224 842 -1224 0 3
rlabel polysilicon 849 -1218 849 -1218 0 1
rlabel polysilicon 849 -1224 849 -1224 0 3
rlabel polysilicon 856 -1218 856 -1218 0 1
rlabel polysilicon 859 -1218 859 -1218 0 2
rlabel polysilicon 856 -1224 856 -1224 0 3
rlabel polysilicon 859 -1224 859 -1224 0 4
rlabel polysilicon 863 -1218 863 -1218 0 1
rlabel polysilicon 863 -1224 863 -1224 0 3
rlabel polysilicon 870 -1218 870 -1218 0 1
rlabel polysilicon 870 -1224 870 -1224 0 3
rlabel polysilicon 877 -1218 877 -1218 0 1
rlabel polysilicon 877 -1224 877 -1224 0 3
rlabel polysilicon 884 -1218 884 -1218 0 1
rlabel polysilicon 884 -1224 884 -1224 0 3
rlabel polysilicon 891 -1218 891 -1218 0 1
rlabel polysilicon 894 -1218 894 -1218 0 2
rlabel polysilicon 891 -1224 891 -1224 0 3
rlabel polysilicon 894 -1224 894 -1224 0 4
rlabel polysilicon 898 -1218 898 -1218 0 1
rlabel polysilicon 898 -1224 898 -1224 0 3
rlabel polysilicon 905 -1218 905 -1218 0 1
rlabel polysilicon 905 -1224 905 -1224 0 3
rlabel polysilicon 912 -1218 912 -1218 0 1
rlabel polysilicon 912 -1224 912 -1224 0 3
rlabel polysilicon 919 -1218 919 -1218 0 1
rlabel polysilicon 919 -1224 919 -1224 0 3
rlabel polysilicon 926 -1218 926 -1218 0 1
rlabel polysilicon 929 -1218 929 -1218 0 2
rlabel polysilicon 926 -1224 926 -1224 0 3
rlabel polysilicon 929 -1224 929 -1224 0 4
rlabel polysilicon 933 -1218 933 -1218 0 1
rlabel polysilicon 933 -1224 933 -1224 0 3
rlabel polysilicon 940 -1218 940 -1218 0 1
rlabel polysilicon 940 -1224 940 -1224 0 3
rlabel polysilicon 947 -1218 947 -1218 0 1
rlabel polysilicon 950 -1218 950 -1218 0 2
rlabel polysilicon 950 -1224 950 -1224 0 4
rlabel polysilicon 954 -1218 954 -1218 0 1
rlabel polysilicon 954 -1224 954 -1224 0 3
rlabel polysilicon 961 -1218 961 -1218 0 1
rlabel polysilicon 961 -1224 961 -1224 0 3
rlabel polysilicon 968 -1218 968 -1218 0 1
rlabel polysilicon 968 -1224 968 -1224 0 3
rlabel polysilicon 975 -1218 975 -1218 0 1
rlabel polysilicon 975 -1224 975 -1224 0 3
rlabel polysilicon 982 -1218 982 -1218 0 1
rlabel polysilicon 982 -1224 982 -1224 0 3
rlabel polysilicon 989 -1218 989 -1218 0 1
rlabel polysilicon 989 -1224 989 -1224 0 3
rlabel polysilicon 996 -1218 996 -1218 0 1
rlabel polysilicon 996 -1224 996 -1224 0 3
rlabel polysilicon 1003 -1218 1003 -1218 0 1
rlabel polysilicon 1003 -1224 1003 -1224 0 3
rlabel polysilicon 1010 -1218 1010 -1218 0 1
rlabel polysilicon 1010 -1224 1010 -1224 0 3
rlabel polysilicon 1017 -1218 1017 -1218 0 1
rlabel polysilicon 1017 -1224 1017 -1224 0 3
rlabel polysilicon 1024 -1218 1024 -1218 0 1
rlabel polysilicon 1024 -1224 1024 -1224 0 3
rlabel polysilicon 1031 -1218 1031 -1218 0 1
rlabel polysilicon 1031 -1224 1031 -1224 0 3
rlabel polysilicon 1038 -1218 1038 -1218 0 1
rlabel polysilicon 1038 -1224 1038 -1224 0 3
rlabel polysilicon 1045 -1218 1045 -1218 0 1
rlabel polysilicon 1045 -1224 1045 -1224 0 3
rlabel polysilicon 1055 -1218 1055 -1218 0 2
rlabel polysilicon 1052 -1224 1052 -1224 0 3
rlabel polysilicon 1055 -1224 1055 -1224 0 4
rlabel polysilicon 1059 -1218 1059 -1218 0 1
rlabel polysilicon 1059 -1224 1059 -1224 0 3
rlabel polysilicon 1066 -1218 1066 -1218 0 1
rlabel polysilicon 1066 -1224 1066 -1224 0 3
rlabel polysilicon 1073 -1218 1073 -1218 0 1
rlabel polysilicon 1073 -1224 1073 -1224 0 3
rlabel polysilicon 1080 -1218 1080 -1218 0 1
rlabel polysilicon 1080 -1224 1080 -1224 0 3
rlabel polysilicon 1087 -1218 1087 -1218 0 1
rlabel polysilicon 1087 -1224 1087 -1224 0 3
rlabel polysilicon 1094 -1218 1094 -1218 0 1
rlabel polysilicon 1094 -1224 1094 -1224 0 3
rlabel polysilicon 1101 -1218 1101 -1218 0 1
rlabel polysilicon 1101 -1224 1101 -1224 0 3
rlabel polysilicon 1108 -1218 1108 -1218 0 1
rlabel polysilicon 1108 -1224 1108 -1224 0 3
rlabel polysilicon 1115 -1218 1115 -1218 0 1
rlabel polysilicon 1115 -1224 1115 -1224 0 3
rlabel polysilicon 1122 -1218 1122 -1218 0 1
rlabel polysilicon 1122 -1224 1122 -1224 0 3
rlabel polysilicon 1129 -1218 1129 -1218 0 1
rlabel polysilicon 1129 -1224 1129 -1224 0 3
rlabel polysilicon 1136 -1218 1136 -1218 0 1
rlabel polysilicon 1136 -1224 1136 -1224 0 3
rlabel polysilicon 1143 -1218 1143 -1218 0 1
rlabel polysilicon 1143 -1224 1143 -1224 0 3
rlabel polysilicon 1150 -1218 1150 -1218 0 1
rlabel polysilicon 1150 -1224 1150 -1224 0 3
rlabel polysilicon 1157 -1218 1157 -1218 0 1
rlabel polysilicon 1157 -1224 1157 -1224 0 3
rlabel polysilicon 1164 -1218 1164 -1218 0 1
rlabel polysilicon 1164 -1224 1164 -1224 0 3
rlabel polysilicon 1171 -1218 1171 -1218 0 1
rlabel polysilicon 1171 -1224 1171 -1224 0 3
rlabel polysilicon 1178 -1218 1178 -1218 0 1
rlabel polysilicon 1178 -1224 1178 -1224 0 3
rlabel polysilicon 1185 -1218 1185 -1218 0 1
rlabel polysilicon 1185 -1224 1185 -1224 0 3
rlabel polysilicon 1192 -1218 1192 -1218 0 1
rlabel polysilicon 1192 -1224 1192 -1224 0 3
rlabel polysilicon 1199 -1218 1199 -1218 0 1
rlabel polysilicon 1199 -1224 1199 -1224 0 3
rlabel polysilicon 1206 -1218 1206 -1218 0 1
rlabel polysilicon 1206 -1224 1206 -1224 0 3
rlabel polysilicon 1213 -1218 1213 -1218 0 1
rlabel polysilicon 1213 -1224 1213 -1224 0 3
rlabel polysilicon 1220 -1218 1220 -1218 0 1
rlabel polysilicon 1220 -1224 1220 -1224 0 3
rlabel polysilicon 1227 -1218 1227 -1218 0 1
rlabel polysilicon 1227 -1224 1227 -1224 0 3
rlabel polysilicon 1234 -1218 1234 -1218 0 1
rlabel polysilicon 1234 -1224 1234 -1224 0 3
rlabel polysilicon 1241 -1218 1241 -1218 0 1
rlabel polysilicon 1241 -1224 1241 -1224 0 3
rlabel polysilicon 1248 -1218 1248 -1218 0 1
rlabel polysilicon 1248 -1224 1248 -1224 0 3
rlabel polysilicon 1255 -1218 1255 -1218 0 1
rlabel polysilicon 1255 -1224 1255 -1224 0 3
rlabel polysilicon 1262 -1218 1262 -1218 0 1
rlabel polysilicon 1262 -1224 1262 -1224 0 3
rlabel polysilicon 1269 -1218 1269 -1218 0 1
rlabel polysilicon 1269 -1224 1269 -1224 0 3
rlabel polysilicon 1276 -1218 1276 -1218 0 1
rlabel polysilicon 1276 -1224 1276 -1224 0 3
rlabel polysilicon 1283 -1218 1283 -1218 0 1
rlabel polysilicon 1283 -1224 1283 -1224 0 3
rlabel polysilicon 1290 -1218 1290 -1218 0 1
rlabel polysilicon 1290 -1224 1290 -1224 0 3
rlabel polysilicon 1297 -1218 1297 -1218 0 1
rlabel polysilicon 1297 -1224 1297 -1224 0 3
rlabel polysilicon 1304 -1218 1304 -1218 0 1
rlabel polysilicon 1311 -1218 1311 -1218 0 1
rlabel polysilicon 1311 -1224 1311 -1224 0 3
rlabel polysilicon 1314 -1224 1314 -1224 0 4
rlabel polysilicon 1318 -1218 1318 -1218 0 1
rlabel polysilicon 1318 -1224 1318 -1224 0 3
rlabel polysilicon 1325 -1218 1325 -1218 0 1
rlabel polysilicon 1325 -1224 1325 -1224 0 3
rlabel polysilicon 1332 -1218 1332 -1218 0 1
rlabel polysilicon 1332 -1224 1332 -1224 0 3
rlabel polysilicon 1339 -1218 1339 -1218 0 1
rlabel polysilicon 1339 -1224 1339 -1224 0 3
rlabel polysilicon 1346 -1218 1346 -1218 0 1
rlabel polysilicon 1346 -1224 1346 -1224 0 3
rlabel polysilicon 1353 -1218 1353 -1218 0 1
rlabel polysilicon 1353 -1224 1353 -1224 0 3
rlabel polysilicon 1360 -1218 1360 -1218 0 1
rlabel polysilicon 1360 -1224 1360 -1224 0 3
rlabel polysilicon 1367 -1218 1367 -1218 0 1
rlabel polysilicon 1367 -1224 1367 -1224 0 3
rlabel polysilicon 1374 -1218 1374 -1218 0 1
rlabel polysilicon 1374 -1224 1374 -1224 0 3
rlabel polysilicon 1381 -1218 1381 -1218 0 1
rlabel polysilicon 1381 -1224 1381 -1224 0 3
rlabel polysilicon 1388 -1218 1388 -1218 0 1
rlabel polysilicon 1388 -1224 1388 -1224 0 3
rlabel polysilicon 1395 -1218 1395 -1218 0 1
rlabel polysilicon 1395 -1224 1395 -1224 0 3
rlabel polysilicon 1402 -1218 1402 -1218 0 1
rlabel polysilicon 1402 -1224 1402 -1224 0 3
rlabel polysilicon 1409 -1218 1409 -1218 0 1
rlabel polysilicon 1409 -1224 1409 -1224 0 3
rlabel polysilicon 1416 -1218 1416 -1218 0 1
rlabel polysilicon 1416 -1224 1416 -1224 0 3
rlabel polysilicon 1423 -1218 1423 -1218 0 1
rlabel polysilicon 1423 -1224 1423 -1224 0 3
rlabel polysilicon 1430 -1218 1430 -1218 0 1
rlabel polysilicon 1430 -1224 1430 -1224 0 3
rlabel polysilicon 1437 -1218 1437 -1218 0 1
rlabel polysilicon 1437 -1224 1437 -1224 0 3
rlabel polysilicon 1444 -1218 1444 -1218 0 1
rlabel polysilicon 1444 -1224 1444 -1224 0 3
rlabel polysilicon 1451 -1218 1451 -1218 0 1
rlabel polysilicon 1451 -1224 1451 -1224 0 3
rlabel polysilicon 1458 -1218 1458 -1218 0 1
rlabel polysilicon 1458 -1224 1458 -1224 0 3
rlabel polysilicon 1465 -1218 1465 -1218 0 1
rlabel polysilicon 1465 -1224 1465 -1224 0 3
rlabel polysilicon 1472 -1218 1472 -1218 0 1
rlabel polysilicon 1472 -1224 1472 -1224 0 3
rlabel polysilicon 1479 -1218 1479 -1218 0 1
rlabel polysilicon 1479 -1224 1479 -1224 0 3
rlabel polysilicon 1486 -1218 1486 -1218 0 1
rlabel polysilicon 1486 -1224 1486 -1224 0 3
rlabel polysilicon 1493 -1218 1493 -1218 0 1
rlabel polysilicon 1493 -1224 1493 -1224 0 3
rlabel polysilicon 1500 -1218 1500 -1218 0 1
rlabel polysilicon 1500 -1224 1500 -1224 0 3
rlabel polysilicon 1507 -1218 1507 -1218 0 1
rlabel polysilicon 1507 -1224 1507 -1224 0 3
rlabel polysilicon 1514 -1218 1514 -1218 0 1
rlabel polysilicon 1514 -1224 1514 -1224 0 3
rlabel polysilicon 1521 -1218 1521 -1218 0 1
rlabel polysilicon 1521 -1224 1521 -1224 0 3
rlabel polysilicon 1528 -1218 1528 -1218 0 1
rlabel polysilicon 1528 -1224 1528 -1224 0 3
rlabel polysilicon 1535 -1218 1535 -1218 0 1
rlabel polysilicon 1535 -1224 1535 -1224 0 3
rlabel polysilicon 1542 -1218 1542 -1218 0 1
rlabel polysilicon 1542 -1224 1542 -1224 0 3
rlabel polysilicon 1549 -1218 1549 -1218 0 1
rlabel polysilicon 1549 -1224 1549 -1224 0 3
rlabel polysilicon 1556 -1218 1556 -1218 0 1
rlabel polysilicon 1556 -1224 1556 -1224 0 3
rlabel polysilicon 1563 -1218 1563 -1218 0 1
rlabel polysilicon 1563 -1224 1563 -1224 0 3
rlabel polysilicon 1570 -1218 1570 -1218 0 1
rlabel polysilicon 1570 -1224 1570 -1224 0 3
rlabel polysilicon 1577 -1218 1577 -1218 0 1
rlabel polysilicon 1577 -1224 1577 -1224 0 3
rlabel polysilicon 1584 -1218 1584 -1218 0 1
rlabel polysilicon 1584 -1224 1584 -1224 0 3
rlabel polysilicon 1591 -1218 1591 -1218 0 1
rlabel polysilicon 1591 -1224 1591 -1224 0 3
rlabel polysilicon 1598 -1218 1598 -1218 0 1
rlabel polysilicon 1598 -1224 1598 -1224 0 3
rlabel polysilicon 1605 -1218 1605 -1218 0 1
rlabel polysilicon 1605 -1224 1605 -1224 0 3
rlabel polysilicon 1612 -1218 1612 -1218 0 1
rlabel polysilicon 1612 -1224 1612 -1224 0 3
rlabel polysilicon 1619 -1218 1619 -1218 0 1
rlabel polysilicon 1619 -1224 1619 -1224 0 3
rlabel polysilicon 1626 -1218 1626 -1218 0 1
rlabel polysilicon 1626 -1224 1626 -1224 0 3
rlabel polysilicon 1633 -1218 1633 -1218 0 1
rlabel polysilicon 1633 -1224 1633 -1224 0 3
rlabel polysilicon 1640 -1218 1640 -1218 0 1
rlabel polysilicon 1640 -1224 1640 -1224 0 3
rlabel polysilicon 1647 -1218 1647 -1218 0 1
rlabel polysilicon 1647 -1224 1647 -1224 0 3
rlabel polysilicon 1654 -1218 1654 -1218 0 1
rlabel polysilicon 1654 -1224 1654 -1224 0 3
rlabel polysilicon 1661 -1218 1661 -1218 0 1
rlabel polysilicon 1661 -1224 1661 -1224 0 3
rlabel polysilicon 1668 -1218 1668 -1218 0 1
rlabel polysilicon 1668 -1224 1668 -1224 0 3
rlabel polysilicon 1675 -1218 1675 -1218 0 1
rlabel polysilicon 1675 -1224 1675 -1224 0 3
rlabel polysilicon 1682 -1218 1682 -1218 0 1
rlabel polysilicon 1682 -1224 1682 -1224 0 3
rlabel polysilicon 1689 -1218 1689 -1218 0 1
rlabel polysilicon 1689 -1224 1689 -1224 0 3
rlabel polysilicon 1696 -1218 1696 -1218 0 1
rlabel polysilicon 1696 -1224 1696 -1224 0 3
rlabel polysilicon 1703 -1218 1703 -1218 0 1
rlabel polysilicon 1703 -1224 1703 -1224 0 3
rlabel polysilicon 1710 -1218 1710 -1218 0 1
rlabel polysilicon 1710 -1224 1710 -1224 0 3
rlabel polysilicon 1717 -1218 1717 -1218 0 1
rlabel polysilicon 1717 -1224 1717 -1224 0 3
rlabel polysilicon 1724 -1218 1724 -1218 0 1
rlabel polysilicon 1724 -1224 1724 -1224 0 3
rlabel polysilicon 1731 -1218 1731 -1218 0 1
rlabel polysilicon 1731 -1224 1731 -1224 0 3
rlabel polysilicon 1738 -1218 1738 -1218 0 1
rlabel polysilicon 1738 -1224 1738 -1224 0 3
rlabel polysilicon 1745 -1218 1745 -1218 0 1
rlabel polysilicon 1748 -1218 1748 -1218 0 2
rlabel polysilicon 1745 -1224 1745 -1224 0 3
rlabel polysilicon 1748 -1224 1748 -1224 0 4
rlabel polysilicon 1752 -1218 1752 -1218 0 1
rlabel polysilicon 1752 -1224 1752 -1224 0 3
rlabel polysilicon 1759 -1218 1759 -1218 0 1
rlabel polysilicon 1759 -1224 1759 -1224 0 3
rlabel polysilicon 1766 -1218 1766 -1218 0 1
rlabel polysilicon 1769 -1218 1769 -1218 0 2
rlabel polysilicon 1766 -1224 1766 -1224 0 3
rlabel polysilicon 1769 -1224 1769 -1224 0 4
rlabel polysilicon 1776 -1224 1776 -1224 0 4
rlabel polysilicon 1780 -1218 1780 -1218 0 1
rlabel polysilicon 1780 -1224 1780 -1224 0 3
rlabel polysilicon 1787 -1218 1787 -1218 0 1
rlabel polysilicon 1787 -1224 1787 -1224 0 3
rlabel polysilicon 16 -1361 16 -1361 0 1
rlabel polysilicon 16 -1367 16 -1367 0 3
rlabel polysilicon 23 -1361 23 -1361 0 1
rlabel polysilicon 23 -1367 23 -1367 0 3
rlabel polysilicon 30 -1361 30 -1361 0 1
rlabel polysilicon 30 -1367 30 -1367 0 3
rlabel polysilicon 44 -1361 44 -1361 0 1
rlabel polysilicon 44 -1367 44 -1367 0 3
rlabel polysilicon 54 -1361 54 -1361 0 2
rlabel polysilicon 51 -1367 51 -1367 0 3
rlabel polysilicon 54 -1367 54 -1367 0 4
rlabel polysilicon 58 -1361 58 -1361 0 1
rlabel polysilicon 61 -1361 61 -1361 0 2
rlabel polysilicon 61 -1367 61 -1367 0 4
rlabel polysilicon 65 -1361 65 -1361 0 1
rlabel polysilicon 65 -1367 65 -1367 0 3
rlabel polysilicon 72 -1361 72 -1361 0 1
rlabel polysilicon 72 -1367 72 -1367 0 3
rlabel polysilicon 82 -1361 82 -1361 0 2
rlabel polysilicon 79 -1367 79 -1367 0 3
rlabel polysilicon 82 -1367 82 -1367 0 4
rlabel polysilicon 86 -1361 86 -1361 0 1
rlabel polysilicon 86 -1367 86 -1367 0 3
rlabel polysilicon 93 -1361 93 -1361 0 1
rlabel polysilicon 93 -1367 93 -1367 0 3
rlabel polysilicon 100 -1361 100 -1361 0 1
rlabel polysilicon 103 -1361 103 -1361 0 2
rlabel polysilicon 100 -1367 100 -1367 0 3
rlabel polysilicon 103 -1367 103 -1367 0 4
rlabel polysilicon 110 -1367 110 -1367 0 4
rlabel polysilicon 114 -1361 114 -1361 0 1
rlabel polysilicon 114 -1367 114 -1367 0 3
rlabel polysilicon 121 -1361 121 -1361 0 1
rlabel polysilicon 121 -1367 121 -1367 0 3
rlabel polysilicon 128 -1367 128 -1367 0 3
rlabel polysilicon 131 -1367 131 -1367 0 4
rlabel polysilicon 135 -1361 135 -1361 0 1
rlabel polysilicon 135 -1367 135 -1367 0 3
rlabel polysilicon 142 -1361 142 -1361 0 1
rlabel polysilicon 142 -1367 142 -1367 0 3
rlabel polysilicon 149 -1361 149 -1361 0 1
rlabel polysilicon 149 -1367 149 -1367 0 3
rlabel polysilicon 156 -1361 156 -1361 0 1
rlabel polysilicon 156 -1367 156 -1367 0 3
rlabel polysilicon 163 -1361 163 -1361 0 1
rlabel polysilicon 163 -1367 163 -1367 0 3
rlabel polysilicon 170 -1361 170 -1361 0 1
rlabel polysilicon 170 -1367 170 -1367 0 3
rlabel polysilicon 177 -1361 177 -1361 0 1
rlabel polysilicon 177 -1367 177 -1367 0 3
rlabel polysilicon 184 -1361 184 -1361 0 1
rlabel polysilicon 187 -1361 187 -1361 0 2
rlabel polysilicon 191 -1361 191 -1361 0 1
rlabel polysilicon 191 -1367 191 -1367 0 3
rlabel polysilicon 198 -1361 198 -1361 0 1
rlabel polysilicon 198 -1367 198 -1367 0 3
rlabel polysilicon 201 -1367 201 -1367 0 4
rlabel polysilicon 205 -1361 205 -1361 0 1
rlabel polysilicon 208 -1361 208 -1361 0 2
rlabel polysilicon 205 -1367 205 -1367 0 3
rlabel polysilicon 208 -1367 208 -1367 0 4
rlabel polysilicon 212 -1361 212 -1361 0 1
rlabel polysilicon 212 -1367 212 -1367 0 3
rlabel polysilicon 222 -1361 222 -1361 0 2
rlabel polysilicon 219 -1367 219 -1367 0 3
rlabel polysilicon 222 -1367 222 -1367 0 4
rlabel polysilicon 226 -1361 226 -1361 0 1
rlabel polysilicon 226 -1367 226 -1367 0 3
rlabel polysilicon 233 -1361 233 -1361 0 1
rlabel polysilicon 233 -1367 233 -1367 0 3
rlabel polysilicon 240 -1361 240 -1361 0 1
rlabel polysilicon 240 -1367 240 -1367 0 3
rlabel polysilicon 247 -1361 247 -1361 0 1
rlabel polysilicon 247 -1367 247 -1367 0 3
rlabel polysilicon 254 -1361 254 -1361 0 1
rlabel polysilicon 254 -1367 254 -1367 0 3
rlabel polysilicon 261 -1361 261 -1361 0 1
rlabel polysilicon 261 -1367 261 -1367 0 3
rlabel polysilicon 268 -1361 268 -1361 0 1
rlabel polysilicon 268 -1367 268 -1367 0 3
rlabel polysilicon 275 -1361 275 -1361 0 1
rlabel polysilicon 275 -1367 275 -1367 0 3
rlabel polysilicon 282 -1361 282 -1361 0 1
rlabel polysilicon 282 -1367 282 -1367 0 3
rlabel polysilicon 292 -1361 292 -1361 0 2
rlabel polysilicon 292 -1367 292 -1367 0 4
rlabel polysilicon 296 -1361 296 -1361 0 1
rlabel polysilicon 296 -1367 296 -1367 0 3
rlabel polysilicon 303 -1361 303 -1361 0 1
rlabel polysilicon 303 -1367 303 -1367 0 3
rlabel polysilicon 310 -1361 310 -1361 0 1
rlabel polysilicon 310 -1367 310 -1367 0 3
rlabel polysilicon 317 -1361 317 -1361 0 1
rlabel polysilicon 317 -1367 317 -1367 0 3
rlabel polysilicon 324 -1361 324 -1361 0 1
rlabel polysilicon 324 -1367 324 -1367 0 3
rlabel polysilicon 331 -1361 331 -1361 0 1
rlabel polysilicon 331 -1367 331 -1367 0 3
rlabel polysilicon 338 -1361 338 -1361 0 1
rlabel polysilicon 338 -1367 338 -1367 0 3
rlabel polysilicon 345 -1361 345 -1361 0 1
rlabel polysilicon 345 -1367 345 -1367 0 3
rlabel polysilicon 352 -1361 352 -1361 0 1
rlabel polysilicon 352 -1367 352 -1367 0 3
rlabel polysilicon 359 -1361 359 -1361 0 1
rlabel polysilicon 359 -1367 359 -1367 0 3
rlabel polysilicon 366 -1361 366 -1361 0 1
rlabel polysilicon 366 -1367 366 -1367 0 3
rlabel polysilicon 373 -1361 373 -1361 0 1
rlabel polysilicon 373 -1367 373 -1367 0 3
rlabel polysilicon 380 -1361 380 -1361 0 1
rlabel polysilicon 380 -1367 380 -1367 0 3
rlabel polysilicon 387 -1361 387 -1361 0 1
rlabel polysilicon 387 -1367 387 -1367 0 3
rlabel polysilicon 394 -1361 394 -1361 0 1
rlabel polysilicon 394 -1367 394 -1367 0 3
rlabel polysilicon 401 -1361 401 -1361 0 1
rlabel polysilicon 401 -1367 401 -1367 0 3
rlabel polysilicon 408 -1361 408 -1361 0 1
rlabel polysilicon 408 -1367 408 -1367 0 3
rlabel polysilicon 415 -1361 415 -1361 0 1
rlabel polysilicon 415 -1367 415 -1367 0 3
rlabel polysilicon 422 -1361 422 -1361 0 1
rlabel polysilicon 422 -1367 422 -1367 0 3
rlabel polysilicon 429 -1361 429 -1361 0 1
rlabel polysilicon 429 -1367 429 -1367 0 3
rlabel polysilicon 436 -1361 436 -1361 0 1
rlabel polysilicon 436 -1367 436 -1367 0 3
rlabel polysilicon 446 -1361 446 -1361 0 2
rlabel polysilicon 443 -1367 443 -1367 0 3
rlabel polysilicon 450 -1361 450 -1361 0 1
rlabel polysilicon 453 -1361 453 -1361 0 2
rlabel polysilicon 453 -1367 453 -1367 0 4
rlabel polysilicon 457 -1361 457 -1361 0 1
rlabel polysilicon 457 -1367 457 -1367 0 3
rlabel polysilicon 464 -1361 464 -1361 0 1
rlabel polysilicon 464 -1367 464 -1367 0 3
rlabel polysilicon 471 -1361 471 -1361 0 1
rlabel polysilicon 471 -1367 471 -1367 0 3
rlabel polysilicon 478 -1361 478 -1361 0 1
rlabel polysilicon 478 -1367 478 -1367 0 3
rlabel polysilicon 485 -1361 485 -1361 0 1
rlabel polysilicon 485 -1367 485 -1367 0 3
rlabel polysilicon 492 -1361 492 -1361 0 1
rlabel polysilicon 492 -1367 492 -1367 0 3
rlabel polysilicon 499 -1361 499 -1361 0 1
rlabel polysilicon 499 -1367 499 -1367 0 3
rlabel polysilicon 506 -1361 506 -1361 0 1
rlabel polysilicon 506 -1367 506 -1367 0 3
rlabel polysilicon 513 -1361 513 -1361 0 1
rlabel polysilicon 513 -1367 513 -1367 0 3
rlabel polysilicon 520 -1361 520 -1361 0 1
rlabel polysilicon 520 -1367 520 -1367 0 3
rlabel polysilicon 527 -1361 527 -1361 0 1
rlabel polysilicon 527 -1367 527 -1367 0 3
rlabel polysilicon 534 -1361 534 -1361 0 1
rlabel polysilicon 534 -1367 534 -1367 0 3
rlabel polysilicon 541 -1361 541 -1361 0 1
rlabel polysilicon 541 -1367 541 -1367 0 3
rlabel polysilicon 548 -1361 548 -1361 0 1
rlabel polysilicon 551 -1361 551 -1361 0 2
rlabel polysilicon 548 -1367 548 -1367 0 3
rlabel polysilicon 551 -1367 551 -1367 0 4
rlabel polysilicon 555 -1361 555 -1361 0 1
rlabel polysilicon 558 -1361 558 -1361 0 2
rlabel polysilicon 555 -1367 555 -1367 0 3
rlabel polysilicon 558 -1367 558 -1367 0 4
rlabel polysilicon 562 -1361 562 -1361 0 1
rlabel polysilicon 565 -1361 565 -1361 0 2
rlabel polysilicon 562 -1367 562 -1367 0 3
rlabel polysilicon 569 -1361 569 -1361 0 1
rlabel polysilicon 572 -1361 572 -1361 0 2
rlabel polysilicon 569 -1367 569 -1367 0 3
rlabel polysilicon 572 -1367 572 -1367 0 4
rlabel polysilicon 576 -1361 576 -1361 0 1
rlabel polysilicon 576 -1367 576 -1367 0 3
rlabel polysilicon 583 -1361 583 -1361 0 1
rlabel polysilicon 583 -1367 583 -1367 0 3
rlabel polysilicon 590 -1361 590 -1361 0 1
rlabel polysilicon 590 -1367 590 -1367 0 3
rlabel polysilicon 597 -1361 597 -1361 0 1
rlabel polysilicon 600 -1361 600 -1361 0 2
rlabel polysilicon 597 -1367 597 -1367 0 3
rlabel polysilicon 604 -1361 604 -1361 0 1
rlabel polysilicon 604 -1367 604 -1367 0 3
rlabel polysilicon 611 -1361 611 -1361 0 1
rlabel polysilicon 611 -1367 611 -1367 0 3
rlabel polysilicon 618 -1361 618 -1361 0 1
rlabel polysilicon 618 -1367 618 -1367 0 3
rlabel polysilicon 625 -1361 625 -1361 0 1
rlabel polysilicon 625 -1367 625 -1367 0 3
rlabel polysilicon 632 -1361 632 -1361 0 1
rlabel polysilicon 632 -1367 632 -1367 0 3
rlabel polysilicon 639 -1361 639 -1361 0 1
rlabel polysilicon 639 -1367 639 -1367 0 3
rlabel polysilicon 646 -1361 646 -1361 0 1
rlabel polysilicon 646 -1367 646 -1367 0 3
rlabel polysilicon 653 -1361 653 -1361 0 1
rlabel polysilicon 653 -1367 653 -1367 0 3
rlabel polysilicon 660 -1361 660 -1361 0 1
rlabel polysilicon 660 -1367 660 -1367 0 3
rlabel polysilicon 667 -1361 667 -1361 0 1
rlabel polysilicon 667 -1367 667 -1367 0 3
rlabel polysilicon 674 -1361 674 -1361 0 1
rlabel polysilicon 674 -1367 674 -1367 0 3
rlabel polysilicon 681 -1361 681 -1361 0 1
rlabel polysilicon 681 -1367 681 -1367 0 3
rlabel polysilicon 688 -1361 688 -1361 0 1
rlabel polysilicon 688 -1367 688 -1367 0 3
rlabel polysilicon 695 -1361 695 -1361 0 1
rlabel polysilicon 695 -1367 695 -1367 0 3
rlabel polysilicon 702 -1361 702 -1361 0 1
rlabel polysilicon 702 -1367 702 -1367 0 3
rlabel polysilicon 709 -1361 709 -1361 0 1
rlabel polysilicon 709 -1367 709 -1367 0 3
rlabel polysilicon 716 -1361 716 -1361 0 1
rlabel polysilicon 716 -1367 716 -1367 0 3
rlabel polysilicon 723 -1361 723 -1361 0 1
rlabel polysilicon 723 -1367 723 -1367 0 3
rlabel polysilicon 730 -1361 730 -1361 0 1
rlabel polysilicon 730 -1367 730 -1367 0 3
rlabel polysilicon 737 -1361 737 -1361 0 1
rlabel polysilicon 740 -1361 740 -1361 0 2
rlabel polysilicon 737 -1367 737 -1367 0 3
rlabel polysilicon 740 -1367 740 -1367 0 4
rlabel polysilicon 744 -1361 744 -1361 0 1
rlabel polysilicon 744 -1367 744 -1367 0 3
rlabel polysilicon 751 -1361 751 -1361 0 1
rlabel polysilicon 754 -1361 754 -1361 0 2
rlabel polysilicon 751 -1367 751 -1367 0 3
rlabel polysilicon 754 -1367 754 -1367 0 4
rlabel polysilicon 758 -1361 758 -1361 0 1
rlabel polysilicon 758 -1367 758 -1367 0 3
rlabel polysilicon 765 -1361 765 -1361 0 1
rlabel polysilicon 765 -1367 765 -1367 0 3
rlabel polysilicon 772 -1361 772 -1361 0 1
rlabel polysilicon 772 -1367 772 -1367 0 3
rlabel polysilicon 779 -1361 779 -1361 0 1
rlabel polysilicon 779 -1367 779 -1367 0 3
rlabel polysilicon 786 -1361 786 -1361 0 1
rlabel polysilicon 789 -1361 789 -1361 0 2
rlabel polysilicon 789 -1367 789 -1367 0 4
rlabel polysilicon 793 -1361 793 -1361 0 1
rlabel polysilicon 793 -1367 793 -1367 0 3
rlabel polysilicon 800 -1361 800 -1361 0 1
rlabel polysilicon 800 -1367 800 -1367 0 3
rlabel polysilicon 807 -1361 807 -1361 0 1
rlabel polysilicon 807 -1367 807 -1367 0 3
rlabel polysilicon 814 -1361 814 -1361 0 1
rlabel polysilicon 817 -1361 817 -1361 0 2
rlabel polysilicon 814 -1367 814 -1367 0 3
rlabel polysilicon 817 -1367 817 -1367 0 4
rlabel polysilicon 821 -1361 821 -1361 0 1
rlabel polysilicon 824 -1361 824 -1361 0 2
rlabel polysilicon 824 -1367 824 -1367 0 4
rlabel polysilicon 831 -1361 831 -1361 0 2
rlabel polysilicon 828 -1367 828 -1367 0 3
rlabel polysilicon 835 -1361 835 -1361 0 1
rlabel polysilicon 835 -1367 835 -1367 0 3
rlabel polysilicon 842 -1361 842 -1361 0 1
rlabel polysilicon 842 -1367 842 -1367 0 3
rlabel polysilicon 849 -1361 849 -1361 0 1
rlabel polysilicon 852 -1361 852 -1361 0 2
rlabel polysilicon 849 -1367 849 -1367 0 3
rlabel polysilicon 852 -1367 852 -1367 0 4
rlabel polysilicon 856 -1361 856 -1361 0 1
rlabel polysilicon 856 -1367 856 -1367 0 3
rlabel polysilicon 863 -1361 863 -1361 0 1
rlabel polysilicon 863 -1367 863 -1367 0 3
rlabel polysilicon 870 -1361 870 -1361 0 1
rlabel polysilicon 870 -1367 870 -1367 0 3
rlabel polysilicon 877 -1361 877 -1361 0 1
rlabel polysilicon 877 -1367 877 -1367 0 3
rlabel polysilicon 884 -1361 884 -1361 0 1
rlabel polysilicon 884 -1367 884 -1367 0 3
rlabel polysilicon 891 -1361 891 -1361 0 1
rlabel polysilicon 891 -1367 891 -1367 0 3
rlabel polysilicon 898 -1361 898 -1361 0 1
rlabel polysilicon 898 -1367 898 -1367 0 3
rlabel polysilicon 905 -1361 905 -1361 0 1
rlabel polysilicon 905 -1367 905 -1367 0 3
rlabel polysilicon 912 -1361 912 -1361 0 1
rlabel polysilicon 912 -1367 912 -1367 0 3
rlabel polysilicon 922 -1361 922 -1361 0 2
rlabel polysilicon 919 -1367 919 -1367 0 3
rlabel polysilicon 922 -1367 922 -1367 0 4
rlabel polysilicon 926 -1361 926 -1361 0 1
rlabel polysilicon 926 -1367 926 -1367 0 3
rlabel polysilicon 933 -1361 933 -1361 0 1
rlabel polysilicon 936 -1361 936 -1361 0 2
rlabel polysilicon 933 -1367 933 -1367 0 3
rlabel polysilicon 936 -1367 936 -1367 0 4
rlabel polysilicon 940 -1361 940 -1361 0 1
rlabel polysilicon 940 -1367 940 -1367 0 3
rlabel polysilicon 947 -1361 947 -1361 0 1
rlabel polysilicon 950 -1361 950 -1361 0 2
rlabel polysilicon 947 -1367 947 -1367 0 3
rlabel polysilicon 950 -1367 950 -1367 0 4
rlabel polysilicon 954 -1361 954 -1361 0 1
rlabel polysilicon 954 -1367 954 -1367 0 3
rlabel polysilicon 961 -1361 961 -1361 0 1
rlabel polysilicon 961 -1367 961 -1367 0 3
rlabel polysilicon 968 -1361 968 -1361 0 1
rlabel polysilicon 968 -1367 968 -1367 0 3
rlabel polysilicon 975 -1361 975 -1361 0 1
rlabel polysilicon 975 -1367 975 -1367 0 3
rlabel polysilicon 982 -1361 982 -1361 0 1
rlabel polysilicon 982 -1367 982 -1367 0 3
rlabel polysilicon 985 -1367 985 -1367 0 4
rlabel polysilicon 989 -1361 989 -1361 0 1
rlabel polysilicon 989 -1367 989 -1367 0 3
rlabel polysilicon 996 -1361 996 -1361 0 1
rlabel polysilicon 996 -1367 996 -1367 0 3
rlabel polysilicon 1003 -1361 1003 -1361 0 1
rlabel polysilicon 1006 -1361 1006 -1361 0 2
rlabel polysilicon 1006 -1367 1006 -1367 0 4
rlabel polysilicon 1010 -1361 1010 -1361 0 1
rlabel polysilicon 1010 -1367 1010 -1367 0 3
rlabel polysilicon 1020 -1361 1020 -1361 0 2
rlabel polysilicon 1017 -1367 1017 -1367 0 3
rlabel polysilicon 1020 -1367 1020 -1367 0 4
rlabel polysilicon 1024 -1361 1024 -1361 0 1
rlabel polysilicon 1024 -1367 1024 -1367 0 3
rlabel polysilicon 1031 -1361 1031 -1361 0 1
rlabel polysilicon 1031 -1367 1031 -1367 0 3
rlabel polysilicon 1038 -1361 1038 -1361 0 1
rlabel polysilicon 1038 -1367 1038 -1367 0 3
rlabel polysilicon 1045 -1361 1045 -1361 0 1
rlabel polysilicon 1045 -1367 1045 -1367 0 3
rlabel polysilicon 1052 -1361 1052 -1361 0 1
rlabel polysilicon 1052 -1367 1052 -1367 0 3
rlabel polysilicon 1059 -1361 1059 -1361 0 1
rlabel polysilicon 1059 -1367 1059 -1367 0 3
rlabel polysilicon 1066 -1361 1066 -1361 0 1
rlabel polysilicon 1066 -1367 1066 -1367 0 3
rlabel polysilicon 1073 -1361 1073 -1361 0 1
rlabel polysilicon 1073 -1367 1073 -1367 0 3
rlabel polysilicon 1080 -1361 1080 -1361 0 1
rlabel polysilicon 1080 -1367 1080 -1367 0 3
rlabel polysilicon 1087 -1361 1087 -1361 0 1
rlabel polysilicon 1087 -1367 1087 -1367 0 3
rlabel polysilicon 1094 -1361 1094 -1361 0 1
rlabel polysilicon 1094 -1367 1094 -1367 0 3
rlabel polysilicon 1101 -1361 1101 -1361 0 1
rlabel polysilicon 1104 -1361 1104 -1361 0 2
rlabel polysilicon 1101 -1367 1101 -1367 0 3
rlabel polysilicon 1104 -1367 1104 -1367 0 4
rlabel polysilicon 1108 -1361 1108 -1361 0 1
rlabel polysilicon 1108 -1367 1108 -1367 0 3
rlabel polysilicon 1115 -1361 1115 -1361 0 1
rlabel polysilicon 1115 -1367 1115 -1367 0 3
rlabel polysilicon 1122 -1361 1122 -1361 0 1
rlabel polysilicon 1122 -1367 1122 -1367 0 3
rlabel polysilicon 1129 -1361 1129 -1361 0 1
rlabel polysilicon 1129 -1367 1129 -1367 0 3
rlabel polysilicon 1136 -1361 1136 -1361 0 1
rlabel polysilicon 1136 -1367 1136 -1367 0 3
rlabel polysilicon 1146 -1361 1146 -1361 0 2
rlabel polysilicon 1143 -1367 1143 -1367 0 3
rlabel polysilicon 1146 -1367 1146 -1367 0 4
rlabel polysilicon 1150 -1361 1150 -1361 0 1
rlabel polysilicon 1150 -1367 1150 -1367 0 3
rlabel polysilicon 1157 -1361 1157 -1361 0 1
rlabel polysilicon 1157 -1367 1157 -1367 0 3
rlabel polysilicon 1164 -1361 1164 -1361 0 1
rlabel polysilicon 1164 -1367 1164 -1367 0 3
rlabel polysilicon 1171 -1361 1171 -1361 0 1
rlabel polysilicon 1171 -1367 1171 -1367 0 3
rlabel polysilicon 1178 -1361 1178 -1361 0 1
rlabel polysilicon 1178 -1367 1178 -1367 0 3
rlabel polysilicon 1185 -1361 1185 -1361 0 1
rlabel polysilicon 1185 -1367 1185 -1367 0 3
rlabel polysilicon 1192 -1361 1192 -1361 0 1
rlabel polysilicon 1192 -1367 1192 -1367 0 3
rlabel polysilicon 1199 -1361 1199 -1361 0 1
rlabel polysilicon 1202 -1361 1202 -1361 0 2
rlabel polysilicon 1202 -1367 1202 -1367 0 4
rlabel polysilicon 1206 -1361 1206 -1361 0 1
rlabel polysilicon 1206 -1367 1206 -1367 0 3
rlabel polysilicon 1213 -1361 1213 -1361 0 1
rlabel polysilicon 1213 -1367 1213 -1367 0 3
rlabel polysilicon 1216 -1367 1216 -1367 0 4
rlabel polysilicon 1220 -1361 1220 -1361 0 1
rlabel polysilicon 1220 -1367 1220 -1367 0 3
rlabel polysilicon 1227 -1361 1227 -1361 0 1
rlabel polysilicon 1227 -1367 1227 -1367 0 3
rlabel polysilicon 1234 -1361 1234 -1361 0 1
rlabel polysilicon 1234 -1367 1234 -1367 0 3
rlabel polysilicon 1241 -1361 1241 -1361 0 1
rlabel polysilicon 1241 -1367 1241 -1367 0 3
rlabel polysilicon 1248 -1361 1248 -1361 0 1
rlabel polysilicon 1248 -1367 1248 -1367 0 3
rlabel polysilicon 1255 -1361 1255 -1361 0 1
rlabel polysilicon 1255 -1367 1255 -1367 0 3
rlabel polysilicon 1262 -1361 1262 -1361 0 1
rlabel polysilicon 1262 -1367 1262 -1367 0 3
rlabel polysilicon 1269 -1361 1269 -1361 0 1
rlabel polysilicon 1269 -1367 1269 -1367 0 3
rlabel polysilicon 1276 -1361 1276 -1361 0 1
rlabel polysilicon 1276 -1367 1276 -1367 0 3
rlabel polysilicon 1283 -1361 1283 -1361 0 1
rlabel polysilicon 1283 -1367 1283 -1367 0 3
rlabel polysilicon 1290 -1361 1290 -1361 0 1
rlabel polysilicon 1290 -1367 1290 -1367 0 3
rlabel polysilicon 1297 -1361 1297 -1361 0 1
rlabel polysilicon 1297 -1367 1297 -1367 0 3
rlabel polysilicon 1304 -1367 1304 -1367 0 3
rlabel polysilicon 1311 -1361 1311 -1361 0 1
rlabel polysilicon 1314 -1361 1314 -1361 0 2
rlabel polysilicon 1311 -1367 1311 -1367 0 3
rlabel polysilicon 1318 -1361 1318 -1361 0 1
rlabel polysilicon 1318 -1367 1318 -1367 0 3
rlabel polysilicon 1325 -1361 1325 -1361 0 1
rlabel polysilicon 1325 -1367 1325 -1367 0 3
rlabel polysilicon 1332 -1361 1332 -1361 0 1
rlabel polysilicon 1332 -1367 1332 -1367 0 3
rlabel polysilicon 1339 -1361 1339 -1361 0 1
rlabel polysilicon 1339 -1367 1339 -1367 0 3
rlabel polysilicon 1346 -1361 1346 -1361 0 1
rlabel polysilicon 1346 -1367 1346 -1367 0 3
rlabel polysilicon 1353 -1361 1353 -1361 0 1
rlabel polysilicon 1353 -1367 1353 -1367 0 3
rlabel polysilicon 1360 -1361 1360 -1361 0 1
rlabel polysilicon 1360 -1367 1360 -1367 0 3
rlabel polysilicon 1367 -1361 1367 -1361 0 1
rlabel polysilicon 1367 -1367 1367 -1367 0 3
rlabel polysilicon 1374 -1361 1374 -1361 0 1
rlabel polysilicon 1374 -1367 1374 -1367 0 3
rlabel polysilicon 1381 -1361 1381 -1361 0 1
rlabel polysilicon 1381 -1367 1381 -1367 0 3
rlabel polysilicon 1388 -1361 1388 -1361 0 1
rlabel polysilicon 1388 -1367 1388 -1367 0 3
rlabel polysilicon 1395 -1361 1395 -1361 0 1
rlabel polysilicon 1395 -1367 1395 -1367 0 3
rlabel polysilicon 1402 -1361 1402 -1361 0 1
rlabel polysilicon 1402 -1367 1402 -1367 0 3
rlabel polysilicon 1409 -1361 1409 -1361 0 1
rlabel polysilicon 1409 -1367 1409 -1367 0 3
rlabel polysilicon 1416 -1361 1416 -1361 0 1
rlabel polysilicon 1416 -1367 1416 -1367 0 3
rlabel polysilicon 1423 -1361 1423 -1361 0 1
rlabel polysilicon 1423 -1367 1423 -1367 0 3
rlabel polysilicon 1430 -1361 1430 -1361 0 1
rlabel polysilicon 1430 -1367 1430 -1367 0 3
rlabel polysilicon 1437 -1361 1437 -1361 0 1
rlabel polysilicon 1437 -1367 1437 -1367 0 3
rlabel polysilicon 1444 -1361 1444 -1361 0 1
rlabel polysilicon 1444 -1367 1444 -1367 0 3
rlabel polysilicon 1451 -1361 1451 -1361 0 1
rlabel polysilicon 1451 -1367 1451 -1367 0 3
rlabel polysilicon 1458 -1361 1458 -1361 0 1
rlabel polysilicon 1458 -1367 1458 -1367 0 3
rlabel polysilicon 1465 -1361 1465 -1361 0 1
rlabel polysilicon 1465 -1367 1465 -1367 0 3
rlabel polysilicon 1472 -1361 1472 -1361 0 1
rlabel polysilicon 1472 -1367 1472 -1367 0 3
rlabel polysilicon 1479 -1361 1479 -1361 0 1
rlabel polysilicon 1479 -1367 1479 -1367 0 3
rlabel polysilicon 1486 -1361 1486 -1361 0 1
rlabel polysilicon 1486 -1367 1486 -1367 0 3
rlabel polysilicon 1493 -1361 1493 -1361 0 1
rlabel polysilicon 1493 -1367 1493 -1367 0 3
rlabel polysilicon 1500 -1361 1500 -1361 0 1
rlabel polysilicon 1500 -1367 1500 -1367 0 3
rlabel polysilicon 1507 -1361 1507 -1361 0 1
rlabel polysilicon 1507 -1367 1507 -1367 0 3
rlabel polysilicon 1514 -1361 1514 -1361 0 1
rlabel polysilicon 1514 -1367 1514 -1367 0 3
rlabel polysilicon 1521 -1361 1521 -1361 0 1
rlabel polysilicon 1521 -1367 1521 -1367 0 3
rlabel polysilicon 1528 -1361 1528 -1361 0 1
rlabel polysilicon 1528 -1367 1528 -1367 0 3
rlabel polysilicon 1535 -1361 1535 -1361 0 1
rlabel polysilicon 1535 -1367 1535 -1367 0 3
rlabel polysilicon 1542 -1361 1542 -1361 0 1
rlabel polysilicon 1542 -1367 1542 -1367 0 3
rlabel polysilicon 1549 -1361 1549 -1361 0 1
rlabel polysilicon 1549 -1367 1549 -1367 0 3
rlabel polysilicon 1556 -1361 1556 -1361 0 1
rlabel polysilicon 1556 -1367 1556 -1367 0 3
rlabel polysilicon 1563 -1361 1563 -1361 0 1
rlabel polysilicon 1563 -1367 1563 -1367 0 3
rlabel polysilicon 1570 -1361 1570 -1361 0 1
rlabel polysilicon 1570 -1367 1570 -1367 0 3
rlabel polysilicon 1577 -1361 1577 -1361 0 1
rlabel polysilicon 1577 -1367 1577 -1367 0 3
rlabel polysilicon 1584 -1361 1584 -1361 0 1
rlabel polysilicon 1584 -1367 1584 -1367 0 3
rlabel polysilicon 1591 -1361 1591 -1361 0 1
rlabel polysilicon 1591 -1367 1591 -1367 0 3
rlabel polysilicon 1598 -1361 1598 -1361 0 1
rlabel polysilicon 1598 -1367 1598 -1367 0 3
rlabel polysilicon 1605 -1361 1605 -1361 0 1
rlabel polysilicon 1605 -1367 1605 -1367 0 3
rlabel polysilicon 1612 -1361 1612 -1361 0 1
rlabel polysilicon 1612 -1367 1612 -1367 0 3
rlabel polysilicon 1619 -1361 1619 -1361 0 1
rlabel polysilicon 1619 -1367 1619 -1367 0 3
rlabel polysilicon 1626 -1361 1626 -1361 0 1
rlabel polysilicon 1626 -1367 1626 -1367 0 3
rlabel polysilicon 1633 -1361 1633 -1361 0 1
rlabel polysilicon 1633 -1367 1633 -1367 0 3
rlabel polysilicon 1640 -1361 1640 -1361 0 1
rlabel polysilicon 1640 -1367 1640 -1367 0 3
rlabel polysilicon 1647 -1361 1647 -1361 0 1
rlabel polysilicon 1647 -1367 1647 -1367 0 3
rlabel polysilicon 1654 -1361 1654 -1361 0 1
rlabel polysilicon 1654 -1367 1654 -1367 0 3
rlabel polysilicon 1661 -1361 1661 -1361 0 1
rlabel polysilicon 1661 -1367 1661 -1367 0 3
rlabel polysilicon 1668 -1361 1668 -1361 0 1
rlabel polysilicon 1668 -1367 1668 -1367 0 3
rlabel polysilicon 1675 -1361 1675 -1361 0 1
rlabel polysilicon 1675 -1367 1675 -1367 0 3
rlabel polysilicon 1682 -1361 1682 -1361 0 1
rlabel polysilicon 1682 -1367 1682 -1367 0 3
rlabel polysilicon 1689 -1361 1689 -1361 0 1
rlabel polysilicon 1689 -1367 1689 -1367 0 3
rlabel polysilicon 1696 -1361 1696 -1361 0 1
rlabel polysilicon 1696 -1367 1696 -1367 0 3
rlabel polysilicon 1703 -1361 1703 -1361 0 1
rlabel polysilicon 1703 -1367 1703 -1367 0 3
rlabel polysilicon 1710 -1361 1710 -1361 0 1
rlabel polysilicon 1710 -1367 1710 -1367 0 3
rlabel polysilicon 1717 -1361 1717 -1361 0 1
rlabel polysilicon 1717 -1367 1717 -1367 0 3
rlabel polysilicon 1724 -1361 1724 -1361 0 1
rlabel polysilicon 1724 -1367 1724 -1367 0 3
rlabel polysilicon 1731 -1361 1731 -1361 0 1
rlabel polysilicon 1731 -1367 1731 -1367 0 3
rlabel polysilicon 1738 -1361 1738 -1361 0 1
rlabel polysilicon 1738 -1367 1738 -1367 0 3
rlabel polysilicon 1745 -1361 1745 -1361 0 1
rlabel polysilicon 1745 -1367 1745 -1367 0 3
rlabel polysilicon 1752 -1361 1752 -1361 0 1
rlabel polysilicon 1752 -1367 1752 -1367 0 3
rlabel polysilicon 23 -1502 23 -1502 0 1
rlabel polysilicon 23 -1508 23 -1508 0 3
rlabel polysilicon 30 -1502 30 -1502 0 1
rlabel polysilicon 30 -1508 30 -1508 0 3
rlabel polysilicon 37 -1502 37 -1502 0 1
rlabel polysilicon 37 -1508 37 -1508 0 3
rlabel polysilicon 44 -1502 44 -1502 0 1
rlabel polysilicon 44 -1508 44 -1508 0 3
rlabel polysilicon 51 -1502 51 -1502 0 1
rlabel polysilicon 51 -1508 51 -1508 0 3
rlabel polysilicon 58 -1502 58 -1502 0 1
rlabel polysilicon 58 -1508 58 -1508 0 3
rlabel polysilicon 65 -1508 65 -1508 0 3
rlabel polysilicon 68 -1508 68 -1508 0 4
rlabel polysilicon 72 -1502 72 -1502 0 1
rlabel polysilicon 72 -1508 72 -1508 0 3
rlabel polysilicon 79 -1502 79 -1502 0 1
rlabel polysilicon 79 -1508 79 -1508 0 3
rlabel polysilicon 86 -1502 86 -1502 0 1
rlabel polysilicon 86 -1508 86 -1508 0 3
rlabel polysilicon 93 -1502 93 -1502 0 1
rlabel polysilicon 93 -1508 93 -1508 0 3
rlabel polysilicon 100 -1502 100 -1502 0 1
rlabel polysilicon 100 -1508 100 -1508 0 3
rlabel polysilicon 107 -1502 107 -1502 0 1
rlabel polysilicon 107 -1508 107 -1508 0 3
rlabel polysilicon 114 -1502 114 -1502 0 1
rlabel polysilicon 114 -1508 114 -1508 0 3
rlabel polysilicon 124 -1502 124 -1502 0 2
rlabel polysilicon 121 -1508 121 -1508 0 3
rlabel polysilicon 124 -1508 124 -1508 0 4
rlabel polysilicon 128 -1502 128 -1502 0 1
rlabel polysilicon 131 -1502 131 -1502 0 2
rlabel polysilicon 128 -1508 128 -1508 0 3
rlabel polysilicon 131 -1508 131 -1508 0 4
rlabel polysilicon 135 -1502 135 -1502 0 1
rlabel polysilicon 135 -1508 135 -1508 0 3
rlabel polysilicon 142 -1502 142 -1502 0 1
rlabel polysilicon 142 -1508 142 -1508 0 3
rlabel polysilicon 149 -1502 149 -1502 0 1
rlabel polysilicon 149 -1508 149 -1508 0 3
rlabel polysilicon 156 -1502 156 -1502 0 1
rlabel polysilicon 159 -1502 159 -1502 0 2
rlabel polysilicon 156 -1508 156 -1508 0 3
rlabel polysilicon 159 -1508 159 -1508 0 4
rlabel polysilicon 163 -1502 163 -1502 0 1
rlabel polysilicon 163 -1508 163 -1508 0 3
rlabel polysilicon 170 -1502 170 -1502 0 1
rlabel polysilicon 170 -1508 170 -1508 0 3
rlabel polysilicon 177 -1502 177 -1502 0 1
rlabel polysilicon 177 -1508 177 -1508 0 3
rlabel polysilicon 184 -1502 184 -1502 0 1
rlabel polysilicon 187 -1502 187 -1502 0 2
rlabel polysilicon 184 -1508 184 -1508 0 3
rlabel polysilicon 191 -1502 191 -1502 0 1
rlabel polysilicon 194 -1502 194 -1502 0 2
rlabel polysilicon 191 -1508 191 -1508 0 3
rlabel polysilicon 194 -1508 194 -1508 0 4
rlabel polysilicon 198 -1502 198 -1502 0 1
rlabel polysilicon 198 -1508 198 -1508 0 3
rlabel polysilicon 205 -1502 205 -1502 0 1
rlabel polysilicon 205 -1508 205 -1508 0 3
rlabel polysilicon 212 -1502 212 -1502 0 1
rlabel polysilicon 215 -1502 215 -1502 0 2
rlabel polysilicon 212 -1508 212 -1508 0 3
rlabel polysilicon 215 -1508 215 -1508 0 4
rlabel polysilicon 219 -1502 219 -1502 0 1
rlabel polysilicon 219 -1508 219 -1508 0 3
rlabel polysilicon 226 -1502 226 -1502 0 1
rlabel polysilicon 229 -1502 229 -1502 0 2
rlabel polysilicon 226 -1508 226 -1508 0 3
rlabel polysilicon 229 -1508 229 -1508 0 4
rlabel polysilicon 233 -1502 233 -1502 0 1
rlabel polysilicon 233 -1508 233 -1508 0 3
rlabel polysilicon 240 -1502 240 -1502 0 1
rlabel polysilicon 240 -1508 240 -1508 0 3
rlabel polysilicon 247 -1502 247 -1502 0 1
rlabel polysilicon 247 -1508 247 -1508 0 3
rlabel polysilicon 254 -1502 254 -1502 0 1
rlabel polysilicon 257 -1502 257 -1502 0 2
rlabel polysilicon 254 -1508 254 -1508 0 3
rlabel polysilicon 261 -1502 261 -1502 0 1
rlabel polysilicon 261 -1508 261 -1508 0 3
rlabel polysilicon 268 -1502 268 -1502 0 1
rlabel polysilicon 268 -1508 268 -1508 0 3
rlabel polysilicon 275 -1502 275 -1502 0 1
rlabel polysilicon 275 -1508 275 -1508 0 3
rlabel polysilicon 282 -1502 282 -1502 0 1
rlabel polysilicon 282 -1508 282 -1508 0 3
rlabel polysilicon 289 -1502 289 -1502 0 1
rlabel polysilicon 289 -1508 289 -1508 0 3
rlabel polysilicon 296 -1502 296 -1502 0 1
rlabel polysilicon 296 -1508 296 -1508 0 3
rlabel polysilicon 303 -1502 303 -1502 0 1
rlabel polysilicon 303 -1508 303 -1508 0 3
rlabel polysilicon 310 -1502 310 -1502 0 1
rlabel polysilicon 310 -1508 310 -1508 0 3
rlabel polysilicon 320 -1508 320 -1508 0 4
rlabel polysilicon 324 -1502 324 -1502 0 1
rlabel polysilicon 324 -1508 324 -1508 0 3
rlabel polysilicon 331 -1502 331 -1502 0 1
rlabel polysilicon 331 -1508 331 -1508 0 3
rlabel polysilicon 338 -1502 338 -1502 0 1
rlabel polysilicon 338 -1508 338 -1508 0 3
rlabel polysilicon 345 -1502 345 -1502 0 1
rlabel polysilicon 345 -1508 345 -1508 0 3
rlabel polysilicon 352 -1502 352 -1502 0 1
rlabel polysilicon 352 -1508 352 -1508 0 3
rlabel polysilicon 359 -1502 359 -1502 0 1
rlabel polysilicon 359 -1508 359 -1508 0 3
rlabel polysilicon 366 -1502 366 -1502 0 1
rlabel polysilicon 366 -1508 366 -1508 0 3
rlabel polysilicon 373 -1502 373 -1502 0 1
rlabel polysilicon 373 -1508 373 -1508 0 3
rlabel polysilicon 380 -1502 380 -1502 0 1
rlabel polysilicon 380 -1508 380 -1508 0 3
rlabel polysilicon 387 -1502 387 -1502 0 1
rlabel polysilicon 387 -1508 387 -1508 0 3
rlabel polysilicon 394 -1502 394 -1502 0 1
rlabel polysilicon 394 -1508 394 -1508 0 3
rlabel polysilicon 401 -1502 401 -1502 0 1
rlabel polysilicon 401 -1508 401 -1508 0 3
rlabel polysilicon 408 -1502 408 -1502 0 1
rlabel polysilicon 408 -1508 408 -1508 0 3
rlabel polysilicon 415 -1502 415 -1502 0 1
rlabel polysilicon 415 -1508 415 -1508 0 3
rlabel polysilicon 418 -1508 418 -1508 0 4
rlabel polysilicon 422 -1502 422 -1502 0 1
rlabel polysilicon 422 -1508 422 -1508 0 3
rlabel polysilicon 429 -1502 429 -1502 0 1
rlabel polysilicon 429 -1508 429 -1508 0 3
rlabel polysilicon 436 -1502 436 -1502 0 1
rlabel polysilicon 436 -1508 436 -1508 0 3
rlabel polysilicon 443 -1502 443 -1502 0 1
rlabel polysilicon 443 -1508 443 -1508 0 3
rlabel polysilicon 450 -1502 450 -1502 0 1
rlabel polysilicon 450 -1508 450 -1508 0 3
rlabel polysilicon 457 -1502 457 -1502 0 1
rlabel polysilicon 460 -1502 460 -1502 0 2
rlabel polysilicon 457 -1508 457 -1508 0 3
rlabel polysilicon 460 -1508 460 -1508 0 4
rlabel polysilicon 464 -1502 464 -1502 0 1
rlabel polysilicon 464 -1508 464 -1508 0 3
rlabel polysilicon 471 -1502 471 -1502 0 1
rlabel polysilicon 471 -1508 471 -1508 0 3
rlabel polysilicon 478 -1502 478 -1502 0 1
rlabel polysilicon 481 -1502 481 -1502 0 2
rlabel polysilicon 478 -1508 478 -1508 0 3
rlabel polysilicon 481 -1508 481 -1508 0 4
rlabel polysilicon 485 -1502 485 -1502 0 1
rlabel polysilicon 492 -1502 492 -1502 0 1
rlabel polysilicon 492 -1508 492 -1508 0 3
rlabel polysilicon 499 -1502 499 -1502 0 1
rlabel polysilicon 499 -1508 499 -1508 0 3
rlabel polysilicon 506 -1502 506 -1502 0 1
rlabel polysilicon 506 -1508 506 -1508 0 3
rlabel polysilicon 513 -1502 513 -1502 0 1
rlabel polysilicon 516 -1502 516 -1502 0 2
rlabel polysilicon 513 -1508 513 -1508 0 3
rlabel polysilicon 520 -1502 520 -1502 0 1
rlabel polysilicon 520 -1508 520 -1508 0 3
rlabel polysilicon 527 -1502 527 -1502 0 1
rlabel polysilicon 527 -1508 527 -1508 0 3
rlabel polysilicon 534 -1502 534 -1502 0 1
rlabel polysilicon 534 -1508 534 -1508 0 3
rlabel polysilicon 541 -1502 541 -1502 0 1
rlabel polysilicon 541 -1508 541 -1508 0 3
rlabel polysilicon 548 -1502 548 -1502 0 1
rlabel polysilicon 548 -1508 548 -1508 0 3
rlabel polysilicon 555 -1502 555 -1502 0 1
rlabel polysilicon 555 -1508 555 -1508 0 3
rlabel polysilicon 562 -1502 562 -1502 0 1
rlabel polysilicon 562 -1508 562 -1508 0 3
rlabel polysilicon 569 -1502 569 -1502 0 1
rlabel polysilicon 569 -1508 569 -1508 0 3
rlabel polysilicon 576 -1502 576 -1502 0 1
rlabel polysilicon 576 -1508 576 -1508 0 3
rlabel polysilicon 583 -1502 583 -1502 0 1
rlabel polysilicon 583 -1508 583 -1508 0 3
rlabel polysilicon 590 -1502 590 -1502 0 1
rlabel polysilicon 590 -1508 590 -1508 0 3
rlabel polysilicon 597 -1502 597 -1502 0 1
rlabel polysilicon 597 -1508 597 -1508 0 3
rlabel polysilicon 604 -1502 604 -1502 0 1
rlabel polysilicon 604 -1508 604 -1508 0 3
rlabel polysilicon 611 -1502 611 -1502 0 1
rlabel polysilicon 611 -1508 611 -1508 0 3
rlabel polysilicon 618 -1502 618 -1502 0 1
rlabel polysilicon 618 -1508 618 -1508 0 3
rlabel polysilicon 625 -1508 625 -1508 0 3
rlabel polysilicon 628 -1508 628 -1508 0 4
rlabel polysilicon 632 -1502 632 -1502 0 1
rlabel polysilicon 632 -1508 632 -1508 0 3
rlabel polysilicon 639 -1502 639 -1502 0 1
rlabel polysilicon 639 -1508 639 -1508 0 3
rlabel polysilicon 646 -1502 646 -1502 0 1
rlabel polysilicon 646 -1508 646 -1508 0 3
rlabel polysilicon 653 -1502 653 -1502 0 1
rlabel polysilicon 653 -1508 653 -1508 0 3
rlabel polysilicon 656 -1508 656 -1508 0 4
rlabel polysilicon 660 -1502 660 -1502 0 1
rlabel polysilicon 660 -1508 660 -1508 0 3
rlabel polysilicon 670 -1502 670 -1502 0 2
rlabel polysilicon 667 -1508 667 -1508 0 3
rlabel polysilicon 670 -1508 670 -1508 0 4
rlabel polysilicon 674 -1502 674 -1502 0 1
rlabel polysilicon 674 -1508 674 -1508 0 3
rlabel polysilicon 681 -1502 681 -1502 0 1
rlabel polysilicon 681 -1508 681 -1508 0 3
rlabel polysilicon 688 -1502 688 -1502 0 1
rlabel polysilicon 688 -1508 688 -1508 0 3
rlabel polysilicon 695 -1502 695 -1502 0 1
rlabel polysilicon 695 -1508 695 -1508 0 3
rlabel polysilicon 702 -1502 702 -1502 0 1
rlabel polysilicon 702 -1508 702 -1508 0 3
rlabel polysilicon 709 -1502 709 -1502 0 1
rlabel polysilicon 709 -1508 709 -1508 0 3
rlabel polysilicon 716 -1502 716 -1502 0 1
rlabel polysilicon 719 -1502 719 -1502 0 2
rlabel polysilicon 716 -1508 716 -1508 0 3
rlabel polysilicon 726 -1502 726 -1502 0 2
rlabel polysilicon 726 -1508 726 -1508 0 4
rlabel polysilicon 730 -1502 730 -1502 0 1
rlabel polysilicon 730 -1508 730 -1508 0 3
rlabel polysilicon 737 -1502 737 -1502 0 1
rlabel polysilicon 740 -1502 740 -1502 0 2
rlabel polysilicon 737 -1508 737 -1508 0 3
rlabel polysilicon 740 -1508 740 -1508 0 4
rlabel polysilicon 744 -1502 744 -1502 0 1
rlabel polysilicon 744 -1508 744 -1508 0 3
rlabel polysilicon 751 -1502 751 -1502 0 1
rlabel polysilicon 751 -1508 751 -1508 0 3
rlabel polysilicon 758 -1502 758 -1502 0 1
rlabel polysilicon 761 -1502 761 -1502 0 2
rlabel polysilicon 758 -1508 758 -1508 0 3
rlabel polysilicon 761 -1508 761 -1508 0 4
rlabel polysilicon 765 -1502 765 -1502 0 1
rlabel polysilicon 765 -1508 765 -1508 0 3
rlabel polysilicon 772 -1502 772 -1502 0 1
rlabel polysilicon 772 -1508 772 -1508 0 3
rlabel polysilicon 779 -1502 779 -1502 0 1
rlabel polysilicon 779 -1508 779 -1508 0 3
rlabel polysilicon 786 -1502 786 -1502 0 1
rlabel polysilicon 786 -1508 786 -1508 0 3
rlabel polysilicon 789 -1508 789 -1508 0 4
rlabel polysilicon 793 -1502 793 -1502 0 1
rlabel polysilicon 793 -1508 793 -1508 0 3
rlabel polysilicon 800 -1502 800 -1502 0 1
rlabel polysilicon 800 -1508 800 -1508 0 3
rlabel polysilicon 807 -1502 807 -1502 0 1
rlabel polysilicon 807 -1508 807 -1508 0 3
rlabel polysilicon 814 -1502 814 -1502 0 1
rlabel polysilicon 814 -1508 814 -1508 0 3
rlabel polysilicon 821 -1502 821 -1502 0 1
rlabel polysilicon 824 -1502 824 -1502 0 2
rlabel polysilicon 821 -1508 821 -1508 0 3
rlabel polysilicon 824 -1508 824 -1508 0 4
rlabel polysilicon 828 -1502 828 -1502 0 1
rlabel polysilicon 831 -1502 831 -1502 0 2
rlabel polysilicon 831 -1508 831 -1508 0 4
rlabel polysilicon 835 -1502 835 -1502 0 1
rlabel polysilicon 835 -1508 835 -1508 0 3
rlabel polysilicon 842 -1502 842 -1502 0 1
rlabel polysilicon 842 -1508 842 -1508 0 3
rlabel polysilicon 849 -1502 849 -1502 0 1
rlabel polysilicon 849 -1508 849 -1508 0 3
rlabel polysilicon 856 -1502 856 -1502 0 1
rlabel polysilicon 856 -1508 856 -1508 0 3
rlabel polysilicon 863 -1502 863 -1502 0 1
rlabel polysilicon 866 -1502 866 -1502 0 2
rlabel polysilicon 863 -1508 863 -1508 0 3
rlabel polysilicon 866 -1508 866 -1508 0 4
rlabel polysilicon 870 -1502 870 -1502 0 1
rlabel polysilicon 870 -1508 870 -1508 0 3
rlabel polysilicon 877 -1502 877 -1502 0 1
rlabel polysilicon 877 -1508 877 -1508 0 3
rlabel polysilicon 884 -1502 884 -1502 0 1
rlabel polysilicon 884 -1508 884 -1508 0 3
rlabel polysilicon 891 -1502 891 -1502 0 1
rlabel polysilicon 891 -1508 891 -1508 0 3
rlabel polysilicon 898 -1502 898 -1502 0 1
rlabel polysilicon 898 -1508 898 -1508 0 3
rlabel polysilicon 905 -1502 905 -1502 0 1
rlabel polysilicon 905 -1508 905 -1508 0 3
rlabel polysilicon 912 -1502 912 -1502 0 1
rlabel polysilicon 912 -1508 912 -1508 0 3
rlabel polysilicon 919 -1502 919 -1502 0 1
rlabel polysilicon 919 -1508 919 -1508 0 3
rlabel polysilicon 926 -1502 926 -1502 0 1
rlabel polysilicon 926 -1508 926 -1508 0 3
rlabel polysilicon 933 -1502 933 -1502 0 1
rlabel polysilicon 936 -1502 936 -1502 0 2
rlabel polysilicon 933 -1508 933 -1508 0 3
rlabel polysilicon 936 -1508 936 -1508 0 4
rlabel polysilicon 940 -1502 940 -1502 0 1
rlabel polysilicon 940 -1508 940 -1508 0 3
rlabel polysilicon 947 -1502 947 -1502 0 1
rlabel polysilicon 950 -1502 950 -1502 0 2
rlabel polysilicon 947 -1508 947 -1508 0 3
rlabel polysilicon 950 -1508 950 -1508 0 4
rlabel polysilicon 954 -1502 954 -1502 0 1
rlabel polysilicon 954 -1508 954 -1508 0 3
rlabel polysilicon 961 -1502 961 -1502 0 1
rlabel polysilicon 961 -1508 961 -1508 0 3
rlabel polysilicon 968 -1502 968 -1502 0 1
rlabel polysilicon 968 -1508 968 -1508 0 3
rlabel polysilicon 978 -1502 978 -1502 0 2
rlabel polysilicon 975 -1508 975 -1508 0 3
rlabel polysilicon 978 -1508 978 -1508 0 4
rlabel polysilicon 982 -1502 982 -1502 0 1
rlabel polysilicon 982 -1508 982 -1508 0 3
rlabel polysilicon 989 -1502 989 -1502 0 1
rlabel polysilicon 989 -1508 989 -1508 0 3
rlabel polysilicon 996 -1502 996 -1502 0 1
rlabel polysilicon 996 -1508 996 -1508 0 3
rlabel polysilicon 1003 -1502 1003 -1502 0 1
rlabel polysilicon 1003 -1508 1003 -1508 0 3
rlabel polysilicon 1010 -1502 1010 -1502 0 1
rlabel polysilicon 1010 -1508 1010 -1508 0 3
rlabel polysilicon 1017 -1502 1017 -1502 0 1
rlabel polysilicon 1017 -1508 1017 -1508 0 3
rlabel polysilicon 1024 -1502 1024 -1502 0 1
rlabel polysilicon 1024 -1508 1024 -1508 0 3
rlabel polysilicon 1031 -1502 1031 -1502 0 1
rlabel polysilicon 1034 -1502 1034 -1502 0 2
rlabel polysilicon 1031 -1508 1031 -1508 0 3
rlabel polysilicon 1034 -1508 1034 -1508 0 4
rlabel polysilicon 1038 -1502 1038 -1502 0 1
rlabel polysilicon 1038 -1508 1038 -1508 0 3
rlabel polysilicon 1045 -1502 1045 -1502 0 1
rlabel polysilicon 1048 -1502 1048 -1502 0 2
rlabel polysilicon 1048 -1508 1048 -1508 0 4
rlabel polysilicon 1052 -1502 1052 -1502 0 1
rlabel polysilicon 1052 -1508 1052 -1508 0 3
rlabel polysilicon 1059 -1502 1059 -1502 0 1
rlabel polysilicon 1059 -1508 1059 -1508 0 3
rlabel polysilicon 1066 -1502 1066 -1502 0 1
rlabel polysilicon 1066 -1508 1066 -1508 0 3
rlabel polysilicon 1073 -1502 1073 -1502 0 1
rlabel polysilicon 1073 -1508 1073 -1508 0 3
rlabel polysilicon 1080 -1502 1080 -1502 0 1
rlabel polysilicon 1080 -1508 1080 -1508 0 3
rlabel polysilicon 1087 -1502 1087 -1502 0 1
rlabel polysilicon 1087 -1508 1087 -1508 0 3
rlabel polysilicon 1094 -1502 1094 -1502 0 1
rlabel polysilicon 1094 -1508 1094 -1508 0 3
rlabel polysilicon 1101 -1502 1101 -1502 0 1
rlabel polysilicon 1101 -1508 1101 -1508 0 3
rlabel polysilicon 1108 -1502 1108 -1502 0 1
rlabel polysilicon 1108 -1508 1108 -1508 0 3
rlabel polysilicon 1115 -1502 1115 -1502 0 1
rlabel polysilicon 1115 -1508 1115 -1508 0 3
rlabel polysilicon 1122 -1502 1122 -1502 0 1
rlabel polysilicon 1122 -1508 1122 -1508 0 3
rlabel polysilicon 1129 -1502 1129 -1502 0 1
rlabel polysilicon 1129 -1508 1129 -1508 0 3
rlabel polysilicon 1136 -1502 1136 -1502 0 1
rlabel polysilicon 1136 -1508 1136 -1508 0 3
rlabel polysilicon 1143 -1502 1143 -1502 0 1
rlabel polysilicon 1143 -1508 1143 -1508 0 3
rlabel polysilicon 1150 -1502 1150 -1502 0 1
rlabel polysilicon 1150 -1508 1150 -1508 0 3
rlabel polysilicon 1157 -1502 1157 -1502 0 1
rlabel polysilicon 1157 -1508 1157 -1508 0 3
rlabel polysilicon 1164 -1502 1164 -1502 0 1
rlabel polysilicon 1164 -1508 1164 -1508 0 3
rlabel polysilicon 1171 -1502 1171 -1502 0 1
rlabel polysilicon 1171 -1508 1171 -1508 0 3
rlabel polysilicon 1178 -1502 1178 -1502 0 1
rlabel polysilicon 1178 -1508 1178 -1508 0 3
rlabel polysilicon 1185 -1502 1185 -1502 0 1
rlabel polysilicon 1185 -1508 1185 -1508 0 3
rlabel polysilicon 1192 -1502 1192 -1502 0 1
rlabel polysilicon 1192 -1508 1192 -1508 0 3
rlabel polysilicon 1199 -1502 1199 -1502 0 1
rlabel polysilicon 1199 -1508 1199 -1508 0 3
rlabel polysilicon 1206 -1502 1206 -1502 0 1
rlabel polysilicon 1206 -1508 1206 -1508 0 3
rlabel polysilicon 1213 -1502 1213 -1502 0 1
rlabel polysilicon 1213 -1508 1213 -1508 0 3
rlabel polysilicon 1220 -1502 1220 -1502 0 1
rlabel polysilicon 1220 -1508 1220 -1508 0 3
rlabel polysilicon 1227 -1502 1227 -1502 0 1
rlabel polysilicon 1227 -1508 1227 -1508 0 3
rlabel polysilicon 1234 -1502 1234 -1502 0 1
rlabel polysilicon 1234 -1508 1234 -1508 0 3
rlabel polysilicon 1241 -1502 1241 -1502 0 1
rlabel polysilicon 1241 -1508 1241 -1508 0 3
rlabel polysilicon 1248 -1502 1248 -1502 0 1
rlabel polysilicon 1248 -1508 1248 -1508 0 3
rlabel polysilicon 1255 -1502 1255 -1502 0 1
rlabel polysilicon 1255 -1508 1255 -1508 0 3
rlabel polysilicon 1262 -1502 1262 -1502 0 1
rlabel polysilicon 1262 -1508 1262 -1508 0 3
rlabel polysilicon 1269 -1502 1269 -1502 0 1
rlabel polysilicon 1269 -1508 1269 -1508 0 3
rlabel polysilicon 1276 -1502 1276 -1502 0 1
rlabel polysilicon 1276 -1508 1276 -1508 0 3
rlabel polysilicon 1283 -1502 1283 -1502 0 1
rlabel polysilicon 1283 -1508 1283 -1508 0 3
rlabel polysilicon 1290 -1502 1290 -1502 0 1
rlabel polysilicon 1290 -1508 1290 -1508 0 3
rlabel polysilicon 1297 -1502 1297 -1502 0 1
rlabel polysilicon 1297 -1508 1297 -1508 0 3
rlabel polysilicon 1304 -1502 1304 -1502 0 1
rlabel polysilicon 1304 -1508 1304 -1508 0 3
rlabel polysilicon 1311 -1502 1311 -1502 0 1
rlabel polysilicon 1311 -1508 1311 -1508 0 3
rlabel polysilicon 1318 -1502 1318 -1502 0 1
rlabel polysilicon 1318 -1508 1318 -1508 0 3
rlabel polysilicon 1325 -1502 1325 -1502 0 1
rlabel polysilicon 1325 -1508 1325 -1508 0 3
rlabel polysilicon 1332 -1502 1332 -1502 0 1
rlabel polysilicon 1332 -1508 1332 -1508 0 3
rlabel polysilicon 1339 -1502 1339 -1502 0 1
rlabel polysilicon 1339 -1508 1339 -1508 0 3
rlabel polysilicon 1346 -1502 1346 -1502 0 1
rlabel polysilicon 1346 -1508 1346 -1508 0 3
rlabel polysilicon 1353 -1502 1353 -1502 0 1
rlabel polysilicon 1353 -1508 1353 -1508 0 3
rlabel polysilicon 1360 -1502 1360 -1502 0 1
rlabel polysilicon 1360 -1508 1360 -1508 0 3
rlabel polysilicon 1367 -1502 1367 -1502 0 1
rlabel polysilicon 1367 -1508 1367 -1508 0 3
rlabel polysilicon 1374 -1502 1374 -1502 0 1
rlabel polysilicon 1374 -1508 1374 -1508 0 3
rlabel polysilicon 1381 -1502 1381 -1502 0 1
rlabel polysilicon 1381 -1508 1381 -1508 0 3
rlabel polysilicon 1388 -1502 1388 -1502 0 1
rlabel polysilicon 1388 -1508 1388 -1508 0 3
rlabel polysilicon 1395 -1502 1395 -1502 0 1
rlabel polysilicon 1395 -1508 1395 -1508 0 3
rlabel polysilicon 1402 -1502 1402 -1502 0 1
rlabel polysilicon 1402 -1508 1402 -1508 0 3
rlabel polysilicon 1409 -1502 1409 -1502 0 1
rlabel polysilicon 1409 -1508 1409 -1508 0 3
rlabel polysilicon 1416 -1502 1416 -1502 0 1
rlabel polysilicon 1416 -1508 1416 -1508 0 3
rlabel polysilicon 1423 -1502 1423 -1502 0 1
rlabel polysilicon 1423 -1508 1423 -1508 0 3
rlabel polysilicon 1430 -1502 1430 -1502 0 1
rlabel polysilicon 1430 -1508 1430 -1508 0 3
rlabel polysilicon 1437 -1502 1437 -1502 0 1
rlabel polysilicon 1437 -1508 1437 -1508 0 3
rlabel polysilicon 1444 -1502 1444 -1502 0 1
rlabel polysilicon 1444 -1508 1444 -1508 0 3
rlabel polysilicon 1451 -1502 1451 -1502 0 1
rlabel polysilicon 1451 -1508 1451 -1508 0 3
rlabel polysilicon 1454 -1508 1454 -1508 0 4
rlabel polysilicon 1458 -1502 1458 -1502 0 1
rlabel polysilicon 1458 -1508 1458 -1508 0 3
rlabel polysilicon 1465 -1502 1465 -1502 0 1
rlabel polysilicon 1465 -1508 1465 -1508 0 3
rlabel polysilicon 1472 -1502 1472 -1502 0 1
rlabel polysilicon 1472 -1508 1472 -1508 0 3
rlabel polysilicon 1479 -1502 1479 -1502 0 1
rlabel polysilicon 1479 -1508 1479 -1508 0 3
rlabel polysilicon 1486 -1502 1486 -1502 0 1
rlabel polysilicon 1486 -1508 1486 -1508 0 3
rlabel polysilicon 1493 -1502 1493 -1502 0 1
rlabel polysilicon 1493 -1508 1493 -1508 0 3
rlabel polysilicon 1500 -1502 1500 -1502 0 1
rlabel polysilicon 1500 -1508 1500 -1508 0 3
rlabel polysilicon 1507 -1502 1507 -1502 0 1
rlabel polysilicon 1507 -1508 1507 -1508 0 3
rlabel polysilicon 1514 -1502 1514 -1502 0 1
rlabel polysilicon 1514 -1508 1514 -1508 0 3
rlabel polysilicon 1521 -1502 1521 -1502 0 1
rlabel polysilicon 1521 -1508 1521 -1508 0 3
rlabel polysilicon 1528 -1502 1528 -1502 0 1
rlabel polysilicon 1528 -1508 1528 -1508 0 3
rlabel polysilicon 1535 -1502 1535 -1502 0 1
rlabel polysilicon 1538 -1502 1538 -1502 0 2
rlabel polysilicon 1535 -1508 1535 -1508 0 3
rlabel polysilicon 1538 -1508 1538 -1508 0 4
rlabel polysilicon 1542 -1502 1542 -1502 0 1
rlabel polysilicon 1542 -1508 1542 -1508 0 3
rlabel polysilicon 1549 -1502 1549 -1502 0 1
rlabel polysilicon 1552 -1502 1552 -1502 0 2
rlabel polysilicon 1549 -1508 1549 -1508 0 3
rlabel polysilicon 1556 -1502 1556 -1502 0 1
rlabel polysilicon 1556 -1508 1556 -1508 0 3
rlabel polysilicon 1563 -1502 1563 -1502 0 1
rlabel polysilicon 1563 -1508 1563 -1508 0 3
rlabel polysilicon 1570 -1502 1570 -1502 0 1
rlabel polysilicon 1570 -1508 1570 -1508 0 3
rlabel polysilicon 1577 -1502 1577 -1502 0 1
rlabel polysilicon 1577 -1508 1577 -1508 0 3
rlabel polysilicon 1584 -1502 1584 -1502 0 1
rlabel polysilicon 1587 -1502 1587 -1502 0 2
rlabel polysilicon 1584 -1508 1584 -1508 0 3
rlabel polysilicon 1591 -1502 1591 -1502 0 1
rlabel polysilicon 1591 -1508 1591 -1508 0 3
rlabel polysilicon 1598 -1502 1598 -1502 0 1
rlabel polysilicon 1598 -1508 1598 -1508 0 3
rlabel polysilicon 1605 -1502 1605 -1502 0 1
rlabel polysilicon 1608 -1502 1608 -1502 0 2
rlabel polysilicon 1605 -1508 1605 -1508 0 3
rlabel polysilicon 1608 -1508 1608 -1508 0 4
rlabel polysilicon 1612 -1502 1612 -1502 0 1
rlabel polysilicon 1612 -1508 1612 -1508 0 3
rlabel polysilicon 1619 -1502 1619 -1502 0 1
rlabel polysilicon 1619 -1508 1619 -1508 0 3
rlabel polysilicon 1626 -1502 1626 -1502 0 1
rlabel polysilicon 1626 -1508 1626 -1508 0 3
rlabel polysilicon 1633 -1502 1633 -1502 0 1
rlabel polysilicon 1633 -1508 1633 -1508 0 3
rlabel polysilicon 1643 -1502 1643 -1502 0 2
rlabel polysilicon 1640 -1508 1640 -1508 0 3
rlabel polysilicon 1643 -1508 1643 -1508 0 4
rlabel polysilicon 1647 -1502 1647 -1502 0 1
rlabel polysilicon 1647 -1508 1647 -1508 0 3
rlabel polysilicon 1654 -1502 1654 -1502 0 1
rlabel polysilicon 1654 -1508 1654 -1508 0 3
rlabel polysilicon 1661 -1502 1661 -1502 0 1
rlabel polysilicon 1661 -1508 1661 -1508 0 3
rlabel polysilicon 1668 -1502 1668 -1502 0 1
rlabel polysilicon 1668 -1508 1668 -1508 0 3
rlabel polysilicon 1675 -1502 1675 -1502 0 1
rlabel polysilicon 1675 -1508 1675 -1508 0 3
rlabel polysilicon 1682 -1502 1682 -1502 0 1
rlabel polysilicon 1682 -1508 1682 -1508 0 3
rlabel polysilicon 1689 -1502 1689 -1502 0 1
rlabel polysilicon 1689 -1508 1689 -1508 0 3
rlabel polysilicon 1696 -1502 1696 -1502 0 1
rlabel polysilicon 1696 -1508 1696 -1508 0 3
rlabel polysilicon 1703 -1502 1703 -1502 0 1
rlabel polysilicon 1703 -1508 1703 -1508 0 3
rlabel polysilicon 1710 -1502 1710 -1502 0 1
rlabel polysilicon 1710 -1508 1710 -1508 0 3
rlabel polysilicon 1717 -1502 1717 -1502 0 1
rlabel polysilicon 1717 -1508 1717 -1508 0 3
rlabel polysilicon 1724 -1502 1724 -1502 0 1
rlabel polysilicon 1724 -1508 1724 -1508 0 3
rlabel polysilicon 1731 -1502 1731 -1502 0 1
rlabel polysilicon 1731 -1508 1731 -1508 0 3
rlabel polysilicon 1801 -1502 1801 -1502 0 1
rlabel polysilicon 1801 -1508 1801 -1508 0 3
rlabel polysilicon 23 -1637 23 -1637 0 1
rlabel polysilicon 23 -1643 23 -1643 0 3
rlabel polysilicon 30 -1637 30 -1637 0 1
rlabel polysilicon 30 -1643 30 -1643 0 3
rlabel polysilicon 37 -1637 37 -1637 0 1
rlabel polysilicon 37 -1643 37 -1643 0 3
rlabel polysilicon 44 -1637 44 -1637 0 1
rlabel polysilicon 44 -1643 44 -1643 0 3
rlabel polysilicon 51 -1637 51 -1637 0 1
rlabel polysilicon 51 -1643 51 -1643 0 3
rlabel polysilicon 61 -1637 61 -1637 0 2
rlabel polysilicon 65 -1637 65 -1637 0 1
rlabel polysilicon 65 -1643 65 -1643 0 3
rlabel polysilicon 72 -1637 72 -1637 0 1
rlabel polysilicon 72 -1643 72 -1643 0 3
rlabel polysilicon 79 -1637 79 -1637 0 1
rlabel polysilicon 79 -1643 79 -1643 0 3
rlabel polysilicon 86 -1637 86 -1637 0 1
rlabel polysilicon 86 -1643 86 -1643 0 3
rlabel polysilicon 93 -1637 93 -1637 0 1
rlabel polysilicon 93 -1643 93 -1643 0 3
rlabel polysilicon 100 -1637 100 -1637 0 1
rlabel polysilicon 100 -1643 100 -1643 0 3
rlabel polysilicon 107 -1637 107 -1637 0 1
rlabel polysilicon 107 -1643 107 -1643 0 3
rlabel polysilicon 114 -1637 114 -1637 0 1
rlabel polysilicon 114 -1643 114 -1643 0 3
rlabel polysilicon 121 -1637 121 -1637 0 1
rlabel polysilicon 124 -1637 124 -1637 0 2
rlabel polysilicon 121 -1643 121 -1643 0 3
rlabel polysilicon 124 -1643 124 -1643 0 4
rlabel polysilicon 128 -1637 128 -1637 0 1
rlabel polysilicon 128 -1643 128 -1643 0 3
rlabel polysilicon 135 -1637 135 -1637 0 1
rlabel polysilicon 135 -1643 135 -1643 0 3
rlabel polysilicon 142 -1637 142 -1637 0 1
rlabel polysilicon 142 -1643 142 -1643 0 3
rlabel polysilicon 149 -1637 149 -1637 0 1
rlabel polysilicon 149 -1643 149 -1643 0 3
rlabel polysilicon 156 -1637 156 -1637 0 1
rlabel polysilicon 156 -1643 156 -1643 0 3
rlabel polysilicon 163 -1637 163 -1637 0 1
rlabel polysilicon 166 -1637 166 -1637 0 2
rlabel polysilicon 163 -1643 163 -1643 0 3
rlabel polysilicon 170 -1637 170 -1637 0 1
rlabel polysilicon 170 -1643 170 -1643 0 3
rlabel polysilicon 177 -1637 177 -1637 0 1
rlabel polysilicon 177 -1643 177 -1643 0 3
rlabel polysilicon 184 -1637 184 -1637 0 1
rlabel polysilicon 187 -1637 187 -1637 0 2
rlabel polysilicon 184 -1643 184 -1643 0 3
rlabel polysilicon 187 -1643 187 -1643 0 4
rlabel polysilicon 191 -1637 191 -1637 0 1
rlabel polysilicon 191 -1643 191 -1643 0 3
rlabel polysilicon 198 -1637 198 -1637 0 1
rlabel polysilicon 198 -1643 198 -1643 0 3
rlabel polysilicon 205 -1637 205 -1637 0 1
rlabel polysilicon 205 -1643 205 -1643 0 3
rlabel polysilicon 212 -1637 212 -1637 0 1
rlabel polysilicon 212 -1643 212 -1643 0 3
rlabel polysilicon 219 -1637 219 -1637 0 1
rlabel polysilicon 222 -1637 222 -1637 0 2
rlabel polysilicon 219 -1643 219 -1643 0 3
rlabel polysilicon 222 -1643 222 -1643 0 4
rlabel polysilicon 226 -1637 226 -1637 0 1
rlabel polysilicon 226 -1643 226 -1643 0 3
rlabel polysilicon 233 -1637 233 -1637 0 1
rlabel polysilicon 233 -1643 233 -1643 0 3
rlabel polysilicon 240 -1637 240 -1637 0 1
rlabel polysilicon 240 -1643 240 -1643 0 3
rlabel polysilicon 247 -1637 247 -1637 0 1
rlabel polysilicon 247 -1643 247 -1643 0 3
rlabel polysilicon 254 -1637 254 -1637 0 1
rlabel polysilicon 254 -1643 254 -1643 0 3
rlabel polysilicon 264 -1637 264 -1637 0 2
rlabel polysilicon 261 -1643 261 -1643 0 3
rlabel polysilicon 268 -1637 268 -1637 0 1
rlabel polysilicon 268 -1643 268 -1643 0 3
rlabel polysilicon 275 -1637 275 -1637 0 1
rlabel polysilicon 275 -1643 275 -1643 0 3
rlabel polysilicon 282 -1637 282 -1637 0 1
rlabel polysilicon 282 -1643 282 -1643 0 3
rlabel polysilicon 289 -1637 289 -1637 0 1
rlabel polysilicon 289 -1643 289 -1643 0 3
rlabel polysilicon 296 -1637 296 -1637 0 1
rlabel polysilicon 296 -1643 296 -1643 0 3
rlabel polysilicon 303 -1637 303 -1637 0 1
rlabel polysilicon 303 -1643 303 -1643 0 3
rlabel polysilicon 310 -1637 310 -1637 0 1
rlabel polysilicon 313 -1637 313 -1637 0 2
rlabel polysilicon 310 -1643 310 -1643 0 3
rlabel polysilicon 317 -1637 317 -1637 0 1
rlabel polysilicon 317 -1643 317 -1643 0 3
rlabel polysilicon 324 -1637 324 -1637 0 1
rlabel polysilicon 324 -1643 324 -1643 0 3
rlabel polysilicon 331 -1637 331 -1637 0 1
rlabel polysilicon 331 -1643 331 -1643 0 3
rlabel polysilicon 338 -1637 338 -1637 0 1
rlabel polysilicon 338 -1643 338 -1643 0 3
rlabel polysilicon 345 -1637 345 -1637 0 1
rlabel polysilicon 345 -1643 345 -1643 0 3
rlabel polysilicon 352 -1637 352 -1637 0 1
rlabel polysilicon 352 -1643 352 -1643 0 3
rlabel polysilicon 359 -1637 359 -1637 0 1
rlabel polysilicon 359 -1643 359 -1643 0 3
rlabel polysilicon 366 -1637 366 -1637 0 1
rlabel polysilicon 366 -1643 366 -1643 0 3
rlabel polysilicon 373 -1637 373 -1637 0 1
rlabel polysilicon 373 -1643 373 -1643 0 3
rlabel polysilicon 380 -1637 380 -1637 0 1
rlabel polysilicon 380 -1643 380 -1643 0 3
rlabel polysilicon 387 -1637 387 -1637 0 1
rlabel polysilicon 387 -1643 387 -1643 0 3
rlabel polysilicon 394 -1637 394 -1637 0 1
rlabel polysilicon 394 -1643 394 -1643 0 3
rlabel polysilicon 401 -1637 401 -1637 0 1
rlabel polysilicon 401 -1643 401 -1643 0 3
rlabel polysilicon 408 -1637 408 -1637 0 1
rlabel polysilicon 408 -1643 408 -1643 0 3
rlabel polysilicon 415 -1637 415 -1637 0 1
rlabel polysilicon 415 -1643 415 -1643 0 3
rlabel polysilicon 422 -1637 422 -1637 0 1
rlabel polysilicon 422 -1643 422 -1643 0 3
rlabel polysilicon 429 -1637 429 -1637 0 1
rlabel polysilicon 429 -1643 429 -1643 0 3
rlabel polysilicon 436 -1637 436 -1637 0 1
rlabel polysilicon 436 -1643 436 -1643 0 3
rlabel polysilicon 443 -1637 443 -1637 0 1
rlabel polysilicon 446 -1637 446 -1637 0 2
rlabel polysilicon 443 -1643 443 -1643 0 3
rlabel polysilicon 446 -1643 446 -1643 0 4
rlabel polysilicon 450 -1637 450 -1637 0 1
rlabel polysilicon 450 -1643 450 -1643 0 3
rlabel polysilicon 453 -1643 453 -1643 0 4
rlabel polysilicon 457 -1637 457 -1637 0 1
rlabel polysilicon 457 -1643 457 -1643 0 3
rlabel polysilicon 464 -1637 464 -1637 0 1
rlabel polysilicon 464 -1643 464 -1643 0 3
rlabel polysilicon 471 -1637 471 -1637 0 1
rlabel polysilicon 471 -1643 471 -1643 0 3
rlabel polysilicon 478 -1637 478 -1637 0 1
rlabel polysilicon 478 -1643 478 -1643 0 3
rlabel polysilicon 485 -1643 485 -1643 0 3
rlabel polysilicon 492 -1637 492 -1637 0 1
rlabel polysilicon 492 -1643 492 -1643 0 3
rlabel polysilicon 499 -1637 499 -1637 0 1
rlabel polysilicon 499 -1643 499 -1643 0 3
rlabel polysilicon 506 -1637 506 -1637 0 1
rlabel polysilicon 506 -1643 506 -1643 0 3
rlabel polysilicon 513 -1637 513 -1637 0 1
rlabel polysilicon 513 -1643 513 -1643 0 3
rlabel polysilicon 520 -1637 520 -1637 0 1
rlabel polysilicon 520 -1643 520 -1643 0 3
rlabel polysilicon 527 -1637 527 -1637 0 1
rlabel polysilicon 527 -1643 527 -1643 0 3
rlabel polysilicon 534 -1637 534 -1637 0 1
rlabel polysilicon 534 -1643 534 -1643 0 3
rlabel polysilicon 541 -1637 541 -1637 0 1
rlabel polysilicon 544 -1637 544 -1637 0 2
rlabel polysilicon 541 -1643 541 -1643 0 3
rlabel polysilicon 544 -1643 544 -1643 0 4
rlabel polysilicon 548 -1637 548 -1637 0 1
rlabel polysilicon 551 -1637 551 -1637 0 2
rlabel polysilicon 548 -1643 548 -1643 0 3
rlabel polysilicon 551 -1643 551 -1643 0 4
rlabel polysilicon 555 -1637 555 -1637 0 1
rlabel polysilicon 555 -1643 555 -1643 0 3
rlabel polysilicon 562 -1637 562 -1637 0 1
rlabel polysilicon 562 -1643 562 -1643 0 3
rlabel polysilicon 569 -1637 569 -1637 0 1
rlabel polysilicon 569 -1643 569 -1643 0 3
rlabel polysilicon 576 -1637 576 -1637 0 1
rlabel polysilicon 576 -1643 576 -1643 0 3
rlabel polysilicon 583 -1637 583 -1637 0 1
rlabel polysilicon 583 -1643 583 -1643 0 3
rlabel polysilicon 590 -1637 590 -1637 0 1
rlabel polysilicon 590 -1643 590 -1643 0 3
rlabel polysilicon 597 -1637 597 -1637 0 1
rlabel polysilicon 597 -1643 597 -1643 0 3
rlabel polysilicon 604 -1637 604 -1637 0 1
rlabel polysilicon 607 -1637 607 -1637 0 2
rlabel polysilicon 607 -1643 607 -1643 0 4
rlabel polysilicon 611 -1637 611 -1637 0 1
rlabel polysilicon 611 -1643 611 -1643 0 3
rlabel polysilicon 618 -1637 618 -1637 0 1
rlabel polysilicon 618 -1643 618 -1643 0 3
rlabel polysilicon 625 -1637 625 -1637 0 1
rlabel polysilicon 625 -1643 625 -1643 0 3
rlabel polysilicon 632 -1637 632 -1637 0 1
rlabel polysilicon 632 -1643 632 -1643 0 3
rlabel polysilicon 639 -1637 639 -1637 0 1
rlabel polysilicon 639 -1643 639 -1643 0 3
rlabel polysilicon 646 -1637 646 -1637 0 1
rlabel polysilicon 646 -1643 646 -1643 0 3
rlabel polysilicon 653 -1637 653 -1637 0 1
rlabel polysilicon 653 -1643 653 -1643 0 3
rlabel polysilicon 660 -1637 660 -1637 0 1
rlabel polysilicon 660 -1643 660 -1643 0 3
rlabel polysilicon 667 -1637 667 -1637 0 1
rlabel polysilicon 667 -1643 667 -1643 0 3
rlabel polysilicon 674 -1637 674 -1637 0 1
rlabel polysilicon 674 -1643 674 -1643 0 3
rlabel polysilicon 681 -1637 681 -1637 0 1
rlabel polysilicon 681 -1643 681 -1643 0 3
rlabel polysilicon 688 -1637 688 -1637 0 1
rlabel polysilicon 688 -1643 688 -1643 0 3
rlabel polysilicon 695 -1637 695 -1637 0 1
rlabel polysilicon 695 -1643 695 -1643 0 3
rlabel polysilicon 702 -1637 702 -1637 0 1
rlabel polysilicon 702 -1643 702 -1643 0 3
rlabel polysilicon 709 -1637 709 -1637 0 1
rlabel polysilicon 709 -1643 709 -1643 0 3
rlabel polysilicon 716 -1637 716 -1637 0 1
rlabel polysilicon 716 -1643 716 -1643 0 3
rlabel polysilicon 723 -1637 723 -1637 0 1
rlabel polysilicon 726 -1637 726 -1637 0 2
rlabel polysilicon 726 -1643 726 -1643 0 4
rlabel polysilicon 730 -1637 730 -1637 0 1
rlabel polysilicon 733 -1637 733 -1637 0 2
rlabel polysilicon 730 -1643 730 -1643 0 3
rlabel polysilicon 733 -1643 733 -1643 0 4
rlabel polysilicon 737 -1637 737 -1637 0 1
rlabel polysilicon 737 -1643 737 -1643 0 3
rlabel polysilicon 747 -1637 747 -1637 0 2
rlabel polysilicon 744 -1643 744 -1643 0 3
rlabel polysilicon 747 -1643 747 -1643 0 4
rlabel polysilicon 751 -1637 751 -1637 0 1
rlabel polysilicon 754 -1637 754 -1637 0 2
rlabel polysilicon 751 -1643 751 -1643 0 3
rlabel polysilicon 754 -1643 754 -1643 0 4
rlabel polysilicon 758 -1637 758 -1637 0 1
rlabel polysilicon 758 -1643 758 -1643 0 3
rlabel polysilicon 765 -1637 765 -1637 0 1
rlabel polysilicon 765 -1643 765 -1643 0 3
rlabel polysilicon 772 -1637 772 -1637 0 1
rlabel polysilicon 772 -1643 772 -1643 0 3
rlabel polysilicon 779 -1637 779 -1637 0 1
rlabel polysilicon 779 -1643 779 -1643 0 3
rlabel polysilicon 786 -1637 786 -1637 0 1
rlabel polysilicon 786 -1643 786 -1643 0 3
rlabel polysilicon 793 -1637 793 -1637 0 1
rlabel polysilicon 793 -1643 793 -1643 0 3
rlabel polysilicon 800 -1637 800 -1637 0 1
rlabel polysilicon 800 -1643 800 -1643 0 3
rlabel polysilicon 807 -1637 807 -1637 0 1
rlabel polysilicon 807 -1643 807 -1643 0 3
rlabel polysilicon 814 -1637 814 -1637 0 1
rlabel polysilicon 817 -1637 817 -1637 0 2
rlabel polysilicon 814 -1643 814 -1643 0 3
rlabel polysilicon 817 -1643 817 -1643 0 4
rlabel polysilicon 821 -1637 821 -1637 0 1
rlabel polysilicon 824 -1637 824 -1637 0 2
rlabel polysilicon 824 -1643 824 -1643 0 4
rlabel polysilicon 828 -1637 828 -1637 0 1
rlabel polysilicon 828 -1643 828 -1643 0 3
rlabel polysilicon 835 -1637 835 -1637 0 1
rlabel polysilicon 835 -1643 835 -1643 0 3
rlabel polysilicon 842 -1637 842 -1637 0 1
rlabel polysilicon 842 -1643 842 -1643 0 3
rlabel polysilicon 849 -1637 849 -1637 0 1
rlabel polysilicon 849 -1643 849 -1643 0 3
rlabel polysilicon 859 -1643 859 -1643 0 4
rlabel polysilicon 863 -1637 863 -1637 0 1
rlabel polysilicon 866 -1637 866 -1637 0 2
rlabel polysilicon 863 -1643 863 -1643 0 3
rlabel polysilicon 866 -1643 866 -1643 0 4
rlabel polysilicon 870 -1637 870 -1637 0 1
rlabel polysilicon 870 -1643 870 -1643 0 3
rlabel polysilicon 877 -1637 877 -1637 0 1
rlabel polysilicon 880 -1637 880 -1637 0 2
rlabel polysilicon 877 -1643 877 -1643 0 3
rlabel polysilicon 880 -1643 880 -1643 0 4
rlabel polysilicon 884 -1637 884 -1637 0 1
rlabel polysilicon 884 -1643 884 -1643 0 3
rlabel polysilicon 891 -1637 891 -1637 0 1
rlabel polysilicon 894 -1637 894 -1637 0 2
rlabel polysilicon 891 -1643 891 -1643 0 3
rlabel polysilicon 898 -1637 898 -1637 0 1
rlabel polysilicon 898 -1643 898 -1643 0 3
rlabel polysilicon 905 -1637 905 -1637 0 1
rlabel polysilicon 905 -1643 905 -1643 0 3
rlabel polysilicon 912 -1637 912 -1637 0 1
rlabel polysilicon 912 -1643 912 -1643 0 3
rlabel polysilicon 919 -1637 919 -1637 0 1
rlabel polysilicon 919 -1643 919 -1643 0 3
rlabel polysilicon 926 -1637 926 -1637 0 1
rlabel polysilicon 926 -1643 926 -1643 0 3
rlabel polysilicon 933 -1637 933 -1637 0 1
rlabel polysilicon 933 -1643 933 -1643 0 3
rlabel polysilicon 940 -1637 940 -1637 0 1
rlabel polysilicon 940 -1643 940 -1643 0 3
rlabel polysilicon 947 -1637 947 -1637 0 1
rlabel polysilicon 947 -1643 947 -1643 0 3
rlabel polysilicon 954 -1637 954 -1637 0 1
rlabel polysilicon 957 -1637 957 -1637 0 2
rlabel polysilicon 957 -1643 957 -1643 0 4
rlabel polysilicon 961 -1637 961 -1637 0 1
rlabel polysilicon 961 -1643 961 -1643 0 3
rlabel polysilicon 968 -1637 968 -1637 0 1
rlabel polysilicon 968 -1643 968 -1643 0 3
rlabel polysilicon 975 -1637 975 -1637 0 1
rlabel polysilicon 975 -1643 975 -1643 0 3
rlabel polysilicon 982 -1637 982 -1637 0 1
rlabel polysilicon 982 -1643 982 -1643 0 3
rlabel polysilicon 989 -1637 989 -1637 0 1
rlabel polysilicon 989 -1643 989 -1643 0 3
rlabel polysilicon 996 -1637 996 -1637 0 1
rlabel polysilicon 996 -1643 996 -1643 0 3
rlabel polysilicon 1003 -1637 1003 -1637 0 1
rlabel polysilicon 1006 -1637 1006 -1637 0 2
rlabel polysilicon 1003 -1643 1003 -1643 0 3
rlabel polysilicon 1006 -1643 1006 -1643 0 4
rlabel polysilicon 1010 -1637 1010 -1637 0 1
rlabel polysilicon 1010 -1643 1010 -1643 0 3
rlabel polysilicon 1017 -1637 1017 -1637 0 1
rlabel polysilicon 1020 -1637 1020 -1637 0 2
rlabel polysilicon 1017 -1643 1017 -1643 0 3
rlabel polysilicon 1020 -1643 1020 -1643 0 4
rlabel polysilicon 1024 -1637 1024 -1637 0 1
rlabel polysilicon 1024 -1643 1024 -1643 0 3
rlabel polysilicon 1031 -1637 1031 -1637 0 1
rlabel polysilicon 1031 -1643 1031 -1643 0 3
rlabel polysilicon 1038 -1637 1038 -1637 0 1
rlabel polysilicon 1038 -1643 1038 -1643 0 3
rlabel polysilicon 1045 -1637 1045 -1637 0 1
rlabel polysilicon 1045 -1643 1045 -1643 0 3
rlabel polysilicon 1052 -1637 1052 -1637 0 1
rlabel polysilicon 1052 -1643 1052 -1643 0 3
rlabel polysilicon 1062 -1637 1062 -1637 0 2
rlabel polysilicon 1059 -1643 1059 -1643 0 3
rlabel polysilicon 1062 -1643 1062 -1643 0 4
rlabel polysilicon 1066 -1637 1066 -1637 0 1
rlabel polysilicon 1066 -1643 1066 -1643 0 3
rlabel polysilicon 1073 -1637 1073 -1637 0 1
rlabel polysilicon 1073 -1643 1073 -1643 0 3
rlabel polysilicon 1080 -1637 1080 -1637 0 1
rlabel polysilicon 1080 -1643 1080 -1643 0 3
rlabel polysilicon 1083 -1643 1083 -1643 0 4
rlabel polysilicon 1087 -1637 1087 -1637 0 1
rlabel polysilicon 1087 -1643 1087 -1643 0 3
rlabel polysilicon 1094 -1637 1094 -1637 0 1
rlabel polysilicon 1094 -1643 1094 -1643 0 3
rlabel polysilicon 1101 -1637 1101 -1637 0 1
rlabel polysilicon 1101 -1643 1101 -1643 0 3
rlabel polysilicon 1108 -1643 1108 -1643 0 3
rlabel polysilicon 1111 -1643 1111 -1643 0 4
rlabel polysilicon 1115 -1637 1115 -1637 0 1
rlabel polysilicon 1115 -1643 1115 -1643 0 3
rlabel polysilicon 1122 -1637 1122 -1637 0 1
rlabel polysilicon 1125 -1637 1125 -1637 0 2
rlabel polysilicon 1122 -1643 1122 -1643 0 3
rlabel polysilicon 1125 -1643 1125 -1643 0 4
rlabel polysilicon 1129 -1637 1129 -1637 0 1
rlabel polysilicon 1129 -1643 1129 -1643 0 3
rlabel polysilicon 1136 -1637 1136 -1637 0 1
rlabel polysilicon 1136 -1643 1136 -1643 0 3
rlabel polysilicon 1143 -1637 1143 -1637 0 1
rlabel polysilicon 1143 -1643 1143 -1643 0 3
rlabel polysilicon 1150 -1637 1150 -1637 0 1
rlabel polysilicon 1150 -1643 1150 -1643 0 3
rlabel polysilicon 1157 -1637 1157 -1637 0 1
rlabel polysilicon 1157 -1643 1157 -1643 0 3
rlabel polysilicon 1164 -1637 1164 -1637 0 1
rlabel polysilicon 1164 -1643 1164 -1643 0 3
rlabel polysilicon 1171 -1637 1171 -1637 0 1
rlabel polysilicon 1171 -1643 1171 -1643 0 3
rlabel polysilicon 1178 -1637 1178 -1637 0 1
rlabel polysilicon 1178 -1643 1178 -1643 0 3
rlabel polysilicon 1185 -1637 1185 -1637 0 1
rlabel polysilicon 1188 -1637 1188 -1637 0 2
rlabel polysilicon 1185 -1643 1185 -1643 0 3
rlabel polysilicon 1192 -1637 1192 -1637 0 1
rlabel polysilicon 1192 -1643 1192 -1643 0 3
rlabel polysilicon 1199 -1637 1199 -1637 0 1
rlabel polysilicon 1199 -1643 1199 -1643 0 3
rlabel polysilicon 1206 -1637 1206 -1637 0 1
rlabel polysilicon 1206 -1643 1206 -1643 0 3
rlabel polysilicon 1209 -1643 1209 -1643 0 4
rlabel polysilicon 1213 -1637 1213 -1637 0 1
rlabel polysilicon 1213 -1643 1213 -1643 0 3
rlabel polysilicon 1220 -1637 1220 -1637 0 1
rlabel polysilicon 1220 -1643 1220 -1643 0 3
rlabel polysilicon 1227 -1637 1227 -1637 0 1
rlabel polysilicon 1227 -1643 1227 -1643 0 3
rlabel polysilicon 1234 -1637 1234 -1637 0 1
rlabel polysilicon 1234 -1643 1234 -1643 0 3
rlabel polysilicon 1241 -1637 1241 -1637 0 1
rlabel polysilicon 1241 -1643 1241 -1643 0 3
rlabel polysilicon 1248 -1637 1248 -1637 0 1
rlabel polysilicon 1248 -1643 1248 -1643 0 3
rlabel polysilicon 1255 -1637 1255 -1637 0 1
rlabel polysilicon 1255 -1643 1255 -1643 0 3
rlabel polysilicon 1262 -1637 1262 -1637 0 1
rlabel polysilicon 1262 -1643 1262 -1643 0 3
rlabel polysilicon 1269 -1637 1269 -1637 0 1
rlabel polysilicon 1269 -1643 1269 -1643 0 3
rlabel polysilicon 1276 -1637 1276 -1637 0 1
rlabel polysilicon 1276 -1643 1276 -1643 0 3
rlabel polysilicon 1283 -1637 1283 -1637 0 1
rlabel polysilicon 1283 -1643 1283 -1643 0 3
rlabel polysilicon 1290 -1637 1290 -1637 0 1
rlabel polysilicon 1290 -1643 1290 -1643 0 3
rlabel polysilicon 1297 -1637 1297 -1637 0 1
rlabel polysilicon 1300 -1643 1300 -1643 0 4
rlabel polysilicon 1304 -1637 1304 -1637 0 1
rlabel polysilicon 1304 -1643 1304 -1643 0 3
rlabel polysilicon 1311 -1637 1311 -1637 0 1
rlabel polysilicon 1311 -1643 1311 -1643 0 3
rlabel polysilicon 1318 -1637 1318 -1637 0 1
rlabel polysilicon 1318 -1643 1318 -1643 0 3
rlabel polysilicon 1325 -1637 1325 -1637 0 1
rlabel polysilicon 1325 -1643 1325 -1643 0 3
rlabel polysilicon 1332 -1637 1332 -1637 0 1
rlabel polysilicon 1332 -1643 1332 -1643 0 3
rlabel polysilicon 1339 -1637 1339 -1637 0 1
rlabel polysilicon 1339 -1643 1339 -1643 0 3
rlabel polysilicon 1346 -1637 1346 -1637 0 1
rlabel polysilicon 1346 -1643 1346 -1643 0 3
rlabel polysilicon 1353 -1637 1353 -1637 0 1
rlabel polysilicon 1353 -1643 1353 -1643 0 3
rlabel polysilicon 1360 -1637 1360 -1637 0 1
rlabel polysilicon 1360 -1643 1360 -1643 0 3
rlabel polysilicon 1367 -1637 1367 -1637 0 1
rlabel polysilicon 1367 -1643 1367 -1643 0 3
rlabel polysilicon 1374 -1637 1374 -1637 0 1
rlabel polysilicon 1374 -1643 1374 -1643 0 3
rlabel polysilicon 1381 -1637 1381 -1637 0 1
rlabel polysilicon 1381 -1643 1381 -1643 0 3
rlabel polysilicon 1388 -1637 1388 -1637 0 1
rlabel polysilicon 1388 -1643 1388 -1643 0 3
rlabel polysilicon 1395 -1637 1395 -1637 0 1
rlabel polysilicon 1395 -1643 1395 -1643 0 3
rlabel polysilicon 1402 -1637 1402 -1637 0 1
rlabel polysilicon 1402 -1643 1402 -1643 0 3
rlabel polysilicon 1409 -1637 1409 -1637 0 1
rlabel polysilicon 1409 -1643 1409 -1643 0 3
rlabel polysilicon 1416 -1637 1416 -1637 0 1
rlabel polysilicon 1416 -1643 1416 -1643 0 3
rlabel polysilicon 1423 -1637 1423 -1637 0 1
rlabel polysilicon 1423 -1643 1423 -1643 0 3
rlabel polysilicon 1430 -1637 1430 -1637 0 1
rlabel polysilicon 1430 -1643 1430 -1643 0 3
rlabel polysilicon 1437 -1637 1437 -1637 0 1
rlabel polysilicon 1437 -1643 1437 -1643 0 3
rlabel polysilicon 1444 -1637 1444 -1637 0 1
rlabel polysilicon 1444 -1643 1444 -1643 0 3
rlabel polysilicon 1451 -1637 1451 -1637 0 1
rlabel polysilicon 1454 -1637 1454 -1637 0 2
rlabel polysilicon 1451 -1643 1451 -1643 0 3
rlabel polysilicon 1458 -1637 1458 -1637 0 1
rlabel polysilicon 1458 -1643 1458 -1643 0 3
rlabel polysilicon 1465 -1637 1465 -1637 0 1
rlabel polysilicon 1465 -1643 1465 -1643 0 3
rlabel polysilicon 1472 -1637 1472 -1637 0 1
rlabel polysilicon 1472 -1643 1472 -1643 0 3
rlabel polysilicon 1479 -1637 1479 -1637 0 1
rlabel polysilicon 1479 -1643 1479 -1643 0 3
rlabel polysilicon 1486 -1637 1486 -1637 0 1
rlabel polysilicon 1486 -1643 1486 -1643 0 3
rlabel polysilicon 1493 -1637 1493 -1637 0 1
rlabel polysilicon 1493 -1643 1493 -1643 0 3
rlabel polysilicon 1500 -1637 1500 -1637 0 1
rlabel polysilicon 1500 -1643 1500 -1643 0 3
rlabel polysilicon 1507 -1637 1507 -1637 0 1
rlabel polysilicon 1507 -1643 1507 -1643 0 3
rlabel polysilicon 1514 -1637 1514 -1637 0 1
rlabel polysilicon 1514 -1643 1514 -1643 0 3
rlabel polysilicon 1521 -1637 1521 -1637 0 1
rlabel polysilicon 1521 -1643 1521 -1643 0 3
rlabel polysilicon 1528 -1637 1528 -1637 0 1
rlabel polysilicon 1528 -1643 1528 -1643 0 3
rlabel polysilicon 1535 -1637 1535 -1637 0 1
rlabel polysilicon 1535 -1643 1535 -1643 0 3
rlabel polysilicon 1542 -1637 1542 -1637 0 1
rlabel polysilicon 1542 -1643 1542 -1643 0 3
rlabel polysilicon 1549 -1637 1549 -1637 0 1
rlabel polysilicon 1549 -1643 1549 -1643 0 3
rlabel polysilicon 1556 -1637 1556 -1637 0 1
rlabel polysilicon 1556 -1643 1556 -1643 0 3
rlabel polysilicon 1563 -1637 1563 -1637 0 1
rlabel polysilicon 1563 -1643 1563 -1643 0 3
rlabel polysilicon 1570 -1637 1570 -1637 0 1
rlabel polysilicon 1570 -1643 1570 -1643 0 3
rlabel polysilicon 1577 -1637 1577 -1637 0 1
rlabel polysilicon 1577 -1643 1577 -1643 0 3
rlabel polysilicon 1584 -1637 1584 -1637 0 1
rlabel polysilicon 1584 -1643 1584 -1643 0 3
rlabel polysilicon 1591 -1637 1591 -1637 0 1
rlabel polysilicon 1591 -1643 1591 -1643 0 3
rlabel polysilicon 1598 -1637 1598 -1637 0 1
rlabel polysilicon 1598 -1643 1598 -1643 0 3
rlabel polysilicon 1605 -1637 1605 -1637 0 1
rlabel polysilicon 1605 -1643 1605 -1643 0 3
rlabel polysilicon 1612 -1637 1612 -1637 0 1
rlabel polysilicon 1612 -1643 1612 -1643 0 3
rlabel polysilicon 1619 -1637 1619 -1637 0 1
rlabel polysilicon 1619 -1643 1619 -1643 0 3
rlabel polysilicon 1626 -1637 1626 -1637 0 1
rlabel polysilicon 1626 -1643 1626 -1643 0 3
rlabel polysilicon 1633 -1637 1633 -1637 0 1
rlabel polysilicon 1633 -1643 1633 -1643 0 3
rlabel polysilicon 1640 -1637 1640 -1637 0 1
rlabel polysilicon 1640 -1643 1640 -1643 0 3
rlabel polysilicon 1647 -1637 1647 -1637 0 1
rlabel polysilicon 1650 -1637 1650 -1637 0 2
rlabel polysilicon 1647 -1643 1647 -1643 0 3
rlabel polysilicon 1650 -1643 1650 -1643 0 4
rlabel polysilicon 1654 -1637 1654 -1637 0 1
rlabel polysilicon 1654 -1643 1654 -1643 0 3
rlabel polysilicon 1661 -1637 1661 -1637 0 1
rlabel polysilicon 1661 -1643 1661 -1643 0 3
rlabel polysilicon 1668 -1637 1668 -1637 0 1
rlabel polysilicon 1668 -1643 1668 -1643 0 3
rlabel polysilicon 1675 -1637 1675 -1637 0 1
rlabel polysilicon 1675 -1643 1675 -1643 0 3
rlabel polysilicon 1682 -1637 1682 -1637 0 1
rlabel polysilicon 1685 -1637 1685 -1637 0 2
rlabel polysilicon 1682 -1643 1682 -1643 0 3
rlabel polysilicon 1685 -1643 1685 -1643 0 4
rlabel polysilicon 1689 -1637 1689 -1637 0 1
rlabel polysilicon 1689 -1643 1689 -1643 0 3
rlabel polysilicon 1696 -1637 1696 -1637 0 1
rlabel polysilicon 1696 -1643 1696 -1643 0 3
rlabel polysilicon 1706 -1637 1706 -1637 0 2
rlabel polysilicon 1710 -1637 1710 -1637 0 1
rlabel polysilicon 1710 -1643 1710 -1643 0 3
rlabel polysilicon 1717 -1637 1717 -1637 0 1
rlabel polysilicon 1717 -1643 1717 -1643 0 3
rlabel polysilicon 1724 -1637 1724 -1637 0 1
rlabel polysilicon 1724 -1643 1724 -1643 0 3
rlabel polysilicon 1822 -1637 1822 -1637 0 1
rlabel polysilicon 1822 -1643 1822 -1643 0 3
rlabel polysilicon 23 -1784 23 -1784 0 1
rlabel polysilicon 23 -1790 23 -1790 0 3
rlabel polysilicon 30 -1784 30 -1784 0 1
rlabel polysilicon 30 -1790 30 -1790 0 3
rlabel polysilicon 37 -1784 37 -1784 0 1
rlabel polysilicon 37 -1790 37 -1790 0 3
rlabel polysilicon 44 -1784 44 -1784 0 1
rlabel polysilicon 44 -1790 44 -1790 0 3
rlabel polysilicon 51 -1784 51 -1784 0 1
rlabel polysilicon 51 -1790 51 -1790 0 3
rlabel polysilicon 58 -1784 58 -1784 0 1
rlabel polysilicon 58 -1790 58 -1790 0 3
rlabel polysilicon 65 -1784 65 -1784 0 1
rlabel polysilicon 65 -1790 65 -1790 0 3
rlabel polysilicon 72 -1784 72 -1784 0 1
rlabel polysilicon 72 -1790 72 -1790 0 3
rlabel polysilicon 75 -1790 75 -1790 0 4
rlabel polysilicon 79 -1784 79 -1784 0 1
rlabel polysilicon 79 -1790 79 -1790 0 3
rlabel polysilicon 86 -1784 86 -1784 0 1
rlabel polysilicon 89 -1784 89 -1784 0 2
rlabel polysilicon 86 -1790 86 -1790 0 3
rlabel polysilicon 89 -1790 89 -1790 0 4
rlabel polysilicon 93 -1784 93 -1784 0 1
rlabel polysilicon 93 -1790 93 -1790 0 3
rlabel polysilicon 100 -1784 100 -1784 0 1
rlabel polysilicon 100 -1790 100 -1790 0 3
rlabel polysilicon 107 -1784 107 -1784 0 1
rlabel polysilicon 107 -1790 107 -1790 0 3
rlabel polysilicon 114 -1784 114 -1784 0 1
rlabel polysilicon 117 -1790 117 -1790 0 4
rlabel polysilicon 121 -1784 121 -1784 0 1
rlabel polysilicon 121 -1790 121 -1790 0 3
rlabel polysilicon 128 -1784 128 -1784 0 1
rlabel polysilicon 128 -1790 128 -1790 0 3
rlabel polysilicon 135 -1784 135 -1784 0 1
rlabel polysilicon 135 -1790 135 -1790 0 3
rlabel polysilicon 145 -1784 145 -1784 0 2
rlabel polysilicon 145 -1790 145 -1790 0 4
rlabel polysilicon 149 -1784 149 -1784 0 1
rlabel polysilicon 149 -1790 149 -1790 0 3
rlabel polysilicon 156 -1784 156 -1784 0 1
rlabel polysilicon 159 -1784 159 -1784 0 2
rlabel polysilicon 156 -1790 156 -1790 0 3
rlabel polysilicon 159 -1790 159 -1790 0 4
rlabel polysilicon 163 -1784 163 -1784 0 1
rlabel polysilicon 163 -1790 163 -1790 0 3
rlabel polysilicon 170 -1784 170 -1784 0 1
rlabel polysilicon 170 -1790 170 -1790 0 3
rlabel polysilicon 177 -1784 177 -1784 0 1
rlabel polysilicon 177 -1790 177 -1790 0 3
rlabel polysilicon 184 -1784 184 -1784 0 1
rlabel polysilicon 184 -1790 184 -1790 0 3
rlabel polysilicon 191 -1784 191 -1784 0 1
rlabel polysilicon 191 -1790 191 -1790 0 3
rlabel polysilicon 198 -1784 198 -1784 0 1
rlabel polysilicon 198 -1790 198 -1790 0 3
rlabel polysilicon 205 -1784 205 -1784 0 1
rlabel polysilicon 205 -1790 205 -1790 0 3
rlabel polysilicon 212 -1784 212 -1784 0 1
rlabel polysilicon 219 -1784 219 -1784 0 1
rlabel polysilicon 222 -1784 222 -1784 0 2
rlabel polysilicon 219 -1790 219 -1790 0 3
rlabel polysilicon 222 -1790 222 -1790 0 4
rlabel polysilicon 226 -1784 226 -1784 0 1
rlabel polysilicon 226 -1790 226 -1790 0 3
rlabel polysilicon 236 -1784 236 -1784 0 2
rlabel polysilicon 233 -1790 233 -1790 0 3
rlabel polysilicon 236 -1790 236 -1790 0 4
rlabel polysilicon 240 -1784 240 -1784 0 1
rlabel polysilicon 240 -1790 240 -1790 0 3
rlabel polysilicon 247 -1784 247 -1784 0 1
rlabel polysilicon 247 -1790 247 -1790 0 3
rlabel polysilicon 254 -1784 254 -1784 0 1
rlabel polysilicon 254 -1790 254 -1790 0 3
rlabel polysilicon 261 -1790 261 -1790 0 3
rlabel polysilicon 264 -1790 264 -1790 0 4
rlabel polysilicon 268 -1784 268 -1784 0 1
rlabel polysilicon 268 -1790 268 -1790 0 3
rlabel polysilicon 275 -1784 275 -1784 0 1
rlabel polysilicon 275 -1790 275 -1790 0 3
rlabel polysilicon 282 -1784 282 -1784 0 1
rlabel polysilicon 282 -1790 282 -1790 0 3
rlabel polysilicon 289 -1784 289 -1784 0 1
rlabel polysilicon 289 -1790 289 -1790 0 3
rlabel polysilicon 296 -1784 296 -1784 0 1
rlabel polysilicon 296 -1790 296 -1790 0 3
rlabel polysilicon 303 -1784 303 -1784 0 1
rlabel polysilicon 303 -1790 303 -1790 0 3
rlabel polysilicon 310 -1784 310 -1784 0 1
rlabel polysilicon 310 -1790 310 -1790 0 3
rlabel polysilicon 317 -1784 317 -1784 0 1
rlabel polysilicon 317 -1790 317 -1790 0 3
rlabel polysilicon 324 -1784 324 -1784 0 1
rlabel polysilicon 324 -1790 324 -1790 0 3
rlabel polysilicon 331 -1784 331 -1784 0 1
rlabel polysilicon 331 -1790 331 -1790 0 3
rlabel polysilicon 338 -1784 338 -1784 0 1
rlabel polysilicon 338 -1790 338 -1790 0 3
rlabel polysilicon 345 -1784 345 -1784 0 1
rlabel polysilicon 345 -1790 345 -1790 0 3
rlabel polysilicon 352 -1784 352 -1784 0 1
rlabel polysilicon 352 -1790 352 -1790 0 3
rlabel polysilicon 362 -1784 362 -1784 0 2
rlabel polysilicon 359 -1790 359 -1790 0 3
rlabel polysilicon 362 -1790 362 -1790 0 4
rlabel polysilicon 366 -1784 366 -1784 0 1
rlabel polysilicon 366 -1790 366 -1790 0 3
rlabel polysilicon 373 -1784 373 -1784 0 1
rlabel polysilicon 373 -1790 373 -1790 0 3
rlabel polysilicon 383 -1784 383 -1784 0 2
rlabel polysilicon 380 -1790 380 -1790 0 3
rlabel polysilicon 383 -1790 383 -1790 0 4
rlabel polysilicon 387 -1784 387 -1784 0 1
rlabel polysilicon 387 -1790 387 -1790 0 3
rlabel polysilicon 394 -1784 394 -1784 0 1
rlabel polysilicon 394 -1790 394 -1790 0 3
rlabel polysilicon 401 -1784 401 -1784 0 1
rlabel polysilicon 401 -1790 401 -1790 0 3
rlabel polysilicon 408 -1784 408 -1784 0 1
rlabel polysilicon 408 -1790 408 -1790 0 3
rlabel polysilicon 415 -1784 415 -1784 0 1
rlabel polysilicon 415 -1790 415 -1790 0 3
rlabel polysilicon 422 -1784 422 -1784 0 1
rlabel polysilicon 422 -1790 422 -1790 0 3
rlabel polysilicon 429 -1784 429 -1784 0 1
rlabel polysilicon 429 -1790 429 -1790 0 3
rlabel polysilicon 436 -1784 436 -1784 0 1
rlabel polysilicon 436 -1790 436 -1790 0 3
rlabel polysilicon 443 -1784 443 -1784 0 1
rlabel polysilicon 443 -1790 443 -1790 0 3
rlabel polysilicon 450 -1784 450 -1784 0 1
rlabel polysilicon 450 -1790 450 -1790 0 3
rlabel polysilicon 457 -1784 457 -1784 0 1
rlabel polysilicon 457 -1790 457 -1790 0 3
rlabel polysilicon 464 -1784 464 -1784 0 1
rlabel polysilicon 464 -1790 464 -1790 0 3
rlabel polysilicon 471 -1784 471 -1784 0 1
rlabel polysilicon 471 -1790 471 -1790 0 3
rlabel polysilicon 478 -1784 478 -1784 0 1
rlabel polysilicon 478 -1790 478 -1790 0 3
rlabel polysilicon 485 -1784 485 -1784 0 1
rlabel polysilicon 485 -1790 485 -1790 0 3
rlabel polysilicon 492 -1784 492 -1784 0 1
rlabel polysilicon 492 -1790 492 -1790 0 3
rlabel polysilicon 499 -1784 499 -1784 0 1
rlabel polysilicon 502 -1784 502 -1784 0 2
rlabel polysilicon 499 -1790 499 -1790 0 3
rlabel polysilicon 502 -1790 502 -1790 0 4
rlabel polysilicon 506 -1784 506 -1784 0 1
rlabel polysilicon 506 -1790 506 -1790 0 3
rlabel polysilicon 513 -1784 513 -1784 0 1
rlabel polysilicon 513 -1790 513 -1790 0 3
rlabel polysilicon 520 -1784 520 -1784 0 1
rlabel polysilicon 520 -1790 520 -1790 0 3
rlabel polysilicon 527 -1784 527 -1784 0 1
rlabel polysilicon 527 -1790 527 -1790 0 3
rlabel polysilicon 534 -1784 534 -1784 0 1
rlabel polysilicon 537 -1784 537 -1784 0 2
rlabel polysilicon 534 -1790 534 -1790 0 3
rlabel polysilicon 537 -1790 537 -1790 0 4
rlabel polysilicon 541 -1784 541 -1784 0 1
rlabel polysilicon 544 -1784 544 -1784 0 2
rlabel polysilicon 544 -1790 544 -1790 0 4
rlabel polysilicon 548 -1784 548 -1784 0 1
rlabel polysilicon 551 -1784 551 -1784 0 2
rlabel polysilicon 548 -1790 548 -1790 0 3
rlabel polysilicon 551 -1790 551 -1790 0 4
rlabel polysilicon 555 -1784 555 -1784 0 1
rlabel polysilicon 555 -1790 555 -1790 0 3
rlabel polysilicon 562 -1784 562 -1784 0 1
rlabel polysilicon 562 -1790 562 -1790 0 3
rlabel polysilicon 569 -1784 569 -1784 0 1
rlabel polysilicon 569 -1790 569 -1790 0 3
rlabel polysilicon 576 -1784 576 -1784 0 1
rlabel polysilicon 579 -1784 579 -1784 0 2
rlabel polysilicon 579 -1790 579 -1790 0 4
rlabel polysilicon 583 -1784 583 -1784 0 1
rlabel polysilicon 583 -1790 583 -1790 0 3
rlabel polysilicon 593 -1784 593 -1784 0 2
rlabel polysilicon 590 -1790 590 -1790 0 3
rlabel polysilicon 593 -1790 593 -1790 0 4
rlabel polysilicon 597 -1784 597 -1784 0 1
rlabel polysilicon 597 -1790 597 -1790 0 3
rlabel polysilicon 604 -1784 604 -1784 0 1
rlabel polysilicon 604 -1790 604 -1790 0 3
rlabel polysilicon 611 -1784 611 -1784 0 1
rlabel polysilicon 611 -1790 611 -1790 0 3
rlabel polysilicon 618 -1784 618 -1784 0 1
rlabel polysilicon 618 -1790 618 -1790 0 3
rlabel polysilicon 625 -1784 625 -1784 0 1
rlabel polysilicon 625 -1790 625 -1790 0 3
rlabel polysilicon 635 -1784 635 -1784 0 2
rlabel polysilicon 632 -1790 632 -1790 0 3
rlabel polysilicon 635 -1790 635 -1790 0 4
rlabel polysilicon 639 -1784 639 -1784 0 1
rlabel polysilicon 639 -1790 639 -1790 0 3
rlabel polysilicon 646 -1784 646 -1784 0 1
rlabel polysilicon 646 -1790 646 -1790 0 3
rlabel polysilicon 653 -1784 653 -1784 0 1
rlabel polysilicon 653 -1790 653 -1790 0 3
rlabel polysilicon 660 -1784 660 -1784 0 1
rlabel polysilicon 660 -1790 660 -1790 0 3
rlabel polysilicon 667 -1784 667 -1784 0 1
rlabel polysilicon 667 -1790 667 -1790 0 3
rlabel polysilicon 674 -1784 674 -1784 0 1
rlabel polysilicon 677 -1784 677 -1784 0 2
rlabel polysilicon 674 -1790 674 -1790 0 3
rlabel polysilicon 677 -1790 677 -1790 0 4
rlabel polysilicon 681 -1784 681 -1784 0 1
rlabel polysilicon 681 -1790 681 -1790 0 3
rlabel polysilicon 688 -1784 688 -1784 0 1
rlabel polysilicon 688 -1790 688 -1790 0 3
rlabel polysilicon 695 -1784 695 -1784 0 1
rlabel polysilicon 695 -1790 695 -1790 0 3
rlabel polysilicon 702 -1784 702 -1784 0 1
rlabel polysilicon 705 -1784 705 -1784 0 2
rlabel polysilicon 702 -1790 702 -1790 0 3
rlabel polysilicon 709 -1784 709 -1784 0 1
rlabel polysilicon 709 -1790 709 -1790 0 3
rlabel polysilicon 716 -1784 716 -1784 0 1
rlabel polysilicon 719 -1784 719 -1784 0 2
rlabel polysilicon 716 -1790 716 -1790 0 3
rlabel polysilicon 719 -1790 719 -1790 0 4
rlabel polysilicon 723 -1784 723 -1784 0 1
rlabel polysilicon 726 -1784 726 -1784 0 2
rlabel polysilicon 726 -1790 726 -1790 0 4
rlabel polysilicon 730 -1784 730 -1784 0 1
rlabel polysilicon 733 -1790 733 -1790 0 4
rlabel polysilicon 737 -1784 737 -1784 0 1
rlabel polysilicon 737 -1790 737 -1790 0 3
rlabel polysilicon 744 -1784 744 -1784 0 1
rlabel polysilicon 744 -1790 744 -1790 0 3
rlabel polysilicon 751 -1784 751 -1784 0 1
rlabel polysilicon 751 -1790 751 -1790 0 3
rlabel polysilicon 758 -1784 758 -1784 0 1
rlabel polysilicon 758 -1790 758 -1790 0 3
rlabel polysilicon 765 -1784 765 -1784 0 1
rlabel polysilicon 765 -1790 765 -1790 0 3
rlabel polysilicon 772 -1784 772 -1784 0 1
rlabel polysilicon 772 -1790 772 -1790 0 3
rlabel polysilicon 779 -1784 779 -1784 0 1
rlabel polysilicon 782 -1784 782 -1784 0 2
rlabel polysilicon 779 -1790 779 -1790 0 3
rlabel polysilicon 782 -1790 782 -1790 0 4
rlabel polysilicon 786 -1784 786 -1784 0 1
rlabel polysilicon 789 -1784 789 -1784 0 2
rlabel polysilicon 786 -1790 786 -1790 0 3
rlabel polysilicon 789 -1790 789 -1790 0 4
rlabel polysilicon 793 -1784 793 -1784 0 1
rlabel polysilicon 793 -1790 793 -1790 0 3
rlabel polysilicon 800 -1784 800 -1784 0 1
rlabel polysilicon 800 -1790 800 -1790 0 3
rlabel polysilicon 807 -1784 807 -1784 0 1
rlabel polysilicon 807 -1790 807 -1790 0 3
rlabel polysilicon 814 -1784 814 -1784 0 1
rlabel polysilicon 814 -1790 814 -1790 0 3
rlabel polysilicon 824 -1784 824 -1784 0 2
rlabel polysilicon 821 -1790 821 -1790 0 3
rlabel polysilicon 824 -1790 824 -1790 0 4
rlabel polysilicon 828 -1784 828 -1784 0 1
rlabel polysilicon 828 -1790 828 -1790 0 3
rlabel polysilicon 835 -1784 835 -1784 0 1
rlabel polysilicon 835 -1790 835 -1790 0 3
rlabel polysilicon 842 -1784 842 -1784 0 1
rlabel polysilicon 842 -1790 842 -1790 0 3
rlabel polysilicon 849 -1784 849 -1784 0 1
rlabel polysilicon 849 -1790 849 -1790 0 3
rlabel polysilicon 856 -1784 856 -1784 0 1
rlabel polysilicon 856 -1790 856 -1790 0 3
rlabel polysilicon 863 -1784 863 -1784 0 1
rlabel polysilicon 863 -1790 863 -1790 0 3
rlabel polysilicon 870 -1784 870 -1784 0 1
rlabel polysilicon 870 -1790 870 -1790 0 3
rlabel polysilicon 877 -1784 877 -1784 0 1
rlabel polysilicon 877 -1790 877 -1790 0 3
rlabel polysilicon 884 -1784 884 -1784 0 1
rlabel polysilicon 887 -1784 887 -1784 0 2
rlabel polysilicon 884 -1790 884 -1790 0 3
rlabel polysilicon 887 -1790 887 -1790 0 4
rlabel polysilicon 891 -1784 891 -1784 0 1
rlabel polysilicon 891 -1790 891 -1790 0 3
rlabel polysilicon 898 -1784 898 -1784 0 1
rlabel polysilicon 901 -1784 901 -1784 0 2
rlabel polysilicon 898 -1790 898 -1790 0 3
rlabel polysilicon 901 -1790 901 -1790 0 4
rlabel polysilicon 905 -1784 905 -1784 0 1
rlabel polysilicon 905 -1790 905 -1790 0 3
rlabel polysilicon 912 -1784 912 -1784 0 1
rlabel polysilicon 912 -1790 912 -1790 0 3
rlabel polysilicon 919 -1784 919 -1784 0 1
rlabel polysilicon 919 -1790 919 -1790 0 3
rlabel polysilicon 926 -1784 926 -1784 0 1
rlabel polysilicon 926 -1790 926 -1790 0 3
rlabel polysilicon 933 -1784 933 -1784 0 1
rlabel polysilicon 933 -1790 933 -1790 0 3
rlabel polysilicon 940 -1784 940 -1784 0 1
rlabel polysilicon 940 -1790 940 -1790 0 3
rlabel polysilicon 947 -1784 947 -1784 0 1
rlabel polysilicon 950 -1784 950 -1784 0 2
rlabel polysilicon 947 -1790 947 -1790 0 3
rlabel polysilicon 954 -1784 954 -1784 0 1
rlabel polysilicon 954 -1790 954 -1790 0 3
rlabel polysilicon 961 -1784 961 -1784 0 1
rlabel polysilicon 961 -1790 961 -1790 0 3
rlabel polysilicon 968 -1784 968 -1784 0 1
rlabel polysilicon 968 -1790 968 -1790 0 3
rlabel polysilicon 978 -1784 978 -1784 0 2
rlabel polysilicon 975 -1790 975 -1790 0 3
rlabel polysilicon 978 -1790 978 -1790 0 4
rlabel polysilicon 982 -1784 982 -1784 0 1
rlabel polysilicon 982 -1790 982 -1790 0 3
rlabel polysilicon 989 -1784 989 -1784 0 1
rlabel polysilicon 989 -1790 989 -1790 0 3
rlabel polysilicon 996 -1784 996 -1784 0 1
rlabel polysilicon 996 -1790 996 -1790 0 3
rlabel polysilicon 1003 -1784 1003 -1784 0 1
rlabel polysilicon 1003 -1790 1003 -1790 0 3
rlabel polysilicon 1010 -1784 1010 -1784 0 1
rlabel polysilicon 1010 -1790 1010 -1790 0 3
rlabel polysilicon 1017 -1784 1017 -1784 0 1
rlabel polysilicon 1017 -1790 1017 -1790 0 3
rlabel polysilicon 1024 -1784 1024 -1784 0 1
rlabel polysilicon 1027 -1784 1027 -1784 0 2
rlabel polysilicon 1024 -1790 1024 -1790 0 3
rlabel polysilicon 1027 -1790 1027 -1790 0 4
rlabel polysilicon 1031 -1784 1031 -1784 0 1
rlabel polysilicon 1031 -1790 1031 -1790 0 3
rlabel polysilicon 1038 -1784 1038 -1784 0 1
rlabel polysilicon 1038 -1790 1038 -1790 0 3
rlabel polysilicon 1045 -1784 1045 -1784 0 1
rlabel polysilicon 1045 -1790 1045 -1790 0 3
rlabel polysilicon 1052 -1784 1052 -1784 0 1
rlabel polysilicon 1055 -1784 1055 -1784 0 2
rlabel polysilicon 1052 -1790 1052 -1790 0 3
rlabel polysilicon 1059 -1784 1059 -1784 0 1
rlabel polysilicon 1059 -1790 1059 -1790 0 3
rlabel polysilicon 1066 -1784 1066 -1784 0 1
rlabel polysilicon 1066 -1790 1066 -1790 0 3
rlabel polysilicon 1073 -1784 1073 -1784 0 1
rlabel polysilicon 1073 -1790 1073 -1790 0 3
rlabel polysilicon 1080 -1784 1080 -1784 0 1
rlabel polysilicon 1080 -1790 1080 -1790 0 3
rlabel polysilicon 1087 -1784 1087 -1784 0 1
rlabel polysilicon 1087 -1790 1087 -1790 0 3
rlabel polysilicon 1094 -1784 1094 -1784 0 1
rlabel polysilicon 1094 -1790 1094 -1790 0 3
rlabel polysilicon 1101 -1784 1101 -1784 0 1
rlabel polysilicon 1101 -1790 1101 -1790 0 3
rlabel polysilicon 1108 -1784 1108 -1784 0 1
rlabel polysilicon 1108 -1790 1108 -1790 0 3
rlabel polysilicon 1115 -1784 1115 -1784 0 1
rlabel polysilicon 1115 -1790 1115 -1790 0 3
rlabel polysilicon 1122 -1784 1122 -1784 0 1
rlabel polysilicon 1122 -1790 1122 -1790 0 3
rlabel polysilicon 1129 -1784 1129 -1784 0 1
rlabel polysilicon 1129 -1790 1129 -1790 0 3
rlabel polysilicon 1136 -1784 1136 -1784 0 1
rlabel polysilicon 1136 -1790 1136 -1790 0 3
rlabel polysilicon 1143 -1784 1143 -1784 0 1
rlabel polysilicon 1146 -1784 1146 -1784 0 2
rlabel polysilicon 1146 -1790 1146 -1790 0 4
rlabel polysilicon 1150 -1784 1150 -1784 0 1
rlabel polysilicon 1150 -1790 1150 -1790 0 3
rlabel polysilicon 1157 -1784 1157 -1784 0 1
rlabel polysilicon 1157 -1790 1157 -1790 0 3
rlabel polysilicon 1164 -1784 1164 -1784 0 1
rlabel polysilicon 1164 -1790 1164 -1790 0 3
rlabel polysilicon 1171 -1784 1171 -1784 0 1
rlabel polysilicon 1171 -1790 1171 -1790 0 3
rlabel polysilicon 1178 -1784 1178 -1784 0 1
rlabel polysilicon 1178 -1790 1178 -1790 0 3
rlabel polysilicon 1185 -1784 1185 -1784 0 1
rlabel polysilicon 1185 -1790 1185 -1790 0 3
rlabel polysilicon 1192 -1784 1192 -1784 0 1
rlabel polysilicon 1192 -1790 1192 -1790 0 3
rlabel polysilicon 1199 -1784 1199 -1784 0 1
rlabel polysilicon 1199 -1790 1199 -1790 0 3
rlabel polysilicon 1206 -1784 1206 -1784 0 1
rlabel polysilicon 1206 -1790 1206 -1790 0 3
rlabel polysilicon 1213 -1784 1213 -1784 0 1
rlabel polysilicon 1213 -1790 1213 -1790 0 3
rlabel polysilicon 1220 -1784 1220 -1784 0 1
rlabel polysilicon 1220 -1790 1220 -1790 0 3
rlabel polysilicon 1227 -1784 1227 -1784 0 1
rlabel polysilicon 1227 -1790 1227 -1790 0 3
rlabel polysilicon 1234 -1784 1234 -1784 0 1
rlabel polysilicon 1234 -1790 1234 -1790 0 3
rlabel polysilicon 1241 -1784 1241 -1784 0 1
rlabel polysilicon 1241 -1790 1241 -1790 0 3
rlabel polysilicon 1248 -1784 1248 -1784 0 1
rlabel polysilicon 1248 -1790 1248 -1790 0 3
rlabel polysilicon 1255 -1784 1255 -1784 0 1
rlabel polysilicon 1255 -1790 1255 -1790 0 3
rlabel polysilicon 1262 -1784 1262 -1784 0 1
rlabel polysilicon 1262 -1790 1262 -1790 0 3
rlabel polysilicon 1269 -1784 1269 -1784 0 1
rlabel polysilicon 1269 -1790 1269 -1790 0 3
rlabel polysilicon 1276 -1784 1276 -1784 0 1
rlabel polysilicon 1276 -1790 1276 -1790 0 3
rlabel polysilicon 1283 -1784 1283 -1784 0 1
rlabel polysilicon 1283 -1790 1283 -1790 0 3
rlabel polysilicon 1290 -1790 1290 -1790 0 3
rlabel polysilicon 1293 -1790 1293 -1790 0 4
rlabel polysilicon 1297 -1784 1297 -1784 0 1
rlabel polysilicon 1297 -1790 1297 -1790 0 3
rlabel polysilicon 1304 -1784 1304 -1784 0 1
rlabel polysilicon 1304 -1790 1304 -1790 0 3
rlabel polysilicon 1311 -1784 1311 -1784 0 1
rlabel polysilicon 1311 -1790 1311 -1790 0 3
rlabel polysilicon 1318 -1784 1318 -1784 0 1
rlabel polysilicon 1318 -1790 1318 -1790 0 3
rlabel polysilicon 1325 -1784 1325 -1784 0 1
rlabel polysilicon 1325 -1790 1325 -1790 0 3
rlabel polysilicon 1332 -1784 1332 -1784 0 1
rlabel polysilicon 1332 -1790 1332 -1790 0 3
rlabel polysilicon 1339 -1784 1339 -1784 0 1
rlabel polysilicon 1339 -1790 1339 -1790 0 3
rlabel polysilicon 1346 -1784 1346 -1784 0 1
rlabel polysilicon 1346 -1790 1346 -1790 0 3
rlabel polysilicon 1353 -1784 1353 -1784 0 1
rlabel polysilicon 1353 -1790 1353 -1790 0 3
rlabel polysilicon 1360 -1784 1360 -1784 0 1
rlabel polysilicon 1360 -1790 1360 -1790 0 3
rlabel polysilicon 1367 -1784 1367 -1784 0 1
rlabel polysilicon 1367 -1790 1367 -1790 0 3
rlabel polysilicon 1374 -1784 1374 -1784 0 1
rlabel polysilicon 1374 -1790 1374 -1790 0 3
rlabel polysilicon 1381 -1784 1381 -1784 0 1
rlabel polysilicon 1381 -1790 1381 -1790 0 3
rlabel polysilicon 1388 -1784 1388 -1784 0 1
rlabel polysilicon 1388 -1790 1388 -1790 0 3
rlabel polysilicon 1395 -1784 1395 -1784 0 1
rlabel polysilicon 1395 -1790 1395 -1790 0 3
rlabel polysilicon 1402 -1784 1402 -1784 0 1
rlabel polysilicon 1402 -1790 1402 -1790 0 3
rlabel polysilicon 1409 -1784 1409 -1784 0 1
rlabel polysilicon 1409 -1790 1409 -1790 0 3
rlabel polysilicon 1416 -1784 1416 -1784 0 1
rlabel polysilicon 1416 -1790 1416 -1790 0 3
rlabel polysilicon 1423 -1784 1423 -1784 0 1
rlabel polysilicon 1423 -1790 1423 -1790 0 3
rlabel polysilicon 1426 -1790 1426 -1790 0 4
rlabel polysilicon 1430 -1784 1430 -1784 0 1
rlabel polysilicon 1430 -1790 1430 -1790 0 3
rlabel polysilicon 1437 -1784 1437 -1784 0 1
rlabel polysilicon 1437 -1790 1437 -1790 0 3
rlabel polysilicon 1444 -1784 1444 -1784 0 1
rlabel polysilicon 1444 -1790 1444 -1790 0 3
rlabel polysilicon 1451 -1784 1451 -1784 0 1
rlabel polysilicon 1451 -1790 1451 -1790 0 3
rlabel polysilicon 1458 -1784 1458 -1784 0 1
rlabel polysilicon 1458 -1790 1458 -1790 0 3
rlabel polysilicon 1465 -1784 1465 -1784 0 1
rlabel polysilicon 1465 -1790 1465 -1790 0 3
rlabel polysilicon 1472 -1784 1472 -1784 0 1
rlabel polysilicon 1472 -1790 1472 -1790 0 3
rlabel polysilicon 1479 -1784 1479 -1784 0 1
rlabel polysilicon 1479 -1790 1479 -1790 0 3
rlabel polysilicon 1486 -1784 1486 -1784 0 1
rlabel polysilicon 1486 -1790 1486 -1790 0 3
rlabel polysilicon 1493 -1784 1493 -1784 0 1
rlabel polysilicon 1493 -1790 1493 -1790 0 3
rlabel polysilicon 1500 -1784 1500 -1784 0 1
rlabel polysilicon 1500 -1790 1500 -1790 0 3
rlabel polysilicon 1507 -1784 1507 -1784 0 1
rlabel polysilicon 1507 -1790 1507 -1790 0 3
rlabel polysilicon 1514 -1784 1514 -1784 0 1
rlabel polysilicon 1514 -1790 1514 -1790 0 3
rlabel polysilicon 1521 -1784 1521 -1784 0 1
rlabel polysilicon 1521 -1790 1521 -1790 0 3
rlabel polysilicon 1528 -1784 1528 -1784 0 1
rlabel polysilicon 1528 -1790 1528 -1790 0 3
rlabel polysilicon 1535 -1784 1535 -1784 0 1
rlabel polysilicon 1535 -1790 1535 -1790 0 3
rlabel polysilicon 1542 -1784 1542 -1784 0 1
rlabel polysilicon 1542 -1790 1542 -1790 0 3
rlabel polysilicon 1549 -1784 1549 -1784 0 1
rlabel polysilicon 1549 -1790 1549 -1790 0 3
rlabel polysilicon 1556 -1784 1556 -1784 0 1
rlabel polysilicon 1556 -1790 1556 -1790 0 3
rlabel polysilicon 1563 -1784 1563 -1784 0 1
rlabel polysilicon 1563 -1790 1563 -1790 0 3
rlabel polysilicon 1570 -1784 1570 -1784 0 1
rlabel polysilicon 1570 -1790 1570 -1790 0 3
rlabel polysilicon 1577 -1784 1577 -1784 0 1
rlabel polysilicon 1577 -1790 1577 -1790 0 3
rlabel polysilicon 1584 -1784 1584 -1784 0 1
rlabel polysilicon 1584 -1790 1584 -1790 0 3
rlabel polysilicon 1591 -1784 1591 -1784 0 1
rlabel polysilicon 1591 -1790 1591 -1790 0 3
rlabel polysilicon 1598 -1784 1598 -1784 0 1
rlabel polysilicon 1598 -1790 1598 -1790 0 3
rlabel polysilicon 1605 -1784 1605 -1784 0 1
rlabel polysilicon 1605 -1790 1605 -1790 0 3
rlabel polysilicon 1612 -1784 1612 -1784 0 1
rlabel polysilicon 1612 -1790 1612 -1790 0 3
rlabel polysilicon 1619 -1784 1619 -1784 0 1
rlabel polysilicon 1619 -1790 1619 -1790 0 3
rlabel polysilicon 1626 -1784 1626 -1784 0 1
rlabel polysilicon 1626 -1790 1626 -1790 0 3
rlabel polysilicon 1633 -1784 1633 -1784 0 1
rlabel polysilicon 1633 -1790 1633 -1790 0 3
rlabel polysilicon 1640 -1784 1640 -1784 0 1
rlabel polysilicon 1640 -1790 1640 -1790 0 3
rlabel polysilicon 1647 -1784 1647 -1784 0 1
rlabel polysilicon 1647 -1790 1647 -1790 0 3
rlabel polysilicon 1654 -1784 1654 -1784 0 1
rlabel polysilicon 1654 -1790 1654 -1790 0 3
rlabel polysilicon 1661 -1784 1661 -1784 0 1
rlabel polysilicon 1661 -1790 1661 -1790 0 3
rlabel polysilicon 1668 -1784 1668 -1784 0 1
rlabel polysilicon 1668 -1790 1668 -1790 0 3
rlabel polysilicon 1675 -1784 1675 -1784 0 1
rlabel polysilicon 1675 -1790 1675 -1790 0 3
rlabel polysilicon 1682 -1784 1682 -1784 0 1
rlabel polysilicon 1682 -1790 1682 -1790 0 3
rlabel polysilicon 1689 -1784 1689 -1784 0 1
rlabel polysilicon 1689 -1790 1689 -1790 0 3
rlabel polysilicon 1696 -1784 1696 -1784 0 1
rlabel polysilicon 1696 -1790 1696 -1790 0 3
rlabel polysilicon 1703 -1784 1703 -1784 0 1
rlabel polysilicon 1703 -1790 1703 -1790 0 3
rlabel polysilicon 1710 -1784 1710 -1784 0 1
rlabel polysilicon 1710 -1790 1710 -1790 0 3
rlabel polysilicon 1717 -1784 1717 -1784 0 1
rlabel polysilicon 1717 -1790 1717 -1790 0 3
rlabel polysilicon 1724 -1784 1724 -1784 0 1
rlabel polysilicon 1724 -1790 1724 -1790 0 3
rlabel polysilicon 1731 -1784 1731 -1784 0 1
rlabel polysilicon 1731 -1790 1731 -1790 0 3
rlabel polysilicon 1738 -1784 1738 -1784 0 1
rlabel polysilicon 1738 -1790 1738 -1790 0 3
rlabel polysilicon 1745 -1784 1745 -1784 0 1
rlabel polysilicon 1745 -1790 1745 -1790 0 3
rlabel polysilicon 1752 -1784 1752 -1784 0 1
rlabel polysilicon 1752 -1790 1752 -1790 0 3
rlabel polysilicon 1759 -1784 1759 -1784 0 1
rlabel polysilicon 1759 -1790 1759 -1790 0 3
rlabel polysilicon 1766 -1784 1766 -1784 0 1
rlabel polysilicon 1766 -1790 1766 -1790 0 3
rlabel polysilicon 1773 -1784 1773 -1784 0 1
rlabel polysilicon 1773 -1790 1773 -1790 0 3
rlabel polysilicon 1780 -1784 1780 -1784 0 1
rlabel polysilicon 1780 -1790 1780 -1790 0 3
rlabel polysilicon 1787 -1784 1787 -1784 0 1
rlabel polysilicon 1787 -1790 1787 -1790 0 3
rlabel polysilicon 1794 -1784 1794 -1784 0 1
rlabel polysilicon 1794 -1790 1794 -1790 0 3
rlabel polysilicon 1801 -1784 1801 -1784 0 1
rlabel polysilicon 1801 -1790 1801 -1790 0 3
rlabel polysilicon 1808 -1784 1808 -1784 0 1
rlabel polysilicon 1808 -1790 1808 -1790 0 3
rlabel polysilicon 1815 -1784 1815 -1784 0 1
rlabel polysilicon 1815 -1790 1815 -1790 0 3
rlabel polysilicon 1822 -1784 1822 -1784 0 1
rlabel polysilicon 1822 -1790 1822 -1790 0 3
rlabel polysilicon 1829 -1784 1829 -1784 0 1
rlabel polysilicon 1829 -1790 1829 -1790 0 3
rlabel polysilicon 1836 -1784 1836 -1784 0 1
rlabel polysilicon 1839 -1784 1839 -1784 0 2
rlabel polysilicon 1836 -1790 1836 -1790 0 3
rlabel polysilicon 1839 -1790 1839 -1790 0 4
rlabel polysilicon 30 -1923 30 -1923 0 1
rlabel polysilicon 30 -1929 30 -1929 0 3
rlabel polysilicon 37 -1923 37 -1923 0 1
rlabel polysilicon 37 -1929 37 -1929 0 3
rlabel polysilicon 44 -1923 44 -1923 0 1
rlabel polysilicon 44 -1929 44 -1929 0 3
rlabel polysilicon 51 -1923 51 -1923 0 1
rlabel polysilicon 51 -1929 51 -1929 0 3
rlabel polysilicon 58 -1923 58 -1923 0 1
rlabel polysilicon 61 -1923 61 -1923 0 2
rlabel polysilicon 61 -1929 61 -1929 0 4
rlabel polysilicon 68 -1923 68 -1923 0 2
rlabel polysilicon 65 -1929 65 -1929 0 3
rlabel polysilicon 68 -1929 68 -1929 0 4
rlabel polysilicon 72 -1923 72 -1923 0 1
rlabel polysilicon 72 -1929 72 -1929 0 3
rlabel polysilicon 79 -1923 79 -1923 0 1
rlabel polysilicon 79 -1929 79 -1929 0 3
rlabel polysilicon 86 -1923 86 -1923 0 1
rlabel polysilicon 86 -1929 86 -1929 0 3
rlabel polysilicon 93 -1923 93 -1923 0 1
rlabel polysilicon 93 -1929 93 -1929 0 3
rlabel polysilicon 100 -1923 100 -1923 0 1
rlabel polysilicon 100 -1929 100 -1929 0 3
rlabel polysilicon 107 -1923 107 -1923 0 1
rlabel polysilicon 110 -1923 110 -1923 0 2
rlabel polysilicon 107 -1929 107 -1929 0 3
rlabel polysilicon 114 -1923 114 -1923 0 1
rlabel polysilicon 114 -1929 114 -1929 0 3
rlabel polysilicon 121 -1923 121 -1923 0 1
rlabel polysilicon 121 -1929 121 -1929 0 3
rlabel polysilicon 128 -1923 128 -1923 0 1
rlabel polysilicon 128 -1929 128 -1929 0 3
rlabel polysilicon 135 -1923 135 -1923 0 1
rlabel polysilicon 135 -1929 135 -1929 0 3
rlabel polysilicon 142 -1923 142 -1923 0 1
rlabel polysilicon 142 -1929 142 -1929 0 3
rlabel polysilicon 149 -1923 149 -1923 0 1
rlabel polysilicon 149 -1929 149 -1929 0 3
rlabel polysilicon 156 -1923 156 -1923 0 1
rlabel polysilicon 156 -1929 156 -1929 0 3
rlabel polysilicon 163 -1923 163 -1923 0 1
rlabel polysilicon 163 -1929 163 -1929 0 3
rlabel polysilicon 173 -1923 173 -1923 0 2
rlabel polysilicon 170 -1929 170 -1929 0 3
rlabel polysilicon 173 -1929 173 -1929 0 4
rlabel polysilicon 177 -1923 177 -1923 0 1
rlabel polysilicon 177 -1929 177 -1929 0 3
rlabel polysilicon 184 -1923 184 -1923 0 1
rlabel polysilicon 184 -1929 184 -1929 0 3
rlabel polysilicon 191 -1923 191 -1923 0 1
rlabel polysilicon 191 -1929 191 -1929 0 3
rlabel polysilicon 198 -1923 198 -1923 0 1
rlabel polysilicon 198 -1929 198 -1929 0 3
rlabel polysilicon 205 -1923 205 -1923 0 1
rlabel polysilicon 205 -1929 205 -1929 0 3
rlabel polysilicon 212 -1929 212 -1929 0 3
rlabel polysilicon 219 -1923 219 -1923 0 1
rlabel polysilicon 222 -1923 222 -1923 0 2
rlabel polysilicon 219 -1929 219 -1929 0 3
rlabel polysilicon 226 -1923 226 -1923 0 1
rlabel polysilicon 226 -1929 226 -1929 0 3
rlabel polysilicon 229 -1929 229 -1929 0 4
rlabel polysilicon 233 -1923 233 -1923 0 1
rlabel polysilicon 233 -1929 233 -1929 0 3
rlabel polysilicon 243 -1923 243 -1923 0 2
rlabel polysilicon 240 -1929 240 -1929 0 3
rlabel polysilicon 243 -1929 243 -1929 0 4
rlabel polysilicon 250 -1923 250 -1923 0 2
rlabel polysilicon 247 -1929 247 -1929 0 3
rlabel polysilicon 250 -1929 250 -1929 0 4
rlabel polysilicon 254 -1923 254 -1923 0 1
rlabel polysilicon 254 -1929 254 -1929 0 3
rlabel polysilicon 261 -1923 261 -1923 0 1
rlabel polysilicon 261 -1929 261 -1929 0 3
rlabel polysilicon 268 -1923 268 -1923 0 1
rlabel polysilicon 268 -1929 268 -1929 0 3
rlabel polysilicon 275 -1923 275 -1923 0 1
rlabel polysilicon 275 -1929 275 -1929 0 3
rlabel polysilicon 282 -1923 282 -1923 0 1
rlabel polysilicon 282 -1929 282 -1929 0 3
rlabel polysilicon 289 -1923 289 -1923 0 1
rlabel polysilicon 289 -1929 289 -1929 0 3
rlabel polysilicon 296 -1923 296 -1923 0 1
rlabel polysilicon 296 -1929 296 -1929 0 3
rlabel polysilicon 303 -1923 303 -1923 0 1
rlabel polysilicon 303 -1929 303 -1929 0 3
rlabel polysilicon 310 -1923 310 -1923 0 1
rlabel polysilicon 310 -1929 310 -1929 0 3
rlabel polysilicon 317 -1923 317 -1923 0 1
rlabel polysilicon 317 -1929 317 -1929 0 3
rlabel polysilicon 324 -1923 324 -1923 0 1
rlabel polysilicon 324 -1929 324 -1929 0 3
rlabel polysilicon 331 -1923 331 -1923 0 1
rlabel polysilicon 331 -1929 331 -1929 0 3
rlabel polysilicon 338 -1923 338 -1923 0 1
rlabel polysilicon 341 -1923 341 -1923 0 2
rlabel polysilicon 338 -1929 338 -1929 0 3
rlabel polysilicon 345 -1923 345 -1923 0 1
rlabel polysilicon 345 -1929 345 -1929 0 3
rlabel polysilicon 352 -1923 352 -1923 0 1
rlabel polysilicon 352 -1929 352 -1929 0 3
rlabel polysilicon 359 -1923 359 -1923 0 1
rlabel polysilicon 359 -1929 359 -1929 0 3
rlabel polysilicon 366 -1923 366 -1923 0 1
rlabel polysilicon 366 -1929 366 -1929 0 3
rlabel polysilicon 373 -1923 373 -1923 0 1
rlabel polysilicon 373 -1929 373 -1929 0 3
rlabel polysilicon 380 -1923 380 -1923 0 1
rlabel polysilicon 380 -1929 380 -1929 0 3
rlabel polysilicon 387 -1923 387 -1923 0 1
rlabel polysilicon 387 -1929 387 -1929 0 3
rlabel polysilicon 394 -1923 394 -1923 0 1
rlabel polysilicon 394 -1929 394 -1929 0 3
rlabel polysilicon 401 -1923 401 -1923 0 1
rlabel polysilicon 404 -1923 404 -1923 0 2
rlabel polysilicon 401 -1929 401 -1929 0 3
rlabel polysilicon 404 -1929 404 -1929 0 4
rlabel polysilicon 408 -1923 408 -1923 0 1
rlabel polysilicon 408 -1929 408 -1929 0 3
rlabel polysilicon 415 -1923 415 -1923 0 1
rlabel polysilicon 415 -1929 415 -1929 0 3
rlabel polysilicon 422 -1923 422 -1923 0 1
rlabel polysilicon 422 -1929 422 -1929 0 3
rlabel polysilicon 432 -1923 432 -1923 0 2
rlabel polysilicon 429 -1929 429 -1929 0 3
rlabel polysilicon 432 -1929 432 -1929 0 4
rlabel polysilicon 436 -1923 436 -1923 0 1
rlabel polysilicon 436 -1929 436 -1929 0 3
rlabel polysilicon 443 -1923 443 -1923 0 1
rlabel polysilicon 443 -1929 443 -1929 0 3
rlabel polysilicon 450 -1923 450 -1923 0 1
rlabel polysilicon 450 -1929 450 -1929 0 3
rlabel polysilicon 457 -1923 457 -1923 0 1
rlabel polysilicon 457 -1929 457 -1929 0 3
rlabel polysilicon 464 -1923 464 -1923 0 1
rlabel polysilicon 464 -1929 464 -1929 0 3
rlabel polysilicon 471 -1923 471 -1923 0 1
rlabel polysilicon 471 -1929 471 -1929 0 3
rlabel polysilicon 478 -1923 478 -1923 0 1
rlabel polysilicon 478 -1929 478 -1929 0 3
rlabel polysilicon 485 -1923 485 -1923 0 1
rlabel polysilicon 485 -1929 485 -1929 0 3
rlabel polysilicon 492 -1923 492 -1923 0 1
rlabel polysilicon 492 -1929 492 -1929 0 3
rlabel polysilicon 499 -1923 499 -1923 0 1
rlabel polysilicon 499 -1929 499 -1929 0 3
rlabel polysilicon 506 -1923 506 -1923 0 1
rlabel polysilicon 506 -1929 506 -1929 0 3
rlabel polysilicon 513 -1923 513 -1923 0 1
rlabel polysilicon 513 -1929 513 -1929 0 3
rlabel polysilicon 520 -1923 520 -1923 0 1
rlabel polysilicon 520 -1929 520 -1929 0 3
rlabel polysilicon 527 -1923 527 -1923 0 1
rlabel polysilicon 527 -1929 527 -1929 0 3
rlabel polysilicon 530 -1929 530 -1929 0 4
rlabel polysilicon 534 -1923 534 -1923 0 1
rlabel polysilicon 534 -1929 534 -1929 0 3
rlabel polysilicon 541 -1923 541 -1923 0 1
rlabel polysilicon 541 -1929 541 -1929 0 3
rlabel polysilicon 548 -1923 548 -1923 0 1
rlabel polysilicon 548 -1929 548 -1929 0 3
rlabel polysilicon 555 -1923 555 -1923 0 1
rlabel polysilicon 555 -1929 555 -1929 0 3
rlabel polysilicon 562 -1923 562 -1923 0 1
rlabel polysilicon 562 -1929 562 -1929 0 3
rlabel polysilicon 569 -1923 569 -1923 0 1
rlabel polysilicon 569 -1929 569 -1929 0 3
rlabel polysilicon 576 -1923 576 -1923 0 1
rlabel polysilicon 576 -1929 576 -1929 0 3
rlabel polysilicon 583 -1923 583 -1923 0 1
rlabel polysilicon 583 -1929 583 -1929 0 3
rlabel polysilicon 590 -1923 590 -1923 0 1
rlabel polysilicon 593 -1923 593 -1923 0 2
rlabel polysilicon 590 -1929 590 -1929 0 3
rlabel polysilicon 593 -1929 593 -1929 0 4
rlabel polysilicon 597 -1923 597 -1923 0 1
rlabel polysilicon 597 -1929 597 -1929 0 3
rlabel polysilicon 604 -1923 604 -1923 0 1
rlabel polysilicon 604 -1929 604 -1929 0 3
rlabel polysilicon 611 -1923 611 -1923 0 1
rlabel polysilicon 611 -1929 611 -1929 0 3
rlabel polysilicon 618 -1923 618 -1923 0 1
rlabel polysilicon 621 -1923 621 -1923 0 2
rlabel polysilicon 618 -1929 618 -1929 0 3
rlabel polysilicon 621 -1929 621 -1929 0 4
rlabel polysilicon 625 -1923 625 -1923 0 1
rlabel polysilicon 625 -1929 625 -1929 0 3
rlabel polysilicon 632 -1923 632 -1923 0 1
rlabel polysilicon 632 -1929 632 -1929 0 3
rlabel polysilicon 639 -1923 639 -1923 0 1
rlabel polysilicon 639 -1929 639 -1929 0 3
rlabel polysilicon 646 -1923 646 -1923 0 1
rlabel polysilicon 646 -1929 646 -1929 0 3
rlabel polysilicon 653 -1923 653 -1923 0 1
rlabel polysilicon 656 -1923 656 -1923 0 2
rlabel polysilicon 653 -1929 653 -1929 0 3
rlabel polysilicon 656 -1929 656 -1929 0 4
rlabel polysilicon 660 -1923 660 -1923 0 1
rlabel polysilicon 660 -1929 660 -1929 0 3
rlabel polysilicon 670 -1923 670 -1923 0 2
rlabel polysilicon 667 -1929 667 -1929 0 3
rlabel polysilicon 670 -1929 670 -1929 0 4
rlabel polysilicon 674 -1923 674 -1923 0 1
rlabel polysilicon 674 -1929 674 -1929 0 3
rlabel polysilicon 681 -1923 681 -1923 0 1
rlabel polysilicon 684 -1923 684 -1923 0 2
rlabel polysilicon 681 -1929 681 -1929 0 3
rlabel polysilicon 684 -1929 684 -1929 0 4
rlabel polysilicon 688 -1923 688 -1923 0 1
rlabel polysilicon 688 -1929 688 -1929 0 3
rlabel polysilicon 695 -1923 695 -1923 0 1
rlabel polysilicon 695 -1929 695 -1929 0 3
rlabel polysilicon 702 -1923 702 -1923 0 1
rlabel polysilicon 702 -1929 702 -1929 0 3
rlabel polysilicon 709 -1923 709 -1923 0 1
rlabel polysilicon 709 -1929 709 -1929 0 3
rlabel polysilicon 716 -1923 716 -1923 0 1
rlabel polysilicon 716 -1929 716 -1929 0 3
rlabel polysilicon 723 -1923 723 -1923 0 1
rlabel polysilicon 726 -1923 726 -1923 0 2
rlabel polysilicon 726 -1929 726 -1929 0 4
rlabel polysilicon 730 -1923 730 -1923 0 1
rlabel polysilicon 730 -1929 730 -1929 0 3
rlabel polysilicon 737 -1923 737 -1923 0 1
rlabel polysilicon 737 -1929 737 -1929 0 3
rlabel polysilicon 744 -1923 744 -1923 0 1
rlabel polysilicon 744 -1929 744 -1929 0 3
rlabel polysilicon 751 -1923 751 -1923 0 1
rlabel polysilicon 751 -1929 751 -1929 0 3
rlabel polysilicon 758 -1923 758 -1923 0 1
rlabel polysilicon 758 -1929 758 -1929 0 3
rlabel polysilicon 765 -1923 765 -1923 0 1
rlabel polysilicon 765 -1929 765 -1929 0 3
rlabel polysilicon 772 -1923 772 -1923 0 1
rlabel polysilicon 772 -1929 772 -1929 0 3
rlabel polysilicon 779 -1923 779 -1923 0 1
rlabel polysilicon 779 -1929 779 -1929 0 3
rlabel polysilicon 786 -1923 786 -1923 0 1
rlabel polysilicon 789 -1923 789 -1923 0 2
rlabel polysilicon 786 -1929 786 -1929 0 3
rlabel polysilicon 789 -1929 789 -1929 0 4
rlabel polysilicon 793 -1923 793 -1923 0 1
rlabel polysilicon 793 -1929 793 -1929 0 3
rlabel polysilicon 800 -1923 800 -1923 0 1
rlabel polysilicon 800 -1929 800 -1929 0 3
rlabel polysilicon 807 -1923 807 -1923 0 1
rlabel polysilicon 810 -1923 810 -1923 0 2
rlabel polysilicon 807 -1929 807 -1929 0 3
rlabel polysilicon 810 -1929 810 -1929 0 4
rlabel polysilicon 814 -1923 814 -1923 0 1
rlabel polysilicon 814 -1929 814 -1929 0 3
rlabel polysilicon 821 -1923 821 -1923 0 1
rlabel polysilicon 821 -1929 821 -1929 0 3
rlabel polysilicon 828 -1923 828 -1923 0 1
rlabel polysilicon 831 -1923 831 -1923 0 2
rlabel polysilicon 828 -1929 828 -1929 0 3
rlabel polysilicon 835 -1923 835 -1923 0 1
rlabel polysilicon 835 -1929 835 -1929 0 3
rlabel polysilicon 842 -1923 842 -1923 0 1
rlabel polysilicon 842 -1929 842 -1929 0 3
rlabel polysilicon 849 -1923 849 -1923 0 1
rlabel polysilicon 856 -1923 856 -1923 0 1
rlabel polysilicon 856 -1929 856 -1929 0 3
rlabel polysilicon 863 -1923 863 -1923 0 1
rlabel polysilicon 863 -1929 863 -1929 0 3
rlabel polysilicon 870 -1923 870 -1923 0 1
rlabel polysilicon 870 -1929 870 -1929 0 3
rlabel polysilicon 873 -1929 873 -1929 0 4
rlabel polysilicon 877 -1923 877 -1923 0 1
rlabel polysilicon 877 -1929 877 -1929 0 3
rlabel polysilicon 884 -1923 884 -1923 0 1
rlabel polysilicon 884 -1929 884 -1929 0 3
rlabel polysilicon 891 -1923 891 -1923 0 1
rlabel polysilicon 891 -1929 891 -1929 0 3
rlabel polysilicon 898 -1923 898 -1923 0 1
rlabel polysilicon 898 -1929 898 -1929 0 3
rlabel polysilicon 905 -1923 905 -1923 0 1
rlabel polysilicon 905 -1929 905 -1929 0 3
rlabel polysilicon 912 -1923 912 -1923 0 1
rlabel polysilicon 915 -1923 915 -1923 0 2
rlabel polysilicon 912 -1929 912 -1929 0 3
rlabel polysilicon 915 -1929 915 -1929 0 4
rlabel polysilicon 919 -1923 919 -1923 0 1
rlabel polysilicon 919 -1929 919 -1929 0 3
rlabel polysilicon 926 -1923 926 -1923 0 1
rlabel polysilicon 926 -1929 926 -1929 0 3
rlabel polysilicon 933 -1923 933 -1923 0 1
rlabel polysilicon 933 -1929 933 -1929 0 3
rlabel polysilicon 940 -1923 940 -1923 0 1
rlabel polysilicon 940 -1929 940 -1929 0 3
rlabel polysilicon 947 -1923 947 -1923 0 1
rlabel polysilicon 947 -1929 947 -1929 0 3
rlabel polysilicon 954 -1923 954 -1923 0 1
rlabel polysilicon 954 -1929 954 -1929 0 3
rlabel polysilicon 961 -1923 961 -1923 0 1
rlabel polysilicon 961 -1929 961 -1929 0 3
rlabel polysilicon 968 -1923 968 -1923 0 1
rlabel polysilicon 968 -1929 968 -1929 0 3
rlabel polysilicon 975 -1923 975 -1923 0 1
rlabel polysilicon 975 -1929 975 -1929 0 3
rlabel polysilicon 985 -1923 985 -1923 0 2
rlabel polysilicon 982 -1929 982 -1929 0 3
rlabel polysilicon 985 -1929 985 -1929 0 4
rlabel polysilicon 989 -1923 989 -1923 0 1
rlabel polysilicon 992 -1923 992 -1923 0 2
rlabel polysilicon 989 -1929 989 -1929 0 3
rlabel polysilicon 996 -1923 996 -1923 0 1
rlabel polysilicon 996 -1929 996 -1929 0 3
rlabel polysilicon 1003 -1923 1003 -1923 0 1
rlabel polysilicon 1003 -1929 1003 -1929 0 3
rlabel polysilicon 1010 -1923 1010 -1923 0 1
rlabel polysilicon 1010 -1929 1010 -1929 0 3
rlabel polysilicon 1017 -1923 1017 -1923 0 1
rlabel polysilicon 1017 -1929 1017 -1929 0 3
rlabel polysilicon 1024 -1923 1024 -1923 0 1
rlabel polysilicon 1024 -1929 1024 -1929 0 3
rlabel polysilicon 1031 -1923 1031 -1923 0 1
rlabel polysilicon 1031 -1929 1031 -1929 0 3
rlabel polysilicon 1038 -1923 1038 -1923 0 1
rlabel polysilicon 1038 -1929 1038 -1929 0 3
rlabel polysilicon 1045 -1923 1045 -1923 0 1
rlabel polysilicon 1045 -1929 1045 -1929 0 3
rlabel polysilicon 1052 -1923 1052 -1923 0 1
rlabel polysilicon 1052 -1929 1052 -1929 0 3
rlabel polysilicon 1059 -1923 1059 -1923 0 1
rlabel polysilicon 1059 -1929 1059 -1929 0 3
rlabel polysilicon 1066 -1923 1066 -1923 0 1
rlabel polysilicon 1066 -1929 1066 -1929 0 3
rlabel polysilicon 1073 -1923 1073 -1923 0 1
rlabel polysilicon 1073 -1929 1073 -1929 0 3
rlabel polysilicon 1080 -1923 1080 -1923 0 1
rlabel polysilicon 1080 -1929 1080 -1929 0 3
rlabel polysilicon 1087 -1923 1087 -1923 0 1
rlabel polysilicon 1087 -1929 1087 -1929 0 3
rlabel polysilicon 1094 -1923 1094 -1923 0 1
rlabel polysilicon 1097 -1923 1097 -1923 0 2
rlabel polysilicon 1094 -1929 1094 -1929 0 3
rlabel polysilicon 1097 -1929 1097 -1929 0 4
rlabel polysilicon 1101 -1923 1101 -1923 0 1
rlabel polysilicon 1101 -1929 1101 -1929 0 3
rlabel polysilicon 1108 -1923 1108 -1923 0 1
rlabel polysilicon 1108 -1929 1108 -1929 0 3
rlabel polysilicon 1115 -1923 1115 -1923 0 1
rlabel polysilicon 1115 -1929 1115 -1929 0 3
rlabel polysilicon 1125 -1923 1125 -1923 0 2
rlabel polysilicon 1122 -1929 1122 -1929 0 3
rlabel polysilicon 1125 -1929 1125 -1929 0 4
rlabel polysilicon 1129 -1923 1129 -1923 0 1
rlabel polysilicon 1129 -1929 1129 -1929 0 3
rlabel polysilicon 1136 -1923 1136 -1923 0 1
rlabel polysilicon 1136 -1929 1136 -1929 0 3
rlabel polysilicon 1143 -1923 1143 -1923 0 1
rlabel polysilicon 1143 -1929 1143 -1929 0 3
rlabel polysilicon 1150 -1923 1150 -1923 0 1
rlabel polysilicon 1150 -1929 1150 -1929 0 3
rlabel polysilicon 1157 -1923 1157 -1923 0 1
rlabel polysilicon 1160 -1923 1160 -1923 0 2
rlabel polysilicon 1157 -1929 1157 -1929 0 3
rlabel polysilicon 1160 -1929 1160 -1929 0 4
rlabel polysilicon 1164 -1923 1164 -1923 0 1
rlabel polysilicon 1167 -1923 1167 -1923 0 2
rlabel polysilicon 1164 -1929 1164 -1929 0 3
rlabel polysilicon 1167 -1929 1167 -1929 0 4
rlabel polysilicon 1171 -1923 1171 -1923 0 1
rlabel polysilicon 1171 -1929 1171 -1929 0 3
rlabel polysilicon 1178 -1923 1178 -1923 0 1
rlabel polysilicon 1178 -1929 1178 -1929 0 3
rlabel polysilicon 1185 -1923 1185 -1923 0 1
rlabel polysilicon 1185 -1929 1185 -1929 0 3
rlabel polysilicon 1192 -1923 1192 -1923 0 1
rlabel polysilicon 1192 -1929 1192 -1929 0 3
rlabel polysilicon 1199 -1923 1199 -1923 0 1
rlabel polysilicon 1199 -1929 1199 -1929 0 3
rlabel polysilicon 1206 -1923 1206 -1923 0 1
rlabel polysilicon 1206 -1929 1206 -1929 0 3
rlabel polysilicon 1213 -1923 1213 -1923 0 1
rlabel polysilicon 1213 -1929 1213 -1929 0 3
rlabel polysilicon 1220 -1923 1220 -1923 0 1
rlabel polysilicon 1220 -1929 1220 -1929 0 3
rlabel polysilicon 1227 -1923 1227 -1923 0 1
rlabel polysilicon 1230 -1923 1230 -1923 0 2
rlabel polysilicon 1227 -1929 1227 -1929 0 3
rlabel polysilicon 1230 -1929 1230 -1929 0 4
rlabel polysilicon 1234 -1923 1234 -1923 0 1
rlabel polysilicon 1234 -1929 1234 -1929 0 3
rlabel polysilicon 1241 -1923 1241 -1923 0 1
rlabel polysilicon 1241 -1929 1241 -1929 0 3
rlabel polysilicon 1248 -1923 1248 -1923 0 1
rlabel polysilicon 1248 -1929 1248 -1929 0 3
rlabel polysilicon 1255 -1923 1255 -1923 0 1
rlabel polysilicon 1255 -1929 1255 -1929 0 3
rlabel polysilicon 1262 -1923 1262 -1923 0 1
rlabel polysilicon 1262 -1929 1262 -1929 0 3
rlabel polysilicon 1269 -1923 1269 -1923 0 1
rlabel polysilicon 1269 -1929 1269 -1929 0 3
rlabel polysilicon 1276 -1923 1276 -1923 0 1
rlabel polysilicon 1276 -1929 1276 -1929 0 3
rlabel polysilicon 1283 -1923 1283 -1923 0 1
rlabel polysilicon 1283 -1929 1283 -1929 0 3
rlabel polysilicon 1290 -1923 1290 -1923 0 1
rlabel polysilicon 1290 -1929 1290 -1929 0 3
rlabel polysilicon 1297 -1923 1297 -1923 0 1
rlabel polysilicon 1297 -1929 1297 -1929 0 3
rlabel polysilicon 1304 -1923 1304 -1923 0 1
rlabel polysilicon 1304 -1929 1304 -1929 0 3
rlabel polysilicon 1311 -1923 1311 -1923 0 1
rlabel polysilicon 1311 -1929 1311 -1929 0 3
rlabel polysilicon 1318 -1923 1318 -1923 0 1
rlabel polysilicon 1318 -1929 1318 -1929 0 3
rlabel polysilicon 1325 -1923 1325 -1923 0 1
rlabel polysilicon 1325 -1929 1325 -1929 0 3
rlabel polysilicon 1332 -1923 1332 -1923 0 1
rlabel polysilicon 1332 -1929 1332 -1929 0 3
rlabel polysilicon 1339 -1923 1339 -1923 0 1
rlabel polysilicon 1339 -1929 1339 -1929 0 3
rlabel polysilicon 1346 -1923 1346 -1923 0 1
rlabel polysilicon 1346 -1929 1346 -1929 0 3
rlabel polysilicon 1353 -1923 1353 -1923 0 1
rlabel polysilicon 1353 -1929 1353 -1929 0 3
rlabel polysilicon 1360 -1923 1360 -1923 0 1
rlabel polysilicon 1360 -1929 1360 -1929 0 3
rlabel polysilicon 1367 -1923 1367 -1923 0 1
rlabel polysilicon 1367 -1929 1367 -1929 0 3
rlabel polysilicon 1374 -1923 1374 -1923 0 1
rlabel polysilicon 1374 -1929 1374 -1929 0 3
rlabel polysilicon 1381 -1923 1381 -1923 0 1
rlabel polysilicon 1384 -1923 1384 -1923 0 2
rlabel polysilicon 1381 -1929 1381 -1929 0 3
rlabel polysilicon 1384 -1929 1384 -1929 0 4
rlabel polysilicon 1388 -1923 1388 -1923 0 1
rlabel polysilicon 1388 -1929 1388 -1929 0 3
rlabel polysilicon 1395 -1923 1395 -1923 0 1
rlabel polysilicon 1395 -1929 1395 -1929 0 3
rlabel polysilicon 1402 -1923 1402 -1923 0 1
rlabel polysilicon 1402 -1929 1402 -1929 0 3
rlabel polysilicon 1409 -1923 1409 -1923 0 1
rlabel polysilicon 1409 -1929 1409 -1929 0 3
rlabel polysilicon 1416 -1923 1416 -1923 0 1
rlabel polysilicon 1416 -1929 1416 -1929 0 3
rlabel polysilicon 1423 -1923 1423 -1923 0 1
rlabel polysilicon 1426 -1923 1426 -1923 0 2
rlabel polysilicon 1423 -1929 1423 -1929 0 3
rlabel polysilicon 1430 -1923 1430 -1923 0 1
rlabel polysilicon 1430 -1929 1430 -1929 0 3
rlabel polysilicon 1437 -1923 1437 -1923 0 1
rlabel polysilicon 1437 -1929 1437 -1929 0 3
rlabel polysilicon 1444 -1923 1444 -1923 0 1
rlabel polysilicon 1444 -1929 1444 -1929 0 3
rlabel polysilicon 1451 -1923 1451 -1923 0 1
rlabel polysilicon 1451 -1929 1451 -1929 0 3
rlabel polysilicon 1458 -1923 1458 -1923 0 1
rlabel polysilicon 1458 -1929 1458 -1929 0 3
rlabel polysilicon 1465 -1923 1465 -1923 0 1
rlabel polysilicon 1465 -1929 1465 -1929 0 3
rlabel polysilicon 1472 -1923 1472 -1923 0 1
rlabel polysilicon 1472 -1929 1472 -1929 0 3
rlabel polysilicon 1479 -1923 1479 -1923 0 1
rlabel polysilicon 1479 -1929 1479 -1929 0 3
rlabel polysilicon 1486 -1923 1486 -1923 0 1
rlabel polysilicon 1486 -1929 1486 -1929 0 3
rlabel polysilicon 1493 -1923 1493 -1923 0 1
rlabel polysilicon 1493 -1929 1493 -1929 0 3
rlabel polysilicon 1500 -1923 1500 -1923 0 1
rlabel polysilicon 1500 -1929 1500 -1929 0 3
rlabel polysilicon 1507 -1923 1507 -1923 0 1
rlabel polysilicon 1507 -1929 1507 -1929 0 3
rlabel polysilicon 1514 -1923 1514 -1923 0 1
rlabel polysilicon 1514 -1929 1514 -1929 0 3
rlabel polysilicon 1521 -1923 1521 -1923 0 1
rlabel polysilicon 1521 -1929 1521 -1929 0 3
rlabel polysilicon 1528 -1923 1528 -1923 0 1
rlabel polysilicon 1528 -1929 1528 -1929 0 3
rlabel polysilicon 1535 -1923 1535 -1923 0 1
rlabel polysilicon 1535 -1929 1535 -1929 0 3
rlabel polysilicon 1542 -1923 1542 -1923 0 1
rlabel polysilicon 1542 -1929 1542 -1929 0 3
rlabel polysilicon 1549 -1923 1549 -1923 0 1
rlabel polysilicon 1549 -1929 1549 -1929 0 3
rlabel polysilicon 1556 -1923 1556 -1923 0 1
rlabel polysilicon 1556 -1929 1556 -1929 0 3
rlabel polysilicon 1563 -1923 1563 -1923 0 1
rlabel polysilicon 1563 -1929 1563 -1929 0 3
rlabel polysilicon 1570 -1923 1570 -1923 0 1
rlabel polysilicon 1570 -1929 1570 -1929 0 3
rlabel polysilicon 1577 -1923 1577 -1923 0 1
rlabel polysilicon 1577 -1929 1577 -1929 0 3
rlabel polysilicon 1584 -1923 1584 -1923 0 1
rlabel polysilicon 1584 -1929 1584 -1929 0 3
rlabel polysilicon 1591 -1923 1591 -1923 0 1
rlabel polysilicon 1591 -1929 1591 -1929 0 3
rlabel polysilicon 1598 -1923 1598 -1923 0 1
rlabel polysilicon 1598 -1929 1598 -1929 0 3
rlabel polysilicon 1605 -1923 1605 -1923 0 1
rlabel polysilicon 1605 -1929 1605 -1929 0 3
rlabel polysilicon 1612 -1923 1612 -1923 0 1
rlabel polysilicon 1612 -1929 1612 -1929 0 3
rlabel polysilicon 1619 -1923 1619 -1923 0 1
rlabel polysilicon 1619 -1929 1619 -1929 0 3
rlabel polysilicon 1626 -1923 1626 -1923 0 1
rlabel polysilicon 1626 -1929 1626 -1929 0 3
rlabel polysilicon 1633 -1923 1633 -1923 0 1
rlabel polysilicon 1633 -1929 1633 -1929 0 3
rlabel polysilicon 1640 -1923 1640 -1923 0 1
rlabel polysilicon 1640 -1929 1640 -1929 0 3
rlabel polysilicon 1647 -1923 1647 -1923 0 1
rlabel polysilicon 1647 -1929 1647 -1929 0 3
rlabel polysilicon 1654 -1923 1654 -1923 0 1
rlabel polysilicon 1654 -1929 1654 -1929 0 3
rlabel polysilicon 1661 -1923 1661 -1923 0 1
rlabel polysilicon 1661 -1929 1661 -1929 0 3
rlabel polysilicon 1668 -1923 1668 -1923 0 1
rlabel polysilicon 1668 -1929 1668 -1929 0 3
rlabel polysilicon 1675 -1923 1675 -1923 0 1
rlabel polysilicon 1675 -1929 1675 -1929 0 3
rlabel polysilicon 1682 -1923 1682 -1923 0 1
rlabel polysilicon 1682 -1929 1682 -1929 0 3
rlabel polysilicon 1689 -1923 1689 -1923 0 1
rlabel polysilicon 1689 -1929 1689 -1929 0 3
rlabel polysilicon 1696 -1923 1696 -1923 0 1
rlabel polysilicon 1696 -1929 1696 -1929 0 3
rlabel polysilicon 1703 -1923 1703 -1923 0 1
rlabel polysilicon 1703 -1929 1703 -1929 0 3
rlabel polysilicon 1710 -1923 1710 -1923 0 1
rlabel polysilicon 1710 -1929 1710 -1929 0 3
rlabel polysilicon 1717 -1923 1717 -1923 0 1
rlabel polysilicon 1717 -1929 1717 -1929 0 3
rlabel polysilicon 1724 -1923 1724 -1923 0 1
rlabel polysilicon 1724 -1929 1724 -1929 0 3
rlabel polysilicon 1731 -1923 1731 -1923 0 1
rlabel polysilicon 1731 -1929 1731 -1929 0 3
rlabel polysilicon 1738 -1923 1738 -1923 0 1
rlabel polysilicon 1738 -1929 1738 -1929 0 3
rlabel polysilicon 1745 -1923 1745 -1923 0 1
rlabel polysilicon 1745 -1929 1745 -1929 0 3
rlabel polysilicon 1755 -1923 1755 -1923 0 2
rlabel polysilicon 1759 -1923 1759 -1923 0 1
rlabel polysilicon 1759 -1929 1759 -1929 0 3
rlabel polysilicon 1766 -1923 1766 -1923 0 1
rlabel polysilicon 1766 -1929 1766 -1929 0 3
rlabel polysilicon 1794 -1923 1794 -1923 0 1
rlabel polysilicon 1794 -1929 1794 -1929 0 3
rlabel polysilicon 23 -2050 23 -2050 0 1
rlabel polysilicon 23 -2056 23 -2056 0 3
rlabel polysilicon 37 -2050 37 -2050 0 1
rlabel polysilicon 37 -2056 37 -2056 0 3
rlabel polysilicon 44 -2050 44 -2050 0 1
rlabel polysilicon 44 -2056 44 -2056 0 3
rlabel polysilicon 51 -2050 51 -2050 0 1
rlabel polysilicon 51 -2056 51 -2056 0 3
rlabel polysilicon 58 -2050 58 -2050 0 1
rlabel polysilicon 58 -2056 58 -2056 0 3
rlabel polysilicon 65 -2050 65 -2050 0 1
rlabel polysilicon 65 -2056 65 -2056 0 3
rlabel polysilicon 72 -2050 72 -2050 0 1
rlabel polysilicon 72 -2056 72 -2056 0 3
rlabel polysilicon 79 -2050 79 -2050 0 1
rlabel polysilicon 79 -2056 79 -2056 0 3
rlabel polysilicon 86 -2050 86 -2050 0 1
rlabel polysilicon 86 -2056 86 -2056 0 3
rlabel polysilicon 93 -2050 93 -2050 0 1
rlabel polysilicon 93 -2056 93 -2056 0 3
rlabel polysilicon 100 -2050 100 -2050 0 1
rlabel polysilicon 100 -2056 100 -2056 0 3
rlabel polysilicon 107 -2050 107 -2050 0 1
rlabel polysilicon 110 -2050 110 -2050 0 2
rlabel polysilicon 107 -2056 107 -2056 0 3
rlabel polysilicon 114 -2050 114 -2050 0 1
rlabel polysilicon 117 -2050 117 -2050 0 2
rlabel polysilicon 114 -2056 114 -2056 0 3
rlabel polysilicon 121 -2050 121 -2050 0 1
rlabel polysilicon 121 -2056 121 -2056 0 3
rlabel polysilicon 128 -2050 128 -2050 0 1
rlabel polysilicon 131 -2050 131 -2050 0 2
rlabel polysilicon 128 -2056 128 -2056 0 3
rlabel polysilicon 135 -2050 135 -2050 0 1
rlabel polysilicon 138 -2050 138 -2050 0 2
rlabel polysilicon 142 -2050 142 -2050 0 1
rlabel polysilicon 142 -2056 142 -2056 0 3
rlabel polysilicon 149 -2050 149 -2050 0 1
rlabel polysilicon 149 -2056 149 -2056 0 3
rlabel polysilicon 156 -2050 156 -2050 0 1
rlabel polysilicon 159 -2050 159 -2050 0 2
rlabel polysilicon 156 -2056 156 -2056 0 3
rlabel polysilicon 163 -2050 163 -2050 0 1
rlabel polysilicon 166 -2050 166 -2050 0 2
rlabel polysilicon 163 -2056 163 -2056 0 3
rlabel polysilicon 166 -2056 166 -2056 0 4
rlabel polysilicon 170 -2050 170 -2050 0 1
rlabel polysilicon 170 -2056 170 -2056 0 3
rlabel polysilicon 177 -2050 177 -2050 0 1
rlabel polysilicon 177 -2056 177 -2056 0 3
rlabel polysilicon 184 -2050 184 -2050 0 1
rlabel polysilicon 184 -2056 184 -2056 0 3
rlabel polysilicon 191 -2050 191 -2050 0 1
rlabel polysilicon 191 -2056 191 -2056 0 3
rlabel polysilicon 198 -2050 198 -2050 0 1
rlabel polysilicon 198 -2056 198 -2056 0 3
rlabel polysilicon 205 -2050 205 -2050 0 1
rlabel polysilicon 208 -2050 208 -2050 0 2
rlabel polysilicon 205 -2056 205 -2056 0 3
rlabel polysilicon 208 -2056 208 -2056 0 4
rlabel polysilicon 212 -2050 212 -2050 0 1
rlabel polysilicon 212 -2056 212 -2056 0 3
rlabel polysilicon 219 -2050 219 -2050 0 1
rlabel polysilicon 219 -2056 219 -2056 0 3
rlabel polysilicon 226 -2050 226 -2050 0 1
rlabel polysilicon 226 -2056 226 -2056 0 3
rlabel polysilicon 233 -2050 233 -2050 0 1
rlabel polysilicon 233 -2056 233 -2056 0 3
rlabel polysilicon 240 -2050 240 -2050 0 1
rlabel polysilicon 240 -2056 240 -2056 0 3
rlabel polysilicon 247 -2050 247 -2050 0 1
rlabel polysilicon 247 -2056 247 -2056 0 3
rlabel polysilicon 254 -2050 254 -2050 0 1
rlabel polysilicon 254 -2056 254 -2056 0 3
rlabel polysilicon 261 -2050 261 -2050 0 1
rlabel polysilicon 261 -2056 261 -2056 0 3
rlabel polysilicon 268 -2050 268 -2050 0 1
rlabel polysilicon 268 -2056 268 -2056 0 3
rlabel polysilicon 275 -2050 275 -2050 0 1
rlabel polysilicon 275 -2056 275 -2056 0 3
rlabel polysilicon 282 -2050 282 -2050 0 1
rlabel polysilicon 282 -2056 282 -2056 0 3
rlabel polysilicon 289 -2050 289 -2050 0 1
rlabel polysilicon 289 -2056 289 -2056 0 3
rlabel polysilicon 296 -2050 296 -2050 0 1
rlabel polysilicon 296 -2056 296 -2056 0 3
rlabel polysilicon 303 -2050 303 -2050 0 1
rlabel polysilicon 303 -2056 303 -2056 0 3
rlabel polysilicon 310 -2050 310 -2050 0 1
rlabel polysilicon 310 -2056 310 -2056 0 3
rlabel polysilicon 317 -2050 317 -2050 0 1
rlabel polysilicon 317 -2056 317 -2056 0 3
rlabel polysilicon 324 -2050 324 -2050 0 1
rlabel polysilicon 324 -2056 324 -2056 0 3
rlabel polysilicon 331 -2050 331 -2050 0 1
rlabel polysilicon 331 -2056 331 -2056 0 3
rlabel polysilicon 338 -2050 338 -2050 0 1
rlabel polysilicon 338 -2056 338 -2056 0 3
rlabel polysilicon 345 -2050 345 -2050 0 1
rlabel polysilicon 345 -2056 345 -2056 0 3
rlabel polysilicon 352 -2050 352 -2050 0 1
rlabel polysilicon 352 -2056 352 -2056 0 3
rlabel polysilicon 359 -2050 359 -2050 0 1
rlabel polysilicon 359 -2056 359 -2056 0 3
rlabel polysilicon 369 -2050 369 -2050 0 2
rlabel polysilicon 366 -2056 366 -2056 0 3
rlabel polysilicon 369 -2056 369 -2056 0 4
rlabel polysilicon 373 -2050 373 -2050 0 1
rlabel polysilicon 373 -2056 373 -2056 0 3
rlabel polysilicon 380 -2050 380 -2050 0 1
rlabel polysilicon 380 -2056 380 -2056 0 3
rlabel polysilicon 387 -2050 387 -2050 0 1
rlabel polysilicon 387 -2056 387 -2056 0 3
rlabel polysilicon 394 -2050 394 -2050 0 1
rlabel polysilicon 394 -2056 394 -2056 0 3
rlabel polysilicon 401 -2050 401 -2050 0 1
rlabel polysilicon 401 -2056 401 -2056 0 3
rlabel polysilicon 408 -2050 408 -2050 0 1
rlabel polysilicon 408 -2056 408 -2056 0 3
rlabel polysilicon 415 -2050 415 -2050 0 1
rlabel polysilicon 415 -2056 415 -2056 0 3
rlabel polysilicon 422 -2050 422 -2050 0 1
rlabel polysilicon 422 -2056 422 -2056 0 3
rlabel polysilicon 429 -2050 429 -2050 0 1
rlabel polysilicon 429 -2056 429 -2056 0 3
rlabel polysilicon 436 -2050 436 -2050 0 1
rlabel polysilicon 436 -2056 436 -2056 0 3
rlabel polysilicon 443 -2050 443 -2050 0 1
rlabel polysilicon 443 -2056 443 -2056 0 3
rlabel polysilicon 450 -2050 450 -2050 0 1
rlabel polysilicon 450 -2056 450 -2056 0 3
rlabel polysilicon 457 -2050 457 -2050 0 1
rlabel polysilicon 457 -2056 457 -2056 0 3
rlabel polysilicon 464 -2050 464 -2050 0 1
rlabel polysilicon 464 -2056 464 -2056 0 3
rlabel polysilicon 471 -2050 471 -2050 0 1
rlabel polysilicon 471 -2056 471 -2056 0 3
rlabel polysilicon 478 -2050 478 -2050 0 1
rlabel polysilicon 478 -2056 478 -2056 0 3
rlabel polysilicon 485 -2050 485 -2050 0 1
rlabel polysilicon 485 -2056 485 -2056 0 3
rlabel polysilicon 492 -2050 492 -2050 0 1
rlabel polysilicon 492 -2056 492 -2056 0 3
rlabel polysilicon 499 -2050 499 -2050 0 1
rlabel polysilicon 499 -2056 499 -2056 0 3
rlabel polysilicon 506 -2050 506 -2050 0 1
rlabel polysilicon 506 -2056 506 -2056 0 3
rlabel polysilicon 513 -2050 513 -2050 0 1
rlabel polysilicon 513 -2056 513 -2056 0 3
rlabel polysilicon 520 -2050 520 -2050 0 1
rlabel polysilicon 520 -2056 520 -2056 0 3
rlabel polysilicon 530 -2050 530 -2050 0 2
rlabel polysilicon 530 -2056 530 -2056 0 4
rlabel polysilicon 534 -2050 534 -2050 0 1
rlabel polysilicon 534 -2056 534 -2056 0 3
rlabel polysilicon 541 -2050 541 -2050 0 1
rlabel polysilicon 541 -2056 541 -2056 0 3
rlabel polysilicon 548 -2050 548 -2050 0 1
rlabel polysilicon 548 -2056 548 -2056 0 3
rlabel polysilicon 555 -2050 555 -2050 0 1
rlabel polysilicon 555 -2056 555 -2056 0 3
rlabel polysilicon 562 -2050 562 -2050 0 1
rlabel polysilicon 562 -2056 562 -2056 0 3
rlabel polysilicon 569 -2050 569 -2050 0 1
rlabel polysilicon 569 -2056 569 -2056 0 3
rlabel polysilicon 576 -2050 576 -2050 0 1
rlabel polysilicon 576 -2056 576 -2056 0 3
rlabel polysilicon 583 -2050 583 -2050 0 1
rlabel polysilicon 583 -2056 583 -2056 0 3
rlabel polysilicon 590 -2050 590 -2050 0 1
rlabel polysilicon 593 -2050 593 -2050 0 2
rlabel polysilicon 593 -2056 593 -2056 0 4
rlabel polysilicon 597 -2050 597 -2050 0 1
rlabel polysilicon 600 -2050 600 -2050 0 2
rlabel polysilicon 600 -2056 600 -2056 0 4
rlabel polysilicon 604 -2050 604 -2050 0 1
rlabel polysilicon 607 -2050 607 -2050 0 2
rlabel polysilicon 607 -2056 607 -2056 0 4
rlabel polysilicon 611 -2050 611 -2050 0 1
rlabel polysilicon 611 -2056 611 -2056 0 3
rlabel polysilicon 618 -2050 618 -2050 0 1
rlabel polysilicon 621 -2050 621 -2050 0 2
rlabel polysilicon 618 -2056 618 -2056 0 3
rlabel polysilicon 621 -2056 621 -2056 0 4
rlabel polysilicon 625 -2050 625 -2050 0 1
rlabel polysilicon 625 -2056 625 -2056 0 3
rlabel polysilicon 632 -2050 632 -2050 0 1
rlabel polysilicon 635 -2050 635 -2050 0 2
rlabel polysilicon 632 -2056 632 -2056 0 3
rlabel polysilicon 635 -2056 635 -2056 0 4
rlabel polysilicon 639 -2050 639 -2050 0 1
rlabel polysilicon 639 -2056 639 -2056 0 3
rlabel polysilicon 646 -2050 646 -2050 0 1
rlabel polysilicon 646 -2056 646 -2056 0 3
rlabel polysilicon 653 -2050 653 -2050 0 1
rlabel polysilicon 653 -2056 653 -2056 0 3
rlabel polysilicon 660 -2050 660 -2050 0 1
rlabel polysilicon 663 -2050 663 -2050 0 2
rlabel polysilicon 660 -2056 660 -2056 0 3
rlabel polysilicon 663 -2056 663 -2056 0 4
rlabel polysilicon 667 -2050 667 -2050 0 1
rlabel polysilicon 670 -2050 670 -2050 0 2
rlabel polysilicon 667 -2056 667 -2056 0 3
rlabel polysilicon 670 -2056 670 -2056 0 4
rlabel polysilicon 674 -2050 674 -2050 0 1
rlabel polysilicon 674 -2056 674 -2056 0 3
rlabel polysilicon 681 -2050 681 -2050 0 1
rlabel polysilicon 681 -2056 681 -2056 0 3
rlabel polysilicon 688 -2050 688 -2050 0 1
rlabel polysilicon 691 -2050 691 -2050 0 2
rlabel polysilicon 688 -2056 688 -2056 0 3
rlabel polysilicon 691 -2056 691 -2056 0 4
rlabel polysilicon 695 -2050 695 -2050 0 1
rlabel polysilicon 695 -2056 695 -2056 0 3
rlabel polysilicon 702 -2050 702 -2050 0 1
rlabel polysilicon 702 -2056 702 -2056 0 3
rlabel polysilicon 709 -2050 709 -2050 0 1
rlabel polysilicon 709 -2056 709 -2056 0 3
rlabel polysilicon 716 -2050 716 -2050 0 1
rlabel polysilicon 716 -2056 716 -2056 0 3
rlabel polysilicon 723 -2050 723 -2050 0 1
rlabel polysilicon 723 -2056 723 -2056 0 3
rlabel polysilicon 730 -2050 730 -2050 0 1
rlabel polysilicon 730 -2056 730 -2056 0 3
rlabel polysilicon 737 -2050 737 -2050 0 1
rlabel polysilicon 737 -2056 737 -2056 0 3
rlabel polysilicon 744 -2050 744 -2050 0 1
rlabel polysilicon 744 -2056 744 -2056 0 3
rlabel polysilicon 751 -2050 751 -2050 0 1
rlabel polysilicon 754 -2050 754 -2050 0 2
rlabel polysilicon 751 -2056 751 -2056 0 3
rlabel polysilicon 754 -2056 754 -2056 0 4
rlabel polysilicon 758 -2050 758 -2050 0 1
rlabel polysilicon 758 -2056 758 -2056 0 3
rlabel polysilicon 765 -2050 765 -2050 0 1
rlabel polysilicon 768 -2050 768 -2050 0 2
rlabel polysilicon 765 -2056 765 -2056 0 3
rlabel polysilicon 772 -2050 772 -2050 0 1
rlabel polysilicon 772 -2056 772 -2056 0 3
rlabel polysilicon 782 -2050 782 -2050 0 2
rlabel polysilicon 779 -2056 779 -2056 0 3
rlabel polysilicon 782 -2056 782 -2056 0 4
rlabel polysilicon 786 -2050 786 -2050 0 1
rlabel polysilicon 786 -2056 786 -2056 0 3
rlabel polysilicon 793 -2050 793 -2050 0 1
rlabel polysilicon 793 -2056 793 -2056 0 3
rlabel polysilicon 800 -2050 800 -2050 0 1
rlabel polysilicon 803 -2050 803 -2050 0 2
rlabel polysilicon 800 -2056 800 -2056 0 3
rlabel polysilicon 803 -2056 803 -2056 0 4
rlabel polysilicon 807 -2050 807 -2050 0 1
rlabel polysilicon 807 -2056 807 -2056 0 3
rlabel polysilicon 814 -2050 814 -2050 0 1
rlabel polysilicon 817 -2050 817 -2050 0 2
rlabel polysilicon 814 -2056 814 -2056 0 3
rlabel polysilicon 817 -2056 817 -2056 0 4
rlabel polysilicon 821 -2050 821 -2050 0 1
rlabel polysilicon 821 -2056 821 -2056 0 3
rlabel polysilicon 828 -2050 828 -2050 0 1
rlabel polysilicon 828 -2056 828 -2056 0 3
rlabel polysilicon 835 -2050 835 -2050 0 1
rlabel polysilicon 835 -2056 835 -2056 0 3
rlabel polysilicon 842 -2050 842 -2050 0 1
rlabel polysilicon 842 -2056 842 -2056 0 3
rlabel polysilicon 849 -2050 849 -2050 0 1
rlabel polysilicon 849 -2056 849 -2056 0 3
rlabel polysilicon 856 -2050 856 -2050 0 1
rlabel polysilicon 856 -2056 856 -2056 0 3
rlabel polysilicon 863 -2050 863 -2050 0 1
rlabel polysilicon 863 -2056 863 -2056 0 3
rlabel polysilicon 870 -2050 870 -2050 0 1
rlabel polysilicon 870 -2056 870 -2056 0 3
rlabel polysilicon 877 -2050 877 -2050 0 1
rlabel polysilicon 877 -2056 877 -2056 0 3
rlabel polysilicon 884 -2050 884 -2050 0 1
rlabel polysilicon 884 -2056 884 -2056 0 3
rlabel polysilicon 891 -2050 891 -2050 0 1
rlabel polysilicon 891 -2056 891 -2056 0 3
rlabel polysilicon 898 -2050 898 -2050 0 1
rlabel polysilicon 898 -2056 898 -2056 0 3
rlabel polysilicon 905 -2050 905 -2050 0 1
rlabel polysilicon 908 -2050 908 -2050 0 2
rlabel polysilicon 905 -2056 905 -2056 0 3
rlabel polysilicon 908 -2056 908 -2056 0 4
rlabel polysilicon 912 -2050 912 -2050 0 1
rlabel polysilicon 912 -2056 912 -2056 0 3
rlabel polysilicon 919 -2050 919 -2050 0 1
rlabel polysilicon 919 -2056 919 -2056 0 3
rlabel polysilicon 926 -2050 926 -2050 0 1
rlabel polysilicon 929 -2050 929 -2050 0 2
rlabel polysilicon 926 -2056 926 -2056 0 3
rlabel polysilicon 933 -2050 933 -2050 0 1
rlabel polysilicon 936 -2050 936 -2050 0 2
rlabel polysilicon 933 -2056 933 -2056 0 3
rlabel polysilicon 936 -2056 936 -2056 0 4
rlabel polysilicon 940 -2050 940 -2050 0 1
rlabel polysilicon 950 -2050 950 -2050 0 2
rlabel polysilicon 947 -2056 947 -2056 0 3
rlabel polysilicon 950 -2056 950 -2056 0 4
rlabel polysilicon 954 -2050 954 -2050 0 1
rlabel polysilicon 954 -2056 954 -2056 0 3
rlabel polysilicon 961 -2050 961 -2050 0 1
rlabel polysilicon 961 -2056 961 -2056 0 3
rlabel polysilicon 968 -2050 968 -2050 0 1
rlabel polysilicon 968 -2056 968 -2056 0 3
rlabel polysilicon 975 -2050 975 -2050 0 1
rlabel polysilicon 975 -2056 975 -2056 0 3
rlabel polysilicon 985 -2050 985 -2050 0 2
rlabel polysilicon 982 -2056 982 -2056 0 3
rlabel polysilicon 985 -2056 985 -2056 0 4
rlabel polysilicon 989 -2050 989 -2050 0 1
rlabel polysilicon 989 -2056 989 -2056 0 3
rlabel polysilicon 996 -2050 996 -2050 0 1
rlabel polysilicon 996 -2056 996 -2056 0 3
rlabel polysilicon 1003 -2050 1003 -2050 0 1
rlabel polysilicon 1003 -2056 1003 -2056 0 3
rlabel polysilicon 1010 -2050 1010 -2050 0 1
rlabel polysilicon 1010 -2056 1010 -2056 0 3
rlabel polysilicon 1017 -2050 1017 -2050 0 1
rlabel polysilicon 1020 -2050 1020 -2050 0 2
rlabel polysilicon 1017 -2056 1017 -2056 0 3
rlabel polysilicon 1020 -2056 1020 -2056 0 4
rlabel polysilicon 1024 -2050 1024 -2050 0 1
rlabel polysilicon 1024 -2056 1024 -2056 0 3
rlabel polysilicon 1031 -2050 1031 -2050 0 1
rlabel polysilicon 1031 -2056 1031 -2056 0 3
rlabel polysilicon 1038 -2050 1038 -2050 0 1
rlabel polysilicon 1038 -2056 1038 -2056 0 3
rlabel polysilicon 1045 -2050 1045 -2050 0 1
rlabel polysilicon 1045 -2056 1045 -2056 0 3
rlabel polysilicon 1052 -2050 1052 -2050 0 1
rlabel polysilicon 1052 -2056 1052 -2056 0 3
rlabel polysilicon 1059 -2050 1059 -2050 0 1
rlabel polysilicon 1059 -2056 1059 -2056 0 3
rlabel polysilicon 1066 -2050 1066 -2050 0 1
rlabel polysilicon 1066 -2056 1066 -2056 0 3
rlabel polysilicon 1073 -2050 1073 -2050 0 1
rlabel polysilicon 1073 -2056 1073 -2056 0 3
rlabel polysilicon 1080 -2050 1080 -2050 0 1
rlabel polysilicon 1080 -2056 1080 -2056 0 3
rlabel polysilicon 1087 -2050 1087 -2050 0 1
rlabel polysilicon 1087 -2056 1087 -2056 0 3
rlabel polysilicon 1090 -2056 1090 -2056 0 4
rlabel polysilicon 1094 -2050 1094 -2050 0 1
rlabel polysilicon 1094 -2056 1094 -2056 0 3
rlabel polysilicon 1101 -2050 1101 -2050 0 1
rlabel polysilicon 1101 -2056 1101 -2056 0 3
rlabel polysilicon 1108 -2050 1108 -2050 0 1
rlabel polysilicon 1108 -2056 1108 -2056 0 3
rlabel polysilicon 1115 -2050 1115 -2050 0 1
rlabel polysilicon 1115 -2056 1115 -2056 0 3
rlabel polysilicon 1122 -2050 1122 -2050 0 1
rlabel polysilicon 1122 -2056 1122 -2056 0 3
rlabel polysilicon 1129 -2050 1129 -2050 0 1
rlabel polysilicon 1129 -2056 1129 -2056 0 3
rlabel polysilicon 1136 -2050 1136 -2050 0 1
rlabel polysilicon 1136 -2056 1136 -2056 0 3
rlabel polysilicon 1143 -2050 1143 -2050 0 1
rlabel polysilicon 1143 -2056 1143 -2056 0 3
rlabel polysilicon 1150 -2050 1150 -2050 0 1
rlabel polysilicon 1150 -2056 1150 -2056 0 3
rlabel polysilicon 1157 -2050 1157 -2050 0 1
rlabel polysilicon 1157 -2056 1157 -2056 0 3
rlabel polysilicon 1164 -2050 1164 -2050 0 1
rlabel polysilicon 1164 -2056 1164 -2056 0 3
rlabel polysilicon 1171 -2050 1171 -2050 0 1
rlabel polysilicon 1171 -2056 1171 -2056 0 3
rlabel polysilicon 1178 -2050 1178 -2050 0 1
rlabel polysilicon 1178 -2056 1178 -2056 0 3
rlabel polysilicon 1185 -2050 1185 -2050 0 1
rlabel polysilicon 1185 -2056 1185 -2056 0 3
rlabel polysilicon 1192 -2050 1192 -2050 0 1
rlabel polysilicon 1192 -2056 1192 -2056 0 3
rlabel polysilicon 1199 -2050 1199 -2050 0 1
rlabel polysilicon 1199 -2056 1199 -2056 0 3
rlabel polysilicon 1206 -2050 1206 -2050 0 1
rlabel polysilicon 1206 -2056 1206 -2056 0 3
rlabel polysilicon 1213 -2050 1213 -2050 0 1
rlabel polysilicon 1213 -2056 1213 -2056 0 3
rlabel polysilicon 1220 -2050 1220 -2050 0 1
rlabel polysilicon 1220 -2056 1220 -2056 0 3
rlabel polysilicon 1227 -2050 1227 -2050 0 1
rlabel polysilicon 1227 -2056 1227 -2056 0 3
rlabel polysilicon 1234 -2050 1234 -2050 0 1
rlabel polysilicon 1234 -2056 1234 -2056 0 3
rlabel polysilicon 1241 -2050 1241 -2050 0 1
rlabel polysilicon 1241 -2056 1241 -2056 0 3
rlabel polysilicon 1248 -2050 1248 -2050 0 1
rlabel polysilicon 1248 -2056 1248 -2056 0 3
rlabel polysilicon 1255 -2050 1255 -2050 0 1
rlabel polysilicon 1258 -2050 1258 -2050 0 2
rlabel polysilicon 1255 -2056 1255 -2056 0 3
rlabel polysilicon 1258 -2056 1258 -2056 0 4
rlabel polysilicon 1262 -2050 1262 -2050 0 1
rlabel polysilicon 1262 -2056 1262 -2056 0 3
rlabel polysilicon 1269 -2050 1269 -2050 0 1
rlabel polysilicon 1269 -2056 1269 -2056 0 3
rlabel polysilicon 1276 -2050 1276 -2050 0 1
rlabel polysilicon 1276 -2056 1276 -2056 0 3
rlabel polysilicon 1283 -2050 1283 -2050 0 1
rlabel polysilicon 1283 -2056 1283 -2056 0 3
rlabel polysilicon 1290 -2050 1290 -2050 0 1
rlabel polysilicon 1290 -2056 1290 -2056 0 3
rlabel polysilicon 1297 -2050 1297 -2050 0 1
rlabel polysilicon 1297 -2056 1297 -2056 0 3
rlabel polysilicon 1304 -2050 1304 -2050 0 1
rlabel polysilicon 1304 -2056 1304 -2056 0 3
rlabel polysilicon 1311 -2050 1311 -2050 0 1
rlabel polysilicon 1311 -2056 1311 -2056 0 3
rlabel polysilicon 1318 -2050 1318 -2050 0 1
rlabel polysilicon 1318 -2056 1318 -2056 0 3
rlabel polysilicon 1325 -2050 1325 -2050 0 1
rlabel polysilicon 1325 -2056 1325 -2056 0 3
rlabel polysilicon 1332 -2050 1332 -2050 0 1
rlabel polysilicon 1332 -2056 1332 -2056 0 3
rlabel polysilicon 1339 -2050 1339 -2050 0 1
rlabel polysilicon 1339 -2056 1339 -2056 0 3
rlabel polysilicon 1346 -2050 1346 -2050 0 1
rlabel polysilicon 1346 -2056 1346 -2056 0 3
rlabel polysilicon 1353 -2050 1353 -2050 0 1
rlabel polysilicon 1353 -2056 1353 -2056 0 3
rlabel polysilicon 1360 -2050 1360 -2050 0 1
rlabel polysilicon 1360 -2056 1360 -2056 0 3
rlabel polysilicon 1367 -2050 1367 -2050 0 1
rlabel polysilicon 1367 -2056 1367 -2056 0 3
rlabel polysilicon 1374 -2050 1374 -2050 0 1
rlabel polysilicon 1374 -2056 1374 -2056 0 3
rlabel polysilicon 1381 -2050 1381 -2050 0 1
rlabel polysilicon 1381 -2056 1381 -2056 0 3
rlabel polysilicon 1388 -2050 1388 -2050 0 1
rlabel polysilicon 1388 -2056 1388 -2056 0 3
rlabel polysilicon 1395 -2050 1395 -2050 0 1
rlabel polysilicon 1395 -2056 1395 -2056 0 3
rlabel polysilicon 1402 -2050 1402 -2050 0 1
rlabel polysilicon 1402 -2056 1402 -2056 0 3
rlabel polysilicon 1409 -2050 1409 -2050 0 1
rlabel polysilicon 1409 -2056 1409 -2056 0 3
rlabel polysilicon 1416 -2050 1416 -2050 0 1
rlabel polysilicon 1416 -2056 1416 -2056 0 3
rlabel polysilicon 1423 -2050 1423 -2050 0 1
rlabel polysilicon 1423 -2056 1423 -2056 0 3
rlabel polysilicon 1430 -2050 1430 -2050 0 1
rlabel polysilicon 1430 -2056 1430 -2056 0 3
rlabel polysilicon 1437 -2050 1437 -2050 0 1
rlabel polysilicon 1437 -2056 1437 -2056 0 3
rlabel polysilicon 1444 -2050 1444 -2050 0 1
rlabel polysilicon 1444 -2056 1444 -2056 0 3
rlabel polysilicon 1451 -2056 1451 -2056 0 3
rlabel polysilicon 1458 -2050 1458 -2050 0 1
rlabel polysilicon 1458 -2056 1458 -2056 0 3
rlabel polysilicon 1465 -2050 1465 -2050 0 1
rlabel polysilicon 1465 -2056 1465 -2056 0 3
rlabel polysilicon 1472 -2050 1472 -2050 0 1
rlabel polysilicon 1472 -2056 1472 -2056 0 3
rlabel polysilicon 1479 -2050 1479 -2050 0 1
rlabel polysilicon 1479 -2056 1479 -2056 0 3
rlabel polysilicon 1486 -2050 1486 -2050 0 1
rlabel polysilicon 1486 -2056 1486 -2056 0 3
rlabel polysilicon 1493 -2050 1493 -2050 0 1
rlabel polysilicon 1493 -2056 1493 -2056 0 3
rlabel polysilicon 1500 -2050 1500 -2050 0 1
rlabel polysilicon 1500 -2056 1500 -2056 0 3
rlabel polysilicon 1507 -2050 1507 -2050 0 1
rlabel polysilicon 1507 -2056 1507 -2056 0 3
rlabel polysilicon 1514 -2050 1514 -2050 0 1
rlabel polysilicon 1514 -2056 1514 -2056 0 3
rlabel polysilicon 1521 -2050 1521 -2050 0 1
rlabel polysilicon 1521 -2056 1521 -2056 0 3
rlabel polysilicon 1528 -2050 1528 -2050 0 1
rlabel polysilicon 1528 -2056 1528 -2056 0 3
rlabel polysilicon 1535 -2050 1535 -2050 0 1
rlabel polysilicon 1535 -2056 1535 -2056 0 3
rlabel polysilicon 1542 -2050 1542 -2050 0 1
rlabel polysilicon 1542 -2056 1542 -2056 0 3
rlabel polysilicon 1549 -2050 1549 -2050 0 1
rlabel polysilicon 1549 -2056 1549 -2056 0 3
rlabel polysilicon 1556 -2050 1556 -2050 0 1
rlabel polysilicon 1556 -2056 1556 -2056 0 3
rlabel polysilicon 1563 -2050 1563 -2050 0 1
rlabel polysilicon 1563 -2056 1563 -2056 0 3
rlabel polysilicon 1570 -2050 1570 -2050 0 1
rlabel polysilicon 1570 -2056 1570 -2056 0 3
rlabel polysilicon 1577 -2050 1577 -2050 0 1
rlabel polysilicon 1577 -2056 1577 -2056 0 3
rlabel polysilicon 1584 -2050 1584 -2050 0 1
rlabel polysilicon 1584 -2056 1584 -2056 0 3
rlabel polysilicon 1591 -2050 1591 -2050 0 1
rlabel polysilicon 1591 -2056 1591 -2056 0 3
rlabel polysilicon 1598 -2050 1598 -2050 0 1
rlabel polysilicon 1598 -2056 1598 -2056 0 3
rlabel polysilicon 1605 -2050 1605 -2050 0 1
rlabel polysilicon 1605 -2056 1605 -2056 0 3
rlabel polysilicon 1612 -2050 1612 -2050 0 1
rlabel polysilicon 1612 -2056 1612 -2056 0 3
rlabel polysilicon 1619 -2050 1619 -2050 0 1
rlabel polysilicon 1619 -2056 1619 -2056 0 3
rlabel polysilicon 1626 -2050 1626 -2050 0 1
rlabel polysilicon 1626 -2056 1626 -2056 0 3
rlabel polysilicon 1629 -2056 1629 -2056 0 4
rlabel polysilicon 1633 -2050 1633 -2050 0 1
rlabel polysilicon 1633 -2056 1633 -2056 0 3
rlabel polysilicon 1640 -2050 1640 -2050 0 1
rlabel polysilicon 1640 -2056 1640 -2056 0 3
rlabel polysilicon 1647 -2050 1647 -2050 0 1
rlabel polysilicon 1647 -2056 1647 -2056 0 3
rlabel polysilicon 1654 -2050 1654 -2050 0 1
rlabel polysilicon 1654 -2056 1654 -2056 0 3
rlabel polysilicon 1661 -2050 1661 -2050 0 1
rlabel polysilicon 1661 -2056 1661 -2056 0 3
rlabel polysilicon 1668 -2050 1668 -2050 0 1
rlabel polysilicon 1668 -2056 1668 -2056 0 3
rlabel polysilicon 1675 -2050 1675 -2050 0 1
rlabel polysilicon 1675 -2056 1675 -2056 0 3
rlabel polysilicon 1682 -2050 1682 -2050 0 1
rlabel polysilicon 1682 -2056 1682 -2056 0 3
rlabel polysilicon 1689 -2050 1689 -2050 0 1
rlabel polysilicon 1689 -2056 1689 -2056 0 3
rlabel polysilicon 1696 -2050 1696 -2050 0 1
rlabel polysilicon 1696 -2056 1696 -2056 0 3
rlabel polysilicon 1703 -2050 1703 -2050 0 1
rlabel polysilicon 1703 -2056 1703 -2056 0 3
rlabel polysilicon 1710 -2050 1710 -2050 0 1
rlabel polysilicon 1710 -2056 1710 -2056 0 3
rlabel polysilicon 1717 -2050 1717 -2050 0 1
rlabel polysilicon 1717 -2056 1717 -2056 0 3
rlabel polysilicon 1724 -2050 1724 -2050 0 1
rlabel polysilicon 1724 -2056 1724 -2056 0 3
rlabel polysilicon 1731 -2050 1731 -2050 0 1
rlabel polysilicon 1731 -2056 1731 -2056 0 3
rlabel polysilicon 1738 -2050 1738 -2050 0 1
rlabel polysilicon 1738 -2056 1738 -2056 0 3
rlabel polysilicon 1745 -2050 1745 -2050 0 1
rlabel polysilicon 1745 -2056 1745 -2056 0 3
rlabel polysilicon 1748 -2056 1748 -2056 0 4
rlabel polysilicon 1752 -2050 1752 -2050 0 1
rlabel polysilicon 1752 -2056 1752 -2056 0 3
rlabel polysilicon 1759 -2050 1759 -2050 0 1
rlabel polysilicon 1762 -2050 1762 -2050 0 2
rlabel polysilicon 1762 -2056 1762 -2056 0 4
rlabel polysilicon 1766 -2050 1766 -2050 0 1
rlabel polysilicon 1766 -2056 1766 -2056 0 3
rlabel polysilicon 1773 -2050 1773 -2050 0 1
rlabel polysilicon 1773 -2056 1773 -2056 0 3
rlabel polysilicon 30 -2189 30 -2189 0 1
rlabel polysilicon 30 -2195 30 -2195 0 3
rlabel polysilicon 40 -2189 40 -2189 0 2
rlabel polysilicon 40 -2195 40 -2195 0 4
rlabel polysilicon 47 -2189 47 -2189 0 2
rlabel polysilicon 44 -2195 44 -2195 0 3
rlabel polysilicon 51 -2189 51 -2189 0 1
rlabel polysilicon 54 -2189 54 -2189 0 2
rlabel polysilicon 51 -2195 51 -2195 0 3
rlabel polysilicon 58 -2189 58 -2189 0 1
rlabel polysilicon 58 -2195 58 -2195 0 3
rlabel polysilicon 65 -2189 65 -2189 0 1
rlabel polysilicon 68 -2189 68 -2189 0 2
rlabel polysilicon 68 -2195 68 -2195 0 4
rlabel polysilicon 72 -2189 72 -2189 0 1
rlabel polysilicon 72 -2195 72 -2195 0 3
rlabel polysilicon 79 -2189 79 -2189 0 1
rlabel polysilicon 79 -2195 79 -2195 0 3
rlabel polysilicon 86 -2189 86 -2189 0 1
rlabel polysilicon 86 -2195 86 -2195 0 3
rlabel polysilicon 89 -2195 89 -2195 0 4
rlabel polysilicon 93 -2189 93 -2189 0 1
rlabel polysilicon 96 -2189 96 -2189 0 2
rlabel polysilicon 96 -2195 96 -2195 0 4
rlabel polysilicon 100 -2189 100 -2189 0 1
rlabel polysilicon 100 -2195 100 -2195 0 3
rlabel polysilicon 107 -2189 107 -2189 0 1
rlabel polysilicon 107 -2195 107 -2195 0 3
rlabel polysilicon 114 -2189 114 -2189 0 1
rlabel polysilicon 114 -2195 114 -2195 0 3
rlabel polysilicon 121 -2189 121 -2189 0 1
rlabel polysilicon 121 -2195 121 -2195 0 3
rlabel polysilicon 128 -2189 128 -2189 0 1
rlabel polysilicon 131 -2189 131 -2189 0 2
rlabel polysilicon 128 -2195 128 -2195 0 3
rlabel polysilicon 131 -2195 131 -2195 0 4
rlabel polysilicon 135 -2189 135 -2189 0 1
rlabel polysilicon 135 -2195 135 -2195 0 3
rlabel polysilicon 142 -2189 142 -2189 0 1
rlabel polysilicon 142 -2195 142 -2195 0 3
rlabel polysilicon 152 -2189 152 -2189 0 2
rlabel polysilicon 149 -2195 149 -2195 0 3
rlabel polysilicon 152 -2195 152 -2195 0 4
rlabel polysilicon 156 -2189 156 -2189 0 1
rlabel polysilicon 156 -2195 156 -2195 0 3
rlabel polysilicon 163 -2189 163 -2189 0 1
rlabel polysilicon 163 -2195 163 -2195 0 3
rlabel polysilicon 170 -2189 170 -2189 0 1
rlabel polysilicon 173 -2189 173 -2189 0 2
rlabel polysilicon 170 -2195 170 -2195 0 3
rlabel polysilicon 173 -2195 173 -2195 0 4
rlabel polysilicon 177 -2189 177 -2189 0 1
rlabel polysilicon 177 -2195 177 -2195 0 3
rlabel polysilicon 184 -2189 184 -2189 0 1
rlabel polysilicon 184 -2195 184 -2195 0 3
rlabel polysilicon 191 -2189 191 -2189 0 1
rlabel polysilicon 191 -2195 191 -2195 0 3
rlabel polysilicon 198 -2189 198 -2189 0 1
rlabel polysilicon 198 -2195 198 -2195 0 3
rlabel polysilicon 205 -2189 205 -2189 0 1
rlabel polysilicon 205 -2195 205 -2195 0 3
rlabel polysilicon 212 -2189 212 -2189 0 1
rlabel polysilicon 212 -2195 212 -2195 0 3
rlabel polysilicon 219 -2189 219 -2189 0 1
rlabel polysilicon 219 -2195 219 -2195 0 3
rlabel polysilicon 226 -2189 226 -2189 0 1
rlabel polysilicon 229 -2189 229 -2189 0 2
rlabel polysilicon 229 -2195 229 -2195 0 4
rlabel polysilicon 233 -2189 233 -2189 0 1
rlabel polysilicon 233 -2195 233 -2195 0 3
rlabel polysilicon 240 -2189 240 -2189 0 1
rlabel polysilicon 240 -2195 240 -2195 0 3
rlabel polysilicon 247 -2189 247 -2189 0 1
rlabel polysilicon 247 -2195 247 -2195 0 3
rlabel polysilicon 254 -2189 254 -2189 0 1
rlabel polysilicon 254 -2195 254 -2195 0 3
rlabel polysilicon 261 -2189 261 -2189 0 1
rlabel polysilicon 261 -2195 261 -2195 0 3
rlabel polysilicon 271 -2195 271 -2195 0 4
rlabel polysilicon 275 -2189 275 -2189 0 1
rlabel polysilicon 275 -2195 275 -2195 0 3
rlabel polysilicon 282 -2189 282 -2189 0 1
rlabel polysilicon 282 -2195 282 -2195 0 3
rlabel polysilicon 289 -2189 289 -2189 0 1
rlabel polysilicon 289 -2195 289 -2195 0 3
rlabel polysilicon 296 -2189 296 -2189 0 1
rlabel polysilicon 296 -2195 296 -2195 0 3
rlabel polysilicon 303 -2189 303 -2189 0 1
rlabel polysilicon 303 -2195 303 -2195 0 3
rlabel polysilicon 310 -2189 310 -2189 0 1
rlabel polysilicon 310 -2195 310 -2195 0 3
rlabel polysilicon 317 -2189 317 -2189 0 1
rlabel polysilicon 317 -2195 317 -2195 0 3
rlabel polysilicon 324 -2189 324 -2189 0 1
rlabel polysilicon 324 -2195 324 -2195 0 3
rlabel polysilicon 331 -2189 331 -2189 0 1
rlabel polysilicon 331 -2195 331 -2195 0 3
rlabel polysilicon 338 -2189 338 -2189 0 1
rlabel polysilicon 338 -2195 338 -2195 0 3
rlabel polysilicon 345 -2189 345 -2189 0 1
rlabel polysilicon 345 -2195 345 -2195 0 3
rlabel polysilicon 352 -2189 352 -2189 0 1
rlabel polysilicon 352 -2195 352 -2195 0 3
rlabel polysilicon 359 -2189 359 -2189 0 1
rlabel polysilicon 362 -2189 362 -2189 0 2
rlabel polysilicon 359 -2195 359 -2195 0 3
rlabel polysilicon 362 -2195 362 -2195 0 4
rlabel polysilicon 366 -2189 366 -2189 0 1
rlabel polysilicon 366 -2195 366 -2195 0 3
rlabel polysilicon 373 -2189 373 -2189 0 1
rlabel polysilicon 373 -2195 373 -2195 0 3
rlabel polysilicon 380 -2189 380 -2189 0 1
rlabel polysilicon 380 -2195 380 -2195 0 3
rlabel polysilicon 387 -2189 387 -2189 0 1
rlabel polysilicon 387 -2195 387 -2195 0 3
rlabel polysilicon 394 -2189 394 -2189 0 1
rlabel polysilicon 394 -2195 394 -2195 0 3
rlabel polysilicon 401 -2189 401 -2189 0 1
rlabel polysilicon 401 -2195 401 -2195 0 3
rlabel polysilicon 408 -2189 408 -2189 0 1
rlabel polysilicon 415 -2189 415 -2189 0 1
rlabel polysilicon 415 -2195 415 -2195 0 3
rlabel polysilicon 422 -2189 422 -2189 0 1
rlabel polysilicon 422 -2195 422 -2195 0 3
rlabel polysilicon 429 -2189 429 -2189 0 1
rlabel polysilicon 429 -2195 429 -2195 0 3
rlabel polysilicon 436 -2189 436 -2189 0 1
rlabel polysilicon 436 -2195 436 -2195 0 3
rlabel polysilicon 443 -2189 443 -2189 0 1
rlabel polysilicon 443 -2195 443 -2195 0 3
rlabel polysilicon 450 -2189 450 -2189 0 1
rlabel polysilicon 453 -2189 453 -2189 0 2
rlabel polysilicon 450 -2195 450 -2195 0 3
rlabel polysilicon 453 -2195 453 -2195 0 4
rlabel polysilicon 457 -2189 457 -2189 0 1
rlabel polysilicon 457 -2195 457 -2195 0 3
rlabel polysilicon 464 -2189 464 -2189 0 1
rlabel polysilicon 464 -2195 464 -2195 0 3
rlabel polysilicon 471 -2189 471 -2189 0 1
rlabel polysilicon 471 -2195 471 -2195 0 3
rlabel polysilicon 478 -2189 478 -2189 0 1
rlabel polysilicon 478 -2195 478 -2195 0 3
rlabel polysilicon 485 -2189 485 -2189 0 1
rlabel polysilicon 485 -2195 485 -2195 0 3
rlabel polysilicon 492 -2189 492 -2189 0 1
rlabel polysilicon 492 -2195 492 -2195 0 3
rlabel polysilicon 499 -2189 499 -2189 0 1
rlabel polysilicon 499 -2195 499 -2195 0 3
rlabel polysilicon 506 -2189 506 -2189 0 1
rlabel polysilicon 506 -2195 506 -2195 0 3
rlabel polysilicon 513 -2189 513 -2189 0 1
rlabel polysilicon 513 -2195 513 -2195 0 3
rlabel polysilicon 520 -2189 520 -2189 0 1
rlabel polysilicon 520 -2195 520 -2195 0 3
rlabel polysilicon 523 -2195 523 -2195 0 4
rlabel polysilicon 527 -2189 527 -2189 0 1
rlabel polysilicon 527 -2195 527 -2195 0 3
rlabel polysilicon 534 -2189 534 -2189 0 1
rlabel polysilicon 534 -2195 534 -2195 0 3
rlabel polysilicon 541 -2189 541 -2189 0 1
rlabel polysilicon 541 -2195 541 -2195 0 3
rlabel polysilicon 548 -2189 548 -2189 0 1
rlabel polysilicon 548 -2195 548 -2195 0 3
rlabel polysilicon 555 -2189 555 -2189 0 1
rlabel polysilicon 555 -2195 555 -2195 0 3
rlabel polysilicon 562 -2189 562 -2189 0 1
rlabel polysilicon 562 -2195 562 -2195 0 3
rlabel polysilicon 569 -2189 569 -2189 0 1
rlabel polysilicon 569 -2195 569 -2195 0 3
rlabel polysilicon 576 -2189 576 -2189 0 1
rlabel polysilicon 576 -2195 576 -2195 0 3
rlabel polysilicon 583 -2189 583 -2189 0 1
rlabel polysilicon 583 -2195 583 -2195 0 3
rlabel polysilicon 590 -2189 590 -2189 0 1
rlabel polysilicon 590 -2195 590 -2195 0 3
rlabel polysilicon 597 -2189 597 -2189 0 1
rlabel polysilicon 597 -2195 597 -2195 0 3
rlabel polysilicon 604 -2195 604 -2195 0 3
rlabel polysilicon 607 -2195 607 -2195 0 4
rlabel polysilicon 611 -2189 611 -2189 0 1
rlabel polysilicon 611 -2195 611 -2195 0 3
rlabel polysilicon 618 -2189 618 -2189 0 1
rlabel polysilicon 621 -2189 621 -2189 0 2
rlabel polysilicon 618 -2195 618 -2195 0 3
rlabel polysilicon 625 -2189 625 -2189 0 1
rlabel polysilicon 625 -2195 625 -2195 0 3
rlabel polysilicon 632 -2189 632 -2189 0 1
rlabel polysilicon 632 -2195 632 -2195 0 3
rlabel polysilicon 639 -2189 639 -2189 0 1
rlabel polysilicon 639 -2195 639 -2195 0 3
rlabel polysilicon 646 -2189 646 -2189 0 1
rlabel polysilicon 646 -2195 646 -2195 0 3
rlabel polysilicon 653 -2189 653 -2189 0 1
rlabel polysilicon 653 -2195 653 -2195 0 3
rlabel polysilicon 660 -2189 660 -2189 0 1
rlabel polysilicon 660 -2195 660 -2195 0 3
rlabel polysilicon 667 -2189 667 -2189 0 1
rlabel polysilicon 667 -2195 667 -2195 0 3
rlabel polysilicon 674 -2189 674 -2189 0 1
rlabel polysilicon 674 -2195 674 -2195 0 3
rlabel polysilicon 681 -2189 681 -2189 0 1
rlabel polysilicon 681 -2195 681 -2195 0 3
rlabel polysilicon 688 -2189 688 -2189 0 1
rlabel polysilicon 688 -2195 688 -2195 0 3
rlabel polysilicon 695 -2189 695 -2189 0 1
rlabel polysilicon 695 -2195 695 -2195 0 3
rlabel polysilicon 702 -2189 702 -2189 0 1
rlabel polysilicon 705 -2189 705 -2189 0 2
rlabel polysilicon 702 -2195 702 -2195 0 3
rlabel polysilicon 705 -2195 705 -2195 0 4
rlabel polysilicon 709 -2189 709 -2189 0 1
rlabel polysilicon 709 -2195 709 -2195 0 3
rlabel polysilicon 716 -2189 716 -2189 0 1
rlabel polysilicon 716 -2195 716 -2195 0 3
rlabel polysilicon 723 -2189 723 -2189 0 1
rlabel polysilicon 726 -2189 726 -2189 0 2
rlabel polysilicon 723 -2195 723 -2195 0 3
rlabel polysilicon 730 -2189 730 -2189 0 1
rlabel polysilicon 733 -2189 733 -2189 0 2
rlabel polysilicon 730 -2195 730 -2195 0 3
rlabel polysilicon 733 -2195 733 -2195 0 4
rlabel polysilicon 737 -2189 737 -2189 0 1
rlabel polysilicon 737 -2195 737 -2195 0 3
rlabel polysilicon 744 -2189 744 -2189 0 1
rlabel polysilicon 747 -2189 747 -2189 0 2
rlabel polysilicon 744 -2195 744 -2195 0 3
rlabel polysilicon 747 -2195 747 -2195 0 4
rlabel polysilicon 751 -2189 751 -2189 0 1
rlabel polysilicon 751 -2195 751 -2195 0 3
rlabel polysilicon 758 -2189 758 -2189 0 1
rlabel polysilicon 761 -2189 761 -2189 0 2
rlabel polysilicon 761 -2195 761 -2195 0 4
rlabel polysilicon 765 -2189 765 -2189 0 1
rlabel polysilicon 765 -2195 765 -2195 0 3
rlabel polysilicon 772 -2189 772 -2189 0 1
rlabel polysilicon 772 -2195 772 -2195 0 3
rlabel polysilicon 775 -2195 775 -2195 0 4
rlabel polysilicon 779 -2189 779 -2189 0 1
rlabel polysilicon 779 -2195 779 -2195 0 3
rlabel polysilicon 786 -2189 786 -2189 0 1
rlabel polysilicon 786 -2195 786 -2195 0 3
rlabel polysilicon 793 -2195 793 -2195 0 3
rlabel polysilicon 796 -2195 796 -2195 0 4
rlabel polysilicon 800 -2189 800 -2189 0 1
rlabel polysilicon 800 -2195 800 -2195 0 3
rlabel polysilicon 807 -2189 807 -2189 0 1
rlabel polysilicon 807 -2195 807 -2195 0 3
rlabel polysilicon 814 -2189 814 -2189 0 1
rlabel polysilicon 817 -2189 817 -2189 0 2
rlabel polysilicon 814 -2195 814 -2195 0 3
rlabel polysilicon 821 -2189 821 -2189 0 1
rlabel polysilicon 821 -2195 821 -2195 0 3
rlabel polysilicon 831 -2189 831 -2189 0 2
rlabel polysilicon 828 -2195 828 -2195 0 3
rlabel polysilicon 831 -2195 831 -2195 0 4
rlabel polysilicon 835 -2189 835 -2189 0 1
rlabel polysilicon 835 -2195 835 -2195 0 3
rlabel polysilicon 842 -2189 842 -2189 0 1
rlabel polysilicon 842 -2195 842 -2195 0 3
rlabel polysilicon 849 -2189 849 -2189 0 1
rlabel polysilicon 849 -2195 849 -2195 0 3
rlabel polysilicon 856 -2189 856 -2189 0 1
rlabel polysilicon 856 -2195 856 -2195 0 3
rlabel polysilicon 863 -2189 863 -2189 0 1
rlabel polysilicon 863 -2195 863 -2195 0 3
rlabel polysilicon 873 -2189 873 -2189 0 2
rlabel polysilicon 870 -2195 870 -2195 0 3
rlabel polysilicon 873 -2195 873 -2195 0 4
rlabel polysilicon 877 -2189 877 -2189 0 1
rlabel polysilicon 877 -2195 877 -2195 0 3
rlabel polysilicon 884 -2189 884 -2189 0 1
rlabel polysilicon 884 -2195 884 -2195 0 3
rlabel polysilicon 891 -2189 891 -2189 0 1
rlabel polysilicon 891 -2195 891 -2195 0 3
rlabel polysilicon 898 -2189 898 -2189 0 1
rlabel polysilicon 898 -2195 898 -2195 0 3
rlabel polysilicon 905 -2189 905 -2189 0 1
rlabel polysilicon 905 -2195 905 -2195 0 3
rlabel polysilicon 912 -2189 912 -2189 0 1
rlabel polysilicon 912 -2195 912 -2195 0 3
rlabel polysilicon 919 -2189 919 -2189 0 1
rlabel polysilicon 919 -2195 919 -2195 0 3
rlabel polysilicon 926 -2189 926 -2189 0 1
rlabel polysilicon 926 -2195 926 -2195 0 3
rlabel polysilicon 933 -2189 933 -2189 0 1
rlabel polysilicon 936 -2189 936 -2189 0 2
rlabel polysilicon 933 -2195 933 -2195 0 3
rlabel polysilicon 936 -2195 936 -2195 0 4
rlabel polysilicon 940 -2195 940 -2195 0 3
rlabel polysilicon 947 -2189 947 -2189 0 1
rlabel polysilicon 947 -2195 947 -2195 0 3
rlabel polysilicon 954 -2189 954 -2189 0 1
rlabel polysilicon 954 -2195 954 -2195 0 3
rlabel polysilicon 961 -2189 961 -2189 0 1
rlabel polysilicon 961 -2195 961 -2195 0 3
rlabel polysilicon 968 -2189 968 -2189 0 1
rlabel polysilicon 968 -2195 968 -2195 0 3
rlabel polysilicon 978 -2189 978 -2189 0 2
rlabel polysilicon 975 -2195 975 -2195 0 3
rlabel polysilicon 978 -2195 978 -2195 0 4
rlabel polysilicon 982 -2189 982 -2189 0 1
rlabel polysilicon 982 -2195 982 -2195 0 3
rlabel polysilicon 989 -2189 989 -2189 0 1
rlabel polysilicon 989 -2195 989 -2195 0 3
rlabel polysilicon 996 -2189 996 -2189 0 1
rlabel polysilicon 996 -2195 996 -2195 0 3
rlabel polysilicon 999 -2195 999 -2195 0 4
rlabel polysilicon 1003 -2189 1003 -2189 0 1
rlabel polysilicon 1003 -2195 1003 -2195 0 3
rlabel polysilicon 1013 -2189 1013 -2189 0 2
rlabel polysilicon 1010 -2195 1010 -2195 0 3
rlabel polysilicon 1013 -2195 1013 -2195 0 4
rlabel polysilicon 1017 -2189 1017 -2189 0 1
rlabel polysilicon 1017 -2195 1017 -2195 0 3
rlabel polysilicon 1024 -2189 1024 -2189 0 1
rlabel polysilicon 1024 -2195 1024 -2195 0 3
rlabel polysilicon 1031 -2189 1031 -2189 0 1
rlabel polysilicon 1031 -2195 1031 -2195 0 3
rlabel polysilicon 1038 -2189 1038 -2189 0 1
rlabel polysilicon 1038 -2195 1038 -2195 0 3
rlabel polysilicon 1045 -2189 1045 -2189 0 1
rlabel polysilicon 1045 -2195 1045 -2195 0 3
rlabel polysilicon 1052 -2189 1052 -2189 0 1
rlabel polysilicon 1052 -2195 1052 -2195 0 3
rlabel polysilicon 1059 -2189 1059 -2189 0 1
rlabel polysilicon 1059 -2195 1059 -2195 0 3
rlabel polysilicon 1066 -2189 1066 -2189 0 1
rlabel polysilicon 1066 -2195 1066 -2195 0 3
rlabel polysilicon 1073 -2189 1073 -2189 0 1
rlabel polysilicon 1073 -2195 1073 -2195 0 3
rlabel polysilicon 1080 -2189 1080 -2189 0 1
rlabel polysilicon 1080 -2195 1080 -2195 0 3
rlabel polysilicon 1087 -2189 1087 -2189 0 1
rlabel polysilicon 1087 -2195 1087 -2195 0 3
rlabel polysilicon 1094 -2189 1094 -2189 0 1
rlabel polysilicon 1094 -2195 1094 -2195 0 3
rlabel polysilicon 1104 -2189 1104 -2189 0 2
rlabel polysilicon 1101 -2195 1101 -2195 0 3
rlabel polysilicon 1104 -2195 1104 -2195 0 4
rlabel polysilicon 1108 -2189 1108 -2189 0 1
rlabel polysilicon 1108 -2195 1108 -2195 0 3
rlabel polysilicon 1115 -2189 1115 -2189 0 1
rlabel polysilicon 1118 -2189 1118 -2189 0 2
rlabel polysilicon 1115 -2195 1115 -2195 0 3
rlabel polysilicon 1118 -2195 1118 -2195 0 4
rlabel polysilicon 1122 -2189 1122 -2189 0 1
rlabel polysilicon 1122 -2195 1122 -2195 0 3
rlabel polysilicon 1129 -2189 1129 -2189 0 1
rlabel polysilicon 1129 -2195 1129 -2195 0 3
rlabel polysilicon 1136 -2189 1136 -2189 0 1
rlabel polysilicon 1136 -2195 1136 -2195 0 3
rlabel polysilicon 1143 -2189 1143 -2189 0 1
rlabel polysilicon 1143 -2195 1143 -2195 0 3
rlabel polysilicon 1150 -2189 1150 -2189 0 1
rlabel polysilicon 1150 -2195 1150 -2195 0 3
rlabel polysilicon 1157 -2189 1157 -2189 0 1
rlabel polysilicon 1157 -2195 1157 -2195 0 3
rlabel polysilicon 1164 -2189 1164 -2189 0 1
rlabel polysilicon 1164 -2195 1164 -2195 0 3
rlabel polysilicon 1171 -2189 1171 -2189 0 1
rlabel polysilicon 1171 -2195 1171 -2195 0 3
rlabel polysilicon 1178 -2189 1178 -2189 0 1
rlabel polysilicon 1178 -2195 1178 -2195 0 3
rlabel polysilicon 1185 -2189 1185 -2189 0 1
rlabel polysilicon 1185 -2195 1185 -2195 0 3
rlabel polysilicon 1192 -2189 1192 -2189 0 1
rlabel polysilicon 1192 -2195 1192 -2195 0 3
rlabel polysilicon 1199 -2189 1199 -2189 0 1
rlabel polysilicon 1199 -2195 1199 -2195 0 3
rlabel polysilicon 1206 -2189 1206 -2189 0 1
rlabel polysilicon 1206 -2195 1206 -2195 0 3
rlabel polysilicon 1213 -2189 1213 -2189 0 1
rlabel polysilicon 1213 -2195 1213 -2195 0 3
rlabel polysilicon 1220 -2189 1220 -2189 0 1
rlabel polysilicon 1220 -2195 1220 -2195 0 3
rlabel polysilicon 1227 -2189 1227 -2189 0 1
rlabel polysilicon 1227 -2195 1227 -2195 0 3
rlabel polysilicon 1234 -2189 1234 -2189 0 1
rlabel polysilicon 1234 -2195 1234 -2195 0 3
rlabel polysilicon 1241 -2189 1241 -2189 0 1
rlabel polysilicon 1241 -2195 1241 -2195 0 3
rlabel polysilicon 1248 -2189 1248 -2189 0 1
rlabel polysilicon 1248 -2195 1248 -2195 0 3
rlabel polysilicon 1255 -2189 1255 -2189 0 1
rlabel polysilicon 1255 -2195 1255 -2195 0 3
rlabel polysilicon 1262 -2189 1262 -2189 0 1
rlabel polysilicon 1262 -2195 1262 -2195 0 3
rlabel polysilicon 1269 -2189 1269 -2189 0 1
rlabel polysilicon 1269 -2195 1269 -2195 0 3
rlabel polysilicon 1276 -2189 1276 -2189 0 1
rlabel polysilicon 1276 -2195 1276 -2195 0 3
rlabel polysilicon 1283 -2189 1283 -2189 0 1
rlabel polysilicon 1283 -2195 1283 -2195 0 3
rlabel polysilicon 1290 -2189 1290 -2189 0 1
rlabel polysilicon 1290 -2195 1290 -2195 0 3
rlabel polysilicon 1297 -2189 1297 -2189 0 1
rlabel polysilicon 1297 -2195 1297 -2195 0 3
rlabel polysilicon 1304 -2189 1304 -2189 0 1
rlabel polysilicon 1304 -2195 1304 -2195 0 3
rlabel polysilicon 1311 -2189 1311 -2189 0 1
rlabel polysilicon 1311 -2195 1311 -2195 0 3
rlabel polysilicon 1318 -2189 1318 -2189 0 1
rlabel polysilicon 1318 -2195 1318 -2195 0 3
rlabel polysilicon 1325 -2189 1325 -2189 0 1
rlabel polysilicon 1325 -2195 1325 -2195 0 3
rlabel polysilicon 1332 -2189 1332 -2189 0 1
rlabel polysilicon 1332 -2195 1332 -2195 0 3
rlabel polysilicon 1339 -2189 1339 -2189 0 1
rlabel polysilicon 1339 -2195 1339 -2195 0 3
rlabel polysilicon 1346 -2189 1346 -2189 0 1
rlabel polysilicon 1346 -2195 1346 -2195 0 3
rlabel polysilicon 1353 -2189 1353 -2189 0 1
rlabel polysilicon 1353 -2195 1353 -2195 0 3
rlabel polysilicon 1360 -2189 1360 -2189 0 1
rlabel polysilicon 1360 -2195 1360 -2195 0 3
rlabel polysilicon 1367 -2189 1367 -2189 0 1
rlabel polysilicon 1367 -2195 1367 -2195 0 3
rlabel polysilicon 1374 -2189 1374 -2189 0 1
rlabel polysilicon 1374 -2195 1374 -2195 0 3
rlabel polysilicon 1381 -2189 1381 -2189 0 1
rlabel polysilicon 1381 -2195 1381 -2195 0 3
rlabel polysilicon 1388 -2189 1388 -2189 0 1
rlabel polysilicon 1388 -2195 1388 -2195 0 3
rlabel polysilicon 1395 -2189 1395 -2189 0 1
rlabel polysilicon 1395 -2195 1395 -2195 0 3
rlabel polysilicon 1402 -2189 1402 -2189 0 1
rlabel polysilicon 1402 -2195 1402 -2195 0 3
rlabel polysilicon 1409 -2189 1409 -2189 0 1
rlabel polysilicon 1409 -2195 1409 -2195 0 3
rlabel polysilicon 1416 -2189 1416 -2189 0 1
rlabel polysilicon 1416 -2195 1416 -2195 0 3
rlabel polysilicon 1423 -2189 1423 -2189 0 1
rlabel polysilicon 1423 -2195 1423 -2195 0 3
rlabel polysilicon 1430 -2189 1430 -2189 0 1
rlabel polysilicon 1430 -2195 1430 -2195 0 3
rlabel polysilicon 1437 -2189 1437 -2189 0 1
rlabel polysilicon 1437 -2195 1437 -2195 0 3
rlabel polysilicon 1444 -2189 1444 -2189 0 1
rlabel polysilicon 1444 -2195 1444 -2195 0 3
rlabel polysilicon 1451 -2189 1451 -2189 0 1
rlabel polysilicon 1451 -2195 1451 -2195 0 3
rlabel polysilicon 1458 -2189 1458 -2189 0 1
rlabel polysilicon 1458 -2195 1458 -2195 0 3
rlabel polysilicon 1465 -2189 1465 -2189 0 1
rlabel polysilicon 1465 -2195 1465 -2195 0 3
rlabel polysilicon 1472 -2189 1472 -2189 0 1
rlabel polysilicon 1472 -2195 1472 -2195 0 3
rlabel polysilicon 1479 -2189 1479 -2189 0 1
rlabel polysilicon 1479 -2195 1479 -2195 0 3
rlabel polysilicon 1486 -2189 1486 -2189 0 1
rlabel polysilicon 1486 -2195 1486 -2195 0 3
rlabel polysilicon 1493 -2189 1493 -2189 0 1
rlabel polysilicon 1493 -2195 1493 -2195 0 3
rlabel polysilicon 1500 -2189 1500 -2189 0 1
rlabel polysilicon 1500 -2195 1500 -2195 0 3
rlabel polysilicon 1507 -2189 1507 -2189 0 1
rlabel polysilicon 1507 -2195 1507 -2195 0 3
rlabel polysilicon 1514 -2189 1514 -2189 0 1
rlabel polysilicon 1514 -2195 1514 -2195 0 3
rlabel polysilicon 1521 -2189 1521 -2189 0 1
rlabel polysilicon 1521 -2195 1521 -2195 0 3
rlabel polysilicon 1528 -2189 1528 -2189 0 1
rlabel polysilicon 1528 -2195 1528 -2195 0 3
rlabel polysilicon 1535 -2189 1535 -2189 0 1
rlabel polysilicon 1535 -2195 1535 -2195 0 3
rlabel polysilicon 1542 -2189 1542 -2189 0 1
rlabel polysilicon 1542 -2195 1542 -2195 0 3
rlabel polysilicon 1549 -2189 1549 -2189 0 1
rlabel polysilicon 1549 -2195 1549 -2195 0 3
rlabel polysilicon 1556 -2189 1556 -2189 0 1
rlabel polysilicon 1556 -2195 1556 -2195 0 3
rlabel polysilicon 1563 -2189 1563 -2189 0 1
rlabel polysilicon 1563 -2195 1563 -2195 0 3
rlabel polysilicon 1570 -2189 1570 -2189 0 1
rlabel polysilicon 1570 -2195 1570 -2195 0 3
rlabel polysilicon 1577 -2189 1577 -2189 0 1
rlabel polysilicon 1577 -2195 1577 -2195 0 3
rlabel polysilicon 1584 -2189 1584 -2189 0 1
rlabel polysilicon 1584 -2195 1584 -2195 0 3
rlabel polysilicon 1591 -2189 1591 -2189 0 1
rlabel polysilicon 1591 -2195 1591 -2195 0 3
rlabel polysilicon 1598 -2189 1598 -2189 0 1
rlabel polysilicon 1598 -2195 1598 -2195 0 3
rlabel polysilicon 1605 -2189 1605 -2189 0 1
rlabel polysilicon 1605 -2195 1605 -2195 0 3
rlabel polysilicon 1612 -2189 1612 -2189 0 1
rlabel polysilicon 1612 -2195 1612 -2195 0 3
rlabel polysilicon 1619 -2189 1619 -2189 0 1
rlabel polysilicon 1619 -2195 1619 -2195 0 3
rlabel polysilicon 1626 -2189 1626 -2189 0 1
rlabel polysilicon 1629 -2189 1629 -2189 0 2
rlabel polysilicon 1626 -2195 1626 -2195 0 3
rlabel polysilicon 1633 -2189 1633 -2189 0 1
rlabel polysilicon 1633 -2195 1633 -2195 0 3
rlabel polysilicon 1640 -2189 1640 -2189 0 1
rlabel polysilicon 1640 -2195 1640 -2195 0 3
rlabel polysilicon 1647 -2189 1647 -2189 0 1
rlabel polysilicon 1647 -2195 1647 -2195 0 3
rlabel polysilicon 1654 -2189 1654 -2189 0 1
rlabel polysilicon 1654 -2195 1654 -2195 0 3
rlabel polysilicon 1661 -2189 1661 -2189 0 1
rlabel polysilicon 1661 -2195 1661 -2195 0 3
rlabel polysilicon 1668 -2189 1668 -2189 0 1
rlabel polysilicon 1668 -2195 1668 -2195 0 3
rlabel polysilicon 1675 -2189 1675 -2189 0 1
rlabel polysilicon 1675 -2195 1675 -2195 0 3
rlabel polysilicon 1682 -2189 1682 -2189 0 1
rlabel polysilicon 1682 -2195 1682 -2195 0 3
rlabel polysilicon 1689 -2189 1689 -2189 0 1
rlabel polysilicon 1689 -2195 1689 -2195 0 3
rlabel polysilicon 1696 -2189 1696 -2189 0 1
rlabel polysilicon 1696 -2195 1696 -2195 0 3
rlabel polysilicon 1703 -2189 1703 -2189 0 1
rlabel polysilicon 1703 -2195 1703 -2195 0 3
rlabel polysilicon 1710 -2189 1710 -2189 0 1
rlabel polysilicon 1710 -2195 1710 -2195 0 3
rlabel polysilicon 1717 -2189 1717 -2189 0 1
rlabel polysilicon 1717 -2195 1717 -2195 0 3
rlabel polysilicon 1724 -2189 1724 -2189 0 1
rlabel polysilicon 1724 -2195 1724 -2195 0 3
rlabel polysilicon 1731 -2189 1731 -2189 0 1
rlabel polysilicon 1731 -2195 1731 -2195 0 3
rlabel polysilicon 1738 -2189 1738 -2189 0 1
rlabel polysilicon 1738 -2195 1738 -2195 0 3
rlabel polysilicon 1745 -2189 1745 -2189 0 1
rlabel polysilicon 1745 -2195 1745 -2195 0 3
rlabel polysilicon 1755 -2189 1755 -2189 0 2
rlabel polysilicon 1752 -2195 1752 -2195 0 3
rlabel polysilicon 1755 -2195 1755 -2195 0 4
rlabel polysilicon 1759 -2189 1759 -2189 0 1
rlabel polysilicon 1759 -2195 1759 -2195 0 3
rlabel polysilicon 1766 -2189 1766 -2189 0 1
rlabel polysilicon 1766 -2195 1766 -2195 0 3
rlabel polysilicon 44 -2324 44 -2324 0 1
rlabel polysilicon 44 -2330 44 -2330 0 3
rlabel polysilicon 51 -2324 51 -2324 0 1
rlabel polysilicon 51 -2330 51 -2330 0 3
rlabel polysilicon 58 -2324 58 -2324 0 1
rlabel polysilicon 58 -2330 58 -2330 0 3
rlabel polysilicon 65 -2324 65 -2324 0 1
rlabel polysilicon 65 -2330 65 -2330 0 3
rlabel polysilicon 72 -2324 72 -2324 0 1
rlabel polysilicon 72 -2330 72 -2330 0 3
rlabel polysilicon 79 -2324 79 -2324 0 1
rlabel polysilicon 79 -2330 79 -2330 0 3
rlabel polysilicon 89 -2324 89 -2324 0 2
rlabel polysilicon 86 -2330 86 -2330 0 3
rlabel polysilicon 93 -2324 93 -2324 0 1
rlabel polysilicon 96 -2324 96 -2324 0 2
rlabel polysilicon 93 -2330 93 -2330 0 3
rlabel polysilicon 96 -2330 96 -2330 0 4
rlabel polysilicon 100 -2324 100 -2324 0 1
rlabel polysilicon 100 -2330 100 -2330 0 3
rlabel polysilicon 107 -2324 107 -2324 0 1
rlabel polysilicon 107 -2330 107 -2330 0 3
rlabel polysilicon 114 -2324 114 -2324 0 1
rlabel polysilicon 117 -2324 117 -2324 0 2
rlabel polysilicon 114 -2330 114 -2330 0 3
rlabel polysilicon 117 -2330 117 -2330 0 4
rlabel polysilicon 121 -2324 121 -2324 0 1
rlabel polysilicon 121 -2330 121 -2330 0 3
rlabel polysilicon 128 -2324 128 -2324 0 1
rlabel polysilicon 128 -2330 128 -2330 0 3
rlabel polysilicon 135 -2324 135 -2324 0 1
rlabel polysilicon 138 -2324 138 -2324 0 2
rlabel polysilicon 135 -2330 135 -2330 0 3
rlabel polysilicon 138 -2330 138 -2330 0 4
rlabel polysilicon 142 -2324 142 -2324 0 1
rlabel polysilicon 142 -2330 142 -2330 0 3
rlabel polysilicon 149 -2324 149 -2324 0 1
rlabel polysilicon 149 -2330 149 -2330 0 3
rlabel polysilicon 156 -2324 156 -2324 0 1
rlabel polysilicon 156 -2330 156 -2330 0 3
rlabel polysilicon 163 -2324 163 -2324 0 1
rlabel polysilicon 163 -2330 163 -2330 0 3
rlabel polysilicon 170 -2324 170 -2324 0 1
rlabel polysilicon 173 -2324 173 -2324 0 2
rlabel polysilicon 170 -2330 170 -2330 0 3
rlabel polysilicon 173 -2330 173 -2330 0 4
rlabel polysilicon 177 -2324 177 -2324 0 1
rlabel polysilicon 177 -2330 177 -2330 0 3
rlabel polysilicon 184 -2324 184 -2324 0 1
rlabel polysilicon 184 -2330 184 -2330 0 3
rlabel polysilicon 191 -2324 191 -2324 0 1
rlabel polysilicon 191 -2330 191 -2330 0 3
rlabel polysilicon 198 -2324 198 -2324 0 1
rlabel polysilicon 198 -2330 198 -2330 0 3
rlabel polysilicon 205 -2324 205 -2324 0 1
rlabel polysilicon 205 -2330 205 -2330 0 3
rlabel polysilicon 215 -2324 215 -2324 0 2
rlabel polysilicon 212 -2330 212 -2330 0 3
rlabel polysilicon 215 -2330 215 -2330 0 4
rlabel polysilicon 219 -2324 219 -2324 0 1
rlabel polysilicon 219 -2330 219 -2330 0 3
rlabel polysilicon 226 -2324 226 -2324 0 1
rlabel polysilicon 226 -2330 226 -2330 0 3
rlabel polysilicon 233 -2324 233 -2324 0 1
rlabel polysilicon 236 -2324 236 -2324 0 2
rlabel polysilicon 236 -2330 236 -2330 0 4
rlabel polysilicon 240 -2324 240 -2324 0 1
rlabel polysilicon 240 -2330 240 -2330 0 3
rlabel polysilicon 247 -2324 247 -2324 0 1
rlabel polysilicon 247 -2330 247 -2330 0 3
rlabel polysilicon 254 -2324 254 -2324 0 1
rlabel polysilicon 254 -2330 254 -2330 0 3
rlabel polysilicon 261 -2324 261 -2324 0 1
rlabel polysilicon 261 -2330 261 -2330 0 3
rlabel polysilicon 268 -2324 268 -2324 0 1
rlabel polysilicon 268 -2330 268 -2330 0 3
rlabel polysilicon 275 -2324 275 -2324 0 1
rlabel polysilicon 275 -2330 275 -2330 0 3
rlabel polysilicon 282 -2324 282 -2324 0 1
rlabel polysilicon 282 -2330 282 -2330 0 3
rlabel polysilicon 289 -2324 289 -2324 0 1
rlabel polysilicon 289 -2330 289 -2330 0 3
rlabel polysilicon 296 -2324 296 -2324 0 1
rlabel polysilicon 296 -2330 296 -2330 0 3
rlabel polysilicon 303 -2324 303 -2324 0 1
rlabel polysilicon 303 -2330 303 -2330 0 3
rlabel polysilicon 310 -2324 310 -2324 0 1
rlabel polysilicon 310 -2330 310 -2330 0 3
rlabel polysilicon 317 -2324 317 -2324 0 1
rlabel polysilicon 317 -2330 317 -2330 0 3
rlabel polysilicon 324 -2324 324 -2324 0 1
rlabel polysilicon 324 -2330 324 -2330 0 3
rlabel polysilicon 331 -2324 331 -2324 0 1
rlabel polysilicon 331 -2330 331 -2330 0 3
rlabel polysilicon 338 -2324 338 -2324 0 1
rlabel polysilicon 338 -2330 338 -2330 0 3
rlabel polysilicon 345 -2324 345 -2324 0 1
rlabel polysilicon 345 -2330 345 -2330 0 3
rlabel polysilicon 352 -2324 352 -2324 0 1
rlabel polysilicon 352 -2330 352 -2330 0 3
rlabel polysilicon 359 -2324 359 -2324 0 1
rlabel polysilicon 359 -2330 359 -2330 0 3
rlabel polysilicon 366 -2324 366 -2324 0 1
rlabel polysilicon 366 -2330 366 -2330 0 3
rlabel polysilicon 373 -2324 373 -2324 0 1
rlabel polysilicon 373 -2330 373 -2330 0 3
rlabel polysilicon 380 -2324 380 -2324 0 1
rlabel polysilicon 380 -2330 380 -2330 0 3
rlabel polysilicon 387 -2324 387 -2324 0 1
rlabel polysilicon 387 -2330 387 -2330 0 3
rlabel polysilicon 394 -2324 394 -2324 0 1
rlabel polysilicon 394 -2330 394 -2330 0 3
rlabel polysilicon 401 -2324 401 -2324 0 1
rlabel polysilicon 401 -2330 401 -2330 0 3
rlabel polysilicon 408 -2324 408 -2324 0 1
rlabel polysilicon 408 -2330 408 -2330 0 3
rlabel polysilicon 415 -2324 415 -2324 0 1
rlabel polysilicon 415 -2330 415 -2330 0 3
rlabel polysilicon 422 -2324 422 -2324 0 1
rlabel polysilicon 422 -2330 422 -2330 0 3
rlabel polysilicon 429 -2324 429 -2324 0 1
rlabel polysilicon 429 -2330 429 -2330 0 3
rlabel polysilicon 436 -2324 436 -2324 0 1
rlabel polysilicon 436 -2330 436 -2330 0 3
rlabel polysilicon 443 -2324 443 -2324 0 1
rlabel polysilicon 443 -2330 443 -2330 0 3
rlabel polysilicon 450 -2324 450 -2324 0 1
rlabel polysilicon 450 -2330 450 -2330 0 3
rlabel polysilicon 457 -2324 457 -2324 0 1
rlabel polysilicon 457 -2330 457 -2330 0 3
rlabel polysilicon 464 -2324 464 -2324 0 1
rlabel polysilicon 464 -2330 464 -2330 0 3
rlabel polysilicon 471 -2324 471 -2324 0 1
rlabel polysilicon 471 -2330 471 -2330 0 3
rlabel polysilicon 478 -2324 478 -2324 0 1
rlabel polysilicon 478 -2330 478 -2330 0 3
rlabel polysilicon 485 -2324 485 -2324 0 1
rlabel polysilicon 485 -2330 485 -2330 0 3
rlabel polysilicon 492 -2324 492 -2324 0 1
rlabel polysilicon 492 -2330 492 -2330 0 3
rlabel polysilicon 499 -2324 499 -2324 0 1
rlabel polysilicon 499 -2330 499 -2330 0 3
rlabel polysilicon 506 -2324 506 -2324 0 1
rlabel polysilicon 506 -2330 506 -2330 0 3
rlabel polysilicon 513 -2324 513 -2324 0 1
rlabel polysilicon 513 -2330 513 -2330 0 3
rlabel polysilicon 520 -2324 520 -2324 0 1
rlabel polysilicon 520 -2330 520 -2330 0 3
rlabel polysilicon 527 -2324 527 -2324 0 1
rlabel polysilicon 527 -2330 527 -2330 0 3
rlabel polysilicon 534 -2324 534 -2324 0 1
rlabel polysilicon 534 -2330 534 -2330 0 3
rlabel polysilicon 537 -2330 537 -2330 0 4
rlabel polysilicon 541 -2324 541 -2324 0 1
rlabel polysilicon 541 -2330 541 -2330 0 3
rlabel polysilicon 548 -2324 548 -2324 0 1
rlabel polysilicon 548 -2330 548 -2330 0 3
rlabel polysilicon 555 -2324 555 -2324 0 1
rlabel polysilicon 555 -2330 555 -2330 0 3
rlabel polysilicon 562 -2324 562 -2324 0 1
rlabel polysilicon 562 -2330 562 -2330 0 3
rlabel polysilicon 569 -2324 569 -2324 0 1
rlabel polysilicon 569 -2330 569 -2330 0 3
rlabel polysilicon 576 -2324 576 -2324 0 1
rlabel polysilicon 576 -2330 576 -2330 0 3
rlabel polysilicon 583 -2324 583 -2324 0 1
rlabel polysilicon 586 -2324 586 -2324 0 2
rlabel polysilicon 583 -2330 583 -2330 0 3
rlabel polysilicon 590 -2324 590 -2324 0 1
rlabel polysilicon 590 -2330 590 -2330 0 3
rlabel polysilicon 597 -2324 597 -2324 0 1
rlabel polysilicon 597 -2330 597 -2330 0 3
rlabel polysilicon 604 -2324 604 -2324 0 1
rlabel polysilicon 604 -2330 604 -2330 0 3
rlabel polysilicon 611 -2324 611 -2324 0 1
rlabel polysilicon 611 -2330 611 -2330 0 3
rlabel polysilicon 618 -2324 618 -2324 0 1
rlabel polysilicon 618 -2330 618 -2330 0 3
rlabel polysilicon 625 -2324 625 -2324 0 1
rlabel polysilicon 625 -2330 625 -2330 0 3
rlabel polysilicon 632 -2324 632 -2324 0 1
rlabel polysilicon 632 -2330 632 -2330 0 3
rlabel polysilicon 639 -2324 639 -2324 0 1
rlabel polysilicon 642 -2330 642 -2330 0 4
rlabel polysilicon 646 -2324 646 -2324 0 1
rlabel polysilicon 646 -2330 646 -2330 0 3
rlabel polysilicon 653 -2324 653 -2324 0 1
rlabel polysilicon 656 -2324 656 -2324 0 2
rlabel polysilicon 653 -2330 653 -2330 0 3
rlabel polysilicon 656 -2330 656 -2330 0 4
rlabel polysilicon 660 -2324 660 -2324 0 1
rlabel polysilicon 660 -2330 660 -2330 0 3
rlabel polysilicon 667 -2324 667 -2324 0 1
rlabel polysilicon 667 -2330 667 -2330 0 3
rlabel polysilicon 674 -2324 674 -2324 0 1
rlabel polysilicon 674 -2330 674 -2330 0 3
rlabel polysilicon 681 -2324 681 -2324 0 1
rlabel polysilicon 681 -2330 681 -2330 0 3
rlabel polysilicon 688 -2324 688 -2324 0 1
rlabel polysilicon 691 -2324 691 -2324 0 2
rlabel polysilicon 688 -2330 688 -2330 0 3
rlabel polysilicon 691 -2330 691 -2330 0 4
rlabel polysilicon 695 -2324 695 -2324 0 1
rlabel polysilicon 695 -2330 695 -2330 0 3
rlabel polysilicon 702 -2324 702 -2324 0 1
rlabel polysilicon 705 -2324 705 -2324 0 2
rlabel polysilicon 702 -2330 702 -2330 0 3
rlabel polysilicon 705 -2330 705 -2330 0 4
rlabel polysilicon 709 -2324 709 -2324 0 1
rlabel polysilicon 709 -2330 709 -2330 0 3
rlabel polysilicon 716 -2324 716 -2324 0 1
rlabel polysilicon 716 -2330 716 -2330 0 3
rlabel polysilicon 723 -2324 723 -2324 0 1
rlabel polysilicon 723 -2330 723 -2330 0 3
rlabel polysilicon 730 -2324 730 -2324 0 1
rlabel polysilicon 733 -2324 733 -2324 0 2
rlabel polysilicon 730 -2330 730 -2330 0 3
rlabel polysilicon 733 -2330 733 -2330 0 4
rlabel polysilicon 737 -2324 737 -2324 0 1
rlabel polysilicon 737 -2330 737 -2330 0 3
rlabel polysilicon 744 -2324 744 -2324 0 1
rlabel polysilicon 747 -2324 747 -2324 0 2
rlabel polysilicon 744 -2330 744 -2330 0 3
rlabel polysilicon 747 -2330 747 -2330 0 4
rlabel polysilicon 751 -2324 751 -2324 0 1
rlabel polysilicon 751 -2330 751 -2330 0 3
rlabel polysilicon 758 -2324 758 -2324 0 1
rlabel polysilicon 758 -2330 758 -2330 0 3
rlabel polysilicon 765 -2324 765 -2324 0 1
rlabel polysilicon 765 -2330 765 -2330 0 3
rlabel polysilicon 772 -2324 772 -2324 0 1
rlabel polysilicon 772 -2330 772 -2330 0 3
rlabel polysilicon 775 -2330 775 -2330 0 4
rlabel polysilicon 779 -2324 779 -2324 0 1
rlabel polysilicon 779 -2330 779 -2330 0 3
rlabel polysilicon 786 -2324 786 -2324 0 1
rlabel polysilicon 786 -2330 786 -2330 0 3
rlabel polysilicon 793 -2324 793 -2324 0 1
rlabel polysilicon 793 -2330 793 -2330 0 3
rlabel polysilicon 800 -2324 800 -2324 0 1
rlabel polysilicon 800 -2330 800 -2330 0 3
rlabel polysilicon 807 -2324 807 -2324 0 1
rlabel polysilicon 807 -2330 807 -2330 0 3
rlabel polysilicon 814 -2324 814 -2324 0 1
rlabel polysilicon 814 -2330 814 -2330 0 3
rlabel polysilicon 821 -2324 821 -2324 0 1
rlabel polysilicon 821 -2330 821 -2330 0 3
rlabel polysilicon 828 -2324 828 -2324 0 1
rlabel polysilicon 828 -2330 828 -2330 0 3
rlabel polysilicon 835 -2324 835 -2324 0 1
rlabel polysilicon 835 -2330 835 -2330 0 3
rlabel polysilicon 842 -2324 842 -2324 0 1
rlabel polysilicon 842 -2330 842 -2330 0 3
rlabel polysilicon 849 -2324 849 -2324 0 1
rlabel polysilicon 852 -2324 852 -2324 0 2
rlabel polysilicon 849 -2330 849 -2330 0 3
rlabel polysilicon 856 -2324 856 -2324 0 1
rlabel polysilicon 856 -2330 856 -2330 0 3
rlabel polysilicon 863 -2324 863 -2324 0 1
rlabel polysilicon 863 -2330 863 -2330 0 3
rlabel polysilicon 870 -2324 870 -2324 0 1
rlabel polysilicon 873 -2324 873 -2324 0 2
rlabel polysilicon 873 -2330 873 -2330 0 4
rlabel polysilicon 877 -2324 877 -2324 0 1
rlabel polysilicon 877 -2330 877 -2330 0 3
rlabel polysilicon 884 -2324 884 -2324 0 1
rlabel polysilicon 884 -2330 884 -2330 0 3
rlabel polysilicon 891 -2324 891 -2324 0 1
rlabel polysilicon 891 -2330 891 -2330 0 3
rlabel polysilicon 898 -2324 898 -2324 0 1
rlabel polysilicon 901 -2324 901 -2324 0 2
rlabel polysilicon 898 -2330 898 -2330 0 3
rlabel polysilicon 901 -2330 901 -2330 0 4
rlabel polysilicon 905 -2324 905 -2324 0 1
rlabel polysilicon 905 -2330 905 -2330 0 3
rlabel polysilicon 912 -2324 912 -2324 0 1
rlabel polysilicon 912 -2330 912 -2330 0 3
rlabel polysilicon 919 -2324 919 -2324 0 1
rlabel polysilicon 919 -2330 919 -2330 0 3
rlabel polysilicon 926 -2324 926 -2324 0 1
rlabel polysilicon 926 -2330 926 -2330 0 3
rlabel polysilicon 933 -2324 933 -2324 0 1
rlabel polysilicon 933 -2330 933 -2330 0 3
rlabel polysilicon 940 -2324 940 -2324 0 1
rlabel polysilicon 940 -2330 940 -2330 0 3
rlabel polysilicon 947 -2324 947 -2324 0 1
rlabel polysilicon 947 -2330 947 -2330 0 3
rlabel polysilicon 954 -2324 954 -2324 0 1
rlabel polysilicon 957 -2324 957 -2324 0 2
rlabel polysilicon 954 -2330 954 -2330 0 3
rlabel polysilicon 957 -2330 957 -2330 0 4
rlabel polysilicon 961 -2324 961 -2324 0 1
rlabel polysilicon 961 -2330 961 -2330 0 3
rlabel polysilicon 968 -2324 968 -2324 0 1
rlabel polysilicon 971 -2330 971 -2330 0 4
rlabel polysilicon 975 -2324 975 -2324 0 1
rlabel polysilicon 975 -2330 975 -2330 0 3
rlabel polysilicon 982 -2324 982 -2324 0 1
rlabel polysilicon 982 -2330 982 -2330 0 3
rlabel polysilicon 989 -2324 989 -2324 0 1
rlabel polysilicon 989 -2330 989 -2330 0 3
rlabel polysilicon 996 -2324 996 -2324 0 1
rlabel polysilicon 999 -2324 999 -2324 0 2
rlabel polysilicon 996 -2330 996 -2330 0 3
rlabel polysilicon 999 -2330 999 -2330 0 4
rlabel polysilicon 1003 -2324 1003 -2324 0 1
rlabel polysilicon 1003 -2330 1003 -2330 0 3
rlabel polysilicon 1010 -2324 1010 -2324 0 1
rlabel polysilicon 1010 -2330 1010 -2330 0 3
rlabel polysilicon 1017 -2324 1017 -2324 0 1
rlabel polysilicon 1017 -2330 1017 -2330 0 3
rlabel polysilicon 1024 -2324 1024 -2324 0 1
rlabel polysilicon 1024 -2330 1024 -2330 0 3
rlabel polysilicon 1031 -2324 1031 -2324 0 1
rlabel polysilicon 1031 -2330 1031 -2330 0 3
rlabel polysilicon 1038 -2324 1038 -2324 0 1
rlabel polysilicon 1038 -2330 1038 -2330 0 3
rlabel polysilicon 1045 -2324 1045 -2324 0 1
rlabel polysilicon 1045 -2330 1045 -2330 0 3
rlabel polysilicon 1052 -2324 1052 -2324 0 1
rlabel polysilicon 1052 -2330 1052 -2330 0 3
rlabel polysilicon 1059 -2324 1059 -2324 0 1
rlabel polysilicon 1059 -2330 1059 -2330 0 3
rlabel polysilicon 1066 -2324 1066 -2324 0 1
rlabel polysilicon 1066 -2330 1066 -2330 0 3
rlabel polysilicon 1073 -2324 1073 -2324 0 1
rlabel polysilicon 1073 -2330 1073 -2330 0 3
rlabel polysilicon 1083 -2324 1083 -2324 0 2
rlabel polysilicon 1080 -2330 1080 -2330 0 3
rlabel polysilicon 1083 -2330 1083 -2330 0 4
rlabel polysilicon 1087 -2324 1087 -2324 0 1
rlabel polysilicon 1087 -2330 1087 -2330 0 3
rlabel polysilicon 1094 -2324 1094 -2324 0 1
rlabel polysilicon 1094 -2330 1094 -2330 0 3
rlabel polysilicon 1097 -2330 1097 -2330 0 4
rlabel polysilicon 1101 -2324 1101 -2324 0 1
rlabel polysilicon 1101 -2330 1101 -2330 0 3
rlabel polysilicon 1108 -2324 1108 -2324 0 1
rlabel polysilicon 1108 -2330 1108 -2330 0 3
rlabel polysilicon 1115 -2324 1115 -2324 0 1
rlabel polysilicon 1115 -2330 1115 -2330 0 3
rlabel polysilicon 1122 -2324 1122 -2324 0 1
rlabel polysilicon 1122 -2330 1122 -2330 0 3
rlabel polysilicon 1125 -2330 1125 -2330 0 4
rlabel polysilicon 1129 -2324 1129 -2324 0 1
rlabel polysilicon 1129 -2330 1129 -2330 0 3
rlabel polysilicon 1136 -2324 1136 -2324 0 1
rlabel polysilicon 1136 -2330 1136 -2330 0 3
rlabel polysilicon 1143 -2324 1143 -2324 0 1
rlabel polysilicon 1146 -2324 1146 -2324 0 2
rlabel polysilicon 1143 -2330 1143 -2330 0 3
rlabel polysilicon 1146 -2330 1146 -2330 0 4
rlabel polysilicon 1150 -2324 1150 -2324 0 1
rlabel polysilicon 1150 -2330 1150 -2330 0 3
rlabel polysilicon 1157 -2324 1157 -2324 0 1
rlabel polysilicon 1157 -2330 1157 -2330 0 3
rlabel polysilicon 1164 -2324 1164 -2324 0 1
rlabel polysilicon 1164 -2330 1164 -2330 0 3
rlabel polysilicon 1171 -2330 1171 -2330 0 3
rlabel polysilicon 1178 -2324 1178 -2324 0 1
rlabel polysilicon 1178 -2330 1178 -2330 0 3
rlabel polysilicon 1185 -2324 1185 -2324 0 1
rlabel polysilicon 1185 -2330 1185 -2330 0 3
rlabel polysilicon 1192 -2324 1192 -2324 0 1
rlabel polysilicon 1192 -2330 1192 -2330 0 3
rlabel polysilicon 1199 -2324 1199 -2324 0 1
rlabel polysilicon 1199 -2330 1199 -2330 0 3
rlabel polysilicon 1206 -2324 1206 -2324 0 1
rlabel polysilicon 1206 -2330 1206 -2330 0 3
rlabel polysilicon 1213 -2324 1213 -2324 0 1
rlabel polysilicon 1213 -2330 1213 -2330 0 3
rlabel polysilicon 1220 -2324 1220 -2324 0 1
rlabel polysilicon 1220 -2330 1220 -2330 0 3
rlabel polysilicon 1227 -2324 1227 -2324 0 1
rlabel polysilicon 1227 -2330 1227 -2330 0 3
rlabel polysilicon 1237 -2324 1237 -2324 0 2
rlabel polysilicon 1234 -2330 1234 -2330 0 3
rlabel polysilicon 1241 -2324 1241 -2324 0 1
rlabel polysilicon 1241 -2330 1241 -2330 0 3
rlabel polysilicon 1248 -2324 1248 -2324 0 1
rlabel polysilicon 1248 -2330 1248 -2330 0 3
rlabel polysilicon 1255 -2324 1255 -2324 0 1
rlabel polysilicon 1255 -2330 1255 -2330 0 3
rlabel polysilicon 1262 -2324 1262 -2324 0 1
rlabel polysilicon 1262 -2330 1262 -2330 0 3
rlabel polysilicon 1269 -2324 1269 -2324 0 1
rlabel polysilicon 1269 -2330 1269 -2330 0 3
rlabel polysilicon 1276 -2324 1276 -2324 0 1
rlabel polysilicon 1276 -2330 1276 -2330 0 3
rlabel polysilicon 1283 -2324 1283 -2324 0 1
rlabel polysilicon 1283 -2330 1283 -2330 0 3
rlabel polysilicon 1290 -2324 1290 -2324 0 1
rlabel polysilicon 1290 -2330 1290 -2330 0 3
rlabel polysilicon 1297 -2324 1297 -2324 0 1
rlabel polysilicon 1297 -2330 1297 -2330 0 3
rlabel polysilicon 1304 -2324 1304 -2324 0 1
rlabel polysilicon 1304 -2330 1304 -2330 0 3
rlabel polysilicon 1307 -2330 1307 -2330 0 4
rlabel polysilicon 1311 -2324 1311 -2324 0 1
rlabel polysilicon 1311 -2330 1311 -2330 0 3
rlabel polysilicon 1318 -2324 1318 -2324 0 1
rlabel polysilicon 1318 -2330 1318 -2330 0 3
rlabel polysilicon 1325 -2324 1325 -2324 0 1
rlabel polysilicon 1325 -2330 1325 -2330 0 3
rlabel polysilicon 1332 -2324 1332 -2324 0 1
rlabel polysilicon 1335 -2324 1335 -2324 0 2
rlabel polysilicon 1332 -2330 1332 -2330 0 3
rlabel polysilicon 1335 -2330 1335 -2330 0 4
rlabel polysilicon 1339 -2324 1339 -2324 0 1
rlabel polysilicon 1339 -2330 1339 -2330 0 3
rlabel polysilicon 1346 -2324 1346 -2324 0 1
rlabel polysilicon 1346 -2330 1346 -2330 0 3
rlabel polysilicon 1353 -2324 1353 -2324 0 1
rlabel polysilicon 1353 -2330 1353 -2330 0 3
rlabel polysilicon 1360 -2324 1360 -2324 0 1
rlabel polysilicon 1360 -2330 1360 -2330 0 3
rlabel polysilicon 1367 -2324 1367 -2324 0 1
rlabel polysilicon 1367 -2330 1367 -2330 0 3
rlabel polysilicon 1374 -2324 1374 -2324 0 1
rlabel polysilicon 1374 -2330 1374 -2330 0 3
rlabel polysilicon 1381 -2324 1381 -2324 0 1
rlabel polysilicon 1381 -2330 1381 -2330 0 3
rlabel polysilicon 1388 -2324 1388 -2324 0 1
rlabel polysilicon 1388 -2330 1388 -2330 0 3
rlabel polysilicon 1395 -2324 1395 -2324 0 1
rlabel polysilicon 1395 -2330 1395 -2330 0 3
rlabel polysilicon 1402 -2324 1402 -2324 0 1
rlabel polysilicon 1402 -2330 1402 -2330 0 3
rlabel polysilicon 1409 -2324 1409 -2324 0 1
rlabel polysilicon 1409 -2330 1409 -2330 0 3
rlabel polysilicon 1416 -2324 1416 -2324 0 1
rlabel polysilicon 1416 -2330 1416 -2330 0 3
rlabel polysilicon 1423 -2324 1423 -2324 0 1
rlabel polysilicon 1423 -2330 1423 -2330 0 3
rlabel polysilicon 1430 -2324 1430 -2324 0 1
rlabel polysilicon 1430 -2330 1430 -2330 0 3
rlabel polysilicon 1437 -2324 1437 -2324 0 1
rlabel polysilicon 1437 -2330 1437 -2330 0 3
rlabel polysilicon 1444 -2324 1444 -2324 0 1
rlabel polysilicon 1444 -2330 1444 -2330 0 3
rlabel polysilicon 1451 -2324 1451 -2324 0 1
rlabel polysilicon 1451 -2330 1451 -2330 0 3
rlabel polysilicon 1458 -2324 1458 -2324 0 1
rlabel polysilicon 1458 -2330 1458 -2330 0 3
rlabel polysilicon 1465 -2324 1465 -2324 0 1
rlabel polysilicon 1465 -2330 1465 -2330 0 3
rlabel polysilicon 1472 -2324 1472 -2324 0 1
rlabel polysilicon 1472 -2330 1472 -2330 0 3
rlabel polysilicon 1479 -2324 1479 -2324 0 1
rlabel polysilicon 1479 -2330 1479 -2330 0 3
rlabel polysilicon 1486 -2324 1486 -2324 0 1
rlabel polysilicon 1486 -2330 1486 -2330 0 3
rlabel polysilicon 1493 -2324 1493 -2324 0 1
rlabel polysilicon 1493 -2330 1493 -2330 0 3
rlabel polysilicon 1500 -2324 1500 -2324 0 1
rlabel polysilicon 1500 -2330 1500 -2330 0 3
rlabel polysilicon 1507 -2324 1507 -2324 0 1
rlabel polysilicon 1507 -2330 1507 -2330 0 3
rlabel polysilicon 1514 -2324 1514 -2324 0 1
rlabel polysilicon 1514 -2330 1514 -2330 0 3
rlabel polysilicon 1521 -2324 1521 -2324 0 1
rlabel polysilicon 1521 -2330 1521 -2330 0 3
rlabel polysilicon 1528 -2324 1528 -2324 0 1
rlabel polysilicon 1528 -2330 1528 -2330 0 3
rlabel polysilicon 1535 -2324 1535 -2324 0 1
rlabel polysilicon 1535 -2330 1535 -2330 0 3
rlabel polysilicon 1542 -2324 1542 -2324 0 1
rlabel polysilicon 1542 -2330 1542 -2330 0 3
rlabel polysilicon 1549 -2324 1549 -2324 0 1
rlabel polysilicon 1549 -2330 1549 -2330 0 3
rlabel polysilicon 1556 -2324 1556 -2324 0 1
rlabel polysilicon 1556 -2330 1556 -2330 0 3
rlabel polysilicon 1563 -2324 1563 -2324 0 1
rlabel polysilicon 1563 -2330 1563 -2330 0 3
rlabel polysilicon 1570 -2324 1570 -2324 0 1
rlabel polysilicon 1570 -2330 1570 -2330 0 3
rlabel polysilicon 1577 -2324 1577 -2324 0 1
rlabel polysilicon 1577 -2330 1577 -2330 0 3
rlabel polysilicon 1584 -2324 1584 -2324 0 1
rlabel polysilicon 1584 -2330 1584 -2330 0 3
rlabel polysilicon 1591 -2324 1591 -2324 0 1
rlabel polysilicon 1591 -2330 1591 -2330 0 3
rlabel polysilicon 1598 -2324 1598 -2324 0 1
rlabel polysilicon 1598 -2330 1598 -2330 0 3
rlabel polysilicon 1605 -2324 1605 -2324 0 1
rlabel polysilicon 1605 -2330 1605 -2330 0 3
rlabel polysilicon 1612 -2324 1612 -2324 0 1
rlabel polysilicon 1612 -2330 1612 -2330 0 3
rlabel polysilicon 1619 -2324 1619 -2324 0 1
rlabel polysilicon 1619 -2330 1619 -2330 0 3
rlabel polysilicon 1626 -2324 1626 -2324 0 1
rlabel polysilicon 1626 -2330 1626 -2330 0 3
rlabel polysilicon 1633 -2324 1633 -2324 0 1
rlabel polysilicon 1633 -2330 1633 -2330 0 3
rlabel polysilicon 1640 -2324 1640 -2324 0 1
rlabel polysilicon 1640 -2330 1640 -2330 0 3
rlabel polysilicon 1647 -2324 1647 -2324 0 1
rlabel polysilicon 1647 -2330 1647 -2330 0 3
rlabel polysilicon 1654 -2324 1654 -2324 0 1
rlabel polysilicon 1654 -2330 1654 -2330 0 3
rlabel polysilicon 1661 -2324 1661 -2324 0 1
rlabel polysilicon 1661 -2330 1661 -2330 0 3
rlabel polysilicon 1668 -2324 1668 -2324 0 1
rlabel polysilicon 1668 -2330 1668 -2330 0 3
rlabel polysilicon 1675 -2324 1675 -2324 0 1
rlabel polysilicon 1675 -2330 1675 -2330 0 3
rlabel polysilicon 1682 -2324 1682 -2324 0 1
rlabel polysilicon 1682 -2330 1682 -2330 0 3
rlabel polysilicon 1689 -2324 1689 -2324 0 1
rlabel polysilicon 1689 -2330 1689 -2330 0 3
rlabel polysilicon 1696 -2324 1696 -2324 0 1
rlabel polysilicon 1696 -2330 1696 -2330 0 3
rlabel polysilicon 1703 -2324 1703 -2324 0 1
rlabel polysilicon 1706 -2324 1706 -2324 0 2
rlabel polysilicon 1703 -2330 1703 -2330 0 3
rlabel polysilicon 1706 -2330 1706 -2330 0 4
rlabel polysilicon 1710 -2324 1710 -2324 0 1
rlabel polysilicon 1713 -2324 1713 -2324 0 2
rlabel polysilicon 1710 -2330 1710 -2330 0 3
rlabel polysilicon 1717 -2324 1717 -2324 0 1
rlabel polysilicon 1717 -2330 1717 -2330 0 3
rlabel polysilicon 1724 -2324 1724 -2324 0 1
rlabel polysilicon 1724 -2330 1724 -2330 0 3
rlabel polysilicon 1731 -2324 1731 -2324 0 1
rlabel polysilicon 1731 -2330 1731 -2330 0 3
rlabel polysilicon 1738 -2324 1738 -2324 0 1
rlabel polysilicon 1738 -2330 1738 -2330 0 3
rlabel polysilicon 51 -2439 51 -2439 0 1
rlabel polysilicon 51 -2445 51 -2445 0 3
rlabel polysilicon 58 -2439 58 -2439 0 1
rlabel polysilicon 58 -2445 58 -2445 0 3
rlabel polysilicon 65 -2439 65 -2439 0 1
rlabel polysilicon 65 -2445 65 -2445 0 3
rlabel polysilicon 72 -2439 72 -2439 0 1
rlabel polysilicon 72 -2445 72 -2445 0 3
rlabel polysilicon 79 -2439 79 -2439 0 1
rlabel polysilicon 79 -2445 79 -2445 0 3
rlabel polysilicon 86 -2439 86 -2439 0 1
rlabel polysilicon 86 -2445 86 -2445 0 3
rlabel polysilicon 93 -2439 93 -2439 0 1
rlabel polysilicon 93 -2445 93 -2445 0 3
rlabel polysilicon 100 -2439 100 -2439 0 1
rlabel polysilicon 100 -2445 100 -2445 0 3
rlabel polysilicon 107 -2439 107 -2439 0 1
rlabel polysilicon 107 -2445 107 -2445 0 3
rlabel polysilicon 114 -2439 114 -2439 0 1
rlabel polysilicon 114 -2445 114 -2445 0 3
rlabel polysilicon 121 -2439 121 -2439 0 1
rlabel polysilicon 121 -2445 121 -2445 0 3
rlabel polysilicon 128 -2439 128 -2439 0 1
rlabel polysilicon 128 -2445 128 -2445 0 3
rlabel polysilicon 135 -2439 135 -2439 0 1
rlabel polysilicon 135 -2445 135 -2445 0 3
rlabel polysilicon 142 -2439 142 -2439 0 1
rlabel polysilicon 142 -2445 142 -2445 0 3
rlabel polysilicon 149 -2439 149 -2439 0 1
rlabel polysilicon 149 -2445 149 -2445 0 3
rlabel polysilicon 156 -2439 156 -2439 0 1
rlabel polysilicon 156 -2445 156 -2445 0 3
rlabel polysilicon 163 -2439 163 -2439 0 1
rlabel polysilicon 163 -2445 163 -2445 0 3
rlabel polysilicon 170 -2439 170 -2439 0 1
rlabel polysilicon 170 -2445 170 -2445 0 3
rlabel polysilicon 177 -2439 177 -2439 0 1
rlabel polysilicon 180 -2439 180 -2439 0 2
rlabel polysilicon 180 -2445 180 -2445 0 4
rlabel polysilicon 184 -2439 184 -2439 0 1
rlabel polysilicon 184 -2445 184 -2445 0 3
rlabel polysilicon 191 -2439 191 -2439 0 1
rlabel polysilicon 191 -2445 191 -2445 0 3
rlabel polysilicon 198 -2439 198 -2439 0 1
rlabel polysilicon 198 -2445 198 -2445 0 3
rlabel polysilicon 205 -2439 205 -2439 0 1
rlabel polysilicon 205 -2445 205 -2445 0 3
rlabel polysilicon 212 -2439 212 -2439 0 1
rlabel polysilicon 215 -2439 215 -2439 0 2
rlabel polysilicon 212 -2445 212 -2445 0 3
rlabel polysilicon 215 -2445 215 -2445 0 4
rlabel polysilicon 219 -2439 219 -2439 0 1
rlabel polysilicon 219 -2445 219 -2445 0 3
rlabel polysilicon 226 -2439 226 -2439 0 1
rlabel polysilicon 226 -2445 226 -2445 0 3
rlabel polysilicon 233 -2439 233 -2439 0 1
rlabel polysilicon 233 -2445 233 -2445 0 3
rlabel polysilicon 240 -2439 240 -2439 0 1
rlabel polysilicon 240 -2445 240 -2445 0 3
rlabel polysilicon 247 -2439 247 -2439 0 1
rlabel polysilicon 247 -2445 247 -2445 0 3
rlabel polysilicon 254 -2439 254 -2439 0 1
rlabel polysilicon 257 -2445 257 -2445 0 4
rlabel polysilicon 261 -2439 261 -2439 0 1
rlabel polysilicon 261 -2445 261 -2445 0 3
rlabel polysilicon 268 -2439 268 -2439 0 1
rlabel polysilicon 268 -2445 268 -2445 0 3
rlabel polysilicon 275 -2439 275 -2439 0 1
rlabel polysilicon 275 -2445 275 -2445 0 3
rlabel polysilicon 282 -2439 282 -2439 0 1
rlabel polysilicon 282 -2445 282 -2445 0 3
rlabel polysilicon 289 -2439 289 -2439 0 1
rlabel polysilicon 289 -2445 289 -2445 0 3
rlabel polysilicon 296 -2439 296 -2439 0 1
rlabel polysilicon 296 -2445 296 -2445 0 3
rlabel polysilicon 303 -2439 303 -2439 0 1
rlabel polysilicon 303 -2445 303 -2445 0 3
rlabel polysilicon 310 -2439 310 -2439 0 1
rlabel polysilicon 313 -2445 313 -2445 0 4
rlabel polysilicon 317 -2439 317 -2439 0 1
rlabel polysilicon 317 -2445 317 -2445 0 3
rlabel polysilicon 324 -2439 324 -2439 0 1
rlabel polysilicon 324 -2445 324 -2445 0 3
rlabel polysilicon 331 -2439 331 -2439 0 1
rlabel polysilicon 331 -2445 331 -2445 0 3
rlabel polysilicon 338 -2439 338 -2439 0 1
rlabel polysilicon 338 -2445 338 -2445 0 3
rlabel polysilicon 345 -2439 345 -2439 0 1
rlabel polysilicon 345 -2445 345 -2445 0 3
rlabel polysilicon 352 -2439 352 -2439 0 1
rlabel polysilicon 352 -2445 352 -2445 0 3
rlabel polysilicon 359 -2439 359 -2439 0 1
rlabel polysilicon 359 -2445 359 -2445 0 3
rlabel polysilicon 366 -2439 366 -2439 0 1
rlabel polysilicon 366 -2445 366 -2445 0 3
rlabel polysilicon 373 -2439 373 -2439 0 1
rlabel polysilicon 373 -2445 373 -2445 0 3
rlabel polysilicon 380 -2439 380 -2439 0 1
rlabel polysilicon 380 -2445 380 -2445 0 3
rlabel polysilicon 387 -2439 387 -2439 0 1
rlabel polysilicon 387 -2445 387 -2445 0 3
rlabel polysilicon 394 -2439 394 -2439 0 1
rlabel polysilicon 394 -2445 394 -2445 0 3
rlabel polysilicon 401 -2439 401 -2439 0 1
rlabel polysilicon 401 -2445 401 -2445 0 3
rlabel polysilicon 408 -2439 408 -2439 0 1
rlabel polysilicon 408 -2445 408 -2445 0 3
rlabel polysilicon 415 -2439 415 -2439 0 1
rlabel polysilicon 415 -2445 415 -2445 0 3
rlabel polysilicon 422 -2439 422 -2439 0 1
rlabel polysilicon 422 -2445 422 -2445 0 3
rlabel polysilicon 432 -2439 432 -2439 0 2
rlabel polysilicon 429 -2445 429 -2445 0 3
rlabel polysilicon 432 -2445 432 -2445 0 4
rlabel polysilicon 436 -2439 436 -2439 0 1
rlabel polysilicon 436 -2445 436 -2445 0 3
rlabel polysilicon 443 -2439 443 -2439 0 1
rlabel polysilicon 443 -2445 443 -2445 0 3
rlabel polysilicon 450 -2439 450 -2439 0 1
rlabel polysilicon 450 -2445 450 -2445 0 3
rlabel polysilicon 457 -2439 457 -2439 0 1
rlabel polysilicon 457 -2445 457 -2445 0 3
rlabel polysilicon 464 -2439 464 -2439 0 1
rlabel polysilicon 464 -2445 464 -2445 0 3
rlabel polysilicon 471 -2439 471 -2439 0 1
rlabel polysilicon 474 -2439 474 -2439 0 2
rlabel polysilicon 474 -2445 474 -2445 0 4
rlabel polysilicon 478 -2439 478 -2439 0 1
rlabel polysilicon 478 -2445 478 -2445 0 3
rlabel polysilicon 485 -2439 485 -2439 0 1
rlabel polysilicon 485 -2445 485 -2445 0 3
rlabel polysilicon 492 -2439 492 -2439 0 1
rlabel polysilicon 492 -2445 492 -2445 0 3
rlabel polysilicon 499 -2439 499 -2439 0 1
rlabel polysilicon 502 -2439 502 -2439 0 2
rlabel polysilicon 499 -2445 499 -2445 0 3
rlabel polysilicon 502 -2445 502 -2445 0 4
rlabel polysilicon 506 -2439 506 -2439 0 1
rlabel polysilicon 506 -2445 506 -2445 0 3
rlabel polysilicon 513 -2439 513 -2439 0 1
rlabel polysilicon 513 -2445 513 -2445 0 3
rlabel polysilicon 520 -2439 520 -2439 0 1
rlabel polysilicon 520 -2445 520 -2445 0 3
rlabel polysilicon 530 -2439 530 -2439 0 2
rlabel polysilicon 527 -2445 527 -2445 0 3
rlabel polysilicon 530 -2445 530 -2445 0 4
rlabel polysilicon 534 -2439 534 -2439 0 1
rlabel polysilicon 534 -2445 534 -2445 0 3
rlabel polysilicon 541 -2439 541 -2439 0 1
rlabel polysilicon 541 -2445 541 -2445 0 3
rlabel polysilicon 548 -2439 548 -2439 0 1
rlabel polysilicon 548 -2445 548 -2445 0 3
rlabel polysilicon 555 -2439 555 -2439 0 1
rlabel polysilicon 555 -2445 555 -2445 0 3
rlabel polysilicon 562 -2439 562 -2439 0 1
rlabel polysilicon 562 -2445 562 -2445 0 3
rlabel polysilicon 569 -2439 569 -2439 0 1
rlabel polysilicon 569 -2445 569 -2445 0 3
rlabel polysilicon 576 -2439 576 -2439 0 1
rlabel polysilicon 576 -2445 576 -2445 0 3
rlabel polysilicon 583 -2439 583 -2439 0 1
rlabel polysilicon 583 -2445 583 -2445 0 3
rlabel polysilicon 590 -2439 590 -2439 0 1
rlabel polysilicon 590 -2445 590 -2445 0 3
rlabel polysilicon 597 -2439 597 -2439 0 1
rlabel polysilicon 597 -2445 597 -2445 0 3
rlabel polysilicon 604 -2439 604 -2439 0 1
rlabel polysilicon 604 -2445 604 -2445 0 3
rlabel polysilicon 611 -2439 611 -2439 0 1
rlabel polysilicon 614 -2439 614 -2439 0 2
rlabel polysilicon 611 -2445 611 -2445 0 3
rlabel polysilicon 618 -2439 618 -2439 0 1
rlabel polysilicon 618 -2445 618 -2445 0 3
rlabel polysilicon 625 -2439 625 -2439 0 1
rlabel polysilicon 625 -2445 625 -2445 0 3
rlabel polysilicon 632 -2439 632 -2439 0 1
rlabel polysilicon 632 -2445 632 -2445 0 3
rlabel polysilicon 639 -2439 639 -2439 0 1
rlabel polysilicon 642 -2445 642 -2445 0 4
rlabel polysilicon 646 -2439 646 -2439 0 1
rlabel polysilicon 646 -2445 646 -2445 0 3
rlabel polysilicon 653 -2439 653 -2439 0 1
rlabel polysilicon 653 -2445 653 -2445 0 3
rlabel polysilicon 660 -2439 660 -2439 0 1
rlabel polysilicon 660 -2445 660 -2445 0 3
rlabel polysilicon 667 -2439 667 -2439 0 1
rlabel polysilicon 667 -2445 667 -2445 0 3
rlabel polysilicon 674 -2439 674 -2439 0 1
rlabel polysilicon 677 -2439 677 -2439 0 2
rlabel polysilicon 674 -2445 674 -2445 0 3
rlabel polysilicon 677 -2445 677 -2445 0 4
rlabel polysilicon 684 -2439 684 -2439 0 2
rlabel polysilicon 681 -2445 681 -2445 0 3
rlabel polysilicon 684 -2445 684 -2445 0 4
rlabel polysilicon 688 -2439 688 -2439 0 1
rlabel polysilicon 688 -2445 688 -2445 0 3
rlabel polysilicon 695 -2439 695 -2439 0 1
rlabel polysilicon 695 -2445 695 -2445 0 3
rlabel polysilicon 705 -2439 705 -2439 0 2
rlabel polysilicon 705 -2445 705 -2445 0 4
rlabel polysilicon 709 -2439 709 -2439 0 1
rlabel polysilicon 709 -2445 709 -2445 0 3
rlabel polysilicon 716 -2439 716 -2439 0 1
rlabel polysilicon 716 -2445 716 -2445 0 3
rlabel polysilicon 723 -2439 723 -2439 0 1
rlabel polysilicon 723 -2445 723 -2445 0 3
rlabel polysilicon 730 -2439 730 -2439 0 1
rlabel polysilicon 733 -2439 733 -2439 0 2
rlabel polysilicon 730 -2445 730 -2445 0 3
rlabel polysilicon 733 -2445 733 -2445 0 4
rlabel polysilicon 737 -2439 737 -2439 0 1
rlabel polysilicon 737 -2445 737 -2445 0 3
rlabel polysilicon 744 -2439 744 -2439 0 1
rlabel polysilicon 747 -2439 747 -2439 0 2
rlabel polysilicon 747 -2445 747 -2445 0 4
rlabel polysilicon 751 -2439 751 -2439 0 1
rlabel polysilicon 751 -2445 751 -2445 0 3
rlabel polysilicon 758 -2439 758 -2439 0 1
rlabel polysilicon 758 -2445 758 -2445 0 3
rlabel polysilicon 765 -2439 765 -2439 0 1
rlabel polysilicon 765 -2445 765 -2445 0 3
rlabel polysilicon 772 -2439 772 -2439 0 1
rlabel polysilicon 772 -2445 772 -2445 0 3
rlabel polysilicon 779 -2439 779 -2439 0 1
rlabel polysilicon 779 -2445 779 -2445 0 3
rlabel polysilicon 786 -2439 786 -2439 0 1
rlabel polysilicon 786 -2445 786 -2445 0 3
rlabel polysilicon 793 -2439 793 -2439 0 1
rlabel polysilicon 793 -2445 793 -2445 0 3
rlabel polysilicon 800 -2439 800 -2439 0 1
rlabel polysilicon 800 -2445 800 -2445 0 3
rlabel polysilicon 807 -2439 807 -2439 0 1
rlabel polysilicon 810 -2439 810 -2439 0 2
rlabel polysilicon 807 -2445 807 -2445 0 3
rlabel polysilicon 810 -2445 810 -2445 0 4
rlabel polysilicon 814 -2439 814 -2439 0 1
rlabel polysilicon 814 -2445 814 -2445 0 3
rlabel polysilicon 821 -2439 821 -2439 0 1
rlabel polysilicon 824 -2439 824 -2439 0 2
rlabel polysilicon 821 -2445 821 -2445 0 3
rlabel polysilicon 824 -2445 824 -2445 0 4
rlabel polysilicon 828 -2439 828 -2439 0 1
rlabel polysilicon 828 -2445 828 -2445 0 3
rlabel polysilicon 835 -2439 835 -2439 0 1
rlabel polysilicon 835 -2445 835 -2445 0 3
rlabel polysilicon 842 -2439 842 -2439 0 1
rlabel polysilicon 845 -2439 845 -2439 0 2
rlabel polysilicon 845 -2445 845 -2445 0 4
rlabel polysilicon 849 -2439 849 -2439 0 1
rlabel polysilicon 852 -2439 852 -2439 0 2
rlabel polysilicon 849 -2445 849 -2445 0 3
rlabel polysilicon 852 -2445 852 -2445 0 4
rlabel polysilicon 856 -2439 856 -2439 0 1
rlabel polysilicon 856 -2445 856 -2445 0 3
rlabel polysilicon 859 -2445 859 -2445 0 4
rlabel polysilicon 863 -2439 863 -2439 0 1
rlabel polysilicon 863 -2445 863 -2445 0 3
rlabel polysilicon 870 -2439 870 -2439 0 1
rlabel polysilicon 870 -2445 870 -2445 0 3
rlabel polysilicon 877 -2439 877 -2439 0 1
rlabel polysilicon 877 -2445 877 -2445 0 3
rlabel polysilicon 884 -2439 884 -2439 0 1
rlabel polysilicon 884 -2445 884 -2445 0 3
rlabel polysilicon 891 -2439 891 -2439 0 1
rlabel polysilicon 891 -2445 891 -2445 0 3
rlabel polysilicon 894 -2445 894 -2445 0 4
rlabel polysilicon 898 -2439 898 -2439 0 1
rlabel polysilicon 901 -2439 901 -2439 0 2
rlabel polysilicon 898 -2445 898 -2445 0 3
rlabel polysilicon 901 -2445 901 -2445 0 4
rlabel polysilicon 905 -2439 905 -2439 0 1
rlabel polysilicon 905 -2445 905 -2445 0 3
rlabel polysilicon 912 -2439 912 -2439 0 1
rlabel polysilicon 912 -2445 912 -2445 0 3
rlabel polysilicon 919 -2439 919 -2439 0 1
rlabel polysilicon 919 -2445 919 -2445 0 3
rlabel polysilicon 926 -2439 926 -2439 0 1
rlabel polysilicon 926 -2445 926 -2445 0 3
rlabel polysilicon 933 -2439 933 -2439 0 1
rlabel polysilicon 933 -2445 933 -2445 0 3
rlabel polysilicon 940 -2439 940 -2439 0 1
rlabel polysilicon 940 -2445 940 -2445 0 3
rlabel polysilicon 947 -2439 947 -2439 0 1
rlabel polysilicon 947 -2445 947 -2445 0 3
rlabel polysilicon 954 -2439 954 -2439 0 1
rlabel polysilicon 954 -2445 954 -2445 0 3
rlabel polysilicon 961 -2439 961 -2439 0 1
rlabel polysilicon 961 -2445 961 -2445 0 3
rlabel polysilicon 968 -2439 968 -2439 0 1
rlabel polysilicon 971 -2439 971 -2439 0 2
rlabel polysilicon 968 -2445 968 -2445 0 3
rlabel polysilicon 971 -2445 971 -2445 0 4
rlabel polysilicon 975 -2439 975 -2439 0 1
rlabel polysilicon 975 -2445 975 -2445 0 3
rlabel polysilicon 982 -2439 982 -2439 0 1
rlabel polysilicon 982 -2445 982 -2445 0 3
rlabel polysilicon 989 -2439 989 -2439 0 1
rlabel polysilicon 989 -2445 989 -2445 0 3
rlabel polysilicon 996 -2439 996 -2439 0 1
rlabel polysilicon 996 -2445 996 -2445 0 3
rlabel polysilicon 1003 -2439 1003 -2439 0 1
rlabel polysilicon 1003 -2445 1003 -2445 0 3
rlabel polysilicon 1010 -2439 1010 -2439 0 1
rlabel polysilicon 1010 -2445 1010 -2445 0 3
rlabel polysilicon 1017 -2439 1017 -2439 0 1
rlabel polysilicon 1017 -2445 1017 -2445 0 3
rlabel polysilicon 1024 -2439 1024 -2439 0 1
rlabel polysilicon 1024 -2445 1024 -2445 0 3
rlabel polysilicon 1031 -2439 1031 -2439 0 1
rlabel polysilicon 1031 -2445 1031 -2445 0 3
rlabel polysilicon 1038 -2439 1038 -2439 0 1
rlabel polysilicon 1038 -2445 1038 -2445 0 3
rlabel polysilicon 1045 -2439 1045 -2439 0 1
rlabel polysilicon 1045 -2445 1045 -2445 0 3
rlabel polysilicon 1052 -2439 1052 -2439 0 1
rlabel polysilicon 1052 -2445 1052 -2445 0 3
rlabel polysilicon 1059 -2439 1059 -2439 0 1
rlabel polysilicon 1059 -2445 1059 -2445 0 3
rlabel polysilicon 1066 -2439 1066 -2439 0 1
rlabel polysilicon 1066 -2445 1066 -2445 0 3
rlabel polysilicon 1073 -2439 1073 -2439 0 1
rlabel polysilicon 1076 -2439 1076 -2439 0 2
rlabel polysilicon 1073 -2445 1073 -2445 0 3
rlabel polysilicon 1076 -2445 1076 -2445 0 4
rlabel polysilicon 1080 -2439 1080 -2439 0 1
rlabel polysilicon 1080 -2445 1080 -2445 0 3
rlabel polysilicon 1087 -2439 1087 -2439 0 1
rlabel polysilicon 1087 -2445 1087 -2445 0 3
rlabel polysilicon 1094 -2439 1094 -2439 0 1
rlabel polysilicon 1094 -2445 1094 -2445 0 3
rlabel polysilicon 1101 -2439 1101 -2439 0 1
rlabel polysilicon 1101 -2445 1101 -2445 0 3
rlabel polysilicon 1108 -2439 1108 -2439 0 1
rlabel polysilicon 1108 -2445 1108 -2445 0 3
rlabel polysilicon 1115 -2439 1115 -2439 0 1
rlabel polysilicon 1115 -2445 1115 -2445 0 3
rlabel polysilicon 1122 -2439 1122 -2439 0 1
rlabel polysilicon 1122 -2445 1122 -2445 0 3
rlabel polysilicon 1129 -2439 1129 -2439 0 1
rlabel polysilicon 1129 -2445 1129 -2445 0 3
rlabel polysilicon 1136 -2439 1136 -2439 0 1
rlabel polysilicon 1136 -2445 1136 -2445 0 3
rlabel polysilicon 1143 -2439 1143 -2439 0 1
rlabel polysilicon 1143 -2445 1143 -2445 0 3
rlabel polysilicon 1150 -2439 1150 -2439 0 1
rlabel polysilicon 1150 -2445 1150 -2445 0 3
rlabel polysilicon 1157 -2439 1157 -2439 0 1
rlabel polysilicon 1157 -2445 1157 -2445 0 3
rlabel polysilicon 1164 -2439 1164 -2439 0 1
rlabel polysilicon 1164 -2445 1164 -2445 0 3
rlabel polysilicon 1171 -2439 1171 -2439 0 1
rlabel polysilicon 1171 -2445 1171 -2445 0 3
rlabel polysilicon 1178 -2439 1178 -2439 0 1
rlabel polysilicon 1178 -2445 1178 -2445 0 3
rlabel polysilicon 1185 -2439 1185 -2439 0 1
rlabel polysilicon 1185 -2445 1185 -2445 0 3
rlabel polysilicon 1192 -2439 1192 -2439 0 1
rlabel polysilicon 1195 -2439 1195 -2439 0 2
rlabel polysilicon 1192 -2445 1192 -2445 0 3
rlabel polysilicon 1195 -2445 1195 -2445 0 4
rlabel polysilicon 1199 -2439 1199 -2439 0 1
rlabel polysilicon 1199 -2445 1199 -2445 0 3
rlabel polysilicon 1206 -2439 1206 -2439 0 1
rlabel polysilicon 1206 -2445 1206 -2445 0 3
rlabel polysilicon 1209 -2445 1209 -2445 0 4
rlabel polysilicon 1213 -2439 1213 -2439 0 1
rlabel polysilicon 1213 -2445 1213 -2445 0 3
rlabel polysilicon 1220 -2439 1220 -2439 0 1
rlabel polysilicon 1220 -2445 1220 -2445 0 3
rlabel polysilicon 1227 -2439 1227 -2439 0 1
rlabel polysilicon 1227 -2445 1227 -2445 0 3
rlabel polysilicon 1234 -2439 1234 -2439 0 1
rlabel polysilicon 1234 -2445 1234 -2445 0 3
rlabel polysilicon 1241 -2439 1241 -2439 0 1
rlabel polysilicon 1244 -2439 1244 -2439 0 2
rlabel polysilicon 1244 -2445 1244 -2445 0 4
rlabel polysilicon 1248 -2439 1248 -2439 0 1
rlabel polysilicon 1248 -2445 1248 -2445 0 3
rlabel polysilicon 1255 -2439 1255 -2439 0 1
rlabel polysilicon 1255 -2445 1255 -2445 0 3
rlabel polysilicon 1262 -2439 1262 -2439 0 1
rlabel polysilicon 1262 -2445 1262 -2445 0 3
rlabel polysilicon 1269 -2439 1269 -2439 0 1
rlabel polysilicon 1269 -2445 1269 -2445 0 3
rlabel polysilicon 1276 -2439 1276 -2439 0 1
rlabel polysilicon 1276 -2445 1276 -2445 0 3
rlabel polysilicon 1283 -2439 1283 -2439 0 1
rlabel polysilicon 1283 -2445 1283 -2445 0 3
rlabel polysilicon 1290 -2439 1290 -2439 0 1
rlabel polysilicon 1290 -2445 1290 -2445 0 3
rlabel polysilicon 1297 -2445 1297 -2445 0 3
rlabel polysilicon 1300 -2445 1300 -2445 0 4
rlabel polysilicon 1304 -2439 1304 -2439 0 1
rlabel polysilicon 1304 -2445 1304 -2445 0 3
rlabel polysilicon 1314 -2439 1314 -2439 0 2
rlabel polysilicon 1311 -2445 1311 -2445 0 3
rlabel polysilicon 1314 -2445 1314 -2445 0 4
rlabel polysilicon 1318 -2439 1318 -2439 0 1
rlabel polysilicon 1318 -2445 1318 -2445 0 3
rlabel polysilicon 1325 -2439 1325 -2439 0 1
rlabel polysilicon 1325 -2445 1325 -2445 0 3
rlabel polysilicon 1332 -2439 1332 -2439 0 1
rlabel polysilicon 1332 -2445 1332 -2445 0 3
rlabel polysilicon 1339 -2439 1339 -2439 0 1
rlabel polysilicon 1339 -2445 1339 -2445 0 3
rlabel polysilicon 1346 -2439 1346 -2439 0 1
rlabel polysilicon 1346 -2445 1346 -2445 0 3
rlabel polysilicon 1353 -2439 1353 -2439 0 1
rlabel polysilicon 1353 -2445 1353 -2445 0 3
rlabel polysilicon 1360 -2439 1360 -2439 0 1
rlabel polysilicon 1360 -2445 1360 -2445 0 3
rlabel polysilicon 1367 -2439 1367 -2439 0 1
rlabel polysilicon 1367 -2445 1367 -2445 0 3
rlabel polysilicon 1374 -2439 1374 -2439 0 1
rlabel polysilicon 1374 -2445 1374 -2445 0 3
rlabel polysilicon 1381 -2439 1381 -2439 0 1
rlabel polysilicon 1384 -2439 1384 -2439 0 2
rlabel polysilicon 1381 -2445 1381 -2445 0 3
rlabel polysilicon 1388 -2439 1388 -2439 0 1
rlabel polysilicon 1388 -2445 1388 -2445 0 3
rlabel polysilicon 1395 -2439 1395 -2439 0 1
rlabel polysilicon 1395 -2445 1395 -2445 0 3
rlabel polysilicon 1402 -2439 1402 -2439 0 1
rlabel polysilicon 1402 -2445 1402 -2445 0 3
rlabel polysilicon 1409 -2439 1409 -2439 0 1
rlabel polysilicon 1409 -2445 1409 -2445 0 3
rlabel polysilicon 1416 -2439 1416 -2439 0 1
rlabel polysilicon 1416 -2445 1416 -2445 0 3
rlabel polysilicon 1423 -2439 1423 -2439 0 1
rlabel polysilicon 1423 -2445 1423 -2445 0 3
rlabel polysilicon 1430 -2439 1430 -2439 0 1
rlabel polysilicon 1430 -2445 1430 -2445 0 3
rlabel polysilicon 1437 -2439 1437 -2439 0 1
rlabel polysilicon 1437 -2445 1437 -2445 0 3
rlabel polysilicon 1444 -2439 1444 -2439 0 1
rlabel polysilicon 1444 -2445 1444 -2445 0 3
rlabel polysilicon 1451 -2439 1451 -2439 0 1
rlabel polysilicon 1451 -2445 1451 -2445 0 3
rlabel polysilicon 1458 -2439 1458 -2439 0 1
rlabel polysilicon 1458 -2445 1458 -2445 0 3
rlabel polysilicon 1465 -2439 1465 -2439 0 1
rlabel polysilicon 1465 -2445 1465 -2445 0 3
rlabel polysilicon 1472 -2439 1472 -2439 0 1
rlabel polysilicon 1472 -2445 1472 -2445 0 3
rlabel polysilicon 1479 -2439 1479 -2439 0 1
rlabel polysilicon 1479 -2445 1479 -2445 0 3
rlabel polysilicon 1486 -2439 1486 -2439 0 1
rlabel polysilicon 1486 -2445 1486 -2445 0 3
rlabel polysilicon 1493 -2439 1493 -2439 0 1
rlabel polysilicon 1493 -2445 1493 -2445 0 3
rlabel polysilicon 1500 -2439 1500 -2439 0 1
rlabel polysilicon 1500 -2445 1500 -2445 0 3
rlabel polysilicon 1507 -2439 1507 -2439 0 1
rlabel polysilicon 1507 -2445 1507 -2445 0 3
rlabel polysilicon 1514 -2439 1514 -2439 0 1
rlabel polysilicon 1514 -2445 1514 -2445 0 3
rlabel polysilicon 1521 -2439 1521 -2439 0 1
rlabel polysilicon 1521 -2445 1521 -2445 0 3
rlabel polysilicon 1528 -2439 1528 -2439 0 1
rlabel polysilicon 1528 -2445 1528 -2445 0 3
rlabel polysilicon 1538 -2439 1538 -2439 0 2
rlabel polysilicon 1535 -2445 1535 -2445 0 3
rlabel polysilicon 1538 -2445 1538 -2445 0 4
rlabel polysilicon 1542 -2439 1542 -2439 0 1
rlabel polysilicon 1542 -2445 1542 -2445 0 3
rlabel polysilicon 1549 -2439 1549 -2439 0 1
rlabel polysilicon 1549 -2445 1549 -2445 0 3
rlabel polysilicon 1556 -2439 1556 -2439 0 1
rlabel polysilicon 1556 -2445 1556 -2445 0 3
rlabel polysilicon 1563 -2439 1563 -2439 0 1
rlabel polysilicon 1563 -2445 1563 -2445 0 3
rlabel polysilicon 1570 -2439 1570 -2439 0 1
rlabel polysilicon 1570 -2445 1570 -2445 0 3
rlabel polysilicon 1577 -2439 1577 -2439 0 1
rlabel polysilicon 1577 -2445 1577 -2445 0 3
rlabel polysilicon 1580 -2445 1580 -2445 0 4
rlabel polysilicon 1584 -2439 1584 -2439 0 1
rlabel polysilicon 1584 -2445 1584 -2445 0 3
rlabel polysilicon 1591 -2439 1591 -2439 0 1
rlabel polysilicon 1591 -2445 1591 -2445 0 3
rlabel polysilicon 1598 -2439 1598 -2439 0 1
rlabel polysilicon 1598 -2445 1598 -2445 0 3
rlabel polysilicon 1605 -2439 1605 -2439 0 1
rlabel polysilicon 1605 -2445 1605 -2445 0 3
rlabel polysilicon 1675 -2439 1675 -2439 0 1
rlabel polysilicon 1675 -2445 1675 -2445 0 3
rlabel polysilicon 44 -2556 44 -2556 0 1
rlabel polysilicon 44 -2562 44 -2562 0 3
rlabel polysilicon 51 -2556 51 -2556 0 1
rlabel polysilicon 51 -2562 51 -2562 0 3
rlabel polysilicon 58 -2556 58 -2556 0 1
rlabel polysilicon 58 -2562 58 -2562 0 3
rlabel polysilicon 65 -2556 65 -2556 0 1
rlabel polysilicon 68 -2556 68 -2556 0 2
rlabel polysilicon 75 -2556 75 -2556 0 2
rlabel polysilicon 72 -2562 72 -2562 0 3
rlabel polysilicon 75 -2562 75 -2562 0 4
rlabel polysilicon 79 -2556 79 -2556 0 1
rlabel polysilicon 79 -2562 79 -2562 0 3
rlabel polysilicon 86 -2556 86 -2556 0 1
rlabel polysilicon 86 -2562 86 -2562 0 3
rlabel polysilicon 93 -2556 93 -2556 0 1
rlabel polysilicon 93 -2562 93 -2562 0 3
rlabel polysilicon 100 -2556 100 -2556 0 1
rlabel polysilicon 103 -2556 103 -2556 0 2
rlabel polysilicon 100 -2562 100 -2562 0 3
rlabel polysilicon 107 -2556 107 -2556 0 1
rlabel polysilicon 107 -2562 107 -2562 0 3
rlabel polysilicon 114 -2556 114 -2556 0 1
rlabel polysilicon 114 -2562 114 -2562 0 3
rlabel polysilicon 121 -2556 121 -2556 0 1
rlabel polysilicon 121 -2562 121 -2562 0 3
rlabel polysilicon 128 -2556 128 -2556 0 1
rlabel polysilicon 128 -2562 128 -2562 0 3
rlabel polysilicon 135 -2556 135 -2556 0 1
rlabel polysilicon 135 -2562 135 -2562 0 3
rlabel polysilicon 142 -2556 142 -2556 0 1
rlabel polysilicon 142 -2562 142 -2562 0 3
rlabel polysilicon 149 -2556 149 -2556 0 1
rlabel polysilicon 152 -2556 152 -2556 0 2
rlabel polysilicon 149 -2562 149 -2562 0 3
rlabel polysilicon 152 -2562 152 -2562 0 4
rlabel polysilicon 156 -2556 156 -2556 0 1
rlabel polysilicon 156 -2562 156 -2562 0 3
rlabel polysilicon 163 -2556 163 -2556 0 1
rlabel polysilicon 166 -2556 166 -2556 0 2
rlabel polysilicon 163 -2562 163 -2562 0 3
rlabel polysilicon 166 -2562 166 -2562 0 4
rlabel polysilicon 173 -2556 173 -2556 0 2
rlabel polysilicon 170 -2562 170 -2562 0 3
rlabel polysilicon 177 -2556 177 -2556 0 1
rlabel polysilicon 177 -2562 177 -2562 0 3
rlabel polysilicon 184 -2556 184 -2556 0 1
rlabel polysilicon 184 -2562 184 -2562 0 3
rlabel polysilicon 191 -2556 191 -2556 0 1
rlabel polysilicon 191 -2562 191 -2562 0 3
rlabel polysilicon 198 -2556 198 -2556 0 1
rlabel polysilicon 198 -2562 198 -2562 0 3
rlabel polysilicon 205 -2556 205 -2556 0 1
rlabel polysilicon 205 -2562 205 -2562 0 3
rlabel polysilicon 212 -2556 212 -2556 0 1
rlabel polysilicon 212 -2562 212 -2562 0 3
rlabel polysilicon 219 -2556 219 -2556 0 1
rlabel polysilicon 219 -2562 219 -2562 0 3
rlabel polysilicon 226 -2556 226 -2556 0 1
rlabel polysilicon 226 -2562 226 -2562 0 3
rlabel polysilicon 233 -2556 233 -2556 0 1
rlabel polysilicon 233 -2562 233 -2562 0 3
rlabel polysilicon 240 -2556 240 -2556 0 1
rlabel polysilicon 240 -2562 240 -2562 0 3
rlabel polysilicon 247 -2556 247 -2556 0 1
rlabel polysilicon 247 -2562 247 -2562 0 3
rlabel polysilicon 254 -2562 254 -2562 0 3
rlabel polysilicon 257 -2562 257 -2562 0 4
rlabel polysilicon 261 -2556 261 -2556 0 1
rlabel polysilicon 261 -2562 261 -2562 0 3
rlabel polysilicon 268 -2556 268 -2556 0 1
rlabel polysilicon 268 -2562 268 -2562 0 3
rlabel polysilicon 275 -2556 275 -2556 0 1
rlabel polysilicon 275 -2562 275 -2562 0 3
rlabel polysilicon 282 -2556 282 -2556 0 1
rlabel polysilicon 282 -2562 282 -2562 0 3
rlabel polysilicon 289 -2556 289 -2556 0 1
rlabel polysilicon 289 -2562 289 -2562 0 3
rlabel polysilicon 296 -2556 296 -2556 0 1
rlabel polysilicon 296 -2562 296 -2562 0 3
rlabel polysilicon 303 -2556 303 -2556 0 1
rlabel polysilicon 303 -2562 303 -2562 0 3
rlabel polysilicon 310 -2556 310 -2556 0 1
rlabel polysilicon 310 -2562 310 -2562 0 3
rlabel polysilicon 317 -2556 317 -2556 0 1
rlabel polysilicon 317 -2562 317 -2562 0 3
rlabel polysilicon 324 -2556 324 -2556 0 1
rlabel polysilicon 324 -2562 324 -2562 0 3
rlabel polysilicon 331 -2556 331 -2556 0 1
rlabel polysilicon 331 -2562 331 -2562 0 3
rlabel polysilicon 338 -2556 338 -2556 0 1
rlabel polysilicon 338 -2562 338 -2562 0 3
rlabel polysilicon 345 -2556 345 -2556 0 1
rlabel polysilicon 345 -2562 345 -2562 0 3
rlabel polysilicon 352 -2556 352 -2556 0 1
rlabel polysilicon 352 -2562 352 -2562 0 3
rlabel polysilicon 359 -2556 359 -2556 0 1
rlabel polysilicon 359 -2562 359 -2562 0 3
rlabel polysilicon 366 -2556 366 -2556 0 1
rlabel polysilicon 366 -2562 366 -2562 0 3
rlabel polysilicon 373 -2556 373 -2556 0 1
rlabel polysilicon 373 -2562 373 -2562 0 3
rlabel polysilicon 380 -2556 380 -2556 0 1
rlabel polysilicon 380 -2562 380 -2562 0 3
rlabel polysilicon 387 -2556 387 -2556 0 1
rlabel polysilicon 387 -2562 387 -2562 0 3
rlabel polysilicon 394 -2556 394 -2556 0 1
rlabel polysilicon 394 -2562 394 -2562 0 3
rlabel polysilicon 401 -2556 401 -2556 0 1
rlabel polysilicon 401 -2562 401 -2562 0 3
rlabel polysilicon 408 -2556 408 -2556 0 1
rlabel polysilicon 411 -2556 411 -2556 0 2
rlabel polysilicon 408 -2562 408 -2562 0 3
rlabel polysilicon 415 -2556 415 -2556 0 1
rlabel polysilicon 415 -2562 415 -2562 0 3
rlabel polysilicon 422 -2556 422 -2556 0 1
rlabel polysilicon 422 -2562 422 -2562 0 3
rlabel polysilicon 432 -2556 432 -2556 0 2
rlabel polysilicon 429 -2562 429 -2562 0 3
rlabel polysilicon 432 -2562 432 -2562 0 4
rlabel polysilicon 436 -2556 436 -2556 0 1
rlabel polysilicon 436 -2562 436 -2562 0 3
rlabel polysilicon 443 -2556 443 -2556 0 1
rlabel polysilicon 446 -2556 446 -2556 0 2
rlabel polysilicon 443 -2562 443 -2562 0 3
rlabel polysilicon 446 -2562 446 -2562 0 4
rlabel polysilicon 450 -2556 450 -2556 0 1
rlabel polysilicon 450 -2562 450 -2562 0 3
rlabel polysilicon 457 -2556 457 -2556 0 1
rlabel polysilicon 457 -2562 457 -2562 0 3
rlabel polysilicon 464 -2556 464 -2556 0 1
rlabel polysilicon 464 -2562 464 -2562 0 3
rlabel polysilicon 471 -2556 471 -2556 0 1
rlabel polysilicon 471 -2562 471 -2562 0 3
rlabel polysilicon 478 -2556 478 -2556 0 1
rlabel polysilicon 478 -2562 478 -2562 0 3
rlabel polysilicon 485 -2556 485 -2556 0 1
rlabel polysilicon 485 -2562 485 -2562 0 3
rlabel polysilicon 492 -2556 492 -2556 0 1
rlabel polysilicon 492 -2562 492 -2562 0 3
rlabel polysilicon 499 -2556 499 -2556 0 1
rlabel polysilicon 499 -2562 499 -2562 0 3
rlabel polysilicon 506 -2556 506 -2556 0 1
rlabel polysilicon 506 -2562 506 -2562 0 3
rlabel polysilicon 513 -2556 513 -2556 0 1
rlabel polysilicon 513 -2562 513 -2562 0 3
rlabel polysilicon 520 -2556 520 -2556 0 1
rlabel polysilicon 520 -2562 520 -2562 0 3
rlabel polysilicon 527 -2556 527 -2556 0 1
rlabel polysilicon 527 -2562 527 -2562 0 3
rlabel polysilicon 534 -2556 534 -2556 0 1
rlabel polysilicon 534 -2562 534 -2562 0 3
rlabel polysilicon 541 -2556 541 -2556 0 1
rlabel polysilicon 541 -2562 541 -2562 0 3
rlabel polysilicon 548 -2556 548 -2556 0 1
rlabel polysilicon 551 -2556 551 -2556 0 2
rlabel polysilicon 548 -2562 548 -2562 0 3
rlabel polysilicon 551 -2562 551 -2562 0 4
rlabel polysilicon 555 -2556 555 -2556 0 1
rlabel polysilicon 555 -2562 555 -2562 0 3
rlabel polysilicon 562 -2556 562 -2556 0 1
rlabel polysilicon 562 -2562 562 -2562 0 3
rlabel polysilicon 569 -2556 569 -2556 0 1
rlabel polysilicon 569 -2562 569 -2562 0 3
rlabel polysilicon 576 -2556 576 -2556 0 1
rlabel polysilicon 576 -2562 576 -2562 0 3
rlabel polysilicon 583 -2556 583 -2556 0 1
rlabel polysilicon 583 -2562 583 -2562 0 3
rlabel polysilicon 590 -2556 590 -2556 0 1
rlabel polysilicon 593 -2556 593 -2556 0 2
rlabel polysilicon 590 -2562 590 -2562 0 3
rlabel polysilicon 593 -2562 593 -2562 0 4
rlabel polysilicon 597 -2556 597 -2556 0 1
rlabel polysilicon 597 -2562 597 -2562 0 3
rlabel polysilicon 604 -2556 604 -2556 0 1
rlabel polysilicon 604 -2562 604 -2562 0 3
rlabel polysilicon 611 -2556 611 -2556 0 1
rlabel polysilicon 611 -2562 611 -2562 0 3
rlabel polysilicon 618 -2556 618 -2556 0 1
rlabel polysilicon 618 -2562 618 -2562 0 3
rlabel polysilicon 625 -2556 625 -2556 0 1
rlabel polysilicon 628 -2556 628 -2556 0 2
rlabel polysilicon 625 -2562 625 -2562 0 3
rlabel polysilicon 632 -2556 632 -2556 0 1
rlabel polysilicon 632 -2562 632 -2562 0 3
rlabel polysilicon 639 -2556 639 -2556 0 1
rlabel polysilicon 639 -2562 639 -2562 0 3
rlabel polysilicon 646 -2556 646 -2556 0 1
rlabel polysilicon 649 -2556 649 -2556 0 2
rlabel polysilicon 646 -2562 646 -2562 0 3
rlabel polysilicon 649 -2562 649 -2562 0 4
rlabel polysilicon 653 -2556 653 -2556 0 1
rlabel polysilicon 653 -2562 653 -2562 0 3
rlabel polysilicon 660 -2556 660 -2556 0 1
rlabel polysilicon 663 -2556 663 -2556 0 2
rlabel polysilicon 660 -2562 660 -2562 0 3
rlabel polysilicon 663 -2562 663 -2562 0 4
rlabel polysilicon 667 -2556 667 -2556 0 1
rlabel polysilicon 667 -2562 667 -2562 0 3
rlabel polysilicon 674 -2556 674 -2556 0 1
rlabel polysilicon 674 -2562 674 -2562 0 3
rlabel polysilicon 681 -2556 681 -2556 0 1
rlabel polysilicon 681 -2562 681 -2562 0 3
rlabel polysilicon 688 -2556 688 -2556 0 1
rlabel polysilicon 688 -2562 688 -2562 0 3
rlabel polysilicon 695 -2556 695 -2556 0 1
rlabel polysilicon 695 -2562 695 -2562 0 3
rlabel polysilicon 702 -2556 702 -2556 0 1
rlabel polysilicon 702 -2562 702 -2562 0 3
rlabel polysilicon 709 -2556 709 -2556 0 1
rlabel polysilicon 709 -2562 709 -2562 0 3
rlabel polysilicon 716 -2556 716 -2556 0 1
rlabel polysilicon 716 -2562 716 -2562 0 3
rlabel polysilicon 723 -2556 723 -2556 0 1
rlabel polysilicon 723 -2562 723 -2562 0 3
rlabel polysilicon 730 -2556 730 -2556 0 1
rlabel polysilicon 733 -2556 733 -2556 0 2
rlabel polysilicon 730 -2562 730 -2562 0 3
rlabel polysilicon 733 -2562 733 -2562 0 4
rlabel polysilicon 737 -2556 737 -2556 0 1
rlabel polysilicon 740 -2556 740 -2556 0 2
rlabel polysilicon 737 -2562 737 -2562 0 3
rlabel polysilicon 740 -2562 740 -2562 0 4
rlabel polysilicon 744 -2556 744 -2556 0 1
rlabel polysilicon 747 -2556 747 -2556 0 2
rlabel polysilicon 747 -2562 747 -2562 0 4
rlabel polysilicon 751 -2556 751 -2556 0 1
rlabel polysilicon 754 -2556 754 -2556 0 2
rlabel polysilicon 751 -2562 751 -2562 0 3
rlabel polysilicon 754 -2562 754 -2562 0 4
rlabel polysilicon 758 -2556 758 -2556 0 1
rlabel polysilicon 758 -2562 758 -2562 0 3
rlabel polysilicon 765 -2556 765 -2556 0 1
rlabel polysilicon 765 -2562 765 -2562 0 3
rlabel polysilicon 772 -2556 772 -2556 0 1
rlabel polysilicon 772 -2562 772 -2562 0 3
rlabel polysilicon 779 -2556 779 -2556 0 1
rlabel polysilicon 779 -2562 779 -2562 0 3
rlabel polysilicon 786 -2556 786 -2556 0 1
rlabel polysilicon 789 -2556 789 -2556 0 2
rlabel polysilicon 786 -2562 786 -2562 0 3
rlabel polysilicon 789 -2562 789 -2562 0 4
rlabel polysilicon 793 -2556 793 -2556 0 1
rlabel polysilicon 793 -2562 793 -2562 0 3
rlabel polysilicon 800 -2556 800 -2556 0 1
rlabel polysilicon 800 -2562 800 -2562 0 3
rlabel polysilicon 807 -2556 807 -2556 0 1
rlabel polysilicon 807 -2562 807 -2562 0 3
rlabel polysilicon 814 -2556 814 -2556 0 1
rlabel polysilicon 814 -2562 814 -2562 0 3
rlabel polysilicon 821 -2556 821 -2556 0 1
rlabel polysilicon 824 -2556 824 -2556 0 2
rlabel polysilicon 821 -2562 821 -2562 0 3
rlabel polysilicon 824 -2562 824 -2562 0 4
rlabel polysilicon 828 -2556 828 -2556 0 1
rlabel polysilicon 828 -2562 828 -2562 0 3
rlabel polysilicon 835 -2556 835 -2556 0 1
rlabel polysilicon 835 -2562 835 -2562 0 3
rlabel polysilicon 842 -2556 842 -2556 0 1
rlabel polysilicon 842 -2562 842 -2562 0 3
rlabel polysilicon 849 -2556 849 -2556 0 1
rlabel polysilicon 849 -2562 849 -2562 0 3
rlabel polysilicon 856 -2556 856 -2556 0 1
rlabel polysilicon 856 -2562 856 -2562 0 3
rlabel polysilicon 863 -2556 863 -2556 0 1
rlabel polysilicon 863 -2562 863 -2562 0 3
rlabel polysilicon 870 -2556 870 -2556 0 1
rlabel polysilicon 873 -2556 873 -2556 0 2
rlabel polysilicon 870 -2562 870 -2562 0 3
rlabel polysilicon 873 -2562 873 -2562 0 4
rlabel polysilicon 877 -2556 877 -2556 0 1
rlabel polysilicon 877 -2562 877 -2562 0 3
rlabel polysilicon 884 -2556 884 -2556 0 1
rlabel polysilicon 884 -2562 884 -2562 0 3
rlabel polysilicon 891 -2556 891 -2556 0 1
rlabel polysilicon 891 -2562 891 -2562 0 3
rlabel polysilicon 898 -2556 898 -2556 0 1
rlabel polysilicon 898 -2562 898 -2562 0 3
rlabel polysilicon 905 -2556 905 -2556 0 1
rlabel polysilicon 905 -2562 905 -2562 0 3
rlabel polysilicon 912 -2556 912 -2556 0 1
rlabel polysilicon 912 -2562 912 -2562 0 3
rlabel polysilicon 919 -2556 919 -2556 0 1
rlabel polysilicon 919 -2562 919 -2562 0 3
rlabel polysilicon 926 -2556 926 -2556 0 1
rlabel polysilicon 929 -2556 929 -2556 0 2
rlabel polysilicon 926 -2562 926 -2562 0 3
rlabel polysilicon 929 -2562 929 -2562 0 4
rlabel polysilicon 933 -2556 933 -2556 0 1
rlabel polysilicon 933 -2562 933 -2562 0 3
rlabel polysilicon 940 -2556 940 -2556 0 1
rlabel polysilicon 940 -2562 940 -2562 0 3
rlabel polysilicon 947 -2556 947 -2556 0 1
rlabel polysilicon 947 -2562 947 -2562 0 3
rlabel polysilicon 954 -2556 954 -2556 0 1
rlabel polysilicon 957 -2556 957 -2556 0 2
rlabel polysilicon 954 -2562 954 -2562 0 3
rlabel polysilicon 957 -2562 957 -2562 0 4
rlabel polysilicon 961 -2556 961 -2556 0 1
rlabel polysilicon 961 -2562 961 -2562 0 3
rlabel polysilicon 968 -2556 968 -2556 0 1
rlabel polysilicon 968 -2562 968 -2562 0 3
rlabel polysilicon 975 -2556 975 -2556 0 1
rlabel polysilicon 975 -2562 975 -2562 0 3
rlabel polysilicon 982 -2556 982 -2556 0 1
rlabel polysilicon 982 -2562 982 -2562 0 3
rlabel polysilicon 989 -2556 989 -2556 0 1
rlabel polysilicon 989 -2562 989 -2562 0 3
rlabel polysilicon 996 -2556 996 -2556 0 1
rlabel polysilicon 996 -2562 996 -2562 0 3
rlabel polysilicon 1003 -2556 1003 -2556 0 1
rlabel polysilicon 1003 -2562 1003 -2562 0 3
rlabel polysilicon 1010 -2556 1010 -2556 0 1
rlabel polysilicon 1010 -2562 1010 -2562 0 3
rlabel polysilicon 1017 -2556 1017 -2556 0 1
rlabel polysilicon 1017 -2562 1017 -2562 0 3
rlabel polysilicon 1024 -2556 1024 -2556 0 1
rlabel polysilicon 1024 -2562 1024 -2562 0 3
rlabel polysilicon 1031 -2556 1031 -2556 0 1
rlabel polysilicon 1031 -2562 1031 -2562 0 3
rlabel polysilicon 1038 -2556 1038 -2556 0 1
rlabel polysilicon 1038 -2562 1038 -2562 0 3
rlabel polysilicon 1045 -2556 1045 -2556 0 1
rlabel polysilicon 1045 -2562 1045 -2562 0 3
rlabel polysilicon 1052 -2556 1052 -2556 0 1
rlabel polysilicon 1052 -2562 1052 -2562 0 3
rlabel polysilicon 1059 -2556 1059 -2556 0 1
rlabel polysilicon 1062 -2556 1062 -2556 0 2
rlabel polysilicon 1059 -2562 1059 -2562 0 3
rlabel polysilicon 1062 -2562 1062 -2562 0 4
rlabel polysilicon 1066 -2556 1066 -2556 0 1
rlabel polysilicon 1066 -2562 1066 -2562 0 3
rlabel polysilicon 1073 -2556 1073 -2556 0 1
rlabel polysilicon 1073 -2562 1073 -2562 0 3
rlabel polysilicon 1080 -2556 1080 -2556 0 1
rlabel polysilicon 1083 -2556 1083 -2556 0 2
rlabel polysilicon 1083 -2562 1083 -2562 0 4
rlabel polysilicon 1087 -2556 1087 -2556 0 1
rlabel polysilicon 1090 -2556 1090 -2556 0 2
rlabel polysilicon 1090 -2562 1090 -2562 0 4
rlabel polysilicon 1094 -2556 1094 -2556 0 1
rlabel polysilicon 1094 -2562 1094 -2562 0 3
rlabel polysilicon 1101 -2556 1101 -2556 0 1
rlabel polysilicon 1101 -2562 1101 -2562 0 3
rlabel polysilicon 1108 -2556 1108 -2556 0 1
rlabel polysilicon 1108 -2562 1108 -2562 0 3
rlabel polysilicon 1115 -2556 1115 -2556 0 1
rlabel polysilicon 1115 -2562 1115 -2562 0 3
rlabel polysilicon 1122 -2556 1122 -2556 0 1
rlabel polysilicon 1122 -2562 1122 -2562 0 3
rlabel polysilicon 1129 -2556 1129 -2556 0 1
rlabel polysilicon 1129 -2562 1129 -2562 0 3
rlabel polysilicon 1136 -2556 1136 -2556 0 1
rlabel polysilicon 1136 -2562 1136 -2562 0 3
rlabel polysilicon 1143 -2556 1143 -2556 0 1
rlabel polysilicon 1143 -2562 1143 -2562 0 3
rlabel polysilicon 1150 -2556 1150 -2556 0 1
rlabel polysilicon 1150 -2562 1150 -2562 0 3
rlabel polysilicon 1157 -2556 1157 -2556 0 1
rlabel polysilicon 1157 -2562 1157 -2562 0 3
rlabel polysilicon 1164 -2556 1164 -2556 0 1
rlabel polysilicon 1167 -2556 1167 -2556 0 2
rlabel polysilicon 1164 -2562 1164 -2562 0 3
rlabel polysilicon 1167 -2562 1167 -2562 0 4
rlabel polysilicon 1171 -2556 1171 -2556 0 1
rlabel polysilicon 1171 -2562 1171 -2562 0 3
rlabel polysilicon 1178 -2556 1178 -2556 0 1
rlabel polysilicon 1178 -2562 1178 -2562 0 3
rlabel polysilicon 1185 -2556 1185 -2556 0 1
rlabel polysilicon 1188 -2556 1188 -2556 0 2
rlabel polysilicon 1185 -2562 1185 -2562 0 3
rlabel polysilicon 1192 -2556 1192 -2556 0 1
rlabel polysilicon 1192 -2562 1192 -2562 0 3
rlabel polysilicon 1199 -2556 1199 -2556 0 1
rlabel polysilicon 1199 -2562 1199 -2562 0 3
rlabel polysilicon 1206 -2556 1206 -2556 0 1
rlabel polysilicon 1206 -2562 1206 -2562 0 3
rlabel polysilicon 1213 -2556 1213 -2556 0 1
rlabel polysilicon 1213 -2562 1213 -2562 0 3
rlabel polysilicon 1220 -2556 1220 -2556 0 1
rlabel polysilicon 1220 -2562 1220 -2562 0 3
rlabel polysilicon 1227 -2556 1227 -2556 0 1
rlabel polysilicon 1227 -2562 1227 -2562 0 3
rlabel polysilicon 1234 -2556 1234 -2556 0 1
rlabel polysilicon 1234 -2562 1234 -2562 0 3
rlabel polysilicon 1241 -2556 1241 -2556 0 1
rlabel polysilicon 1241 -2562 1241 -2562 0 3
rlabel polysilicon 1248 -2556 1248 -2556 0 1
rlabel polysilicon 1248 -2562 1248 -2562 0 3
rlabel polysilicon 1255 -2556 1255 -2556 0 1
rlabel polysilicon 1255 -2562 1255 -2562 0 3
rlabel polysilicon 1262 -2556 1262 -2556 0 1
rlabel polysilicon 1262 -2562 1262 -2562 0 3
rlabel polysilicon 1269 -2556 1269 -2556 0 1
rlabel polysilicon 1269 -2562 1269 -2562 0 3
rlabel polysilicon 1276 -2556 1276 -2556 0 1
rlabel polysilicon 1276 -2562 1276 -2562 0 3
rlabel polysilicon 1283 -2556 1283 -2556 0 1
rlabel polysilicon 1283 -2562 1283 -2562 0 3
rlabel polysilicon 1290 -2556 1290 -2556 0 1
rlabel polysilicon 1290 -2562 1290 -2562 0 3
rlabel polysilicon 1297 -2556 1297 -2556 0 1
rlabel polysilicon 1297 -2562 1297 -2562 0 3
rlabel polysilicon 1304 -2556 1304 -2556 0 1
rlabel polysilicon 1304 -2562 1304 -2562 0 3
rlabel polysilicon 1311 -2556 1311 -2556 0 1
rlabel polysilicon 1311 -2562 1311 -2562 0 3
rlabel polysilicon 1318 -2556 1318 -2556 0 1
rlabel polysilicon 1318 -2562 1318 -2562 0 3
rlabel polysilicon 1325 -2556 1325 -2556 0 1
rlabel polysilicon 1325 -2562 1325 -2562 0 3
rlabel polysilicon 1332 -2556 1332 -2556 0 1
rlabel polysilicon 1332 -2562 1332 -2562 0 3
rlabel polysilicon 1339 -2556 1339 -2556 0 1
rlabel polysilicon 1339 -2562 1339 -2562 0 3
rlabel polysilicon 1346 -2556 1346 -2556 0 1
rlabel polysilicon 1346 -2562 1346 -2562 0 3
rlabel polysilicon 1353 -2556 1353 -2556 0 1
rlabel polysilicon 1353 -2562 1353 -2562 0 3
rlabel polysilicon 1360 -2556 1360 -2556 0 1
rlabel polysilicon 1360 -2562 1360 -2562 0 3
rlabel polysilicon 1367 -2556 1367 -2556 0 1
rlabel polysilicon 1367 -2562 1367 -2562 0 3
rlabel polysilicon 1374 -2556 1374 -2556 0 1
rlabel polysilicon 1374 -2562 1374 -2562 0 3
rlabel polysilicon 1381 -2556 1381 -2556 0 1
rlabel polysilicon 1381 -2562 1381 -2562 0 3
rlabel polysilicon 1388 -2556 1388 -2556 0 1
rlabel polysilicon 1388 -2562 1388 -2562 0 3
rlabel polysilicon 1395 -2556 1395 -2556 0 1
rlabel polysilicon 1395 -2562 1395 -2562 0 3
rlabel polysilicon 1402 -2556 1402 -2556 0 1
rlabel polysilicon 1402 -2562 1402 -2562 0 3
rlabel polysilicon 1409 -2556 1409 -2556 0 1
rlabel polysilicon 1409 -2562 1409 -2562 0 3
rlabel polysilicon 1416 -2556 1416 -2556 0 1
rlabel polysilicon 1416 -2562 1416 -2562 0 3
rlabel polysilicon 1423 -2556 1423 -2556 0 1
rlabel polysilicon 1423 -2562 1423 -2562 0 3
rlabel polysilicon 1430 -2556 1430 -2556 0 1
rlabel polysilicon 1430 -2562 1430 -2562 0 3
rlabel polysilicon 1437 -2556 1437 -2556 0 1
rlabel polysilicon 1437 -2562 1437 -2562 0 3
rlabel polysilicon 1444 -2556 1444 -2556 0 1
rlabel polysilicon 1444 -2562 1444 -2562 0 3
rlabel polysilicon 1451 -2556 1451 -2556 0 1
rlabel polysilicon 1451 -2562 1451 -2562 0 3
rlabel polysilicon 1458 -2556 1458 -2556 0 1
rlabel polysilicon 1458 -2562 1458 -2562 0 3
rlabel polysilicon 1465 -2556 1465 -2556 0 1
rlabel polysilicon 1465 -2562 1465 -2562 0 3
rlabel polysilicon 1472 -2556 1472 -2556 0 1
rlabel polysilicon 1472 -2562 1472 -2562 0 3
rlabel polysilicon 1479 -2556 1479 -2556 0 1
rlabel polysilicon 1479 -2562 1479 -2562 0 3
rlabel polysilicon 1486 -2556 1486 -2556 0 1
rlabel polysilicon 1486 -2562 1486 -2562 0 3
rlabel polysilicon 1493 -2556 1493 -2556 0 1
rlabel polysilicon 1493 -2562 1493 -2562 0 3
rlabel polysilicon 1500 -2556 1500 -2556 0 1
rlabel polysilicon 1500 -2562 1500 -2562 0 3
rlabel polysilicon 1507 -2556 1507 -2556 0 1
rlabel polysilicon 1507 -2562 1507 -2562 0 3
rlabel polysilicon 1514 -2556 1514 -2556 0 1
rlabel polysilicon 1514 -2562 1514 -2562 0 3
rlabel polysilicon 1521 -2556 1521 -2556 0 1
rlabel polysilicon 1521 -2562 1521 -2562 0 3
rlabel polysilicon 1528 -2556 1528 -2556 0 1
rlabel polysilicon 1528 -2562 1528 -2562 0 3
rlabel polysilicon 1535 -2556 1535 -2556 0 1
rlabel polysilicon 1535 -2562 1535 -2562 0 3
rlabel polysilicon 1542 -2556 1542 -2556 0 1
rlabel polysilicon 1542 -2562 1542 -2562 0 3
rlabel polysilicon 1549 -2556 1549 -2556 0 1
rlabel polysilicon 1549 -2562 1549 -2562 0 3
rlabel polysilicon 1556 -2556 1556 -2556 0 1
rlabel polysilicon 1556 -2562 1556 -2562 0 3
rlabel polysilicon 1563 -2556 1563 -2556 0 1
rlabel polysilicon 1563 -2562 1563 -2562 0 3
rlabel polysilicon 1570 -2556 1570 -2556 0 1
rlabel polysilicon 1570 -2562 1570 -2562 0 3
rlabel polysilicon 1577 -2556 1577 -2556 0 1
rlabel polysilicon 1577 -2562 1577 -2562 0 3
rlabel polysilicon 1584 -2556 1584 -2556 0 1
rlabel polysilicon 1584 -2562 1584 -2562 0 3
rlabel polysilicon 1591 -2556 1591 -2556 0 1
rlabel polysilicon 1591 -2562 1591 -2562 0 3
rlabel polysilicon 1598 -2556 1598 -2556 0 1
rlabel polysilicon 1598 -2562 1598 -2562 0 3
rlabel polysilicon 1605 -2556 1605 -2556 0 1
rlabel polysilicon 1605 -2562 1605 -2562 0 3
rlabel polysilicon 1612 -2556 1612 -2556 0 1
rlabel polysilicon 1612 -2562 1612 -2562 0 3
rlabel polysilicon 1619 -2556 1619 -2556 0 1
rlabel polysilicon 1619 -2562 1619 -2562 0 3
rlabel polysilicon 1626 -2556 1626 -2556 0 1
rlabel polysilicon 1626 -2562 1626 -2562 0 3
rlabel polysilicon 1633 -2556 1633 -2556 0 1
rlabel polysilicon 1633 -2562 1633 -2562 0 3
rlabel polysilicon 1640 -2556 1640 -2556 0 1
rlabel polysilicon 1640 -2562 1640 -2562 0 3
rlabel polysilicon 1647 -2556 1647 -2556 0 1
rlabel polysilicon 1647 -2562 1647 -2562 0 3
rlabel polysilicon 1654 -2556 1654 -2556 0 1
rlabel polysilicon 1654 -2562 1654 -2562 0 3
rlabel polysilicon 1661 -2556 1661 -2556 0 1
rlabel polysilicon 1661 -2562 1661 -2562 0 3
rlabel polysilicon 1668 -2556 1668 -2556 0 1
rlabel polysilicon 1668 -2562 1668 -2562 0 3
rlabel polysilicon 1678 -2556 1678 -2556 0 2
rlabel polysilicon 1675 -2562 1675 -2562 0 3
rlabel polysilicon 1678 -2562 1678 -2562 0 4
rlabel polysilicon 1682 -2556 1682 -2556 0 1
rlabel polysilicon 1682 -2562 1682 -2562 0 3
rlabel polysilicon 1689 -2556 1689 -2556 0 1
rlabel polysilicon 1689 -2562 1689 -2562 0 3
rlabel polysilicon 1696 -2556 1696 -2556 0 1
rlabel polysilicon 1696 -2562 1696 -2562 0 3
rlabel polysilicon 1706 -2556 1706 -2556 0 2
rlabel polysilicon 1703 -2562 1703 -2562 0 3
rlabel polysilicon 1710 -2556 1710 -2556 0 1
rlabel polysilicon 1710 -2562 1710 -2562 0 3
rlabel polysilicon 1717 -2556 1717 -2556 0 1
rlabel polysilicon 1717 -2562 1717 -2562 0 3
rlabel polysilicon 1724 -2556 1724 -2556 0 1
rlabel polysilicon 1724 -2562 1724 -2562 0 3
rlabel polysilicon 1731 -2556 1731 -2556 0 1
rlabel polysilicon 1731 -2562 1731 -2562 0 3
rlabel polysilicon 1738 -2556 1738 -2556 0 1
rlabel polysilicon 1738 -2562 1738 -2562 0 3
rlabel polysilicon 44 -2685 44 -2685 0 1
rlabel polysilicon 44 -2691 44 -2691 0 3
rlabel polysilicon 51 -2685 51 -2685 0 1
rlabel polysilicon 51 -2691 51 -2691 0 3
rlabel polysilicon 58 -2685 58 -2685 0 1
rlabel polysilicon 58 -2691 58 -2691 0 3
rlabel polysilicon 65 -2685 65 -2685 0 1
rlabel polysilicon 68 -2685 68 -2685 0 2
rlabel polysilicon 65 -2691 65 -2691 0 3
rlabel polysilicon 68 -2691 68 -2691 0 4
rlabel polysilicon 72 -2685 72 -2685 0 1
rlabel polysilicon 72 -2691 72 -2691 0 3
rlabel polysilicon 82 -2685 82 -2685 0 2
rlabel polysilicon 79 -2691 79 -2691 0 3
rlabel polysilicon 82 -2691 82 -2691 0 4
rlabel polysilicon 86 -2685 86 -2685 0 1
rlabel polysilicon 89 -2685 89 -2685 0 2
rlabel polysilicon 86 -2691 86 -2691 0 3
rlabel polysilicon 89 -2691 89 -2691 0 4
rlabel polysilicon 93 -2685 93 -2685 0 1
rlabel polysilicon 93 -2691 93 -2691 0 3
rlabel polysilicon 100 -2685 100 -2685 0 1
rlabel polysilicon 100 -2691 100 -2691 0 3
rlabel polysilicon 107 -2685 107 -2685 0 1
rlabel polysilicon 107 -2691 107 -2691 0 3
rlabel polysilicon 117 -2685 117 -2685 0 2
rlabel polysilicon 114 -2691 114 -2691 0 3
rlabel polysilicon 117 -2691 117 -2691 0 4
rlabel polysilicon 121 -2685 121 -2685 0 1
rlabel polysilicon 121 -2691 121 -2691 0 3
rlabel polysilicon 128 -2685 128 -2685 0 1
rlabel polysilicon 128 -2691 128 -2691 0 3
rlabel polysilicon 135 -2685 135 -2685 0 1
rlabel polysilicon 135 -2691 135 -2691 0 3
rlabel polysilicon 142 -2685 142 -2685 0 1
rlabel polysilicon 142 -2691 142 -2691 0 3
rlabel polysilicon 149 -2685 149 -2685 0 1
rlabel polysilicon 149 -2691 149 -2691 0 3
rlabel polysilicon 156 -2685 156 -2685 0 1
rlabel polysilicon 156 -2691 156 -2691 0 3
rlabel polysilicon 163 -2685 163 -2685 0 1
rlabel polysilicon 166 -2685 166 -2685 0 2
rlabel polysilicon 163 -2691 163 -2691 0 3
rlabel polysilicon 166 -2691 166 -2691 0 4
rlabel polysilicon 170 -2685 170 -2685 0 1
rlabel polysilicon 170 -2691 170 -2691 0 3
rlabel polysilicon 177 -2685 177 -2685 0 1
rlabel polysilicon 177 -2691 177 -2691 0 3
rlabel polysilicon 184 -2685 184 -2685 0 1
rlabel polysilicon 184 -2691 184 -2691 0 3
rlabel polysilicon 191 -2685 191 -2685 0 1
rlabel polysilicon 201 -2685 201 -2685 0 2
rlabel polysilicon 198 -2691 198 -2691 0 3
rlabel polysilicon 201 -2691 201 -2691 0 4
rlabel polysilicon 205 -2685 205 -2685 0 1
rlabel polysilicon 205 -2691 205 -2691 0 3
rlabel polysilicon 212 -2685 212 -2685 0 1
rlabel polysilicon 212 -2691 212 -2691 0 3
rlabel polysilicon 219 -2685 219 -2685 0 1
rlabel polysilicon 219 -2691 219 -2691 0 3
rlabel polysilicon 226 -2685 226 -2685 0 1
rlabel polysilicon 226 -2691 226 -2691 0 3
rlabel polysilicon 233 -2685 233 -2685 0 1
rlabel polysilicon 233 -2691 233 -2691 0 3
rlabel polysilicon 240 -2685 240 -2685 0 1
rlabel polysilicon 240 -2691 240 -2691 0 3
rlabel polysilicon 247 -2691 247 -2691 0 3
rlabel polysilicon 250 -2691 250 -2691 0 4
rlabel polysilicon 254 -2685 254 -2685 0 1
rlabel polysilicon 254 -2691 254 -2691 0 3
rlabel polysilicon 261 -2685 261 -2685 0 1
rlabel polysilicon 261 -2691 261 -2691 0 3
rlabel polysilicon 268 -2685 268 -2685 0 1
rlabel polysilicon 268 -2691 268 -2691 0 3
rlabel polysilicon 275 -2685 275 -2685 0 1
rlabel polysilicon 275 -2691 275 -2691 0 3
rlabel polysilicon 278 -2691 278 -2691 0 4
rlabel polysilicon 282 -2685 282 -2685 0 1
rlabel polysilicon 282 -2691 282 -2691 0 3
rlabel polysilicon 289 -2685 289 -2685 0 1
rlabel polysilicon 289 -2691 289 -2691 0 3
rlabel polysilicon 296 -2685 296 -2685 0 1
rlabel polysilicon 296 -2691 296 -2691 0 3
rlabel polysilicon 303 -2685 303 -2685 0 1
rlabel polysilicon 303 -2691 303 -2691 0 3
rlabel polysilicon 310 -2685 310 -2685 0 1
rlabel polysilicon 310 -2691 310 -2691 0 3
rlabel polysilicon 317 -2685 317 -2685 0 1
rlabel polysilicon 317 -2691 317 -2691 0 3
rlabel polysilicon 324 -2685 324 -2685 0 1
rlabel polysilicon 324 -2691 324 -2691 0 3
rlabel polysilicon 331 -2685 331 -2685 0 1
rlabel polysilicon 331 -2691 331 -2691 0 3
rlabel polysilicon 338 -2685 338 -2685 0 1
rlabel polysilicon 338 -2691 338 -2691 0 3
rlabel polysilicon 345 -2685 345 -2685 0 1
rlabel polysilicon 345 -2691 345 -2691 0 3
rlabel polysilicon 352 -2685 352 -2685 0 1
rlabel polysilicon 352 -2691 352 -2691 0 3
rlabel polysilicon 359 -2685 359 -2685 0 1
rlabel polysilicon 359 -2691 359 -2691 0 3
rlabel polysilicon 366 -2685 366 -2685 0 1
rlabel polysilicon 366 -2691 366 -2691 0 3
rlabel polysilicon 373 -2685 373 -2685 0 1
rlabel polysilicon 373 -2691 373 -2691 0 3
rlabel polysilicon 380 -2685 380 -2685 0 1
rlabel polysilicon 380 -2691 380 -2691 0 3
rlabel polysilicon 387 -2685 387 -2685 0 1
rlabel polysilicon 387 -2691 387 -2691 0 3
rlabel polysilicon 394 -2685 394 -2685 0 1
rlabel polysilicon 394 -2691 394 -2691 0 3
rlabel polysilicon 401 -2685 401 -2685 0 1
rlabel polysilicon 401 -2691 401 -2691 0 3
rlabel polysilicon 408 -2685 408 -2685 0 1
rlabel polysilicon 411 -2685 411 -2685 0 2
rlabel polysilicon 411 -2691 411 -2691 0 4
rlabel polysilicon 418 -2685 418 -2685 0 2
rlabel polysilicon 415 -2691 415 -2691 0 3
rlabel polysilicon 418 -2691 418 -2691 0 4
rlabel polysilicon 422 -2685 422 -2685 0 1
rlabel polysilicon 422 -2691 422 -2691 0 3
rlabel polysilicon 429 -2685 429 -2685 0 1
rlabel polysilicon 429 -2691 429 -2691 0 3
rlabel polysilicon 436 -2685 436 -2685 0 1
rlabel polysilicon 436 -2691 436 -2691 0 3
rlabel polysilicon 443 -2685 443 -2685 0 1
rlabel polysilicon 443 -2691 443 -2691 0 3
rlabel polysilicon 450 -2685 450 -2685 0 1
rlabel polysilicon 450 -2691 450 -2691 0 3
rlabel polysilicon 453 -2691 453 -2691 0 4
rlabel polysilicon 457 -2685 457 -2685 0 1
rlabel polysilicon 460 -2685 460 -2685 0 2
rlabel polysilicon 457 -2691 457 -2691 0 3
rlabel polysilicon 464 -2685 464 -2685 0 1
rlabel polysilicon 464 -2691 464 -2691 0 3
rlabel polysilicon 467 -2691 467 -2691 0 4
rlabel polysilicon 471 -2685 471 -2685 0 1
rlabel polysilicon 471 -2691 471 -2691 0 3
rlabel polysilicon 478 -2685 478 -2685 0 1
rlabel polysilicon 481 -2691 481 -2691 0 4
rlabel polysilicon 485 -2685 485 -2685 0 1
rlabel polysilicon 485 -2691 485 -2691 0 3
rlabel polysilicon 492 -2685 492 -2685 0 1
rlabel polysilicon 492 -2691 492 -2691 0 3
rlabel polysilicon 499 -2685 499 -2685 0 1
rlabel polysilicon 499 -2691 499 -2691 0 3
rlabel polysilicon 506 -2685 506 -2685 0 1
rlabel polysilicon 506 -2691 506 -2691 0 3
rlabel polysilicon 513 -2685 513 -2685 0 1
rlabel polysilicon 513 -2691 513 -2691 0 3
rlabel polysilicon 520 -2685 520 -2685 0 1
rlabel polysilicon 520 -2691 520 -2691 0 3
rlabel polysilicon 527 -2685 527 -2685 0 1
rlabel polysilicon 527 -2691 527 -2691 0 3
rlabel polysilicon 534 -2685 534 -2685 0 1
rlabel polysilicon 534 -2691 534 -2691 0 3
rlabel polysilicon 541 -2685 541 -2685 0 1
rlabel polysilicon 541 -2691 541 -2691 0 3
rlabel polysilicon 548 -2685 548 -2685 0 1
rlabel polysilicon 548 -2691 548 -2691 0 3
rlabel polysilicon 555 -2685 555 -2685 0 1
rlabel polysilicon 555 -2691 555 -2691 0 3
rlabel polysilicon 562 -2685 562 -2685 0 1
rlabel polysilicon 562 -2691 562 -2691 0 3
rlabel polysilicon 569 -2685 569 -2685 0 1
rlabel polysilicon 569 -2691 569 -2691 0 3
rlabel polysilicon 576 -2685 576 -2685 0 1
rlabel polysilicon 579 -2691 579 -2691 0 4
rlabel polysilicon 583 -2685 583 -2685 0 1
rlabel polysilicon 583 -2691 583 -2691 0 3
rlabel polysilicon 590 -2685 590 -2685 0 1
rlabel polysilicon 590 -2691 590 -2691 0 3
rlabel polysilicon 597 -2685 597 -2685 0 1
rlabel polysilicon 600 -2685 600 -2685 0 2
rlabel polysilicon 597 -2691 597 -2691 0 3
rlabel polysilicon 600 -2691 600 -2691 0 4
rlabel polysilicon 604 -2685 604 -2685 0 1
rlabel polysilicon 604 -2691 604 -2691 0 3
rlabel polysilicon 611 -2685 611 -2685 0 1
rlabel polysilicon 611 -2691 611 -2691 0 3
rlabel polysilicon 618 -2685 618 -2685 0 1
rlabel polysilicon 618 -2691 618 -2691 0 3
rlabel polysilicon 625 -2685 625 -2685 0 1
rlabel polysilicon 628 -2685 628 -2685 0 2
rlabel polysilicon 625 -2691 625 -2691 0 3
rlabel polysilicon 628 -2691 628 -2691 0 4
rlabel polysilicon 632 -2685 632 -2685 0 1
rlabel polysilicon 632 -2691 632 -2691 0 3
rlabel polysilicon 639 -2685 639 -2685 0 1
rlabel polysilicon 639 -2691 639 -2691 0 3
rlabel polysilicon 646 -2685 646 -2685 0 1
rlabel polysilicon 646 -2691 646 -2691 0 3
rlabel polysilicon 653 -2685 653 -2685 0 1
rlabel polysilicon 653 -2691 653 -2691 0 3
rlabel polysilicon 660 -2685 660 -2685 0 1
rlabel polysilicon 660 -2691 660 -2691 0 3
rlabel polysilicon 667 -2685 667 -2685 0 1
rlabel polysilicon 670 -2685 670 -2685 0 2
rlabel polysilicon 667 -2691 667 -2691 0 3
rlabel polysilicon 670 -2691 670 -2691 0 4
rlabel polysilicon 674 -2685 674 -2685 0 1
rlabel polysilicon 677 -2685 677 -2685 0 2
rlabel polysilicon 674 -2691 674 -2691 0 3
rlabel polysilicon 677 -2691 677 -2691 0 4
rlabel polysilicon 681 -2685 681 -2685 0 1
rlabel polysilicon 681 -2691 681 -2691 0 3
rlabel polysilicon 688 -2685 688 -2685 0 1
rlabel polysilicon 691 -2685 691 -2685 0 2
rlabel polysilicon 688 -2691 688 -2691 0 3
rlabel polysilicon 695 -2685 695 -2685 0 1
rlabel polysilicon 695 -2691 695 -2691 0 3
rlabel polysilicon 702 -2685 702 -2685 0 1
rlabel polysilicon 702 -2691 702 -2691 0 3
rlabel polysilicon 709 -2685 709 -2685 0 1
rlabel polysilicon 709 -2691 709 -2691 0 3
rlabel polysilicon 716 -2685 716 -2685 0 1
rlabel polysilicon 716 -2691 716 -2691 0 3
rlabel polysilicon 723 -2685 723 -2685 0 1
rlabel polysilicon 723 -2691 723 -2691 0 3
rlabel polysilicon 733 -2685 733 -2685 0 2
rlabel polysilicon 730 -2691 730 -2691 0 3
rlabel polysilicon 733 -2691 733 -2691 0 4
rlabel polysilicon 737 -2685 737 -2685 0 1
rlabel polysilicon 737 -2691 737 -2691 0 3
rlabel polysilicon 744 -2685 744 -2685 0 1
rlabel polysilicon 744 -2691 744 -2691 0 3
rlabel polysilicon 751 -2685 751 -2685 0 1
rlabel polysilicon 751 -2691 751 -2691 0 3
rlabel polysilicon 754 -2691 754 -2691 0 4
rlabel polysilicon 758 -2685 758 -2685 0 1
rlabel polysilicon 758 -2691 758 -2691 0 3
rlabel polysilicon 765 -2685 765 -2685 0 1
rlabel polysilicon 768 -2685 768 -2685 0 2
rlabel polysilicon 765 -2691 765 -2691 0 3
rlabel polysilicon 768 -2691 768 -2691 0 4
rlabel polysilicon 772 -2685 772 -2685 0 1
rlabel polysilicon 772 -2691 772 -2691 0 3
rlabel polysilicon 779 -2685 779 -2685 0 1
rlabel polysilicon 779 -2691 779 -2691 0 3
rlabel polysilicon 786 -2685 786 -2685 0 1
rlabel polysilicon 786 -2691 786 -2691 0 3
rlabel polysilicon 793 -2685 793 -2685 0 1
rlabel polysilicon 793 -2691 793 -2691 0 3
rlabel polysilicon 800 -2685 800 -2685 0 1
rlabel polysilicon 803 -2685 803 -2685 0 2
rlabel polysilicon 800 -2691 800 -2691 0 3
rlabel polysilicon 803 -2691 803 -2691 0 4
rlabel polysilicon 807 -2685 807 -2685 0 1
rlabel polysilicon 807 -2691 807 -2691 0 3
rlabel polysilicon 814 -2685 814 -2685 0 1
rlabel polysilicon 814 -2691 814 -2691 0 3
rlabel polysilicon 821 -2685 821 -2685 0 1
rlabel polysilicon 821 -2691 821 -2691 0 3
rlabel polysilicon 828 -2685 828 -2685 0 1
rlabel polysilicon 828 -2691 828 -2691 0 3
rlabel polysilicon 838 -2685 838 -2685 0 2
rlabel polysilicon 835 -2691 835 -2691 0 3
rlabel polysilicon 838 -2691 838 -2691 0 4
rlabel polysilicon 842 -2685 842 -2685 0 1
rlabel polysilicon 845 -2685 845 -2685 0 2
rlabel polysilicon 842 -2691 842 -2691 0 3
rlabel polysilicon 845 -2691 845 -2691 0 4
rlabel polysilicon 849 -2685 849 -2685 0 1
rlabel polysilicon 849 -2691 849 -2691 0 3
rlabel polysilicon 856 -2685 856 -2685 0 1
rlabel polysilicon 856 -2691 856 -2691 0 3
rlabel polysilicon 863 -2685 863 -2685 0 1
rlabel polysilicon 863 -2691 863 -2691 0 3
rlabel polysilicon 870 -2685 870 -2685 0 1
rlabel polysilicon 873 -2685 873 -2685 0 2
rlabel polysilicon 870 -2691 870 -2691 0 3
rlabel polysilicon 873 -2691 873 -2691 0 4
rlabel polysilicon 877 -2685 877 -2685 0 1
rlabel polysilicon 877 -2691 877 -2691 0 3
rlabel polysilicon 884 -2685 884 -2685 0 1
rlabel polysilicon 884 -2691 884 -2691 0 3
rlabel polysilicon 891 -2685 891 -2685 0 1
rlabel polysilicon 894 -2685 894 -2685 0 2
rlabel polysilicon 894 -2691 894 -2691 0 4
rlabel polysilicon 898 -2685 898 -2685 0 1
rlabel polysilicon 898 -2691 898 -2691 0 3
rlabel polysilicon 905 -2685 905 -2685 0 1
rlabel polysilicon 905 -2691 905 -2691 0 3
rlabel polysilicon 912 -2685 912 -2685 0 1
rlabel polysilicon 912 -2691 912 -2691 0 3
rlabel polysilicon 919 -2685 919 -2685 0 1
rlabel polysilicon 919 -2691 919 -2691 0 3
rlabel polysilicon 926 -2685 926 -2685 0 1
rlabel polysilicon 926 -2691 926 -2691 0 3
rlabel polysilicon 933 -2685 933 -2685 0 1
rlabel polysilicon 933 -2691 933 -2691 0 3
rlabel polysilicon 940 -2685 940 -2685 0 1
rlabel polysilicon 940 -2691 940 -2691 0 3
rlabel polysilicon 947 -2685 947 -2685 0 1
rlabel polysilicon 947 -2691 947 -2691 0 3
rlabel polysilicon 954 -2685 954 -2685 0 1
rlabel polysilicon 957 -2685 957 -2685 0 2
rlabel polysilicon 954 -2691 954 -2691 0 3
rlabel polysilicon 957 -2691 957 -2691 0 4
rlabel polysilicon 961 -2685 961 -2685 0 1
rlabel polysilicon 961 -2691 961 -2691 0 3
rlabel polysilicon 968 -2685 968 -2685 0 1
rlabel polysilicon 968 -2691 968 -2691 0 3
rlabel polysilicon 975 -2685 975 -2685 0 1
rlabel polysilicon 975 -2691 975 -2691 0 3
rlabel polysilicon 982 -2685 982 -2685 0 1
rlabel polysilicon 982 -2691 982 -2691 0 3
rlabel polysilicon 989 -2685 989 -2685 0 1
rlabel polysilicon 989 -2691 989 -2691 0 3
rlabel polysilicon 996 -2685 996 -2685 0 1
rlabel polysilicon 996 -2691 996 -2691 0 3
rlabel polysilicon 1003 -2685 1003 -2685 0 1
rlabel polysilicon 1003 -2691 1003 -2691 0 3
rlabel polysilicon 1010 -2685 1010 -2685 0 1
rlabel polysilicon 1010 -2691 1010 -2691 0 3
rlabel polysilicon 1017 -2685 1017 -2685 0 1
rlabel polysilicon 1017 -2691 1017 -2691 0 3
rlabel polysilicon 1024 -2685 1024 -2685 0 1
rlabel polysilicon 1024 -2691 1024 -2691 0 3
rlabel polysilicon 1031 -2685 1031 -2685 0 1
rlabel polysilicon 1034 -2685 1034 -2685 0 2
rlabel polysilicon 1031 -2691 1031 -2691 0 3
rlabel polysilicon 1034 -2691 1034 -2691 0 4
rlabel polysilicon 1038 -2685 1038 -2685 0 1
rlabel polysilicon 1038 -2691 1038 -2691 0 3
rlabel polysilicon 1045 -2685 1045 -2685 0 1
rlabel polysilicon 1045 -2691 1045 -2691 0 3
rlabel polysilicon 1052 -2685 1052 -2685 0 1
rlabel polysilicon 1052 -2691 1052 -2691 0 3
rlabel polysilicon 1059 -2685 1059 -2685 0 1
rlabel polysilicon 1059 -2691 1059 -2691 0 3
rlabel polysilicon 1066 -2685 1066 -2685 0 1
rlabel polysilicon 1066 -2691 1066 -2691 0 3
rlabel polysilicon 1073 -2685 1073 -2685 0 1
rlabel polysilicon 1073 -2691 1073 -2691 0 3
rlabel polysilicon 1080 -2685 1080 -2685 0 1
rlabel polysilicon 1080 -2691 1080 -2691 0 3
rlabel polysilicon 1087 -2685 1087 -2685 0 1
rlabel polysilicon 1087 -2691 1087 -2691 0 3
rlabel polysilicon 1094 -2685 1094 -2685 0 1
rlabel polysilicon 1097 -2685 1097 -2685 0 2
rlabel polysilicon 1094 -2691 1094 -2691 0 3
rlabel polysilicon 1101 -2685 1101 -2685 0 1
rlabel polysilicon 1101 -2691 1101 -2691 0 3
rlabel polysilicon 1108 -2685 1108 -2685 0 1
rlabel polysilicon 1108 -2691 1108 -2691 0 3
rlabel polysilicon 1115 -2685 1115 -2685 0 1
rlabel polysilicon 1115 -2691 1115 -2691 0 3
rlabel polysilicon 1122 -2685 1122 -2685 0 1
rlabel polysilicon 1122 -2691 1122 -2691 0 3
rlabel polysilicon 1129 -2685 1129 -2685 0 1
rlabel polysilicon 1129 -2691 1129 -2691 0 3
rlabel polysilicon 1136 -2685 1136 -2685 0 1
rlabel polysilicon 1136 -2691 1136 -2691 0 3
rlabel polysilicon 1143 -2685 1143 -2685 0 1
rlabel polysilicon 1143 -2691 1143 -2691 0 3
rlabel polysilicon 1150 -2685 1150 -2685 0 1
rlabel polysilicon 1150 -2691 1150 -2691 0 3
rlabel polysilicon 1157 -2685 1157 -2685 0 1
rlabel polysilicon 1157 -2691 1157 -2691 0 3
rlabel polysilicon 1164 -2685 1164 -2685 0 1
rlabel polysilicon 1164 -2691 1164 -2691 0 3
rlabel polysilicon 1171 -2685 1171 -2685 0 1
rlabel polysilicon 1171 -2691 1171 -2691 0 3
rlabel polysilicon 1178 -2685 1178 -2685 0 1
rlabel polysilicon 1178 -2691 1178 -2691 0 3
rlabel polysilicon 1185 -2685 1185 -2685 0 1
rlabel polysilicon 1185 -2691 1185 -2691 0 3
rlabel polysilicon 1192 -2685 1192 -2685 0 1
rlabel polysilicon 1192 -2691 1192 -2691 0 3
rlabel polysilicon 1199 -2685 1199 -2685 0 1
rlabel polysilicon 1199 -2691 1199 -2691 0 3
rlabel polysilicon 1206 -2685 1206 -2685 0 1
rlabel polysilicon 1206 -2691 1206 -2691 0 3
rlabel polysilicon 1213 -2685 1213 -2685 0 1
rlabel polysilicon 1213 -2691 1213 -2691 0 3
rlabel polysilicon 1220 -2685 1220 -2685 0 1
rlabel polysilicon 1220 -2691 1220 -2691 0 3
rlabel polysilicon 1227 -2685 1227 -2685 0 1
rlabel polysilicon 1227 -2691 1227 -2691 0 3
rlabel polysilicon 1234 -2685 1234 -2685 0 1
rlabel polysilicon 1234 -2691 1234 -2691 0 3
rlabel polysilicon 1241 -2685 1241 -2685 0 1
rlabel polysilicon 1241 -2691 1241 -2691 0 3
rlabel polysilicon 1248 -2685 1248 -2685 0 1
rlabel polysilicon 1248 -2691 1248 -2691 0 3
rlabel polysilicon 1255 -2685 1255 -2685 0 1
rlabel polysilicon 1255 -2691 1255 -2691 0 3
rlabel polysilicon 1262 -2685 1262 -2685 0 1
rlabel polysilicon 1262 -2691 1262 -2691 0 3
rlabel polysilicon 1269 -2685 1269 -2685 0 1
rlabel polysilicon 1269 -2691 1269 -2691 0 3
rlabel polysilicon 1276 -2685 1276 -2685 0 1
rlabel polysilicon 1276 -2691 1276 -2691 0 3
rlabel polysilicon 1283 -2685 1283 -2685 0 1
rlabel polysilicon 1283 -2691 1283 -2691 0 3
rlabel polysilicon 1290 -2685 1290 -2685 0 1
rlabel polysilicon 1290 -2691 1290 -2691 0 3
rlabel polysilicon 1297 -2685 1297 -2685 0 1
rlabel polysilicon 1297 -2691 1297 -2691 0 3
rlabel polysilicon 1304 -2685 1304 -2685 0 1
rlabel polysilicon 1304 -2691 1304 -2691 0 3
rlabel polysilicon 1311 -2685 1311 -2685 0 1
rlabel polysilicon 1311 -2691 1311 -2691 0 3
rlabel polysilicon 1318 -2685 1318 -2685 0 1
rlabel polysilicon 1318 -2691 1318 -2691 0 3
rlabel polysilicon 1325 -2685 1325 -2685 0 1
rlabel polysilicon 1325 -2691 1325 -2691 0 3
rlabel polysilicon 1332 -2685 1332 -2685 0 1
rlabel polysilicon 1332 -2691 1332 -2691 0 3
rlabel polysilicon 1339 -2685 1339 -2685 0 1
rlabel polysilicon 1339 -2691 1339 -2691 0 3
rlabel polysilicon 1346 -2685 1346 -2685 0 1
rlabel polysilicon 1346 -2691 1346 -2691 0 3
rlabel polysilicon 1353 -2685 1353 -2685 0 1
rlabel polysilicon 1353 -2691 1353 -2691 0 3
rlabel polysilicon 1360 -2685 1360 -2685 0 1
rlabel polysilicon 1360 -2691 1360 -2691 0 3
rlabel polysilicon 1367 -2685 1367 -2685 0 1
rlabel polysilicon 1367 -2691 1367 -2691 0 3
rlabel polysilicon 1374 -2685 1374 -2685 0 1
rlabel polysilicon 1374 -2691 1374 -2691 0 3
rlabel polysilicon 1381 -2685 1381 -2685 0 1
rlabel polysilicon 1381 -2691 1381 -2691 0 3
rlabel polysilicon 1388 -2685 1388 -2685 0 1
rlabel polysilicon 1388 -2691 1388 -2691 0 3
rlabel polysilicon 1395 -2685 1395 -2685 0 1
rlabel polysilicon 1395 -2691 1395 -2691 0 3
rlabel polysilicon 1402 -2685 1402 -2685 0 1
rlabel polysilicon 1402 -2691 1402 -2691 0 3
rlabel polysilicon 1409 -2685 1409 -2685 0 1
rlabel polysilicon 1409 -2691 1409 -2691 0 3
rlabel polysilicon 1416 -2685 1416 -2685 0 1
rlabel polysilicon 1416 -2691 1416 -2691 0 3
rlabel polysilicon 1423 -2685 1423 -2685 0 1
rlabel polysilicon 1423 -2691 1423 -2691 0 3
rlabel polysilicon 1430 -2685 1430 -2685 0 1
rlabel polysilicon 1430 -2691 1430 -2691 0 3
rlabel polysilicon 1437 -2685 1437 -2685 0 1
rlabel polysilicon 1437 -2691 1437 -2691 0 3
rlabel polysilicon 1444 -2685 1444 -2685 0 1
rlabel polysilicon 1444 -2691 1444 -2691 0 3
rlabel polysilicon 1451 -2685 1451 -2685 0 1
rlabel polysilicon 1451 -2691 1451 -2691 0 3
rlabel polysilicon 1458 -2685 1458 -2685 0 1
rlabel polysilicon 1458 -2691 1458 -2691 0 3
rlabel polysilicon 1465 -2685 1465 -2685 0 1
rlabel polysilicon 1465 -2691 1465 -2691 0 3
rlabel polysilicon 1472 -2685 1472 -2685 0 1
rlabel polysilicon 1472 -2691 1472 -2691 0 3
rlabel polysilicon 1479 -2685 1479 -2685 0 1
rlabel polysilicon 1479 -2691 1479 -2691 0 3
rlabel polysilicon 1486 -2685 1486 -2685 0 1
rlabel polysilicon 1486 -2691 1486 -2691 0 3
rlabel polysilicon 1493 -2685 1493 -2685 0 1
rlabel polysilicon 1493 -2691 1493 -2691 0 3
rlabel polysilicon 1500 -2685 1500 -2685 0 1
rlabel polysilicon 1500 -2691 1500 -2691 0 3
rlabel polysilicon 1507 -2685 1507 -2685 0 1
rlabel polysilicon 1507 -2691 1507 -2691 0 3
rlabel polysilicon 1514 -2685 1514 -2685 0 1
rlabel polysilicon 1514 -2691 1514 -2691 0 3
rlabel polysilicon 1521 -2685 1521 -2685 0 1
rlabel polysilicon 1521 -2691 1521 -2691 0 3
rlabel polysilicon 1528 -2685 1528 -2685 0 1
rlabel polysilicon 1528 -2691 1528 -2691 0 3
rlabel polysilicon 1535 -2685 1535 -2685 0 1
rlabel polysilicon 1535 -2691 1535 -2691 0 3
rlabel polysilicon 1542 -2685 1542 -2685 0 1
rlabel polysilicon 1542 -2691 1542 -2691 0 3
rlabel polysilicon 1549 -2685 1549 -2685 0 1
rlabel polysilicon 1549 -2691 1549 -2691 0 3
rlabel polysilicon 1556 -2685 1556 -2685 0 1
rlabel polysilicon 1556 -2691 1556 -2691 0 3
rlabel polysilicon 1563 -2685 1563 -2685 0 1
rlabel polysilicon 1563 -2691 1563 -2691 0 3
rlabel polysilicon 1570 -2685 1570 -2685 0 1
rlabel polysilicon 1570 -2691 1570 -2691 0 3
rlabel polysilicon 1577 -2685 1577 -2685 0 1
rlabel polysilicon 1577 -2691 1577 -2691 0 3
rlabel polysilicon 1584 -2685 1584 -2685 0 1
rlabel polysilicon 1584 -2691 1584 -2691 0 3
rlabel polysilicon 1591 -2685 1591 -2685 0 1
rlabel polysilicon 1591 -2691 1591 -2691 0 3
rlabel polysilicon 1598 -2685 1598 -2685 0 1
rlabel polysilicon 1598 -2691 1598 -2691 0 3
rlabel polysilicon 1605 -2685 1605 -2685 0 1
rlabel polysilicon 1605 -2691 1605 -2691 0 3
rlabel polysilicon 1612 -2685 1612 -2685 0 1
rlabel polysilicon 1612 -2691 1612 -2691 0 3
rlabel polysilicon 1619 -2685 1619 -2685 0 1
rlabel polysilicon 1619 -2691 1619 -2691 0 3
rlabel polysilicon 1626 -2685 1626 -2685 0 1
rlabel polysilicon 1626 -2691 1626 -2691 0 3
rlabel polysilicon 1633 -2685 1633 -2685 0 1
rlabel polysilicon 1633 -2691 1633 -2691 0 3
rlabel polysilicon 1640 -2685 1640 -2685 0 1
rlabel polysilicon 1640 -2691 1640 -2691 0 3
rlabel polysilicon 1647 -2685 1647 -2685 0 1
rlabel polysilicon 1647 -2691 1647 -2691 0 3
rlabel polysilicon 1654 -2685 1654 -2685 0 1
rlabel polysilicon 1654 -2691 1654 -2691 0 3
rlabel polysilicon 1661 -2685 1661 -2685 0 1
rlabel polysilicon 1661 -2691 1661 -2691 0 3
rlabel polysilicon 1668 -2685 1668 -2685 0 1
rlabel polysilicon 1668 -2691 1668 -2691 0 3
rlabel polysilicon 1675 -2685 1675 -2685 0 1
rlabel polysilicon 1675 -2691 1675 -2691 0 3
rlabel polysilicon 1682 -2685 1682 -2685 0 1
rlabel polysilicon 1682 -2691 1682 -2691 0 3
rlabel polysilicon 1689 -2685 1689 -2685 0 1
rlabel polysilicon 1689 -2691 1689 -2691 0 3
rlabel polysilicon 1696 -2685 1696 -2685 0 1
rlabel polysilicon 1696 -2691 1696 -2691 0 3
rlabel polysilicon 1703 -2685 1703 -2685 0 1
rlabel polysilicon 1703 -2691 1703 -2691 0 3
rlabel polysilicon 37 -2834 37 -2834 0 1
rlabel polysilicon 37 -2840 37 -2840 0 3
rlabel polysilicon 44 -2834 44 -2834 0 1
rlabel polysilicon 44 -2840 44 -2840 0 3
rlabel polysilicon 51 -2834 51 -2834 0 1
rlabel polysilicon 51 -2840 51 -2840 0 3
rlabel polysilicon 58 -2834 58 -2834 0 1
rlabel polysilicon 58 -2840 58 -2840 0 3
rlabel polysilicon 65 -2834 65 -2834 0 1
rlabel polysilicon 65 -2840 65 -2840 0 3
rlabel polysilicon 72 -2834 72 -2834 0 1
rlabel polysilicon 72 -2840 72 -2840 0 3
rlabel polysilicon 79 -2834 79 -2834 0 1
rlabel polysilicon 79 -2840 79 -2840 0 3
rlabel polysilicon 86 -2834 86 -2834 0 1
rlabel polysilicon 89 -2834 89 -2834 0 2
rlabel polysilicon 93 -2834 93 -2834 0 1
rlabel polysilicon 96 -2834 96 -2834 0 2
rlabel polysilicon 93 -2840 93 -2840 0 3
rlabel polysilicon 96 -2840 96 -2840 0 4
rlabel polysilicon 100 -2834 100 -2834 0 1
rlabel polysilicon 100 -2840 100 -2840 0 3
rlabel polysilicon 107 -2834 107 -2834 0 1
rlabel polysilicon 110 -2834 110 -2834 0 2
rlabel polysilicon 107 -2840 107 -2840 0 3
rlabel polysilicon 110 -2840 110 -2840 0 4
rlabel polysilicon 114 -2834 114 -2834 0 1
rlabel polysilicon 114 -2840 114 -2840 0 3
rlabel polysilicon 121 -2834 121 -2834 0 1
rlabel polysilicon 121 -2840 121 -2840 0 3
rlabel polysilicon 128 -2834 128 -2834 0 1
rlabel polysilicon 131 -2834 131 -2834 0 2
rlabel polysilicon 128 -2840 128 -2840 0 3
rlabel polysilicon 135 -2834 135 -2834 0 1
rlabel polysilicon 135 -2840 135 -2840 0 3
rlabel polysilicon 142 -2834 142 -2834 0 1
rlabel polysilicon 142 -2840 142 -2840 0 3
rlabel polysilicon 149 -2834 149 -2834 0 1
rlabel polysilicon 149 -2840 149 -2840 0 3
rlabel polysilicon 156 -2834 156 -2834 0 1
rlabel polysilicon 156 -2840 156 -2840 0 3
rlabel polysilicon 163 -2834 163 -2834 0 1
rlabel polysilicon 166 -2834 166 -2834 0 2
rlabel polysilicon 163 -2840 163 -2840 0 3
rlabel polysilicon 170 -2834 170 -2834 0 1
rlabel polysilicon 170 -2840 170 -2840 0 3
rlabel polysilicon 180 -2834 180 -2834 0 2
rlabel polysilicon 177 -2840 177 -2840 0 3
rlabel polysilicon 180 -2840 180 -2840 0 4
rlabel polysilicon 184 -2834 184 -2834 0 1
rlabel polysilicon 184 -2840 184 -2840 0 3
rlabel polysilicon 191 -2840 191 -2840 0 3
rlabel polysilicon 198 -2834 198 -2834 0 1
rlabel polysilicon 198 -2840 198 -2840 0 3
rlabel polysilicon 205 -2834 205 -2834 0 1
rlabel polysilicon 205 -2840 205 -2840 0 3
rlabel polysilicon 212 -2834 212 -2834 0 1
rlabel polysilicon 212 -2840 212 -2840 0 3
rlabel polysilicon 219 -2834 219 -2834 0 1
rlabel polysilicon 219 -2840 219 -2840 0 3
rlabel polysilicon 226 -2834 226 -2834 0 1
rlabel polysilicon 229 -2834 229 -2834 0 2
rlabel polysilicon 226 -2840 226 -2840 0 3
rlabel polysilicon 229 -2840 229 -2840 0 4
rlabel polysilicon 233 -2834 233 -2834 0 1
rlabel polysilicon 233 -2840 233 -2840 0 3
rlabel polysilicon 240 -2834 240 -2834 0 1
rlabel polysilicon 240 -2840 240 -2840 0 3
rlabel polysilicon 247 -2834 247 -2834 0 1
rlabel polysilicon 250 -2834 250 -2834 0 2
rlabel polysilicon 250 -2840 250 -2840 0 4
rlabel polysilicon 254 -2834 254 -2834 0 1
rlabel polysilicon 254 -2840 254 -2840 0 3
rlabel polysilicon 261 -2834 261 -2834 0 1
rlabel polysilicon 261 -2840 261 -2840 0 3
rlabel polysilicon 268 -2834 268 -2834 0 1
rlabel polysilicon 268 -2840 268 -2840 0 3
rlabel polysilicon 275 -2834 275 -2834 0 1
rlabel polysilicon 278 -2834 278 -2834 0 2
rlabel polysilicon 275 -2840 275 -2840 0 3
rlabel polysilicon 282 -2834 282 -2834 0 1
rlabel polysilicon 282 -2840 282 -2840 0 3
rlabel polysilicon 289 -2834 289 -2834 0 1
rlabel polysilicon 289 -2840 289 -2840 0 3
rlabel polysilicon 296 -2834 296 -2834 0 1
rlabel polysilicon 296 -2840 296 -2840 0 3
rlabel polysilicon 303 -2834 303 -2834 0 1
rlabel polysilicon 303 -2840 303 -2840 0 3
rlabel polysilicon 310 -2834 310 -2834 0 1
rlabel polysilicon 310 -2840 310 -2840 0 3
rlabel polysilicon 317 -2834 317 -2834 0 1
rlabel polysilicon 317 -2840 317 -2840 0 3
rlabel polysilicon 324 -2834 324 -2834 0 1
rlabel polysilicon 324 -2840 324 -2840 0 3
rlabel polysilicon 331 -2834 331 -2834 0 1
rlabel polysilicon 331 -2840 331 -2840 0 3
rlabel polysilicon 338 -2834 338 -2834 0 1
rlabel polysilicon 338 -2840 338 -2840 0 3
rlabel polysilicon 345 -2834 345 -2834 0 1
rlabel polysilicon 345 -2840 345 -2840 0 3
rlabel polysilicon 352 -2834 352 -2834 0 1
rlabel polysilicon 352 -2840 352 -2840 0 3
rlabel polysilicon 359 -2834 359 -2834 0 1
rlabel polysilicon 359 -2840 359 -2840 0 3
rlabel polysilicon 366 -2834 366 -2834 0 1
rlabel polysilicon 366 -2840 366 -2840 0 3
rlabel polysilicon 373 -2834 373 -2834 0 1
rlabel polysilicon 373 -2840 373 -2840 0 3
rlabel polysilicon 380 -2834 380 -2834 0 1
rlabel polysilicon 383 -2834 383 -2834 0 2
rlabel polysilicon 380 -2840 380 -2840 0 3
rlabel polysilicon 387 -2834 387 -2834 0 1
rlabel polysilicon 387 -2840 387 -2840 0 3
rlabel polysilicon 394 -2834 394 -2834 0 1
rlabel polysilicon 394 -2840 394 -2840 0 3
rlabel polysilicon 401 -2834 401 -2834 0 1
rlabel polysilicon 401 -2840 401 -2840 0 3
rlabel polysilicon 408 -2834 408 -2834 0 1
rlabel polysilicon 408 -2840 408 -2840 0 3
rlabel polysilicon 415 -2834 415 -2834 0 1
rlabel polysilicon 415 -2840 415 -2840 0 3
rlabel polysilicon 422 -2834 422 -2834 0 1
rlabel polysilicon 422 -2840 422 -2840 0 3
rlabel polysilicon 429 -2834 429 -2834 0 1
rlabel polysilicon 429 -2840 429 -2840 0 3
rlabel polysilicon 436 -2834 436 -2834 0 1
rlabel polysilicon 436 -2840 436 -2840 0 3
rlabel polysilicon 443 -2834 443 -2834 0 1
rlabel polysilicon 443 -2840 443 -2840 0 3
rlabel polysilicon 450 -2834 450 -2834 0 1
rlabel polysilicon 450 -2840 450 -2840 0 3
rlabel polysilicon 457 -2834 457 -2834 0 1
rlabel polysilicon 457 -2840 457 -2840 0 3
rlabel polysilicon 464 -2834 464 -2834 0 1
rlabel polysilicon 464 -2840 464 -2840 0 3
rlabel polysilicon 471 -2834 471 -2834 0 1
rlabel polysilicon 471 -2840 471 -2840 0 3
rlabel polysilicon 478 -2834 478 -2834 0 1
rlabel polysilicon 478 -2840 478 -2840 0 3
rlabel polysilicon 485 -2834 485 -2834 0 1
rlabel polysilicon 485 -2840 485 -2840 0 3
rlabel polysilicon 492 -2834 492 -2834 0 1
rlabel polysilicon 492 -2840 492 -2840 0 3
rlabel polysilicon 499 -2834 499 -2834 0 1
rlabel polysilicon 499 -2840 499 -2840 0 3
rlabel polysilicon 506 -2834 506 -2834 0 1
rlabel polysilicon 506 -2840 506 -2840 0 3
rlabel polysilicon 513 -2834 513 -2834 0 1
rlabel polysilicon 513 -2840 513 -2840 0 3
rlabel polysilicon 520 -2834 520 -2834 0 1
rlabel polysilicon 523 -2834 523 -2834 0 2
rlabel polysilicon 520 -2840 520 -2840 0 3
rlabel polysilicon 523 -2840 523 -2840 0 4
rlabel polysilicon 527 -2834 527 -2834 0 1
rlabel polysilicon 527 -2840 527 -2840 0 3
rlabel polysilicon 534 -2834 534 -2834 0 1
rlabel polysilicon 534 -2840 534 -2840 0 3
rlabel polysilicon 541 -2834 541 -2834 0 1
rlabel polysilicon 541 -2840 541 -2840 0 3
rlabel polysilicon 548 -2834 548 -2834 0 1
rlabel polysilicon 548 -2840 548 -2840 0 3
rlabel polysilicon 555 -2834 555 -2834 0 1
rlabel polysilicon 555 -2840 555 -2840 0 3
rlabel polysilicon 562 -2834 562 -2834 0 1
rlabel polysilicon 562 -2840 562 -2840 0 3
rlabel polysilicon 569 -2834 569 -2834 0 1
rlabel polysilicon 569 -2840 569 -2840 0 3
rlabel polysilicon 576 -2834 576 -2834 0 1
rlabel polysilicon 576 -2840 576 -2840 0 3
rlabel polysilicon 583 -2834 583 -2834 0 1
rlabel polysilicon 583 -2840 583 -2840 0 3
rlabel polysilicon 590 -2834 590 -2834 0 1
rlabel polysilicon 593 -2834 593 -2834 0 2
rlabel polysilicon 590 -2840 590 -2840 0 3
rlabel polysilicon 593 -2840 593 -2840 0 4
rlabel polysilicon 597 -2834 597 -2834 0 1
rlabel polysilicon 597 -2840 597 -2840 0 3
rlabel polysilicon 604 -2834 604 -2834 0 1
rlabel polysilicon 604 -2840 604 -2840 0 3
rlabel polysilicon 611 -2834 611 -2834 0 1
rlabel polysilicon 611 -2840 611 -2840 0 3
rlabel polysilicon 618 -2834 618 -2834 0 1
rlabel polysilicon 618 -2840 618 -2840 0 3
rlabel polysilicon 625 -2834 625 -2834 0 1
rlabel polysilicon 625 -2840 625 -2840 0 3
rlabel polysilicon 632 -2834 632 -2834 0 1
rlabel polysilicon 632 -2840 632 -2840 0 3
rlabel polysilicon 639 -2834 639 -2834 0 1
rlabel polysilicon 639 -2840 639 -2840 0 3
rlabel polysilicon 649 -2834 649 -2834 0 2
rlabel polysilicon 646 -2840 646 -2840 0 3
rlabel polysilicon 649 -2840 649 -2840 0 4
rlabel polysilicon 653 -2834 653 -2834 0 1
rlabel polysilicon 653 -2840 653 -2840 0 3
rlabel polysilicon 656 -2840 656 -2840 0 4
rlabel polysilicon 660 -2834 660 -2834 0 1
rlabel polysilicon 660 -2840 660 -2840 0 3
rlabel polysilicon 667 -2834 667 -2834 0 1
rlabel polysilicon 667 -2840 667 -2840 0 3
rlabel polysilicon 674 -2834 674 -2834 0 1
rlabel polysilicon 674 -2840 674 -2840 0 3
rlabel polysilicon 681 -2834 681 -2834 0 1
rlabel polysilicon 684 -2834 684 -2834 0 2
rlabel polysilicon 684 -2840 684 -2840 0 4
rlabel polysilicon 688 -2834 688 -2834 0 1
rlabel polysilicon 688 -2840 688 -2840 0 3
rlabel polysilicon 695 -2834 695 -2834 0 1
rlabel polysilicon 695 -2840 695 -2840 0 3
rlabel polysilicon 702 -2834 702 -2834 0 1
rlabel polysilicon 702 -2840 702 -2840 0 3
rlabel polysilicon 709 -2834 709 -2834 0 1
rlabel polysilicon 709 -2840 709 -2840 0 3
rlabel polysilicon 716 -2834 716 -2834 0 1
rlabel polysilicon 716 -2840 716 -2840 0 3
rlabel polysilicon 723 -2834 723 -2834 0 1
rlabel polysilicon 723 -2840 723 -2840 0 3
rlabel polysilicon 730 -2834 730 -2834 0 1
rlabel polysilicon 730 -2840 730 -2840 0 3
rlabel polysilicon 737 -2834 737 -2834 0 1
rlabel polysilicon 737 -2840 737 -2840 0 3
rlabel polysilicon 744 -2834 744 -2834 0 1
rlabel polysilicon 744 -2840 744 -2840 0 3
rlabel polysilicon 751 -2834 751 -2834 0 1
rlabel polysilicon 751 -2840 751 -2840 0 3
rlabel polysilicon 758 -2834 758 -2834 0 1
rlabel polysilicon 761 -2834 761 -2834 0 2
rlabel polysilicon 758 -2840 758 -2840 0 3
rlabel polysilicon 761 -2840 761 -2840 0 4
rlabel polysilicon 765 -2834 765 -2834 0 1
rlabel polysilicon 768 -2834 768 -2834 0 2
rlabel polysilicon 765 -2840 765 -2840 0 3
rlabel polysilicon 768 -2840 768 -2840 0 4
rlabel polysilicon 772 -2834 772 -2834 0 1
rlabel polysilicon 775 -2834 775 -2834 0 2
rlabel polysilicon 775 -2840 775 -2840 0 4
rlabel polysilicon 779 -2834 779 -2834 0 1
rlabel polysilicon 779 -2840 779 -2840 0 3
rlabel polysilicon 786 -2834 786 -2834 0 1
rlabel polysilicon 786 -2840 786 -2840 0 3
rlabel polysilicon 793 -2834 793 -2834 0 1
rlabel polysilicon 793 -2840 793 -2840 0 3
rlabel polysilicon 800 -2834 800 -2834 0 1
rlabel polysilicon 803 -2834 803 -2834 0 2
rlabel polysilicon 800 -2840 800 -2840 0 3
rlabel polysilicon 803 -2840 803 -2840 0 4
rlabel polysilicon 807 -2834 807 -2834 0 1
rlabel polysilicon 807 -2840 807 -2840 0 3
rlabel polysilicon 814 -2834 814 -2834 0 1
rlabel polysilicon 814 -2840 814 -2840 0 3
rlabel polysilicon 821 -2834 821 -2834 0 1
rlabel polysilicon 821 -2840 821 -2840 0 3
rlabel polysilicon 828 -2834 828 -2834 0 1
rlabel polysilicon 828 -2840 828 -2840 0 3
rlabel polysilicon 835 -2834 835 -2834 0 1
rlabel polysilicon 835 -2840 835 -2840 0 3
rlabel polysilicon 842 -2834 842 -2834 0 1
rlabel polysilicon 842 -2840 842 -2840 0 3
rlabel polysilicon 849 -2834 849 -2834 0 1
rlabel polysilicon 849 -2840 849 -2840 0 3
rlabel polysilicon 856 -2834 856 -2834 0 1
rlabel polysilicon 856 -2840 856 -2840 0 3
rlabel polysilicon 863 -2834 863 -2834 0 1
rlabel polysilicon 863 -2840 863 -2840 0 3
rlabel polysilicon 870 -2834 870 -2834 0 1
rlabel polysilicon 870 -2840 870 -2840 0 3
rlabel polysilicon 877 -2834 877 -2834 0 1
rlabel polysilicon 877 -2840 877 -2840 0 3
rlabel polysilicon 884 -2834 884 -2834 0 1
rlabel polysilicon 887 -2834 887 -2834 0 2
rlabel polysilicon 884 -2840 884 -2840 0 3
rlabel polysilicon 887 -2840 887 -2840 0 4
rlabel polysilicon 891 -2834 891 -2834 0 1
rlabel polysilicon 894 -2834 894 -2834 0 2
rlabel polysilicon 891 -2840 891 -2840 0 3
rlabel polysilicon 898 -2834 898 -2834 0 1
rlabel polysilicon 901 -2834 901 -2834 0 2
rlabel polysilicon 898 -2840 898 -2840 0 3
rlabel polysilicon 901 -2840 901 -2840 0 4
rlabel polysilicon 905 -2834 905 -2834 0 1
rlabel polysilicon 905 -2840 905 -2840 0 3
rlabel polysilicon 912 -2834 912 -2834 0 1
rlabel polysilicon 912 -2840 912 -2840 0 3
rlabel polysilicon 919 -2834 919 -2834 0 1
rlabel polysilicon 919 -2840 919 -2840 0 3
rlabel polysilicon 926 -2834 926 -2834 0 1
rlabel polysilicon 926 -2840 926 -2840 0 3
rlabel polysilicon 933 -2834 933 -2834 0 1
rlabel polysilicon 933 -2840 933 -2840 0 3
rlabel polysilicon 940 -2834 940 -2834 0 1
rlabel polysilicon 940 -2840 940 -2840 0 3
rlabel polysilicon 947 -2834 947 -2834 0 1
rlabel polysilicon 947 -2840 947 -2840 0 3
rlabel polysilicon 954 -2834 954 -2834 0 1
rlabel polysilicon 954 -2840 954 -2840 0 3
rlabel polysilicon 961 -2834 961 -2834 0 1
rlabel polysilicon 961 -2840 961 -2840 0 3
rlabel polysilicon 968 -2834 968 -2834 0 1
rlabel polysilicon 968 -2840 968 -2840 0 3
rlabel polysilicon 975 -2834 975 -2834 0 1
rlabel polysilicon 975 -2840 975 -2840 0 3
rlabel polysilicon 982 -2834 982 -2834 0 1
rlabel polysilicon 985 -2834 985 -2834 0 2
rlabel polysilicon 982 -2840 982 -2840 0 3
rlabel polysilicon 989 -2834 989 -2834 0 1
rlabel polysilicon 989 -2840 989 -2840 0 3
rlabel polysilicon 996 -2834 996 -2834 0 1
rlabel polysilicon 999 -2834 999 -2834 0 2
rlabel polysilicon 996 -2840 996 -2840 0 3
rlabel polysilicon 999 -2840 999 -2840 0 4
rlabel polysilicon 1003 -2834 1003 -2834 0 1
rlabel polysilicon 1003 -2840 1003 -2840 0 3
rlabel polysilicon 1010 -2834 1010 -2834 0 1
rlabel polysilicon 1010 -2840 1010 -2840 0 3
rlabel polysilicon 1017 -2834 1017 -2834 0 1
rlabel polysilicon 1017 -2840 1017 -2840 0 3
rlabel polysilicon 1024 -2834 1024 -2834 0 1
rlabel polysilicon 1024 -2840 1024 -2840 0 3
rlabel polysilicon 1031 -2834 1031 -2834 0 1
rlabel polysilicon 1031 -2840 1031 -2840 0 3
rlabel polysilicon 1038 -2834 1038 -2834 0 1
rlabel polysilicon 1038 -2840 1038 -2840 0 3
rlabel polysilicon 1045 -2834 1045 -2834 0 1
rlabel polysilicon 1048 -2834 1048 -2834 0 2
rlabel polysilicon 1045 -2840 1045 -2840 0 3
rlabel polysilicon 1048 -2840 1048 -2840 0 4
rlabel polysilicon 1052 -2834 1052 -2834 0 1
rlabel polysilicon 1052 -2840 1052 -2840 0 3
rlabel polysilicon 1059 -2834 1059 -2834 0 1
rlabel polysilicon 1059 -2840 1059 -2840 0 3
rlabel polysilicon 1066 -2834 1066 -2834 0 1
rlabel polysilicon 1066 -2840 1066 -2840 0 3
rlabel polysilicon 1073 -2834 1073 -2834 0 1
rlabel polysilicon 1073 -2840 1073 -2840 0 3
rlabel polysilicon 1080 -2834 1080 -2834 0 1
rlabel polysilicon 1080 -2840 1080 -2840 0 3
rlabel polysilicon 1087 -2834 1087 -2834 0 1
rlabel polysilicon 1087 -2840 1087 -2840 0 3
rlabel polysilicon 1094 -2834 1094 -2834 0 1
rlabel polysilicon 1097 -2834 1097 -2834 0 2
rlabel polysilicon 1097 -2840 1097 -2840 0 4
rlabel polysilicon 1101 -2834 1101 -2834 0 1
rlabel polysilicon 1101 -2840 1101 -2840 0 3
rlabel polysilicon 1108 -2834 1108 -2834 0 1
rlabel polysilicon 1108 -2840 1108 -2840 0 3
rlabel polysilicon 1115 -2834 1115 -2834 0 1
rlabel polysilicon 1115 -2840 1115 -2840 0 3
rlabel polysilicon 1118 -2840 1118 -2840 0 4
rlabel polysilicon 1122 -2834 1122 -2834 0 1
rlabel polysilicon 1122 -2840 1122 -2840 0 3
rlabel polysilicon 1129 -2834 1129 -2834 0 1
rlabel polysilicon 1129 -2840 1129 -2840 0 3
rlabel polysilicon 1136 -2834 1136 -2834 0 1
rlabel polysilicon 1136 -2840 1136 -2840 0 3
rlabel polysilicon 1143 -2834 1143 -2834 0 1
rlabel polysilicon 1143 -2840 1143 -2840 0 3
rlabel polysilicon 1150 -2834 1150 -2834 0 1
rlabel polysilicon 1150 -2840 1150 -2840 0 3
rlabel polysilicon 1157 -2834 1157 -2834 0 1
rlabel polysilicon 1157 -2840 1157 -2840 0 3
rlabel polysilicon 1164 -2834 1164 -2834 0 1
rlabel polysilicon 1164 -2840 1164 -2840 0 3
rlabel polysilicon 1171 -2834 1171 -2834 0 1
rlabel polysilicon 1171 -2840 1171 -2840 0 3
rlabel polysilicon 1178 -2834 1178 -2834 0 1
rlabel polysilicon 1178 -2840 1178 -2840 0 3
rlabel polysilicon 1185 -2834 1185 -2834 0 1
rlabel polysilicon 1188 -2834 1188 -2834 0 2
rlabel polysilicon 1185 -2840 1185 -2840 0 3
rlabel polysilicon 1188 -2840 1188 -2840 0 4
rlabel polysilicon 1192 -2834 1192 -2834 0 1
rlabel polysilicon 1192 -2840 1192 -2840 0 3
rlabel polysilicon 1199 -2834 1199 -2834 0 1
rlabel polysilicon 1199 -2840 1199 -2840 0 3
rlabel polysilicon 1206 -2834 1206 -2834 0 1
rlabel polysilicon 1206 -2840 1206 -2840 0 3
rlabel polysilicon 1213 -2834 1213 -2834 0 1
rlabel polysilicon 1213 -2840 1213 -2840 0 3
rlabel polysilicon 1220 -2834 1220 -2834 0 1
rlabel polysilicon 1220 -2840 1220 -2840 0 3
rlabel polysilicon 1227 -2834 1227 -2834 0 1
rlabel polysilicon 1227 -2840 1227 -2840 0 3
rlabel polysilicon 1234 -2834 1234 -2834 0 1
rlabel polysilicon 1234 -2840 1234 -2840 0 3
rlabel polysilicon 1241 -2834 1241 -2834 0 1
rlabel polysilicon 1241 -2840 1241 -2840 0 3
rlabel polysilicon 1248 -2834 1248 -2834 0 1
rlabel polysilicon 1248 -2840 1248 -2840 0 3
rlabel polysilicon 1255 -2834 1255 -2834 0 1
rlabel polysilicon 1255 -2840 1255 -2840 0 3
rlabel polysilicon 1262 -2834 1262 -2834 0 1
rlabel polysilicon 1262 -2840 1262 -2840 0 3
rlabel polysilicon 1269 -2834 1269 -2834 0 1
rlabel polysilicon 1269 -2840 1269 -2840 0 3
rlabel polysilicon 1276 -2834 1276 -2834 0 1
rlabel polysilicon 1279 -2834 1279 -2834 0 2
rlabel polysilicon 1279 -2840 1279 -2840 0 4
rlabel polysilicon 1283 -2834 1283 -2834 0 1
rlabel polysilicon 1283 -2840 1283 -2840 0 3
rlabel polysilicon 1290 -2834 1290 -2834 0 1
rlabel polysilicon 1290 -2840 1290 -2840 0 3
rlabel polysilicon 1297 -2834 1297 -2834 0 1
rlabel polysilicon 1297 -2840 1297 -2840 0 3
rlabel polysilicon 1304 -2834 1304 -2834 0 1
rlabel polysilicon 1304 -2840 1304 -2840 0 3
rlabel polysilicon 1311 -2834 1311 -2834 0 1
rlabel polysilicon 1311 -2840 1311 -2840 0 3
rlabel polysilicon 1318 -2834 1318 -2834 0 1
rlabel polysilicon 1318 -2840 1318 -2840 0 3
rlabel polysilicon 1325 -2834 1325 -2834 0 1
rlabel polysilicon 1325 -2840 1325 -2840 0 3
rlabel polysilicon 1332 -2834 1332 -2834 0 1
rlabel polysilicon 1332 -2840 1332 -2840 0 3
rlabel polysilicon 1339 -2834 1339 -2834 0 1
rlabel polysilicon 1339 -2840 1339 -2840 0 3
rlabel polysilicon 1346 -2834 1346 -2834 0 1
rlabel polysilicon 1346 -2840 1346 -2840 0 3
rlabel polysilicon 1353 -2834 1353 -2834 0 1
rlabel polysilicon 1353 -2840 1353 -2840 0 3
rlabel polysilicon 1360 -2834 1360 -2834 0 1
rlabel polysilicon 1360 -2840 1360 -2840 0 3
rlabel polysilicon 1367 -2834 1367 -2834 0 1
rlabel polysilicon 1367 -2840 1367 -2840 0 3
rlabel polysilicon 1374 -2834 1374 -2834 0 1
rlabel polysilicon 1374 -2840 1374 -2840 0 3
rlabel polysilicon 1381 -2834 1381 -2834 0 1
rlabel polysilicon 1381 -2840 1381 -2840 0 3
rlabel polysilicon 1388 -2834 1388 -2834 0 1
rlabel polysilicon 1388 -2840 1388 -2840 0 3
rlabel polysilicon 1395 -2834 1395 -2834 0 1
rlabel polysilicon 1395 -2840 1395 -2840 0 3
rlabel polysilicon 1402 -2834 1402 -2834 0 1
rlabel polysilicon 1402 -2840 1402 -2840 0 3
rlabel polysilicon 1409 -2834 1409 -2834 0 1
rlabel polysilicon 1409 -2840 1409 -2840 0 3
rlabel polysilicon 1416 -2834 1416 -2834 0 1
rlabel polysilicon 1416 -2840 1416 -2840 0 3
rlabel polysilicon 1423 -2834 1423 -2834 0 1
rlabel polysilicon 1423 -2840 1423 -2840 0 3
rlabel polysilicon 1430 -2834 1430 -2834 0 1
rlabel polysilicon 1430 -2840 1430 -2840 0 3
rlabel polysilicon 1437 -2834 1437 -2834 0 1
rlabel polysilicon 1437 -2840 1437 -2840 0 3
rlabel polysilicon 1444 -2834 1444 -2834 0 1
rlabel polysilicon 1444 -2840 1444 -2840 0 3
rlabel polysilicon 1451 -2834 1451 -2834 0 1
rlabel polysilicon 1451 -2840 1451 -2840 0 3
rlabel polysilicon 1458 -2834 1458 -2834 0 1
rlabel polysilicon 1458 -2840 1458 -2840 0 3
rlabel polysilicon 1465 -2834 1465 -2834 0 1
rlabel polysilicon 1465 -2840 1465 -2840 0 3
rlabel polysilicon 1472 -2834 1472 -2834 0 1
rlabel polysilicon 1472 -2840 1472 -2840 0 3
rlabel polysilicon 1479 -2834 1479 -2834 0 1
rlabel polysilicon 1479 -2840 1479 -2840 0 3
rlabel polysilicon 1486 -2834 1486 -2834 0 1
rlabel polysilicon 1486 -2840 1486 -2840 0 3
rlabel polysilicon 1493 -2834 1493 -2834 0 1
rlabel polysilicon 1493 -2840 1493 -2840 0 3
rlabel polysilicon 1500 -2834 1500 -2834 0 1
rlabel polysilicon 1500 -2840 1500 -2840 0 3
rlabel polysilicon 1507 -2834 1507 -2834 0 1
rlabel polysilicon 1510 -2834 1510 -2834 0 2
rlabel polysilicon 1507 -2840 1507 -2840 0 3
rlabel polysilicon 1510 -2840 1510 -2840 0 4
rlabel polysilicon 1514 -2834 1514 -2834 0 1
rlabel polysilicon 1514 -2840 1514 -2840 0 3
rlabel polysilicon 1521 -2834 1521 -2834 0 1
rlabel polysilicon 1521 -2840 1521 -2840 0 3
rlabel polysilicon 1528 -2834 1528 -2834 0 1
rlabel polysilicon 1528 -2840 1528 -2840 0 3
rlabel polysilicon 1535 -2834 1535 -2834 0 1
rlabel polysilicon 1535 -2840 1535 -2840 0 3
rlabel polysilicon 1542 -2834 1542 -2834 0 1
rlabel polysilicon 1542 -2840 1542 -2840 0 3
rlabel polysilicon 1549 -2834 1549 -2834 0 1
rlabel polysilicon 1549 -2840 1549 -2840 0 3
rlabel polysilicon 1556 -2834 1556 -2834 0 1
rlabel polysilicon 1556 -2840 1556 -2840 0 3
rlabel polysilicon 30 -2945 30 -2945 0 1
rlabel polysilicon 30 -2951 30 -2951 0 3
rlabel polysilicon 37 -2945 37 -2945 0 1
rlabel polysilicon 37 -2951 37 -2951 0 3
rlabel polysilicon 44 -2945 44 -2945 0 1
rlabel polysilicon 44 -2951 44 -2951 0 3
rlabel polysilicon 51 -2945 51 -2945 0 1
rlabel polysilicon 51 -2951 51 -2951 0 3
rlabel polysilicon 58 -2945 58 -2945 0 1
rlabel polysilicon 58 -2951 58 -2951 0 3
rlabel polysilicon 65 -2945 65 -2945 0 1
rlabel polysilicon 65 -2951 65 -2951 0 3
rlabel polysilicon 72 -2945 72 -2945 0 1
rlabel polysilicon 75 -2945 75 -2945 0 2
rlabel polysilicon 79 -2945 79 -2945 0 1
rlabel polysilicon 79 -2951 79 -2951 0 3
rlabel polysilicon 86 -2945 86 -2945 0 1
rlabel polysilicon 86 -2951 86 -2951 0 3
rlabel polysilicon 93 -2945 93 -2945 0 1
rlabel polysilicon 93 -2951 93 -2951 0 3
rlabel polysilicon 100 -2945 100 -2945 0 1
rlabel polysilicon 100 -2951 100 -2951 0 3
rlabel polysilicon 107 -2945 107 -2945 0 1
rlabel polysilicon 107 -2951 107 -2951 0 3
rlabel polysilicon 114 -2945 114 -2945 0 1
rlabel polysilicon 117 -2945 117 -2945 0 2
rlabel polysilicon 114 -2951 114 -2951 0 3
rlabel polysilicon 121 -2945 121 -2945 0 1
rlabel polysilicon 121 -2951 121 -2951 0 3
rlabel polysilicon 128 -2945 128 -2945 0 1
rlabel polysilicon 128 -2951 128 -2951 0 3
rlabel polysilicon 135 -2945 135 -2945 0 1
rlabel polysilicon 135 -2951 135 -2951 0 3
rlabel polysilicon 142 -2945 142 -2945 0 1
rlabel polysilicon 142 -2951 142 -2951 0 3
rlabel polysilicon 149 -2945 149 -2945 0 1
rlabel polysilicon 149 -2951 149 -2951 0 3
rlabel polysilicon 159 -2951 159 -2951 0 4
rlabel polysilicon 163 -2945 163 -2945 0 1
rlabel polysilicon 163 -2951 163 -2951 0 3
rlabel polysilicon 170 -2945 170 -2945 0 1
rlabel polysilicon 170 -2951 170 -2951 0 3
rlabel polysilicon 177 -2945 177 -2945 0 1
rlabel polysilicon 177 -2951 177 -2951 0 3
rlabel polysilicon 180 -2951 180 -2951 0 4
rlabel polysilicon 184 -2945 184 -2945 0 1
rlabel polysilicon 184 -2951 184 -2951 0 3
rlabel polysilicon 191 -2945 191 -2945 0 1
rlabel polysilicon 191 -2951 191 -2951 0 3
rlabel polysilicon 198 -2945 198 -2945 0 1
rlabel polysilicon 198 -2951 198 -2951 0 3
rlabel polysilicon 205 -2945 205 -2945 0 1
rlabel polysilicon 205 -2951 205 -2951 0 3
rlabel polysilicon 212 -2945 212 -2945 0 1
rlabel polysilicon 212 -2951 212 -2951 0 3
rlabel polysilicon 219 -2945 219 -2945 0 1
rlabel polysilicon 219 -2951 219 -2951 0 3
rlabel polysilicon 226 -2945 226 -2945 0 1
rlabel polysilicon 226 -2951 226 -2951 0 3
rlabel polysilicon 233 -2945 233 -2945 0 1
rlabel polysilicon 233 -2951 233 -2951 0 3
rlabel polysilicon 240 -2945 240 -2945 0 1
rlabel polysilicon 240 -2951 240 -2951 0 3
rlabel polysilicon 247 -2945 247 -2945 0 1
rlabel polysilicon 250 -2945 250 -2945 0 2
rlabel polysilicon 250 -2951 250 -2951 0 4
rlabel polysilicon 254 -2945 254 -2945 0 1
rlabel polysilicon 257 -2945 257 -2945 0 2
rlabel polysilicon 254 -2951 254 -2951 0 3
rlabel polysilicon 257 -2951 257 -2951 0 4
rlabel polysilicon 264 -2945 264 -2945 0 2
rlabel polysilicon 261 -2951 261 -2951 0 3
rlabel polysilicon 264 -2951 264 -2951 0 4
rlabel polysilicon 268 -2945 268 -2945 0 1
rlabel polysilicon 268 -2951 268 -2951 0 3
rlabel polysilicon 275 -2945 275 -2945 0 1
rlabel polysilicon 275 -2951 275 -2951 0 3
rlabel polysilicon 282 -2945 282 -2945 0 1
rlabel polysilicon 282 -2951 282 -2951 0 3
rlabel polysilicon 289 -2945 289 -2945 0 1
rlabel polysilicon 289 -2951 289 -2951 0 3
rlabel polysilicon 296 -2945 296 -2945 0 1
rlabel polysilicon 296 -2951 296 -2951 0 3
rlabel polysilicon 303 -2945 303 -2945 0 1
rlabel polysilicon 303 -2951 303 -2951 0 3
rlabel polysilicon 310 -2945 310 -2945 0 1
rlabel polysilicon 310 -2951 310 -2951 0 3
rlabel polysilicon 317 -2945 317 -2945 0 1
rlabel polysilicon 317 -2951 317 -2951 0 3
rlabel polysilicon 324 -2945 324 -2945 0 1
rlabel polysilicon 324 -2951 324 -2951 0 3
rlabel polysilicon 331 -2945 331 -2945 0 1
rlabel polysilicon 331 -2951 331 -2951 0 3
rlabel polysilicon 338 -2945 338 -2945 0 1
rlabel polysilicon 338 -2951 338 -2951 0 3
rlabel polysilicon 345 -2945 345 -2945 0 1
rlabel polysilicon 345 -2951 345 -2951 0 3
rlabel polysilicon 352 -2945 352 -2945 0 1
rlabel polysilicon 352 -2951 352 -2951 0 3
rlabel polysilicon 359 -2945 359 -2945 0 1
rlabel polysilicon 359 -2951 359 -2951 0 3
rlabel polysilicon 366 -2945 366 -2945 0 1
rlabel polysilicon 366 -2951 366 -2951 0 3
rlabel polysilicon 373 -2951 373 -2951 0 3
rlabel polysilicon 376 -2951 376 -2951 0 4
rlabel polysilicon 380 -2945 380 -2945 0 1
rlabel polysilicon 380 -2951 380 -2951 0 3
rlabel polysilicon 387 -2945 387 -2945 0 1
rlabel polysilicon 387 -2951 387 -2951 0 3
rlabel polysilicon 394 -2945 394 -2945 0 1
rlabel polysilicon 394 -2951 394 -2951 0 3
rlabel polysilicon 401 -2945 401 -2945 0 1
rlabel polysilicon 404 -2945 404 -2945 0 2
rlabel polysilicon 401 -2951 401 -2951 0 3
rlabel polysilicon 404 -2951 404 -2951 0 4
rlabel polysilicon 408 -2945 408 -2945 0 1
rlabel polysilicon 411 -2945 411 -2945 0 2
rlabel polysilicon 408 -2951 408 -2951 0 3
rlabel polysilicon 415 -2945 415 -2945 0 1
rlabel polysilicon 415 -2951 415 -2951 0 3
rlabel polysilicon 422 -2945 422 -2945 0 1
rlabel polysilicon 422 -2951 422 -2951 0 3
rlabel polysilicon 429 -2945 429 -2945 0 1
rlabel polysilicon 429 -2951 429 -2951 0 3
rlabel polysilicon 436 -2945 436 -2945 0 1
rlabel polysilicon 436 -2951 436 -2951 0 3
rlabel polysilicon 443 -2945 443 -2945 0 1
rlabel polysilicon 443 -2951 443 -2951 0 3
rlabel polysilicon 450 -2945 450 -2945 0 1
rlabel polysilicon 450 -2951 450 -2951 0 3
rlabel polysilicon 457 -2945 457 -2945 0 1
rlabel polysilicon 457 -2951 457 -2951 0 3
rlabel polysilicon 464 -2945 464 -2945 0 1
rlabel polysilicon 464 -2951 464 -2951 0 3
rlabel polysilicon 471 -2945 471 -2945 0 1
rlabel polysilicon 474 -2945 474 -2945 0 2
rlabel polysilicon 471 -2951 471 -2951 0 3
rlabel polysilicon 474 -2951 474 -2951 0 4
rlabel polysilicon 478 -2945 478 -2945 0 1
rlabel polysilicon 478 -2951 478 -2951 0 3
rlabel polysilicon 481 -2951 481 -2951 0 4
rlabel polysilicon 485 -2945 485 -2945 0 1
rlabel polysilicon 485 -2951 485 -2951 0 3
rlabel polysilicon 492 -2945 492 -2945 0 1
rlabel polysilicon 492 -2951 492 -2951 0 3
rlabel polysilicon 499 -2945 499 -2945 0 1
rlabel polysilicon 502 -2945 502 -2945 0 2
rlabel polysilicon 502 -2951 502 -2951 0 4
rlabel polysilicon 506 -2945 506 -2945 0 1
rlabel polysilicon 506 -2951 506 -2951 0 3
rlabel polysilicon 513 -2945 513 -2945 0 1
rlabel polysilicon 513 -2951 513 -2951 0 3
rlabel polysilicon 520 -2945 520 -2945 0 1
rlabel polysilicon 520 -2951 520 -2951 0 3
rlabel polysilicon 527 -2945 527 -2945 0 1
rlabel polysilicon 527 -2951 527 -2951 0 3
rlabel polysilicon 534 -2945 534 -2945 0 1
rlabel polysilicon 534 -2951 534 -2951 0 3
rlabel polysilicon 541 -2945 541 -2945 0 1
rlabel polysilicon 541 -2951 541 -2951 0 3
rlabel polysilicon 548 -2945 548 -2945 0 1
rlabel polysilicon 548 -2951 548 -2951 0 3
rlabel polysilicon 555 -2945 555 -2945 0 1
rlabel polysilicon 555 -2951 555 -2951 0 3
rlabel polysilicon 562 -2945 562 -2945 0 1
rlabel polysilicon 565 -2945 565 -2945 0 2
rlabel polysilicon 565 -2951 565 -2951 0 4
rlabel polysilicon 569 -2945 569 -2945 0 1
rlabel polysilicon 569 -2951 569 -2951 0 3
rlabel polysilicon 576 -2945 576 -2945 0 1
rlabel polysilicon 576 -2951 576 -2951 0 3
rlabel polysilicon 583 -2945 583 -2945 0 1
rlabel polysilicon 583 -2951 583 -2951 0 3
rlabel polysilicon 590 -2945 590 -2945 0 1
rlabel polysilicon 590 -2951 590 -2951 0 3
rlabel polysilicon 597 -2945 597 -2945 0 1
rlabel polysilicon 597 -2951 597 -2951 0 3
rlabel polysilicon 607 -2945 607 -2945 0 2
rlabel polysilicon 604 -2951 604 -2951 0 3
rlabel polysilicon 607 -2951 607 -2951 0 4
rlabel polysilicon 611 -2945 611 -2945 0 1
rlabel polysilicon 611 -2951 611 -2951 0 3
rlabel polysilicon 618 -2945 618 -2945 0 1
rlabel polysilicon 618 -2951 618 -2951 0 3
rlabel polysilicon 625 -2945 625 -2945 0 1
rlabel polysilicon 625 -2951 625 -2951 0 3
rlabel polysilicon 632 -2945 632 -2945 0 1
rlabel polysilicon 632 -2951 632 -2951 0 3
rlabel polysilicon 635 -2951 635 -2951 0 4
rlabel polysilicon 639 -2945 639 -2945 0 1
rlabel polysilicon 639 -2951 639 -2951 0 3
rlabel polysilicon 646 -2945 646 -2945 0 1
rlabel polysilicon 646 -2951 646 -2951 0 3
rlabel polysilicon 653 -2945 653 -2945 0 1
rlabel polysilicon 653 -2951 653 -2951 0 3
rlabel polysilicon 660 -2945 660 -2945 0 1
rlabel polysilicon 660 -2951 660 -2951 0 3
rlabel polysilicon 667 -2945 667 -2945 0 1
rlabel polysilicon 670 -2945 670 -2945 0 2
rlabel polysilicon 667 -2951 667 -2951 0 3
rlabel polysilicon 670 -2951 670 -2951 0 4
rlabel polysilicon 674 -2945 674 -2945 0 1
rlabel polysilicon 674 -2951 674 -2951 0 3
rlabel polysilicon 681 -2945 681 -2945 0 1
rlabel polysilicon 681 -2951 681 -2951 0 3
rlabel polysilicon 688 -2951 688 -2951 0 3
rlabel polysilicon 691 -2951 691 -2951 0 4
rlabel polysilicon 695 -2945 695 -2945 0 1
rlabel polysilicon 695 -2951 695 -2951 0 3
rlabel polysilicon 702 -2945 702 -2945 0 1
rlabel polysilicon 702 -2951 702 -2951 0 3
rlabel polysilicon 705 -2951 705 -2951 0 4
rlabel polysilicon 709 -2945 709 -2945 0 1
rlabel polysilicon 709 -2951 709 -2951 0 3
rlabel polysilicon 716 -2945 716 -2945 0 1
rlabel polysilicon 716 -2951 716 -2951 0 3
rlabel polysilicon 723 -2945 723 -2945 0 1
rlabel polysilicon 723 -2951 723 -2951 0 3
rlabel polysilicon 730 -2945 730 -2945 0 1
rlabel polysilicon 733 -2945 733 -2945 0 2
rlabel polysilicon 730 -2951 730 -2951 0 3
rlabel polysilicon 733 -2951 733 -2951 0 4
rlabel polysilicon 737 -2945 737 -2945 0 1
rlabel polysilicon 737 -2951 737 -2951 0 3
rlabel polysilicon 744 -2945 744 -2945 0 1
rlabel polysilicon 744 -2951 744 -2951 0 3
rlabel polysilicon 751 -2945 751 -2945 0 1
rlabel polysilicon 751 -2951 751 -2951 0 3
rlabel polysilicon 761 -2945 761 -2945 0 2
rlabel polysilicon 758 -2951 758 -2951 0 3
rlabel polysilicon 761 -2951 761 -2951 0 4
rlabel polysilicon 765 -2945 765 -2945 0 1
rlabel polysilicon 765 -2951 765 -2951 0 3
rlabel polysilicon 772 -2945 772 -2945 0 1
rlabel polysilicon 772 -2951 772 -2951 0 3
rlabel polysilicon 779 -2945 779 -2945 0 1
rlabel polysilicon 779 -2951 779 -2951 0 3
rlabel polysilicon 786 -2945 786 -2945 0 1
rlabel polysilicon 786 -2951 786 -2951 0 3
rlabel polysilicon 793 -2945 793 -2945 0 1
rlabel polysilicon 793 -2951 793 -2951 0 3
rlabel polysilicon 800 -2945 800 -2945 0 1
rlabel polysilicon 800 -2951 800 -2951 0 3
rlabel polysilicon 807 -2945 807 -2945 0 1
rlabel polysilicon 807 -2951 807 -2951 0 3
rlabel polysilicon 814 -2945 814 -2945 0 1
rlabel polysilicon 814 -2951 814 -2951 0 3
rlabel polysilicon 821 -2945 821 -2945 0 1
rlabel polysilicon 821 -2951 821 -2951 0 3
rlabel polysilicon 828 -2945 828 -2945 0 1
rlabel polysilicon 828 -2951 828 -2951 0 3
rlabel polysilicon 835 -2945 835 -2945 0 1
rlabel polysilicon 835 -2951 835 -2951 0 3
rlabel polysilicon 842 -2945 842 -2945 0 1
rlabel polysilicon 842 -2951 842 -2951 0 3
rlabel polysilicon 849 -2945 849 -2945 0 1
rlabel polysilicon 849 -2951 849 -2951 0 3
rlabel polysilicon 856 -2945 856 -2945 0 1
rlabel polysilicon 856 -2951 856 -2951 0 3
rlabel polysilicon 863 -2945 863 -2945 0 1
rlabel polysilicon 866 -2945 866 -2945 0 2
rlabel polysilicon 863 -2951 863 -2951 0 3
rlabel polysilicon 866 -2951 866 -2951 0 4
rlabel polysilicon 870 -2945 870 -2945 0 1
rlabel polysilicon 870 -2951 870 -2951 0 3
rlabel polysilicon 877 -2945 877 -2945 0 1
rlabel polysilicon 877 -2951 877 -2951 0 3
rlabel polysilicon 884 -2945 884 -2945 0 1
rlabel polysilicon 884 -2951 884 -2951 0 3
rlabel polysilicon 891 -2945 891 -2945 0 1
rlabel polysilicon 891 -2951 891 -2951 0 3
rlabel polysilicon 898 -2945 898 -2945 0 1
rlabel polysilicon 898 -2951 898 -2951 0 3
rlabel polysilicon 905 -2945 905 -2945 0 1
rlabel polysilicon 905 -2951 905 -2951 0 3
rlabel polysilicon 912 -2945 912 -2945 0 1
rlabel polysilicon 915 -2945 915 -2945 0 2
rlabel polysilicon 912 -2951 912 -2951 0 3
rlabel polysilicon 919 -2945 919 -2945 0 1
rlabel polysilicon 919 -2951 919 -2951 0 3
rlabel polysilicon 926 -2945 926 -2945 0 1
rlabel polysilicon 929 -2945 929 -2945 0 2
rlabel polysilicon 926 -2951 926 -2951 0 3
rlabel polysilicon 929 -2951 929 -2951 0 4
rlabel polysilicon 936 -2945 936 -2945 0 2
rlabel polysilicon 933 -2951 933 -2951 0 3
rlabel polysilicon 936 -2951 936 -2951 0 4
rlabel polysilicon 940 -2945 940 -2945 0 1
rlabel polysilicon 940 -2951 940 -2951 0 3
rlabel polysilicon 947 -2945 947 -2945 0 1
rlabel polysilicon 947 -2951 947 -2951 0 3
rlabel polysilicon 954 -2945 954 -2945 0 1
rlabel polysilicon 954 -2951 954 -2951 0 3
rlabel polysilicon 961 -2945 961 -2945 0 1
rlabel polysilicon 961 -2951 961 -2951 0 3
rlabel polysilicon 968 -2945 968 -2945 0 1
rlabel polysilicon 968 -2951 968 -2951 0 3
rlabel polysilicon 975 -2945 975 -2945 0 1
rlabel polysilicon 975 -2951 975 -2951 0 3
rlabel polysilicon 982 -2945 982 -2945 0 1
rlabel polysilicon 982 -2951 982 -2951 0 3
rlabel polysilicon 989 -2945 989 -2945 0 1
rlabel polysilicon 989 -2951 989 -2951 0 3
rlabel polysilicon 996 -2945 996 -2945 0 1
rlabel polysilicon 996 -2951 996 -2951 0 3
rlabel polysilicon 999 -2951 999 -2951 0 4
rlabel polysilicon 1003 -2945 1003 -2945 0 1
rlabel polysilicon 1003 -2951 1003 -2951 0 3
rlabel polysilicon 1010 -2945 1010 -2945 0 1
rlabel polysilicon 1010 -2951 1010 -2951 0 3
rlabel polysilicon 1017 -2945 1017 -2945 0 1
rlabel polysilicon 1017 -2951 1017 -2951 0 3
rlabel polysilicon 1020 -2951 1020 -2951 0 4
rlabel polysilicon 1024 -2945 1024 -2945 0 1
rlabel polysilicon 1027 -2945 1027 -2945 0 2
rlabel polysilicon 1024 -2951 1024 -2951 0 3
rlabel polysilicon 1031 -2945 1031 -2945 0 1
rlabel polysilicon 1031 -2951 1031 -2951 0 3
rlabel polysilicon 1038 -2945 1038 -2945 0 1
rlabel polysilicon 1038 -2951 1038 -2951 0 3
rlabel polysilicon 1045 -2945 1045 -2945 0 1
rlabel polysilicon 1045 -2951 1045 -2951 0 3
rlabel polysilicon 1052 -2945 1052 -2945 0 1
rlabel polysilicon 1052 -2951 1052 -2951 0 3
rlabel polysilicon 1059 -2945 1059 -2945 0 1
rlabel polysilicon 1059 -2951 1059 -2951 0 3
rlabel polysilicon 1066 -2945 1066 -2945 0 1
rlabel polysilicon 1066 -2951 1066 -2951 0 3
rlabel polysilicon 1073 -2945 1073 -2945 0 1
rlabel polysilicon 1073 -2951 1073 -2951 0 3
rlabel polysilicon 1080 -2945 1080 -2945 0 1
rlabel polysilicon 1080 -2951 1080 -2951 0 3
rlabel polysilicon 1087 -2945 1087 -2945 0 1
rlabel polysilicon 1087 -2951 1087 -2951 0 3
rlabel polysilicon 1094 -2945 1094 -2945 0 1
rlabel polysilicon 1094 -2951 1094 -2951 0 3
rlabel polysilicon 1101 -2945 1101 -2945 0 1
rlabel polysilicon 1101 -2951 1101 -2951 0 3
rlabel polysilicon 1108 -2945 1108 -2945 0 1
rlabel polysilicon 1108 -2951 1108 -2951 0 3
rlabel polysilicon 1115 -2945 1115 -2945 0 1
rlabel polysilicon 1115 -2951 1115 -2951 0 3
rlabel polysilicon 1122 -2945 1122 -2945 0 1
rlabel polysilicon 1122 -2951 1122 -2951 0 3
rlabel polysilicon 1129 -2945 1129 -2945 0 1
rlabel polysilicon 1129 -2951 1129 -2951 0 3
rlabel polysilicon 1136 -2945 1136 -2945 0 1
rlabel polysilicon 1136 -2951 1136 -2951 0 3
rlabel polysilicon 1143 -2945 1143 -2945 0 1
rlabel polysilicon 1143 -2951 1143 -2951 0 3
rlabel polysilicon 1150 -2945 1150 -2945 0 1
rlabel polysilicon 1150 -2951 1150 -2951 0 3
rlabel polysilicon 1157 -2945 1157 -2945 0 1
rlabel polysilicon 1157 -2951 1157 -2951 0 3
rlabel polysilicon 1164 -2945 1164 -2945 0 1
rlabel polysilicon 1164 -2951 1164 -2951 0 3
rlabel polysilicon 1171 -2945 1171 -2945 0 1
rlabel polysilicon 1171 -2951 1171 -2951 0 3
rlabel polysilicon 1178 -2945 1178 -2945 0 1
rlabel polysilicon 1178 -2951 1178 -2951 0 3
rlabel polysilicon 1185 -2945 1185 -2945 0 1
rlabel polysilicon 1185 -2951 1185 -2951 0 3
rlabel polysilicon 1192 -2945 1192 -2945 0 1
rlabel polysilicon 1192 -2951 1192 -2951 0 3
rlabel polysilicon 1199 -2945 1199 -2945 0 1
rlabel polysilicon 1202 -2945 1202 -2945 0 2
rlabel polysilicon 1206 -2945 1206 -2945 0 1
rlabel polysilicon 1206 -2951 1206 -2951 0 3
rlabel polysilicon 1213 -2945 1213 -2945 0 1
rlabel polysilicon 1213 -2951 1213 -2951 0 3
rlabel polysilicon 1220 -2945 1220 -2945 0 1
rlabel polysilicon 1220 -2951 1220 -2951 0 3
rlabel polysilicon 1227 -2945 1227 -2945 0 1
rlabel polysilicon 1227 -2951 1227 -2951 0 3
rlabel polysilicon 1234 -2945 1234 -2945 0 1
rlabel polysilicon 1234 -2951 1234 -2951 0 3
rlabel polysilicon 1241 -2945 1241 -2945 0 1
rlabel polysilicon 1241 -2951 1241 -2951 0 3
rlabel polysilicon 1248 -2945 1248 -2945 0 1
rlabel polysilicon 1248 -2951 1248 -2951 0 3
rlabel polysilicon 1255 -2945 1255 -2945 0 1
rlabel polysilicon 1255 -2951 1255 -2951 0 3
rlabel polysilicon 1262 -2945 1262 -2945 0 1
rlabel polysilicon 1262 -2951 1262 -2951 0 3
rlabel polysilicon 1269 -2945 1269 -2945 0 1
rlabel polysilicon 1269 -2951 1269 -2951 0 3
rlabel polysilicon 1276 -2945 1276 -2945 0 1
rlabel polysilicon 1276 -2951 1276 -2951 0 3
rlabel polysilicon 1283 -2945 1283 -2945 0 1
rlabel polysilicon 1283 -2951 1283 -2951 0 3
rlabel polysilicon 1290 -2945 1290 -2945 0 1
rlabel polysilicon 1290 -2951 1290 -2951 0 3
rlabel polysilicon 1297 -2945 1297 -2945 0 1
rlabel polysilicon 1297 -2951 1297 -2951 0 3
rlabel polysilicon 1304 -2945 1304 -2945 0 1
rlabel polysilicon 1304 -2951 1304 -2951 0 3
rlabel polysilicon 1311 -2945 1311 -2945 0 1
rlabel polysilicon 1311 -2951 1311 -2951 0 3
rlabel polysilicon 1318 -2945 1318 -2945 0 1
rlabel polysilicon 1318 -2951 1318 -2951 0 3
rlabel polysilicon 1325 -2945 1325 -2945 0 1
rlabel polysilicon 1325 -2951 1325 -2951 0 3
rlabel polysilicon 1332 -2945 1332 -2945 0 1
rlabel polysilicon 1332 -2951 1332 -2951 0 3
rlabel polysilicon 1339 -2945 1339 -2945 0 1
rlabel polysilicon 1339 -2951 1339 -2951 0 3
rlabel polysilicon 1346 -2945 1346 -2945 0 1
rlabel polysilicon 1346 -2951 1346 -2951 0 3
rlabel polysilicon 1353 -2945 1353 -2945 0 1
rlabel polysilicon 1353 -2951 1353 -2951 0 3
rlabel polysilicon 1360 -2945 1360 -2945 0 1
rlabel polysilicon 1360 -2951 1360 -2951 0 3
rlabel polysilicon 1367 -2945 1367 -2945 0 1
rlabel polysilicon 1367 -2951 1367 -2951 0 3
rlabel polysilicon 1374 -2945 1374 -2945 0 1
rlabel polysilicon 1374 -2951 1374 -2951 0 3
rlabel polysilicon 1381 -2945 1381 -2945 0 1
rlabel polysilicon 1381 -2951 1381 -2951 0 3
rlabel polysilicon 1388 -2945 1388 -2945 0 1
rlabel polysilicon 1388 -2951 1388 -2951 0 3
rlabel polysilicon 1395 -2945 1395 -2945 0 1
rlabel polysilicon 1395 -2951 1395 -2951 0 3
rlabel polysilicon 1402 -2945 1402 -2945 0 1
rlabel polysilicon 1402 -2951 1402 -2951 0 3
rlabel polysilicon 1409 -2945 1409 -2945 0 1
rlabel polysilicon 1409 -2951 1409 -2951 0 3
rlabel polysilicon 1416 -2945 1416 -2945 0 1
rlabel polysilicon 1416 -2951 1416 -2951 0 3
rlabel polysilicon 1423 -2945 1423 -2945 0 1
rlabel polysilicon 1423 -2951 1423 -2951 0 3
rlabel polysilicon 1430 -2945 1430 -2945 0 1
rlabel polysilicon 1430 -2951 1430 -2951 0 3
rlabel polysilicon 1437 -2945 1437 -2945 0 1
rlabel polysilicon 1437 -2951 1437 -2951 0 3
rlabel polysilicon 1447 -2945 1447 -2945 0 2
rlabel polysilicon 1444 -2951 1444 -2951 0 3
rlabel polysilicon 1447 -2951 1447 -2951 0 4
rlabel polysilicon 1451 -2945 1451 -2945 0 1
rlabel polysilicon 1451 -2951 1451 -2951 0 3
rlabel polysilicon 1458 -2945 1458 -2945 0 1
rlabel polysilicon 1458 -2951 1458 -2951 0 3
rlabel polysilicon 1465 -2945 1465 -2945 0 1
rlabel polysilicon 1465 -2951 1465 -2951 0 3
rlabel polysilicon 1479 -2945 1479 -2945 0 1
rlabel polysilicon 1479 -2951 1479 -2951 0 3
rlabel polysilicon 1486 -2945 1486 -2945 0 1
rlabel polysilicon 1486 -2951 1486 -2951 0 3
rlabel polysilicon 1493 -2945 1493 -2945 0 1
rlabel polysilicon 1493 -2951 1493 -2951 0 3
rlabel polysilicon 1500 -2945 1500 -2945 0 1
rlabel polysilicon 1500 -2951 1500 -2951 0 3
rlabel polysilicon 37 -3064 37 -3064 0 1
rlabel polysilicon 37 -3070 37 -3070 0 3
rlabel polysilicon 44 -3064 44 -3064 0 1
rlabel polysilicon 44 -3070 44 -3070 0 3
rlabel polysilicon 51 -3064 51 -3064 0 1
rlabel polysilicon 51 -3070 51 -3070 0 3
rlabel polysilicon 58 -3064 58 -3064 0 1
rlabel polysilicon 58 -3070 58 -3070 0 3
rlabel polysilicon 65 -3064 65 -3064 0 1
rlabel polysilicon 65 -3070 65 -3070 0 3
rlabel polysilicon 72 -3064 72 -3064 0 1
rlabel polysilicon 72 -3070 72 -3070 0 3
rlabel polysilicon 79 -3064 79 -3064 0 1
rlabel polysilicon 79 -3070 79 -3070 0 3
rlabel polysilicon 86 -3064 86 -3064 0 1
rlabel polysilicon 86 -3070 86 -3070 0 3
rlabel polysilicon 96 -3064 96 -3064 0 2
rlabel polysilicon 93 -3070 93 -3070 0 3
rlabel polysilicon 96 -3070 96 -3070 0 4
rlabel polysilicon 100 -3064 100 -3064 0 1
rlabel polysilicon 100 -3070 100 -3070 0 3
rlabel polysilicon 107 -3064 107 -3064 0 1
rlabel polysilicon 107 -3070 107 -3070 0 3
rlabel polysilicon 114 -3064 114 -3064 0 1
rlabel polysilicon 114 -3070 114 -3070 0 3
rlabel polysilicon 121 -3064 121 -3064 0 1
rlabel polysilicon 124 -3064 124 -3064 0 2
rlabel polysilicon 121 -3070 121 -3070 0 3
rlabel polysilicon 128 -3064 128 -3064 0 1
rlabel polysilicon 128 -3070 128 -3070 0 3
rlabel polysilicon 135 -3064 135 -3064 0 1
rlabel polysilicon 135 -3070 135 -3070 0 3
rlabel polysilicon 142 -3064 142 -3064 0 1
rlabel polysilicon 142 -3070 142 -3070 0 3
rlabel polysilicon 149 -3064 149 -3064 0 1
rlabel polysilicon 149 -3070 149 -3070 0 3
rlabel polysilicon 156 -3064 156 -3064 0 1
rlabel polysilicon 156 -3070 156 -3070 0 3
rlabel polysilicon 163 -3064 163 -3064 0 1
rlabel polysilicon 163 -3070 163 -3070 0 3
rlabel polysilicon 170 -3064 170 -3064 0 1
rlabel polysilicon 170 -3070 170 -3070 0 3
rlabel polysilicon 177 -3064 177 -3064 0 1
rlabel polysilicon 177 -3070 177 -3070 0 3
rlabel polysilicon 180 -3070 180 -3070 0 4
rlabel polysilicon 184 -3064 184 -3064 0 1
rlabel polysilicon 184 -3070 184 -3070 0 3
rlabel polysilicon 191 -3064 191 -3064 0 1
rlabel polysilicon 191 -3070 191 -3070 0 3
rlabel polysilicon 201 -3064 201 -3064 0 2
rlabel polysilicon 198 -3070 198 -3070 0 3
rlabel polysilicon 201 -3070 201 -3070 0 4
rlabel polysilicon 205 -3064 205 -3064 0 1
rlabel polysilicon 205 -3070 205 -3070 0 3
rlabel polysilicon 212 -3064 212 -3064 0 1
rlabel polysilicon 212 -3070 212 -3070 0 3
rlabel polysilicon 222 -3070 222 -3070 0 4
rlabel polysilicon 226 -3064 226 -3064 0 1
rlabel polysilicon 226 -3070 226 -3070 0 3
rlabel polysilicon 233 -3064 233 -3064 0 1
rlabel polysilicon 233 -3070 233 -3070 0 3
rlabel polysilicon 243 -3064 243 -3064 0 2
rlabel polysilicon 240 -3070 240 -3070 0 3
rlabel polysilicon 243 -3070 243 -3070 0 4
rlabel polysilicon 247 -3064 247 -3064 0 1
rlabel polysilicon 250 -3064 250 -3064 0 2
rlabel polysilicon 247 -3070 247 -3070 0 3
rlabel polysilicon 250 -3070 250 -3070 0 4
rlabel polysilicon 254 -3064 254 -3064 0 1
rlabel polysilicon 254 -3070 254 -3070 0 3
rlabel polysilicon 261 -3064 261 -3064 0 1
rlabel polysilicon 264 -3064 264 -3064 0 2
rlabel polysilicon 261 -3070 261 -3070 0 3
rlabel polysilicon 268 -3064 268 -3064 0 1
rlabel polysilicon 268 -3070 268 -3070 0 3
rlabel polysilicon 275 -3064 275 -3064 0 1
rlabel polysilicon 275 -3070 275 -3070 0 3
rlabel polysilicon 282 -3064 282 -3064 0 1
rlabel polysilicon 282 -3070 282 -3070 0 3
rlabel polysilicon 289 -3064 289 -3064 0 1
rlabel polysilicon 289 -3070 289 -3070 0 3
rlabel polysilicon 296 -3064 296 -3064 0 1
rlabel polysilicon 296 -3070 296 -3070 0 3
rlabel polysilicon 299 -3070 299 -3070 0 4
rlabel polysilicon 303 -3064 303 -3064 0 1
rlabel polysilicon 303 -3070 303 -3070 0 3
rlabel polysilicon 310 -3064 310 -3064 0 1
rlabel polysilicon 310 -3070 310 -3070 0 3
rlabel polysilicon 317 -3064 317 -3064 0 1
rlabel polysilicon 317 -3070 317 -3070 0 3
rlabel polysilicon 324 -3064 324 -3064 0 1
rlabel polysilicon 324 -3070 324 -3070 0 3
rlabel polysilicon 331 -3064 331 -3064 0 1
rlabel polysilicon 331 -3070 331 -3070 0 3
rlabel polysilicon 338 -3064 338 -3064 0 1
rlabel polysilicon 338 -3070 338 -3070 0 3
rlabel polysilicon 345 -3064 345 -3064 0 1
rlabel polysilicon 345 -3070 345 -3070 0 3
rlabel polysilicon 352 -3064 352 -3064 0 1
rlabel polysilicon 355 -3064 355 -3064 0 2
rlabel polysilicon 352 -3070 352 -3070 0 3
rlabel polysilicon 355 -3070 355 -3070 0 4
rlabel polysilicon 359 -3064 359 -3064 0 1
rlabel polysilicon 359 -3070 359 -3070 0 3
rlabel polysilicon 366 -3064 366 -3064 0 1
rlabel polysilicon 366 -3070 366 -3070 0 3
rlabel polysilicon 373 -3064 373 -3064 0 1
rlabel polysilicon 373 -3070 373 -3070 0 3
rlabel polysilicon 380 -3064 380 -3064 0 1
rlabel polysilicon 380 -3070 380 -3070 0 3
rlabel polysilicon 387 -3064 387 -3064 0 1
rlabel polysilicon 387 -3070 387 -3070 0 3
rlabel polysilicon 394 -3064 394 -3064 0 1
rlabel polysilicon 394 -3070 394 -3070 0 3
rlabel polysilicon 401 -3064 401 -3064 0 1
rlabel polysilicon 401 -3070 401 -3070 0 3
rlabel polysilicon 408 -3064 408 -3064 0 1
rlabel polysilicon 411 -3064 411 -3064 0 2
rlabel polysilicon 408 -3070 408 -3070 0 3
rlabel polysilicon 415 -3064 415 -3064 0 1
rlabel polysilicon 415 -3070 415 -3070 0 3
rlabel polysilicon 422 -3064 422 -3064 0 1
rlabel polysilicon 422 -3070 422 -3070 0 3
rlabel polysilicon 429 -3064 429 -3064 0 1
rlabel polysilicon 429 -3070 429 -3070 0 3
rlabel polysilicon 436 -3064 436 -3064 0 1
rlabel polysilicon 436 -3070 436 -3070 0 3
rlabel polysilicon 443 -3064 443 -3064 0 1
rlabel polysilicon 443 -3070 443 -3070 0 3
rlabel polysilicon 450 -3064 450 -3064 0 1
rlabel polysilicon 450 -3070 450 -3070 0 3
rlabel polysilicon 457 -3064 457 -3064 0 1
rlabel polysilicon 457 -3070 457 -3070 0 3
rlabel polysilicon 464 -3064 464 -3064 0 1
rlabel polysilicon 464 -3070 464 -3070 0 3
rlabel polysilicon 471 -3064 471 -3064 0 1
rlabel polysilicon 471 -3070 471 -3070 0 3
rlabel polysilicon 478 -3064 478 -3064 0 1
rlabel polysilicon 478 -3070 478 -3070 0 3
rlabel polysilicon 485 -3064 485 -3064 0 1
rlabel polysilicon 485 -3070 485 -3070 0 3
rlabel polysilicon 492 -3064 492 -3064 0 1
rlabel polysilicon 492 -3070 492 -3070 0 3
rlabel polysilicon 499 -3064 499 -3064 0 1
rlabel polysilicon 499 -3070 499 -3070 0 3
rlabel polysilicon 506 -3064 506 -3064 0 1
rlabel polysilicon 506 -3070 506 -3070 0 3
rlabel polysilicon 513 -3064 513 -3064 0 1
rlabel polysilicon 513 -3070 513 -3070 0 3
rlabel polysilicon 520 -3064 520 -3064 0 1
rlabel polysilicon 523 -3064 523 -3064 0 2
rlabel polysilicon 520 -3070 520 -3070 0 3
rlabel polysilicon 523 -3070 523 -3070 0 4
rlabel polysilicon 527 -3064 527 -3064 0 1
rlabel polysilicon 527 -3070 527 -3070 0 3
rlabel polysilicon 534 -3064 534 -3064 0 1
rlabel polysilicon 534 -3070 534 -3070 0 3
rlabel polysilicon 541 -3064 541 -3064 0 1
rlabel polysilicon 541 -3070 541 -3070 0 3
rlabel polysilicon 548 -3064 548 -3064 0 1
rlabel polysilicon 548 -3070 548 -3070 0 3
rlabel polysilicon 555 -3064 555 -3064 0 1
rlabel polysilicon 555 -3070 555 -3070 0 3
rlabel polysilicon 562 -3064 562 -3064 0 1
rlabel polysilicon 562 -3070 562 -3070 0 3
rlabel polysilicon 569 -3064 569 -3064 0 1
rlabel polysilicon 569 -3070 569 -3070 0 3
rlabel polysilicon 576 -3064 576 -3064 0 1
rlabel polysilicon 576 -3070 576 -3070 0 3
rlabel polysilicon 583 -3064 583 -3064 0 1
rlabel polysilicon 583 -3070 583 -3070 0 3
rlabel polysilicon 590 -3064 590 -3064 0 1
rlabel polysilicon 590 -3070 590 -3070 0 3
rlabel polysilicon 597 -3064 597 -3064 0 1
rlabel polysilicon 597 -3070 597 -3070 0 3
rlabel polysilicon 604 -3064 604 -3064 0 1
rlabel polysilicon 607 -3064 607 -3064 0 2
rlabel polysilicon 604 -3070 604 -3070 0 3
rlabel polysilicon 611 -3064 611 -3064 0 1
rlabel polysilicon 611 -3070 611 -3070 0 3
rlabel polysilicon 618 -3064 618 -3064 0 1
rlabel polysilicon 621 -3064 621 -3064 0 2
rlabel polysilicon 618 -3070 618 -3070 0 3
rlabel polysilicon 621 -3070 621 -3070 0 4
rlabel polysilicon 625 -3064 625 -3064 0 1
rlabel polysilicon 625 -3070 625 -3070 0 3
rlabel polysilicon 632 -3064 632 -3064 0 1
rlabel polysilicon 632 -3070 632 -3070 0 3
rlabel polysilicon 639 -3064 639 -3064 0 1
rlabel polysilicon 642 -3064 642 -3064 0 2
rlabel polysilicon 642 -3070 642 -3070 0 4
rlabel polysilicon 646 -3064 646 -3064 0 1
rlabel polysilicon 646 -3070 646 -3070 0 3
rlabel polysilicon 653 -3064 653 -3064 0 1
rlabel polysilicon 653 -3070 653 -3070 0 3
rlabel polysilicon 660 -3064 660 -3064 0 1
rlabel polysilicon 660 -3070 660 -3070 0 3
rlabel polysilicon 667 -3064 667 -3064 0 1
rlabel polysilicon 667 -3070 667 -3070 0 3
rlabel polysilicon 674 -3064 674 -3064 0 1
rlabel polysilicon 674 -3070 674 -3070 0 3
rlabel polysilicon 681 -3064 681 -3064 0 1
rlabel polysilicon 684 -3064 684 -3064 0 2
rlabel polysilicon 681 -3070 681 -3070 0 3
rlabel polysilicon 684 -3070 684 -3070 0 4
rlabel polysilicon 688 -3064 688 -3064 0 1
rlabel polysilicon 688 -3070 688 -3070 0 3
rlabel polysilicon 695 -3064 695 -3064 0 1
rlabel polysilicon 695 -3070 695 -3070 0 3
rlabel polysilicon 702 -3064 702 -3064 0 1
rlabel polysilicon 705 -3064 705 -3064 0 2
rlabel polysilicon 702 -3070 702 -3070 0 3
rlabel polysilicon 705 -3070 705 -3070 0 4
rlabel polysilicon 709 -3064 709 -3064 0 1
rlabel polysilicon 709 -3070 709 -3070 0 3
rlabel polysilicon 716 -3064 716 -3064 0 1
rlabel polysilicon 716 -3070 716 -3070 0 3
rlabel polysilicon 723 -3064 723 -3064 0 1
rlabel polysilicon 723 -3070 723 -3070 0 3
rlabel polysilicon 730 -3064 730 -3064 0 1
rlabel polysilicon 730 -3070 730 -3070 0 3
rlabel polysilicon 740 -3064 740 -3064 0 2
rlabel polysilicon 737 -3070 737 -3070 0 3
rlabel polysilicon 740 -3070 740 -3070 0 4
rlabel polysilicon 744 -3064 744 -3064 0 1
rlabel polysilicon 744 -3070 744 -3070 0 3
rlabel polysilicon 751 -3064 751 -3064 0 1
rlabel polysilicon 751 -3070 751 -3070 0 3
rlabel polysilicon 758 -3064 758 -3064 0 1
rlabel polysilicon 758 -3070 758 -3070 0 3
rlabel polysilicon 765 -3064 765 -3064 0 1
rlabel polysilicon 765 -3070 765 -3070 0 3
rlabel polysilicon 772 -3064 772 -3064 0 1
rlabel polysilicon 772 -3070 772 -3070 0 3
rlabel polysilicon 779 -3064 779 -3064 0 1
rlabel polysilicon 779 -3070 779 -3070 0 3
rlabel polysilicon 786 -3064 786 -3064 0 1
rlabel polysilicon 786 -3070 786 -3070 0 3
rlabel polysilicon 796 -3064 796 -3064 0 2
rlabel polysilicon 793 -3070 793 -3070 0 3
rlabel polysilicon 796 -3070 796 -3070 0 4
rlabel polysilicon 800 -3064 800 -3064 0 1
rlabel polysilicon 800 -3070 800 -3070 0 3
rlabel polysilicon 807 -3064 807 -3064 0 1
rlabel polysilicon 807 -3070 807 -3070 0 3
rlabel polysilicon 814 -3064 814 -3064 0 1
rlabel polysilicon 814 -3070 814 -3070 0 3
rlabel polysilicon 821 -3064 821 -3064 0 1
rlabel polysilicon 821 -3070 821 -3070 0 3
rlabel polysilicon 828 -3064 828 -3064 0 1
rlabel polysilicon 828 -3070 828 -3070 0 3
rlabel polysilicon 835 -3064 835 -3064 0 1
rlabel polysilicon 835 -3070 835 -3070 0 3
rlabel polysilicon 842 -3064 842 -3064 0 1
rlabel polysilicon 842 -3070 842 -3070 0 3
rlabel polysilicon 849 -3064 849 -3064 0 1
rlabel polysilicon 852 -3064 852 -3064 0 2
rlabel polysilicon 849 -3070 849 -3070 0 3
rlabel polysilicon 856 -3064 856 -3064 0 1
rlabel polysilicon 856 -3070 856 -3070 0 3
rlabel polysilicon 863 -3064 863 -3064 0 1
rlabel polysilicon 863 -3070 863 -3070 0 3
rlabel polysilicon 870 -3064 870 -3064 0 1
rlabel polysilicon 873 -3064 873 -3064 0 2
rlabel polysilicon 870 -3070 870 -3070 0 3
rlabel polysilicon 873 -3070 873 -3070 0 4
rlabel polysilicon 877 -3064 877 -3064 0 1
rlabel polysilicon 877 -3070 877 -3070 0 3
rlabel polysilicon 884 -3064 884 -3064 0 1
rlabel polysilicon 884 -3070 884 -3070 0 3
rlabel polysilicon 891 -3064 891 -3064 0 1
rlabel polysilicon 891 -3070 891 -3070 0 3
rlabel polysilicon 898 -3064 898 -3064 0 1
rlabel polysilicon 898 -3070 898 -3070 0 3
rlabel polysilicon 905 -3064 905 -3064 0 1
rlabel polysilicon 905 -3070 905 -3070 0 3
rlabel polysilicon 912 -3064 912 -3064 0 1
rlabel polysilicon 912 -3070 912 -3070 0 3
rlabel polysilicon 919 -3064 919 -3064 0 1
rlabel polysilicon 922 -3064 922 -3064 0 2
rlabel polysilicon 919 -3070 919 -3070 0 3
rlabel polysilicon 926 -3064 926 -3064 0 1
rlabel polysilicon 926 -3070 926 -3070 0 3
rlabel polysilicon 929 -3070 929 -3070 0 4
rlabel polysilicon 933 -3064 933 -3064 0 1
rlabel polysilicon 933 -3070 933 -3070 0 3
rlabel polysilicon 940 -3064 940 -3064 0 1
rlabel polysilicon 940 -3070 940 -3070 0 3
rlabel polysilicon 947 -3064 947 -3064 0 1
rlabel polysilicon 947 -3070 947 -3070 0 3
rlabel polysilicon 954 -3064 954 -3064 0 1
rlabel polysilicon 954 -3070 954 -3070 0 3
rlabel polysilicon 961 -3064 961 -3064 0 1
rlabel polysilicon 961 -3070 961 -3070 0 3
rlabel polysilicon 964 -3070 964 -3070 0 4
rlabel polysilicon 968 -3064 968 -3064 0 1
rlabel polysilicon 968 -3070 968 -3070 0 3
rlabel polysilicon 975 -3064 975 -3064 0 1
rlabel polysilicon 975 -3070 975 -3070 0 3
rlabel polysilicon 982 -3064 982 -3064 0 1
rlabel polysilicon 982 -3070 982 -3070 0 3
rlabel polysilicon 989 -3064 989 -3064 0 1
rlabel polysilicon 989 -3070 989 -3070 0 3
rlabel polysilicon 996 -3064 996 -3064 0 1
rlabel polysilicon 999 -3064 999 -3064 0 2
rlabel polysilicon 996 -3070 996 -3070 0 3
rlabel polysilicon 1003 -3064 1003 -3064 0 1
rlabel polysilicon 1003 -3070 1003 -3070 0 3
rlabel polysilicon 1010 -3064 1010 -3064 0 1
rlabel polysilicon 1010 -3070 1010 -3070 0 3
rlabel polysilicon 1017 -3064 1017 -3064 0 1
rlabel polysilicon 1017 -3070 1017 -3070 0 3
rlabel polysilicon 1024 -3064 1024 -3064 0 1
rlabel polysilicon 1024 -3070 1024 -3070 0 3
rlabel polysilicon 1031 -3064 1031 -3064 0 1
rlabel polysilicon 1031 -3070 1031 -3070 0 3
rlabel polysilicon 1038 -3064 1038 -3064 0 1
rlabel polysilicon 1038 -3070 1038 -3070 0 3
rlabel polysilicon 1045 -3064 1045 -3064 0 1
rlabel polysilicon 1045 -3070 1045 -3070 0 3
rlabel polysilicon 1052 -3064 1052 -3064 0 1
rlabel polysilicon 1052 -3070 1052 -3070 0 3
rlabel polysilicon 1062 -3064 1062 -3064 0 2
rlabel polysilicon 1062 -3070 1062 -3070 0 4
rlabel polysilicon 1066 -3064 1066 -3064 0 1
rlabel polysilicon 1066 -3070 1066 -3070 0 3
rlabel polysilicon 1073 -3064 1073 -3064 0 1
rlabel polysilicon 1073 -3070 1073 -3070 0 3
rlabel polysilicon 1080 -3064 1080 -3064 0 1
rlabel polysilicon 1080 -3070 1080 -3070 0 3
rlabel polysilicon 1087 -3064 1087 -3064 0 1
rlabel polysilicon 1090 -3064 1090 -3064 0 2
rlabel polysilicon 1087 -3070 1087 -3070 0 3
rlabel polysilicon 1094 -3064 1094 -3064 0 1
rlabel polysilicon 1094 -3070 1094 -3070 0 3
rlabel polysilicon 1101 -3064 1101 -3064 0 1
rlabel polysilicon 1101 -3070 1101 -3070 0 3
rlabel polysilicon 1108 -3064 1108 -3064 0 1
rlabel polysilicon 1108 -3070 1108 -3070 0 3
rlabel polysilicon 1115 -3064 1115 -3064 0 1
rlabel polysilicon 1115 -3070 1115 -3070 0 3
rlabel polysilicon 1122 -3064 1122 -3064 0 1
rlabel polysilicon 1122 -3070 1122 -3070 0 3
rlabel polysilicon 1129 -3064 1129 -3064 0 1
rlabel polysilicon 1129 -3070 1129 -3070 0 3
rlabel polysilicon 1136 -3064 1136 -3064 0 1
rlabel polysilicon 1136 -3070 1136 -3070 0 3
rlabel polysilicon 1143 -3064 1143 -3064 0 1
rlabel polysilicon 1143 -3070 1143 -3070 0 3
rlabel polysilicon 1150 -3064 1150 -3064 0 1
rlabel polysilicon 1150 -3070 1150 -3070 0 3
rlabel polysilicon 1157 -3064 1157 -3064 0 1
rlabel polysilicon 1157 -3070 1157 -3070 0 3
rlabel polysilicon 1164 -3064 1164 -3064 0 1
rlabel polysilicon 1164 -3070 1164 -3070 0 3
rlabel polysilicon 1171 -3064 1171 -3064 0 1
rlabel polysilicon 1171 -3070 1171 -3070 0 3
rlabel polysilicon 1178 -3064 1178 -3064 0 1
rlabel polysilicon 1178 -3070 1178 -3070 0 3
rlabel polysilicon 1185 -3064 1185 -3064 0 1
rlabel polysilicon 1185 -3070 1185 -3070 0 3
rlabel polysilicon 1192 -3064 1192 -3064 0 1
rlabel polysilicon 1192 -3070 1192 -3070 0 3
rlabel polysilicon 1199 -3064 1199 -3064 0 1
rlabel polysilicon 1199 -3070 1199 -3070 0 3
rlabel polysilicon 1206 -3064 1206 -3064 0 1
rlabel polysilicon 1206 -3070 1206 -3070 0 3
rlabel polysilicon 1213 -3064 1213 -3064 0 1
rlabel polysilicon 1213 -3070 1213 -3070 0 3
rlabel polysilicon 1220 -3064 1220 -3064 0 1
rlabel polysilicon 1223 -3064 1223 -3064 0 2
rlabel polysilicon 1220 -3070 1220 -3070 0 3
rlabel polysilicon 1223 -3070 1223 -3070 0 4
rlabel polysilicon 1227 -3064 1227 -3064 0 1
rlabel polysilicon 1227 -3070 1227 -3070 0 3
rlabel polysilicon 1234 -3064 1234 -3064 0 1
rlabel polysilicon 1234 -3070 1234 -3070 0 3
rlabel polysilicon 1241 -3064 1241 -3064 0 1
rlabel polysilicon 1241 -3070 1241 -3070 0 3
rlabel polysilicon 1248 -3064 1248 -3064 0 1
rlabel polysilicon 1248 -3070 1248 -3070 0 3
rlabel polysilicon 1255 -3064 1255 -3064 0 1
rlabel polysilicon 1255 -3070 1255 -3070 0 3
rlabel polysilicon 1262 -3064 1262 -3064 0 1
rlabel polysilicon 1262 -3070 1262 -3070 0 3
rlabel polysilicon 1269 -3064 1269 -3064 0 1
rlabel polysilicon 1269 -3070 1269 -3070 0 3
rlabel polysilicon 1276 -3064 1276 -3064 0 1
rlabel polysilicon 1276 -3070 1276 -3070 0 3
rlabel polysilicon 1283 -3064 1283 -3064 0 1
rlabel polysilicon 1283 -3070 1283 -3070 0 3
rlabel polysilicon 1286 -3070 1286 -3070 0 4
rlabel polysilicon 1290 -3064 1290 -3064 0 1
rlabel polysilicon 1290 -3070 1290 -3070 0 3
rlabel polysilicon 1297 -3064 1297 -3064 0 1
rlabel polysilicon 1297 -3070 1297 -3070 0 3
rlabel polysilicon 1304 -3064 1304 -3064 0 1
rlabel polysilicon 1304 -3070 1304 -3070 0 3
rlabel polysilicon 1311 -3064 1311 -3064 0 1
rlabel polysilicon 1311 -3070 1311 -3070 0 3
rlabel polysilicon 1318 -3064 1318 -3064 0 1
rlabel polysilicon 1318 -3070 1318 -3070 0 3
rlabel polysilicon 1325 -3064 1325 -3064 0 1
rlabel polysilicon 1325 -3070 1325 -3070 0 3
rlabel polysilicon 1332 -3064 1332 -3064 0 1
rlabel polysilicon 1332 -3070 1332 -3070 0 3
rlabel polysilicon 1339 -3064 1339 -3064 0 1
rlabel polysilicon 1339 -3070 1339 -3070 0 3
rlabel polysilicon 1346 -3064 1346 -3064 0 1
rlabel polysilicon 1346 -3070 1346 -3070 0 3
rlabel polysilicon 1374 -3064 1374 -3064 0 1
rlabel polysilicon 1374 -3070 1374 -3070 0 3
rlabel polysilicon 1381 -3064 1381 -3064 0 1
rlabel polysilicon 1381 -3070 1381 -3070 0 3
rlabel polysilicon 1416 -3064 1416 -3064 0 1
rlabel polysilicon 1416 -3070 1416 -3070 0 3
rlabel polysilicon 1458 -3064 1458 -3064 0 1
rlabel polysilicon 1458 -3070 1458 -3070 0 3
rlabel polysilicon 1465 -3064 1465 -3064 0 1
rlabel polysilicon 1465 -3070 1465 -3070 0 3
rlabel polysilicon 1472 -3064 1472 -3064 0 1
rlabel polysilicon 1472 -3070 1472 -3070 0 3
rlabel polysilicon 79 -3153 79 -3153 0 1
rlabel polysilicon 79 -3159 79 -3159 0 3
rlabel polysilicon 86 -3153 86 -3153 0 1
rlabel polysilicon 86 -3159 86 -3159 0 3
rlabel polysilicon 93 -3153 93 -3153 0 1
rlabel polysilicon 93 -3159 93 -3159 0 3
rlabel polysilicon 100 -3153 100 -3153 0 1
rlabel polysilicon 100 -3159 100 -3159 0 3
rlabel polysilicon 107 -3153 107 -3153 0 1
rlabel polysilicon 107 -3159 107 -3159 0 3
rlabel polysilicon 114 -3153 114 -3153 0 1
rlabel polysilicon 114 -3159 114 -3159 0 3
rlabel polysilicon 121 -3153 121 -3153 0 1
rlabel polysilicon 121 -3159 121 -3159 0 3
rlabel polysilicon 128 -3153 128 -3153 0 1
rlabel polysilicon 128 -3159 128 -3159 0 3
rlabel polysilicon 135 -3153 135 -3153 0 1
rlabel polysilicon 135 -3159 135 -3159 0 3
rlabel polysilicon 142 -3153 142 -3153 0 1
rlabel polysilicon 142 -3159 142 -3159 0 3
rlabel polysilicon 149 -3153 149 -3153 0 1
rlabel polysilicon 149 -3159 149 -3159 0 3
rlabel polysilicon 156 -3153 156 -3153 0 1
rlabel polysilicon 156 -3159 156 -3159 0 3
rlabel polysilicon 163 -3153 163 -3153 0 1
rlabel polysilicon 163 -3159 163 -3159 0 3
rlabel polysilicon 170 -3153 170 -3153 0 1
rlabel polysilicon 170 -3159 170 -3159 0 3
rlabel polysilicon 177 -3153 177 -3153 0 1
rlabel polysilicon 177 -3159 177 -3159 0 3
rlabel polysilicon 187 -3153 187 -3153 0 2
rlabel polysilicon 187 -3159 187 -3159 0 4
rlabel polysilicon 191 -3153 191 -3153 0 1
rlabel polysilicon 191 -3159 191 -3159 0 3
rlabel polysilicon 198 -3153 198 -3153 0 1
rlabel polysilicon 198 -3159 198 -3159 0 3
rlabel polysilicon 205 -3153 205 -3153 0 1
rlabel polysilicon 205 -3159 205 -3159 0 3
rlabel polysilicon 215 -3153 215 -3153 0 2
rlabel polysilicon 212 -3159 212 -3159 0 3
rlabel polysilicon 215 -3159 215 -3159 0 4
rlabel polysilicon 219 -3153 219 -3153 0 1
rlabel polysilicon 222 -3153 222 -3153 0 2
rlabel polysilicon 222 -3159 222 -3159 0 4
rlabel polysilicon 226 -3153 226 -3153 0 1
rlabel polysilicon 226 -3159 226 -3159 0 3
rlabel polysilicon 233 -3153 233 -3153 0 1
rlabel polysilicon 233 -3159 233 -3159 0 3
rlabel polysilicon 240 -3153 240 -3153 0 1
rlabel polysilicon 240 -3159 240 -3159 0 3
rlabel polysilicon 247 -3153 247 -3153 0 1
rlabel polysilicon 247 -3159 247 -3159 0 3
rlabel polysilicon 254 -3153 254 -3153 0 1
rlabel polysilicon 254 -3159 254 -3159 0 3
rlabel polysilicon 261 -3153 261 -3153 0 1
rlabel polysilicon 261 -3159 261 -3159 0 3
rlabel polysilicon 268 -3153 268 -3153 0 1
rlabel polysilicon 268 -3159 268 -3159 0 3
rlabel polysilicon 275 -3153 275 -3153 0 1
rlabel polysilicon 275 -3159 275 -3159 0 3
rlabel polysilicon 282 -3153 282 -3153 0 1
rlabel polysilicon 282 -3159 282 -3159 0 3
rlabel polysilicon 289 -3153 289 -3153 0 1
rlabel polysilicon 289 -3159 289 -3159 0 3
rlabel polysilicon 296 -3153 296 -3153 0 1
rlabel polysilicon 296 -3159 296 -3159 0 3
rlabel polysilicon 303 -3153 303 -3153 0 1
rlabel polysilicon 306 -3159 306 -3159 0 4
rlabel polysilicon 310 -3153 310 -3153 0 1
rlabel polysilicon 310 -3159 310 -3159 0 3
rlabel polysilicon 317 -3153 317 -3153 0 1
rlabel polysilicon 317 -3159 317 -3159 0 3
rlabel polysilicon 324 -3153 324 -3153 0 1
rlabel polysilicon 324 -3159 324 -3159 0 3
rlabel polysilicon 331 -3153 331 -3153 0 1
rlabel polysilicon 331 -3159 331 -3159 0 3
rlabel polysilicon 338 -3153 338 -3153 0 1
rlabel polysilicon 338 -3159 338 -3159 0 3
rlabel polysilicon 345 -3153 345 -3153 0 1
rlabel polysilicon 345 -3159 345 -3159 0 3
rlabel polysilicon 352 -3153 352 -3153 0 1
rlabel polysilicon 352 -3159 352 -3159 0 3
rlabel polysilicon 359 -3153 359 -3153 0 1
rlabel polysilicon 362 -3153 362 -3153 0 2
rlabel polysilicon 359 -3159 359 -3159 0 3
rlabel polysilicon 362 -3159 362 -3159 0 4
rlabel polysilicon 366 -3153 366 -3153 0 1
rlabel polysilicon 366 -3159 366 -3159 0 3
rlabel polysilicon 373 -3153 373 -3153 0 1
rlabel polysilicon 373 -3159 373 -3159 0 3
rlabel polysilicon 380 -3153 380 -3153 0 1
rlabel polysilicon 380 -3159 380 -3159 0 3
rlabel polysilicon 387 -3153 387 -3153 0 1
rlabel polysilicon 387 -3159 387 -3159 0 3
rlabel polysilicon 394 -3153 394 -3153 0 1
rlabel polysilicon 394 -3159 394 -3159 0 3
rlabel polysilicon 401 -3153 401 -3153 0 1
rlabel polysilicon 401 -3159 401 -3159 0 3
rlabel polysilicon 408 -3153 408 -3153 0 1
rlabel polysilicon 408 -3159 408 -3159 0 3
rlabel polysilicon 415 -3153 415 -3153 0 1
rlabel polysilicon 415 -3159 415 -3159 0 3
rlabel polysilicon 422 -3153 422 -3153 0 1
rlabel polysilicon 422 -3159 422 -3159 0 3
rlabel polysilicon 432 -3159 432 -3159 0 4
rlabel polysilicon 436 -3153 436 -3153 0 1
rlabel polysilicon 436 -3159 436 -3159 0 3
rlabel polysilicon 443 -3153 443 -3153 0 1
rlabel polysilicon 443 -3159 443 -3159 0 3
rlabel polysilicon 450 -3153 450 -3153 0 1
rlabel polysilicon 450 -3159 450 -3159 0 3
rlabel polysilicon 457 -3153 457 -3153 0 1
rlabel polysilicon 457 -3159 457 -3159 0 3
rlabel polysilicon 464 -3153 464 -3153 0 1
rlabel polysilicon 464 -3159 464 -3159 0 3
rlabel polysilicon 471 -3153 471 -3153 0 1
rlabel polysilicon 471 -3159 471 -3159 0 3
rlabel polysilicon 478 -3153 478 -3153 0 1
rlabel polysilicon 478 -3159 478 -3159 0 3
rlabel polysilicon 485 -3153 485 -3153 0 1
rlabel polysilicon 485 -3159 485 -3159 0 3
rlabel polysilicon 492 -3153 492 -3153 0 1
rlabel polysilicon 492 -3159 492 -3159 0 3
rlabel polysilicon 499 -3153 499 -3153 0 1
rlabel polysilicon 499 -3159 499 -3159 0 3
rlabel polysilicon 506 -3153 506 -3153 0 1
rlabel polysilicon 506 -3159 506 -3159 0 3
rlabel polysilicon 513 -3153 513 -3153 0 1
rlabel polysilicon 513 -3159 513 -3159 0 3
rlabel polysilicon 520 -3153 520 -3153 0 1
rlabel polysilicon 527 -3153 527 -3153 0 1
rlabel polysilicon 527 -3159 527 -3159 0 3
rlabel polysilicon 534 -3153 534 -3153 0 1
rlabel polysilicon 534 -3159 534 -3159 0 3
rlabel polysilicon 541 -3153 541 -3153 0 1
rlabel polysilicon 541 -3159 541 -3159 0 3
rlabel polysilicon 548 -3153 548 -3153 0 1
rlabel polysilicon 548 -3159 548 -3159 0 3
rlabel polysilicon 555 -3153 555 -3153 0 1
rlabel polysilicon 555 -3159 555 -3159 0 3
rlabel polysilicon 562 -3153 562 -3153 0 1
rlabel polysilicon 562 -3159 562 -3159 0 3
rlabel polysilicon 569 -3153 569 -3153 0 1
rlabel polysilicon 569 -3159 569 -3159 0 3
rlabel polysilicon 576 -3153 576 -3153 0 1
rlabel polysilicon 579 -3153 579 -3153 0 2
rlabel polysilicon 579 -3159 579 -3159 0 4
rlabel polysilicon 583 -3153 583 -3153 0 1
rlabel polysilicon 583 -3159 583 -3159 0 3
rlabel polysilicon 590 -3153 590 -3153 0 1
rlabel polysilicon 590 -3159 590 -3159 0 3
rlabel polysilicon 597 -3153 597 -3153 0 1
rlabel polysilicon 597 -3159 597 -3159 0 3
rlabel polysilicon 604 -3153 604 -3153 0 1
rlabel polysilicon 607 -3153 607 -3153 0 2
rlabel polysilicon 604 -3159 604 -3159 0 3
rlabel polysilicon 611 -3153 611 -3153 0 1
rlabel polysilicon 611 -3159 611 -3159 0 3
rlabel polysilicon 621 -3153 621 -3153 0 2
rlabel polysilicon 618 -3159 618 -3159 0 3
rlabel polysilicon 625 -3153 625 -3153 0 1
rlabel polysilicon 625 -3159 625 -3159 0 3
rlabel polysilicon 632 -3153 632 -3153 0 1
rlabel polysilicon 635 -3153 635 -3153 0 2
rlabel polysilicon 632 -3159 632 -3159 0 3
rlabel polysilicon 639 -3153 639 -3153 0 1
rlabel polysilicon 639 -3159 639 -3159 0 3
rlabel polysilicon 646 -3153 646 -3153 0 1
rlabel polysilicon 646 -3159 646 -3159 0 3
rlabel polysilicon 653 -3153 653 -3153 0 1
rlabel polysilicon 656 -3153 656 -3153 0 2
rlabel polysilicon 656 -3159 656 -3159 0 4
rlabel polysilicon 660 -3153 660 -3153 0 1
rlabel polysilicon 660 -3159 660 -3159 0 3
rlabel polysilicon 663 -3159 663 -3159 0 4
rlabel polysilicon 667 -3153 667 -3153 0 1
rlabel polysilicon 667 -3159 667 -3159 0 3
rlabel polysilicon 674 -3153 674 -3153 0 1
rlabel polysilicon 674 -3159 674 -3159 0 3
rlabel polysilicon 681 -3153 681 -3153 0 1
rlabel polysilicon 681 -3159 681 -3159 0 3
rlabel polysilicon 688 -3159 688 -3159 0 3
rlabel polysilicon 695 -3153 695 -3153 0 1
rlabel polysilicon 695 -3159 695 -3159 0 3
rlabel polysilicon 705 -3153 705 -3153 0 2
rlabel polysilicon 702 -3159 702 -3159 0 3
rlabel polysilicon 705 -3159 705 -3159 0 4
rlabel polysilicon 709 -3153 709 -3153 0 1
rlabel polysilicon 709 -3159 709 -3159 0 3
rlabel polysilicon 716 -3153 716 -3153 0 1
rlabel polysilicon 716 -3159 716 -3159 0 3
rlabel polysilicon 723 -3153 723 -3153 0 1
rlabel polysilicon 723 -3159 723 -3159 0 3
rlabel polysilicon 730 -3153 730 -3153 0 1
rlabel polysilicon 730 -3159 730 -3159 0 3
rlabel polysilicon 733 -3159 733 -3159 0 4
rlabel polysilicon 737 -3153 737 -3153 0 1
rlabel polysilicon 737 -3159 737 -3159 0 3
rlabel polysilicon 744 -3153 744 -3153 0 1
rlabel polysilicon 744 -3159 744 -3159 0 3
rlabel polysilicon 751 -3153 751 -3153 0 1
rlabel polysilicon 751 -3159 751 -3159 0 3
rlabel polysilicon 758 -3153 758 -3153 0 1
rlabel polysilicon 758 -3159 758 -3159 0 3
rlabel polysilicon 765 -3153 765 -3153 0 1
rlabel polysilicon 765 -3159 765 -3159 0 3
rlabel polysilicon 772 -3153 772 -3153 0 1
rlabel polysilicon 775 -3153 775 -3153 0 2
rlabel polysilicon 772 -3159 772 -3159 0 3
rlabel polysilicon 775 -3159 775 -3159 0 4
rlabel polysilicon 779 -3153 779 -3153 0 1
rlabel polysilicon 782 -3153 782 -3153 0 2
rlabel polysilicon 779 -3159 779 -3159 0 3
rlabel polysilicon 782 -3159 782 -3159 0 4
rlabel polysilicon 786 -3153 786 -3153 0 1
rlabel polysilicon 786 -3159 786 -3159 0 3
rlabel polysilicon 793 -3153 793 -3153 0 1
rlabel polysilicon 793 -3159 793 -3159 0 3
rlabel polysilicon 800 -3153 800 -3153 0 1
rlabel polysilicon 800 -3159 800 -3159 0 3
rlabel polysilicon 807 -3153 807 -3153 0 1
rlabel polysilicon 807 -3159 807 -3159 0 3
rlabel polysilicon 814 -3153 814 -3153 0 1
rlabel polysilicon 814 -3159 814 -3159 0 3
rlabel polysilicon 821 -3153 821 -3153 0 1
rlabel polysilicon 821 -3159 821 -3159 0 3
rlabel polysilicon 828 -3153 828 -3153 0 1
rlabel polysilicon 828 -3159 828 -3159 0 3
rlabel polysilicon 835 -3153 835 -3153 0 1
rlabel polysilicon 835 -3159 835 -3159 0 3
rlabel polysilicon 842 -3153 842 -3153 0 1
rlabel polysilicon 845 -3153 845 -3153 0 2
rlabel polysilicon 845 -3159 845 -3159 0 4
rlabel polysilicon 849 -3153 849 -3153 0 1
rlabel polysilicon 849 -3159 849 -3159 0 3
rlabel polysilicon 856 -3153 856 -3153 0 1
rlabel polysilicon 856 -3159 856 -3159 0 3
rlabel polysilicon 863 -3153 863 -3153 0 1
rlabel polysilicon 863 -3159 863 -3159 0 3
rlabel polysilicon 870 -3153 870 -3153 0 1
rlabel polysilicon 870 -3159 870 -3159 0 3
rlabel polysilicon 877 -3153 877 -3153 0 1
rlabel polysilicon 880 -3153 880 -3153 0 2
rlabel polysilicon 880 -3159 880 -3159 0 4
rlabel polysilicon 884 -3153 884 -3153 0 1
rlabel polysilicon 884 -3159 884 -3159 0 3
rlabel polysilicon 891 -3153 891 -3153 0 1
rlabel polysilicon 891 -3159 891 -3159 0 3
rlabel polysilicon 898 -3153 898 -3153 0 1
rlabel polysilicon 898 -3159 898 -3159 0 3
rlabel polysilicon 905 -3153 905 -3153 0 1
rlabel polysilicon 905 -3159 905 -3159 0 3
rlabel polysilicon 912 -3153 912 -3153 0 1
rlabel polysilicon 912 -3159 912 -3159 0 3
rlabel polysilicon 919 -3153 919 -3153 0 1
rlabel polysilicon 919 -3159 919 -3159 0 3
rlabel polysilicon 926 -3153 926 -3153 0 1
rlabel polysilicon 926 -3159 926 -3159 0 3
rlabel polysilicon 933 -3153 933 -3153 0 1
rlabel polysilicon 933 -3159 933 -3159 0 3
rlabel polysilicon 940 -3153 940 -3153 0 1
rlabel polysilicon 940 -3159 940 -3159 0 3
rlabel polysilicon 947 -3153 947 -3153 0 1
rlabel polysilicon 947 -3159 947 -3159 0 3
rlabel polysilicon 954 -3153 954 -3153 0 1
rlabel polysilicon 954 -3159 954 -3159 0 3
rlabel polysilicon 961 -3153 961 -3153 0 1
rlabel polysilicon 964 -3153 964 -3153 0 2
rlabel polysilicon 961 -3159 961 -3159 0 3
rlabel polysilicon 964 -3159 964 -3159 0 4
rlabel polysilicon 968 -3153 968 -3153 0 1
rlabel polysilicon 968 -3159 968 -3159 0 3
rlabel polysilicon 975 -3153 975 -3153 0 1
rlabel polysilicon 975 -3159 975 -3159 0 3
rlabel polysilicon 982 -3153 982 -3153 0 1
rlabel polysilicon 982 -3159 982 -3159 0 3
rlabel polysilicon 989 -3153 989 -3153 0 1
rlabel polysilicon 989 -3159 989 -3159 0 3
rlabel polysilicon 996 -3159 996 -3159 0 3
rlabel polysilicon 999 -3159 999 -3159 0 4
rlabel polysilicon 1003 -3153 1003 -3153 0 1
rlabel polysilicon 1003 -3159 1003 -3159 0 3
rlabel polysilicon 1010 -3153 1010 -3153 0 1
rlabel polysilicon 1010 -3159 1010 -3159 0 3
rlabel polysilicon 1017 -3153 1017 -3153 0 1
rlabel polysilicon 1017 -3159 1017 -3159 0 3
rlabel polysilicon 1024 -3153 1024 -3153 0 1
rlabel polysilicon 1024 -3159 1024 -3159 0 3
rlabel polysilicon 1031 -3153 1031 -3153 0 1
rlabel polysilicon 1031 -3159 1031 -3159 0 3
rlabel polysilicon 1038 -3153 1038 -3153 0 1
rlabel polysilicon 1038 -3159 1038 -3159 0 3
rlabel polysilicon 1045 -3153 1045 -3153 0 1
rlabel polysilicon 1045 -3159 1045 -3159 0 3
rlabel polysilicon 1052 -3153 1052 -3153 0 1
rlabel polysilicon 1052 -3159 1052 -3159 0 3
rlabel polysilicon 1059 -3153 1059 -3153 0 1
rlabel polysilicon 1059 -3159 1059 -3159 0 3
rlabel polysilicon 1066 -3153 1066 -3153 0 1
rlabel polysilicon 1066 -3159 1066 -3159 0 3
rlabel polysilicon 1073 -3153 1073 -3153 0 1
rlabel polysilicon 1073 -3159 1073 -3159 0 3
rlabel polysilicon 1080 -3153 1080 -3153 0 1
rlabel polysilicon 1080 -3159 1080 -3159 0 3
rlabel polysilicon 1090 -3153 1090 -3153 0 2
rlabel polysilicon 1094 -3153 1094 -3153 0 1
rlabel polysilicon 1094 -3159 1094 -3159 0 3
rlabel polysilicon 1097 -3159 1097 -3159 0 4
rlabel polysilicon 1101 -3153 1101 -3153 0 1
rlabel polysilicon 1101 -3159 1101 -3159 0 3
rlabel polysilicon 1108 -3153 1108 -3153 0 1
rlabel polysilicon 1108 -3159 1108 -3159 0 3
rlabel polysilicon 1115 -3153 1115 -3153 0 1
rlabel polysilicon 1115 -3159 1115 -3159 0 3
rlabel polysilicon 1122 -3153 1122 -3153 0 1
rlabel polysilicon 1122 -3159 1122 -3159 0 3
rlabel polysilicon 1129 -3153 1129 -3153 0 1
rlabel polysilicon 1129 -3159 1129 -3159 0 3
rlabel polysilicon 1136 -3153 1136 -3153 0 1
rlabel polysilicon 1136 -3159 1136 -3159 0 3
rlabel polysilicon 1143 -3153 1143 -3153 0 1
rlabel polysilicon 1143 -3159 1143 -3159 0 3
rlabel polysilicon 1150 -3153 1150 -3153 0 1
rlabel polysilicon 1150 -3159 1150 -3159 0 3
rlabel polysilicon 1157 -3153 1157 -3153 0 1
rlabel polysilicon 1157 -3159 1157 -3159 0 3
rlabel polysilicon 1164 -3153 1164 -3153 0 1
rlabel polysilicon 1164 -3159 1164 -3159 0 3
rlabel polysilicon 1171 -3153 1171 -3153 0 1
rlabel polysilicon 1171 -3159 1171 -3159 0 3
rlabel polysilicon 1178 -3153 1178 -3153 0 1
rlabel polysilicon 1178 -3159 1178 -3159 0 3
rlabel polysilicon 1188 -3153 1188 -3153 0 2
rlabel polysilicon 1185 -3159 1185 -3159 0 3
rlabel polysilicon 1188 -3159 1188 -3159 0 4
rlabel polysilicon 1192 -3153 1192 -3153 0 1
rlabel polysilicon 1192 -3159 1192 -3159 0 3
rlabel polysilicon 1199 -3153 1199 -3153 0 1
rlabel polysilicon 1199 -3159 1199 -3159 0 3
rlabel polysilicon 1206 -3153 1206 -3153 0 1
rlabel polysilicon 1206 -3159 1206 -3159 0 3
rlabel polysilicon 1213 -3153 1213 -3153 0 1
rlabel polysilicon 1213 -3159 1213 -3159 0 3
rlabel polysilicon 1220 -3153 1220 -3153 0 1
rlabel polysilicon 1220 -3159 1220 -3159 0 3
rlabel polysilicon 1227 -3153 1227 -3153 0 1
rlabel polysilicon 1230 -3153 1230 -3153 0 2
rlabel polysilicon 1227 -3159 1227 -3159 0 3
rlabel polysilicon 1237 -3159 1237 -3159 0 4
rlabel polysilicon 1241 -3153 1241 -3153 0 1
rlabel polysilicon 1241 -3159 1241 -3159 0 3
rlabel polysilicon 1244 -3159 1244 -3159 0 4
rlabel polysilicon 1262 -3153 1262 -3153 0 1
rlabel polysilicon 1262 -3159 1262 -3159 0 3
rlabel polysilicon 1276 -3153 1276 -3153 0 1
rlabel polysilicon 1276 -3159 1276 -3159 0 3
rlabel polysilicon 1290 -3153 1290 -3153 0 1
rlabel polysilicon 1293 -3153 1293 -3153 0 2
rlabel polysilicon 1293 -3159 1293 -3159 0 4
rlabel polysilicon 1346 -3153 1346 -3153 0 1
rlabel polysilicon 1346 -3159 1346 -3159 0 3
rlabel polysilicon 1353 -3153 1353 -3153 0 1
rlabel polysilicon 1353 -3159 1353 -3159 0 3
rlabel polysilicon 1367 -3153 1367 -3153 0 1
rlabel polysilicon 1367 -3159 1367 -3159 0 3
rlabel polysilicon 1409 -3153 1409 -3153 0 1
rlabel polysilicon 1409 -3159 1409 -3159 0 3
rlabel polysilicon 1451 -3153 1451 -3153 0 1
rlabel polysilicon 1451 -3159 1451 -3159 0 3
rlabel polysilicon 1458 -3153 1458 -3153 0 1
rlabel polysilicon 1458 -3159 1458 -3159 0 3
rlabel polysilicon 1465 -3153 1465 -3153 0 1
rlabel polysilicon 1465 -3159 1465 -3159 0 3
rlabel polysilicon 58 -3214 58 -3214 0 1
rlabel polysilicon 58 -3220 58 -3220 0 3
rlabel polysilicon 65 -3214 65 -3214 0 1
rlabel polysilicon 65 -3220 65 -3220 0 3
rlabel polysilicon 72 -3214 72 -3214 0 1
rlabel polysilicon 72 -3220 72 -3220 0 3
rlabel polysilicon 79 -3214 79 -3214 0 1
rlabel polysilicon 79 -3220 79 -3220 0 3
rlabel polysilicon 86 -3214 86 -3214 0 1
rlabel polysilicon 86 -3220 86 -3220 0 3
rlabel polysilicon 93 -3214 93 -3214 0 1
rlabel polysilicon 93 -3220 93 -3220 0 3
rlabel polysilicon 100 -3214 100 -3214 0 1
rlabel polysilicon 100 -3220 100 -3220 0 3
rlabel polysilicon 107 -3214 107 -3214 0 1
rlabel polysilicon 107 -3220 107 -3220 0 3
rlabel polysilicon 114 -3220 114 -3220 0 3
rlabel polysilicon 117 -3220 117 -3220 0 4
rlabel polysilicon 121 -3214 121 -3214 0 1
rlabel polysilicon 121 -3220 121 -3220 0 3
rlabel polysilicon 128 -3214 128 -3214 0 1
rlabel polysilicon 131 -3214 131 -3214 0 2
rlabel polysilicon 128 -3220 128 -3220 0 3
rlabel polysilicon 131 -3220 131 -3220 0 4
rlabel polysilicon 135 -3214 135 -3214 0 1
rlabel polysilicon 135 -3220 135 -3220 0 3
rlabel polysilicon 142 -3214 142 -3214 0 1
rlabel polysilicon 145 -3214 145 -3214 0 2
rlabel polysilicon 152 -3214 152 -3214 0 2
rlabel polysilicon 149 -3220 149 -3220 0 3
rlabel polysilicon 152 -3220 152 -3220 0 4
rlabel polysilicon 156 -3214 156 -3214 0 1
rlabel polysilicon 156 -3220 156 -3220 0 3
rlabel polysilicon 163 -3214 163 -3214 0 1
rlabel polysilicon 163 -3220 163 -3220 0 3
rlabel polysilicon 173 -3214 173 -3214 0 2
rlabel polysilicon 173 -3220 173 -3220 0 4
rlabel polysilicon 180 -3214 180 -3214 0 2
rlabel polysilicon 180 -3220 180 -3220 0 4
rlabel polysilicon 184 -3214 184 -3214 0 1
rlabel polysilicon 184 -3220 184 -3220 0 3
rlabel polysilicon 191 -3214 191 -3214 0 1
rlabel polysilicon 194 -3214 194 -3214 0 2
rlabel polysilicon 191 -3220 191 -3220 0 3
rlabel polysilicon 198 -3214 198 -3214 0 1
rlabel polysilicon 201 -3214 201 -3214 0 2
rlabel polysilicon 198 -3220 198 -3220 0 3
rlabel polysilicon 201 -3220 201 -3220 0 4
rlabel polysilicon 205 -3214 205 -3214 0 1
rlabel polysilicon 208 -3214 208 -3214 0 2
rlabel polysilicon 208 -3220 208 -3220 0 4
rlabel polysilicon 212 -3214 212 -3214 0 1
rlabel polysilicon 212 -3220 212 -3220 0 3
rlabel polysilicon 219 -3214 219 -3214 0 1
rlabel polysilicon 219 -3220 219 -3220 0 3
rlabel polysilicon 226 -3214 226 -3214 0 1
rlabel polysilicon 226 -3220 226 -3220 0 3
rlabel polysilicon 233 -3214 233 -3214 0 1
rlabel polysilicon 233 -3220 233 -3220 0 3
rlabel polysilicon 240 -3214 240 -3214 0 1
rlabel polysilicon 240 -3220 240 -3220 0 3
rlabel polysilicon 247 -3214 247 -3214 0 1
rlabel polysilicon 250 -3214 250 -3214 0 2
rlabel polysilicon 247 -3220 247 -3220 0 3
rlabel polysilicon 250 -3220 250 -3220 0 4
rlabel polysilicon 254 -3214 254 -3214 0 1
rlabel polysilicon 261 -3214 261 -3214 0 1
rlabel polysilicon 264 -3214 264 -3214 0 2
rlabel polysilicon 261 -3220 261 -3220 0 3
rlabel polysilicon 264 -3220 264 -3220 0 4
rlabel polysilicon 268 -3214 268 -3214 0 1
rlabel polysilicon 268 -3220 268 -3220 0 3
rlabel polysilicon 275 -3214 275 -3214 0 1
rlabel polysilicon 275 -3220 275 -3220 0 3
rlabel polysilicon 282 -3214 282 -3214 0 1
rlabel polysilicon 282 -3220 282 -3220 0 3
rlabel polysilicon 289 -3214 289 -3214 0 1
rlabel polysilicon 289 -3220 289 -3220 0 3
rlabel polysilicon 296 -3214 296 -3214 0 1
rlabel polysilicon 296 -3220 296 -3220 0 3
rlabel polysilicon 303 -3214 303 -3214 0 1
rlabel polysilicon 303 -3220 303 -3220 0 3
rlabel polysilicon 310 -3214 310 -3214 0 1
rlabel polysilicon 310 -3220 310 -3220 0 3
rlabel polysilicon 317 -3214 317 -3214 0 1
rlabel polysilicon 317 -3220 317 -3220 0 3
rlabel polysilicon 324 -3214 324 -3214 0 1
rlabel polysilicon 327 -3214 327 -3214 0 2
rlabel polysilicon 324 -3220 324 -3220 0 3
rlabel polysilicon 331 -3214 331 -3214 0 1
rlabel polysilicon 331 -3220 331 -3220 0 3
rlabel polysilicon 338 -3214 338 -3214 0 1
rlabel polysilicon 338 -3220 338 -3220 0 3
rlabel polysilicon 345 -3214 345 -3214 0 1
rlabel polysilicon 352 -3214 352 -3214 0 1
rlabel polysilicon 352 -3220 352 -3220 0 3
rlabel polysilicon 359 -3214 359 -3214 0 1
rlabel polysilicon 359 -3220 359 -3220 0 3
rlabel polysilicon 366 -3214 366 -3214 0 1
rlabel polysilicon 366 -3220 366 -3220 0 3
rlabel polysilicon 373 -3214 373 -3214 0 1
rlabel polysilicon 373 -3220 373 -3220 0 3
rlabel polysilicon 380 -3214 380 -3214 0 1
rlabel polysilicon 380 -3220 380 -3220 0 3
rlabel polysilicon 387 -3214 387 -3214 0 1
rlabel polysilicon 387 -3220 387 -3220 0 3
rlabel polysilicon 394 -3214 394 -3214 0 1
rlabel polysilicon 394 -3220 394 -3220 0 3
rlabel polysilicon 401 -3214 401 -3214 0 1
rlabel polysilicon 401 -3220 401 -3220 0 3
rlabel polysilicon 408 -3214 408 -3214 0 1
rlabel polysilicon 408 -3220 408 -3220 0 3
rlabel polysilicon 415 -3214 415 -3214 0 1
rlabel polysilicon 415 -3220 415 -3220 0 3
rlabel polysilicon 422 -3214 422 -3214 0 1
rlabel polysilicon 422 -3220 422 -3220 0 3
rlabel polysilicon 429 -3214 429 -3214 0 1
rlabel polysilicon 429 -3220 429 -3220 0 3
rlabel polysilicon 436 -3214 436 -3214 0 1
rlabel polysilicon 436 -3220 436 -3220 0 3
rlabel polysilicon 443 -3214 443 -3214 0 1
rlabel polysilicon 443 -3220 443 -3220 0 3
rlabel polysilicon 450 -3214 450 -3214 0 1
rlabel polysilicon 450 -3220 450 -3220 0 3
rlabel polysilicon 457 -3214 457 -3214 0 1
rlabel polysilicon 457 -3220 457 -3220 0 3
rlabel polysilicon 464 -3214 464 -3214 0 1
rlabel polysilicon 464 -3220 464 -3220 0 3
rlabel polysilicon 471 -3214 471 -3214 0 1
rlabel polysilicon 471 -3220 471 -3220 0 3
rlabel polysilicon 478 -3214 478 -3214 0 1
rlabel polysilicon 478 -3220 478 -3220 0 3
rlabel polysilicon 485 -3214 485 -3214 0 1
rlabel polysilicon 485 -3220 485 -3220 0 3
rlabel polysilicon 492 -3214 492 -3214 0 1
rlabel polysilicon 492 -3220 492 -3220 0 3
rlabel polysilicon 499 -3214 499 -3214 0 1
rlabel polysilicon 499 -3220 499 -3220 0 3
rlabel polysilicon 506 -3214 506 -3214 0 1
rlabel polysilicon 506 -3220 506 -3220 0 3
rlabel polysilicon 513 -3214 513 -3214 0 1
rlabel polysilicon 513 -3220 513 -3220 0 3
rlabel polysilicon 520 -3220 520 -3220 0 3
rlabel polysilicon 527 -3214 527 -3214 0 1
rlabel polysilicon 527 -3220 527 -3220 0 3
rlabel polysilicon 534 -3214 534 -3214 0 1
rlabel polysilicon 534 -3220 534 -3220 0 3
rlabel polysilicon 537 -3220 537 -3220 0 4
rlabel polysilicon 541 -3214 541 -3214 0 1
rlabel polysilicon 541 -3220 541 -3220 0 3
rlabel polysilicon 548 -3214 548 -3214 0 1
rlabel polysilicon 548 -3220 548 -3220 0 3
rlabel polysilicon 555 -3214 555 -3214 0 1
rlabel polysilicon 555 -3220 555 -3220 0 3
rlabel polysilicon 558 -3220 558 -3220 0 4
rlabel polysilicon 562 -3214 562 -3214 0 1
rlabel polysilicon 562 -3220 562 -3220 0 3
rlabel polysilicon 569 -3214 569 -3214 0 1
rlabel polysilicon 569 -3220 569 -3220 0 3
rlabel polysilicon 576 -3220 576 -3220 0 3
rlabel polysilicon 579 -3220 579 -3220 0 4
rlabel polysilicon 583 -3214 583 -3214 0 1
rlabel polysilicon 583 -3220 583 -3220 0 3
rlabel polysilicon 590 -3214 590 -3214 0 1
rlabel polysilicon 590 -3220 590 -3220 0 3
rlabel polysilicon 597 -3214 597 -3214 0 1
rlabel polysilicon 597 -3220 597 -3220 0 3
rlabel polysilicon 604 -3214 604 -3214 0 1
rlabel polysilicon 607 -3214 607 -3214 0 2
rlabel polysilicon 604 -3220 604 -3220 0 3
rlabel polysilicon 607 -3220 607 -3220 0 4
rlabel polysilicon 611 -3214 611 -3214 0 1
rlabel polysilicon 611 -3220 611 -3220 0 3
rlabel polysilicon 618 -3214 618 -3214 0 1
rlabel polysilicon 618 -3220 618 -3220 0 3
rlabel polysilicon 625 -3214 625 -3214 0 1
rlabel polysilicon 628 -3220 628 -3220 0 4
rlabel polysilicon 632 -3214 632 -3214 0 1
rlabel polysilicon 635 -3214 635 -3214 0 2
rlabel polysilicon 632 -3220 632 -3220 0 3
rlabel polysilicon 635 -3220 635 -3220 0 4
rlabel polysilicon 639 -3214 639 -3214 0 1
rlabel polysilicon 639 -3220 639 -3220 0 3
rlabel polysilicon 646 -3214 646 -3214 0 1
rlabel polysilicon 646 -3220 646 -3220 0 3
rlabel polysilicon 653 -3214 653 -3214 0 1
rlabel polysilicon 653 -3220 653 -3220 0 3
rlabel polysilicon 660 -3214 660 -3214 0 1
rlabel polysilicon 660 -3220 660 -3220 0 3
rlabel polysilicon 663 -3220 663 -3220 0 4
rlabel polysilicon 667 -3214 667 -3214 0 1
rlabel polysilicon 667 -3220 667 -3220 0 3
rlabel polysilicon 674 -3214 674 -3214 0 1
rlabel polysilicon 674 -3220 674 -3220 0 3
rlabel polysilicon 681 -3214 681 -3214 0 1
rlabel polysilicon 681 -3220 681 -3220 0 3
rlabel polysilicon 688 -3214 688 -3214 0 1
rlabel polysilicon 688 -3220 688 -3220 0 3
rlabel polysilicon 695 -3214 695 -3214 0 1
rlabel polysilicon 695 -3220 695 -3220 0 3
rlabel polysilicon 702 -3214 702 -3214 0 1
rlabel polysilicon 702 -3220 702 -3220 0 3
rlabel polysilicon 709 -3214 709 -3214 0 1
rlabel polysilicon 709 -3220 709 -3220 0 3
rlabel polysilicon 716 -3214 716 -3214 0 1
rlabel polysilicon 716 -3220 716 -3220 0 3
rlabel polysilicon 723 -3214 723 -3214 0 1
rlabel polysilicon 723 -3220 723 -3220 0 3
rlabel polysilicon 730 -3214 730 -3214 0 1
rlabel polysilicon 730 -3220 730 -3220 0 3
rlabel polysilicon 737 -3214 737 -3214 0 1
rlabel polysilicon 737 -3220 737 -3220 0 3
rlabel polysilicon 744 -3214 744 -3214 0 1
rlabel polysilicon 744 -3220 744 -3220 0 3
rlabel polysilicon 751 -3214 751 -3214 0 1
rlabel polysilicon 751 -3220 751 -3220 0 3
rlabel polysilicon 758 -3214 758 -3214 0 1
rlabel polysilicon 761 -3214 761 -3214 0 2
rlabel polysilicon 758 -3220 758 -3220 0 3
rlabel polysilicon 765 -3214 765 -3214 0 1
rlabel polysilicon 765 -3220 765 -3220 0 3
rlabel polysilicon 772 -3214 772 -3214 0 1
rlabel polysilicon 772 -3220 772 -3220 0 3
rlabel polysilicon 779 -3214 779 -3214 0 1
rlabel polysilicon 779 -3220 779 -3220 0 3
rlabel polysilicon 786 -3214 786 -3214 0 1
rlabel polysilicon 786 -3220 786 -3220 0 3
rlabel polysilicon 793 -3214 793 -3214 0 1
rlabel polysilicon 793 -3220 793 -3220 0 3
rlabel polysilicon 800 -3214 800 -3214 0 1
rlabel polysilicon 800 -3220 800 -3220 0 3
rlabel polysilicon 807 -3214 807 -3214 0 1
rlabel polysilicon 807 -3220 807 -3220 0 3
rlabel polysilicon 814 -3214 814 -3214 0 1
rlabel polysilicon 814 -3220 814 -3220 0 3
rlabel polysilicon 821 -3214 821 -3214 0 1
rlabel polysilicon 821 -3220 821 -3220 0 3
rlabel polysilicon 828 -3214 828 -3214 0 1
rlabel polysilicon 828 -3220 828 -3220 0 3
rlabel polysilicon 835 -3214 835 -3214 0 1
rlabel polysilicon 835 -3220 835 -3220 0 3
rlabel polysilicon 842 -3214 842 -3214 0 1
rlabel polysilicon 842 -3220 842 -3220 0 3
rlabel polysilicon 849 -3214 849 -3214 0 1
rlabel polysilicon 849 -3220 849 -3220 0 3
rlabel polysilicon 856 -3214 856 -3214 0 1
rlabel polysilicon 856 -3220 856 -3220 0 3
rlabel polysilicon 863 -3214 863 -3214 0 1
rlabel polysilicon 866 -3214 866 -3214 0 2
rlabel polysilicon 863 -3220 863 -3220 0 3
rlabel polysilicon 866 -3220 866 -3220 0 4
rlabel polysilicon 870 -3214 870 -3214 0 1
rlabel polysilicon 870 -3220 870 -3220 0 3
rlabel polysilicon 877 -3214 877 -3214 0 1
rlabel polysilicon 877 -3220 877 -3220 0 3
rlabel polysilicon 884 -3214 884 -3214 0 1
rlabel polysilicon 884 -3220 884 -3220 0 3
rlabel polysilicon 891 -3214 891 -3214 0 1
rlabel polysilicon 891 -3220 891 -3220 0 3
rlabel polysilicon 898 -3214 898 -3214 0 1
rlabel polysilicon 898 -3220 898 -3220 0 3
rlabel polysilicon 905 -3214 905 -3214 0 1
rlabel polysilicon 905 -3220 905 -3220 0 3
rlabel polysilicon 912 -3214 912 -3214 0 1
rlabel polysilicon 912 -3220 912 -3220 0 3
rlabel polysilicon 919 -3214 919 -3214 0 1
rlabel polysilicon 919 -3220 919 -3220 0 3
rlabel polysilicon 926 -3214 926 -3214 0 1
rlabel polysilicon 926 -3220 926 -3220 0 3
rlabel polysilicon 933 -3214 933 -3214 0 1
rlabel polysilicon 933 -3220 933 -3220 0 3
rlabel polysilicon 940 -3214 940 -3214 0 1
rlabel polysilicon 940 -3220 940 -3220 0 3
rlabel polysilicon 947 -3214 947 -3214 0 1
rlabel polysilicon 947 -3220 947 -3220 0 3
rlabel polysilicon 954 -3214 954 -3214 0 1
rlabel polysilicon 954 -3220 954 -3220 0 3
rlabel polysilicon 961 -3214 961 -3214 0 1
rlabel polysilicon 961 -3220 961 -3220 0 3
rlabel polysilicon 968 -3214 968 -3214 0 1
rlabel polysilicon 968 -3220 968 -3220 0 3
rlabel polysilicon 975 -3214 975 -3214 0 1
rlabel polysilicon 975 -3220 975 -3220 0 3
rlabel polysilicon 982 -3214 982 -3214 0 1
rlabel polysilicon 985 -3214 985 -3214 0 2
rlabel polysilicon 982 -3220 982 -3220 0 3
rlabel polysilicon 985 -3220 985 -3220 0 4
rlabel polysilicon 989 -3214 989 -3214 0 1
rlabel polysilicon 989 -3220 989 -3220 0 3
rlabel polysilicon 996 -3214 996 -3214 0 1
rlabel polysilicon 996 -3220 996 -3220 0 3
rlabel polysilicon 1003 -3214 1003 -3214 0 1
rlabel polysilicon 1006 -3214 1006 -3214 0 2
rlabel polysilicon 1003 -3220 1003 -3220 0 3
rlabel polysilicon 1010 -3214 1010 -3214 0 1
rlabel polysilicon 1010 -3220 1010 -3220 0 3
rlabel polysilicon 1017 -3214 1017 -3214 0 1
rlabel polysilicon 1017 -3220 1017 -3220 0 3
rlabel polysilicon 1024 -3214 1024 -3214 0 1
rlabel polysilicon 1024 -3220 1024 -3220 0 3
rlabel polysilicon 1031 -3214 1031 -3214 0 1
rlabel polysilicon 1031 -3220 1031 -3220 0 3
rlabel polysilicon 1038 -3214 1038 -3214 0 1
rlabel polysilicon 1038 -3220 1038 -3220 0 3
rlabel polysilicon 1045 -3214 1045 -3214 0 1
rlabel polysilicon 1045 -3220 1045 -3220 0 3
rlabel polysilicon 1052 -3214 1052 -3214 0 1
rlabel polysilicon 1052 -3220 1052 -3220 0 3
rlabel polysilicon 1059 -3214 1059 -3214 0 1
rlabel polysilicon 1059 -3220 1059 -3220 0 3
rlabel polysilicon 1062 -3220 1062 -3220 0 4
rlabel polysilicon 1073 -3214 1073 -3214 0 1
rlabel polysilicon 1073 -3220 1073 -3220 0 3
rlabel polysilicon 1080 -3214 1080 -3214 0 1
rlabel polysilicon 1080 -3220 1080 -3220 0 3
rlabel polysilicon 1087 -3214 1087 -3214 0 1
rlabel polysilicon 1087 -3220 1087 -3220 0 3
rlabel polysilicon 1094 -3214 1094 -3214 0 1
rlabel polysilicon 1097 -3214 1097 -3214 0 2
rlabel polysilicon 1094 -3220 1094 -3220 0 3
rlabel polysilicon 1101 -3214 1101 -3214 0 1
rlabel polysilicon 1101 -3220 1101 -3220 0 3
rlabel polysilicon 1111 -3214 1111 -3214 0 2
rlabel polysilicon 1108 -3220 1108 -3220 0 3
rlabel polysilicon 1111 -3220 1111 -3220 0 4
rlabel polysilicon 1115 -3214 1115 -3214 0 1
rlabel polysilicon 1115 -3220 1115 -3220 0 3
rlabel polysilicon 1122 -3214 1122 -3214 0 1
rlabel polysilicon 1122 -3220 1122 -3220 0 3
rlabel polysilicon 1129 -3214 1129 -3214 0 1
rlabel polysilicon 1129 -3220 1129 -3220 0 3
rlabel polysilicon 1136 -3214 1136 -3214 0 1
rlabel polysilicon 1136 -3220 1136 -3220 0 3
rlabel polysilicon 1143 -3214 1143 -3214 0 1
rlabel polysilicon 1143 -3220 1143 -3220 0 3
rlabel polysilicon 1150 -3214 1150 -3214 0 1
rlabel polysilicon 1150 -3220 1150 -3220 0 3
rlabel polysilicon 1157 -3214 1157 -3214 0 1
rlabel polysilicon 1157 -3220 1157 -3220 0 3
rlabel polysilicon 1164 -3214 1164 -3214 0 1
rlabel polysilicon 1167 -3214 1167 -3214 0 2
rlabel polysilicon 1164 -3220 1164 -3220 0 3
rlabel polysilicon 1167 -3220 1167 -3220 0 4
rlabel polysilicon 1171 -3214 1171 -3214 0 1
rlabel polysilicon 1171 -3220 1171 -3220 0 3
rlabel polysilicon 1185 -3214 1185 -3214 0 1
rlabel polysilicon 1185 -3220 1185 -3220 0 3
rlabel polysilicon 1192 -3214 1192 -3214 0 1
rlabel polysilicon 1192 -3220 1192 -3220 0 3
rlabel polysilicon 1199 -3214 1199 -3214 0 1
rlabel polysilicon 1199 -3220 1199 -3220 0 3
rlabel polysilicon 1206 -3214 1206 -3214 0 1
rlabel polysilicon 1206 -3220 1206 -3220 0 3
rlabel polysilicon 1213 -3214 1213 -3214 0 1
rlabel polysilicon 1213 -3220 1213 -3220 0 3
rlabel polysilicon 1234 -3214 1234 -3214 0 1
rlabel polysilicon 1234 -3220 1234 -3220 0 3
rlabel polysilicon 1332 -3214 1332 -3214 0 1
rlabel polysilicon 1332 -3220 1332 -3220 0 3
rlabel polysilicon 1360 -3214 1360 -3214 0 1
rlabel polysilicon 1360 -3220 1360 -3220 0 3
rlabel polysilicon 1367 -3214 1367 -3214 0 1
rlabel polysilicon 1367 -3220 1367 -3220 0 3
rlabel polysilicon 1409 -3214 1409 -3214 0 1
rlabel polysilicon 1409 -3220 1409 -3220 0 3
rlabel polysilicon 1451 -3214 1451 -3214 0 1
rlabel polysilicon 1451 -3220 1451 -3220 0 3
rlabel polysilicon 1454 -3220 1454 -3220 0 4
rlabel polysilicon 1458 -3214 1458 -3214 0 1
rlabel polysilicon 1458 -3220 1458 -3220 0 3
rlabel polysilicon 1465 -3214 1465 -3214 0 1
rlabel polysilicon 1465 -3220 1465 -3220 0 3
rlabel polysilicon 156 -3269 156 -3269 0 1
rlabel polysilicon 156 -3275 156 -3275 0 3
rlabel polysilicon 163 -3269 163 -3269 0 1
rlabel polysilicon 163 -3275 163 -3275 0 3
rlabel polysilicon 170 -3269 170 -3269 0 1
rlabel polysilicon 170 -3275 170 -3275 0 3
rlabel polysilicon 177 -3269 177 -3269 0 1
rlabel polysilicon 177 -3275 177 -3275 0 3
rlabel polysilicon 187 -3269 187 -3269 0 2
rlabel polysilicon 184 -3275 184 -3275 0 3
rlabel polysilicon 187 -3275 187 -3275 0 4
rlabel polysilicon 191 -3269 191 -3269 0 1
rlabel polysilicon 191 -3275 191 -3275 0 3
rlabel polysilicon 198 -3269 198 -3269 0 1
rlabel polysilicon 198 -3275 198 -3275 0 3
rlabel polysilicon 208 -3269 208 -3269 0 2
rlabel polysilicon 208 -3275 208 -3275 0 4
rlabel polysilicon 212 -3269 212 -3269 0 1
rlabel polysilicon 212 -3275 212 -3275 0 3
rlabel polysilicon 219 -3269 219 -3269 0 1
rlabel polysilicon 219 -3275 219 -3275 0 3
rlabel polysilicon 226 -3269 226 -3269 0 1
rlabel polysilicon 226 -3275 226 -3275 0 3
rlabel polysilicon 233 -3269 233 -3269 0 1
rlabel polysilicon 233 -3275 233 -3275 0 3
rlabel polysilicon 240 -3269 240 -3269 0 1
rlabel polysilicon 243 -3269 243 -3269 0 2
rlabel polysilicon 243 -3275 243 -3275 0 4
rlabel polysilicon 247 -3269 247 -3269 0 1
rlabel polysilicon 250 -3269 250 -3269 0 2
rlabel polysilicon 254 -3275 254 -3275 0 3
rlabel polysilicon 261 -3269 261 -3269 0 1
rlabel polysilicon 264 -3269 264 -3269 0 2
rlabel polysilicon 268 -3269 268 -3269 0 1
rlabel polysilicon 268 -3275 268 -3275 0 3
rlabel polysilicon 275 -3269 275 -3269 0 1
rlabel polysilicon 275 -3275 275 -3275 0 3
rlabel polysilicon 282 -3269 282 -3269 0 1
rlabel polysilicon 282 -3275 282 -3275 0 3
rlabel polysilicon 289 -3269 289 -3269 0 1
rlabel polysilicon 289 -3275 289 -3275 0 3
rlabel polysilicon 296 -3269 296 -3269 0 1
rlabel polysilicon 296 -3275 296 -3275 0 3
rlabel polysilicon 303 -3269 303 -3269 0 1
rlabel polysilicon 303 -3275 303 -3275 0 3
rlabel polysilicon 310 -3269 310 -3269 0 1
rlabel polysilicon 310 -3275 310 -3275 0 3
rlabel polysilicon 317 -3269 317 -3269 0 1
rlabel polysilicon 317 -3275 317 -3275 0 3
rlabel polysilicon 324 -3269 324 -3269 0 1
rlabel polysilicon 324 -3275 324 -3275 0 3
rlabel polysilicon 331 -3269 331 -3269 0 1
rlabel polysilicon 331 -3275 331 -3275 0 3
rlabel polysilicon 338 -3269 338 -3269 0 1
rlabel polysilicon 338 -3275 338 -3275 0 3
rlabel polysilicon 345 -3275 345 -3275 0 3
rlabel polysilicon 352 -3269 352 -3269 0 1
rlabel polysilicon 352 -3275 352 -3275 0 3
rlabel polysilicon 359 -3269 359 -3269 0 1
rlabel polysilicon 359 -3275 359 -3275 0 3
rlabel polysilicon 366 -3269 366 -3269 0 1
rlabel polysilicon 366 -3275 366 -3275 0 3
rlabel polysilicon 373 -3269 373 -3269 0 1
rlabel polysilicon 373 -3275 373 -3275 0 3
rlabel polysilicon 380 -3269 380 -3269 0 1
rlabel polysilicon 380 -3275 380 -3275 0 3
rlabel polysilicon 387 -3269 387 -3269 0 1
rlabel polysilicon 387 -3275 387 -3275 0 3
rlabel polysilicon 394 -3269 394 -3269 0 1
rlabel polysilicon 397 -3269 397 -3269 0 2
rlabel polysilicon 394 -3275 394 -3275 0 3
rlabel polysilicon 401 -3269 401 -3269 0 1
rlabel polysilicon 404 -3269 404 -3269 0 2
rlabel polysilicon 401 -3275 401 -3275 0 3
rlabel polysilicon 408 -3269 408 -3269 0 1
rlabel polysilicon 408 -3275 408 -3275 0 3
rlabel polysilicon 415 -3269 415 -3269 0 1
rlabel polysilicon 415 -3275 415 -3275 0 3
rlabel polysilicon 422 -3269 422 -3269 0 1
rlabel polysilicon 422 -3275 422 -3275 0 3
rlabel polysilicon 429 -3269 429 -3269 0 1
rlabel polysilicon 429 -3275 429 -3275 0 3
rlabel polysilicon 436 -3269 436 -3269 0 1
rlabel polysilicon 436 -3275 436 -3275 0 3
rlabel polysilicon 443 -3269 443 -3269 0 1
rlabel polysilicon 443 -3275 443 -3275 0 3
rlabel polysilicon 450 -3269 450 -3269 0 1
rlabel polysilicon 450 -3275 450 -3275 0 3
rlabel polysilicon 457 -3269 457 -3269 0 1
rlabel polysilicon 457 -3275 457 -3275 0 3
rlabel polysilicon 464 -3269 464 -3269 0 1
rlabel polysilicon 464 -3275 464 -3275 0 3
rlabel polysilicon 471 -3269 471 -3269 0 1
rlabel polysilicon 474 -3269 474 -3269 0 2
rlabel polysilicon 474 -3275 474 -3275 0 4
rlabel polysilicon 478 -3269 478 -3269 0 1
rlabel polysilicon 478 -3275 478 -3275 0 3
rlabel polysilicon 485 -3269 485 -3269 0 1
rlabel polysilicon 488 -3269 488 -3269 0 2
rlabel polysilicon 485 -3275 485 -3275 0 3
rlabel polysilicon 488 -3275 488 -3275 0 4
rlabel polysilicon 492 -3269 492 -3269 0 1
rlabel polysilicon 492 -3275 492 -3275 0 3
rlabel polysilicon 499 -3269 499 -3269 0 1
rlabel polysilicon 499 -3275 499 -3275 0 3
rlabel polysilicon 506 -3269 506 -3269 0 1
rlabel polysilicon 506 -3275 506 -3275 0 3
rlabel polysilicon 513 -3269 513 -3269 0 1
rlabel polysilicon 513 -3275 513 -3275 0 3
rlabel polysilicon 520 -3269 520 -3269 0 1
rlabel polysilicon 520 -3275 520 -3275 0 3
rlabel polysilicon 527 -3269 527 -3269 0 1
rlabel polysilicon 527 -3275 527 -3275 0 3
rlabel polysilicon 534 -3269 534 -3269 0 1
rlabel polysilicon 537 -3269 537 -3269 0 2
rlabel polysilicon 534 -3275 534 -3275 0 3
rlabel polysilicon 541 -3269 541 -3269 0 1
rlabel polysilicon 541 -3275 541 -3275 0 3
rlabel polysilicon 548 -3269 548 -3269 0 1
rlabel polysilicon 548 -3275 548 -3275 0 3
rlabel polysilicon 555 -3269 555 -3269 0 1
rlabel polysilicon 555 -3275 555 -3275 0 3
rlabel polysilicon 562 -3269 562 -3269 0 1
rlabel polysilicon 562 -3275 562 -3275 0 3
rlabel polysilicon 569 -3269 569 -3269 0 1
rlabel polysilicon 569 -3275 569 -3275 0 3
rlabel polysilicon 576 -3269 576 -3269 0 1
rlabel polysilicon 576 -3275 576 -3275 0 3
rlabel polysilicon 583 -3269 583 -3269 0 1
rlabel polysilicon 583 -3275 583 -3275 0 3
rlabel polysilicon 590 -3275 590 -3275 0 3
rlabel polysilicon 593 -3275 593 -3275 0 4
rlabel polysilicon 597 -3269 597 -3269 0 1
rlabel polysilicon 597 -3275 597 -3275 0 3
rlabel polysilicon 604 -3269 604 -3269 0 1
rlabel polysilicon 604 -3275 604 -3275 0 3
rlabel polysilicon 611 -3269 611 -3269 0 1
rlabel polysilicon 611 -3275 611 -3275 0 3
rlabel polysilicon 618 -3269 618 -3269 0 1
rlabel polysilicon 618 -3275 618 -3275 0 3
rlabel polysilicon 625 -3269 625 -3269 0 1
rlabel polysilicon 625 -3275 625 -3275 0 3
rlabel polysilicon 632 -3269 632 -3269 0 1
rlabel polysilicon 635 -3269 635 -3269 0 2
rlabel polysilicon 632 -3275 632 -3275 0 3
rlabel polysilicon 635 -3275 635 -3275 0 4
rlabel polysilicon 639 -3269 639 -3269 0 1
rlabel polysilicon 639 -3275 639 -3275 0 3
rlabel polysilicon 646 -3269 646 -3269 0 1
rlabel polysilicon 646 -3275 646 -3275 0 3
rlabel polysilicon 653 -3269 653 -3269 0 1
rlabel polysilicon 653 -3275 653 -3275 0 3
rlabel polysilicon 660 -3269 660 -3269 0 1
rlabel polysilicon 660 -3275 660 -3275 0 3
rlabel polysilicon 667 -3269 667 -3269 0 1
rlabel polysilicon 667 -3275 667 -3275 0 3
rlabel polysilicon 674 -3269 674 -3269 0 1
rlabel polysilicon 674 -3275 674 -3275 0 3
rlabel polysilicon 681 -3269 681 -3269 0 1
rlabel polysilicon 681 -3275 681 -3275 0 3
rlabel polysilicon 688 -3269 688 -3269 0 1
rlabel polysilicon 688 -3275 688 -3275 0 3
rlabel polysilicon 695 -3269 695 -3269 0 1
rlabel polysilicon 695 -3275 695 -3275 0 3
rlabel polysilicon 702 -3269 702 -3269 0 1
rlabel polysilicon 702 -3275 702 -3275 0 3
rlabel polysilicon 709 -3269 709 -3269 0 1
rlabel polysilicon 709 -3275 709 -3275 0 3
rlabel polysilicon 716 -3269 716 -3269 0 1
rlabel polysilicon 716 -3275 716 -3275 0 3
rlabel polysilicon 726 -3269 726 -3269 0 2
rlabel polysilicon 723 -3275 723 -3275 0 3
rlabel polysilicon 733 -3269 733 -3269 0 2
rlabel polysilicon 730 -3275 730 -3275 0 3
rlabel polysilicon 737 -3269 737 -3269 0 1
rlabel polysilicon 737 -3275 737 -3275 0 3
rlabel polysilicon 744 -3269 744 -3269 0 1
rlabel polysilicon 744 -3275 744 -3275 0 3
rlabel polysilicon 751 -3269 751 -3269 0 1
rlabel polysilicon 751 -3275 751 -3275 0 3
rlabel polysilicon 758 -3269 758 -3269 0 1
rlabel polysilicon 758 -3275 758 -3275 0 3
rlabel polysilicon 765 -3269 765 -3269 0 1
rlabel polysilicon 765 -3275 765 -3275 0 3
rlabel polysilicon 772 -3269 772 -3269 0 1
rlabel polysilicon 772 -3275 772 -3275 0 3
rlabel polysilicon 782 -3269 782 -3269 0 2
rlabel polysilicon 779 -3275 779 -3275 0 3
rlabel polysilicon 782 -3275 782 -3275 0 4
rlabel polysilicon 786 -3269 786 -3269 0 1
rlabel polysilicon 786 -3275 786 -3275 0 3
rlabel polysilicon 793 -3269 793 -3269 0 1
rlabel polysilicon 793 -3275 793 -3275 0 3
rlabel polysilicon 800 -3269 800 -3269 0 1
rlabel polysilicon 800 -3275 800 -3275 0 3
rlabel polysilicon 807 -3269 807 -3269 0 1
rlabel polysilicon 807 -3275 807 -3275 0 3
rlabel polysilicon 814 -3269 814 -3269 0 1
rlabel polysilicon 814 -3275 814 -3275 0 3
rlabel polysilicon 821 -3269 821 -3269 0 1
rlabel polysilicon 821 -3275 821 -3275 0 3
rlabel polysilicon 828 -3269 828 -3269 0 1
rlabel polysilicon 828 -3275 828 -3275 0 3
rlabel polysilicon 842 -3269 842 -3269 0 1
rlabel polysilicon 842 -3275 842 -3275 0 3
rlabel polysilicon 870 -3269 870 -3269 0 1
rlabel polysilicon 870 -3275 870 -3275 0 3
rlabel polysilicon 877 -3269 877 -3269 0 1
rlabel polysilicon 880 -3269 880 -3269 0 2
rlabel polysilicon 877 -3275 877 -3275 0 3
rlabel polysilicon 880 -3275 880 -3275 0 4
rlabel polysilicon 884 -3269 884 -3269 0 1
rlabel polysilicon 884 -3275 884 -3275 0 3
rlabel polysilicon 891 -3269 891 -3269 0 1
rlabel polysilicon 891 -3275 891 -3275 0 3
rlabel polysilicon 898 -3269 898 -3269 0 1
rlabel polysilicon 898 -3275 898 -3275 0 3
rlabel polysilicon 905 -3269 905 -3269 0 1
rlabel polysilicon 905 -3275 905 -3275 0 3
rlabel polysilicon 912 -3269 912 -3269 0 1
rlabel polysilicon 912 -3275 912 -3275 0 3
rlabel polysilicon 919 -3269 919 -3269 0 1
rlabel polysilicon 919 -3275 919 -3275 0 3
rlabel polysilicon 926 -3269 926 -3269 0 1
rlabel polysilicon 926 -3275 926 -3275 0 3
rlabel polysilicon 933 -3269 933 -3269 0 1
rlabel polysilicon 933 -3275 933 -3275 0 3
rlabel polysilicon 940 -3269 940 -3269 0 1
rlabel polysilicon 940 -3275 940 -3275 0 3
rlabel polysilicon 947 -3269 947 -3269 0 1
rlabel polysilicon 947 -3275 947 -3275 0 3
rlabel polysilicon 954 -3269 954 -3269 0 1
rlabel polysilicon 954 -3275 954 -3275 0 3
rlabel polysilicon 961 -3269 961 -3269 0 1
rlabel polysilicon 961 -3275 961 -3275 0 3
rlabel polysilicon 982 -3269 982 -3269 0 1
rlabel polysilicon 982 -3275 982 -3275 0 3
rlabel polysilicon 992 -3269 992 -3269 0 2
rlabel polysilicon 992 -3275 992 -3275 0 4
rlabel polysilicon 996 -3269 996 -3269 0 1
rlabel polysilicon 996 -3275 996 -3275 0 3
rlabel polysilicon 1003 -3269 1003 -3269 0 1
rlabel polysilicon 1003 -3275 1003 -3275 0 3
rlabel polysilicon 1066 -3269 1066 -3269 0 1
rlabel polysilicon 1066 -3275 1066 -3275 0 3
rlabel polysilicon 1073 -3269 1073 -3269 0 1
rlabel polysilicon 1073 -3275 1073 -3275 0 3
rlabel polysilicon 1080 -3269 1080 -3269 0 1
rlabel polysilicon 1080 -3275 1080 -3275 0 3
rlabel polysilicon 1094 -3269 1094 -3269 0 1
rlabel polysilicon 1094 -3275 1094 -3275 0 3
rlabel polysilicon 1101 -3269 1101 -3269 0 1
rlabel polysilicon 1101 -3275 1101 -3275 0 3
rlabel polysilicon 1108 -3269 1108 -3269 0 1
rlabel polysilicon 1108 -3275 1108 -3275 0 3
rlabel polysilicon 1122 -3269 1122 -3269 0 1
rlabel polysilicon 1125 -3269 1125 -3269 0 2
rlabel polysilicon 1122 -3275 1122 -3275 0 3
rlabel polysilicon 1125 -3275 1125 -3275 0 4
rlabel polysilicon 1129 -3269 1129 -3269 0 1
rlabel polysilicon 1129 -3275 1129 -3275 0 3
rlabel polysilicon 1136 -3269 1136 -3269 0 1
rlabel polysilicon 1136 -3275 1136 -3275 0 3
rlabel polysilicon 1143 -3269 1143 -3269 0 1
rlabel polysilicon 1143 -3275 1143 -3275 0 3
rlabel polysilicon 1150 -3269 1150 -3269 0 1
rlabel polysilicon 1150 -3275 1150 -3275 0 3
rlabel polysilicon 1160 -3269 1160 -3269 0 2
rlabel polysilicon 1157 -3275 1157 -3275 0 3
rlabel polysilicon 1164 -3269 1164 -3269 0 1
rlabel polysilicon 1164 -3275 1164 -3275 0 3
rlabel polysilicon 1171 -3269 1171 -3269 0 1
rlabel polysilicon 1171 -3275 1171 -3275 0 3
rlabel polysilicon 1185 -3269 1185 -3269 0 1
rlabel polysilicon 1188 -3269 1188 -3269 0 2
rlabel polysilicon 1185 -3275 1185 -3275 0 3
rlabel polysilicon 1206 -3269 1206 -3269 0 1
rlabel polysilicon 1206 -3275 1206 -3275 0 3
rlabel polysilicon 1216 -3269 1216 -3269 0 2
rlabel polysilicon 1216 -3275 1216 -3275 0 4
rlabel polysilicon 1220 -3269 1220 -3269 0 1
rlabel polysilicon 1220 -3275 1220 -3275 0 3
rlabel polysilicon 1234 -3269 1234 -3269 0 1
rlabel polysilicon 1251 -3269 1251 -3269 0 2
rlabel polysilicon 1251 -3275 1251 -3275 0 4
rlabel polysilicon 1290 -3269 1290 -3269 0 1
rlabel polysilicon 1290 -3275 1290 -3275 0 3
rlabel polysilicon 1325 -3269 1325 -3269 0 1
rlabel polysilicon 1328 -3269 1328 -3269 0 2
rlabel polysilicon 1360 -3269 1360 -3269 0 1
rlabel polysilicon 1360 -3275 1360 -3275 0 3
rlabel polysilicon 1367 -3269 1367 -3269 0 1
rlabel polysilicon 1367 -3275 1367 -3275 0 3
rlabel polysilicon 1409 -3269 1409 -3269 0 1
rlabel polysilicon 1409 -3275 1409 -3275 0 3
rlabel polysilicon 1451 -3269 1451 -3269 0 1
rlabel polysilicon 1454 -3269 1454 -3269 0 2
rlabel polysilicon 1451 -3275 1451 -3275 0 3
rlabel polysilicon 1458 -3269 1458 -3269 0 1
rlabel polysilicon 1458 -3275 1458 -3275 0 3
rlabel polysilicon 1461 -3275 1461 -3275 0 4
rlabel polysilicon 1465 -3269 1465 -3269 0 1
rlabel polysilicon 1465 -3275 1465 -3275 0 3
rlabel polysilicon 177 -3332 177 -3332 0 1
rlabel polysilicon 177 -3338 177 -3338 0 3
rlabel polysilicon 184 -3332 184 -3332 0 1
rlabel polysilicon 184 -3338 184 -3338 0 3
rlabel polysilicon 191 -3332 191 -3332 0 1
rlabel polysilicon 191 -3338 191 -3338 0 3
rlabel polysilicon 198 -3332 198 -3332 0 1
rlabel polysilicon 198 -3338 198 -3338 0 3
rlabel polysilicon 205 -3332 205 -3332 0 1
rlabel polysilicon 205 -3338 205 -3338 0 3
rlabel polysilicon 212 -3332 212 -3332 0 1
rlabel polysilicon 212 -3338 212 -3338 0 3
rlabel polysilicon 219 -3332 219 -3332 0 1
rlabel polysilicon 219 -3338 219 -3338 0 3
rlabel polysilicon 226 -3332 226 -3332 0 1
rlabel polysilicon 229 -3332 229 -3332 0 2
rlabel polysilicon 233 -3332 233 -3332 0 1
rlabel polysilicon 240 -3332 240 -3332 0 1
rlabel polysilicon 240 -3338 240 -3338 0 3
rlabel polysilicon 247 -3332 247 -3332 0 1
rlabel polysilicon 247 -3338 247 -3338 0 3
rlabel polysilicon 254 -3332 254 -3332 0 1
rlabel polysilicon 254 -3338 254 -3338 0 3
rlabel polysilicon 261 -3338 261 -3338 0 3
rlabel polysilicon 264 -3338 264 -3338 0 4
rlabel polysilicon 268 -3332 268 -3332 0 1
rlabel polysilicon 268 -3338 268 -3338 0 3
rlabel polysilicon 275 -3332 275 -3332 0 1
rlabel polysilicon 275 -3338 275 -3338 0 3
rlabel polysilicon 282 -3332 282 -3332 0 1
rlabel polysilicon 282 -3338 282 -3338 0 3
rlabel polysilicon 289 -3332 289 -3332 0 1
rlabel polysilicon 289 -3338 289 -3338 0 3
rlabel polysilicon 296 -3332 296 -3332 0 1
rlabel polysilicon 296 -3338 296 -3338 0 3
rlabel polysilicon 303 -3332 303 -3332 0 1
rlabel polysilicon 303 -3338 303 -3338 0 3
rlabel polysilicon 306 -3338 306 -3338 0 4
rlabel polysilicon 310 -3332 310 -3332 0 1
rlabel polysilicon 310 -3338 310 -3338 0 3
rlabel polysilicon 317 -3332 317 -3332 0 1
rlabel polysilicon 317 -3338 317 -3338 0 3
rlabel polysilicon 324 -3332 324 -3332 0 1
rlabel polysilicon 324 -3338 324 -3338 0 3
rlabel polysilicon 331 -3332 331 -3332 0 1
rlabel polysilicon 331 -3338 331 -3338 0 3
rlabel polysilicon 338 -3332 338 -3332 0 1
rlabel polysilicon 338 -3338 338 -3338 0 3
rlabel polysilicon 345 -3332 345 -3332 0 1
rlabel polysilicon 345 -3338 345 -3338 0 3
rlabel polysilicon 352 -3332 352 -3332 0 1
rlabel polysilicon 352 -3338 352 -3338 0 3
rlabel polysilicon 359 -3332 359 -3332 0 1
rlabel polysilicon 359 -3338 359 -3338 0 3
rlabel polysilicon 366 -3332 366 -3332 0 1
rlabel polysilicon 366 -3338 366 -3338 0 3
rlabel polysilicon 373 -3332 373 -3332 0 1
rlabel polysilicon 373 -3338 373 -3338 0 3
rlabel polysilicon 380 -3332 380 -3332 0 1
rlabel polysilicon 383 -3332 383 -3332 0 2
rlabel polysilicon 383 -3338 383 -3338 0 4
rlabel polysilicon 387 -3332 387 -3332 0 1
rlabel polysilicon 387 -3338 387 -3338 0 3
rlabel polysilicon 394 -3332 394 -3332 0 1
rlabel polysilicon 394 -3338 394 -3338 0 3
rlabel polysilicon 401 -3332 401 -3332 0 1
rlabel polysilicon 401 -3338 401 -3338 0 3
rlabel polysilicon 408 -3332 408 -3332 0 1
rlabel polysilicon 411 -3332 411 -3332 0 2
rlabel polysilicon 408 -3338 408 -3338 0 3
rlabel polysilicon 411 -3338 411 -3338 0 4
rlabel polysilicon 415 -3332 415 -3332 0 1
rlabel polysilicon 415 -3338 415 -3338 0 3
rlabel polysilicon 422 -3332 422 -3332 0 1
rlabel polysilicon 422 -3338 422 -3338 0 3
rlabel polysilicon 429 -3332 429 -3332 0 1
rlabel polysilicon 429 -3338 429 -3338 0 3
rlabel polysilicon 436 -3332 436 -3332 0 1
rlabel polysilicon 436 -3338 436 -3338 0 3
rlabel polysilicon 443 -3332 443 -3332 0 1
rlabel polysilicon 446 -3332 446 -3332 0 2
rlabel polysilicon 443 -3338 443 -3338 0 3
rlabel polysilicon 446 -3338 446 -3338 0 4
rlabel polysilicon 450 -3332 450 -3332 0 1
rlabel polysilicon 450 -3338 450 -3338 0 3
rlabel polysilicon 457 -3332 457 -3332 0 1
rlabel polysilicon 457 -3338 457 -3338 0 3
rlabel polysilicon 464 -3332 464 -3332 0 1
rlabel polysilicon 467 -3332 467 -3332 0 2
rlabel polysilicon 467 -3338 467 -3338 0 4
rlabel polysilicon 471 -3332 471 -3332 0 1
rlabel polysilicon 471 -3338 471 -3338 0 3
rlabel polysilicon 478 -3332 478 -3332 0 1
rlabel polysilicon 478 -3338 478 -3338 0 3
rlabel polysilicon 485 -3332 485 -3332 0 1
rlabel polysilicon 485 -3338 485 -3338 0 3
rlabel polysilicon 492 -3332 492 -3332 0 1
rlabel polysilicon 492 -3338 492 -3338 0 3
rlabel polysilicon 499 -3332 499 -3332 0 1
rlabel polysilicon 499 -3338 499 -3338 0 3
rlabel polysilicon 506 -3332 506 -3332 0 1
rlabel polysilicon 506 -3338 506 -3338 0 3
rlabel polysilicon 513 -3332 513 -3332 0 1
rlabel polysilicon 513 -3338 513 -3338 0 3
rlabel polysilicon 520 -3332 520 -3332 0 1
rlabel polysilicon 520 -3338 520 -3338 0 3
rlabel polysilicon 527 -3332 527 -3332 0 1
rlabel polysilicon 527 -3338 527 -3338 0 3
rlabel polysilicon 534 -3332 534 -3332 0 1
rlabel polysilicon 534 -3338 534 -3338 0 3
rlabel polysilicon 541 -3332 541 -3332 0 1
rlabel polysilicon 544 -3338 544 -3338 0 4
rlabel polysilicon 548 -3332 548 -3332 0 1
rlabel polysilicon 548 -3338 548 -3338 0 3
rlabel polysilicon 555 -3332 555 -3332 0 1
rlabel polysilicon 555 -3338 555 -3338 0 3
rlabel polysilicon 562 -3332 562 -3332 0 1
rlabel polysilicon 562 -3338 562 -3338 0 3
rlabel polysilicon 572 -3332 572 -3332 0 2
rlabel polysilicon 569 -3338 569 -3338 0 3
rlabel polysilicon 572 -3338 572 -3338 0 4
rlabel polysilicon 576 -3332 576 -3332 0 1
rlabel polysilicon 576 -3338 576 -3338 0 3
rlabel polysilicon 583 -3332 583 -3332 0 1
rlabel polysilicon 583 -3338 583 -3338 0 3
rlabel polysilicon 590 -3332 590 -3332 0 1
rlabel polysilicon 593 -3332 593 -3332 0 2
rlabel polysilicon 593 -3338 593 -3338 0 4
rlabel polysilicon 597 -3332 597 -3332 0 1
rlabel polysilicon 597 -3338 597 -3338 0 3
rlabel polysilicon 604 -3332 604 -3332 0 1
rlabel polysilicon 604 -3338 604 -3338 0 3
rlabel polysilicon 611 -3332 611 -3332 0 1
rlabel polysilicon 611 -3338 611 -3338 0 3
rlabel polysilicon 618 -3332 618 -3332 0 1
rlabel polysilicon 618 -3338 618 -3338 0 3
rlabel polysilicon 621 -3338 621 -3338 0 4
rlabel polysilicon 625 -3332 625 -3332 0 1
rlabel polysilicon 625 -3338 625 -3338 0 3
rlabel polysilicon 632 -3332 632 -3332 0 1
rlabel polysilicon 632 -3338 632 -3338 0 3
rlabel polysilicon 639 -3332 639 -3332 0 1
rlabel polysilicon 639 -3338 639 -3338 0 3
rlabel polysilicon 646 -3332 646 -3332 0 1
rlabel polysilicon 646 -3338 646 -3338 0 3
rlabel polysilicon 653 -3332 653 -3332 0 1
rlabel polysilicon 653 -3338 653 -3338 0 3
rlabel polysilicon 660 -3332 660 -3332 0 1
rlabel polysilicon 660 -3338 660 -3338 0 3
rlabel polysilicon 667 -3332 667 -3332 0 1
rlabel polysilicon 670 -3332 670 -3332 0 2
rlabel polysilicon 667 -3338 667 -3338 0 3
rlabel polysilicon 674 -3332 674 -3332 0 1
rlabel polysilicon 674 -3338 674 -3338 0 3
rlabel polysilicon 681 -3332 681 -3332 0 1
rlabel polysilicon 684 -3332 684 -3332 0 2
rlabel polysilicon 681 -3338 681 -3338 0 3
rlabel polysilicon 688 -3332 688 -3332 0 1
rlabel polysilicon 688 -3338 688 -3338 0 3
rlabel polysilicon 695 -3332 695 -3332 0 1
rlabel polysilicon 695 -3338 695 -3338 0 3
rlabel polysilicon 702 -3332 702 -3332 0 1
rlabel polysilicon 702 -3338 702 -3338 0 3
rlabel polysilicon 709 -3332 709 -3332 0 1
rlabel polysilicon 712 -3332 712 -3332 0 2
rlabel polysilicon 709 -3338 709 -3338 0 3
rlabel polysilicon 712 -3338 712 -3338 0 4
rlabel polysilicon 716 -3332 716 -3332 0 1
rlabel polysilicon 716 -3338 716 -3338 0 3
rlabel polysilicon 723 -3332 723 -3332 0 1
rlabel polysilicon 723 -3338 723 -3338 0 3
rlabel polysilicon 730 -3332 730 -3332 0 1
rlabel polysilicon 730 -3338 730 -3338 0 3
rlabel polysilicon 737 -3332 737 -3332 0 1
rlabel polysilicon 737 -3338 737 -3338 0 3
rlabel polysilicon 740 -3338 740 -3338 0 4
rlabel polysilicon 744 -3332 744 -3332 0 1
rlabel polysilicon 744 -3338 744 -3338 0 3
rlabel polysilicon 751 -3332 751 -3332 0 1
rlabel polysilicon 751 -3338 751 -3338 0 3
rlabel polysilicon 758 -3332 758 -3332 0 1
rlabel polysilicon 758 -3338 758 -3338 0 3
rlabel polysilicon 765 -3332 765 -3332 0 1
rlabel polysilicon 765 -3338 765 -3338 0 3
rlabel polysilicon 772 -3332 772 -3332 0 1
rlabel polysilicon 772 -3338 772 -3338 0 3
rlabel polysilicon 779 -3332 779 -3332 0 1
rlabel polysilicon 779 -3338 779 -3338 0 3
rlabel polysilicon 786 -3332 786 -3332 0 1
rlabel polysilicon 786 -3338 786 -3338 0 3
rlabel polysilicon 793 -3332 793 -3332 0 1
rlabel polysilicon 793 -3338 793 -3338 0 3
rlabel polysilicon 800 -3332 800 -3332 0 1
rlabel polysilicon 800 -3338 800 -3338 0 3
rlabel polysilicon 807 -3332 807 -3332 0 1
rlabel polysilicon 807 -3338 807 -3338 0 3
rlabel polysilicon 814 -3332 814 -3332 0 1
rlabel polysilicon 814 -3338 814 -3338 0 3
rlabel polysilicon 821 -3332 821 -3332 0 1
rlabel polysilicon 821 -3338 821 -3338 0 3
rlabel polysilicon 828 -3332 828 -3332 0 1
rlabel polysilicon 828 -3338 828 -3338 0 3
rlabel polysilicon 835 -3332 835 -3332 0 1
rlabel polysilicon 838 -3332 838 -3332 0 2
rlabel polysilicon 842 -3332 842 -3332 0 1
rlabel polysilicon 845 -3332 845 -3332 0 2
rlabel polysilicon 842 -3338 842 -3338 0 3
rlabel polysilicon 845 -3338 845 -3338 0 4
rlabel polysilicon 849 -3332 849 -3332 0 1
rlabel polysilicon 849 -3338 849 -3338 0 3
rlabel polysilicon 856 -3332 856 -3332 0 1
rlabel polysilicon 856 -3338 856 -3338 0 3
rlabel polysilicon 863 -3332 863 -3332 0 1
rlabel polysilicon 863 -3338 863 -3338 0 3
rlabel polysilicon 870 -3332 870 -3332 0 1
rlabel polysilicon 870 -3338 870 -3338 0 3
rlabel polysilicon 877 -3332 877 -3332 0 1
rlabel polysilicon 877 -3338 877 -3338 0 3
rlabel polysilicon 884 -3332 884 -3332 0 1
rlabel polysilicon 884 -3338 884 -3338 0 3
rlabel polysilicon 891 -3332 891 -3332 0 1
rlabel polysilicon 891 -3338 891 -3338 0 3
rlabel polysilicon 898 -3332 898 -3332 0 1
rlabel polysilicon 898 -3338 898 -3338 0 3
rlabel polysilicon 905 -3332 905 -3332 0 1
rlabel polysilicon 905 -3338 905 -3338 0 3
rlabel polysilicon 912 -3332 912 -3332 0 1
rlabel polysilicon 912 -3338 912 -3338 0 3
rlabel polysilicon 919 -3332 919 -3332 0 1
rlabel polysilicon 919 -3338 919 -3338 0 3
rlabel polysilicon 926 -3332 926 -3332 0 1
rlabel polysilicon 926 -3338 926 -3338 0 3
rlabel polysilicon 933 -3332 933 -3332 0 1
rlabel polysilicon 936 -3332 936 -3332 0 2
rlabel polysilicon 933 -3338 933 -3338 0 3
rlabel polysilicon 936 -3338 936 -3338 0 4
rlabel polysilicon 940 -3332 940 -3332 0 1
rlabel polysilicon 940 -3338 940 -3338 0 3
rlabel polysilicon 947 -3338 947 -3338 0 3
rlabel polysilicon 954 -3332 954 -3332 0 1
rlabel polysilicon 954 -3338 954 -3338 0 3
rlabel polysilicon 961 -3332 961 -3332 0 1
rlabel polysilicon 961 -3338 961 -3338 0 3
rlabel polysilicon 975 -3332 975 -3332 0 1
rlabel polysilicon 975 -3338 975 -3338 0 3
rlabel polysilicon 989 -3332 989 -3332 0 1
rlabel polysilicon 989 -3338 989 -3338 0 3
rlabel polysilicon 1059 -3332 1059 -3332 0 1
rlabel polysilicon 1059 -3338 1059 -3338 0 3
rlabel polysilicon 1062 -3338 1062 -3338 0 4
rlabel polysilicon 1066 -3332 1066 -3332 0 1
rlabel polysilicon 1066 -3338 1066 -3338 0 3
rlabel polysilicon 1073 -3332 1073 -3332 0 1
rlabel polysilicon 1073 -3338 1073 -3338 0 3
rlabel polysilicon 1080 -3332 1080 -3332 0 1
rlabel polysilicon 1080 -3338 1080 -3338 0 3
rlabel polysilicon 1094 -3332 1094 -3332 0 1
rlabel polysilicon 1097 -3332 1097 -3332 0 2
rlabel polysilicon 1097 -3338 1097 -3338 0 4
rlabel polysilicon 1108 -3332 1108 -3332 0 1
rlabel polysilicon 1108 -3338 1108 -3338 0 3
rlabel polysilicon 1115 -3332 1115 -3332 0 1
rlabel polysilicon 1115 -3338 1115 -3338 0 3
rlabel polysilicon 1136 -3332 1136 -3332 0 1
rlabel polysilicon 1139 -3338 1139 -3338 0 4
rlabel polysilicon 1143 -3332 1143 -3332 0 1
rlabel polysilicon 1143 -3338 1143 -3338 0 3
rlabel polysilicon 1213 -3332 1213 -3332 0 1
rlabel polysilicon 1213 -3338 1213 -3338 0 3
rlabel polysilicon 1290 -3332 1290 -3332 0 1
rlabel polysilicon 1290 -3338 1290 -3338 0 3
rlabel polysilicon 1360 -3332 1360 -3332 0 1
rlabel polysilicon 1360 -3338 1360 -3338 0 3
rlabel polysilicon 1367 -3332 1367 -3332 0 1
rlabel polysilicon 1367 -3338 1367 -3338 0 3
rlabel polysilicon 1409 -3332 1409 -3332 0 1
rlabel polysilicon 1409 -3338 1409 -3338 0 3
rlabel polysilicon 177 -3397 177 -3397 0 1
rlabel polysilicon 177 -3403 177 -3403 0 3
rlabel polysilicon 184 -3397 184 -3397 0 1
rlabel polysilicon 184 -3403 184 -3403 0 3
rlabel polysilicon 191 -3397 191 -3397 0 1
rlabel polysilicon 191 -3403 191 -3403 0 3
rlabel polysilicon 198 -3397 198 -3397 0 1
rlabel polysilicon 198 -3403 198 -3403 0 3
rlabel polysilicon 205 -3397 205 -3397 0 1
rlabel polysilicon 205 -3403 205 -3403 0 3
rlabel polysilicon 212 -3397 212 -3397 0 1
rlabel polysilicon 212 -3403 212 -3403 0 3
rlabel polysilicon 219 -3397 219 -3397 0 1
rlabel polysilicon 219 -3403 219 -3403 0 3
rlabel polysilicon 226 -3397 226 -3397 0 1
rlabel polysilicon 229 -3397 229 -3397 0 2
rlabel polysilicon 226 -3403 226 -3403 0 3
rlabel polysilicon 229 -3403 229 -3403 0 4
rlabel polysilicon 233 -3403 233 -3403 0 3
rlabel polysilicon 240 -3397 240 -3397 0 1
rlabel polysilicon 240 -3403 240 -3403 0 3
rlabel polysilicon 247 -3397 247 -3397 0 1
rlabel polysilicon 247 -3403 247 -3403 0 3
rlabel polysilicon 254 -3397 254 -3397 0 1
rlabel polysilicon 254 -3403 254 -3403 0 3
rlabel polysilicon 261 -3397 261 -3397 0 1
rlabel polysilicon 261 -3403 261 -3403 0 3
rlabel polysilicon 268 -3397 268 -3397 0 1
rlabel polysilicon 268 -3403 268 -3403 0 3
rlabel polysilicon 275 -3397 275 -3397 0 1
rlabel polysilicon 275 -3403 275 -3403 0 3
rlabel polysilicon 282 -3397 282 -3397 0 1
rlabel polysilicon 282 -3403 282 -3403 0 3
rlabel polysilicon 289 -3397 289 -3397 0 1
rlabel polysilicon 289 -3403 289 -3403 0 3
rlabel polysilicon 296 -3397 296 -3397 0 1
rlabel polysilicon 296 -3403 296 -3403 0 3
rlabel polysilicon 303 -3397 303 -3397 0 1
rlabel polysilicon 306 -3397 306 -3397 0 2
rlabel polysilicon 303 -3403 303 -3403 0 3
rlabel polysilicon 310 -3397 310 -3397 0 1
rlabel polysilicon 310 -3403 310 -3403 0 3
rlabel polysilicon 317 -3397 317 -3397 0 1
rlabel polysilicon 317 -3403 317 -3403 0 3
rlabel polysilicon 324 -3397 324 -3397 0 1
rlabel polysilicon 324 -3403 324 -3403 0 3
rlabel polysilicon 331 -3397 331 -3397 0 1
rlabel polysilicon 331 -3403 331 -3403 0 3
rlabel polysilicon 341 -3403 341 -3403 0 4
rlabel polysilicon 345 -3397 345 -3397 0 1
rlabel polysilicon 345 -3403 345 -3403 0 3
rlabel polysilicon 352 -3397 352 -3397 0 1
rlabel polysilicon 355 -3397 355 -3397 0 2
rlabel polysilicon 355 -3403 355 -3403 0 4
rlabel polysilicon 359 -3397 359 -3397 0 1
rlabel polysilicon 359 -3403 359 -3403 0 3
rlabel polysilicon 366 -3397 366 -3397 0 1
rlabel polysilicon 366 -3403 366 -3403 0 3
rlabel polysilicon 373 -3397 373 -3397 0 1
rlabel polysilicon 373 -3403 373 -3403 0 3
rlabel polysilicon 380 -3397 380 -3397 0 1
rlabel polysilicon 383 -3403 383 -3403 0 4
rlabel polysilicon 387 -3397 387 -3397 0 1
rlabel polysilicon 387 -3403 387 -3403 0 3
rlabel polysilicon 394 -3397 394 -3397 0 1
rlabel polysilicon 397 -3397 397 -3397 0 2
rlabel polysilicon 394 -3403 394 -3403 0 3
rlabel polysilicon 401 -3397 401 -3397 0 1
rlabel polysilicon 401 -3403 401 -3403 0 3
rlabel polysilicon 408 -3397 408 -3397 0 1
rlabel polysilicon 408 -3403 408 -3403 0 3
rlabel polysilicon 415 -3397 415 -3397 0 1
rlabel polysilicon 415 -3403 415 -3403 0 3
rlabel polysilicon 422 -3397 422 -3397 0 1
rlabel polysilicon 422 -3403 422 -3403 0 3
rlabel polysilicon 429 -3397 429 -3397 0 1
rlabel polysilicon 429 -3403 429 -3403 0 3
rlabel polysilicon 436 -3397 436 -3397 0 1
rlabel polysilicon 436 -3403 436 -3403 0 3
rlabel polysilicon 443 -3397 443 -3397 0 1
rlabel polysilicon 443 -3403 443 -3403 0 3
rlabel polysilicon 450 -3397 450 -3397 0 1
rlabel polysilicon 450 -3403 450 -3403 0 3
rlabel polysilicon 457 -3397 457 -3397 0 1
rlabel polysilicon 457 -3403 457 -3403 0 3
rlabel polysilicon 464 -3397 464 -3397 0 1
rlabel polysilicon 467 -3403 467 -3403 0 4
rlabel polysilicon 471 -3397 471 -3397 0 1
rlabel polysilicon 471 -3403 471 -3403 0 3
rlabel polysilicon 478 -3397 478 -3397 0 1
rlabel polysilicon 478 -3403 478 -3403 0 3
rlabel polysilicon 485 -3397 485 -3397 0 1
rlabel polysilicon 488 -3397 488 -3397 0 2
rlabel polysilicon 488 -3403 488 -3403 0 4
rlabel polysilicon 495 -3397 495 -3397 0 2
rlabel polysilicon 495 -3403 495 -3403 0 4
rlabel polysilicon 499 -3397 499 -3397 0 1
rlabel polysilicon 499 -3403 499 -3403 0 3
rlabel polysilicon 506 -3403 506 -3403 0 3
rlabel polysilicon 513 -3397 513 -3397 0 1
rlabel polysilicon 513 -3403 513 -3403 0 3
rlabel polysilicon 520 -3397 520 -3397 0 1
rlabel polysilicon 520 -3403 520 -3403 0 3
rlabel polysilicon 527 -3397 527 -3397 0 1
rlabel polysilicon 527 -3403 527 -3403 0 3
rlabel polysilicon 534 -3397 534 -3397 0 1
rlabel polysilicon 537 -3397 537 -3397 0 2
rlabel polysilicon 534 -3403 534 -3403 0 3
rlabel polysilicon 541 -3397 541 -3397 0 1
rlabel polysilicon 541 -3403 541 -3403 0 3
rlabel polysilicon 548 -3397 548 -3397 0 1
rlabel polysilicon 548 -3403 548 -3403 0 3
rlabel polysilicon 558 -3397 558 -3397 0 2
rlabel polysilicon 558 -3403 558 -3403 0 4
rlabel polysilicon 562 -3397 562 -3397 0 1
rlabel polysilicon 562 -3403 562 -3403 0 3
rlabel polysilicon 569 -3397 569 -3397 0 1
rlabel polysilicon 569 -3403 569 -3403 0 3
rlabel polysilicon 576 -3397 576 -3397 0 1
rlabel polysilicon 576 -3403 576 -3403 0 3
rlabel polysilicon 583 -3397 583 -3397 0 1
rlabel polysilicon 583 -3403 583 -3403 0 3
rlabel polysilicon 590 -3397 590 -3397 0 1
rlabel polysilicon 590 -3403 590 -3403 0 3
rlabel polysilicon 597 -3397 597 -3397 0 1
rlabel polysilicon 597 -3403 597 -3403 0 3
rlabel polysilicon 604 -3397 604 -3397 0 1
rlabel polysilicon 604 -3403 604 -3403 0 3
rlabel polysilicon 611 -3397 611 -3397 0 1
rlabel polysilicon 611 -3403 611 -3403 0 3
rlabel polysilicon 618 -3397 618 -3397 0 1
rlabel polysilicon 618 -3403 618 -3403 0 3
rlabel polysilicon 625 -3397 625 -3397 0 1
rlabel polysilicon 625 -3403 625 -3403 0 3
rlabel polysilicon 632 -3397 632 -3397 0 1
rlabel polysilicon 632 -3403 632 -3403 0 3
rlabel polysilicon 639 -3397 639 -3397 0 1
rlabel polysilicon 639 -3403 639 -3403 0 3
rlabel polysilicon 646 -3397 646 -3397 0 1
rlabel polysilicon 646 -3403 646 -3403 0 3
rlabel polysilicon 653 -3397 653 -3397 0 1
rlabel polysilicon 653 -3403 653 -3403 0 3
rlabel polysilicon 660 -3397 660 -3397 0 1
rlabel polysilicon 660 -3403 660 -3403 0 3
rlabel polysilicon 667 -3397 667 -3397 0 1
rlabel polysilicon 674 -3397 674 -3397 0 1
rlabel polysilicon 674 -3403 674 -3403 0 3
rlabel polysilicon 681 -3397 681 -3397 0 1
rlabel polysilicon 681 -3403 681 -3403 0 3
rlabel polysilicon 688 -3397 688 -3397 0 1
rlabel polysilicon 688 -3403 688 -3403 0 3
rlabel polysilicon 695 -3397 695 -3397 0 1
rlabel polysilicon 695 -3403 695 -3403 0 3
rlabel polysilicon 702 -3397 702 -3397 0 1
rlabel polysilicon 709 -3397 709 -3397 0 1
rlabel polysilicon 709 -3403 709 -3403 0 3
rlabel polysilicon 716 -3397 716 -3397 0 1
rlabel polysilicon 716 -3403 716 -3403 0 3
rlabel polysilicon 723 -3397 723 -3397 0 1
rlabel polysilicon 723 -3403 723 -3403 0 3
rlabel polysilicon 730 -3397 730 -3397 0 1
rlabel polysilicon 730 -3403 730 -3403 0 3
rlabel polysilicon 733 -3403 733 -3403 0 4
rlabel polysilicon 737 -3397 737 -3397 0 1
rlabel polysilicon 737 -3403 737 -3403 0 3
rlabel polysilicon 744 -3397 744 -3397 0 1
rlabel polysilicon 744 -3403 744 -3403 0 3
rlabel polysilicon 751 -3397 751 -3397 0 1
rlabel polysilicon 751 -3403 751 -3403 0 3
rlabel polysilicon 758 -3397 758 -3397 0 1
rlabel polysilicon 758 -3403 758 -3403 0 3
rlabel polysilicon 765 -3397 765 -3397 0 1
rlabel polysilicon 765 -3403 765 -3403 0 3
rlabel polysilicon 775 -3397 775 -3397 0 2
rlabel polysilicon 772 -3403 772 -3403 0 3
rlabel polysilicon 775 -3403 775 -3403 0 4
rlabel polysilicon 779 -3397 779 -3397 0 1
rlabel polysilicon 779 -3403 779 -3403 0 3
rlabel polysilicon 814 -3397 814 -3397 0 1
rlabel polysilicon 814 -3403 814 -3403 0 3
rlabel polysilicon 821 -3397 821 -3397 0 1
rlabel polysilicon 821 -3403 821 -3403 0 3
rlabel polysilicon 828 -3397 828 -3397 0 1
rlabel polysilicon 831 -3397 831 -3397 0 2
rlabel polysilicon 835 -3397 835 -3397 0 1
rlabel polysilicon 835 -3403 835 -3403 0 3
rlabel polysilicon 845 -3397 845 -3397 0 2
rlabel polysilicon 842 -3403 842 -3403 0 3
rlabel polysilicon 845 -3403 845 -3403 0 4
rlabel polysilicon 849 -3397 849 -3397 0 1
rlabel polysilicon 849 -3403 849 -3403 0 3
rlabel polysilicon 856 -3397 856 -3397 0 1
rlabel polysilicon 856 -3403 856 -3403 0 3
rlabel polysilicon 863 -3397 863 -3397 0 1
rlabel polysilicon 866 -3397 866 -3397 0 2
rlabel polysilicon 863 -3403 863 -3403 0 3
rlabel polysilicon 870 -3397 870 -3397 0 1
rlabel polysilicon 870 -3403 870 -3403 0 3
rlabel polysilicon 877 -3397 877 -3397 0 1
rlabel polysilicon 877 -3403 877 -3403 0 3
rlabel polysilicon 884 -3397 884 -3397 0 1
rlabel polysilicon 884 -3403 884 -3403 0 3
rlabel polysilicon 894 -3397 894 -3397 0 2
rlabel polysilicon 891 -3403 891 -3403 0 3
rlabel polysilicon 905 -3397 905 -3397 0 1
rlabel polysilicon 905 -3403 905 -3403 0 3
rlabel polysilicon 912 -3397 912 -3397 0 1
rlabel polysilicon 912 -3403 912 -3403 0 3
rlabel polysilicon 919 -3397 919 -3397 0 1
rlabel polysilicon 919 -3403 919 -3403 0 3
rlabel polysilicon 926 -3397 926 -3397 0 1
rlabel polysilicon 926 -3403 926 -3403 0 3
rlabel polysilicon 940 -3397 940 -3397 0 1
rlabel polysilicon 940 -3403 940 -3403 0 3
rlabel polysilicon 989 -3397 989 -3397 0 1
rlabel polysilicon 989 -3403 989 -3403 0 3
rlabel polysilicon 996 -3397 996 -3397 0 1
rlabel polysilicon 996 -3403 996 -3403 0 3
rlabel polysilicon 1073 -3397 1073 -3397 0 1
rlabel polysilicon 1073 -3403 1073 -3403 0 3
rlabel polysilicon 1115 -3397 1115 -3397 0 1
rlabel polysilicon 1115 -3403 1115 -3403 0 3
rlabel polysilicon 1122 -3397 1122 -3397 0 1
rlabel polysilicon 1122 -3403 1122 -3403 0 3
rlabel polysilicon 1213 -3397 1213 -3397 0 1
rlabel polysilicon 1213 -3403 1213 -3403 0 3
rlabel polysilicon 1353 -3397 1353 -3397 0 1
rlabel polysilicon 1353 -3403 1353 -3403 0 3
rlabel polysilicon 1360 -3397 1360 -3397 0 1
rlabel polysilicon 1360 -3403 1360 -3403 0 3
rlabel polysilicon 1367 -3397 1367 -3397 0 1
rlabel polysilicon 1367 -3403 1367 -3403 0 3
rlabel polysilicon 1409 -3397 1409 -3397 0 1
rlabel polysilicon 1409 -3403 1409 -3403 0 3
rlabel polysilicon 222 -3440 222 -3440 0 2
rlabel polysilicon 222 -3446 222 -3446 0 4
rlabel polysilicon 240 -3440 240 -3440 0 1
rlabel polysilicon 240 -3446 240 -3446 0 3
rlabel polysilicon 254 -3440 254 -3440 0 1
rlabel polysilicon 254 -3446 254 -3446 0 3
rlabel polysilicon 264 -3440 264 -3440 0 2
rlabel polysilicon 264 -3446 264 -3446 0 4
rlabel polysilicon 268 -3440 268 -3440 0 1
rlabel polysilicon 268 -3446 268 -3446 0 3
rlabel polysilicon 275 -3440 275 -3440 0 1
rlabel polysilicon 275 -3446 275 -3446 0 3
rlabel polysilicon 282 -3440 282 -3440 0 1
rlabel polysilicon 282 -3446 282 -3446 0 3
rlabel polysilicon 289 -3446 289 -3446 0 3
rlabel polysilicon 292 -3446 292 -3446 0 4
rlabel polysilicon 296 -3440 296 -3440 0 1
rlabel polysilicon 296 -3446 296 -3446 0 3
rlabel polysilicon 303 -3440 303 -3440 0 1
rlabel polysilicon 306 -3446 306 -3446 0 4
rlabel polysilicon 310 -3440 310 -3440 0 1
rlabel polysilicon 310 -3446 310 -3446 0 3
rlabel polysilicon 317 -3440 317 -3440 0 1
rlabel polysilicon 317 -3446 317 -3446 0 3
rlabel polysilicon 324 -3440 324 -3440 0 1
rlabel polysilicon 327 -3440 327 -3440 0 2
rlabel polysilicon 327 -3446 327 -3446 0 4
rlabel polysilicon 338 -3440 338 -3440 0 1
rlabel polysilicon 341 -3440 341 -3440 0 2
rlabel polysilicon 345 -3440 345 -3440 0 1
rlabel polysilicon 345 -3446 345 -3446 0 3
rlabel polysilicon 352 -3440 352 -3440 0 1
rlabel polysilicon 352 -3446 352 -3446 0 3
rlabel polysilicon 359 -3440 359 -3440 0 1
rlabel polysilicon 359 -3446 359 -3446 0 3
rlabel polysilicon 373 -3440 373 -3440 0 1
rlabel polysilicon 373 -3446 373 -3446 0 3
rlabel polysilicon 387 -3440 387 -3440 0 1
rlabel polysilicon 387 -3446 387 -3446 0 3
rlabel polysilicon 394 -3440 394 -3440 0 1
rlabel polysilicon 394 -3446 394 -3446 0 3
rlabel polysilicon 401 -3440 401 -3440 0 1
rlabel polysilicon 401 -3446 401 -3446 0 3
rlabel polysilicon 408 -3440 408 -3440 0 1
rlabel polysilicon 408 -3446 408 -3446 0 3
rlabel polysilicon 422 -3440 422 -3440 0 1
rlabel polysilicon 422 -3446 422 -3446 0 3
rlabel polysilicon 429 -3440 429 -3440 0 1
rlabel polysilicon 429 -3446 429 -3446 0 3
rlabel polysilicon 436 -3440 436 -3440 0 1
rlabel polysilicon 436 -3446 436 -3446 0 3
rlabel polysilicon 443 -3440 443 -3440 0 1
rlabel polysilicon 443 -3446 443 -3446 0 3
rlabel polysilicon 450 -3440 450 -3440 0 1
rlabel polysilicon 450 -3446 450 -3446 0 3
rlabel polysilicon 471 -3440 471 -3440 0 1
rlabel polysilicon 471 -3446 471 -3446 0 3
rlabel polysilicon 485 -3440 485 -3440 0 1
rlabel polysilicon 485 -3446 485 -3446 0 3
rlabel polysilicon 492 -3440 492 -3440 0 1
rlabel polysilicon 492 -3446 492 -3446 0 3
rlabel polysilicon 499 -3440 499 -3440 0 1
rlabel polysilicon 502 -3446 502 -3446 0 4
rlabel polysilicon 534 -3440 534 -3440 0 1
rlabel polysilicon 534 -3446 534 -3446 0 3
rlabel polysilicon 541 -3440 541 -3440 0 1
rlabel polysilicon 541 -3446 541 -3446 0 3
rlabel polysilicon 548 -3440 548 -3440 0 1
rlabel polysilicon 548 -3446 548 -3446 0 3
rlabel polysilicon 555 -3440 555 -3440 0 1
rlabel polysilicon 555 -3446 555 -3446 0 3
rlabel polysilicon 562 -3440 562 -3440 0 1
rlabel polysilicon 562 -3446 562 -3446 0 3
rlabel polysilicon 569 -3440 569 -3440 0 1
rlabel polysilicon 569 -3446 569 -3446 0 3
rlabel polysilicon 572 -3446 572 -3446 0 4
rlabel polysilicon 576 -3440 576 -3440 0 1
rlabel polysilicon 576 -3446 576 -3446 0 3
rlabel polysilicon 583 -3440 583 -3440 0 1
rlabel polysilicon 583 -3446 583 -3446 0 3
rlabel polysilicon 597 -3440 597 -3440 0 1
rlabel polysilicon 597 -3446 597 -3446 0 3
rlabel polysilicon 625 -3440 625 -3440 0 1
rlabel polysilicon 625 -3446 625 -3446 0 3
rlabel polysilicon 632 -3440 632 -3440 0 1
rlabel polysilicon 632 -3446 632 -3446 0 3
rlabel polysilicon 639 -3440 639 -3440 0 1
rlabel polysilicon 642 -3440 642 -3440 0 2
rlabel polysilicon 639 -3446 639 -3446 0 3
rlabel polysilicon 642 -3446 642 -3446 0 4
rlabel polysilicon 646 -3440 646 -3440 0 1
rlabel polysilicon 646 -3446 646 -3446 0 3
rlabel polysilicon 653 -3440 653 -3440 0 1
rlabel polysilicon 653 -3446 653 -3446 0 3
rlabel polysilicon 660 -3440 660 -3440 0 1
rlabel polysilicon 660 -3446 660 -3446 0 3
rlabel polysilicon 667 -3446 667 -3446 0 3
rlabel polysilicon 674 -3440 674 -3440 0 1
rlabel polysilicon 674 -3446 674 -3446 0 3
rlabel polysilicon 681 -3440 681 -3440 0 1
rlabel polysilicon 681 -3446 681 -3446 0 3
rlabel polysilicon 688 -3440 688 -3440 0 1
rlabel polysilicon 688 -3446 688 -3446 0 3
rlabel polysilicon 695 -3440 695 -3440 0 1
rlabel polysilicon 695 -3446 695 -3446 0 3
rlabel polysilicon 702 -3440 702 -3440 0 1
rlabel polysilicon 702 -3446 702 -3446 0 3
rlabel polysilicon 709 -3440 709 -3440 0 1
rlabel polysilicon 709 -3446 709 -3446 0 3
rlabel polysilicon 719 -3440 719 -3440 0 2
rlabel polysilicon 716 -3446 716 -3446 0 3
rlabel polysilicon 719 -3446 719 -3446 0 4
rlabel polysilicon 723 -3440 723 -3440 0 1
rlabel polysilicon 723 -3446 723 -3446 0 3
rlabel polysilicon 726 -3446 726 -3446 0 4
rlabel polysilicon 730 -3440 730 -3440 0 1
rlabel polysilicon 733 -3440 733 -3440 0 2
rlabel polysilicon 730 -3446 730 -3446 0 3
rlabel polysilicon 737 -3446 737 -3446 0 3
rlabel polysilicon 740 -3446 740 -3446 0 4
rlabel polysilicon 744 -3440 744 -3440 0 1
rlabel polysilicon 744 -3446 744 -3446 0 3
rlabel polysilicon 751 -3440 751 -3440 0 1
rlabel polysilicon 751 -3446 751 -3446 0 3
rlabel polysilicon 758 -3440 758 -3440 0 1
rlabel polysilicon 758 -3446 758 -3446 0 3
rlabel polysilicon 765 -3440 765 -3440 0 1
rlabel polysilicon 765 -3446 765 -3446 0 3
rlabel polysilicon 772 -3440 772 -3440 0 1
rlabel polysilicon 779 -3440 779 -3440 0 1
rlabel polysilicon 782 -3440 782 -3440 0 2
rlabel polysilicon 779 -3446 779 -3446 0 3
rlabel polysilicon 782 -3446 782 -3446 0 4
rlabel polysilicon 821 -3440 821 -3440 0 1
rlabel polysilicon 821 -3446 821 -3446 0 3
rlabel polysilicon 831 -3440 831 -3440 0 2
rlabel polysilicon 828 -3446 828 -3446 0 3
rlabel polysilicon 831 -3446 831 -3446 0 4
rlabel polysilicon 835 -3440 835 -3440 0 1
rlabel polysilicon 835 -3446 835 -3446 0 3
rlabel polysilicon 842 -3440 842 -3440 0 1
rlabel polysilicon 842 -3446 842 -3446 0 3
rlabel polysilicon 849 -3440 849 -3440 0 1
rlabel polysilicon 849 -3446 849 -3446 0 3
rlabel polysilicon 856 -3440 856 -3440 0 1
rlabel polysilicon 856 -3446 856 -3446 0 3
rlabel polysilicon 863 -3440 863 -3440 0 1
rlabel polysilicon 863 -3446 863 -3446 0 3
rlabel polysilicon 870 -3440 870 -3440 0 1
rlabel polysilicon 870 -3446 870 -3446 0 3
rlabel polysilicon 884 -3440 884 -3440 0 1
rlabel polysilicon 884 -3446 884 -3446 0 3
rlabel polysilicon 912 -3440 912 -3440 0 1
rlabel polysilicon 912 -3446 912 -3446 0 3
rlabel polysilicon 919 -3440 919 -3440 0 1
rlabel polysilicon 919 -3446 919 -3446 0 3
rlabel polysilicon 926 -3440 926 -3440 0 1
rlabel polysilicon 926 -3446 926 -3446 0 3
rlabel polysilicon 940 -3440 940 -3440 0 1
rlabel polysilicon 940 -3446 940 -3446 0 3
rlabel polysilicon 947 -3440 947 -3440 0 1
rlabel polysilicon 947 -3446 947 -3446 0 3
rlabel polysilicon 954 -3440 954 -3440 0 1
rlabel polysilicon 954 -3446 954 -3446 0 3
rlabel polysilicon 957 -3446 957 -3446 0 4
rlabel polysilicon 961 -3440 961 -3440 0 1
rlabel polysilicon 964 -3440 964 -3440 0 2
rlabel polysilicon 961 -3446 961 -3446 0 3
rlabel polysilicon 964 -3446 964 -3446 0 4
rlabel polysilicon 968 -3440 968 -3440 0 1
rlabel polysilicon 968 -3446 968 -3446 0 3
rlabel polysilicon 975 -3440 975 -3440 0 1
rlabel polysilicon 975 -3446 975 -3446 0 3
rlabel polysilicon 982 -3440 982 -3440 0 1
rlabel polysilicon 982 -3446 982 -3446 0 3
rlabel polysilicon 989 -3440 989 -3440 0 1
rlabel polysilicon 989 -3446 989 -3446 0 3
rlabel polysilicon 996 -3440 996 -3440 0 1
rlabel polysilicon 996 -3446 996 -3446 0 3
rlabel polysilicon 1010 -3440 1010 -3440 0 1
rlabel polysilicon 1010 -3446 1010 -3446 0 3
rlabel polysilicon 1073 -3440 1073 -3440 0 1
rlabel polysilicon 1073 -3446 1073 -3446 0 3
rlabel polysilicon 1094 -3440 1094 -3440 0 1
rlabel polysilicon 1094 -3446 1094 -3446 0 3
rlabel polysilicon 1115 -3440 1115 -3440 0 1
rlabel polysilicon 1115 -3446 1115 -3446 0 3
rlabel polysilicon 1122 -3440 1122 -3440 0 1
rlabel polysilicon 1122 -3446 1122 -3446 0 3
rlabel polysilicon 1213 -3440 1213 -3440 0 1
rlabel polysilicon 1213 -3446 1213 -3446 0 3
rlabel polysilicon 1353 -3440 1353 -3440 0 1
rlabel polysilicon 1353 -3446 1353 -3446 0 3
rlabel polysilicon 1360 -3440 1360 -3440 0 1
rlabel polysilicon 1360 -3446 1360 -3446 0 3
rlabel polysilicon 1395 -3440 1395 -3440 0 1
rlabel polysilicon 1395 -3446 1395 -3446 0 3
rlabel polysilicon 1409 -3440 1409 -3440 0 1
rlabel polysilicon 1409 -3446 1409 -3446 0 3
rlabel polysilicon 254 -3467 254 -3467 0 1
rlabel polysilicon 254 -3473 254 -3473 0 3
rlabel polysilicon 261 -3467 261 -3467 0 1
rlabel polysilicon 261 -3473 261 -3473 0 3
rlabel polysilicon 303 -3467 303 -3467 0 1
rlabel polysilicon 303 -3473 303 -3473 0 3
rlabel polysilicon 317 -3467 317 -3467 0 1
rlabel polysilicon 317 -3473 317 -3473 0 3
rlabel polysilicon 327 -3467 327 -3467 0 2
rlabel polysilicon 327 -3473 327 -3473 0 4
rlabel polysilicon 331 -3467 331 -3467 0 1
rlabel polysilicon 331 -3473 331 -3473 0 3
rlabel polysilicon 338 -3467 338 -3467 0 1
rlabel polysilicon 338 -3473 338 -3473 0 3
rlabel polysilicon 352 -3467 352 -3467 0 1
rlabel polysilicon 352 -3473 352 -3473 0 3
rlabel polysilicon 359 -3467 359 -3467 0 1
rlabel polysilicon 359 -3473 359 -3473 0 3
rlabel polysilicon 380 -3467 380 -3467 0 1
rlabel polysilicon 380 -3473 380 -3473 0 3
rlabel polysilicon 394 -3467 394 -3467 0 1
rlabel polysilicon 394 -3473 394 -3473 0 3
rlabel polysilicon 401 -3467 401 -3467 0 1
rlabel polysilicon 401 -3473 401 -3473 0 3
rlabel polysilicon 408 -3473 408 -3473 0 3
rlabel polysilicon 411 -3473 411 -3473 0 4
rlabel polysilicon 415 -3467 415 -3467 0 1
rlabel polysilicon 415 -3473 415 -3473 0 3
rlabel polysilicon 422 -3467 422 -3467 0 1
rlabel polysilicon 425 -3467 425 -3467 0 2
rlabel polysilicon 429 -3467 429 -3467 0 1
rlabel polysilicon 429 -3473 429 -3473 0 3
rlabel polysilicon 436 -3473 436 -3473 0 3
rlabel polysilicon 439 -3473 439 -3473 0 4
rlabel polysilicon 443 -3467 443 -3467 0 1
rlabel polysilicon 443 -3473 443 -3473 0 3
rlabel polysilicon 457 -3467 457 -3467 0 1
rlabel polysilicon 460 -3467 460 -3467 0 2
rlabel polysilicon 464 -3467 464 -3467 0 1
rlabel polysilicon 467 -3473 467 -3473 0 4
rlabel polysilicon 471 -3467 471 -3467 0 1
rlabel polysilicon 471 -3473 471 -3473 0 3
rlabel polysilicon 478 -3467 478 -3467 0 1
rlabel polysilicon 478 -3473 478 -3473 0 3
rlabel polysilicon 485 -3467 485 -3467 0 1
rlabel polysilicon 485 -3473 485 -3473 0 3
rlabel polysilicon 492 -3467 492 -3467 0 1
rlabel polysilicon 492 -3473 492 -3473 0 3
rlabel polysilicon 499 -3473 499 -3473 0 3
rlabel polysilicon 502 -3473 502 -3473 0 4
rlabel polysilicon 506 -3467 506 -3467 0 1
rlabel polysilicon 506 -3473 506 -3473 0 3
rlabel polysilicon 513 -3473 513 -3473 0 3
rlabel polysilicon 516 -3473 516 -3473 0 4
rlabel polysilicon 520 -3467 520 -3467 0 1
rlabel polysilicon 520 -3473 520 -3473 0 3
rlabel polysilicon 541 -3467 541 -3467 0 1
rlabel polysilicon 541 -3473 541 -3473 0 3
rlabel polysilicon 548 -3467 548 -3467 0 1
rlabel polysilicon 548 -3473 548 -3473 0 3
rlabel polysilicon 555 -3467 555 -3467 0 1
rlabel polysilicon 562 -3467 562 -3467 0 1
rlabel polysilicon 562 -3473 562 -3473 0 3
rlabel polysilicon 569 -3467 569 -3467 0 1
rlabel polysilicon 569 -3473 569 -3473 0 3
rlabel polysilicon 576 -3467 576 -3467 0 1
rlabel polysilicon 576 -3473 576 -3473 0 3
rlabel polysilicon 583 -3467 583 -3467 0 1
rlabel polysilicon 583 -3473 583 -3473 0 3
rlabel polysilicon 604 -3467 604 -3467 0 1
rlabel polysilicon 604 -3473 604 -3473 0 3
rlabel polysilicon 614 -3467 614 -3467 0 2
rlabel polysilicon 611 -3473 611 -3473 0 3
rlabel polysilicon 614 -3473 614 -3473 0 4
rlabel polysilicon 621 -3467 621 -3467 0 2
rlabel polysilicon 621 -3473 621 -3473 0 4
rlabel polysilicon 625 -3467 625 -3467 0 1
rlabel polysilicon 625 -3473 625 -3473 0 3
rlabel polysilicon 646 -3467 646 -3467 0 1
rlabel polysilicon 646 -3473 646 -3473 0 3
rlabel polysilicon 653 -3467 653 -3467 0 1
rlabel polysilicon 653 -3473 653 -3473 0 3
rlabel polysilicon 660 -3467 660 -3467 0 1
rlabel polysilicon 660 -3473 660 -3473 0 3
rlabel polysilicon 674 -3467 674 -3467 0 1
rlabel polysilicon 674 -3473 674 -3473 0 3
rlabel polysilicon 681 -3467 681 -3467 0 1
rlabel polysilicon 681 -3473 681 -3473 0 3
rlabel polysilicon 688 -3467 688 -3467 0 1
rlabel polysilicon 691 -3467 691 -3467 0 2
rlabel polysilicon 695 -3467 695 -3467 0 1
rlabel polysilicon 698 -3467 698 -3467 0 2
rlabel polysilicon 695 -3473 695 -3473 0 3
rlabel polysilicon 698 -3473 698 -3473 0 4
rlabel polysilicon 709 -3467 709 -3467 0 1
rlabel polysilicon 709 -3473 709 -3473 0 3
rlabel polysilicon 737 -3467 737 -3467 0 1
rlabel polysilicon 737 -3473 737 -3473 0 3
rlabel polysilicon 758 -3467 758 -3467 0 1
rlabel polysilicon 758 -3473 758 -3473 0 3
rlabel polysilicon 821 -3467 821 -3467 0 1
rlabel polysilicon 824 -3467 824 -3467 0 2
rlabel polysilicon 821 -3473 821 -3473 0 3
rlabel polysilicon 835 -3467 835 -3467 0 1
rlabel polysilicon 835 -3473 835 -3473 0 3
rlabel polysilicon 842 -3467 842 -3467 0 1
rlabel polysilicon 842 -3473 842 -3473 0 3
rlabel polysilicon 849 -3467 849 -3467 0 1
rlabel polysilicon 852 -3473 852 -3473 0 4
rlabel polysilicon 856 -3467 856 -3467 0 1
rlabel polysilicon 856 -3473 856 -3473 0 3
rlabel polysilicon 870 -3467 870 -3467 0 1
rlabel polysilicon 870 -3473 870 -3473 0 3
rlabel polysilicon 884 -3467 884 -3467 0 1
rlabel polysilicon 884 -3473 884 -3473 0 3
rlabel polysilicon 891 -3467 891 -3467 0 1
rlabel polysilicon 891 -3473 891 -3473 0 3
rlabel polysilicon 912 -3467 912 -3467 0 1
rlabel polysilicon 912 -3473 912 -3473 0 3
rlabel polysilicon 919 -3467 919 -3467 0 1
rlabel polysilicon 919 -3473 919 -3473 0 3
rlabel polysilicon 926 -3467 926 -3467 0 1
rlabel polysilicon 926 -3473 926 -3473 0 3
rlabel polysilicon 933 -3467 933 -3467 0 1
rlabel polysilicon 933 -3473 933 -3473 0 3
rlabel polysilicon 940 -3467 940 -3467 0 1
rlabel polysilicon 940 -3473 940 -3473 0 3
rlabel polysilicon 989 -3467 989 -3467 0 1
rlabel polysilicon 989 -3473 989 -3473 0 3
rlabel polysilicon 996 -3467 996 -3467 0 1
rlabel polysilicon 996 -3473 996 -3473 0 3
rlabel polysilicon 1066 -3467 1066 -3467 0 1
rlabel polysilicon 1066 -3473 1066 -3473 0 3
rlabel polysilicon 1073 -3467 1073 -3467 0 1
rlabel polysilicon 1076 -3467 1076 -3467 0 2
rlabel polysilicon 1115 -3467 1115 -3467 0 1
rlabel polysilicon 1115 -3473 1115 -3473 0 3
rlabel polysilicon 1122 -3467 1122 -3467 0 1
rlabel polysilicon 1122 -3473 1122 -3473 0 3
rlabel polysilicon 1213 -3467 1213 -3467 0 1
rlabel polysilicon 1213 -3473 1213 -3473 0 3
rlabel polysilicon 1220 -3467 1220 -3467 0 1
rlabel polysilicon 1223 -3467 1223 -3467 0 2
rlabel polysilicon 1220 -3473 1220 -3473 0 3
rlabel polysilicon 1227 -3467 1227 -3467 0 1
rlabel polysilicon 1227 -3473 1227 -3473 0 3
rlabel polysilicon 1353 -3467 1353 -3467 0 1
rlabel polysilicon 1353 -3473 1353 -3473 0 3
rlabel polysilicon 1360 -3467 1360 -3467 0 1
rlabel polysilicon 1360 -3473 1360 -3473 0 3
rlabel polysilicon 1409 -3467 1409 -3467 0 1
rlabel polysilicon 1409 -3473 1409 -3473 0 3
rlabel polysilicon 1412 -3473 1412 -3473 0 4
rlabel polysilicon 1416 -3467 1416 -3467 0 1
rlabel polysilicon 1416 -3473 1416 -3473 0 3
rlabel polysilicon 261 -3490 261 -3490 0 1
rlabel polysilicon 261 -3496 261 -3496 0 3
rlabel polysilicon 268 -3490 268 -3490 0 1
rlabel polysilicon 268 -3496 268 -3496 0 3
rlabel polysilicon 310 -3490 310 -3490 0 1
rlabel polysilicon 310 -3496 310 -3496 0 3
rlabel polysilicon 331 -3490 331 -3490 0 1
rlabel polysilicon 331 -3496 331 -3496 0 3
rlabel polysilicon 338 -3490 338 -3490 0 1
rlabel polysilicon 338 -3496 338 -3496 0 3
rlabel polysilicon 345 -3496 345 -3496 0 3
rlabel polysilicon 352 -3490 352 -3490 0 1
rlabel polysilicon 352 -3496 352 -3496 0 3
rlabel polysilicon 408 -3490 408 -3490 0 1
rlabel polysilicon 408 -3496 408 -3496 0 3
rlabel polysilicon 418 -3490 418 -3490 0 2
rlabel polysilicon 418 -3496 418 -3496 0 4
rlabel polysilicon 429 -3490 429 -3490 0 1
rlabel polysilicon 429 -3496 429 -3496 0 3
rlabel polysilicon 436 -3490 436 -3490 0 1
rlabel polysilicon 436 -3496 436 -3496 0 3
rlabel polysilicon 478 -3490 478 -3490 0 1
rlabel polysilicon 478 -3496 478 -3496 0 3
rlabel polysilicon 541 -3490 541 -3490 0 1
rlabel polysilicon 541 -3496 541 -3496 0 3
rlabel polysilicon 548 -3490 548 -3490 0 1
rlabel polysilicon 548 -3496 548 -3496 0 3
rlabel polysilicon 555 -3496 555 -3496 0 3
rlabel polysilicon 569 -3490 569 -3490 0 1
rlabel polysilicon 569 -3496 569 -3496 0 3
rlabel polysilicon 576 -3490 576 -3490 0 1
rlabel polysilicon 576 -3496 576 -3496 0 3
rlabel polysilicon 583 -3490 583 -3490 0 1
rlabel polysilicon 583 -3496 583 -3496 0 3
rlabel polysilicon 590 -3490 590 -3490 0 1
rlabel polysilicon 590 -3496 590 -3496 0 3
rlabel polysilicon 597 -3490 597 -3490 0 1
rlabel polysilicon 597 -3496 597 -3496 0 3
rlabel polysilicon 646 -3490 646 -3490 0 1
rlabel polysilicon 646 -3496 646 -3496 0 3
rlabel polysilicon 653 -3490 653 -3490 0 1
rlabel polysilicon 653 -3496 653 -3496 0 3
rlabel polysilicon 660 -3490 660 -3490 0 1
rlabel polysilicon 660 -3496 660 -3496 0 3
rlabel polysilicon 681 -3490 681 -3490 0 1
rlabel polysilicon 681 -3496 681 -3496 0 3
rlabel polysilicon 688 -3490 688 -3490 0 1
rlabel polysilicon 688 -3496 688 -3496 0 3
rlabel polysilicon 716 -3490 716 -3490 0 1
rlabel polysilicon 716 -3496 716 -3496 0 3
rlabel polysilicon 726 -3490 726 -3490 0 2
rlabel polysilicon 723 -3496 723 -3496 0 3
rlabel polysilicon 828 -3490 828 -3490 0 1
rlabel polysilicon 828 -3496 828 -3496 0 3
rlabel polysilicon 835 -3490 835 -3490 0 1
rlabel polysilicon 835 -3496 835 -3496 0 3
rlabel polysilicon 842 -3496 842 -3496 0 3
rlabel polysilicon 849 -3490 849 -3490 0 1
rlabel polysilicon 849 -3496 849 -3496 0 3
rlabel polysilicon 877 -3490 877 -3490 0 1
rlabel polysilicon 877 -3496 877 -3496 0 3
rlabel polysilicon 884 -3490 884 -3490 0 1
rlabel polysilicon 887 -3490 887 -3490 0 2
rlabel polysilicon 898 -3490 898 -3490 0 1
rlabel polysilicon 898 -3496 898 -3496 0 3
rlabel polysilicon 905 -3490 905 -3490 0 1
rlabel polysilicon 905 -3496 905 -3496 0 3
rlabel polysilicon 912 -3490 912 -3490 0 1
rlabel polysilicon 912 -3496 912 -3496 0 3
rlabel polysilicon 919 -3490 919 -3490 0 1
rlabel polysilicon 919 -3496 919 -3496 0 3
rlabel polysilicon 926 -3490 926 -3490 0 1
rlabel polysilicon 926 -3496 926 -3496 0 3
rlabel polysilicon 940 -3490 940 -3490 0 1
rlabel polysilicon 940 -3496 940 -3496 0 3
rlabel polysilicon 950 -3490 950 -3490 0 2
rlabel polysilicon 950 -3496 950 -3496 0 4
rlabel polysilicon 992 -3490 992 -3490 0 2
rlabel polysilicon 989 -3496 989 -3496 0 3
rlabel polysilicon 996 -3490 996 -3490 0 1
rlabel polysilicon 996 -3496 996 -3496 0 3
rlabel polysilicon 1094 -3490 1094 -3490 0 1
rlabel polysilicon 1094 -3496 1094 -3496 0 3
rlabel polysilicon 1115 -3490 1115 -3490 0 1
rlabel polysilicon 1115 -3496 1115 -3496 0 3
rlabel polysilicon 1118 -3496 1118 -3496 0 4
rlabel polysilicon 1122 -3490 1122 -3490 0 1
rlabel polysilicon 1122 -3496 1122 -3496 0 3
rlabel polysilicon 1220 -3490 1220 -3490 0 1
rlabel polysilicon 1353 -3490 1353 -3490 0 1
rlabel polysilicon 1353 -3496 1353 -3496 0 3
rlabel polysilicon 1360 -3490 1360 -3490 0 1
rlabel polysilicon 1360 -3496 1360 -3496 0 3
rlabel polysilicon 1409 -3490 1409 -3490 0 1
rlabel polysilicon 1412 -3490 1412 -3490 0 2
rlabel polysilicon 1412 -3496 1412 -3496 0 4
rlabel polysilicon 1416 -3490 1416 -3490 0 1
rlabel polysilicon 1416 -3496 1416 -3496 0 3
rlabel polysilicon 271 -3505 271 -3505 0 2
rlabel polysilicon 271 -3511 271 -3511 0 4
rlabel polysilicon 275 -3505 275 -3505 0 1
rlabel polysilicon 275 -3511 275 -3511 0 3
rlabel polysilicon 324 -3505 324 -3505 0 1
rlabel polysilicon 327 -3511 327 -3511 0 4
rlabel polysilicon 331 -3505 331 -3505 0 1
rlabel polysilicon 331 -3511 331 -3511 0 3
rlabel polysilicon 355 -3505 355 -3505 0 2
rlabel polysilicon 355 -3511 355 -3511 0 4
rlabel polysilicon 359 -3505 359 -3505 0 1
rlabel polysilicon 359 -3511 359 -3511 0 3
rlabel polysilicon 541 -3505 541 -3505 0 1
rlabel polysilicon 541 -3511 541 -3511 0 3
rlabel polysilicon 551 -3505 551 -3505 0 2
rlabel polysilicon 555 -3511 555 -3511 0 3
rlabel polysilicon 565 -3505 565 -3505 0 2
rlabel polysilicon 565 -3511 565 -3511 0 4
rlabel polysilicon 569 -3505 569 -3505 0 1
rlabel polysilicon 569 -3511 569 -3511 0 3
rlabel polysilicon 576 -3505 576 -3505 0 1
rlabel polysilicon 579 -3511 579 -3511 0 4
rlabel polysilicon 583 -3505 583 -3505 0 1
rlabel polysilicon 583 -3511 583 -3511 0 3
rlabel polysilicon 660 -3511 660 -3511 0 3
rlabel polysilicon 667 -3505 667 -3505 0 1
rlabel polysilicon 667 -3511 667 -3511 0 3
rlabel polysilicon 688 -3505 688 -3505 0 1
rlabel polysilicon 691 -3505 691 -3505 0 2
rlabel polysilicon 859 -3505 859 -3505 0 2
rlabel polysilicon 856 -3511 856 -3511 0 3
rlabel polysilicon 870 -3505 870 -3505 0 1
rlabel polysilicon 870 -3511 870 -3511 0 3
rlabel polysilicon 877 -3505 877 -3505 0 1
rlabel polysilicon 877 -3511 877 -3511 0 3
rlabel polysilicon 912 -3505 912 -3505 0 1
rlabel polysilicon 915 -3511 915 -3511 0 4
rlabel polysilicon 919 -3505 919 -3505 0 1
rlabel polysilicon 922 -3505 922 -3505 0 2
rlabel polysilicon 1353 -3505 1353 -3505 0 1
rlabel polysilicon 1353 -3511 1353 -3511 0 3
rlabel polysilicon 1360 -3511 1360 -3511 0 3
rlabel polysilicon 1363 -3511 1363 -3511 0 4
rlabel polysilicon 1367 -3505 1367 -3505 0 1
rlabel polysilicon 1367 -3511 1367 -3511 0 3
rlabel metal2 282 1 282 1 0 net=10991
rlabel metal2 425 1 425 1 0 net=6739
rlabel metal2 464 1 464 1 0 net=5629
rlabel metal2 905 1 905 1 0 net=12253
rlabel metal2 317 -1 317 -1 0 net=11673
rlabel metal2 436 -1 436 -1 0 net=8305
rlabel metal2 947 -1 947 -1 0 net=12025
rlabel metal2 443 -3 443 -3 0 net=2547
rlabel metal2 226 -14 226 -14 0 net=5715
rlabel metal2 303 -14 303 -14 0 net=11675
rlabel metal2 338 -14 338 -14 0 net=7909
rlabel metal2 366 -14 366 -14 0 net=2681
rlabel metal2 450 -14 450 -14 0 net=6741
rlabel metal2 478 -14 478 -14 0 net=3673
rlabel metal2 506 -14 506 -14 0 net=11241
rlabel metal2 618 -14 618 -14 0 net=5919
rlabel metal2 891 -14 891 -14 0 net=12255
rlabel metal2 989 -14 989 -14 0 net=12027
rlabel metal2 345 -16 345 -16 0 net=10993
rlabel metal2 380 -16 380 -16 0 net=3317
rlabel metal2 436 -16 436 -16 0 net=2549
rlabel metal2 450 -16 450 -16 0 net=5631
rlabel metal2 513 -16 513 -16 0 net=8307
rlabel metal2 579 -16 579 -16 0 net=10117
rlabel metal2 597 -16 597 -16 0 net=12171
rlabel metal2 289 -18 289 -18 0 net=1959
rlabel metal2 348 -18 348 -18 0 net=4217
rlabel metal2 422 -18 422 -18 0 net=5755
rlabel metal2 527 -18 527 -18 0 net=8327
rlabel metal2 583 -18 583 -18 0 net=9699
rlabel metal2 352 -20 352 -20 0 net=1827
rlabel metal2 394 -20 394 -20 0 net=2519
rlabel metal2 460 -20 460 -20 0 net=11333
rlabel metal2 509 -20 509 -20 0 net=9393
rlabel metal2 537 -20 537 -20 0 net=8009
rlabel metal2 352 -22 352 -22 0 net=4929
rlabel metal2 219 -33 219 -33 0 net=5717
rlabel metal2 275 -33 275 -33 0 net=1961
rlabel metal2 303 -33 303 -33 0 net=11677
rlabel metal2 303 -33 303 -33 0 net=11677
rlabel metal2 324 -33 324 -33 0 net=2683
rlabel metal2 373 -33 373 -33 0 net=10995
rlabel metal2 373 -33 373 -33 0 net=10995
rlabel metal2 387 -33 387 -33 0 net=1829
rlabel metal2 415 -33 415 -33 0 net=2551
rlabel metal2 443 -33 443 -33 0 net=6743
rlabel metal2 464 -33 464 -33 0 net=11335
rlabel metal2 492 -33 492 -33 0 net=6351
rlabel metal2 576 -33 576 -33 0 net=12173
rlabel metal2 604 -33 604 -33 0 net=9701
rlabel metal2 604 -33 604 -33 0 net=9701
rlabel metal2 611 -33 611 -33 0 net=11243
rlabel metal2 674 -33 674 -33 0 net=8011
rlabel metal2 758 -33 758 -33 0 net=6213
rlabel metal2 884 -33 884 -33 0 net=12257
rlabel metal2 1003 -33 1003 -33 0 net=12029
rlabel metal2 282 -35 282 -35 0 net=3599
rlabel metal2 331 -35 331 -35 0 net=4111
rlabel metal2 352 -35 352 -35 0 net=4931
rlabel metal2 352 -35 352 -35 0 net=4931
rlabel metal2 359 -35 359 -35 0 net=3919
rlabel metal2 436 -35 436 -35 0 net=6827
rlabel metal2 499 -35 499 -35 0 net=3675
rlabel metal2 513 -35 513 -35 0 net=9394
rlabel metal2 541 -35 541 -35 0 net=8329
rlabel metal2 583 -35 583 -35 0 net=5013
rlabel metal2 625 -35 625 -35 0 net=5921
rlabel metal2 639 -35 639 -35 0 net=8291
rlabel metal2 338 -37 338 -37 0 net=7911
rlabel metal2 366 -37 366 -37 0 net=3319
rlabel metal2 387 -37 387 -37 0 net=2573
rlabel metal2 499 -37 499 -37 0 net=6793
rlabel metal2 520 -37 520 -37 0 net=4517
rlabel metal2 551 -37 551 -37 0 net=12625
rlabel metal2 338 -39 338 -39 0 net=5756
rlabel metal2 450 -39 450 -39 0 net=5633
rlabel metal2 523 -39 523 -39 0 net=7967
rlabel metal2 590 -39 590 -39 0 net=10119
rlabel metal2 625 -39 625 -39 0 net=5397
rlabel metal2 380 -41 380 -41 0 net=2521
rlabel metal2 408 -41 408 -41 0 net=4219
rlabel metal2 548 -41 548 -41 0 net=8309
rlabel metal2 635 -41 635 -41 0 net=9711
rlabel metal2 394 -43 394 -43 0 net=3295
rlabel metal2 408 -45 408 -45 0 net=1889
rlabel metal2 422 -45 422 -45 0 net=6171
rlabel metal2 191 -56 191 -56 0 net=10807
rlabel metal2 278 -56 278 -56 0 net=3600
rlabel metal2 289 -56 289 -56 0 net=5635
rlabel metal2 506 -56 506 -56 0 net=3676
rlabel metal2 523 -56 523 -56 0 net=10633
rlabel metal2 789 -56 789 -56 0 net=10827
rlabel metal2 884 -56 884 -56 0 net=12259
rlabel metal2 1010 -56 1010 -56 0 net=12031
rlabel metal2 205 -58 205 -58 0 net=4119
rlabel metal2 243 -58 243 -58 0 net=1643
rlabel metal2 275 -58 275 -58 0 net=1963
rlabel metal2 296 -58 296 -58 0 net=11678
rlabel metal2 317 -58 317 -58 0 net=7913
rlabel metal2 401 -58 401 -58 0 net=1831
rlabel metal2 401 -58 401 -58 0 net=1831
rlabel metal2 408 -58 408 -58 0 net=1891
rlabel metal2 408 -58 408 -58 0 net=1891
rlabel metal2 464 -58 464 -58 0 net=6795
rlabel metal2 513 -58 513 -58 0 net=4518
rlabel metal2 527 -58 527 -58 0 net=4423
rlabel metal2 597 -58 597 -58 0 net=10121
rlabel metal2 709 -58 709 -58 0 net=6215
rlabel metal2 793 -58 793 -58 0 net=12065
rlabel metal2 828 -58 828 -58 0 net=12387
rlabel metal2 219 -60 219 -60 0 net=5719
rlabel metal2 275 -60 275 -60 0 net=3837
rlabel metal2 341 -60 341 -60 0 net=7912
rlabel metal2 390 -60 390 -60 0 net=9545
rlabel metal2 562 -60 562 -60 0 net=546
rlabel metal2 233 -62 233 -62 0 net=1805
rlabel metal2 345 -62 345 -62 0 net=2523
rlabel metal2 471 -62 471 -62 0 net=11337
rlabel metal2 569 -62 569 -62 0 net=5398
rlabel metal2 632 -62 632 -62 0 net=5923
rlabel metal2 653 -62 653 -62 0 net=11245
rlabel metal2 730 -62 730 -62 0 net=12627
rlabel metal2 299 -64 299 -64 0 net=147
rlabel metal2 373 -64 373 -64 0 net=10996
rlabel metal2 471 -64 471 -64 0 net=4055
rlabel metal2 569 -64 569 -64 0 net=5015
rlabel metal2 590 -64 590 -64 0 net=8311
rlabel metal2 604 -64 604 -64 0 net=9703
rlabel metal2 639 -64 639 -64 0 net=9713
rlabel metal2 723 -64 723 -64 0 net=8013
rlabel metal2 219 -66 219 -66 0 net=2271
rlabel metal2 303 -66 303 -66 0 net=2685
rlabel metal2 338 -66 338 -66 0 net=3963
rlabel metal2 576 -66 576 -66 0 net=12175
rlabel metal2 604 -66 604 -66 0 net=8325
rlabel metal2 681 -66 681 -66 0 net=9625
rlabel metal2 324 -68 324 -68 0 net=2323
rlabel metal2 555 -68 555 -68 0 net=8331
rlabel metal2 611 -68 611 -68 0 net=10929
rlabel metal2 621 -68 621 -68 0 net=11823
rlabel metal2 373 -70 373 -70 0 net=6745
rlabel metal2 485 -70 485 -70 0 net=2575
rlabel metal2 572 -70 572 -70 0 net=10159
rlabel metal2 614 -70 614 -70 0 net=6723
rlabel metal2 674 -70 674 -70 0 net=8293
rlabel metal2 436 -72 436 -72 0 net=6829
rlabel metal2 457 -72 457 -72 0 net=5083
rlabel metal2 520 -72 520 -72 0 net=10409
rlabel metal2 383 -74 383 -74 0 net=4867
rlabel metal2 541 -74 541 -74 0 net=7969
rlabel metal2 422 -76 422 -76 0 net=6173
rlabel metal2 422 -78 422 -78 0 net=6353
rlabel metal2 429 -80 429 -80 0 net=6405
rlabel metal2 415 -82 415 -82 0 net=2553
rlabel metal2 415 -84 415 -84 0 net=4221
rlabel metal2 331 -86 331 -86 0 net=4113
rlabel metal2 331 -88 331 -88 0 net=3921
rlabel metal2 352 -90 352 -90 0 net=4933
rlabel metal2 352 -92 352 -92 0 net=3321
rlabel metal2 366 -94 366 -94 0 net=3297
rlabel metal2 394 -96 394 -96 0 net=5619
rlabel metal2 114 -107 114 -107 0 net=10809
rlabel metal2 198 -107 198 -107 0 net=10507
rlabel metal2 299 -107 299 -107 0 net=35
rlabel metal2 471 -107 471 -107 0 net=4056
rlabel metal2 565 -107 565 -107 0 net=9801
rlabel metal2 723 -107 723 -107 0 net=9626
rlabel metal2 793 -107 793 -107 0 net=12067
rlabel metal2 891 -107 891 -107 0 net=12261
rlabel metal2 1010 -107 1010 -107 0 net=10379
rlabel metal2 121 -109 121 -109 0 net=9495
rlabel metal2 387 -109 387 -109 0 net=4114
rlabel metal2 509 -109 509 -109 0 net=8519
rlabel metal2 569 -109 569 -109 0 net=5016
rlabel metal2 569 -109 569 -109 0 net=5016
rlabel metal2 572 -109 572 -109 0 net=9955
rlabel metal2 782 -109 782 -109 0 net=11537
rlabel metal2 135 -111 135 -111 0 net=2157
rlabel metal2 334 -111 334 -111 0 net=10061
rlabel metal2 737 -111 737 -111 0 net=10635
rlabel metal2 898 -111 898 -111 0 net=12389
rlabel metal2 1017 -111 1017 -111 0 net=12033
rlabel metal2 142 -113 142 -113 0 net=4485
rlabel metal2 537 -113 537 -113 0 net=11891
rlabel metal2 863 -113 863 -113 0 net=10829
rlabel metal2 149 -115 149 -115 0 net=6747
rlabel metal2 380 -115 380 -115 0 net=2973
rlabel metal2 558 -115 558 -115 0 net=8326
rlabel metal2 611 -115 611 -115 0 net=10161
rlabel metal2 800 -115 800 -115 0 net=8169
rlabel metal2 156 -117 156 -117 0 net=3839
rlabel metal2 369 -117 369 -117 0 net=6119
rlabel metal2 583 -117 583 -117 0 net=12176
rlabel metal2 593 -117 593 -117 0 net=7093
rlabel metal2 807 -117 807 -117 0 net=12629
rlabel metal2 163 -119 163 -119 0 net=4121
rlabel metal2 212 -119 212 -119 0 net=3795
rlabel metal2 516 -119 516 -119 0 net=11097
rlabel metal2 863 -119 863 -119 0 net=8465
rlabel metal2 170 -121 170 -121 0 net=5637
rlabel metal2 310 -121 310 -121 0 net=1893
rlabel metal2 443 -121 443 -121 0 net=6831
rlabel metal2 614 -121 614 -121 0 net=9401
rlabel metal2 177 -123 177 -123 0 net=1587
rlabel metal2 240 -123 240 -123 0 net=2687
rlabel metal2 408 -123 408 -123 0 net=3591
rlabel metal2 618 -123 618 -123 0 net=10931
rlabel metal2 184 -125 184 -125 0 net=2273
rlabel metal2 226 -125 226 -125 0 net=275
rlabel metal2 586 -125 586 -125 0 net=9743
rlabel metal2 625 -125 625 -125 0 net=6971
rlabel metal2 191 -127 191 -127 0 net=5621
rlabel metal2 415 -127 415 -127 0 net=4223
rlabel metal2 450 -127 450 -127 0 net=11338
rlabel metal2 513 -127 513 -127 0 net=8039
rlabel metal2 576 -127 576 -127 0 net=8333
rlabel metal2 628 -127 628 -127 0 net=10045
rlabel metal2 205 -129 205 -129 0 net=1807
rlabel metal2 247 -129 247 -129 0 net=5721
rlabel metal2 394 -129 394 -129 0 net=2577
rlabel metal2 639 -129 639 -129 0 net=10411
rlabel metal2 219 -131 219 -131 0 net=2325
rlabel metal2 415 -131 415 -131 0 net=7509
rlabel metal2 639 -131 639 -131 0 net=5925
rlabel metal2 660 -131 660 -131 0 net=10123
rlabel metal2 233 -133 233 -133 0 net=3511
rlabel metal2 667 -133 667 -133 0 net=6725
rlabel metal2 247 -135 247 -135 0 net=1525
rlabel metal2 261 -135 261 -135 0 net=1645
rlabel metal2 261 -135 261 -135 0 net=1645
rlabel metal2 268 -135 268 -135 0 net=6355
rlabel metal2 464 -135 464 -135 0 net=6796
rlabel metal2 597 -135 597 -135 0 net=8313
rlabel metal2 681 -135 681 -135 0 net=8295
rlabel metal2 681 -135 681 -135 0 net=8295
rlabel metal2 688 -135 688 -135 0 net=11825
rlabel metal2 271 -137 271 -137 0 net=1055
rlabel metal2 282 -137 282 -137 0 net=1965
rlabel metal2 282 -137 282 -137 0 net=1965
rlabel metal2 289 -137 289 -137 0 net=1689
rlabel metal2 555 -137 555 -137 0 net=7971
rlabel metal2 632 -137 632 -137 0 net=9705
rlabel metal2 702 -137 702 -137 0 net=11247
rlabel metal2 275 -139 275 -139 0 net=3965
rlabel metal2 390 -139 390 -139 0 net=4551
rlabel metal2 464 -139 464 -139 0 net=4425
rlabel metal2 555 -139 555 -139 0 net=11219
rlabel metal2 702 -139 702 -139 0 net=8015
rlabel metal2 303 -141 303 -141 0 net=6381
rlabel metal2 527 -141 527 -141 0 net=10567
rlabel metal2 324 -143 324 -143 0 net=3323
rlabel metal2 478 -143 478 -143 0 net=9547
rlabel metal2 730 -143 730 -143 0 net=11207
rlabel metal2 338 -145 338 -145 0 net=3299
rlabel metal2 478 -145 478 -145 0 net=5085
rlabel metal2 492 -145 492 -145 0 net=6407
rlabel metal2 632 -145 632 -145 0 net=6217
rlabel metal2 128 -147 128 -147 0 net=4215
rlabel metal2 457 -147 457 -147 0 net=4869
rlabel metal2 492 -147 492 -147 0 net=4895
rlabel metal2 653 -147 653 -147 0 net=9715
rlabel metal2 345 -149 345 -149 0 net=2525
rlabel metal2 436 -149 436 -149 0 net=6175
rlabel metal2 499 -149 499 -149 0 net=9123
rlabel metal2 583 -149 583 -149 0 net=7269
rlabel metal2 656 -149 656 -149 0 net=8079
rlabel metal2 345 -151 345 -151 0 net=1833
rlabel metal2 359 -153 359 -153 0 net=4935
rlabel metal2 359 -155 359 -155 0 net=2555
rlabel metal2 317 -157 317 -157 0 net=7915
rlabel metal2 254 -159 254 -159 0 net=2103
rlabel metal2 401 -159 401 -159 0 net=10533
rlabel metal2 254 -161 254 -161 0 net=3923
rlabel metal2 331 -163 331 -163 0 net=7019
rlabel metal2 72 -174 72 -174 0 net=6009
rlabel metal2 597 -174 597 -174 0 net=7973
rlabel metal2 709 -174 709 -174 0 net=8081
rlabel metal2 898 -174 898 -174 0 net=10831
rlabel metal2 940 -174 940 -174 0 net=12391
rlabel metal2 1024 -174 1024 -174 0 net=12035
rlabel metal2 1136 -174 1136 -174 0 net=10381
rlabel metal2 86 -176 86 -176 0 net=11905
rlabel metal2 751 -176 751 -176 0 net=6727
rlabel metal2 1171 -176 1171 -176 0 net=11539
rlabel metal2 93 -178 93 -178 0 net=6357
rlabel metal2 275 -178 275 -178 0 net=3966
rlabel metal2 310 -178 310 -178 0 net=1894
rlabel metal2 457 -178 457 -178 0 net=6177
rlabel metal2 457 -178 457 -178 0 net=6177
rlabel metal2 478 -178 478 -178 0 net=5086
rlabel metal2 548 -178 548 -178 0 net=6409
rlabel metal2 597 -178 597 -178 0 net=6219
rlabel metal2 772 -178 772 -178 0 net=10163
rlabel metal2 919 -178 919 -178 0 net=12263
rlabel metal2 100 -180 100 -180 0 net=10509
rlabel metal2 205 -180 205 -180 0 net=1808
rlabel metal2 446 -180 446 -180 0 net=11319
rlabel metal2 107 -182 107 -182 0 net=7511
rlabel metal2 513 -182 513 -182 0 net=9399
rlabel metal2 793 -182 793 -182 0 net=10933
rlabel metal2 114 -184 114 -184 0 net=10810
rlabel metal2 222 -184 222 -184 0 net=10903
rlabel metal2 121 -186 121 -186 0 net=9496
rlabel metal2 240 -186 240 -186 0 net=2688
rlabel metal2 401 -186 401 -186 0 net=3429
rlabel metal2 520 -186 520 -186 0 net=9675
rlabel metal2 800 -186 800 -186 0 net=11099
rlabel metal2 121 -188 121 -188 0 net=4487
rlabel metal2 149 -188 149 -188 0 net=6749
rlabel metal2 576 -188 576 -188 0 net=9125
rlabel metal2 716 -188 716 -188 0 net=10047
rlabel metal2 807 -188 807 -188 0 net=11249
rlabel metal2 142 -190 142 -190 0 net=7021
rlabel metal2 523 -190 523 -190 0 net=46
rlabel metal2 674 -190 674 -190 0 net=11221
rlabel metal2 149 -192 149 -192 0 net=2275
rlabel metal2 191 -192 191 -192 0 net=5623
rlabel metal2 534 -192 534 -192 0 net=6121
rlabel metal2 625 -192 625 -192 0 net=8335
rlabel metal2 681 -192 681 -192 0 net=8297
rlabel metal2 737 -192 737 -192 0 net=9403
rlabel metal2 814 -192 814 -192 0 net=11827
rlabel metal2 79 -194 79 -194 0 net=8637
rlabel metal2 681 -194 681 -194 0 net=9717
rlabel metal2 702 -194 702 -194 0 net=8017
rlabel metal2 744 -194 744 -194 0 net=9957
rlabel metal2 821 -194 821 -194 0 net=11893
rlabel metal2 163 -196 163 -196 0 net=4123
rlabel metal2 282 -196 282 -196 0 net=1967
rlabel metal2 282 -196 282 -196 0 net=1967
rlabel metal2 289 -196 289 -196 0 net=1691
rlabel metal2 310 -196 310 -196 0 net=1935
rlabel metal2 422 -196 422 -196 0 net=4553
rlabel metal2 555 -196 555 -196 0 net=5263
rlabel metal2 667 -196 667 -196 0 net=9707
rlabel metal2 828 -196 828 -196 0 net=10569
rlabel metal2 163 -198 163 -198 0 net=1589
rlabel metal2 184 -198 184 -198 0 net=2327
rlabel metal2 233 -198 233 -198 0 net=3513
rlabel metal2 432 -198 432 -198 0 net=11703
rlabel metal2 835 -198 835 -198 0 net=11209
rlabel metal2 114 -200 114 -200 0 net=7787
rlabel metal2 233 -200 233 -200 0 net=1387
rlabel metal2 436 -200 436 -200 0 net=4937
rlabel metal2 558 -200 558 -200 0 net=7295
rlabel metal2 688 -200 688 -200 0 net=4631
rlabel metal2 765 -200 765 -200 0 net=10125
rlabel metal2 856 -200 856 -200 0 net=12069
rlabel metal2 170 -202 170 -202 0 net=5639
rlabel metal2 243 -202 243 -202 0 net=4455
rlabel metal2 464 -202 464 -202 0 net=4427
rlabel metal2 562 -202 562 -202 0 net=8521
rlabel metal2 618 -202 618 -202 0 net=9745
rlabel metal2 870 -202 870 -202 0 net=12631
rlabel metal2 156 -204 156 -204 0 net=3841
rlabel metal2 177 -204 177 -204 0 net=5401
rlabel metal2 443 -204 443 -204 0 net=4225
rlabel metal2 471 -204 471 -204 0 net=6833
rlabel metal2 702 -204 702 -204 0 net=7095
rlabel metal2 786 -204 786 -204 0 net=10535
rlabel metal2 877 -204 877 -204 0 net=8171
rlabel metal2 128 -206 128 -206 0 net=4216
rlabel metal2 471 -206 471 -206 0 net=4897
rlabel metal2 607 -206 607 -206 0 net=9337
rlabel metal2 842 -206 842 -206 0 net=10637
rlabel metal2 128 -208 128 -208 0 net=7471
rlabel metal2 229 -208 229 -208 0 net=10283
rlabel metal2 191 -210 191 -210 0 net=2909
rlabel metal2 261 -210 261 -210 0 net=1647
rlabel metal2 289 -210 289 -210 0 net=2527
rlabel metal2 387 -210 387 -210 0 net=9865
rlabel metal2 247 -212 247 -212 0 net=1527
rlabel metal2 331 -212 331 -212 0 net=3300
rlabel metal2 352 -212 352 -212 0 net=4917
rlabel metal2 380 -212 380 -212 0 net=2975
rlabel metal2 394 -212 394 -212 0 net=2579
rlabel metal2 485 -212 485 -212 0 net=4871
rlabel metal2 618 -212 618 -212 0 net=8315
rlabel metal2 660 -212 660 -212 0 net=9549
rlabel metal2 212 -214 212 -214 0 net=3797
rlabel metal2 373 -214 373 -214 0 net=5723
rlabel metal2 394 -214 394 -214 0 net=3905
rlabel metal2 611 -214 611 -214 0 net=8877
rlabel metal2 723 -214 723 -214 0 net=10063
rlabel metal2 212 -216 212 -216 0 net=1985
rlabel metal2 611 -216 611 -216 0 net=11811
rlabel metal2 247 -218 247 -218 0 net=3325
rlabel metal2 359 -218 359 -218 0 net=2557
rlabel metal2 429 -218 429 -218 0 net=7917
rlabel metal2 723 -218 723 -218 0 net=8467
rlabel metal2 135 -220 135 -220 0 net=2158
rlabel metal2 492 -220 492 -220 0 net=8041
rlabel metal2 779 -220 779 -220 0 net=10413
rlabel metal2 135 -222 135 -222 0 net=3925
rlabel metal2 317 -222 317 -222 0 net=2105
rlabel metal2 345 -222 345 -222 0 net=1835
rlabel metal2 499 -222 499 -222 0 net=6013
rlabel metal2 695 -222 695 -222 0 net=9803
rlabel metal2 254 -224 254 -224 0 net=6382
rlabel metal2 317 -224 317 -224 0 net=3593
rlabel metal2 541 -224 541 -224 0 net=5927
rlabel metal2 695 -224 695 -224 0 net=7815
rlabel metal2 303 -226 303 -226 0 net=9721
rlabel metal2 583 -226 583 -226 0 net=7271
rlabel metal2 324 -228 324 -228 0 net=2737
rlabel metal2 583 -228 583 -228 0 net=6973
rlabel metal2 345 -230 345 -230 0 net=1553
rlabel metal2 450 -230 450 -230 0 net=133
rlabel metal2 849 -230 849 -230 0 net=12499
rlabel metal2 93 -241 93 -241 0 net=6358
rlabel metal2 488 -241 488 -241 0 net=9550
rlabel metal2 884 -241 884 -241 0 net=8083
rlabel metal2 1185 -241 1185 -241 0 net=10383
rlabel metal2 1307 -241 1307 -241 0 net=11571
rlabel metal2 93 -243 93 -243 0 net=7023
rlabel metal2 145 -243 145 -243 0 net=3430
rlabel metal2 446 -243 446 -243 0 net=8042
rlabel metal2 502 -243 502 -243 0 net=10164
rlabel metal2 919 -243 919 -243 0 net=11223
rlabel metal2 1325 -243 1325 -243 0 net=11541
rlabel metal2 100 -245 100 -245 0 net=10510
rlabel metal2 177 -245 177 -245 0 net=5402
rlabel metal2 485 -245 485 -245 0 net=4433
rlabel metal2 754 -245 754 -245 0 net=11585
rlabel metal2 100 -247 100 -247 0 net=4677
rlabel metal2 247 -247 247 -247 0 net=3327
rlabel metal2 453 -247 453 -247 0 net=10934
rlabel metal2 1038 -247 1038 -247 0 net=12037
rlabel metal2 107 -249 107 -249 0 net=7512
rlabel metal2 492 -249 492 -249 0 net=4873
rlabel metal2 537 -249 537 -249 0 net=12719
rlabel metal2 107 -251 107 -251 0 net=7595
rlabel metal2 159 -251 159 -251 0 net=679
rlabel metal2 268 -251 268 -251 0 net=1649
rlabel metal2 268 -251 268 -251 0 net=1649
rlabel metal2 303 -251 303 -251 0 net=9722
rlabel metal2 600 -251 600 -251 0 net=12203
rlabel metal2 954 -251 954 -251 0 net=11813
rlabel metal2 128 -253 128 -253 0 net=7473
rlabel metal2 247 -253 247 -253 0 net=7331
rlabel metal2 369 -253 369 -253 0 net=6178
rlabel metal2 506 -253 506 -253 0 net=5625
rlabel metal2 551 -253 551 -253 0 net=8316
rlabel metal2 628 -253 628 -253 0 net=10219
rlabel metal2 968 -253 968 -253 0 net=12071
rlabel metal2 79 -255 79 -255 0 net=8639
rlabel metal2 138 -255 138 -255 0 net=4632
rlabel metal2 737 -255 737 -255 0 net=8019
rlabel metal2 765 -255 765 -255 0 net=9747
rlabel metal2 79 -257 79 -257 0 net=2277
rlabel metal2 163 -257 163 -257 0 net=1591
rlabel metal2 191 -257 191 -257 0 net=2911
rlabel metal2 205 -257 205 -257 0 net=777
rlabel metal2 233 -257 233 -257 0 net=2529
rlabel metal2 303 -257 303 -257 0 net=6123
rlabel metal2 618 -257 618 -257 0 net=3755
rlabel metal2 632 -257 632 -257 0 net=7975
rlabel metal2 716 -257 716 -257 0 net=8299
rlabel metal2 786 -257 786 -257 0 net=9867
rlabel metal2 877 -257 877 -257 0 net=10639
rlabel metal2 975 -257 975 -257 0 net=12633
rlabel metal2 114 -259 114 -259 0 net=7789
rlabel metal2 163 -259 163 -259 0 net=2329
rlabel metal2 191 -259 191 -259 0 net=6379
rlabel metal2 226 -259 226 -259 0 net=6015
rlabel metal2 632 -259 632 -259 0 net=6729
rlabel metal2 114 -261 114 -261 0 net=4489
rlabel metal2 170 -261 170 -261 0 net=3842
rlabel metal2 541 -261 541 -261 0 net=5929
rlabel metal2 670 -261 670 -261 0 net=11704
rlabel metal2 821 -261 821 -261 0 net=10065
rlabel metal2 891 -261 891 -261 0 net=10905
rlabel metal2 121 -263 121 -263 0 net=4919
rlabel metal2 366 -263 366 -263 0 net=2559
rlabel metal2 376 -263 376 -263 0 net=4938
rlabel metal2 541 -263 541 -263 0 net=5265
rlabel metal2 674 -263 674 -263 0 net=8337
rlabel metal2 982 -263 982 -263 0 net=12265
rlabel metal2 289 -265 289 -265 0 net=3907
rlabel metal2 450 -265 450 -265 0 net=4177
rlabel metal2 646 -265 646 -265 0 net=7919
rlabel metal2 695 -265 695 -265 0 net=7817
rlabel metal2 779 -265 779 -265 0 net=9805
rlabel metal2 835 -265 835 -265 0 net=10127
rlabel metal2 905 -265 905 -265 0 net=11211
rlabel metal2 198 -267 198 -267 0 net=5641
rlabel metal2 625 -267 625 -267 0 net=9065
rlabel metal2 793 -267 793 -267 0 net=10049
rlabel metal2 905 -267 905 -267 0 net=8173
rlabel metal2 198 -269 198 -269 0 net=1529
rlabel metal2 331 -269 331 -269 0 net=2107
rlabel metal2 380 -269 380 -269 0 net=5725
rlabel metal2 646 -269 646 -269 0 net=10849
rlabel metal2 989 -269 989 -269 0 net=12393
rlabel metal2 208 -271 208 -271 0 net=3029
rlabel metal2 380 -271 380 -271 0 net=8913
rlabel metal2 86 -273 86 -273 0 net=11906
rlabel metal2 212 -273 212 -273 0 net=1987
rlabel metal2 383 -273 383 -273 0 net=8522
rlabel metal2 709 -273 709 -273 0 net=9127
rlabel metal2 898 -273 898 -273 0 net=11101
rlabel metal2 996 -273 996 -273 0 net=12501
rlabel metal2 86 -275 86 -275 0 net=2269
rlabel metal2 450 -275 450 -275 0 net=2279
rlabel metal2 604 -275 604 -275 0 net=11828
rlabel metal2 184 -277 184 -277 0 net=1743
rlabel metal2 387 -277 387 -277 0 net=2977
rlabel metal2 415 -277 415 -277 0 net=3515
rlabel metal2 457 -277 457 -277 0 net=4227
rlabel metal2 478 -277 478 -277 0 net=9023
rlabel metal2 926 -277 926 -277 0 net=11251
rlabel metal2 187 -279 187 -279 0 net=6685
rlabel metal2 499 -279 499 -279 0 net=6221
rlabel metal2 607 -279 607 -279 0 net=10233
rlabel metal2 933 -279 933 -279 0 net=10833
rlabel metal2 317 -281 317 -281 0 net=3595
rlabel metal2 513 -281 513 -281 0 net=4555
rlabel metal2 534 -281 534 -281 0 net=4428
rlabel metal2 611 -281 611 -281 0 net=8501
rlabel metal2 723 -281 723 -281 0 net=8469
rlabel metal2 842 -281 842 -281 0 net=10285
rlabel metal2 940 -281 940 -281 0 net=11321
rlabel metal2 65 -283 65 -283 0 net=9663
rlabel metal2 590 -283 590 -283 0 net=6411
rlabel metal2 660 -283 660 -283 0 net=8879
rlabel metal2 744 -283 744 -283 0 net=9709
rlabel metal2 947 -283 947 -283 0 net=10571
rlabel metal2 317 -285 317 -285 0 net=2739
rlabel metal2 387 -285 387 -285 0 net=812
rlabel metal2 863 -285 863 -285 0 net=10415
rlabel metal2 961 -285 961 -285 0 net=11895
rlabel metal2 324 -287 324 -287 0 net=1555
rlabel metal2 390 -287 390 -287 0 net=6834
rlabel metal2 744 -287 744 -287 0 net=9847
rlabel metal2 870 -287 870 -287 0 net=10537
rlabel metal2 72 -289 72 -289 0 net=6011
rlabel metal2 394 -289 394 -289 0 net=4899
rlabel metal2 590 -289 590 -289 0 net=9993
rlabel metal2 72 -291 72 -291 0 net=1452
rlabel metal2 275 -291 275 -291 0 net=4125
rlabel metal2 653 -291 653 -291 0 net=7297
rlabel metal2 667 -291 667 -291 0 net=9400
rlabel metal2 800 -291 800 -291 0 net=9405
rlabel metal2 156 -293 156 -293 0 net=12435
rlabel metal2 275 -293 275 -293 0 net=1693
rlabel metal2 411 -293 411 -293 0 net=9267
rlabel metal2 170 -295 170 -295 0 net=9585
rlabel metal2 814 -295 814 -295 0 net=9959
rlabel metal2 254 -297 254 -297 0 net=3627
rlabel metal2 422 -297 422 -297 0 net=4457
rlabel metal2 639 -297 639 -297 0 net=7273
rlabel metal2 730 -297 730 -297 0 net=9677
rlabel metal2 828 -297 828 -297 0 net=10685
rlabel metal2 282 -299 282 -299 0 net=1969
rlabel metal2 422 -299 422 -299 0 net=2581
rlabel metal2 481 -299 481 -299 0 net=10601
rlabel metal2 135 -301 135 -301 0 net=3927
rlabel metal2 583 -301 583 -301 0 net=6975
rlabel metal2 681 -301 681 -301 0 net=9719
rlabel metal2 758 -301 758 -301 0 net=9339
rlabel metal2 243 -303 243 -303 0 net=3655
rlabel metal2 446 -303 446 -303 0 net=8955
rlabel metal2 569 -305 569 -305 0 net=6751
rlabel metal2 681 -305 681 -305 0 net=7097
rlabel metal2 338 -307 338 -307 0 net=3799
rlabel metal2 695 -307 695 -307 0 net=8565
rlabel metal2 338 -309 338 -309 0 net=1837
rlabel metal2 310 -311 310 -311 0 net=1937
rlabel metal2 310 -313 310 -313 0 net=9633
rlabel metal2 65 -324 65 -324 0 net=9664
rlabel metal2 446 -324 446 -324 0 net=5642
rlabel metal2 590 -324 590 -324 0 net=9748
rlabel metal2 1101 -324 1101 -324 0 net=12721
rlabel metal2 1381 -324 1381 -324 0 net=11543
rlabel metal2 1458 -324 1458 -324 0 net=11573
rlabel metal2 72 -326 72 -326 0 net=1286
rlabel metal2 369 -326 369 -326 0 net=3800
rlabel metal2 597 -326 597 -326 0 net=9710
rlabel metal2 912 -326 912 -326 0 net=12205
rlabel metal2 1171 -326 1171 -326 0 net=12461
rlabel metal2 72 -328 72 -328 0 net=4921
rlabel metal2 135 -328 135 -328 0 net=3909
rlabel metal2 345 -328 345 -328 0 net=6012
rlabel metal2 548 -328 548 -328 0 net=11224
rlabel metal2 1059 -328 1059 -328 0 net=12395
rlabel metal2 1199 -328 1199 -328 0 net=12725
rlabel metal2 79 -330 79 -330 0 net=2278
rlabel metal2 205 -330 205 -330 0 net=11814
rlabel metal2 1122 -330 1122 -330 0 net=8915
rlabel metal2 58 -332 58 -332 0 net=4855
rlabel metal2 250 -332 250 -332 0 net=7087
rlabel metal2 541 -332 541 -332 0 net=5267
rlabel metal2 551 -332 551 -332 0 net=8338
rlabel metal2 989 -332 989 -332 0 net=11103
rlabel metal2 1206 -332 1206 -332 0 net=10385
rlabel metal2 1206 -332 1206 -332 0 net=10385
rlabel metal2 79 -334 79 -334 0 net=7791
rlabel metal2 166 -334 166 -334 0 net=7383
rlabel metal2 597 -334 597 -334 0 net=7513
rlabel metal2 807 -334 807 -334 0 net=9635
rlabel metal2 926 -334 926 -334 0 net=10235
rlabel metal2 1003 -334 1003 -334 0 net=11213
rlabel metal2 86 -336 86 -336 0 net=2270
rlabel metal2 478 -336 478 -336 0 net=4691
rlabel metal2 565 -336 565 -336 0 net=11463
rlabel metal2 86 -338 86 -338 0 net=5241
rlabel metal2 604 -338 604 -338 0 net=3756
rlabel metal2 625 -338 625 -338 0 net=10906
rlabel metal2 1066 -338 1066 -338 0 net=12039
rlabel metal2 93 -340 93 -340 0 net=7024
rlabel metal2 618 -340 618 -340 0 net=7299
rlabel metal2 667 -340 667 -340 0 net=7977
rlabel metal2 702 -340 702 -340 0 net=8567
rlabel metal2 821 -340 821 -340 0 net=9807
rlabel metal2 975 -340 975 -340 0 net=10835
rlabel metal2 1073 -340 1073 -340 0 net=12635
rlabel metal2 93 -342 93 -342 0 net=7681
rlabel metal2 464 -342 464 -342 0 net=6687
rlabel metal2 625 -342 625 -342 0 net=8853
rlabel metal2 835 -342 835 -342 0 net=9849
rlabel metal2 961 -342 961 -342 0 net=10687
rlabel metal2 1017 -342 1017 -342 0 net=11323
rlabel metal2 100 -344 100 -344 0 net=4678
rlabel metal2 191 -344 191 -344 0 net=6380
rlabel metal2 464 -344 464 -344 0 net=5727
rlabel metal2 583 -344 583 -344 0 net=6753
rlabel metal2 702 -344 702 -344 0 net=9129
rlabel metal2 856 -344 856 -344 0 net=9869
rlabel metal2 947 -344 947 -344 0 net=10539
rlabel metal2 1024 -344 1024 -344 0 net=11897
rlabel metal2 100 -346 100 -346 0 net=12437
rlabel metal2 170 -346 170 -346 0 net=9268
rlabel metal2 856 -346 856 -346 0 net=8175
rlabel metal2 947 -346 947 -346 0 net=11253
rlabel metal2 1031 -346 1031 -346 0 net=12073
rlabel metal2 121 -348 121 -348 0 net=8641
rlabel metal2 149 -348 149 -348 0 net=55
rlabel metal2 345 -348 345 -348 0 net=2281
rlabel metal2 495 -348 495 -348 0 net=4458
rlabel metal2 555 -348 555 -348 0 net=7275
rlabel metal2 758 -348 758 -348 0 net=8957
rlabel metal2 870 -348 870 -348 0 net=9995
rlabel metal2 1080 -348 1080 -348 0 net=11587
rlabel metal2 128 -350 128 -350 0 net=6125
rlabel metal2 310 -350 310 -350 0 net=1939
rlabel metal2 373 -350 373 -350 0 net=4435
rlabel metal2 506 -350 506 -350 0 net=5627
rlabel metal2 628 -350 628 -350 0 net=9720
rlabel metal2 765 -350 765 -350 0 net=9025
rlabel metal2 884 -350 884 -350 0 net=10067
rlabel metal2 982 -350 982 -350 0 net=10851
rlabel metal2 1080 -350 1080 -350 0 net=8085
rlabel metal2 173 -352 173 -352 0 net=1483
rlabel metal2 583 -352 583 -352 0 net=8379
rlabel metal2 772 -352 772 -352 0 net=10603
rlabel metal2 1038 -352 1038 -352 0 net=12267
rlabel metal2 1087 -352 1087 -352 0 net=12503
rlabel metal2 107 -354 107 -354 0 net=7597
rlabel metal2 107 -356 107 -356 0 net=4491
rlabel metal2 173 -356 173 -356 0 net=5445
rlabel metal2 513 -356 513 -356 0 net=4179
rlabel metal2 632 -356 632 -356 0 net=6730
rlabel metal2 709 -356 709 -356 0 net=8503
rlabel metal2 786 -356 786 -356 0 net=11951
rlabel metal2 114 -358 114 -358 0 net=4127
rlabel metal2 481 -358 481 -358 0 net=7669
rlabel metal2 730 -358 730 -358 0 net=9587
rlabel metal2 814 -358 814 -358 0 net=9679
rlabel metal2 919 -358 919 -358 0 net=10221
rlabel metal2 996 -358 996 -358 0 net=10573
rlabel metal2 184 -360 184 -360 0 net=11453
rlabel metal2 138 -362 138 -362 0 net=793
rlabel metal2 194 -362 194 -362 0 net=5747
rlabel metal2 520 -362 520 -362 0 net=4557
rlabel metal2 572 -362 572 -362 0 net=9001
rlabel metal2 828 -362 828 -362 0 net=9341
rlabel metal2 891 -362 891 -362 0 net=10129
rlabel metal2 247 -364 247 -364 0 net=7333
rlabel metal2 793 -364 793 -364 0 net=8471
rlabel metal2 842 -364 842 -364 0 net=9407
rlabel metal2 940 -364 940 -364 0 net=10417
rlabel metal2 156 -366 156 -366 0 net=2123
rlabel metal2 282 -366 282 -366 0 net=3928
rlabel metal2 415 -366 415 -366 0 net=3597
rlabel metal2 646 -366 646 -366 0 net=6641
rlabel metal2 842 -366 842 -366 0 net=10287
rlabel metal2 954 -366 954 -366 0 net=10641
rlabel metal2 142 -368 142 -368 0 net=452
rlabel metal2 436 -368 436 -368 0 net=3657
rlabel metal2 586 -368 586 -368 0 net=9943
rlabel metal2 142 -370 142 -370 0 net=2331
rlabel metal2 233 -370 233 -370 0 net=2531
rlabel metal2 289 -370 289 -370 0 net=4861
rlabel metal2 723 -370 723 -370 0 net=8881
rlabel metal2 863 -370 863 -370 0 net=9961
rlabel metal2 233 -372 233 -372 0 net=3183
rlabel metal2 670 -372 670 -372 0 net=10307
rlabel metal2 303 -374 303 -374 0 net=1839
rlabel metal2 376 -374 376 -374 0 net=5353
rlabel metal2 737 -374 737 -374 0 net=8301
rlabel metal2 261 -376 261 -376 0 net=3031
rlabel metal2 387 -376 387 -376 0 net=8809
rlabel metal2 877 -376 877 -376 0 net=10051
rlabel metal2 212 -378 212 -378 0 net=1745
rlabel metal2 313 -378 313 -378 0 net=2725
rlabel metal2 408 -378 408 -378 0 net=2978
rlabel metal2 747 -378 747 -378 0 net=12059
rlabel metal2 212 -380 212 -380 0 net=2913
rlabel metal2 366 -380 366 -380 0 net=2561
rlabel metal2 436 -380 436 -380 0 net=6413
rlabel metal2 716 -380 716 -380 0 net=7819
rlabel metal2 779 -380 779 -380 0 net=9067
rlabel metal2 177 -382 177 -382 0 net=1593
rlabel metal2 443 -382 443 -382 0 net=8761
rlabel metal2 716 -382 716 -382 0 net=9281
rlabel metal2 177 -384 177 -384 0 net=3629
rlabel metal2 422 -384 422 -384 0 net=2583
rlabel metal2 562 -384 562 -384 0 net=5931
rlabel metal2 751 -384 751 -384 0 net=8021
rlabel metal2 240 -386 240 -386 0 net=7475
rlabel metal2 600 -386 600 -386 0 net=8695
rlabel metal2 240 -388 240 -388 0 net=4901
rlabel metal2 632 -388 632 -388 0 net=8273
rlabel metal2 254 -390 254 -390 0 net=1651
rlabel metal2 394 -390 394 -390 0 net=3329
rlabel metal2 198 -392 198 -392 0 net=1531
rlabel metal2 401 -392 401 -392 0 net=5317
rlabel metal2 198 -394 198 -394 0 net=4875
rlabel metal2 681 -394 681 -394 0 net=7099
rlabel metal2 275 -396 275 -396 0 net=1694
rlabel metal2 639 -396 639 -396 0 net=6977
rlabel metal2 275 -398 275 -398 0 net=1557
rlabel metal2 639 -398 639 -398 0 net=7921
rlabel metal2 324 -400 324 -400 0 net=1989
rlabel metal2 499 -400 499 -400 0 net=6223
rlabel metal2 226 -402 226 -402 0 net=6017
rlabel metal2 226 -404 226 -404 0 net=2741
rlabel metal2 331 -404 331 -404 0 net=2109
rlabel metal2 296 -406 296 -406 0 net=1971
rlabel metal2 352 -406 352 -406 0 net=4229
rlabel metal2 208 -408 208 -408 0 net=3777
rlabel metal2 296 -410 296 -410 0 net=3517
rlabel metal2 429 -412 429 -412 0 net=2693
rlabel metal2 51 -423 51 -423 0 net=4567
rlabel metal2 194 -423 194 -423 0 net=7334
rlabel metal2 838 -423 838 -423 0 net=12722
rlabel metal2 1388 -423 1388 -423 0 net=8917
rlabel metal2 1521 -423 1521 -423 0 net=11575
rlabel metal2 58 -425 58 -425 0 net=9941
rlabel metal2 149 -425 149 -425 0 net=2914
rlabel metal2 250 -425 250 -425 0 net=1972
rlabel metal2 359 -425 359 -425 0 net=5628
rlabel metal2 611 -425 611 -425 0 net=5932
rlabel metal2 656 -425 656 -425 0 net=9588
rlabel metal2 754 -425 754 -425 0 net=11104
rlabel metal2 1157 -425 1157 -425 0 net=12505
rlabel metal2 1409 -425 1409 -425 0 net=11545
rlabel metal2 65 -427 65 -427 0 net=8643
rlabel metal2 124 -427 124 -427 0 net=11324
rlabel metal2 1185 -427 1185 -427 0 net=12637
rlabel metal2 72 -429 72 -429 0 net=4922
rlabel metal2 450 -429 450 -429 0 net=3658
rlabel metal2 544 -429 544 -429 0 net=8882
rlabel metal2 856 -429 856 -429 0 net=8177
rlabel metal2 856 -429 856 -429 0 net=8177
rlabel metal2 891 -429 891 -429 0 net=9409
rlabel metal2 891 -429 891 -429 0 net=9409
rlabel metal2 919 -429 919 -429 0 net=8303
rlabel metal2 72 -431 72 -431 0 net=3929
rlabel metal2 572 -431 572 -431 0 net=9130
rlabel metal2 737 -431 737 -431 0 net=7821
rlabel metal2 870 -431 870 -431 0 net=9283
rlabel metal2 996 -431 996 -431 0 net=10309
rlabel metal2 996 -431 996 -431 0 net=10309
rlabel metal2 1073 -431 1073 -431 0 net=11455
rlabel metal2 1192 -431 1192 -431 0 net=11589
rlabel metal2 79 -433 79 -433 0 net=7793
rlabel metal2 79 -433 79 -433 0 net=7793
rlabel metal2 86 -433 86 -433 0 net=5242
rlabel metal2 177 -433 177 -433 0 net=3630
rlabel metal2 415 -433 415 -433 0 net=3598
rlabel metal2 541 -433 541 -433 0 net=6225
rlabel metal2 688 -433 688 -433 0 net=10288
rlabel metal2 1031 -433 1031 -433 0 net=10605
rlabel metal2 1080 -433 1080 -433 0 net=8087
rlabel metal2 86 -435 86 -435 0 net=4493
rlabel metal2 114 -435 114 -435 0 net=4129
rlabel metal2 163 -435 163 -435 0 net=7476
rlabel metal2 450 -435 450 -435 0 net=3439
rlabel metal2 558 -435 558 -435 0 net=7300
rlabel metal2 628 -435 628 -435 0 net=6781
rlabel metal2 821 -435 821 -435 0 net=9027
rlabel metal2 1108 -435 1108 -435 0 net=12041
rlabel metal2 1206 -435 1206 -435 0 net=10386
rlabel metal2 93 -437 93 -437 0 net=7682
rlabel metal2 691 -437 691 -437 0 net=11214
rlabel metal2 1136 -437 1136 -437 0 net=12075
rlabel metal2 1164 -437 1164 -437 0 net=12397
rlabel metal2 93 -439 93 -439 0 net=12439
rlabel metal2 114 -439 114 -439 0 net=6415
rlabel metal2 464 -439 464 -439 0 net=5729
rlabel metal2 548 -439 548 -439 0 net=5269
rlabel metal2 583 -439 583 -439 0 net=9808
rlabel metal2 1101 -439 1101 -439 0 net=11953
rlabel metal2 1164 -439 1164 -439 0 net=12727
rlabel metal2 100 -441 100 -441 0 net=4877
rlabel metal2 212 -441 212 -441 0 net=1559
rlabel metal2 296 -441 296 -441 0 net=3518
rlabel metal2 590 -441 590 -441 0 net=6642
rlabel metal2 663 -441 663 -441 0 net=7133
rlabel metal2 824 -441 824 -441 0 net=11229
rlabel metal2 1115 -441 1115 -441 0 net=12061
rlabel metal2 1171 -441 1171 -441 0 net=12463
rlabel metal2 121 -443 121 -443 0 net=7598
rlabel metal2 1094 -443 1094 -443 0 net=11899
rlabel metal2 1150 -443 1150 -443 0 net=12207
rlabel metal2 135 -445 135 -445 0 net=3911
rlabel metal2 495 -445 495 -445 0 net=11705
rlabel metal2 107 -447 107 -447 0 net=3277
rlabel metal2 138 -447 138 -447 0 net=302
rlabel metal2 852 -447 852 -447 0 net=10353
rlabel metal2 1045 -447 1045 -447 0 net=10837
rlabel metal2 142 -449 142 -449 0 net=2332
rlabel metal2 166 -449 166 -449 0 net=73
rlabel metal2 257 -449 257 -449 0 net=3032
rlabel metal2 359 -449 359 -449 0 net=4181
rlabel metal2 548 -449 548 -449 0 net=6688
rlabel metal2 632 -449 632 -449 0 net=12141
rlabel metal2 152 -451 152 -451 0 net=2003
rlabel metal2 366 -451 366 -451 0 net=5081
rlabel metal2 947 -451 947 -451 0 net=11255
rlabel metal2 166 -453 166 -453 0 net=608
rlabel metal2 170 -455 170 -455 0 net=7025
rlabel metal2 317 -455 317 -455 0 net=1991
rlabel metal2 366 -455 366 -455 0 net=5789
rlabel metal2 632 -455 632 -455 0 net=5735
rlabel metal2 177 -457 177 -457 0 net=6475
rlabel metal2 667 -457 667 -457 0 net=7979
rlabel metal2 905 -457 905 -457 0 net=9681
rlabel metal2 968 -457 968 -457 0 net=10223
rlabel metal2 1024 -457 1024 -457 0 net=10575
rlabel metal2 184 -459 184 -459 0 net=1595
rlabel metal2 247 -459 247 -459 0 net=5683
rlabel metal2 667 -459 667 -459 0 net=8275
rlabel metal2 835 -459 835 -459 0 net=9949
rlabel metal2 961 -459 961 -459 0 net=10069
rlabel metal2 989 -459 989 -459 0 net=10237
rlabel metal2 1038 -459 1038 -459 0 net=10643
rlabel metal2 191 -461 191 -461 0 net=869
rlabel metal2 219 -461 219 -461 0 net=4231
rlabel metal2 380 -461 380 -461 0 net=6183
rlabel metal2 695 -461 695 -461 0 net=7101
rlabel metal2 779 -461 779 -461 0 net=8023
rlabel metal2 898 -461 898 -461 0 net=9637
rlabel metal2 1017 -461 1017 -461 0 net=10541
rlabel metal2 142 -463 142 -463 0 net=9599
rlabel metal2 814 -463 814 -463 0 net=9003
rlabel metal2 954 -463 954 -463 0 net=10053
rlabel metal2 1010 -463 1010 -463 0 net=10419
rlabel metal2 191 -465 191 -465 0 net=6625
rlabel metal2 698 -465 698 -465 0 net=9996
rlabel metal2 261 -467 261 -467 0 net=1747
rlabel metal2 331 -467 331 -467 0 net=2111
rlabel metal2 383 -467 383 -467 0 net=3330
rlabel metal2 401 -467 401 -467 0 net=5319
rlabel metal2 464 -467 464 -467 0 net=6754
rlabel metal2 723 -467 723 -467 0 net=12453
rlabel metal2 261 -469 261 -469 0 net=1941
rlabel metal2 345 -469 345 -469 0 net=2283
rlabel metal2 394 -469 394 -469 0 net=2563
rlabel metal2 415 -469 415 -469 0 net=3105
rlabel metal2 726 -469 726 -469 0 net=12303
rlabel metal2 275 -471 275 -471 0 net=2533
rlabel metal2 296 -471 296 -471 0 net=2726
rlabel metal2 408 -471 408 -471 0 net=3033
rlabel metal2 877 -471 877 -471 0 net=8697
rlabel metal2 156 -473 156 -473 0 net=2125
rlabel metal2 303 -473 303 -473 0 net=1841
rlabel metal2 345 -473 345 -473 0 net=3493
rlabel metal2 471 -473 471 -473 0 net=5355
rlabel metal2 569 -473 569 -473 0 net=2667
rlabel metal2 765 -473 765 -473 0 net=8381
rlabel metal2 940 -473 940 -473 0 net=9963
rlabel metal2 1003 -473 1003 -473 0 net=10689
rlabel metal2 198 -475 198 -475 0 net=2353
rlabel metal2 418 -475 418 -475 0 net=7255
rlabel metal2 744 -475 744 -475 0 net=8569
rlabel metal2 800 -475 800 -475 0 net=8811
rlabel metal2 912 -475 912 -475 0 net=9851
rlabel metal2 303 -477 303 -477 0 net=5893
rlabel metal2 653 -477 653 -477 0 net=7671
rlabel metal2 772 -477 772 -477 0 net=8505
rlabel metal2 863 -477 863 -477 0 net=9069
rlabel metal2 310 -479 310 -479 0 net=2653
rlabel metal2 422 -479 422 -479 0 net=6978
rlabel metal2 807 -479 807 -479 0 net=8855
rlabel metal2 884 -479 884 -479 0 net=9343
rlabel metal2 429 -481 429 -481 0 net=2695
rlabel metal2 478 -481 478 -481 0 net=4693
rlabel metal2 653 -481 653 -481 0 net=6879
rlabel metal2 709 -481 709 -481 0 net=8763
rlabel metal2 828 -481 828 -481 0 net=8473
rlabel metal2 226 -483 226 -483 0 net=2743
rlabel metal2 478 -483 478 -483 0 net=6019
rlabel metal2 506 -483 506 -483 0 net=5447
rlabel metal2 597 -483 597 -483 0 net=7515
rlabel metal2 226 -485 226 -485 0 net=4903
rlabel metal2 373 -485 373 -485 0 net=4437
rlabel metal2 534 -485 534 -485 0 net=7089
rlabel metal2 205 -487 205 -487 0 net=4857
rlabel metal2 373 -487 373 -487 0 net=2585
rlabel metal2 485 -487 485 -487 0 net=5749
rlabel metal2 681 -487 681 -487 0 net=11464
rlabel metal2 128 -489 128 -489 0 net=6127
rlabel metal2 499 -489 499 -489 0 net=5565
rlabel metal2 1059 -489 1059 -489 0 net=12269
rlabel metal2 128 -491 128 -491 0 net=4565
rlabel metal2 443 -491 443 -491 0 net=3779
rlabel metal2 527 -491 527 -491 0 net=4559
rlabel metal2 555 -491 555 -491 0 net=7277
rlabel metal2 1059 -491 1059 -491 0 net=10853
rlabel metal2 205 -493 205 -493 0 net=3185
rlabel metal2 289 -493 289 -493 0 net=4863
rlabel metal2 555 -493 555 -493 0 net=6243
rlabel metal2 975 -493 975 -493 0 net=10131
rlabel metal2 268 -495 268 -495 0 net=1533
rlabel metal2 457 -495 457 -495 0 net=3395
rlabel metal2 933 -495 933 -495 0 net=9945
rlabel metal2 254 -497 254 -497 0 net=1653
rlabel metal2 576 -497 576 -497 0 net=7385
rlabel metal2 926 -497 926 -497 0 net=9871
rlabel metal2 156 -499 156 -499 0 net=2893
rlabel metal2 576 -499 576 -499 0 net=7923
rlabel metal2 849 -499 849 -499 0 net=8959
rlabel metal2 369 -501 369 -501 0 net=6433
rlabel metal2 44 -512 44 -512 0 net=4495
rlabel metal2 93 -512 93 -512 0 net=12441
rlabel metal2 1419 -512 1419 -512 0 net=7745
rlabel metal2 58 -514 58 -514 0 net=9942
rlabel metal2 649 -514 649 -514 0 net=11257
rlabel metal2 1430 -514 1430 -514 0 net=11547
rlabel metal2 1486 -514 1486 -514 0 net=8919
rlabel metal2 1542 -514 1542 -514 0 net=11577
rlabel metal2 58 -516 58 -516 0 net=5827
rlabel metal2 751 -516 751 -516 0 net=10606
rlabel metal2 1087 -516 1087 -516 0 net=10839
rlabel metal2 1227 -516 1227 -516 0 net=12507
rlabel metal2 65 -518 65 -518 0 net=8644
rlabel metal2 254 -518 254 -518 0 net=2285
rlabel metal2 387 -518 387 -518 0 net=11456
rlabel metal2 1178 -518 1178 -518 0 net=12271
rlabel metal2 65 -520 65 -520 0 net=2853
rlabel metal2 264 -520 264 -520 0 net=12127
rlabel metal2 72 -522 72 -522 0 net=3930
rlabel metal2 401 -522 401 -522 0 net=2669
rlabel metal2 590 -522 590 -522 0 net=7633
rlabel metal2 863 -522 863 -522 0 net=8857
rlabel metal2 72 -524 72 -524 0 net=6997
rlabel metal2 663 -524 663 -524 0 net=9004
rlabel metal2 905 -524 905 -524 0 net=9951
rlabel metal2 86 -526 86 -526 0 net=4131
rlabel metal2 156 -526 156 -526 0 net=2895
rlabel metal2 425 -526 425 -526 0 net=4475
rlabel metal2 593 -526 593 -526 0 net=10132
rlabel metal2 1115 -526 1115 -526 0 net=11901
rlabel metal2 93 -528 93 -528 0 net=4733
rlabel metal2 268 -528 268 -528 0 net=1654
rlabel metal2 296 -528 296 -528 0 net=849
rlabel metal2 450 -528 450 -528 0 net=3441
rlabel metal2 618 -528 618 -528 0 net=12521
rlabel metal2 121 -530 121 -530 0 net=2075
rlabel metal2 429 -530 429 -530 0 net=2745
rlabel metal2 520 -530 520 -530 0 net=5731
rlabel metal2 520 -530 520 -530 0 net=5731
rlabel metal2 527 -530 527 -530 0 net=4865
rlabel metal2 621 -530 621 -530 0 net=10527
rlabel metal2 128 -532 128 -532 0 net=4566
rlabel metal2 730 -532 730 -532 0 net=5082
rlabel metal2 821 -532 821 -532 0 net=7995
rlabel metal2 128 -534 128 -534 0 net=3187
rlabel metal2 296 -534 296 -534 0 net=3091
rlabel metal2 646 -534 646 -534 0 net=10420
rlabel metal2 1024 -534 1024 -534 0 net=10239
rlabel metal2 124 -536 124 -536 0 net=4793
rlabel metal2 299 -536 299 -536 0 net=4438
rlabel metal2 534 -536 534 -536 0 net=4561
rlabel metal2 555 -536 555 -536 0 net=8570
rlabel metal2 789 -536 789 -536 0 net=11777
rlabel metal2 135 -538 135 -538 0 net=4079
rlabel metal2 660 -538 660 -538 0 net=5981
rlabel metal2 1241 -538 1241 -538 0 net=11590
rlabel metal2 142 -540 142 -540 0 net=1596
rlabel metal2 191 -540 191 -540 0 net=4905
rlabel metal2 359 -540 359 -540 0 net=4183
rlabel metal2 555 -540 555 -540 0 net=7091
rlabel metal2 716 -540 716 -540 0 net=7257
rlabel metal2 856 -540 856 -540 0 net=8179
rlabel metal2 933 -540 933 -540 0 net=9873
rlabel metal2 142 -542 142 -542 0 net=3397
rlabel metal2 471 -542 471 -542 0 net=2697
rlabel metal2 625 -542 625 -542 0 net=6245
rlabel metal2 744 -542 744 -542 0 net=7673
rlabel metal2 873 -542 873 -542 0 net=9638
rlabel metal2 1010 -542 1010 -542 0 net=8699
rlabel metal2 1122 -542 1122 -542 0 net=12063
rlabel metal2 114 -544 114 -544 0 net=6417
rlabel metal2 653 -544 653 -544 0 net=11256
rlabel metal2 1129 -544 1129 -544 0 net=11955
rlabel metal2 100 -546 100 -546 0 net=4879
rlabel metal2 145 -546 145 -546 0 net=12471
rlabel metal2 100 -548 100 -548 0 net=3279
rlabel metal2 149 -548 149 -548 0 net=1535
rlabel metal2 359 -548 359 -548 0 net=2565
rlabel metal2 471 -548 471 -548 0 net=5449
rlabel metal2 632 -548 632 -548 0 net=5737
rlabel metal2 667 -548 667 -548 0 net=8277
rlabel metal2 919 -548 919 -548 0 net=9285
rlabel metal2 1017 -548 1017 -548 0 net=12728
rlabel metal2 1185 -548 1185 -548 0 net=12043
rlabel metal2 156 -550 156 -550 0 net=2357
rlabel metal2 674 -550 674 -550 0 net=6627
rlabel metal2 754 -550 754 -550 0 net=9009
rlabel metal2 110 -552 110 -552 0 net=10561
rlabel metal2 684 -552 684 -552 0 net=10843
rlabel metal2 163 -554 163 -554 0 net=11701
rlabel metal2 163 -556 163 -556 0 net=3813
rlabel metal2 268 -556 268 -556 0 net=3197
rlabel metal2 478 -556 478 -556 0 net=6021
rlabel metal2 684 -556 684 -556 0 net=9852
rlabel metal2 1024 -556 1024 -556 0 net=8089
rlabel metal2 166 -558 166 -558 0 net=5684
rlabel metal2 355 -558 355 -558 0 net=4801
rlabel metal2 611 -558 611 -558 0 net=4695
rlabel metal2 688 -558 688 -558 0 net=6881
rlabel metal2 800 -558 800 -558 0 net=8507
rlabel metal2 1143 -558 1143 -558 0 net=12077
rlabel metal2 177 -560 177 -560 0 net=6477
rlabel metal2 177 -560 177 -560 0 net=6477
rlabel metal2 184 -560 184 -560 0 net=5895
rlabel metal2 373 -560 373 -560 0 net=2587
rlabel metal2 443 -560 443 -560 0 net=3781
rlabel metal2 698 -560 698 -560 0 net=8304
rlabel metal2 194 -562 194 -562 0 net=11339
rlabel metal2 219 -564 219 -564 0 net=4233
rlabel metal2 394 -564 394 -564 0 net=5751
rlabel metal2 702 -564 702 -564 0 net=6783
rlabel metal2 744 -564 744 -564 0 net=11373
rlabel metal2 219 -566 219 -566 0 net=3495
rlabel metal2 366 -566 366 -566 0 net=5791
rlabel metal2 478 -566 478 -566 0 net=10421
rlabel metal2 198 -568 198 -568 0 net=2355
rlabel metal2 366 -568 366 -568 0 net=3107
rlabel metal2 485 -568 485 -568 0 net=6129
rlabel metal2 758 -568 758 -568 0 net=7981
rlabel metal2 884 -568 884 -568 0 net=8475
rlabel metal2 954 -568 954 -568 0 net=9965
rlabel metal2 1034 -568 1034 -568 0 net=10295
rlabel metal2 1108 -568 1108 -568 0 net=11707
rlabel metal2 1171 -568 1171 -568 0 net=12209
rlabel metal2 1192 -568 1192 -568 0 net=12399
rlabel metal2 226 -570 226 -570 0 net=1749
rlabel metal2 495 -570 495 -570 0 net=6107
rlabel metal2 761 -570 761 -570 0 net=10753
rlabel metal2 1199 -570 1199 -570 0 net=12455
rlabel metal2 247 -572 247 -572 0 net=1843
rlabel metal2 506 -572 506 -572 0 net=5357
rlabel metal2 562 -572 562 -572 0 net=5271
rlabel metal2 828 -572 828 -572 0 net=7517
rlabel metal2 891 -572 891 -572 0 net=9411
rlabel metal2 1031 -572 1031 -572 0 net=10355
rlabel metal2 1206 -572 1206 -572 0 net=12465
rlabel metal2 303 -574 303 -574 0 net=1905
rlabel metal2 786 -574 786 -574 0 net=7135
rlabel metal2 835 -574 835 -574 0 net=8025
rlabel metal2 926 -574 926 -574 0 net=8961
rlabel metal2 961 -574 961 -574 0 net=10055
rlabel metal2 1080 -574 1080 -574 0 net=11231
rlabel metal2 310 -576 310 -576 0 net=2655
rlabel metal2 481 -576 481 -576 0 net=8395
rlabel metal2 968 -576 968 -576 0 net=10225
rlabel metal2 1213 -576 1213 -576 0 net=12639
rlabel metal2 240 -578 240 -578 0 net=4859
rlabel metal2 324 -578 324 -578 0 net=10997
rlabel metal2 1136 -578 1136 -578 0 net=12305
rlabel metal2 240 -580 240 -580 0 net=2126
rlabel metal2 331 -580 331 -580 0 net=1879
rlabel metal2 492 -580 492 -580 0 net=3913
rlabel metal2 723 -580 723 -580 0 net=7387
rlabel metal2 842 -580 842 -580 0 net=7719
rlabel metal2 940 -580 940 -580 0 net=9071
rlabel metal2 975 -580 975 -580 0 net=9947
rlabel metal2 1150 -580 1150 -580 0 net=12143
rlabel metal2 261 -582 261 -582 0 net=1943
rlabel metal2 317 -582 317 -582 0 net=1992
rlabel metal2 499 -582 499 -582 0 net=5567
rlabel metal2 79 -584 79 -584 0 net=7794
rlabel metal2 275 -584 275 -584 0 net=2535
rlabel metal2 576 -584 576 -584 0 net=7925
rlabel metal2 982 -584 982 -584 0 net=10071
rlabel metal2 79 -586 79 -586 0 net=5811
rlabel metal2 639 -586 639 -586 0 net=6435
rlabel metal2 824 -586 824 -586 0 net=10173
rlabel metal2 1101 -586 1101 -586 0 net=10577
rlabel metal2 275 -588 275 -588 0 net=1873
rlabel metal2 436 -588 436 -588 0 net=5321
rlabel metal2 639 -588 639 -588 0 net=7278
rlabel metal2 870 -588 870 -588 0 net=9029
rlabel metal2 996 -588 996 -588 0 net=10311
rlabel metal2 51 -590 51 -590 0 net=4568
rlabel metal2 467 -590 467 -590 0 net=9901
rlabel metal2 51 -592 51 -592 0 net=7027
rlabel metal2 289 -592 289 -592 0 net=4613
rlabel metal2 562 -592 562 -592 0 net=4519
rlabel metal2 912 -592 912 -592 0 net=9345
rlabel metal2 1038 -592 1038 -592 0 net=10543
rlabel metal2 107 -594 107 -594 0 net=4577
rlabel metal2 681 -594 681 -594 0 net=9589
rlabel metal2 1045 -594 1045 -594 0 net=10645
rlabel metal2 170 -596 170 -596 0 net=4355
rlabel metal2 390 -596 390 -596 0 net=9423
rlabel metal2 1052 -596 1052 -596 0 net=10691
rlabel metal2 772 -598 772 -598 0 net=8765
rlabel metal2 814 -598 814 -598 0 net=8383
rlabel metal2 947 -598 947 -598 0 net=9683
rlabel metal2 1059 -598 1059 -598 0 net=10855
rlabel metal2 607 -600 607 -600 0 net=6891
rlabel metal2 845 -600 845 -600 0 net=10783
rlabel metal2 695 -602 695 -602 0 net=9777
rlabel metal2 695 -604 695 -604 0 net=9907
rlabel metal2 737 -606 737 -606 0 net=7103
rlabel metal2 845 -606 845 -606 0 net=9775
rlabel metal2 604 -608 604 -608 0 net=6185
rlabel metal2 779 -608 779 -608 0 net=9601
rlabel metal2 464 -610 464 -610 0 net=284
rlabel metal2 779 -610 779 -610 0 net=5795
rlabel metal2 877 -610 877 -610 0 net=8813
rlabel metal2 408 -612 408 -612 0 net=3035
rlabel metal2 793 -612 793 -612 0 net=7823
rlabel metal2 338 -614 338 -614 0 net=2005
rlabel metal2 338 -616 338 -616 0 net=2113
rlabel metal2 404 -616 404 -616 0 net=6807
rlabel metal2 212 -618 212 -618 0 net=1560
rlabel metal2 212 -620 212 -620 0 net=6227
rlabel metal2 387 -622 387 -622 0 net=4253
rlabel metal2 65 -633 65 -633 0 net=2854
rlabel metal2 310 -633 310 -633 0 net=4860
rlabel metal2 334 -633 334 -633 0 net=215
rlabel metal2 523 -633 523 -633 0 net=3782
rlabel metal2 618 -633 618 -633 0 net=4866
rlabel metal2 691 -633 691 -633 0 net=5796
rlabel metal2 786 -633 786 -633 0 net=11702
rlabel metal2 1419 -633 1419 -633 0 net=11548
rlabel metal2 1549 -633 1549 -633 0 net=11579
rlabel metal2 1619 -633 1619 -633 0 net=7747
rlabel metal2 72 -635 72 -635 0 net=6999
rlabel metal2 646 -635 646 -635 0 net=4421
rlabel metal2 1528 -635 1528 -635 0 net=8921
rlabel metal2 68 -637 68 -637 0 net=4651
rlabel metal2 100 -637 100 -637 0 net=3281
rlabel metal2 100 -637 100 -637 0 net=3281
rlabel metal2 121 -637 121 -637 0 net=2076
rlabel metal2 649 -637 649 -637 0 net=8766
rlabel metal2 831 -637 831 -637 0 net=12640
rlabel metal2 1444 -637 1444 -637 0 net=12523
rlabel metal2 1465 -637 1465 -637 0 net=7997
rlabel metal2 121 -639 121 -639 0 net=6229
rlabel metal2 222 -639 222 -639 0 net=10422
rlabel metal2 1276 -639 1276 -639 0 net=11375
rlabel metal2 128 -641 128 -641 0 net=3188
rlabel metal2 240 -641 240 -641 0 net=493
rlabel metal2 485 -641 485 -641 0 net=5813
rlabel metal2 838 -641 838 -641 0 net=9948
rlabel metal2 1360 -641 1360 -641 0 net=12273
rlabel metal2 1437 -641 1437 -641 0 net=12509
rlabel metal2 128 -643 128 -643 0 net=1945
rlabel metal2 296 -643 296 -643 0 net=3093
rlabel metal2 429 -643 429 -643 0 net=2589
rlabel metal2 548 -643 548 -643 0 net=4563
rlabel metal2 548 -643 548 -643 0 net=4563
rlabel metal2 555 -643 555 -643 0 net=7092
rlabel metal2 674 -643 674 -643 0 net=10563
rlabel metal2 1423 -643 1423 -643 0 net=12473
rlabel metal2 159 -645 159 -645 0 net=7926
rlabel metal2 982 -645 982 -645 0 net=9425
rlabel metal2 1164 -645 1164 -645 0 net=11709
rlabel metal2 117 -647 117 -647 0 net=7949
rlabel metal2 1017 -647 1017 -647 0 net=10528
rlabel metal2 79 -649 79 -649 0 net=8455
rlabel metal2 1052 -649 1052 -649 0 net=10785
rlabel metal2 1318 -649 1318 -649 0 net=12129
rlabel metal2 58 -651 58 -651 0 net=5829
rlabel metal2 191 -651 191 -651 0 net=4907
rlabel metal2 674 -651 674 -651 0 net=9776
rlabel metal2 93 -653 93 -653 0 net=4735
rlabel metal2 198 -653 198 -653 0 net=9010
rlabel metal2 93 -655 93 -655 0 net=2359
rlabel metal2 198 -655 198 -655 0 net=2567
rlabel metal2 394 -655 394 -655 0 net=5752
rlabel metal2 492 -655 492 -655 0 net=7883
rlabel metal2 1066 -655 1066 -655 0 net=9909
rlabel metal2 1192 -655 1192 -655 0 net=10755
rlabel metal2 114 -657 114 -657 0 net=4880
rlabel metal2 555 -657 555 -657 0 net=7982
rlabel metal2 870 -657 870 -657 0 net=10240
rlabel metal2 44 -659 44 -659 0 net=4496
rlabel metal2 201 -659 201 -659 0 net=11340
rlabel metal2 1255 -659 1255 -659 0 net=11233
rlabel metal2 44 -661 44 -661 0 net=4235
rlabel metal2 457 -661 457 -661 0 net=5043
rlabel metal2 845 -661 845 -661 0 net=12466
rlabel metal2 205 -663 205 -663 0 net=4795
rlabel metal2 247 -663 247 -663 0 net=1845
rlabel metal2 345 -663 345 -663 0 net=2356
rlabel metal2 590 -663 590 -663 0 net=3443
rlabel metal2 709 -663 709 -663 0 net=6785
rlabel metal2 800 -663 800 -663 0 net=11481
rlabel metal2 149 -665 149 -665 0 net=1537
rlabel metal2 282 -665 282 -665 0 net=3389
rlabel metal2 296 -665 296 -665 0 net=1881
rlabel metal2 345 -665 345 -665 0 net=2303
rlabel metal2 677 -665 677 -665 0 net=9874
rlabel metal2 149 -667 149 -667 0 net=6629
rlabel metal2 758 -667 758 -667 0 net=8858
rlabel metal2 212 -669 212 -669 0 net=3497
rlabel metal2 226 -669 226 -669 0 net=1750
rlabel metal2 495 -669 495 -669 0 net=6697
rlabel metal2 926 -669 926 -669 0 net=8397
rlabel metal2 1108 -669 1108 -669 0 net=10313
rlabel metal2 219 -671 219 -671 0 net=109
rlabel metal2 803 -671 803 -671 0 net=12123
rlabel metal2 1395 -671 1395 -671 0 net=12457
rlabel metal2 226 -673 226 -673 0 net=3631
rlabel metal2 275 -673 275 -673 0 net=1875
rlabel metal2 310 -673 310 -673 0 net=3109
rlabel metal2 478 -673 478 -673 0 net=2699
rlabel metal2 569 -673 569 -673 0 net=4477
rlabel metal2 653 -673 653 -673 0 net=5739
rlabel metal2 828 -673 828 -673 0 net=7137
rlabel metal2 933 -673 933 -673 0 net=8477
rlabel metal2 1038 -673 1038 -673 0 net=9603
rlabel metal2 1206 -673 1206 -673 0 net=12307
rlabel metal2 1283 -673 1283 -673 0 net=11779
rlabel metal2 1304 -673 1304 -673 0 net=11903
rlabel metal2 170 -675 170 -675 0 net=4357
rlabel metal2 471 -675 471 -675 0 net=5451
rlabel metal2 681 -675 681 -675 0 net=6187
rlabel metal2 744 -675 744 -675 0 net=10226
rlabel metal2 1220 -675 1220 -675 0 net=10841
rlabel metal2 142 -677 142 -677 0 net=3399
rlabel metal2 527 -677 527 -677 0 net=4185
rlabel metal2 590 -677 590 -677 0 net=6419
rlabel metal2 632 -677 632 -677 0 net=6023
rlabel metal2 751 -677 751 -677 0 net=8279
rlabel metal2 912 -677 912 -677 0 net=8385
rlabel metal2 961 -677 961 -677 0 net=9031
rlabel metal2 1122 -677 1122 -677 0 net=10999
rlabel metal2 142 -679 142 -679 0 net=4579
rlabel metal2 527 -679 527 -679 0 net=9590
rlabel metal2 1059 -679 1059 -679 0 net=9779
rlabel metal2 1248 -679 1248 -679 0 net=10845
rlabel metal2 156 -681 156 -681 0 net=8629
rlabel metal2 1080 -681 1080 -681 0 net=10175
rlabel metal2 1262 -681 1262 -681 0 net=11259
rlabel metal2 170 -683 170 -683 0 net=2747
rlabel metal2 597 -683 597 -683 0 net=5273
rlabel metal2 632 -683 632 -683 0 net=8508
rlabel metal2 1129 -683 1129 -683 0 net=10545
rlabel metal2 184 -685 184 -685 0 net=5896
rlabel metal2 604 -685 604 -685 0 net=5568
rlabel metal2 184 -687 184 -687 0 net=1907
rlabel metal2 317 -687 317 -687 0 net=2536
rlabel metal2 425 -687 425 -687 0 net=5197
rlabel metal2 761 -687 761 -687 0 net=8869
rlabel metal2 1087 -687 1087 -687 0 net=8701
rlabel metal2 1136 -687 1136 -687 0 net=10857
rlabel metal2 86 -689 86 -689 0 net=4133
rlabel metal2 558 -689 558 -689 0 net=4359
rlabel metal2 604 -689 604 -689 0 net=9952
rlabel metal2 86 -691 86 -691 0 net=4417
rlabel metal2 233 -691 233 -691 0 net=2475
rlabel metal2 355 -691 355 -691 0 net=3533
rlabel metal2 530 -691 530 -691 0 net=11521
rlabel metal2 107 -693 107 -693 0 net=3843
rlabel metal2 821 -693 821 -693 0 net=7259
rlabel metal2 1094 -693 1094 -693 0 net=10297
rlabel metal2 254 -695 254 -695 0 net=2287
rlabel metal2 359 -695 359 -695 0 net=3037
rlabel metal2 688 -695 688 -695 0 net=6109
rlabel metal2 814 -695 814 -695 0 net=7105
rlabel metal2 828 -695 828 -695 0 net=12669
rlabel metal2 177 -697 177 -697 0 net=6479
rlabel metal2 849 -697 849 -697 0 net=7635
rlabel metal2 954 -697 954 -697 0 net=8963
rlabel metal2 1150 -697 1150 -697 0 net=10579
rlabel metal2 177 -699 177 -699 0 net=2499
rlabel metal2 380 -699 380 -699 0 net=2897
rlabel metal2 464 -699 464 -699 0 net=842
rlabel metal2 254 -701 254 -701 0 net=2503
rlabel metal2 429 -701 429 -701 0 net=7683
rlabel metal2 968 -701 968 -701 0 net=9073
rlabel metal2 1178 -701 1178 -701 0 net=10693
rlabel metal2 1388 -701 1388 -701 0 net=12443
rlabel metal2 261 -703 261 -703 0 net=2115
rlabel metal2 467 -703 467 -703 0 net=7771
rlabel metal2 989 -703 989 -703 0 net=9287
rlabel metal2 1178 -703 1178 -703 0 net=12401
rlabel metal2 268 -705 268 -705 0 net=3199
rlabel metal2 702 -705 702 -705 0 net=6131
rlabel metal2 719 -705 719 -705 0 net=12078
rlabel metal2 268 -707 268 -707 0 net=2671
rlabel metal2 460 -707 460 -707 0 net=8197
rlabel metal2 730 -707 730 -707 0 net=8509
rlabel metal2 1185 -707 1185 -707 0 net=12211
rlabel metal2 135 -709 135 -709 0 net=4081
rlabel metal2 684 -709 684 -709 0 net=10033
rlabel metal2 1311 -709 1311 -709 0 net=12045
rlabel metal2 135 -711 135 -711 0 net=4057
rlabel metal2 303 -711 303 -711 0 net=2657
rlabel metal2 733 -711 733 -711 0 net=9902
rlabel metal2 1346 -711 1346 -711 0 net=12145
rlabel metal2 317 -713 317 -713 0 net=2007
rlabel metal2 415 -713 415 -713 0 net=4615
rlabel metal2 733 -713 733 -713 0 net=10072
rlabel metal2 163 -715 163 -715 0 net=3815
rlabel metal2 499 -715 499 -715 0 net=5323
rlabel metal2 793 -715 793 -715 0 net=6809
rlabel metal2 873 -715 873 -715 0 net=11465
rlabel metal2 58 -717 58 -717 0 net=2211
rlabel metal2 331 -717 331 -717 0 net=3759
rlabel metal2 576 -717 576 -717 0 net=6247
rlabel metal2 884 -717 884 -717 0 net=7519
rlabel metal2 919 -717 919 -717 0 net=7721
rlabel metal2 989 -717 989 -717 0 net=8091
rlabel metal2 1045 -717 1045 -717 0 net=9685
rlabel metal2 1171 -717 1171 -717 0 net=10647
rlabel metal2 275 -719 275 -719 0 net=1777
rlabel metal2 877 -719 877 -719 0 net=7825
rlabel metal2 432 -721 432 -721 0 net=6951
rlabel metal2 891 -721 891 -721 0 net=8027
rlabel metal2 929 -721 929 -721 0 net=9005
rlabel metal2 51 -723 51 -723 0 net=7029
rlabel metal2 905 -723 905 -723 0 net=10356
rlabel metal2 51 -725 51 -725 0 net=5381
rlabel metal2 436 -725 436 -725 0 net=3049
rlabel metal2 1073 -725 1073 -725 0 net=10057
rlabel metal2 642 -727 642 -727 0 net=8665
rlabel metal2 807 -729 807 -729 0 net=6893
rlabel metal2 908 -729 908 -729 0 net=11683
rlabel metal2 723 -731 723 -731 0 net=6437
rlabel metal2 996 -731 996 -731 0 net=9347
rlabel metal2 506 -733 506 -733 0 net=5359
rlabel metal2 947 -733 947 -733 0 net=8815
rlabel metal2 1003 -733 1003 -733 0 net=9967
rlabel metal2 257 -735 257 -735 0 net=3607
rlabel metal2 520 -735 520 -735 0 net=5733
rlabel metal2 1010 -735 1010 -735 0 net=9413
rlabel metal2 863 -737 863 -737 0 net=7675
rlabel metal2 1020 -737 1020 -737 0 net=10671
rlabel metal2 765 -739 765 -739 0 net=6883
rlabel metal2 898 -739 898 -739 0 net=8181
rlabel metal2 443 -741 443 -741 0 net=5793
rlabel metal2 835 -741 835 -741 0 net=7389
rlabel metal2 443 -743 443 -743 0 net=5983
rlabel metal2 835 -743 835 -743 0 net=12064
rlabel metal2 660 -745 660 -745 0 net=4697
rlabel metal2 1241 -745 1241 -745 0 net=11957
rlabel metal2 583 -747 583 -747 0 net=4803
rlabel metal2 698 -747 698 -747 0 net=10591
rlabel metal2 541 -749 541 -749 0 net=4255
rlabel metal2 513 -751 513 -751 0 net=3915
rlabel metal2 513 -753 513 -753 0 net=4521
rlabel metal2 562 -755 562 -755 0 net=5523
rlabel metal2 37 -766 37 -766 0 net=5383
rlabel metal2 58 -766 58 -766 0 net=5525
rlabel metal2 572 -766 572 -766 0 net=12130
rlabel metal2 1430 -766 1430 -766 0 net=11001
rlabel metal2 1696 -766 1696 -766 0 net=7749
rlabel metal2 44 -768 44 -768 0 net=4236
rlabel metal2 485 -768 485 -768 0 net=2590
rlabel metal2 551 -768 551 -768 0 net=5198
rlabel metal2 793 -768 793 -768 0 net=9604
rlabel metal2 1255 -768 1255 -768 0 net=12309
rlabel metal2 1549 -768 1549 -768 0 net=8923
rlabel metal2 44 -770 44 -770 0 net=3415
rlabel metal2 65 -770 65 -770 0 net=2304
rlabel metal2 366 -770 366 -770 0 net=4358
rlabel metal2 667 -770 667 -770 0 net=4804
rlabel metal2 737 -770 737 -770 0 net=7677
rlabel metal2 954 -770 954 -770 0 net=7685
rlabel metal2 954 -770 954 -770 0 net=7685
rlabel metal2 961 -770 961 -770 0 net=7723
rlabel metal2 1297 -770 1297 -770 0 net=11235
rlabel metal2 1297 -770 1297 -770 0 net=11235
rlabel metal2 1332 -770 1332 -770 0 net=11523
rlabel metal2 1332 -770 1332 -770 0 net=11523
rlabel metal2 1353 -770 1353 -770 0 net=11959
rlabel metal2 1437 -770 1437 -770 0 net=12475
rlabel metal2 1528 -770 1528 -770 0 net=7999
rlabel metal2 65 -772 65 -772 0 net=4653
rlabel metal2 114 -772 114 -772 0 net=3039
rlabel metal2 366 -772 366 -772 0 net=4523
rlabel metal2 530 -772 530 -772 0 net=4564
rlabel metal2 558 -772 558 -772 0 net=7260
rlabel metal2 1108 -772 1108 -772 0 net=9033
rlabel metal2 1108 -772 1108 -772 0 net=9033
rlabel metal2 1115 -772 1115 -772 0 net=9075
rlabel metal2 1262 -772 1262 -772 0 net=10695
rlabel metal2 1409 -772 1409 -772 0 net=12275
rlabel metal2 1556 -772 1556 -772 0 net=11580
rlabel metal2 1556 -772 1556 -772 0 net=11580
rlabel metal2 72 -774 72 -774 0 net=2361
rlabel metal2 124 -774 124 -774 0 net=1876
rlabel metal2 296 -774 296 -774 0 net=1882
rlabel metal2 607 -774 607 -774 0 net=5814
rlabel metal2 793 -774 793 -774 0 net=6895
rlabel metal2 905 -774 905 -774 0 net=11479
rlabel metal2 1444 -774 1444 -774 0 net=12511
rlabel metal2 93 -776 93 -776 0 net=1909
rlabel metal2 187 -776 187 -776 0 net=3110
rlabel metal2 324 -776 324 -776 0 net=1847
rlabel metal2 380 -776 380 -776 0 net=3761
rlabel metal2 604 -776 604 -776 0 net=7217
rlabel metal2 908 -776 908 -776 0 net=10842
rlabel metal2 1367 -776 1367 -776 0 net=12047
rlabel metal2 1458 -776 1458 -776 0 net=12525
rlabel metal2 135 -778 135 -778 0 net=4058
rlabel metal2 345 -778 345 -778 0 net=2289
rlabel metal2 380 -778 380 -778 0 net=5045
rlabel metal2 478 -778 478 -778 0 net=2701
rlabel metal2 534 -778 534 -778 0 net=4187
rlabel metal2 611 -778 611 -778 0 net=4478
rlabel metal2 684 -778 684 -778 0 net=500
rlabel metal2 926 -778 926 -778 0 net=12402
rlabel metal2 1220 -778 1220 -778 0 net=10547
rlabel metal2 1290 -778 1290 -778 0 net=11781
rlabel metal2 1416 -778 1416 -778 0 net=12445
rlabel metal2 135 -780 135 -780 0 net=1735
rlabel metal2 163 -780 163 -780 0 net=2213
rlabel metal2 394 -780 394 -780 0 net=3535
rlabel metal2 506 -780 506 -780 0 net=3608
rlabel metal2 835 -780 835 -780 0 net=7138
rlabel metal2 926 -780 926 -780 0 net=8093
rlabel metal2 1017 -780 1017 -780 0 net=8457
rlabel metal2 1115 -780 1115 -780 0 net=10593
rlabel metal2 1346 -780 1346 -780 0 net=11685
rlabel metal2 1374 -780 1374 -780 0 net=12125
rlabel metal2 1472 -780 1472 -780 0 net=12671
rlabel metal2 163 -782 163 -782 0 net=1106
rlabel metal2 796 -782 796 -782 0 net=9414
rlabel metal2 1150 -782 1150 -782 0 net=9687
rlabel metal2 1150 -782 1150 -782 0 net=9687
rlabel metal2 1157 -782 1157 -782 0 net=9781
rlabel metal2 1157 -782 1157 -782 0 net=9781
rlabel metal2 1171 -782 1171 -782 0 net=9969
rlabel metal2 1171 -782 1171 -782 0 net=9969
rlabel metal2 1178 -782 1178 -782 0 net=10177
rlabel metal2 1213 -782 1213 -782 0 net=10299
rlabel metal2 1227 -782 1227 -782 0 net=10565
rlabel metal2 1479 -782 1479 -782 0 net=4422
rlabel metal2 117 -784 117 -784 0 net=9447
rlabel metal2 1241 -784 1241 -784 0 net=10787
rlabel metal2 1311 -784 1311 -784 0 net=11467
rlabel metal2 1486 -784 1486 -784 0 net=11377
rlabel metal2 166 -786 166 -786 0 net=1402
rlabel metal2 688 -786 688 -786 0 net=7826
rlabel metal2 1059 -786 1059 -786 0 net=8631
rlabel metal2 184 -788 184 -788 0 net=5734
rlabel metal2 1024 -788 1024 -788 0 net=10815
rlabel metal2 191 -790 191 -790 0 net=4736
rlabel metal2 485 -790 485 -790 0 net=3263
rlabel metal2 849 -790 849 -790 0 net=6811
rlabel metal2 929 -790 929 -790 0 net=8398
rlabel metal2 1094 -790 1094 -790 0 net=9007
rlabel metal2 1248 -790 1248 -790 0 net=10673
rlabel metal2 191 -792 191 -792 0 net=3067
rlabel metal2 569 -792 569 -792 0 net=3825
rlabel metal2 1080 -792 1080 -792 0 net=8871
rlabel metal2 1199 -792 1199 -792 0 net=10059
rlabel metal2 205 -794 205 -794 0 net=5794
rlabel metal2 772 -794 772 -794 0 net=6439
rlabel metal2 828 -794 828 -794 0 net=12331
rlabel metal2 208 -796 208 -796 0 net=10327
rlabel metal2 1248 -796 1248 -796 0 net=11261
rlabel metal2 208 -798 208 -798 0 net=5360
rlabel metal2 751 -798 751 -798 0 net=8281
rlabel metal2 1027 -798 1027 -798 0 net=12233
rlabel metal2 226 -800 226 -800 0 net=3633
rlabel metal2 352 -800 352 -800 0 net=3079
rlabel metal2 527 -800 527 -800 0 net=10241
rlabel metal2 212 -802 212 -802 0 net=3499
rlabel metal2 240 -802 240 -802 0 net=4797
rlabel metal2 296 -802 296 -802 0 net=2265
rlabel metal2 534 -802 534 -802 0 net=5740
rlabel metal2 800 -802 800 -802 0 net=8897
rlabel metal2 212 -804 212 -804 0 net=3051
rlabel metal2 457 -804 457 -804 0 net=5087
rlabel metal2 541 -804 541 -804 0 net=3917
rlabel metal2 1045 -804 1045 -804 0 net=8965
rlabel metal2 233 -806 233 -806 0 net=2477
rlabel metal2 464 -806 464 -806 0 net=3401
rlabel metal2 576 -806 576 -806 0 net=6249
rlabel metal2 786 -806 786 -806 0 net=6111
rlabel metal2 807 -806 807 -806 0 net=6885
rlabel metal2 940 -806 940 -806 0 net=7637
rlabel metal2 961 -806 961 -806 0 net=10858
rlabel metal2 121 -808 121 -808 0 net=6231
rlabel metal2 821 -808 821 -808 0 net=7107
rlabel metal2 975 -808 975 -808 0 net=7885
rlabel metal2 1059 -808 1059 -808 0 net=9289
rlabel metal2 233 -810 233 -810 0 net=5753
rlabel metal2 415 -810 415 -810 0 net=4616
rlabel metal2 583 -810 583 -810 0 net=4257
rlabel metal2 632 -810 632 -810 0 net=4605
rlabel metal2 702 -810 702 -810 0 net=8199
rlabel metal2 814 -810 814 -810 0 net=6481
rlabel metal2 838 -810 838 -810 0 net=11271
rlabel metal2 142 -812 142 -812 0 net=4580
rlabel metal2 583 -812 583 -812 0 net=6189
rlabel metal2 709 -812 709 -812 0 net=6133
rlabel metal2 814 -812 814 -812 0 net=12089
rlabel metal2 142 -814 142 -814 0 net=7031
rlabel metal2 968 -814 968 -814 0 net=7773
rlabel metal2 982 -814 982 -814 0 net=7951
rlabel metal2 996 -814 996 -814 0 net=8817
rlabel metal2 1122 -814 1122 -814 0 net=8703
rlabel metal2 79 -816 79 -816 0 net=5831
rlabel metal2 919 -816 919 -816 0 net=8029
rlabel metal2 1073 -816 1073 -816 0 net=8667
rlabel metal2 1122 -816 1122 -816 0 net=9349
rlabel metal2 79 -818 79 -818 0 net=4419
rlabel metal2 156 -818 156 -818 0 net=2801
rlabel metal2 716 -818 716 -818 0 net=7243
rlabel metal2 982 -818 982 -818 0 net=8183
rlabel metal2 1052 -818 1052 -818 0 net=8511
rlabel metal2 1136 -818 1136 -818 0 net=9427
rlabel metal2 86 -820 86 -820 0 net=3283
rlabel metal2 240 -820 240 -820 0 net=4135
rlabel metal2 401 -820 401 -820 0 net=4083
rlabel metal2 590 -820 590 -820 0 net=6421
rlabel metal2 863 -820 863 -820 0 net=6953
rlabel metal2 933 -820 933 -820 0 net=8387
rlabel metal2 1031 -820 1031 -820 0 net=8479
rlabel metal2 100 -822 100 -822 0 net=5985
rlabel metal2 509 -822 509 -822 0 net=11581
rlabel metal2 152 -824 152 -824 0 net=5115
rlabel metal2 590 -824 590 -824 0 net=7001
rlabel metal2 646 -824 646 -824 0 net=10314
rlabel metal2 149 -826 149 -826 0 net=6631
rlabel metal2 649 -826 649 -826 0 net=12321
rlabel metal2 51 -828 51 -828 0 net=6835
rlabel metal2 261 -828 261 -828 0 net=2117
rlabel metal2 338 -828 338 -828 0 net=3201
rlabel metal2 401 -828 401 -828 0 net=3095
rlabel metal2 429 -828 429 -828 0 net=1
rlabel metal2 744 -828 744 -828 0 net=6025
rlabel metal2 912 -828 912 -828 0 net=7521
rlabel metal2 1381 -828 1381 -828 0 net=12147
rlabel metal2 170 -830 170 -830 0 net=2749
rlabel metal2 373 -830 373 -830 0 net=2505
rlabel metal2 499 -830 499 -830 0 net=5325
rlabel metal2 838 -830 838 -830 0 net=10648
rlabel metal2 170 -832 170 -832 0 net=2569
rlabel metal2 247 -832 247 -832 0 net=1539
rlabel metal2 282 -832 282 -832 0 net=3391
rlabel metal2 408 -832 408 -832 0 net=3817
rlabel metal2 625 -832 625 -832 0 net=5275
rlabel metal2 1283 -832 1283 -832 0 net=10847
rlabel metal2 121 -834 121 -834 0 net=4197
rlabel metal2 303 -834 303 -834 0 net=2659
rlabel metal2 422 -834 422 -834 0 net=4509
rlabel metal2 877 -834 877 -834 0 net=9557
rlabel metal2 1269 -834 1269 -834 0 net=10757
rlabel metal2 1360 -834 1360 -834 0 net=11711
rlabel metal2 128 -836 128 -836 0 net=1947
rlabel metal2 268 -836 268 -836 0 net=2673
rlabel metal2 317 -836 317 -836 0 net=2009
rlabel metal2 499 -836 499 -836 0 net=11185
rlabel metal2 128 -838 128 -838 0 net=2501
rlabel metal2 198 -838 198 -838 0 net=3387
rlabel metal2 268 -838 268 -838 0 net=4005
rlabel metal2 873 -838 873 -838 0 net=12458
rlabel metal2 177 -840 177 -840 0 net=1779
rlabel metal2 317 -840 317 -840 0 net=2899
rlabel metal2 635 -840 635 -840 0 net=5573
rlabel metal2 831 -840 831 -840 0 net=11904
rlabel metal2 107 -842 107 -842 0 net=3845
rlabel metal2 649 -842 649 -842 0 net=5337
rlabel metal2 880 -842 880 -842 0 net=11121
rlabel metal2 107 -844 107 -844 0 net=9697
rlabel metal2 254 -846 254 -846 0 net=2789
rlabel metal2 373 -846 373 -846 0 net=1789
rlabel metal2 898 -846 898 -846 0 net=7391
rlabel metal2 919 -846 919 -846 0 net=8391
rlabel metal2 1164 -846 1164 -846 0 net=9911
rlabel metal2 1388 -846 1388 -846 0 net=12213
rlabel metal2 159 -848 159 -848 0 net=7157
rlabel metal2 1185 -848 1185 -848 0 net=10035
rlabel metal2 520 -850 520 -850 0 net=10195
rlabel metal2 1234 -850 1234 -850 0 net=10581
rlabel metal2 520 -852 520 -852 0 net=3635
rlabel metal2 653 -852 653 -852 0 net=5453
rlabel metal2 870 -852 870 -852 0 net=9929
rlabel metal2 1234 -852 1234 -852 0 net=11483
rlabel metal2 653 -854 653 -854 0 net=5027
rlabel metal2 691 -854 691 -854 0 net=11307
rlabel metal2 660 -856 660 -856 0 net=4699
rlabel metal2 751 -856 751 -856 0 net=5161
rlabel metal2 660 -858 660 -858 0 net=3445
rlabel metal2 618 -860 618 -860 0 net=4909
rlabel metal2 597 -862 597 -862 0 net=4361
rlabel metal2 597 -864 597 -864 0 net=6699
rlabel metal2 779 -866 779 -866 0 net=6787
rlabel metal2 471 -868 471 -868 0 net=3161
rlabel metal2 30 -879 30 -879 0 net=7033
rlabel metal2 149 -879 149 -879 0 net=5832
rlabel metal2 919 -879 919 -879 0 net=12214
rlabel metal2 1458 -879 1458 -879 0 net=12091
rlabel metal2 1458 -879 1458 -879 0 net=12091
rlabel metal2 1500 -879 1500 -879 0 net=12447
rlabel metal2 1500 -879 1500 -879 0 net=12447
rlabel metal2 1542 -879 1542 -879 0 net=11378
rlabel metal2 1570 -879 1570 -879 0 net=8001
rlabel metal2 1724 -879 1724 -879 0 net=7751
rlabel metal2 44 -881 44 -881 0 net=3416
rlabel metal2 656 -881 656 -881 0 net=454
rlabel metal2 1577 -881 1577 -881 0 net=8925
rlabel metal2 44 -883 44 -883 0 net=6837
rlabel metal2 79 -883 79 -883 0 net=4420
rlabel metal2 660 -883 660 -883 0 net=3446
rlabel metal2 838 -883 838 -883 0 net=1418
rlabel metal2 873 -883 873 -883 0 net=9076
rlabel metal2 1318 -883 1318 -883 0 net=11309
rlabel metal2 51 -885 51 -885 0 net=4655
rlabel metal2 79 -885 79 -885 0 net=2502
rlabel metal2 135 -885 135 -885 0 net=1737
rlabel metal2 166 -885 166 -885 0 net=9912
rlabel metal2 1521 -885 1521 -885 0 net=12673
rlabel metal2 1573 -885 1573 -885 0 net=4173
rlabel metal2 1584 -885 1584 -885 0 net=11003
rlabel metal2 65 -887 65 -887 0 net=2363
rlabel metal2 82 -887 82 -887 0 net=5754
rlabel metal2 257 -887 257 -887 0 net=11480
rlabel metal2 1479 -887 1479 -887 0 net=11469
rlabel metal2 72 -889 72 -889 0 net=3285
rlabel metal2 93 -889 93 -889 0 net=1910
rlabel metal2 208 -889 208 -889 0 net=3080
rlabel metal2 408 -889 408 -889 0 net=890
rlabel metal2 660 -889 660 -889 0 net=6813
rlabel metal2 880 -889 880 -889 0 net=12276
rlabel metal2 58 -891 58 -891 0 net=5527
rlabel metal2 93 -891 93 -891 0 net=3827
rlabel metal2 667 -891 667 -891 0 net=7108
rlabel metal2 964 -891 964 -891 0 net=12126
rlabel metal2 1437 -891 1437 -891 0 net=12049
rlabel metal2 1479 -891 1479 -891 0 net=12323
rlabel metal2 1493 -891 1493 -891 0 net=12333
rlabel metal2 58 -893 58 -893 0 net=4511
rlabel metal2 436 -893 436 -893 0 net=2478
rlabel metal2 667 -893 667 -893 0 net=4701
rlabel metal2 775 -893 775 -893 0 net=9008
rlabel metal2 1346 -893 1346 -893 0 net=8632
rlabel metal2 100 -895 100 -895 0 net=5986
rlabel metal2 985 -895 985 -895 0 net=10848
rlabel metal2 1388 -895 1388 -895 0 net=10037
rlabel metal2 1465 -895 1465 -895 0 net=12149
rlabel metal2 1514 -895 1514 -895 0 net=12527
rlabel metal2 100 -897 100 -897 0 net=4155
rlabel metal2 891 -897 891 -897 0 net=7687
rlabel metal2 961 -897 961 -897 0 net=12697
rlabel metal2 107 -899 107 -899 0 net=2266
rlabel metal2 317 -899 317 -899 0 net=2901
rlabel metal2 331 -899 331 -899 0 net=2215
rlabel metal2 331 -899 331 -899 0 net=2215
rlabel metal2 338 -899 338 -899 0 net=2750
rlabel metal2 502 -899 502 -899 0 net=5276
rlabel metal2 992 -899 992 -899 0 net=12079
rlabel metal2 1465 -899 1465 -899 0 net=12477
rlabel metal2 107 -901 107 -901 0 net=3053
rlabel metal2 219 -901 219 -901 0 net=7839
rlabel metal2 548 -901 548 -901 0 net=7002
rlabel metal2 674 -901 674 -901 0 net=6026
rlabel metal2 905 -901 905 -901 0 net=7219
rlabel metal2 926 -901 926 -901 0 net=8095
rlabel metal2 940 -901 940 -901 0 net=8389
rlabel metal2 1069 -901 1069 -901 0 net=12512
rlabel metal2 110 -903 110 -903 0 net=3634
rlabel metal2 317 -903 317 -903 0 net=2119
rlabel metal2 352 -903 352 -903 0 net=3847
rlabel metal2 502 -903 502 -903 0 net=9698
rlabel metal2 1472 -903 1472 -903 0 net=12235
rlabel metal2 1549 -903 1549 -903 0 net=985
rlabel metal2 121 -905 121 -905 0 net=4524
rlabel metal2 408 -905 408 -905 0 net=8201
rlabel metal2 779 -905 779 -905 0 net=6789
rlabel metal2 856 -905 856 -905 0 net=7775
rlabel metal2 1111 -905 1111 -905 0 net=12361
rlabel metal2 1563 -905 1563 -905 0 net=2369
rlabel metal2 121 -907 121 -907 0 net=9593
rlabel metal2 128 -907 128 -907 0 net=2790
rlabel metal2 289 -907 289 -907 0 net=4799
rlabel metal2 310 -907 310 -907 0 net=3393
rlabel metal2 411 -907 411 -907 0 net=1081
rlabel metal2 926 -907 926 -907 0 net=7523
rlabel metal2 968 -907 968 -907 0 net=7953
rlabel metal2 1129 -907 1129 -907 0 net=8705
rlabel metal2 1129 -907 1129 -907 0 net=8705
rlabel metal2 1171 -907 1171 -907 0 net=9971
rlabel metal2 1248 -907 1248 -907 0 net=11263
rlabel metal2 1409 -907 1409 -907 0 net=11783
rlabel metal2 138 -909 138 -909 0 net=5046
rlabel metal2 394 -909 394 -909 0 net=5339
rlabel metal2 723 -909 723 -909 0 net=6135
rlabel metal2 782 -909 782 -909 0 net=11122
rlabel metal2 163 -911 163 -911 0 net=3667
rlabel metal2 222 -911 222 -911 0 net=1032
rlabel metal2 268 -911 268 -911 0 net=4007
rlabel metal2 446 -911 446 -911 0 net=8767
rlabel metal2 877 -911 877 -911 0 net=7725
rlabel metal2 1248 -911 1248 -911 0 net=10549
rlabel metal2 1290 -911 1290 -911 0 net=11187
rlabel metal2 1367 -911 1367 -911 0 net=11687
rlabel metal2 163 -913 163 -913 0 net=1781
rlabel metal2 191 -913 191 -913 0 net=3069
rlabel metal2 380 -913 380 -913 0 net=6441
rlabel metal2 828 -913 828 -913 0 net=11865
rlabel metal2 1374 -913 1374 -913 0 net=10817
rlabel metal2 177 -915 177 -915 0 net=3203
rlabel metal2 450 -915 450 -915 0 net=2507
rlabel metal2 506 -915 506 -915 0 net=3918
rlabel metal2 1164 -915 1164 -915 0 net=9931
rlabel metal2 1241 -915 1241 -915 0 net=10789
rlabel metal2 1269 -915 1269 -915 0 net=10583
rlabel metal2 1297 -915 1297 -915 0 net=11237
rlabel metal2 1395 -915 1395 -915 0 net=11961
rlabel metal2 191 -917 191 -917 0 net=2703
rlabel metal2 520 -917 520 -917 0 net=11059
rlabel metal2 135 -919 135 -919 0 net=4703
rlabel metal2 523 -919 523 -919 0 net=4910
rlabel metal2 698 -919 698 -919 0 net=8139
rlabel metal2 975 -919 975 -919 0 net=10663
rlabel metal2 1304 -919 1304 -919 0 net=11273
rlabel metal2 198 -921 198 -921 0 net=3388
rlabel metal2 425 -921 425 -921 0 net=3583
rlabel metal2 530 -921 530 -921 0 net=7886
rlabel metal2 1115 -921 1115 -921 0 net=10595
rlabel metal2 198 -923 198 -923 0 net=1541
rlabel metal2 268 -923 268 -923 0 net=2675
rlabel metal2 387 -923 387 -923 0 net=4607
rlabel metal2 670 -923 670 -923 0 net=9361
rlabel metal2 845 -923 845 -923 0 net=12087
rlabel metal2 205 -925 205 -925 0 net=2479
rlabel metal2 492 -925 492 -925 0 net=9021
rlabel metal2 688 -925 688 -925 0 net=10674
rlabel metal2 205 -927 205 -927 0 net=1791
rlabel metal2 509 -927 509 -927 0 net=7199
rlabel metal2 534 -927 534 -927 0 net=3763
rlabel metal2 569 -927 569 -927 0 net=4363
rlabel metal2 625 -927 625 -927 0 net=12237
rlabel metal2 184 -929 184 -929 0 net=6087
rlabel metal2 586 -929 586 -929 0 net=8321
rlabel metal2 1157 -929 1157 -929 0 net=9783
rlabel metal2 1171 -929 1171 -929 0 net=10179
rlabel metal2 1227 -929 1227 -929 0 net=10329
rlabel metal2 1283 -929 1283 -929 0 net=10759
rlabel metal2 149 -931 149 -931 0 net=1579
rlabel metal2 226 -931 226 -931 0 net=3501
rlabel metal2 373 -931 373 -931 0 net=3097
rlabel metal2 506 -931 506 -931 0 net=10555
rlabel metal2 233 -933 233 -933 0 net=3537
rlabel metal2 509 -933 509 -933 0 net=1045
rlabel metal2 590 -933 590 -933 0 net=6483
rlabel metal2 898 -933 898 -933 0 net=7159
rlabel metal2 933 -933 933 -933 0 net=7639
rlabel metal2 999 -933 999 -933 0 net=10735
rlabel metal2 1234 -933 1234 -933 0 net=11485
rlabel metal2 250 -935 250 -935 0 net=3953
rlabel metal2 611 -935 611 -935 0 net=4259
rlabel metal2 674 -935 674 -935 0 net=5455
rlabel metal2 758 -935 758 -935 0 net=6233
rlabel metal2 898 -935 898 -935 0 net=10696
rlabel metal2 254 -937 254 -937 0 net=4199
rlabel metal2 303 -937 303 -937 0 net=2661
rlabel metal2 478 -937 478 -937 0 net=3265
rlabel metal2 527 -937 527 -937 0 net=2779
rlabel metal2 835 -937 835 -937 0 net=11975
rlabel metal2 170 -939 170 -939 0 net=2571
rlabel metal2 401 -939 401 -939 0 net=2011
rlabel metal2 485 -939 485 -939 0 net=5029
rlabel metal2 677 -939 677 -939 0 net=10566
rlabel metal2 156 -941 156 -941 0 net=2803
rlabel metal2 261 -941 261 -941 0 net=2291
rlabel metal2 415 -941 415 -941 0 net=3637
rlabel metal2 604 -941 604 -941 0 net=4189
rlabel metal2 625 -941 625 -941 0 net=8821
rlabel metal2 684 -941 684 -941 0 net=2665
rlabel metal2 800 -941 800 -941 0 net=6113
rlabel metal2 901 -941 901 -941 0 net=10811
rlabel metal2 1325 -941 1325 -941 0 net=11583
rlabel metal2 156 -943 156 -943 0 net=1949
rlabel metal2 275 -943 275 -943 0 net=3163
rlabel metal2 541 -943 541 -943 0 net=3819
rlabel metal2 695 -943 695 -943 0 net=5326
rlabel metal2 768 -943 768 -943 0 net=11071
rlabel metal2 345 -945 345 -945 0 net=1849
rlabel metal2 429 -945 429 -945 0 net=4085
rlabel metal2 597 -945 597 -945 0 net=6701
rlabel metal2 772 -945 772 -945 0 net=5815
rlabel metal2 114 -947 114 -947 0 net=3041
rlabel metal2 457 -947 457 -947 0 net=5089
rlabel metal2 702 -947 702 -947 0 net=5163
rlabel metal2 793 -947 793 -947 0 net=6897
rlabel metal2 1017 -947 1017 -947 0 net=8459
rlabel metal2 1150 -947 1150 -947 0 net=9689
rlabel metal2 1220 -947 1220 -947 0 net=10301
rlabel metal2 114 -949 114 -949 0 net=4137
rlabel metal2 443 -949 443 -949 0 net=5117
rlabel metal2 464 -949 464 -949 0 net=3403
rlabel metal2 562 -949 562 -949 0 net=6251
rlabel metal2 793 -949 793 -949 0 net=6887
rlabel metal2 1024 -949 1024 -949 0 net=8481
rlabel metal2 1108 -949 1108 -949 0 net=9035
rlabel metal2 37 -951 37 -951 0 net=5385
rlabel metal2 443 -951 443 -951 0 net=12139
rlabel metal2 37 -953 37 -953 0 net=6955
rlabel metal2 929 -953 929 -953 0 net=1
rlabel metal2 1038 -953 1038 -953 0 net=8873
rlabel metal2 1150 -953 1150 -953 0 net=11525
rlabel metal2 464 -955 464 -955 0 net=4947
rlabel metal2 1052 -955 1052 -955 0 net=8899
rlabel metal2 1332 -955 1332 -955 0 net=11713
rlabel metal2 576 -957 576 -957 0 net=7679
rlabel metal2 765 -957 765 -957 0 net=5819
rlabel metal2 583 -959 583 -959 0 net=6191
rlabel metal2 842 -959 842 -959 0 net=11591
rlabel metal2 583 -961 583 -961 0 net=6422
rlabel metal2 1059 -961 1059 -961 0 net=9291
rlabel metal2 597 -963 597 -963 0 net=8283
rlabel metal2 1031 -963 1031 -963 0 net=8393
rlabel metal2 1094 -963 1094 -963 0 net=10197
rlabel metal2 639 -965 639 -965 0 net=6633
rlabel metal2 639 -967 639 -967 0 net=12001
rlabel metal2 646 -969 646 -969 0 net=6821
rlabel metal2 982 -969 982 -969 0 net=8185
rlabel metal2 1031 -969 1031 -969 0 net=8513
rlabel metal2 646 -971 646 -971 0 net=10060
rlabel metal2 716 -973 716 -973 0 net=7245
rlabel metal2 849 -973 849 -973 0 net=7393
rlabel metal2 978 -973 978 -973 0 net=10451
rlabel metal2 681 -975 681 -975 0 net=7561
rlabel metal2 982 -975 982 -975 0 net=9448
rlabel metal2 226 -977 226 -977 0 net=2625
rlabel metal2 709 -977 709 -977 0 net=5575
rlabel metal2 730 -977 730 -977 0 net=10289
rlabel metal2 499 -979 499 -979 0 net=4465
rlabel metal2 733 -979 733 -979 0 net=6691
rlabel metal2 1073 -979 1073 -979 0 net=8669
rlabel metal2 1199 -979 1199 -979 0 net=10243
rlabel metal2 737 -981 737 -981 0 net=8031
rlabel metal2 1045 -981 1045 -981 0 net=8967
rlabel metal2 996 -983 996 -983 0 net=12310
rlabel metal2 653 -985 653 -985 0 net=12581
rlabel metal2 1045 -987 1045 -987 0 net=9559
rlabel metal2 1080 -989 1080 -989 0 net=8819
rlabel metal2 1136 -989 1136 -989 0 net=9429
rlabel metal2 884 -991 884 -991 0 net=9177
rlabel metal2 1122 -991 1122 -991 0 net=9351
rlabel metal2 1066 -993 1066 -993 0 net=10133
rlabel metal2 537 -995 537 -995 0 net=9055
rlabel metal2 23 -1006 23 -1006 0 net=12103
rlabel metal2 628 -1006 628 -1006 0 net=6136
rlabel metal2 751 -1006 751 -1006 0 net=6193
rlabel metal2 751 -1006 751 -1006 0 net=6193
rlabel metal2 768 -1006 768 -1006 0 net=8390
rlabel metal2 961 -1006 961 -1006 0 net=11714
rlabel metal2 1339 -1006 1339 -1006 0 net=11073
rlabel metal2 1339 -1006 1339 -1006 0 net=11073
rlabel metal2 1374 -1006 1374 -1006 0 net=12088
rlabel metal2 1570 -1006 1570 -1006 0 net=12485
rlabel metal2 1738 -1006 1738 -1006 0 net=7753
rlabel metal2 30 -1008 30 -1008 0 net=7034
rlabel metal2 149 -1008 149 -1008 0 net=1793
rlabel metal2 250 -1008 250 -1008 0 net=4800
rlabel metal2 310 -1008 310 -1008 0 net=3394
rlabel metal2 555 -1008 555 -1008 0 net=6089
rlabel metal2 786 -1008 786 -1008 0 net=2666
rlabel metal2 919 -1008 919 -1008 0 net=7220
rlabel metal2 1528 -1008 1528 -1008 0 net=12529
rlabel metal2 1591 -1008 1591 -1008 0 net=5817
rlabel metal2 30 -1010 30 -1010 0 net=8285
rlabel metal2 611 -1010 611 -1010 0 net=4190
rlabel metal2 667 -1010 667 -1010 0 net=4702
rlabel metal2 786 -1010 786 -1010 0 net=6899
rlabel metal2 845 -1010 845 -1010 0 net=8968
rlabel metal2 1241 -1010 1241 -1010 0 net=11487
rlabel metal2 1486 -1010 1486 -1010 0 net=12363
rlabel metal2 1535 -1010 1535 -1010 0 net=12583
rlabel metal2 37 -1012 37 -1012 0 net=6956
rlabel metal2 698 -1012 698 -1012 0 net=12683
rlabel metal2 1626 -1012 1626 -1012 0 net=8003
rlabel metal2 44 -1014 44 -1014 0 net=6838
rlabel metal2 82 -1014 82 -1014 0 net=3054
rlabel metal2 114 -1014 114 -1014 0 net=4138
rlabel metal2 275 -1014 275 -1014 0 net=3164
rlabel metal2 1010 -1014 1010 -1014 0 net=12334
rlabel metal2 1552 -1014 1552 -1014 0 net=8926
rlabel metal2 1633 -1014 1633 -1014 0 net=11311
rlabel metal2 1633 -1014 1633 -1014 0 net=11311
rlabel metal2 44 -1016 44 -1016 0 net=5529
rlabel metal2 89 -1016 89 -1016 0 net=8202
rlabel metal2 422 -1016 422 -1016 0 net=2370
rlabel metal2 58 -1018 58 -1018 0 net=4513
rlabel metal2 72 -1018 72 -1018 0 net=3286
rlabel metal2 100 -1018 100 -1018 0 net=4156
rlabel metal2 485 -1018 485 -1018 0 net=5031
rlabel metal2 618 -1018 618 -1018 0 net=4261
rlabel metal2 684 -1018 684 -1018 0 net=9036
rlabel metal2 1241 -1018 1241 -1018 0 net=10597
rlabel metal2 1360 -1018 1360 -1018 0 net=11867
rlabel metal2 1500 -1018 1500 -1018 0 net=12449
rlabel metal2 1556 -1018 1556 -1018 0 net=12699
rlabel metal2 51 -1020 51 -1020 0 net=4656
rlabel metal2 100 -1020 100 -1020 0 net=4009
rlabel metal2 492 -1020 492 -1020 0 net=9022
rlabel metal2 800 -1020 800 -1020 0 net=10550
rlabel metal2 1269 -1020 1269 -1020 0 net=10331
rlabel metal2 1269 -1020 1269 -1020 0 net=10331
rlabel metal2 1297 -1020 1297 -1020 0 net=10813
rlabel metal2 1395 -1020 1395 -1020 0 net=11963
rlabel metal2 1563 -1020 1563 -1020 0 net=7167
rlabel metal2 51 -1022 51 -1022 0 net=9595
rlabel metal2 128 -1022 128 -1022 0 net=859
rlabel metal2 268 -1022 268 -1022 0 net=2677
rlabel metal2 492 -1022 492 -1022 0 net=3623
rlabel metal2 996 -1022 996 -1022 0 net=11584
rlabel metal2 1381 -1022 1381 -1022 0 net=11265
rlabel metal2 1423 -1022 1423 -1022 0 net=12239
rlabel metal2 1577 -1022 1577 -1022 0 net=4175
rlabel metal2 58 -1024 58 -1024 0 net=2365
rlabel metal2 107 -1024 107 -1024 0 net=8859
rlabel metal2 499 -1024 499 -1024 0 net=5090
rlabel metal2 632 -1024 632 -1024 0 net=5165
rlabel metal2 730 -1024 730 -1024 0 net=6234
rlabel metal2 835 -1024 835 -1024 0 net=6693
rlabel metal2 1003 -1024 1003 -1024 0 net=8187
rlabel metal2 1013 -1024 1013 -1024 0 net=8514
rlabel metal2 1108 -1024 1108 -1024 0 net=12495
rlabel metal2 1584 -1024 1584 -1024 0 net=11471
rlabel metal2 114 -1026 114 -1026 0 net=3669
rlabel metal2 275 -1026 275 -1026 0 net=6307
rlabel metal2 849 -1026 849 -1026 0 net=7395
rlabel metal2 849 -1026 849 -1026 0 net=7395
rlabel metal2 856 -1026 856 -1026 0 net=7777
rlabel metal2 933 -1026 933 -1026 0 net=7641
rlabel metal2 975 -1026 975 -1026 0 net=9057
rlabel metal2 1111 -1026 1111 -1026 0 net=12150
rlabel metal2 1507 -1026 1507 -1026 0 net=10819
rlabel metal2 121 -1028 121 -1028 0 net=2121
rlabel metal2 324 -1028 324 -1028 0 net=2902
rlabel metal2 520 -1028 520 -1028 0 net=3585
rlabel metal2 733 -1028 733 -1028 0 net=11363
rlabel metal2 1409 -1028 1409 -1028 0 net=11689
rlabel metal2 1430 -1028 1430 -1028 0 net=12003
rlabel metal2 1542 -1028 1542 -1028 0 net=12675
rlabel metal2 128 -1030 128 -1030 0 net=3539
rlabel metal2 282 -1030 282 -1030 0 net=2572
rlabel metal2 541 -1030 541 -1030 0 net=3821
rlabel metal2 688 -1030 688 -1030 0 net=6634
rlabel metal2 1220 -1030 1220 -1030 0 net=10664
rlabel metal2 1318 -1030 1318 -1030 0 net=11061
rlabel metal2 1409 -1030 1409 -1030 0 net=12051
rlabel metal2 1444 -1030 1444 -1030 0 net=10039
rlabel metal2 138 -1032 138 -1032 0 net=5741
rlabel metal2 506 -1032 506 -1032 0 net=11009
rlabel metal2 1416 -1032 1416 -1032 0 net=11785
rlabel metal2 1444 -1032 1444 -1032 0 net=12081
rlabel metal2 138 -1034 138 -1034 0 net=12140
rlabel metal2 156 -1036 156 -1036 0 net=1951
rlabel metal2 331 -1036 331 -1036 0 net=2216
rlabel metal2 541 -1036 541 -1036 0 net=4365
rlabel metal2 576 -1036 576 -1036 0 net=7680
rlabel metal2 737 -1036 737 -1036 0 net=8033
rlabel metal2 863 -1036 863 -1036 0 net=6822
rlabel metal2 891 -1036 891 -1036 0 net=7689
rlabel metal2 954 -1036 954 -1036 0 net=8141
rlabel metal2 1066 -1036 1066 -1036 0 net=9293
rlabel metal2 1115 -1036 1115 -1036 0 net=8323
rlabel metal2 1402 -1036 1402 -1036 0 net=11593
rlabel metal2 1472 -1036 1472 -1036 0 net=11004
rlabel metal2 156 -1038 156 -1038 0 net=4609
rlabel metal2 394 -1038 394 -1038 0 net=5341
rlabel metal2 548 -1038 548 -1038 0 net=3955
rlabel metal2 562 -1038 562 -1038 0 net=6253
rlabel metal2 660 -1038 660 -1038 0 net=6815
rlabel metal2 793 -1038 793 -1038 0 net=6889
rlabel metal2 866 -1038 866 -1038 0 net=11526
rlabel metal2 1157 -1038 1157 -1038 0 net=10737
rlabel metal2 1388 -1038 1388 -1038 0 net=11275
rlabel metal2 1598 -1038 1598 -1038 0 net=5821
rlabel metal2 170 -1040 170 -1040 0 net=2805
rlabel metal2 177 -1040 177 -1040 0 net=3205
rlabel metal2 296 -1040 296 -1040 0 net=6065
rlabel metal2 891 -1040 891 -1040 0 net=9553
rlabel metal2 1129 -1040 1129 -1040 0 net=8707
rlabel metal2 1157 -1040 1157 -1040 0 net=10859
rlabel metal2 1388 -1040 1388 -1040 0 net=11215
rlabel metal2 170 -1042 170 -1042 0 net=5387
rlabel metal2 310 -1042 310 -1042 0 net=1863
rlabel metal2 401 -1042 401 -1042 0 net=2013
rlabel metal2 457 -1042 457 -1042 0 net=5119
rlabel metal2 548 -1042 548 -1042 0 net=6235
rlabel metal2 691 -1042 691 -1042 0 net=2791
rlabel metal2 894 -1042 894 -1042 0 net=8820
rlabel metal2 1090 -1042 1090 -1042 0 net=11763
rlabel metal2 177 -1044 177 -1044 0 net=4339
rlabel metal2 219 -1044 219 -1044 0 net=7841
rlabel metal2 331 -1044 331 -1044 0 net=2509
rlabel metal2 457 -1044 457 -1044 0 net=3405
rlabel metal2 562 -1044 562 -1044 0 net=4309
rlabel metal2 184 -1046 184 -1046 0 net=1581
rlabel metal2 219 -1046 219 -1046 0 net=3765
rlabel metal2 569 -1046 569 -1046 0 net=5457
rlabel metal2 716 -1046 716 -1046 0 net=5577
rlabel metal2 870 -1046 870 -1046 0 net=8769
rlabel metal2 1129 -1046 1129 -1046 0 net=9785
rlabel metal2 1185 -1046 1185 -1046 0 net=9973
rlabel metal2 1234 -1046 1234 -1046 0 net=10303
rlabel metal2 1255 -1046 1255 -1046 0 net=10761
rlabel metal2 142 -1048 142 -1048 0 net=1739
rlabel metal2 191 -1048 191 -1048 0 net=2704
rlabel metal2 660 -1048 660 -1048 0 net=3973
rlabel metal2 821 -1048 821 -1048 0 net=7247
rlabel metal2 877 -1048 877 -1048 0 net=7727
rlabel metal2 142 -1050 142 -1050 0 net=3447
rlabel metal2 733 -1050 733 -1050 0 net=10611
rlabel metal2 191 -1052 191 -1052 0 net=4201
rlabel metal2 338 -1052 338 -1052 0 net=2481
rlabel metal2 394 -1052 394 -1052 0 net=11976
rlabel metal2 198 -1054 198 -1054 0 net=1543
rlabel metal2 345 -1054 345 -1054 0 net=1851
rlabel metal2 345 -1054 345 -1054 0 net=1851
rlabel metal2 352 -1054 352 -1054 0 net=3848
rlabel metal2 625 -1054 625 -1054 0 net=8823
rlabel metal2 744 -1054 744 -1054 0 net=6703
rlabel metal2 877 -1054 877 -1054 0 net=10259
rlabel metal2 1206 -1054 1206 -1054 0 net=8571
rlabel metal2 163 -1056 163 -1056 0 net=1783
rlabel metal2 254 -1056 254 -1056 0 net=3639
rlabel metal2 446 -1056 446 -1056 0 net=908
rlabel metal2 744 -1056 744 -1056 0 net=6791
rlabel metal2 912 -1056 912 -1056 0 net=7563
rlabel metal2 163 -1058 163 -1058 0 net=6443
rlabel metal2 401 -1058 401 -1058 0 net=6485
rlabel metal2 597 -1058 597 -1058 0 net=4145
rlabel metal2 1073 -1058 1073 -1058 0 net=8671
rlabel metal2 1227 -1058 1227 -1058 0 net=10291
rlabel metal2 1353 -1058 1353 -1058 0 net=11239
rlabel metal2 1465 -1058 1465 -1058 0 net=12479
rlabel metal2 261 -1060 261 -1060 0 net=2293
rlabel metal2 359 -1060 359 -1060 0 net=3043
rlabel metal2 450 -1060 450 -1060 0 net=3941
rlabel metal2 653 -1060 653 -1060 0 net=11081
rlabel metal2 926 -1060 926 -1060 0 net=7525
rlabel metal2 982 -1060 982 -1060 0 net=9473
rlabel metal2 1213 -1060 1213 -1060 0 net=10245
rlabel metal2 1346 -1060 1346 -1060 0 net=11189
rlabel metal2 1465 -1060 1465 -1060 0 net=12325
rlabel metal2 359 -1062 359 -1062 0 net=2487
rlabel metal2 905 -1062 905 -1062 0 net=7161
rlabel metal2 985 -1062 985 -1062 0 net=12236
rlabel metal2 366 -1064 366 -1064 0 net=3503
rlabel metal2 366 -1064 366 -1064 0 net=3503
rlabel metal2 373 -1064 373 -1064 0 net=3099
rlabel metal2 464 -1064 464 -1064 0 net=4949
rlabel metal2 649 -1064 649 -1064 0 net=7425
rlabel metal2 933 -1064 933 -1064 0 net=8461
rlabel metal2 1024 -1064 1024 -1064 0 net=8483
rlabel metal2 1073 -1064 1073 -1064 0 net=9353
rlabel metal2 1171 -1064 1171 -1064 0 net=10181
rlabel metal2 1458 -1064 1458 -1064 0 net=12093
rlabel metal2 226 -1066 226 -1066 0 net=2627
rlabel metal2 380 -1066 380 -1066 0 net=4087
rlabel metal2 471 -1066 471 -1066 0 net=7403
rlabel metal2 968 -1066 968 -1066 0 net=7955
rlabel metal2 1024 -1066 1024 -1066 0 net=8875
rlabel metal2 1136 -1066 1136 -1066 0 net=9691
rlabel metal2 226 -1068 226 -1068 0 net=2663
rlabel metal2 429 -1068 429 -1068 0 net=3267
rlabel metal2 534 -1068 534 -1068 0 net=3359
rlabel metal2 863 -1068 863 -1068 0 net=11847
rlabel metal2 289 -1070 289 -1070 0 net=3071
rlabel metal2 576 -1070 576 -1070 0 net=5363
rlabel metal2 289 -1072 289 -1072 0 net=2781
rlabel metal2 583 -1072 583 -1072 0 net=7207
rlabel metal2 905 -1072 905 -1072 0 net=7221
rlabel metal2 1122 -1072 1122 -1072 0 net=10135
rlabel metal2 250 -1074 250 -1074 0 net=4031
rlabel metal2 586 -1074 586 -1074 0 net=7169
rlabel metal2 947 -1074 947 -1074 0 net=8097
rlabel metal2 989 -1074 989 -1074 0 net=10790
rlabel metal2 303 -1076 303 -1076 0 net=4015
rlabel metal2 947 -1076 947 -1076 0 net=8901
rlabel metal2 1132 -1076 1132 -1076 0 net=1
rlabel metal2 1171 -1076 1171 -1076 0 net=9933
rlabel metal2 1262 -1076 1262 -1076 0 net=10585
rlabel metal2 131 -1078 131 -1078 0 net=4431
rlabel metal2 1045 -1078 1045 -1078 0 net=9561
rlabel metal2 1143 -1078 1143 -1078 0 net=9431
rlabel metal2 1283 -1078 1283 -1078 0 net=10557
rlabel metal2 338 -1080 338 -1080 0 net=11443
rlabel metal2 1045 -1080 1045 -1080 0 net=8394
rlabel metal2 1094 -1080 1094 -1080 0 net=10199
rlabel metal2 1276 -1080 1276 -1080 0 net=10453
rlabel metal2 513 -1082 513 -1082 0 net=4705
rlabel metal2 642 -1082 642 -1082 0 net=11829
rlabel metal2 513 -1084 513 -1084 0 net=486
rlabel metal2 828 -1084 828 -1084 0 net=9363
rlabel metal2 79 -1086 79 -1086 0 net=5757
rlabel metal2 814 -1086 814 -1086 0 net=6115
rlabel metal2 978 -1086 978 -1086 0 net=8263
rlabel metal2 79 -1088 79 -1088 0 net=3829
rlabel metal2 653 -1088 653 -1088 0 net=4467
rlabel metal2 807 -1088 807 -1088 0 net=7201
rlabel metal2 1006 -1088 1006 -1088 0 net=10387
rlabel metal2 93 -1090 93 -1090 0 net=4029
rlabel metal2 674 -1090 674 -1090 0 net=12301
rlabel metal2 499 -1092 499 -1092 0 net=9927
rlabel metal2 709 -1092 709 -1092 0 net=5473
rlabel metal2 807 -1094 807 -1094 0 net=3967
rlabel metal2 898 -1094 898 -1094 0 net=9179
rlabel metal2 1087 -1096 1087 -1096 0 net=9221
rlabel metal2 23 -1107 23 -1107 0 net=12104
rlabel metal2 471 -1107 471 -1107 0 net=3586
rlabel metal2 730 -1107 730 -1107 0 net=10598
rlabel metal2 1255 -1107 1255 -1107 0 net=10762
rlabel metal2 1384 -1107 1384 -1107 0 net=4176
rlabel metal2 1640 -1107 1640 -1107 0 net=12585
rlabel metal2 1745 -1107 1745 -1107 0 net=7755
rlabel metal2 23 -1109 23 -1109 0 net=3871
rlabel metal2 275 -1109 275 -1109 0 net=6309
rlabel metal2 499 -1109 499 -1109 0 net=9928
rlabel metal2 649 -1109 649 -1109 0 net=6792
rlabel metal2 765 -1109 765 -1109 0 net=4432
rlabel metal2 887 -1109 887 -1109 0 net=11488
rlabel metal2 1423 -1109 1423 -1109 0 net=11691
rlabel metal2 1423 -1109 1423 -1109 0 net=11691
rlabel metal2 1444 -1109 1444 -1109 0 net=12083
rlabel metal2 1675 -1109 1675 -1109 0 net=12487
rlabel metal2 37 -1111 37 -1111 0 net=5461
rlabel metal2 219 -1111 219 -1111 0 net=3766
rlabel metal2 275 -1111 275 -1111 0 net=4017
rlabel metal2 324 -1111 324 -1111 0 net=1544
rlabel metal2 366 -1111 366 -1111 0 net=3505
rlabel metal2 366 -1111 366 -1111 0 net=3505
rlabel metal2 401 -1111 401 -1111 0 net=6486
rlabel metal2 681 -1111 681 -1111 0 net=5759
rlabel metal2 817 -1111 817 -1111 0 net=9974
rlabel metal2 1213 -1111 1213 -1111 0 net=10183
rlabel metal2 1444 -1111 1444 -1111 0 net=10977
rlabel metal2 72 -1113 72 -1113 0 net=4367
rlabel metal2 656 -1113 656 -1113 0 net=12302
rlabel metal2 1451 -1113 1451 -1113 0 net=10040
rlabel metal2 1570 -1113 1570 -1113 0 net=12531
rlabel metal2 75 -1115 75 -1115 0 net=12115
rlabel metal2 1682 -1115 1682 -1115 0 net=5818
rlabel metal2 89 -1117 89 -1117 0 net=5765
rlabel metal2 516 -1117 516 -1117 0 net=4146
rlabel metal2 681 -1117 681 -1117 0 net=2793
rlabel metal2 835 -1117 835 -1117 0 net=6890
rlabel metal2 929 -1117 929 -1117 0 net=10814
rlabel metal2 1318 -1117 1318 -1117 0 net=11011
rlabel metal2 1465 -1117 1465 -1117 0 net=12327
rlabel metal2 93 -1119 93 -1119 0 net=4030
rlabel metal2 548 -1119 548 -1119 0 net=6237
rlabel metal2 933 -1119 933 -1119 0 net=8463
rlabel metal2 1437 -1119 1437 -1119 0 net=11787
rlabel metal2 1570 -1119 1570 -1119 0 net=11473
rlabel metal2 1612 -1119 1612 -1119 0 net=12701
rlabel metal2 93 -1121 93 -1121 0 net=1725
rlabel metal2 173 -1121 173 -1121 0 net=3822
rlabel metal2 688 -1121 688 -1121 0 net=945
rlabel metal2 859 -1121 859 -1121 0 net=9180
rlabel metal2 912 -1121 912 -1121 0 net=7405
rlabel metal2 950 -1121 950 -1121 0 net=7728
rlabel metal2 1311 -1121 1311 -1121 0 net=10739
rlabel metal2 1479 -1121 1479 -1121 0 net=11849
rlabel metal2 1654 -1121 1654 -1121 0 net=8005
rlabel metal2 100 -1123 100 -1123 0 net=4011
rlabel metal2 506 -1123 506 -1123 0 net=5121
rlabel metal2 737 -1123 737 -1123 0 net=5579
rlabel metal2 758 -1123 758 -1123 0 net=6817
rlabel metal2 1045 -1123 1045 -1123 0 net=10292
rlabel metal2 1248 -1123 1248 -1123 0 net=10305
rlabel metal2 58 -1125 58 -1125 0 net=2367
rlabel metal2 107 -1125 107 -1125 0 net=8860
rlabel metal2 236 -1125 236 -1125 0 net=11183
rlabel metal2 1493 -1125 1493 -1125 0 net=5822
rlabel metal2 58 -1127 58 -1127 0 net=5389
rlabel metal2 177 -1127 177 -1127 0 net=4341
rlabel metal2 653 -1127 653 -1127 0 net=4469
rlabel metal2 891 -1127 891 -1127 0 net=9533
rlabel metal2 1332 -1127 1332 -1127 0 net=8324
rlabel metal2 1496 -1127 1496 -1127 0 net=7168
rlabel metal2 68 -1129 68 -1129 0 net=9241
rlabel metal2 1290 -1129 1290 -1129 0 net=10559
rlabel metal2 89 -1131 89 -1131 0 net=8759
rlabel metal2 1500 -1131 1500 -1131 0 net=11965
rlabel metal2 110 -1133 110 -1133 0 net=5249
rlabel metal2 380 -1133 380 -1133 0 net=4089
rlabel metal2 698 -1133 698 -1133 0 net=6900
rlabel metal2 891 -1133 891 -1133 0 net=9515
rlabel metal2 1325 -1133 1325 -1133 0 net=11063
rlabel metal2 1507 -1133 1507 -1133 0 net=12005
rlabel metal2 114 -1135 114 -1135 0 net=3671
rlabel metal2 114 -1135 114 -1135 0 net=3671
rlabel metal2 121 -1135 121 -1135 0 net=2122
rlabel metal2 401 -1135 401 -1135 0 net=2679
rlabel metal2 415 -1135 415 -1135 0 net=3044
rlabel metal2 716 -1135 716 -1135 0 net=8825
rlabel metal2 1220 -1135 1220 -1135 0 net=12513
rlabel metal2 121 -1137 121 -1137 0 net=11857
rlabel metal2 128 -1139 128 -1139 0 net=3541
rlabel metal2 180 -1139 180 -1139 0 net=1864
rlabel metal2 380 -1139 380 -1139 0 net=5459
rlabel metal2 649 -1139 649 -1139 0 net=9117
rlabel metal2 1325 -1139 1325 -1139 0 net=11765
rlabel metal2 1514 -1139 1514 -1139 0 net=12095
rlabel metal2 128 -1141 128 -1141 0 net=1599
rlabel metal2 233 -1141 233 -1141 0 net=3269
rlabel metal2 485 -1141 485 -1141 0 net=5743
rlabel metal2 919 -1141 919 -1141 0 net=7779
rlabel metal2 1048 -1141 1048 -1141 0 net=10260
rlabel metal2 1339 -1141 1339 -1141 0 net=11075
rlabel metal2 1528 -1141 1528 -1141 0 net=12365
rlabel metal2 184 -1143 184 -1143 0 net=1741
rlabel metal2 387 -1143 387 -1143 0 net=2483
rlabel metal2 415 -1143 415 -1143 0 net=3943
rlabel metal2 492 -1143 492 -1143 0 net=3625
rlabel metal2 723 -1143 723 -1143 0 net=6091
rlabel metal2 968 -1143 968 -1143 0 net=8099
rlabel metal2 1367 -1143 1367 -1143 0 net=11191
rlabel metal2 1549 -1143 1549 -1143 0 net=12481
rlabel metal2 79 -1145 79 -1145 0 net=3831
rlabel metal2 443 -1145 443 -1145 0 net=3101
rlabel metal2 499 -1145 499 -1145 0 net=4965
rlabel metal2 758 -1145 758 -1145 0 net=5237
rlabel metal2 1055 -1145 1055 -1145 0 net=11240
rlabel metal2 1402 -1145 1402 -1145 0 net=11277
rlabel metal2 1556 -1145 1556 -1145 0 net=12497
rlabel metal2 51 -1147 51 -1147 0 net=9597
rlabel metal2 1409 -1147 1409 -1147 0 net=12053
rlabel metal2 51 -1149 51 -1149 0 net=6679
rlabel metal2 611 -1149 611 -1149 0 net=5033
rlabel metal2 765 -1149 765 -1149 0 net=6755
rlabel metal2 1055 -1149 1055 -1149 0 net=8597
rlabel metal2 1269 -1149 1269 -1149 0 net=10333
rlabel metal2 1416 -1149 1416 -1149 0 net=11595
rlabel metal2 1577 -1149 1577 -1149 0 net=12677
rlabel metal2 65 -1151 65 -1151 0 net=4515
rlabel metal2 124 -1151 124 -1151 0 net=7139
rlabel metal2 1066 -1151 1066 -1151 0 net=9295
rlabel metal2 1276 -1151 1276 -1151 0 net=10389
rlabel metal2 1416 -1151 1416 -1151 0 net=10469
rlabel metal2 65 -1153 65 -1153 0 net=11043
rlabel metal2 1535 -1153 1535 -1153 0 net=12451
rlabel metal2 1577 -1153 1577 -1153 0 net=11313
rlabel metal2 142 -1155 142 -1155 0 net=3449
rlabel metal2 520 -1155 520 -1155 0 net=5343
rlabel metal2 768 -1155 768 -1155 0 net=8034
rlabel metal2 905 -1155 905 -1155 0 net=7223
rlabel metal2 1283 -1155 1283 -1155 0 net=10455
rlabel metal2 1486 -1155 1486 -1155 0 net=11869
rlabel metal2 184 -1157 184 -1157 0 net=4707
rlabel metal2 779 -1157 779 -1157 0 net=11083
rlabel metal2 1598 -1157 1598 -1157 0 net=10613
rlabel metal2 191 -1159 191 -1159 0 net=4203
rlabel metal2 191 -1159 191 -1159 0 net=4203
rlabel metal2 198 -1159 198 -1159 0 net=1785
rlabel metal2 338 -1159 338 -1159 0 net=6159
rlabel metal2 880 -1159 880 -1159 0 net=9417
rlabel metal2 1388 -1159 1388 -1159 0 net=11217
rlabel metal2 198 -1161 198 -1161 0 net=3641
rlabel metal2 282 -1161 282 -1161 0 net=7842
rlabel metal2 793 -1161 793 -1161 0 net=7171
rlabel metal2 1003 -1161 1003 -1161 0 net=9307
rlabel metal2 1458 -1161 1458 -1161 0 net=11831
rlabel metal2 177 -1163 177 -1163 0 net=2591
rlabel metal2 261 -1163 261 -1163 0 net=7555
rlabel metal2 1052 -1163 1052 -1163 0 net=11561
rlabel metal2 212 -1165 212 -1165 0 net=1545
rlabel metal2 821 -1165 821 -1165 0 net=6705
rlabel metal2 1066 -1165 1066 -1165 0 net=7565
rlabel metal2 219 -1167 219 -1167 0 net=2751
rlabel metal2 282 -1167 282 -1167 0 net=3573
rlabel metal2 443 -1167 443 -1167 0 net=5199
rlabel metal2 793 -1167 793 -1167 0 net=9354
rlabel metal2 1087 -1167 1087 -1167 0 net=9786
rlabel metal2 1143 -1167 1143 -1167 0 net=10201
rlabel metal2 1458 -1167 1458 -1167 0 net=12685
rlabel metal2 226 -1169 226 -1169 0 net=2664
rlabel metal2 688 -1169 688 -1169 0 net=4671
rlabel metal2 961 -1169 961 -1169 0 net=7643
rlabel metal2 1094 -1169 1094 -1169 0 net=9365
rlabel metal2 1521 -1169 1521 -1169 0 net=12241
rlabel metal2 1584 -1169 1584 -1169 0 net=10821
rlabel metal2 30 -1171 30 -1171 0 net=8286
rlabel metal2 247 -1171 247 -1171 0 net=3417
rlabel metal2 520 -1171 520 -1171 0 net=3663
rlabel metal2 996 -1171 996 -1171 0 net=6695
rlabel metal2 1101 -1171 1101 -1171 0 net=8673
rlabel metal2 1395 -1171 1395 -1171 0 net=11267
rlabel metal2 30 -1173 30 -1173 0 net=5677
rlabel metal2 205 -1173 205 -1173 0 net=1583
rlabel metal2 296 -1173 296 -1173 0 net=6067
rlabel metal2 471 -1173 471 -1173 0 net=3173
rlabel metal2 1010 -1173 1010 -1173 0 net=8189
rlabel metal2 1150 -1173 1150 -1173 0 net=9223
rlabel metal2 86 -1175 86 -1175 0 net=6444
rlabel metal2 205 -1175 205 -1175 0 net=3407
rlabel metal2 527 -1175 527 -1175 0 net=4033
rlabel metal2 618 -1175 618 -1175 0 net=4263
rlabel metal2 695 -1175 695 -1175 0 net=11364
rlabel metal2 149 -1177 149 -1177 0 net=1795
rlabel metal2 289 -1177 289 -1177 0 net=2783
rlabel metal2 338 -1177 338 -1177 0 net=2015
rlabel metal2 457 -1177 457 -1177 0 net=3361
rlabel metal2 569 -1177 569 -1177 0 net=5475
rlabel metal2 828 -1177 828 -1177 0 net=6117
rlabel metal2 982 -1177 982 -1177 0 net=7163
rlabel metal2 1017 -1177 1017 -1177 0 net=7957
rlabel metal2 1101 -1177 1101 -1177 0 net=9693
rlabel metal2 1157 -1177 1157 -1177 0 net=10861
rlabel metal2 1360 -1177 1360 -1177 0 net=10165
rlabel metal2 145 -1179 145 -1179 0 net=3559
rlabel metal2 170 -1179 170 -1179 0 net=8137
rlabel metal2 1164 -1179 1164 -1179 0 net=8709
rlabel metal2 268 -1181 268 -1181 0 net=3206
rlabel metal2 464 -1181 464 -1181 0 net=3073
rlabel metal2 562 -1181 562 -1181 0 net=4311
rlabel metal2 740 -1181 740 -1181 0 net=8359
rlabel metal2 1171 -1181 1171 -1181 0 net=9935
rlabel metal2 142 -1183 142 -1183 0 net=3045
rlabel metal2 331 -1183 331 -1183 0 net=2511
rlabel metal2 562 -1183 562 -1183 0 net=961
rlabel metal2 849 -1183 849 -1183 0 net=7397
rlabel metal2 1038 -1183 1038 -1183 0 net=8485
rlabel metal2 1178 -1183 1178 -1183 0 net=10137
rlabel metal2 331 -1185 331 -1185 0 net=2489
rlabel metal2 576 -1185 576 -1185 0 net=5365
rlabel metal2 856 -1185 856 -1185 0 net=7209
rlabel metal2 1059 -1185 1059 -1185 0 net=8265
rlabel metal2 1178 -1185 1178 -1185 0 net=8573
rlabel metal2 1227 -1185 1227 -1185 0 net=10247
rlabel metal2 345 -1187 345 -1187 0 net=1853
rlabel metal2 555 -1187 555 -1187 0 net=3957
rlabel metal2 583 -1187 583 -1187 0 net=6137
rlabel metal2 751 -1187 751 -1187 0 net=6195
rlabel metal2 856 -1187 856 -1187 0 net=7307
rlabel metal2 1080 -1187 1080 -1187 0 net=8771
rlabel metal2 1227 -1187 1227 -1187 0 net=10587
rlabel metal2 345 -1189 345 -1189 0 net=2267
rlabel metal2 555 -1189 555 -1189 0 net=5167
rlabel metal2 674 -1189 674 -1189 0 net=3969
rlabel metal2 926 -1189 926 -1189 0 net=7427
rlabel metal2 1108 -1189 1108 -1189 0 net=9475
rlabel metal2 1192 -1189 1192 -1189 0 net=9433
rlabel metal2 394 -1191 394 -1191 0 net=7853
rlabel metal2 1115 -1191 1115 -1191 0 net=9555
rlabel metal2 352 -1193 352 -1193 0 net=2295
rlabel metal2 618 -1193 618 -1193 0 net=4439
rlabel metal2 898 -1193 898 -1193 0 net=6447
rlabel metal2 940 -1193 940 -1193 0 net=7691
rlabel metal2 1122 -1193 1122 -1193 0 net=9563
rlabel metal2 352 -1195 352 -1195 0 net=2629
rlabel metal2 691 -1195 691 -1195 0 net=7887
rlabel metal2 1262 -1195 1262 -1195 0 net=5471
rlabel metal2 317 -1197 317 -1197 0 net=1953
rlabel metal2 702 -1197 702 -1197 0 net=7901
rlabel metal2 44 -1199 44 -1199 0 net=5531
rlabel metal2 751 -1199 751 -1199 0 net=5231
rlabel metal2 947 -1199 947 -1199 0 net=8903
rlabel metal2 44 -1201 44 -1201 0 net=4611
rlabel metal2 541 -1201 541 -1201 0 net=9037
rlabel metal2 947 -1201 947 -1201 0 net=8876
rlabel metal2 1031 -1201 1031 -1201 0 net=8143
rlabel metal2 156 -1203 156 -1203 0 net=4951
rlabel metal2 796 -1203 796 -1203 0 net=5847
rlabel metal2 954 -1203 954 -1203 0 net=7527
rlabel metal2 590 -1205 590 -1205 0 net=3975
rlabel metal2 698 -1205 698 -1205 0 net=6931
rlabel metal2 975 -1205 975 -1205 0 net=9059
rlabel metal2 604 -1207 604 -1207 0 net=6255
rlabel metal2 814 -1207 814 -1207 0 net=7203
rlabel metal2 989 -1207 989 -1207 0 net=11445
rlabel metal2 527 -1209 527 -1209 0 net=4991
rlabel metal2 814 -1209 814 -1209 0 net=6839
rlabel metal2 870 -1211 870 -1211 0 net=7249
rlabel metal2 240 -1213 240 -1213 0 net=2807
rlabel metal2 240 -1215 240 -1215 0 net=1717
rlabel metal2 16 -1226 16 -1226 0 net=2545
rlabel metal2 471 -1226 471 -1226 0 net=3175
rlabel metal2 471 -1226 471 -1226 0 net=3175
rlabel metal2 506 -1226 506 -1226 0 net=9038
rlabel metal2 891 -1226 891 -1226 0 net=7958
rlabel metal2 1094 -1226 1094 -1226 0 net=6696
rlabel metal2 1276 -1226 1276 -1226 0 net=9309
rlabel metal2 1276 -1226 1276 -1226 0 net=9309
rlabel metal2 1283 -1226 1283 -1226 0 net=9419
rlabel metal2 1283 -1226 1283 -1226 0 net=9419
rlabel metal2 1290 -1226 1290 -1226 0 net=9517
rlabel metal2 1311 -1226 1311 -1226 0 net=9535
rlabel metal2 1451 -1226 1451 -1226 0 net=11013
rlabel metal2 1451 -1226 1451 -1226 0 net=11013
rlabel metal2 1661 -1226 1661 -1226 0 net=12085
rlabel metal2 1661 -1226 1661 -1226 0 net=12085
rlabel metal2 1703 -1226 1703 -1226 0 net=12488
rlabel metal2 1766 -1226 1766 -1226 0 net=10614
rlabel metal2 44 -1228 44 -1228 0 net=4612
rlabel metal2 289 -1228 289 -1228 0 net=1718
rlabel metal2 548 -1228 548 -1228 0 net=4090
rlabel metal2 590 -1228 590 -1228 0 net=3976
rlabel metal2 607 -1228 607 -1228 0 net=7224
rlabel metal2 1290 -1228 1290 -1228 0 net=9565
rlabel metal2 1311 -1228 1311 -1228 0 net=9937
rlabel metal2 1696 -1228 1696 -1228 0 net=12483
rlabel metal2 1745 -1228 1745 -1228 0 net=7756
rlabel metal2 44 -1230 44 -1230 0 net=3331
rlabel metal2 93 -1230 93 -1230 0 net=1727
rlabel metal2 93 -1230 93 -1230 0 net=1727
rlabel metal2 103 -1230 103 -1230 0 net=1742
rlabel metal2 345 -1230 345 -1230 0 net=2268
rlabel metal2 800 -1230 800 -1230 0 net=5761
rlabel metal2 894 -1230 894 -1230 0 net=10306
rlabel metal2 1745 -1230 1745 -1230 0 net=11109
rlabel metal2 65 -1232 65 -1232 0 net=9598
rlabel metal2 1612 -1232 1612 -1232 0 net=12533
rlabel metal2 54 -1234 54 -1234 0 net=1983
rlabel metal2 68 -1234 68 -1234 0 net=4516
rlabel metal2 107 -1234 107 -1234 0 net=3672
rlabel metal2 121 -1234 121 -1234 0 net=8464
rlabel metal2 1717 -1234 1717 -1234 0 net=12679
rlabel metal2 72 -1236 72 -1236 0 net=4369
rlabel metal2 709 -1236 709 -1236 0 net=4312
rlabel metal2 817 -1236 817 -1236 0 net=6118
rlabel metal2 1010 -1236 1010 -1236 0 net=7165
rlabel metal2 1146 -1236 1146 -1236 0 net=8710
rlabel metal2 51 -1238 51 -1238 0 net=6681
rlabel metal2 110 -1238 110 -1238 0 net=6256
rlabel metal2 667 -1238 667 -1238 0 net=5345
rlabel metal2 821 -1238 821 -1238 0 net=10560
rlabel metal2 114 -1240 114 -1240 0 net=6841
rlabel metal2 947 -1240 947 -1240 0 net=11218
rlabel metal2 121 -1242 121 -1242 0 net=6453
rlabel metal2 551 -1242 551 -1242 0 net=8138
rlabel metal2 1178 -1242 1178 -1242 0 net=8575
rlabel metal2 1178 -1242 1178 -1242 0 net=8575
rlabel metal2 1248 -1242 1248 -1242 0 net=9243
rlabel metal2 1314 -1242 1314 -1242 0 net=1
rlabel metal2 1353 -1242 1353 -1242 0 net=11045
rlabel metal2 1486 -1242 1486 -1242 0 net=11563
rlabel metal2 124 -1244 124 -1244 0 net=6310
rlabel metal2 565 -1244 565 -1244 0 net=3626
rlabel metal2 737 -1244 737 -1244 0 net=5580
rlabel metal2 751 -1244 751 -1244 0 net=5233
rlabel metal2 779 -1244 779 -1244 0 net=5367
rlabel metal2 821 -1244 821 -1244 0 net=12242
rlabel metal2 61 -1246 61 -1246 0 net=872
rlabel metal2 740 -1246 740 -1246 0 net=8100
rlabel metal2 1360 -1246 1360 -1246 0 net=10167
rlabel metal2 1458 -1246 1458 -1246 0 net=12687
rlabel metal2 145 -1248 145 -1248 0 net=12452
rlabel metal2 170 -1250 170 -1250 0 net=182
rlabel metal2 180 -1250 180 -1250 0 net=12498
rlabel metal2 142 -1252 142 -1252 0 net=5287
rlabel metal2 177 -1252 177 -1252 0 net=3643
rlabel metal2 208 -1252 208 -1252 0 net=4167
rlabel metal2 243 -1252 243 -1252 0 net=8904
rlabel metal2 1220 -1252 1220 -1252 0 net=9119
rlabel metal2 1325 -1252 1325 -1252 0 net=11767
rlabel metal2 142 -1254 142 -1254 0 net=1547
rlabel metal2 226 -1254 226 -1254 0 net=7556
rlabel metal2 1010 -1254 1010 -1254 0 net=7781
rlabel metal2 1052 -1254 1052 -1254 0 net=9434
rlabel metal2 128 -1256 128 -1256 0 net=1601
rlabel metal2 226 -1256 226 -1256 0 net=2593
rlabel metal2 261 -1256 261 -1256 0 net=2167
rlabel metal2 443 -1256 443 -1256 0 net=5200
rlabel metal2 1059 -1256 1059 -1256 0 net=7429
rlabel metal2 1171 -1256 1171 -1256 0 net=8487
rlabel metal2 1325 -1256 1325 -1256 0 net=9571
rlabel metal2 163 -1258 163 -1258 0 net=1797
rlabel metal2 292 -1258 292 -1258 0 net=2808
rlabel metal2 933 -1258 933 -1258 0 net=7407
rlabel metal2 1087 -1258 1087 -1258 0 net=11065
rlabel metal2 1542 -1258 1542 -1258 0 net=11597
rlabel metal2 1584 -1258 1584 -1258 0 net=10823
rlabel metal2 163 -1260 163 -1260 0 net=3349
rlabel metal2 723 -1260 723 -1260 0 net=5035
rlabel metal2 751 -1260 751 -1260 0 net=937
rlabel metal2 824 -1260 824 -1260 0 net=578
rlabel metal2 1101 -1260 1101 -1260 0 net=9695
rlabel metal2 1402 -1260 1402 -1260 0 net=10391
rlabel metal2 1465 -1260 1465 -1260 0 net=11077
rlabel metal2 1549 -1260 1549 -1260 0 net=11833
rlabel metal2 184 -1262 184 -1262 0 net=4709
rlabel metal2 740 -1262 740 -1262 0 net=11084
rlabel metal2 1479 -1262 1479 -1262 0 net=11967
rlabel metal2 184 -1264 184 -1264 0 net=4440
rlabel metal2 632 -1264 632 -1264 0 net=9366
rlabel metal2 1402 -1264 1402 -1264 0 net=10979
rlabel metal2 1486 -1264 1486 -1264 0 net=11279
rlabel metal2 1570 -1264 1570 -1264 0 net=11475
rlabel metal2 1598 -1264 1598 -1264 0 net=11871
rlabel metal2 1640 -1264 1640 -1264 0 net=12055
rlabel metal2 198 -1266 198 -1266 0 net=7937
rlabel metal2 828 -1266 828 -1266 0 net=10073
rlabel metal2 1423 -1266 1423 -1266 0 net=11693
rlabel metal2 1528 -1266 1528 -1266 0 net=11315
rlabel metal2 1633 -1266 1633 -1266 0 net=12007
rlabel metal2 1654 -1266 1654 -1266 0 net=12117
rlabel metal2 296 -1268 296 -1268 0 net=2784
rlabel metal2 611 -1268 611 -1268 0 net=4035
rlabel metal2 639 -1268 639 -1268 0 net=4265
rlabel metal2 831 -1268 831 -1268 0 net=9296
rlabel metal2 1339 -1268 1339 -1268 0 net=10139
rlabel metal2 1423 -1268 1423 -1268 0 net=11193
rlabel metal2 1577 -1268 1577 -1268 0 net=11859
rlabel metal2 1647 -1268 1647 -1268 0 net=12097
rlabel metal2 1675 -1268 1675 -1268 0 net=12367
rlabel metal2 58 -1270 58 -1270 0 net=5391
rlabel metal2 611 -1270 611 -1270 0 net=6819
rlabel metal2 922 -1270 922 -1270 0 net=11863
rlabel metal2 1682 -1270 1682 -1270 0 net=12329
rlabel metal2 58 -1272 58 -1272 0 net=2368
rlabel metal2 296 -1272 296 -1272 0 net=2631
rlabel metal2 380 -1272 380 -1272 0 net=5460
rlabel metal2 702 -1272 702 -1272 0 net=10031
rlabel metal2 1500 -1272 1500 -1272 0 net=11269
rlabel metal2 1682 -1272 1682 -1272 0 net=12515
rlabel metal2 205 -1274 205 -1274 0 net=3409
rlabel metal2 380 -1274 380 -1274 0 net=3215
rlabel metal2 600 -1274 600 -1274 0 net=4147
rlabel metal2 688 -1274 688 -1274 0 net=4673
rlabel metal2 831 -1274 831 -1274 0 net=5472
rlabel metal2 1710 -1274 1710 -1274 0 net=12587
rlabel metal2 23 -1276 23 -1276 0 net=3872
rlabel metal2 303 -1276 303 -1276 0 net=2491
rlabel metal2 345 -1276 345 -1276 0 net=1955
rlabel metal2 387 -1276 387 -1276 0 net=3833
rlabel metal2 681 -1276 681 -1276 0 net=2795
rlabel metal2 835 -1276 835 -1276 0 net=6093
rlabel metal2 912 -1276 912 -1276 0 net=7211
rlabel metal2 996 -1276 996 -1276 0 net=7309
rlabel metal2 1101 -1276 1101 -1276 0 net=11184
rlabel metal2 1724 -1276 1724 -1276 0 net=12703
rlabel metal2 23 -1278 23 -1278 0 net=2825
rlabel metal2 548 -1278 548 -1278 0 net=9173
rlabel metal2 1752 -1278 1752 -1278 0 net=8007
rlabel metal2 310 -1280 310 -1280 0 net=1787
rlabel metal2 852 -1280 852 -1280 0 net=7172
rlabel metal2 929 -1280 929 -1280 0 net=12215
rlabel metal2 156 -1282 156 -1282 0 net=4953
rlabel metal2 317 -1282 317 -1282 0 net=5533
rlabel metal2 415 -1282 415 -1282 0 net=3945
rlabel metal2 513 -1282 513 -1282 0 net=5767
rlabel metal2 933 -1282 933 -1282 0 net=12609
rlabel metal2 149 -1284 149 -1284 0 net=3561
rlabel metal2 317 -1284 317 -1284 0 net=4981
rlabel metal2 856 -1284 856 -1284 0 net=8760
rlabel metal2 100 -1286 100 -1286 0 net=11283
rlabel metal2 149 -1288 149 -1288 0 net=6239
rlabel metal2 936 -1288 936 -1288 0 net=9556
rlabel metal2 331 -1290 331 -1290 0 net=1855
rlabel metal2 366 -1290 366 -1290 0 net=3507
rlabel metal2 625 -1290 625 -1290 0 net=4343
rlabel metal2 807 -1290 807 -1290 0 net=5849
rlabel metal2 940 -1290 940 -1290 0 net=6493
rlabel metal2 1017 -1290 1017 -1290 0 net=7399
rlabel metal2 1104 -1290 1104 -1290 0 net=11987
rlabel metal2 275 -1292 275 -1292 0 net=4019
rlabel metal2 667 -1292 667 -1292 0 net=4285
rlabel metal2 1038 -1292 1038 -1292 0 net=7693
rlabel metal2 135 -1294 135 -1294 0 net=3543
rlabel metal2 282 -1294 282 -1294 0 net=3575
rlabel metal2 373 -1294 373 -1294 0 net=2513
rlabel metal2 499 -1294 499 -1294 0 net=4967
rlabel metal2 772 -1294 772 -1294 0 net=4471
rlabel metal2 842 -1294 842 -1294 0 net=6161
rlabel metal2 859 -1294 859 -1294 0 net=7644
rlabel metal2 1115 -1294 1115 -1294 0 net=7903
rlabel metal2 82 -1296 82 -1296 0 net=1613
rlabel metal2 187 -1296 187 -1296 0 net=8043
rlabel metal2 635 -1296 635 -1296 0 net=7261
rlabel metal2 1108 -1296 1108 -1296 0 net=7889
rlabel metal2 1129 -1296 1129 -1296 0 net=8191
rlabel metal2 1150 -1296 1150 -1296 0 net=9477
rlabel metal2 191 -1298 191 -1298 0 net=4205
rlabel metal2 558 -1298 558 -1298 0 net=8055
rlabel metal2 1143 -1298 1143 -1298 0 net=8267
rlabel metal2 1164 -1298 1164 -1298 0 net=8361
rlabel metal2 1192 -1298 1192 -1298 0 net=11447
rlabel metal2 191 -1300 191 -1300 0 net=7205
rlabel metal2 1031 -1300 1031 -1300 0 net=7529
rlabel metal2 1080 -1300 1080 -1300 0 net=7855
rlabel metal2 1164 -1300 1164 -1300 0 net=8773
rlabel metal2 1227 -1300 1227 -1300 0 net=10589
rlabel metal2 247 -1302 247 -1302 0 net=1585
rlabel metal2 338 -1302 338 -1302 0 net=2017
rlabel metal2 422 -1302 422 -1302 0 net=4013
rlabel metal2 950 -1302 950 -1302 0 net=11345
rlabel metal2 173 -1304 173 -1304 0 net=1913
rlabel metal2 359 -1304 359 -1304 0 net=3207
rlabel metal2 674 -1304 674 -1304 0 net=3971
rlabel metal2 950 -1304 950 -1304 0 net=6715
rlabel metal2 989 -1304 989 -1304 0 net=7251
rlabel metal2 1080 -1304 1080 -1304 0 net=8599
rlabel metal2 1206 -1304 1206 -1304 0 net=8827
rlabel metal2 1234 -1304 1234 -1304 0 net=10863
rlabel metal2 86 -1306 86 -1306 0 net=3461
rlabel metal2 695 -1306 695 -1306 0 net=5373
rlabel metal2 1241 -1306 1241 -1306 0 net=9225
rlabel metal2 86 -1308 86 -1308 0 net=4993
rlabel metal2 562 -1308 562 -1308 0 net=8645
rlabel metal2 247 -1310 247 -1310 0 net=3047
rlabel metal2 408 -1310 408 -1310 0 net=2485
rlabel metal2 926 -1310 926 -1310 0 net=9355
rlabel metal2 222 -1312 222 -1312 0 net=1517
rlabel metal2 324 -1312 324 -1312 0 net=5251
rlabel metal2 422 -1312 422 -1312 0 net=1809
rlabel metal2 898 -1312 898 -1312 0 net=6449
rlabel metal2 954 -1312 954 -1312 0 net=6933
rlabel metal2 1003 -1312 1003 -1312 0 net=8991
rlabel metal2 324 -1314 324 -1314 0 net=7141
rlabel metal2 1024 -1314 1024 -1314 0 net=9061
rlabel metal2 436 -1316 436 -1316 0 net=5239
rlabel metal2 849 -1316 849 -1316 0 net=6197
rlabel metal2 450 -1318 450 -1318 0 net=3103
rlabel metal2 485 -1318 485 -1318 0 net=3418
rlabel metal2 572 -1318 572 -1318 0 net=8883
rlabel metal2 450 -1320 450 -1320 0 net=7039
rlabel metal2 457 -1322 457 -1322 0 net=3363
rlabel metal2 555 -1322 555 -1322 0 net=5169
rlabel metal2 884 -1322 884 -1322 0 net=6757
rlabel metal2 401 -1324 401 -1324 0 net=2680
rlabel metal2 583 -1324 583 -1324 0 net=6139
rlabel metal2 905 -1324 905 -1324 0 net=6707
rlabel metal2 394 -1326 394 -1326 0 net=2297
rlabel metal2 429 -1326 429 -1326 0 net=6069
rlabel metal2 219 -1328 219 -1328 0 net=2753
rlabel metal2 457 -1328 457 -1328 0 net=3075
rlabel metal2 618 -1328 618 -1328 0 net=5501
rlabel metal2 394 -1330 394 -1330 0 net=3959
rlabel metal2 698 -1330 698 -1330 0 net=7843
rlabel metal2 37 -1332 37 -1332 0 net=5463
rlabel metal2 786 -1332 786 -1332 0 net=5745
rlabel metal2 492 -1334 492 -1334 0 net=3451
rlabel metal2 534 -1334 534 -1334 0 net=4317
rlabel metal2 233 -1336 233 -1336 0 net=3271
rlabel metal2 520 -1336 520 -1336 0 net=3665
rlabel metal2 646 -1336 646 -1336 0 net=3545
rlabel metal2 30 -1338 30 -1338 0 net=5679
rlabel metal2 520 -1338 520 -1338 0 net=5123
rlabel metal2 786 -1338 786 -1338 0 net=10334
rlabel metal2 30 -1340 30 -1340 0 net=5477
rlabel metal2 730 -1340 730 -1340 0 net=7567
rlabel metal2 1367 -1340 1367 -1340 0 net=10185
rlabel metal2 485 -1342 485 -1342 0 net=2373
rlabel metal2 1066 -1342 1066 -1342 0 net=8145
rlabel metal2 1381 -1342 1381 -1342 0 net=10203
rlabel metal2 1122 -1344 1122 -1344 0 net=8675
rlabel metal2 1388 -1344 1388 -1344 0 net=10249
rlabel metal2 1199 -1346 1199 -1346 0 net=10945
rlabel metal2 1395 -1348 1395 -1348 0 net=10457
rlabel metal2 1409 -1350 1409 -1350 0 net=10471
rlabel metal2 1416 -1352 1416 -1352 0 net=10741
rlabel metal2 1437 -1354 1437 -1354 0 net=11789
rlabel metal2 1563 -1356 1563 -1356 0 net=11851
rlabel metal2 817 -1358 817 -1358 0 net=11977
rlabel metal2 16 -1369 16 -1369 0 net=2546
rlabel metal2 121 -1369 121 -1369 0 net=6454
rlabel metal2 219 -1369 219 -1369 0 net=7262
rlabel metal2 1048 -1369 1048 -1369 0 net=7166
rlabel metal2 1104 -1369 1104 -1369 0 net=12330
rlabel metal2 1738 -1369 1738 -1369 0 net=7905
rlabel metal2 51 -1371 51 -1371 0 net=1728
rlabel metal2 100 -1371 100 -1371 0 net=5699
rlabel metal2 100 -1371 100 -1371 0 net=5699
rlabel metal2 107 -1371 107 -1371 0 net=3547
rlabel metal2 688 -1371 688 -1371 0 net=2797
rlabel metal2 688 -1371 688 -1371 0 net=2797
rlabel metal2 719 -1371 719 -1371 0 net=6198
rlabel metal2 1038 -1371 1038 -1371 0 net=7857
rlabel metal2 1146 -1371 1146 -1371 0 net=12086
rlabel metal2 1689 -1371 1689 -1371 0 net=12611
rlabel metal2 51 -1373 51 -1373 0 net=6241
rlabel metal2 159 -1373 159 -1373 0 net=3644
rlabel metal2 187 -1373 187 -1373 0 net=5234
rlabel metal2 814 -1373 814 -1373 0 net=8192
rlabel metal2 1164 -1373 1164 -1373 0 net=8775
rlabel metal2 1164 -1373 1164 -1373 0 net=8775
rlabel metal2 1199 -1373 1199 -1373 0 net=10141
rlabel metal2 1591 -1373 1591 -1373 0 net=11477
rlabel metal2 58 -1375 58 -1375 0 net=5503
rlabel metal2 646 -1375 646 -1375 0 net=4267
rlabel metal2 744 -1375 744 -1375 0 net=5037
rlabel metal2 744 -1375 744 -1375 0 net=5037
rlabel metal2 751 -1375 751 -1375 0 net=9566
rlabel metal2 1346 -1375 1346 -1375 0 net=10459
rlabel metal2 1591 -1375 1591 -1375 0 net=12009
rlabel metal2 65 -1377 65 -1377 0 net=1984
rlabel metal2 82 -1377 82 -1377 0 net=10168
rlabel metal2 1395 -1377 1395 -1377 0 net=10981
rlabel metal2 1528 -1377 1528 -1377 0 net=11317
rlabel metal2 79 -1379 79 -1379 0 net=6495
rlabel metal2 978 -1379 978 -1379 0 net=11270
rlabel metal2 1612 -1379 1612 -1379 0 net=12535
rlabel metal2 93 -1381 93 -1381 0 net=5125
rlabel metal2 551 -1381 551 -1381 0 net=4014
rlabel metal2 849 -1381 849 -1381 0 net=9572
rlabel metal2 1374 -1381 1374 -1381 0 net=10473
rlabel metal2 1437 -1381 1437 -1381 0 net=11791
rlabel metal2 1612 -1381 1612 -1381 0 net=12099
rlabel metal2 124 -1383 124 -1383 0 net=1788
rlabel metal2 751 -1383 751 -1383 0 net=5171
rlabel metal2 761 -1383 761 -1383 0 net=7694
rlabel metal2 1647 -1383 1647 -1383 0 net=12517
rlabel metal2 149 -1385 149 -1385 0 net=4347
rlabel metal2 831 -1385 831 -1385 0 net=8488
rlabel metal2 1227 -1385 1227 -1385 0 net=8885
rlabel metal2 1500 -1385 1500 -1385 0 net=11769
rlabel metal2 1626 -1385 1626 -1385 0 net=12369
rlabel metal2 156 -1387 156 -1387 0 net=3563
rlabel metal2 194 -1387 194 -1387 0 net=1586
rlabel metal2 289 -1387 289 -1387 0 net=3177
rlabel metal2 478 -1387 478 -1387 0 net=3104
rlabel metal2 520 -1387 520 -1387 0 net=7253
rlabel metal2 1034 -1387 1034 -1387 0 net=12595
rlabel metal2 103 -1389 103 -1389 0 net=259
rlabel metal2 1066 -1389 1066 -1389 0 net=8147
rlabel metal2 1108 -1389 1108 -1389 0 net=9121
rlabel metal2 1402 -1389 1402 -1389 0 net=10365
rlabel metal2 156 -1391 156 -1391 0 net=1490
rlabel metal2 317 -1391 317 -1391 0 net=4983
rlabel metal2 625 -1391 625 -1391 0 net=4021
rlabel metal2 758 -1391 758 -1391 0 net=10261
rlabel metal2 1556 -1391 1556 -1391 0 net=11853
rlabel metal2 170 -1393 170 -1393 0 net=5288
rlabel metal2 219 -1393 219 -1393 0 net=4955
rlabel metal2 324 -1393 324 -1393 0 net=7142
rlabel metal2 786 -1393 786 -1393 0 net=8557
rlabel metal2 1202 -1393 1202 -1393 0 net=12484
rlabel metal2 114 -1395 114 -1395 0 net=6843
rlabel metal2 222 -1395 222 -1395 0 net=10032
rlabel metal2 1563 -1395 1563 -1395 0 net=12217
rlabel metal2 114 -1397 114 -1397 0 net=2761
rlabel metal2 789 -1397 789 -1397 0 net=1685
rlabel metal2 982 -1397 982 -1397 0 net=12688
rlabel metal2 170 -1399 170 -1399 0 net=4149
rlabel metal2 817 -1399 817 -1399 0 net=9131
rlabel metal2 1227 -1399 1227 -1399 0 net=9175
rlabel metal2 1339 -1399 1339 -1399 0 net=10205
rlabel metal2 1584 -1399 1584 -1399 0 net=10825
rlabel metal2 1731 -1399 1731 -1399 0 net=11111
rlabel metal2 163 -1401 163 -1401 0 net=3351
rlabel metal2 821 -1401 821 -1401 0 net=9696
rlabel metal2 1381 -1401 1381 -1401 0 net=10865
rlabel metal2 1584 -1401 1584 -1401 0 net=4943
rlabel metal2 163 -1403 163 -1403 0 net=1799
rlabel metal2 257 -1403 257 -1403 0 net=6820
rlabel metal2 849 -1403 849 -1403 0 net=6095
rlabel metal2 919 -1403 919 -1403 0 net=860
rlabel metal2 198 -1405 198 -1405 0 net=3508
rlabel metal2 555 -1405 555 -1405 0 net=5746
rlabel metal2 919 -1405 919 -1405 0 net=6451
rlabel metal2 982 -1405 982 -1405 0 net=7041
rlabel metal2 1003 -1405 1003 -1405 0 net=5777
rlabel metal2 1216 -1405 1216 -1405 0 net=11694
rlabel metal2 54 -1407 54 -1407 0 net=7279
rlabel metal2 1006 -1407 1006 -1407 0 net=10590
rlabel metal2 1507 -1407 1507 -1407 0 net=11873
rlabel metal2 135 -1409 135 -1409 0 net=1615
rlabel metal2 201 -1409 201 -1409 0 net=11127
rlabel metal2 1472 -1409 1472 -1409 0 net=11979
rlabel metal2 135 -1411 135 -1411 0 net=1549
rlabel metal2 226 -1411 226 -1411 0 net=2595
rlabel metal2 310 -1411 310 -1411 0 net=3077
rlabel metal2 471 -1411 471 -1411 0 net=2375
rlabel metal2 506 -1411 506 -1411 0 net=3947
rlabel metal2 558 -1411 558 -1411 0 net=11864
rlabel metal2 1598 -1411 1598 -1411 0 net=12705
rlabel metal2 142 -1413 142 -1413 0 net=1603
rlabel metal2 229 -1413 229 -1413 0 net=2492
rlabel metal2 366 -1413 366 -1413 0 net=3577
rlabel metal2 541 -1413 541 -1413 0 net=3711
rlabel metal2 1010 -1413 1010 -1413 0 net=7783
rlabel metal2 1066 -1413 1066 -1413 0 net=7891
rlabel metal2 1157 -1413 1157 -1413 0 net=7430
rlabel metal2 191 -1415 191 -1415 0 net=7206
rlabel metal2 215 -1415 215 -1415 0 net=3055
rlabel metal2 380 -1415 380 -1415 0 net=3217
rlabel metal2 562 -1415 562 -1415 0 net=6903
rlabel metal2 891 -1415 891 -1415 0 net=6709
rlabel metal2 1010 -1415 1010 -1415 0 net=7409
rlabel metal2 1115 -1415 1115 -1415 0 net=8269
rlabel metal2 1157 -1415 1157 -1415 0 net=8647
rlabel metal2 1213 -1415 1213 -1415 0 net=9227
rlabel metal2 1332 -1415 1332 -1415 0 net=11565
rlabel metal2 37 -1417 37 -1417 0 net=8841
rlabel metal2 240 -1417 240 -1417 0 net=4169
rlabel metal2 380 -1417 380 -1417 0 net=3365
rlabel metal2 562 -1417 562 -1417 0 net=4345
rlabel metal2 730 -1417 730 -1417 0 net=7569
rlabel metal2 933 -1417 933 -1417 0 net=10191
rlabel metal2 1318 -1417 1318 -1417 0 net=9536
rlabel metal2 86 -1419 86 -1419 0 net=4995
rlabel metal2 922 -1419 922 -1419 0 net=9356
rlabel metal2 1248 -1419 1248 -1419 0 net=9311
rlabel metal2 1318 -1419 1318 -1419 0 net=10743
rlabel metal2 1430 -1419 1430 -1419 0 net=11015
rlabel metal2 1479 -1419 1479 -1419 0 net=11969
rlabel metal2 86 -1421 86 -1421 0 net=5347
rlabel metal2 950 -1421 950 -1421 0 net=11327
rlabel metal2 1479 -1421 1479 -1421 0 net=12119
rlabel metal2 254 -1423 254 -1423 0 net=2861
rlabel metal2 387 -1423 387 -1423 0 net=5535
rlabel metal2 954 -1423 954 -1423 0 net=6759
rlabel metal2 1017 -1423 1017 -1423 0 net=12547
rlabel metal2 61 -1425 61 -1425 0 net=2727
rlabel metal2 408 -1425 408 -1425 0 net=5253
rlabel metal2 793 -1425 793 -1425 0 net=5369
rlabel metal2 968 -1425 968 -1425 0 net=7311
rlabel metal2 1059 -1425 1059 -1425 0 net=8057
rlabel metal2 1192 -1425 1192 -1425 0 net=9245
rlabel metal2 1276 -1425 1276 -1425 0 net=11861
rlabel metal2 268 -1427 268 -1427 0 net=1518
rlabel metal2 1129 -1427 1129 -1427 0 net=8363
rlabel metal2 1255 -1427 1255 -1427 0 net=9479
rlabel metal2 1416 -1427 1416 -1427 0 net=11347
rlabel metal2 1538 -1427 1538 -1427 0 net=4099
rlabel metal2 268 -1429 268 -1429 0 net=2633
rlabel metal2 408 -1429 408 -1429 0 net=5393
rlabel metal2 611 -1429 611 -1429 0 net=4115
rlabel metal2 1017 -1429 1017 -1429 0 net=7531
rlabel metal2 1080 -1429 1080 -1429 0 net=8601
rlabel metal2 1171 -1429 1171 -1429 0 net=8829
rlabel metal2 1262 -1429 1262 -1429 0 net=9519
rlabel metal2 1577 -1429 1577 -1429 0 net=11989
rlabel metal2 184 -1431 184 -1431 0 net=12161
rlabel metal2 275 -1433 275 -1433 0 net=3544
rlabel metal2 499 -1433 499 -1433 0 net=8045
rlabel metal2 975 -1433 975 -1433 0 net=7845
rlabel metal2 1143 -1433 1143 -1433 0 net=12181
rlabel metal2 275 -1435 275 -1435 0 net=4925
rlabel metal2 1020 -1435 1020 -1435 0 net=8676
rlabel metal2 1143 -1435 1143 -1435 0 net=8577
rlabel metal2 1297 -1435 1297 -1435 0 net=11285
rlabel metal2 296 -1437 296 -1437 0 net=4207
rlabel metal2 478 -1437 478 -1437 0 net=9297
rlabel metal2 1304 -1437 1304 -1437 0 net=11047
rlabel metal2 1360 -1437 1360 -1437 0 net=10075
rlabel metal2 44 -1439 44 -1439 0 net=3333
rlabel metal2 499 -1439 499 -1439 0 net=4319
rlabel metal2 569 -1439 569 -1439 0 net=7400
rlabel metal2 1178 -1439 1178 -1439 0 net=8993
rlabel metal2 1353 -1439 1353 -1439 0 net=10947
rlabel metal2 44 -1441 44 -1441 0 net=6683
rlabel metal2 415 -1441 415 -1441 0 net=2018
rlabel metal2 597 -1441 597 -1441 0 net=34
rlabel metal2 779 -1441 779 -1441 0 net=7939
rlabel metal2 1185 -1441 1185 -1441 0 net=9939
rlabel metal2 1360 -1441 1360 -1441 0 net=11079
rlabel metal2 72 -1443 72 -1443 0 net=11149
rlabel metal2 240 -1443 240 -1443 0 net=1611
rlabel metal2 1045 -1443 1045 -1443 0 net=10392
rlabel metal2 1465 -1443 1465 -1443 0 net=12057
rlabel metal2 247 -1445 247 -1445 0 net=3048
rlabel metal2 436 -1445 436 -1445 0 net=5240
rlabel metal2 1052 -1445 1052 -1445 0 net=9063
rlabel metal2 1444 -1445 1444 -1445 0 net=11281
rlabel metal2 247 -1447 247 -1447 0 net=1915
rlabel metal2 436 -1447 436 -1447 0 net=4053
rlabel metal2 947 -1447 947 -1447 0 net=12680
rlabel metal2 261 -1449 261 -1449 0 net=2169
rlabel metal2 450 -1449 450 -1449 0 net=4287
rlabel metal2 674 -1449 674 -1449 0 net=3463
rlabel metal2 261 -1451 261 -1451 0 net=1857
rlabel metal2 453 -1451 453 -1451 0 net=2486
rlabel metal2 1241 -1451 1241 -1451 0 net=9421
rlabel metal2 1458 -1451 1458 -1451 0 net=11599
rlabel metal2 1710 -1451 1710 -1451 0 net=12589
rlabel metal2 233 -1453 233 -1453 0 net=5681
rlabel metal2 1283 -1453 1283 -1453 0 net=10187
rlabel metal2 1486 -1453 1486 -1453 0 net=11449
rlabel metal2 1542 -1453 1542 -1453 0 net=11835
rlabel metal2 1643 -1453 1643 -1453 0 net=11119
rlabel metal2 233 -1455 233 -1455 0 net=1811
rlabel metal2 457 -1455 457 -1455 0 net=6647
rlabel metal2 1367 -1455 1367 -1455 0 net=11195
rlabel metal2 1549 -1455 1549 -1455 0 net=8008
rlabel metal2 331 -1457 331 -1457 0 net=2183
rlabel metal2 569 -1457 569 -1457 0 net=3835
rlabel metal2 604 -1457 604 -1457 0 net=5769
rlabel metal2 1388 -1457 1388 -1457 0 net=10251
rlabel metal2 422 -1459 422 -1459 0 net=2979
rlabel metal2 460 -1461 460 -1461 0 net=9357
rlabel metal2 513 -1463 513 -1463 0 net=9751
rlabel metal2 527 -1465 527 -1465 0 net=3453
rlabel metal2 653 -1465 653 -1465 0 net=4371
rlabel metal2 681 -1465 681 -1465 0 net=4473
rlabel metal2 852 -1465 852 -1465 0 net=12723
rlabel metal2 373 -1467 373 -1467 0 net=2515
rlabel metal2 534 -1467 534 -1467 0 net=2931
rlabel metal2 870 -1467 870 -1467 0 net=5851
rlabel metal2 373 -1469 373 -1469 0 net=3273
rlabel metal2 548 -1469 548 -1469 0 net=4835
rlabel metal2 30 -1471 30 -1471 0 net=5479
rlabel metal2 576 -1471 576 -1471 0 net=5465
rlabel metal2 877 -1471 877 -1471 0 net=6071
rlabel metal2 30 -1473 30 -1473 0 net=9537
rlabel metal2 576 -1473 576 -1473 0 net=4037
rlabel metal2 653 -1473 653 -1473 0 net=11066
rlabel metal2 131 -1475 131 -1475 0 net=3666
rlabel metal2 590 -1475 590 -1475 0 net=5243
rlabel metal2 394 -1477 394 -1477 0 net=3961
rlabel metal2 632 -1477 632 -1477 0 net=6935
rlabel metal2 394 -1479 394 -1479 0 net=2755
rlabel metal2 443 -1479 443 -1479 0 net=7945
rlabel metal2 359 -1481 359 -1481 0 net=3209
rlabel metal2 443 -1481 443 -1481 0 net=4675
rlabel metal2 726 -1481 726 -1481 0 net=8317
rlabel metal2 352 -1483 352 -1483 0 net=3411
rlabel metal2 695 -1483 695 -1483 0 net=5375
rlabel metal2 352 -1485 352 -1485 0 net=2299
rlabel metal2 695 -1485 695 -1485 0 net=4969
rlabel metal2 740 -1485 740 -1485 0 net=10919
rlabel metal2 345 -1487 345 -1487 0 net=1957
rlabel metal2 702 -1487 702 -1487 0 net=3603
rlabel metal2 884 -1487 884 -1487 0 net=6141
rlabel metal2 912 -1487 912 -1487 0 net=7213
rlabel metal2 23 -1489 23 -1489 0 net=2827
rlabel metal2 754 -1489 754 -1489 0 net=6575
rlabel metal2 856 -1489 856 -1489 0 net=6163
rlabel metal2 912 -1489 912 -1489 0 net=6717
rlabel metal2 23 -1491 23 -1491 0 net=10599
rlabel metal2 856 -1491 856 -1491 0 net=5763
rlabel metal2 961 -1491 961 -1491 0 net=6981
rlabel metal2 128 -1493 128 -1493 0 net=10207
rlabel metal2 772 -1495 772 -1495 0 net=3972
rlabel metal2 709 -1497 709 -1497 0 net=4711
rlabel metal2 709 -1499 709 -1499 0 net=7445
rlabel metal2 23 -1510 23 -1510 0 net=10600
rlabel metal2 240 -1510 240 -1510 0 net=1612
rlabel metal2 352 -1510 352 -1510 0 net=2301
rlabel metal2 352 -1510 352 -1510 0 net=2301
rlabel metal2 373 -1510 373 -1510 0 net=3275
rlabel metal2 401 -1510 401 -1510 0 net=1958
rlabel metal2 460 -1510 460 -1510 0 net=9176
rlabel metal2 1248 -1510 1248 -1510 0 net=9313
rlabel metal2 1248 -1510 1248 -1510 0 net=9313
rlabel metal2 1374 -1510 1374 -1510 0 net=10475
rlabel metal2 1374 -1510 1374 -1510 0 net=10475
rlabel metal2 1437 -1510 1437 -1510 0 net=11129
rlabel metal2 1437 -1510 1437 -1510 0 net=11129
rlabel metal2 1451 -1510 1451 -1510 0 net=11329
rlabel metal2 1486 -1510 1486 -1510 0 net=11451
rlabel metal2 1486 -1510 1486 -1510 0 net=11451
rlabel metal2 1521 -1510 1521 -1510 0 net=12724
rlabel metal2 1584 -1510 1584 -1510 0 net=10826
rlabel metal2 1706 -1510 1706 -1510 0 net=11120
rlabel metal2 1801 -1510 1801 -1510 0 net=7907
rlabel metal2 23 -1512 23 -1512 0 net=5897
rlabel metal2 436 -1512 436 -1512 0 net=4054
rlabel metal2 779 -1512 779 -1512 0 net=5467
rlabel metal2 866 -1512 866 -1512 0 net=10252
rlabel metal2 1451 -1512 1451 -1512 0 net=11981
rlabel metal2 1521 -1512 1521 -1512 0 net=11379
rlabel metal2 1619 -1512 1619 -1512 0 net=12163
rlabel metal2 1619 -1512 1619 -1512 0 net=12163
rlabel metal2 1640 -1512 1640 -1512 0 net=11112
rlabel metal2 37 -1514 37 -1514 0 net=8842
rlabel metal2 737 -1514 737 -1514 0 net=9132
rlabel metal2 1227 -1514 1227 -1514 0 net=9481
rlabel metal2 1304 -1514 1304 -1514 0 net=11049
rlabel metal2 1528 -1514 1528 -1514 0 net=11793
rlabel metal2 1528 -1514 1528 -1514 0 net=11793
rlabel metal2 1535 -1514 1535 -1514 0 net=11478
rlabel metal2 37 -1516 37 -1516 0 net=11557
rlabel metal2 93 -1516 93 -1516 0 net=5127
rlabel metal2 373 -1516 373 -1516 0 net=3579
rlabel metal2 492 -1516 492 -1516 0 net=5480
rlabel metal2 681 -1516 681 -1516 0 net=4474
rlabel metal2 1020 -1516 1020 -1516 0 net=12058
rlabel metal2 1535 -1516 1535 -1516 0 net=11837
rlabel metal2 1577 -1516 1577 -1516 0 net=11991
rlabel metal2 1598 -1516 1598 -1516 0 net=12707
rlabel metal2 51 -1518 51 -1518 0 net=6242
rlabel metal2 646 -1518 646 -1518 0 net=4269
rlabel metal2 646 -1518 646 -1518 0 net=4269
rlabel metal2 688 -1518 688 -1518 0 net=2798
rlabel metal2 961 -1518 961 -1518 0 net=6983
rlabel metal2 961 -1518 961 -1518 0 net=6983
rlabel metal2 1031 -1518 1031 -1518 0 net=10142
rlabel metal2 1255 -1518 1255 -1518 0 net=9521
rlabel metal2 1454 -1518 1454 -1518 0 net=1
rlabel metal2 1507 -1518 1507 -1518 0 net=11875
rlabel metal2 1577 -1518 1577 -1518 0 net=12101
rlabel metal2 1640 -1518 1640 -1518 0 net=12519
rlabel metal2 1650 -1518 1650 -1518 0 net=3464
rlabel metal2 51 -1520 51 -1520 0 net=1859
rlabel metal2 264 -1520 264 -1520 0 net=7254
rlabel metal2 527 -1520 527 -1520 0 net=2516
rlabel metal2 695 -1520 695 -1520 0 net=4971
rlabel metal2 695 -1520 695 -1520 0 net=4971
rlabel metal2 716 -1520 716 -1520 0 net=8943
rlabel metal2 1311 -1520 1311 -1520 0 net=10209
rlabel metal2 1591 -1520 1591 -1520 0 net=12011
rlabel metal2 1612 -1520 1612 -1520 0 net=12371
rlabel metal2 1643 -1520 1643 -1520 0 net=2155
rlabel metal2 1717 -1520 1717 -1520 0 net=12591
rlabel metal2 58 -1522 58 -1522 0 net=5504
rlabel metal2 989 -1522 989 -1522 0 net=7215
rlabel metal2 1034 -1522 1034 -1522 0 net=9122
rlabel metal2 1157 -1522 1157 -1522 0 net=8649
rlabel metal2 1311 -1522 1311 -1522 0 net=10745
rlabel metal2 1479 -1522 1479 -1522 0 net=12121
rlabel metal2 1668 -1522 1668 -1522 0 net=12597
rlabel metal2 1703 -1522 1703 -1522 0 net=4945
rlabel metal2 65 -1524 65 -1524 0 net=5853
rlabel metal2 880 -1524 880 -1524 0 net=7532
rlabel metal2 1045 -1524 1045 -1524 0 net=7893
rlabel metal2 1171 -1524 1171 -1524 0 net=8831
rlabel metal2 1171 -1524 1171 -1524 0 net=8831
rlabel metal2 1188 -1524 1188 -1524 0 net=11600
rlabel metal2 1514 -1524 1514 -1524 0 net=12183
rlabel metal2 1633 -1524 1633 -1524 0 net=11318
rlabel metal2 93 -1526 93 -1526 0 net=3713
rlabel metal2 607 -1526 607 -1526 0 net=6452
rlabel metal2 936 -1526 936 -1526 0 net=9940
rlabel metal2 1192 -1526 1192 -1526 0 net=9247
rlabel metal2 1318 -1526 1318 -1526 0 net=7335
rlabel metal2 124 -1528 124 -1528 0 net=206
rlabel metal2 380 -1528 380 -1528 0 net=3367
rlabel metal2 481 -1528 481 -1528 0 net=1328
rlabel metal2 44 -1530 44 -1530 0 net=6684
rlabel metal2 128 -1530 128 -1530 0 net=1616
rlabel metal2 212 -1530 212 -1530 0 net=3165
rlabel metal2 303 -1530 303 -1530 0 net=2863
rlabel metal2 303 -1530 303 -1530 0 net=2863
rlabel metal2 310 -1530 310 -1530 0 net=3078
rlabel metal2 737 -1530 737 -1530 0 net=5039
rlabel metal2 747 -1530 747 -1530 0 net=1150
rlabel metal2 947 -1530 947 -1530 0 net=9358
rlabel metal2 1332 -1530 1332 -1530 0 net=11567
rlabel metal2 1563 -1530 1563 -1530 0 net=12219
rlabel metal2 44 -1532 44 -1532 0 net=4429
rlabel metal2 79 -1532 79 -1532 0 net=6497
rlabel metal2 131 -1532 131 -1532 0 net=4208
rlabel metal2 415 -1532 415 -1532 0 net=3836
rlabel metal2 611 -1532 611 -1532 0 net=4117
rlabel metal2 702 -1532 702 -1532 0 net=3605
rlabel metal2 723 -1532 723 -1532 0 net=11080
rlabel metal2 1416 -1532 1416 -1532 0 net=11349
rlabel metal2 1556 -1532 1556 -1532 0 net=11855
rlabel metal2 79 -1534 79 -1534 0 net=2493
rlabel metal2 1048 -1534 1048 -1534 0 net=10188
rlabel metal2 1325 -1534 1325 -1534 0 net=10263
rlabel metal2 1395 -1534 1395 -1534 0 net=10983
rlabel metal2 1430 -1534 1430 -1534 0 net=11017
rlabel metal2 1556 -1534 1556 -1534 0 net=11971
rlabel metal2 149 -1536 149 -1536 0 net=4349
rlabel metal2 625 -1536 625 -1536 0 net=4497
rlabel metal2 831 -1536 831 -1536 0 net=12151
rlabel metal2 135 -1538 135 -1538 0 net=1551
rlabel metal2 156 -1538 156 -1538 0 net=11941
rlabel metal2 159 -1540 159 -1540 0 net=5427
rlabel metal2 415 -1540 415 -1540 0 net=2377
rlabel metal2 506 -1540 506 -1540 0 net=3219
rlabel metal2 569 -1540 569 -1540 0 net=4101
rlabel metal2 177 -1542 177 -1542 0 net=3565
rlabel metal2 177 -1542 177 -1542 0 net=3565
rlabel metal2 184 -1542 184 -1542 0 net=4676
rlabel metal2 506 -1542 506 -1542 0 net=3949
rlabel metal2 604 -1542 604 -1542 0 net=5771
rlabel metal2 709 -1542 709 -1542 0 net=7447
rlabel metal2 1073 -1542 1073 -1542 0 net=7847
rlabel metal2 1206 -1542 1206 -1542 0 net=9299
rlabel metal2 1290 -1542 1290 -1542 0 net=10193
rlabel metal2 1381 -1542 1381 -1542 0 net=10867
rlabel metal2 1493 -1542 1493 -1542 0 net=10077
rlabel metal2 1654 -1542 1654 -1542 0 net=12537
rlabel metal2 184 -1544 184 -1544 0 net=11085
rlabel metal2 1661 -1544 1661 -1544 0 net=12549
rlabel metal2 191 -1546 191 -1546 0 net=3979
rlabel metal2 422 -1546 422 -1546 0 net=2981
rlabel metal2 544 -1546 544 -1546 0 net=10701
rlabel metal2 1675 -1546 1675 -1546 0 net=12613
rlabel metal2 86 -1548 86 -1548 0 net=5349
rlabel metal2 436 -1548 436 -1548 0 net=7281
rlabel metal2 1059 -1548 1059 -1548 0 net=8059
rlabel metal2 1164 -1548 1164 -1548 0 net=8777
rlabel metal2 1269 -1548 1269 -1548 0 net=9753
rlabel metal2 1685 -1548 1685 -1548 0 net=7059
rlabel metal2 68 -1550 68 -1550 0 net=1639
rlabel metal2 191 -1550 191 -1550 0 net=1917
rlabel metal2 387 -1550 387 -1550 0 net=2729
rlabel metal2 478 -1550 478 -1550 0 net=11553
rlabel metal2 194 -1552 194 -1552 0 net=11137
rlabel metal2 198 -1554 198 -1554 0 net=4289
rlabel metal2 653 -1554 653 -1554 0 net=6333
rlabel metal2 947 -1554 947 -1554 0 net=6605
rlabel metal2 205 -1556 205 -1556 0 net=6845
rlabel metal2 968 -1556 968 -1556 0 net=7313
rlabel metal2 996 -1556 996 -1556 0 net=8319
rlabel metal2 1178 -1556 1178 -1556 0 net=8995
rlabel metal2 121 -1558 121 -1558 0 net=9759
rlabel metal2 212 -1558 212 -1558 0 net=4171
rlabel metal2 387 -1558 387 -1558 0 net=3335
rlabel metal2 541 -1558 541 -1558 0 net=170
rlabel metal2 1136 -1558 1136 -1558 0 net=8559
rlabel metal2 1185 -1558 1185 -1558 0 net=10087
rlabel metal2 121 -1560 121 -1560 0 net=2333
rlabel metal2 215 -1560 215 -1560 0 net=5394
rlabel metal2 443 -1560 443 -1560 0 net=4346
rlabel metal2 632 -1560 632 -1560 0 net=6937
rlabel metal2 1062 -1560 1062 -1560 0 net=11282
rlabel metal2 219 -1562 219 -1562 0 net=4957
rlabel metal2 709 -1562 709 -1562 0 net=6905
rlabel metal2 863 -1562 863 -1562 0 net=11007
rlabel metal2 1367 -1562 1367 -1562 0 net=11197
rlabel metal2 30 -1564 30 -1564 0 net=9538
rlabel metal2 222 -1564 222 -1564 0 net=1097
rlabel metal2 740 -1564 740 -1564 0 net=5376
rlabel metal2 1136 -1564 1136 -1564 0 net=8579
rlabel metal2 1346 -1564 1346 -1564 0 net=10461
rlabel metal2 30 -1566 30 -1566 0 net=4817
rlabel metal2 653 -1566 653 -1566 0 net=4373
rlabel metal2 754 -1566 754 -1566 0 net=9064
rlabel metal2 1101 -1566 1101 -1566 0 net=8603
rlabel metal2 1346 -1566 1346 -1566 0 net=10367
rlabel metal2 233 -1568 233 -1568 0 net=1813
rlabel metal2 324 -1568 324 -1568 0 net=2101
rlabel metal2 863 -1568 863 -1568 0 net=8287
rlabel metal2 1388 -1568 1388 -1568 0 net=10921
rlabel metal2 233 -1570 233 -1570 0 net=3211
rlabel metal2 446 -1570 446 -1570 0 net=4617
rlabel metal2 499 -1570 499 -1570 0 net=4321
rlabel metal2 667 -1570 667 -1570 0 net=8547
rlabel metal2 1388 -1570 1388 -1570 0 net=11771
rlabel metal2 247 -1572 247 -1572 0 net=4717
rlabel metal2 429 -1572 429 -1572 0 net=7983
rlabel metal2 870 -1572 870 -1572 0 net=5779
rlabel metal2 1094 -1572 1094 -1572 0 net=8149
rlabel metal2 1409 -1572 1409 -1572 0 net=8887
rlabel metal2 275 -1574 275 -1574 0 net=4927
rlabel metal2 464 -1574 464 -1574 0 net=7151
rlabel metal2 758 -1574 758 -1574 0 net=5764
rlabel metal2 894 -1574 894 -1574 0 net=9422
rlabel metal2 1353 -1574 1353 -1574 0 net=10949
rlabel metal2 142 -1576 142 -1576 0 net=1605
rlabel metal2 499 -1576 499 -1576 0 net=3353
rlabel metal2 730 -1576 730 -1576 0 net=4997
rlabel metal2 779 -1576 779 -1576 0 net=4721
rlabel metal2 1094 -1576 1094 -1576 0 net=8365
rlabel metal2 1297 -1576 1297 -1576 0 net=11287
rlabel metal2 142 -1578 142 -1578 0 net=1801
rlabel metal2 548 -1578 548 -1578 0 net=4837
rlabel metal2 730 -1578 730 -1578 0 net=10206
rlabel metal2 163 -1580 163 -1580 0 net=8927
rlabel metal2 1297 -1580 1297 -1580 0 net=10423
rlabel metal2 548 -1582 548 -1582 0 net=3962
rlabel metal2 590 -1582 590 -1582 0 net=5245
rlabel metal2 786 -1582 786 -1582 0 net=7570
rlabel metal2 940 -1582 940 -1582 0 net=1686
rlabel metal2 1115 -1582 1115 -1582 0 net=8271
rlabel metal2 187 -1584 187 -1584 0 net=5017
rlabel metal2 639 -1584 639 -1584 0 net=6711
rlabel metal2 905 -1584 905 -1584 0 net=6649
rlabel metal2 905 -1584 905 -1584 0 net=6649
rlabel metal2 912 -1584 912 -1584 0 net=6719
rlabel metal2 940 -1584 940 -1584 0 net=7941
rlabel metal2 1087 -1584 1087 -1584 0 net=7947
rlabel metal2 1125 -1584 1125 -1584 0 net=8109
rlabel metal2 492 -1586 492 -1586 0 net=2599
rlabel metal2 898 -1586 898 -1586 0 net=6165
rlabel metal2 975 -1586 975 -1586 0 net=7599
rlabel metal2 1080 -1586 1080 -1586 0 net=636
rlabel metal2 562 -1588 562 -1588 0 net=4039
rlabel metal2 583 -1588 583 -1588 0 net=4023
rlabel metal2 786 -1588 786 -1588 0 net=5289
rlabel metal2 884 -1588 884 -1588 0 net=6143
rlabel metal2 954 -1588 954 -1588 0 net=6761
rlabel metal2 1024 -1588 1024 -1588 0 net=7785
rlabel metal2 135 -1590 135 -1590 0 net=11651
rlabel metal2 849 -1590 849 -1590 0 net=6097
rlabel metal2 954 -1590 954 -1590 0 net=11862
rlabel metal2 450 -1592 450 -1592 0 net=5823
rlabel metal2 1010 -1592 1010 -1592 0 net=7411
rlabel metal2 1213 -1592 1213 -1592 0 net=9229
rlabel metal2 551 -1594 551 -1594 0 net=8677
rlabel metal2 576 -1596 576 -1596 0 net=5255
rlabel metal2 789 -1596 789 -1596 0 net=5682
rlabel metal2 982 -1596 982 -1596 0 net=7043
rlabel metal2 597 -1598 597 -1598 0 net=3455
rlabel metal2 800 -1598 800 -1598 0 net=8047
rlabel metal2 982 -1598 982 -1598 0 net=7859
rlabel metal2 72 -1600 72 -1600 0 net=11151
rlabel metal2 72 -1602 72 -1602 0 net=3431
rlabel metal2 618 -1602 618 -1602 0 net=4985
rlabel metal2 793 -1602 793 -1602 0 net=5371
rlabel metal2 807 -1602 807 -1602 0 net=6576
rlabel metal2 100 -1604 100 -1604 0 net=5701
rlabel metal2 772 -1604 772 -1604 0 net=4713
rlabel metal2 814 -1604 814 -1604 0 net=5537
rlabel metal2 100 -1606 100 -1606 0 net=8425
rlabel metal2 513 -1606 513 -1606 0 net=5403
rlabel metal2 114 -1608 114 -1608 0 net=2763
rlabel metal2 359 -1608 359 -1608 0 net=3413
rlabel metal2 555 -1608 555 -1608 0 net=4581
rlabel metal2 114 -1610 114 -1610 0 net=2185
rlabel metal2 359 -1610 359 -1610 0 net=3057
rlabel metal2 751 -1610 751 -1610 0 net=5173
rlabel metal2 166 -1612 166 -1612 0 net=1635
rlabel metal2 366 -1612 366 -1612 0 net=5803
rlabel metal2 170 -1614 170 -1614 0 net=4151
rlabel metal2 170 -1616 170 -1616 0 net=3179
rlabel metal2 107 -1618 107 -1618 0 net=3549
rlabel metal2 107 -1620 107 -1620 0 net=2757
rlabel metal2 268 -1622 268 -1622 0 net=2635
rlabel metal2 268 -1624 268 -1624 0 net=2597
rlabel metal2 282 -1626 282 -1626 0 net=2171
rlabel metal2 338 -1628 338 -1628 0 net=2829
rlabel metal2 345 -1630 345 -1630 0 net=2933
rlabel metal2 534 -1632 534 -1632 0 net=6073
rlabel metal2 331 -1634 331 -1634 0 net=7617
rlabel metal2 30 -1645 30 -1645 0 net=4818
rlabel metal2 324 -1645 324 -1645 0 net=2102
rlabel metal2 387 -1645 387 -1645 0 net=3336
rlabel metal2 660 -1645 660 -1645 0 net=3456
rlabel metal2 789 -1645 789 -1645 0 net=8843
rlabel metal2 1300 -1645 1300 -1645 0 net=11018
rlabel metal2 1549 -1645 1549 -1645 0 net=11943
rlabel metal2 1822 -1645 1822 -1645 0 net=7908
rlabel metal2 30 -1647 30 -1647 0 net=4291
rlabel metal2 219 -1647 219 -1647 0 net=865
rlabel metal2 548 -1647 548 -1647 0 net=2156
rlabel metal2 23 -1649 23 -1649 0 net=5899
rlabel metal2 236 -1649 236 -1649 0 net=12319
rlabel metal2 23 -1651 23 -1651 0 net=3213
rlabel metal2 275 -1651 275 -1651 0 net=1607
rlabel metal2 338 -1651 338 -1651 0 net=2831
rlabel metal2 338 -1651 338 -1651 0 net=2831
rlabel metal2 345 -1651 345 -1651 0 net=2935
rlabel metal2 345 -1651 345 -1651 0 net=2935
rlabel metal2 352 -1651 352 -1651 0 net=2302
rlabel metal2 551 -1651 551 -1651 0 net=7948
rlabel metal2 1122 -1651 1122 -1651 0 net=10315
rlabel metal2 1598 -1651 1598 -1651 0 net=12013
rlabel metal2 58 -1653 58 -1653 0 net=1503
rlabel metal2 800 -1653 800 -1653 0 net=5372
rlabel metal2 856 -1653 856 -1653 0 net=6099
rlabel metal2 891 -1653 891 -1653 0 net=12467
rlabel metal2 107 -1655 107 -1655 0 net=2759
rlabel metal2 954 -1655 954 -1655 0 net=5833
rlabel metal2 1125 -1655 1125 -1655 0 net=9522
rlabel metal2 1423 -1655 1423 -1655 0 net=11051
rlabel metal2 1605 -1655 1605 -1655 0 net=12153
rlabel metal2 93 -1657 93 -1657 0 net=3715
rlabel metal2 121 -1657 121 -1657 0 net=8832
rlabel metal2 1185 -1657 1185 -1657 0 net=1388
rlabel metal2 93 -1659 93 -1659 0 net=3255
rlabel metal2 576 -1659 576 -1659 0 net=5257
rlabel metal2 814 -1659 814 -1659 0 net=12520
rlabel metal2 1647 -1659 1647 -1659 0 net=12231
rlabel metal2 121 -1661 121 -1661 0 net=3977
rlabel metal2 782 -1661 782 -1661 0 net=11203
rlabel metal2 1619 -1661 1619 -1661 0 net=12165
rlabel metal2 124 -1663 124 -1663 0 net=1175
rlabel metal2 957 -1663 957 -1663 0 net=12105
rlabel metal2 135 -1665 135 -1665 0 net=11652
rlabel metal2 681 -1665 681 -1665 0 net=4118
rlabel metal2 835 -1665 835 -1665 0 net=8049
rlabel metal2 1185 -1665 1185 -1665 0 net=8779
rlabel metal2 1304 -1665 1304 -1665 0 net=10089
rlabel metal2 1451 -1665 1451 -1665 0 net=11983
rlabel metal2 135 -1667 135 -1667 0 net=2447
rlabel metal2 1066 -1667 1066 -1667 0 net=7448
rlabel metal2 1101 -1667 1101 -1667 0 net=8605
rlabel metal2 1332 -1667 1332 -1667 0 net=10265
rlabel metal2 1479 -1667 1479 -1667 0 net=11351
rlabel metal2 1626 -1667 1626 -1667 0 net=12185
rlabel metal2 159 -1669 159 -1669 0 net=996
rlabel metal2 590 -1669 590 -1669 0 net=5019
rlabel metal2 835 -1669 835 -1669 0 net=5825
rlabel metal2 859 -1669 859 -1669 0 net=8320
rlabel metal2 1003 -1669 1003 -1669 0 net=11856
rlabel metal2 1633 -1669 1633 -1669 0 net=12221
rlabel metal2 184 -1671 184 -1671 0 net=4172
rlabel metal2 275 -1671 275 -1671 0 net=2983
rlabel metal2 604 -1671 604 -1671 0 net=3235
rlabel metal2 863 -1671 863 -1671 0 net=7786
rlabel metal2 1101 -1671 1101 -1671 0 net=7061
rlabel metal2 1696 -1671 1696 -1671 0 net=12709
rlabel metal2 145 -1673 145 -1673 0 net=2371
rlabel metal2 187 -1673 187 -1673 0 net=6074
rlabel metal2 611 -1673 611 -1673 0 net=4351
rlabel metal2 674 -1673 674 -1673 0 net=5247
rlabel metal2 828 -1673 828 -1673 0 net=5469
rlabel metal2 877 -1673 877 -1673 0 net=11008
rlabel metal2 1374 -1673 1374 -1673 0 net=10477
rlabel metal2 1521 -1673 1521 -1673 0 net=11381
rlabel metal2 1650 -1673 1650 -1673 0 net=12592
rlabel metal2 44 -1675 44 -1675 0 net=4430
rlabel metal2 681 -1675 681 -1675 0 net=4723
rlabel metal2 786 -1675 786 -1675 0 net=5291
rlabel metal2 877 -1675 877 -1675 0 net=6651
rlabel metal2 950 -1675 950 -1675 0 net=11715
rlabel metal2 1654 -1675 1654 -1675 0 net=12539
rlabel metal2 44 -1677 44 -1677 0 net=6713
rlabel metal2 716 -1677 716 -1677 0 net=3606
rlabel metal2 779 -1677 779 -1677 0 net=827
rlabel metal2 880 -1677 880 -1677 0 net=10194
rlabel metal2 1395 -1677 1395 -1677 0 net=10869
rlabel metal2 1528 -1677 1528 -1677 0 net=11795
rlabel metal2 212 -1679 212 -1679 0 net=4583
rlabel metal2 611 -1679 611 -1679 0 net=5539
rlabel metal2 901 -1679 901 -1679 0 net=6391
rlabel metal2 1017 -1679 1017 -1679 0 net=8272
rlabel metal2 1146 -1679 1146 -1679 0 net=12102
rlabel metal2 1584 -1679 1584 -1679 0 net=11993
rlabel metal2 282 -1681 282 -1681 0 net=2173
rlabel metal2 282 -1681 282 -1681 0 net=2173
rlabel metal2 303 -1681 303 -1681 0 net=2865
rlabel metal2 352 -1681 352 -1681 0 net=2349
rlabel metal2 618 -1681 618 -1681 0 net=5703
rlabel metal2 947 -1681 947 -1681 0 net=6607
rlabel metal2 1020 -1681 1020 -1681 0 net=11093
rlabel metal2 1262 -1681 1262 -1681 0 net=8945
rlabel metal2 1402 -1681 1402 -1681 0 net=10923
rlabel metal2 1542 -1681 1542 -1681 0 net=11877
rlabel metal2 205 -1683 205 -1683 0 net=9761
rlabel metal2 1416 -1683 1416 -1683 0 net=10985
rlabel metal2 1661 -1683 1661 -1683 0 net=12551
rlabel metal2 37 -1685 37 -1685 0 net=11559
rlabel metal2 1668 -1685 1668 -1685 0 net=12599
rlabel metal2 37 -1687 37 -1687 0 net=3951
rlabel metal2 534 -1687 534 -1687 0 net=5361
rlabel metal2 1108 -1687 1108 -1687 0 net=12122
rlabel metal2 1675 -1687 1675 -1687 0 net=12615
rlabel metal2 79 -1689 79 -1689 0 net=2495
rlabel metal2 254 -1689 254 -1689 0 net=1637
rlabel metal2 331 -1689 331 -1689 0 net=7619
rlabel metal2 639 -1689 639 -1689 0 net=4271
rlabel metal2 716 -1689 716 -1689 0 net=7216
rlabel metal2 1038 -1689 1038 -1689 0 net=11153
rlabel metal2 1682 -1689 1682 -1689 0 net=4946
rlabel metal2 79 -1691 79 -1691 0 net=5805
rlabel metal2 387 -1691 387 -1691 0 net=2601
rlabel metal2 499 -1691 499 -1691 0 net=3355
rlabel metal2 646 -1691 646 -1691 0 net=4375
rlabel metal2 723 -1691 723 -1691 0 net=6801
rlabel metal2 1080 -1691 1080 -1691 0 net=9809
rlabel metal2 1437 -1691 1437 -1691 0 net=11131
rlabel metal2 1570 -1691 1570 -1691 0 net=10079
rlabel metal2 254 -1693 254 -1693 0 net=7153
rlabel metal2 485 -1693 485 -1693 0 net=3276
rlabel metal2 632 -1693 632 -1693 0 net=4323
rlabel metal2 747 -1693 747 -1693 0 net=9529
rlabel metal2 1444 -1693 1444 -1693 0 net=11199
rlabel metal2 331 -1695 331 -1695 0 net=3059
rlabel metal2 362 -1695 362 -1695 0 net=6459
rlabel metal2 1010 -1695 1010 -1695 0 net=7045
rlabel metal2 1129 -1695 1129 -1695 0 net=9315
rlabel metal2 1269 -1695 1269 -1695 0 net=8997
rlabel metal2 1388 -1695 1388 -1695 0 net=11773
rlabel metal2 366 -1697 366 -1697 0 net=5429
rlabel metal2 394 -1697 394 -1697 0 net=2636
rlabel metal2 807 -1697 807 -1697 0 net=5405
rlabel metal2 975 -1697 975 -1697 0 net=6763
rlabel metal2 1038 -1697 1038 -1697 0 net=5521
rlabel metal2 1136 -1697 1136 -1697 0 net=8581
rlabel metal2 1290 -1697 1290 -1697 0 net=9755
rlabel metal2 1472 -1697 1472 -1697 0 net=11331
rlabel metal2 394 -1699 394 -1699 0 net=4153
rlabel metal2 754 -1699 754 -1699 0 net=7835
rlabel metal2 1157 -1699 1157 -1699 0 net=8289
rlabel metal2 1493 -1699 1493 -1699 0 net=11555
rlabel metal2 401 -1701 401 -1701 0 net=3981
rlabel metal2 726 -1701 726 -1701 0 net=10675
rlabel metal2 1500 -1701 1500 -1701 0 net=8889
rlabel metal2 240 -1703 240 -1703 0 net=3167
rlabel metal2 408 -1703 408 -1703 0 net=4928
rlabel metal2 765 -1703 765 -1703 0 net=4987
rlabel metal2 824 -1703 824 -1703 0 net=6938
rlabel metal2 978 -1703 978 -1703 0 net=11385
rlabel metal2 114 -1705 114 -1705 0 net=2187
rlabel metal2 408 -1705 408 -1705 0 net=5581
rlabel metal2 898 -1705 898 -1705 0 net=6145
rlabel metal2 989 -1705 989 -1705 0 net=7315
rlabel metal2 1157 -1705 1157 -1705 0 net=7337
rlabel metal2 1339 -1705 1339 -1705 0 net=10425
rlabel metal2 1507 -1705 1507 -1705 0 net=10211
rlabel metal2 415 -1707 415 -1707 0 net=2379
rlabel metal2 457 -1707 457 -1707 0 net=3369
rlabel metal2 506 -1707 506 -1707 0 net=3489
rlabel metal2 758 -1707 758 -1707 0 net=4999
rlabel metal2 919 -1707 919 -1707 0 net=6335
rlabel metal2 1010 -1707 1010 -1707 0 net=8111
rlabel metal2 1164 -1707 1164 -1707 0 net=8549
rlabel metal2 1276 -1707 1276 -1707 0 net=9231
rlabel metal2 1381 -1707 1381 -1707 0 net=10703
rlabel metal2 1514 -1707 1514 -1707 0 net=11569
rlabel metal2 219 -1709 219 -1709 0 net=10771
rlabel metal2 1535 -1709 1535 -1709 0 net=11839
rlabel metal2 415 -1711 415 -1711 0 net=1993
rlabel metal2 635 -1711 635 -1711 0 net=9523
rlabel metal2 1409 -1711 1409 -1711 0 net=10951
rlabel metal2 1556 -1711 1556 -1711 0 net=11973
rlabel metal2 429 -1713 429 -1713 0 net=7985
rlabel metal2 1311 -1713 1311 -1713 0 net=10747
rlabel metal2 436 -1715 436 -1715 0 net=7282
rlabel metal2 758 -1715 758 -1715 0 net=5175
rlabel metal2 786 -1715 786 -1715 0 net=8633
rlabel metal2 1430 -1715 1430 -1715 0 net=11087
rlabel metal2 114 -1717 114 -1717 0 net=5065
rlabel metal2 849 -1717 849 -1717 0 net=5423
rlabel metal2 1178 -1717 1178 -1717 0 net=8561
rlabel metal2 1367 -1717 1367 -1717 0 net=10463
rlabel metal2 436 -1719 436 -1719 0 net=4103
rlabel metal2 695 -1719 695 -1719 0 net=4973
rlabel metal2 870 -1719 870 -1719 0 net=5781
rlabel metal2 933 -1719 933 -1719 0 net=6847
rlabel metal2 1206 -1719 1206 -1719 0 net=12372
rlabel metal2 89 -1721 89 -1721 0 net=6457
rlabel metal2 1220 -1721 1220 -1721 0 net=9249
rlabel metal2 1353 -1721 1353 -1721 0 net=11289
rlabel metal2 443 -1723 443 -1723 0 net=5603
rlabel metal2 443 -1723 443 -1723 0 net=5603
rlabel metal2 446 -1723 446 -1723 0 net=3414
rlabel metal2 541 -1723 541 -1723 0 net=3801
rlabel metal2 562 -1723 562 -1723 0 net=4041
rlabel metal2 695 -1723 695 -1723 0 net=4715
rlabel metal2 870 -1723 870 -1723 0 net=5505
rlabel metal2 1006 -1723 1006 -1723 0 net=9767
rlabel metal2 317 -1725 317 -1725 0 net=5129
rlabel metal2 933 -1725 933 -1725 0 net=6985
rlabel metal2 1024 -1725 1024 -1725 0 net=7413
rlabel metal2 268 -1727 268 -1727 0 net=2598
rlabel metal2 1027 -1727 1027 -1727 0 net=9181
rlabel metal2 1227 -1727 1227 -1727 0 net=9483
rlabel metal2 268 -1729 268 -1729 0 net=4737
rlabel metal2 562 -1729 562 -1729 0 net=3867
rlabel metal2 940 -1729 940 -1729 0 net=7943
rlabel metal2 1241 -1729 1241 -1729 0 net=8929
rlabel metal2 1283 -1729 1283 -1729 0 net=9301
rlabel metal2 100 -1731 100 -1731 0 net=8427
rlabel metal2 100 -1733 100 -1733 0 net=3181
rlabel metal2 261 -1733 261 -1733 0 net=5951
rlabel metal2 1045 -1733 1045 -1733 0 net=7895
rlabel metal2 1213 -1733 1213 -1733 0 net=8679
rlabel metal2 317 -1735 317 -1735 0 net=2077
rlabel metal2 453 -1737 453 -1737 0 net=8219
rlabel metal2 457 -1739 457 -1739 0 net=4619
rlabel metal2 485 -1739 485 -1739 0 net=3221
rlabel metal2 1045 -1739 1045 -1739 0 net=8651
rlabel metal2 163 -1741 163 -1741 0 net=8213
rlabel metal2 163 -1743 163 -1743 0 net=1919
rlabel metal2 289 -1743 289 -1743 0 net=3551
rlabel metal2 1052 -1743 1052 -1743 0 net=7601
rlabel metal2 1150 -1743 1150 -1743 0 net=8151
rlabel metal2 156 -1745 156 -1745 0 net=2335
rlabel metal2 222 -1745 222 -1745 0 net=2917
rlabel metal2 464 -1745 464 -1745 0 net=2731
rlabel metal2 478 -1745 478 -1745 0 net=4025
rlabel metal2 982 -1745 982 -1745 0 net=7861
rlabel metal2 156 -1747 156 -1747 0 net=4881
rlabel metal2 471 -1747 471 -1747 0 net=4499
rlabel metal2 912 -1747 912 -1747 0 net=6167
rlabel metal2 1052 -1747 1052 -1747 0 net=11452
rlabel metal2 170 -1749 170 -1749 0 net=5063
rlabel metal2 499 -1749 499 -1749 0 net=5971
rlabel metal2 1055 -1749 1055 -1749 0 net=11113
rlabel metal2 1465 -1749 1465 -1749 0 net=11139
rlabel metal2 513 -1751 513 -1751 0 net=4839
rlabel metal2 702 -1751 702 -1751 0 net=5773
rlabel metal2 1094 -1751 1094 -1751 0 net=8367
rlabel metal2 1346 -1751 1346 -1751 0 net=10369
rlabel metal2 296 -1753 296 -1753 0 net=1815
rlabel metal2 1192 -1753 1192 -1753 0 net=7849
rlabel metal2 226 -1755 226 -1755 0 net=2765
rlabel metal2 422 -1755 422 -1755 0 net=5350
rlabel metal2 1073 -1755 1073 -1755 0 net=8061
rlabel metal2 51 -1757 51 -1757 0 net=1861
rlabel metal2 422 -1757 422 -1757 0 net=5041
rlabel metal2 51 -1759 51 -1759 0 net=6721
rlabel metal2 65 -1761 65 -1761 0 net=5855
rlabel metal2 65 -1763 65 -1763 0 net=3581
rlabel metal2 583 -1763 583 -1763 0 net=10227
rlabel metal2 247 -1765 247 -1765 0 net=4719
rlabel metal2 625 -1765 625 -1765 0 net=4109
rlabel metal2 72 -1767 72 -1767 0 net=3433
rlabel metal2 667 -1767 667 -1767 0 net=3931
rlabel metal2 709 -1767 709 -1767 0 net=6907
rlabel metal2 72 -1769 72 -1769 0 net=12277
rlabel metal2 688 -1771 688 -1771 0 net=4959
rlabel metal2 128 -1773 128 -1773 0 net=6499
rlabel metal2 709 -1773 709 -1773 0 net=4743
rlabel metal2 86 -1775 86 -1775 0 net=1641
rlabel metal2 86 -1777 86 -1777 0 net=1552
rlabel metal2 149 -1779 149 -1779 0 net=3567
rlabel metal2 142 -1781 142 -1781 0 net=1803
rlabel metal2 37 -1792 37 -1792 0 net=3952
rlabel metal2 541 -1792 541 -1792 0 net=1565
rlabel metal2 695 -1792 695 -1792 0 net=4716
rlabel metal2 947 -1792 947 -1792 0 net=6458
rlabel metal2 1230 -1792 1230 -1792 0 net=11382
rlabel metal2 37 -1794 37 -1794 0 net=5541
rlabel metal2 621 -1794 621 -1794 0 net=5362
rlabel metal2 1143 -1794 1143 -1794 0 net=8063
rlabel metal2 1395 -1794 1395 -1794 0 net=9530
rlabel metal2 30 -1796 30 -1796 0 net=4293
rlabel metal2 635 -1796 635 -1796 0 net=4376
rlabel metal2 656 -1796 656 -1796 0 net=2760
rlabel metal2 898 -1796 898 -1796 0 net=8152
rlabel metal2 1423 -1796 1423 -1796 0 net=10091
rlabel metal2 1451 -1796 1451 -1796 0 net=10267
rlabel metal2 1451 -1796 1451 -1796 0 net=10267
rlabel metal2 1563 -1796 1563 -1796 0 net=11133
rlabel metal2 1563 -1796 1563 -1796 0 net=11133
rlabel metal2 1640 -1796 1640 -1796 0 net=12711
rlabel metal2 30 -1798 30 -1798 0 net=3257
rlabel metal2 100 -1798 100 -1798 0 net=3182
rlabel metal2 142 -1798 142 -1798 0 net=1773
rlabel metal2 1192 -1798 1192 -1798 0 net=8947
rlabel metal2 1423 -1798 1423 -1798 0 net=10953
rlabel metal2 65 -1800 65 -1800 0 net=3582
rlabel metal2 268 -1800 268 -1800 0 net=4739
rlabel metal2 674 -1800 674 -1800 0 net=4811
rlabel metal2 716 -1800 716 -1800 0 net=8290
rlabel metal2 68 -1802 68 -1802 0 net=4720
rlabel metal2 387 -1802 387 -1802 0 net=2603
rlabel metal2 387 -1802 387 -1802 0 net=2603
rlabel metal2 394 -1802 394 -1802 0 net=4154
rlabel metal2 548 -1802 548 -1802 0 net=7944
rlabel metal2 1213 -1802 1213 -1802 0 net=8681
rlabel metal2 1325 -1802 1325 -1802 0 net=10677
rlabel metal2 72 -1804 72 -1804 0 net=1642
rlabel metal2 145 -1804 145 -1804 0 net=1118
rlabel metal2 373 -1804 373 -1804 0 net=4745
rlabel metal2 723 -1804 723 -1804 0 net=382
rlabel metal2 1024 -1804 1024 -1804 0 net=11796
rlabel metal2 72 -1806 72 -1806 0 net=4621
rlabel metal2 499 -1806 499 -1806 0 net=7062
rlabel metal2 1178 -1806 1178 -1806 0 net=8369
rlabel metal2 1234 -1806 1234 -1806 0 net=11095
rlabel metal2 1689 -1806 1689 -1806 0 net=12469
rlabel metal2 75 -1808 75 -1808 0 net=5248
rlabel metal2 821 -1808 821 -1808 0 net=5826
rlabel metal2 884 -1808 884 -1808 0 net=11570
rlabel metal2 79 -1810 79 -1810 0 net=5807
rlabel metal2 89 -1810 89 -1810 0 net=1804
rlabel metal2 184 -1810 184 -1810 0 net=2372
rlabel metal2 250 -1810 250 -1810 0 net=3081
rlabel metal2 548 -1810 548 -1810 0 net=3983
rlabel metal2 674 -1810 674 -1810 0 net=5067
rlabel metal2 782 -1810 782 -1810 0 net=12320
rlabel metal2 58 -1812 58 -1812 0 net=1505
rlabel metal2 184 -1812 184 -1812 0 net=2079
rlabel metal2 338 -1812 338 -1812 0 net=2832
rlabel metal2 576 -1812 576 -1812 0 net=3933
rlabel metal2 677 -1812 677 -1812 0 net=6802
rlabel metal2 1101 -1812 1101 -1812 0 net=7897
rlabel metal2 1283 -1812 1283 -1812 0 net=8999
rlabel metal2 1444 -1812 1444 -1812 0 net=11995
rlabel metal2 1794 -1812 1794 -1812 0 net=10189
rlabel metal2 58 -1814 58 -1814 0 net=11560
rlabel metal2 1668 -1814 1668 -1814 0 net=12155
rlabel metal2 79 -1816 79 -1816 0 net=5605
rlabel metal2 583 -1816 583 -1816 0 net=4110
rlabel metal2 726 -1816 726 -1816 0 net=200
rlabel metal2 1332 -1816 1332 -1816 0 net=9525
rlabel metal2 1661 -1816 1661 -1816 0 net=12107
rlabel metal2 1745 -1816 1745 -1816 0 net=12601
rlabel metal2 93 -1818 93 -1818 0 net=4027
rlabel metal2 534 -1818 534 -1818 0 net=4091
rlabel metal2 597 -1818 597 -1818 0 net=6505
rlabel metal2 786 -1818 786 -1818 0 net=7414
rlabel metal2 1381 -1818 1381 -1818 0 net=12540
rlabel metal2 100 -1820 100 -1820 0 net=1995
rlabel metal2 422 -1820 422 -1820 0 net=5042
rlabel metal2 726 -1820 726 -1820 0 net=522
rlabel metal2 1052 -1820 1052 -1820 0 net=7863
rlabel metal2 1374 -1820 1374 -1820 0 net=9811
rlabel metal2 1577 -1820 1577 -1820 0 net=8891
rlabel metal2 110 -1822 110 -1822 0 net=8711
rlabel metal2 1416 -1822 1416 -1822 0 net=11201
rlabel metal2 128 -1824 128 -1824 0 net=3569
rlabel metal2 159 -1824 159 -1824 0 net=252
rlabel metal2 149 -1826 149 -1826 0 net=3357
rlabel metal2 527 -1826 527 -1826 0 net=3553
rlabel metal2 730 -1826 730 -1826 0 net=5177
rlabel metal2 765 -1826 765 -1826 0 net=5000
rlabel metal2 891 -1826 891 -1826 0 net=5835
rlabel metal2 975 -1826 975 -1826 0 net=8582
rlabel metal2 1293 -1826 1293 -1826 0 net=11663
rlabel metal2 170 -1828 170 -1828 0 net=5064
rlabel metal2 1150 -1828 1150 -1828 0 net=7875
rlabel metal2 1269 -1828 1269 -1828 0 net=10317
rlabel metal2 1577 -1828 1577 -1828 0 net=11353
rlabel metal2 471 -1830 471 -1830 0 net=4501
rlabel metal2 733 -1830 733 -1830 0 net=5292
rlabel metal2 831 -1830 831 -1830 0 net=12232
rlabel metal2 114 -1832 114 -1832 0 net=2419
rlabel metal2 856 -1832 856 -1832 0 net=6101
rlabel metal2 898 -1832 898 -1832 0 net=5783
rlabel metal2 947 -1832 947 -1832 0 net=6383
rlabel metal2 1426 -1832 1426 -1832 0 net=1
rlabel metal2 219 -1834 219 -1834 0 net=2866
rlabel metal2 341 -1834 341 -1834 0 net=1816
rlabel metal2 1290 -1834 1290 -1834 0 net=11695
rlabel metal2 135 -1836 135 -1836 0 net=2449
rlabel metal2 352 -1836 352 -1836 0 net=2351
rlabel metal2 352 -1836 352 -1836 0 net=2351
rlabel metal2 359 -1836 359 -1836 0 net=3869
rlabel metal2 758 -1836 758 -1836 0 net=5131
rlabel metal2 810 -1836 810 -1836 0 net=8562
rlabel metal2 1458 -1836 1458 -1836 0 net=10371
rlabel metal2 135 -1838 135 -1838 0 net=1921
rlabel metal2 222 -1838 222 -1838 0 net=4923
rlabel metal2 765 -1838 765 -1838 0 net=6849
rlabel metal2 1066 -1838 1066 -1838 0 net=7339
rlabel metal2 1311 -1838 1311 -1838 0 net=9303
rlabel metal2 1465 -1838 1465 -1838 0 net=10427
rlabel metal2 163 -1840 163 -1840 0 net=2337
rlabel metal2 222 -1840 222 -1840 0 net=11154
rlabel metal2 191 -1842 191 -1842 0 net=7155
rlabel metal2 261 -1842 261 -1842 0 net=8193
rlabel metal2 527 -1842 527 -1842 0 net=8621
rlabel metal2 1353 -1842 1353 -1842 0 net=9763
rlabel metal2 1430 -1842 1430 -1842 0 net=10465
rlabel metal2 1570 -1842 1570 -1842 0 net=10213
rlabel metal2 61 -1844 61 -1844 0 net=2867
rlabel metal2 268 -1844 268 -1844 0 net=3223
rlabel metal2 544 -1844 544 -1844 0 net=9749
rlabel metal2 1297 -1844 1297 -1844 0 net=8845
rlabel metal2 1570 -1844 1570 -1844 0 net=12617
rlabel metal2 173 -1846 173 -1846 0 net=10019
rlabel metal2 226 -1848 226 -1848 0 net=1862
rlabel metal2 415 -1848 415 -1848 0 net=2217
rlabel metal2 786 -1848 786 -1848 0 net=11386
rlabel metal2 23 -1850 23 -1850 0 net=3214
rlabel metal2 793 -1850 793 -1850 0 net=5407
rlabel metal2 856 -1850 856 -1850 0 net=5875
rlabel metal2 1157 -1850 1157 -1850 0 net=11974
rlabel metal2 226 -1852 226 -1852 0 net=1078
rlabel metal2 814 -1852 814 -1852 0 net=5507
rlabel metal2 901 -1852 901 -1852 0 net=11556
rlabel metal2 233 -1854 233 -1854 0 net=2918
rlabel metal2 303 -1854 303 -1854 0 net=1638
rlabel metal2 394 -1854 394 -1854 0 net=2651
rlabel metal2 821 -1854 821 -1854 0 net=7837
rlabel metal2 1297 -1854 1297 -1854 0 net=9233
rlabel metal2 1605 -1854 1605 -1854 0 net=11205
rlabel metal2 44 -1856 44 -1856 0 net=6714
rlabel metal2 824 -1856 824 -1856 0 net=7533
rlabel metal2 1080 -1856 1080 -1856 0 net=7047
rlabel metal2 1605 -1856 1605 -1856 0 net=12223
rlabel metal2 44 -1858 44 -1858 0 net=4975
rlabel metal2 842 -1858 842 -1858 0 net=5705
rlabel metal2 919 -1858 919 -1858 0 net=6147
rlabel metal2 975 -1858 975 -1858 0 net=6609
rlabel metal2 1024 -1858 1024 -1858 0 net=9769
rlabel metal2 1647 -1858 1647 -1858 0 net=11985
rlabel metal2 219 -1860 219 -1860 0 net=1883
rlabel metal2 317 -1860 317 -1860 0 net=3491
rlabel metal2 562 -1860 562 -1860 0 net=5259
rlabel metal2 870 -1860 870 -1860 0 net=7807
rlabel metal2 1094 -1860 1094 -1860 0 net=11332
rlabel metal2 1654 -1860 1654 -1860 0 net=11945
rlabel metal2 1710 -1860 1710 -1860 0 net=12279
rlabel metal2 198 -1862 198 -1862 0 net=5901
rlabel metal2 632 -1862 632 -1862 0 net=4273
rlabel metal2 702 -1862 702 -1862 0 net=5219
rlabel metal2 800 -1862 800 -1862 0 net=5425
rlabel metal2 877 -1862 877 -1862 0 net=6653
rlabel metal2 1017 -1862 1017 -1862 0 net=6909
rlabel metal2 1080 -1862 1080 -1862 0 net=7603
rlabel metal2 1346 -1862 1346 -1862 0 net=7851
rlabel metal2 86 -1864 86 -1864 0 net=7547
rlabel metal2 1409 -1864 1409 -1864 0 net=10229
rlabel metal2 1626 -1864 1626 -1864 0 net=11841
rlabel metal2 1703 -1864 1703 -1864 0 net=12187
rlabel metal2 86 -1866 86 -1866 0 net=5583
rlabel metal2 422 -1866 422 -1866 0 net=2381
rlabel metal2 471 -1866 471 -1866 0 net=3153
rlabel metal2 1045 -1866 1045 -1866 0 net=8653
rlabel metal2 1437 -1866 1437 -1866 0 net=10871
rlabel metal2 1591 -1866 1591 -1866 0 net=10081
rlabel metal2 156 -1868 156 -1868 0 net=9729
rlabel metal2 1521 -1868 1521 -1868 0 net=10987
rlabel metal2 1591 -1868 1591 -1868 0 net=11291
rlabel metal2 1633 -1868 1633 -1868 0 net=11717
rlabel metal2 156 -1870 156 -1870 0 net=3435
rlabel metal2 254 -1870 254 -1870 0 net=2811
rlabel metal2 849 -1870 849 -1870 0 net=7986
rlabel metal2 1542 -1870 1542 -1870 0 net=11053
rlabel metal2 1612 -1870 1612 -1870 0 net=11775
rlabel metal2 198 -1872 198 -1872 0 net=2937
rlabel metal2 366 -1872 366 -1872 0 net=5431
rlabel metal2 877 -1872 877 -1872 0 net=8113
rlabel metal2 1045 -1872 1045 -1872 0 net=8051
rlabel metal2 1304 -1872 1304 -1872 0 net=9251
rlabel metal2 1549 -1872 1549 -1872 0 net=11089
rlabel metal2 1633 -1872 1633 -1872 0 net=11879
rlabel metal2 240 -1874 240 -1874 0 net=2189
rlabel metal2 296 -1874 296 -1874 0 net=2767
rlabel metal2 429 -1874 429 -1874 0 net=4883
rlabel metal2 905 -1874 905 -1874 0 net=2809
rlabel metal2 1171 -1874 1171 -1874 0 net=8221
rlabel metal2 1318 -1874 1318 -1874 0 net=9485
rlabel metal2 1675 -1874 1675 -1874 0 net=12015
rlabel metal2 275 -1876 275 -1876 0 net=2985
rlabel metal2 618 -1876 618 -1876 0 net=7621
rlabel metal2 702 -1876 702 -1876 0 net=5973
rlabel metal2 1010 -1876 1010 -1876 0 net=6765
rlabel metal2 1360 -1876 1360 -1876 0 net=11115
rlabel metal2 1696 -1876 1696 -1876 0 net=12167
rlabel metal2 275 -1878 275 -1878 0 net=4353
rlabel metal2 688 -1878 688 -1878 0 net=6501
rlabel metal2 1360 -1878 1360 -1878 0 net=9757
rlabel metal2 1731 -1878 1731 -1878 0 net=12553
rlabel metal2 282 -1880 282 -1880 0 net=2174
rlabel metal2 366 -1880 366 -1880 0 net=3237
rlabel metal2 618 -1880 618 -1880 0 net=9609
rlabel metal2 1367 -1880 1367 -1880 0 net=10479
rlabel metal2 282 -1882 282 -1882 0 net=1609
rlabel metal2 331 -1882 331 -1882 0 net=3061
rlabel metal2 478 -1882 478 -1882 0 net=3371
rlabel metal2 579 -1882 579 -1882 0 net=9853
rlabel metal2 1479 -1882 1479 -1882 0 net=10705
rlabel metal2 205 -1884 205 -1884 0 net=2497
rlabel metal2 331 -1884 331 -1884 0 net=1729
rlabel metal2 345 -1884 345 -1884 0 net=5135
rlabel metal2 1500 -1884 1500 -1884 0 net=10749
rlabel metal2 205 -1886 205 -1886 0 net=5953
rlabel metal2 954 -1886 954 -1886 0 net=6461
rlabel metal2 1507 -1886 1507 -1886 0 net=10773
rlabel metal2 296 -1888 296 -1888 0 net=2733
rlabel metal2 485 -1888 485 -1888 0 net=4325
rlabel metal2 660 -1888 660 -1888 0 net=4725
rlabel metal2 688 -1888 688 -1888 0 net=6601
rlabel metal2 1514 -1888 1514 -1888 0 net=10925
rlabel metal2 121 -1890 121 -1890 0 net=3978
rlabel metal2 681 -1890 681 -1890 0 net=5522
rlabel metal2 1486 -1890 1486 -1890 0 net=11141
rlabel metal2 121 -1892 121 -1892 0 net=4961
rlabel metal2 779 -1892 779 -1892 0 net=8985
rlabel metal2 380 -1894 380 -1894 0 net=5845
rlabel metal2 401 -1894 401 -1894 0 net=3169
rlabel metal2 492 -1894 492 -1894 0 net=5775
rlabel metal2 933 -1894 933 -1894 0 net=6987
rlabel metal2 1038 -1894 1038 -1894 0 net=7317
rlabel metal2 1129 -1894 1129 -1894 0 net=9317
rlabel metal2 401 -1896 401 -1896 0 net=12489
rlabel metal2 436 -1898 436 -1898 0 net=4105
rlabel metal2 737 -1898 737 -1898 0 net=4989
rlabel metal2 912 -1898 912 -1898 0 net=9875
rlabel metal2 51 -1900 51 -1900 0 net=6722
rlabel metal2 933 -1900 933 -1900 0 net=6169
rlabel metal2 1108 -1900 1108 -1900 0 net=8635
rlabel metal2 51 -1902 51 -1902 0 net=3721
rlabel metal2 436 -1902 436 -1902 0 net=3803
rlabel metal2 751 -1902 751 -1902 0 net=5021
rlabel metal2 940 -1902 940 -1902 0 net=6393
rlabel metal2 1122 -1902 1122 -1902 0 net=9183
rlabel metal2 551 -1904 551 -1904 0 net=6731
rlabel metal2 1129 -1904 1129 -1904 0 net=8215
rlabel metal2 555 -1906 555 -1906 0 net=4043
rlabel metal2 751 -1906 751 -1906 0 net=5857
rlabel metal2 1199 -1906 1199 -1906 0 net=8607
rlabel metal2 513 -1908 513 -1908 0 net=4841
rlabel metal2 926 -1908 926 -1908 0 net=6337
rlabel metal2 1241 -1908 1241 -1908 0 net=8429
rlabel metal2 107 -1910 107 -1910 0 net=3717
rlabel metal2 1185 -1910 1185 -1910 0 net=8781
rlabel metal2 107 -1912 107 -1912 0 net=5470
rlabel metal2 1185 -1912 1185 -1912 0 net=8551
rlabel metal2 233 -1914 233 -1914 0 net=4755
rlabel metal2 1248 -1914 1248 -1914 0 net=8931
rlabel metal2 590 -1916 590 -1916 0 net=10093
rlabel metal2 590 -1918 590 -1918 0 net=6661
rlabel metal2 863 -1920 863 -1920 0 net=3147
rlabel metal2 23 -1931 23 -1931 0 net=6803
rlabel metal2 950 -1931 950 -1931 0 net=7048
rlabel metal2 1143 -1931 1143 -1931 0 net=8065
rlabel metal2 1143 -1931 1143 -1931 0 net=8065
rlabel metal2 1157 -1931 1157 -1931 0 net=7852
rlabel metal2 30 -1933 30 -1933 0 net=3258
rlabel metal2 65 -1933 65 -1933 0 net=5902
rlabel metal2 534 -1933 534 -1933 0 net=3554
rlabel metal2 618 -1933 618 -1933 0 net=9750
rlabel metal2 1297 -1933 1297 -1933 0 net=9235
rlabel metal2 1297 -1933 1297 -1933 0 net=9235
rlabel metal2 1304 -1933 1304 -1933 0 net=9253
rlabel metal2 1304 -1933 1304 -1933 0 net=9253
rlabel metal2 1318 -1933 1318 -1933 0 net=9487
rlabel metal2 1318 -1933 1318 -1933 0 net=9487
rlabel metal2 1381 -1933 1381 -1933 0 net=12016
rlabel metal2 1738 -1933 1738 -1933 0 net=8893
rlabel metal2 37 -1935 37 -1935 0 net=5542
rlabel metal2 219 -1935 219 -1935 0 net=2652
rlabel metal2 408 -1935 408 -1935 0 net=2768
rlabel metal2 656 -1935 656 -1935 0 net=11206
rlabel metal2 37 -1937 37 -1937 0 net=5585
rlabel metal2 93 -1937 93 -1937 0 net=4028
rlabel metal2 772 -1937 772 -1937 0 net=6170
rlabel metal2 968 -1937 968 -1937 0 net=6655
rlabel metal2 968 -1937 968 -1937 0 net=6655
rlabel metal2 985 -1937 985 -1937 0 net=9758
rlabel metal2 1381 -1937 1381 -1937 0 net=9877
rlabel metal2 1619 -1937 1619 -1937 0 net=11697
rlabel metal2 1619 -1937 1619 -1937 0 net=11697
rlabel metal2 1626 -1937 1626 -1937 0 net=11843
rlabel metal2 1626 -1937 1626 -1937 0 net=11843
rlabel metal2 1633 -1937 1633 -1937 0 net=11881
rlabel metal2 1633 -1937 1633 -1937 0 net=11881
rlabel metal2 1640 -1937 1640 -1937 0 net=12713
rlabel metal2 58 -1939 58 -1939 0 net=4107
rlabel metal2 716 -1939 716 -1939 0 net=4924
rlabel metal2 849 -1939 849 -1939 0 net=5785
rlabel metal2 912 -1939 912 -1939 0 net=11292
rlabel metal2 1640 -1939 1640 -1939 0 net=11947
rlabel metal2 1675 -1939 1675 -1939 0 net=12281
rlabel metal2 1717 -1939 1717 -1939 0 net=12603
rlabel metal2 68 -1941 68 -1941 0 net=12470
rlabel metal2 1710 -1941 1710 -1941 0 net=12491
rlabel metal2 79 -1943 79 -1943 0 net=5607
rlabel metal2 100 -1943 100 -1943 0 net=1997
rlabel metal2 583 -1943 583 -1943 0 net=4093
rlabel metal2 583 -1943 583 -1943 0 net=4093
rlabel metal2 604 -1943 604 -1943 0 net=1443
rlabel metal2 716 -1943 716 -1943 0 net=5179
rlabel metal2 744 -1943 744 -1943 0 net=5221
rlabel metal2 744 -1943 744 -1943 0 net=5221
rlabel metal2 754 -1943 754 -1943 0 net=7838
rlabel metal2 873 -1943 873 -1943 0 net=8636
rlabel metal2 1122 -1943 1122 -1943 0 net=11096
rlabel metal2 1500 -1943 1500 -1943 0 net=10751
rlabel metal2 79 -1945 79 -1945 0 net=1923
rlabel metal2 138 -1945 138 -1945 0 net=7622
rlabel metal2 646 -1945 646 -1945 0 net=4741
rlabel metal2 723 -1945 723 -1945 0 net=3849
rlabel metal2 989 -1945 989 -1945 0 net=10480
rlabel metal2 1384 -1945 1384 -1945 0 net=11142
rlabel metal2 1549 -1945 1549 -1945 0 net=11091
rlabel metal2 1654 -1945 1654 -1945 0 net=12109
rlabel metal2 1682 -1945 1682 -1945 0 net=10082
rlabel metal2 100 -1947 100 -1947 0 net=1775
rlabel metal2 149 -1947 149 -1947 0 net=3358
rlabel metal2 912 -1947 912 -1947 0 net=6463
rlabel metal2 1059 -1947 1059 -1947 0 net=7535
rlabel metal2 107 -1949 107 -1949 0 net=3492
rlabel metal2 359 -1949 359 -1949 0 net=3870
rlabel metal2 884 -1949 884 -1949 0 net=6103
rlabel metal2 884 -1949 884 -1949 0 net=6103
rlabel metal2 898 -1949 898 -1949 0 net=6395
rlabel metal2 947 -1949 947 -1949 0 net=6385
rlabel metal2 1080 -1949 1080 -1949 0 net=7605
rlabel metal2 1157 -1949 1157 -1949 0 net=8223
rlabel metal2 1185 -1949 1185 -1949 0 net=8553
rlabel metal2 1199 -1949 1199 -1949 0 net=8609
rlabel metal2 1199 -1949 1199 -1949 0 net=8609
rlabel metal2 1227 -1949 1227 -1949 0 net=11202
rlabel metal2 1423 -1949 1423 -1949 0 net=10955
rlabel metal2 1528 -1949 1528 -1949 0 net=11143
rlabel metal2 135 -1951 135 -1951 0 net=8986
rlabel metal2 1234 -1951 1234 -1951 0 net=8713
rlabel metal2 1234 -1951 1234 -1951 0 net=8713
rlabel metal2 1269 -1951 1269 -1951 0 net=10319
rlabel metal2 1269 -1951 1269 -1951 0 net=10319
rlabel metal2 1290 -1951 1290 -1951 0 net=10467
rlabel metal2 1570 -1951 1570 -1951 0 net=12619
rlabel metal2 142 -1953 142 -1953 0 net=1567
rlabel metal2 597 -1953 597 -1953 0 net=6507
rlabel metal2 1066 -1953 1066 -1953 0 net=7341
rlabel metal2 1087 -1953 1087 -1953 0 net=7809
rlabel metal2 1160 -1953 1160 -1953 0 net=11718
rlabel metal2 149 -1955 149 -1955 0 net=2339
rlabel metal2 166 -1955 166 -1955 0 net=4884
rlabel metal2 730 -1955 730 -1955 0 net=4819
rlabel metal2 1097 -1955 1097 -1955 0 net=10872
rlabel metal2 1661 -1955 1661 -1955 0 net=12157
rlabel metal2 1682 -1955 1682 -1955 0 net=12373
rlabel metal2 1759 -1955 1759 -1955 0 net=10190
rlabel metal2 65 -1957 65 -1957 0 net=4805
rlabel metal2 170 -1957 170 -1957 0 net=2219
rlabel metal2 432 -1957 432 -1957 0 net=7869
rlabel metal2 1167 -1957 1167 -1957 0 net=11986
rlabel metal2 1668 -1957 1668 -1957 0 net=12189
rlabel metal2 159 -1959 159 -1959 0 net=2352
rlabel metal2 359 -1959 359 -1959 0 net=1715
rlabel metal2 639 -1959 639 -1959 0 net=6149
rlabel metal2 929 -1959 929 -1959 0 net=11489
rlabel metal2 1696 -1959 1696 -1959 0 net=12169
rlabel metal2 72 -1961 72 -1961 0 net=4623
rlabel metal2 380 -1961 380 -1961 0 net=5846
rlabel metal2 646 -1961 646 -1961 0 net=4727
rlabel metal2 670 -1961 670 -1961 0 net=12425
rlabel metal2 72 -1963 72 -1963 0 net=6423
rlabel metal2 219 -1963 219 -1963 0 net=4747
rlabel metal2 394 -1963 394 -1963 0 net=3805
rlabel metal2 471 -1963 471 -1963 0 net=3155
rlabel metal2 621 -1963 621 -1963 0 net=10092
rlabel metal2 51 -1965 51 -1965 0 net=3723
rlabel metal2 492 -1965 492 -1965 0 net=5776
rlabel metal2 660 -1965 660 -1965 0 net=7876
rlabel metal2 1171 -1965 1171 -1965 0 net=8371
rlabel metal2 1185 -1965 1185 -1965 0 net=8783
rlabel metal2 1325 -1965 1325 -1965 0 net=10679
rlabel metal2 51 -1967 51 -1967 0 net=5137
rlabel metal2 373 -1967 373 -1967 0 net=5277
rlabel metal2 821 -1967 821 -1967 0 net=5877
rlabel metal2 877 -1967 877 -1967 0 net=8115
rlabel metal2 1178 -1967 1178 -1967 0 net=11135
rlabel metal2 117 -1969 117 -1969 0 net=3381
rlabel metal2 450 -1969 450 -1969 0 net=3063
rlabel metal2 506 -1969 506 -1969 0 net=4843
rlabel metal2 593 -1969 593 -1969 0 net=10105
rlabel metal2 1444 -1969 1444 -1969 0 net=11997
rlabel metal2 226 -1971 226 -1971 0 net=2498
rlabel metal2 324 -1971 324 -1971 0 net=2451
rlabel metal2 401 -1971 401 -1971 0 net=7173
rlabel metal2 1101 -1971 1101 -1971 0 net=7899
rlabel metal2 1444 -1971 1444 -1971 0 net=10429
rlabel metal2 1514 -1971 1514 -1971 0 net=10927
rlabel metal2 177 -1973 177 -1973 0 net=1507
rlabel metal2 240 -1973 240 -1973 0 net=1301
rlabel metal2 345 -1973 345 -1973 0 net=3719
rlabel metal2 555 -1973 555 -1973 0 net=4045
rlabel metal2 670 -1973 670 -1973 0 net=2810
rlabel metal2 915 -1973 915 -1973 0 net=8932
rlabel metal2 1353 -1973 1353 -1973 0 net=9765
rlabel metal2 156 -1975 156 -1975 0 net=3437
rlabel metal2 691 -1975 691 -1975 0 net=9531
rlabel metal2 156 -1977 156 -1977 0 net=488
rlabel metal2 765 -1977 765 -1977 0 net=6851
rlabel metal2 177 -1979 177 -1979 0 net=4209
rlabel metal2 1024 -1979 1024 -1979 0 net=9771
rlabel metal2 1360 -1979 1360 -1979 0 net=9813
rlabel metal2 1388 -1979 1388 -1979 0 net=9855
rlabel metal2 184 -1981 184 -1981 0 net=2081
rlabel metal2 401 -1981 401 -1981 0 net=2647
rlabel metal2 695 -1981 695 -1981 0 net=4813
rlabel metal2 765 -1981 765 -1981 0 net=10615
rlabel metal2 1073 -1981 1073 -1981 0 net=7549
rlabel metal2 1115 -1981 1115 -1981 0 net=8655
rlabel metal2 1230 -1981 1230 -1981 0 net=8969
rlabel metal2 1367 -1981 1367 -1981 0 net=10269
rlabel metal2 184 -1983 184 -1983 0 net=5433
rlabel metal2 856 -1983 856 -1983 0 net=8623
rlabel metal2 1213 -1983 1213 -1983 0 net=8683
rlabel metal2 1374 -1983 1374 -1983 0 net=10707
rlabel metal2 205 -1985 205 -1985 0 net=5955
rlabel metal2 905 -1985 905 -1985 0 net=11776
rlabel metal2 205 -1987 205 -1987 0 net=515
rlabel metal2 233 -1987 233 -1987 0 net=4757
rlabel metal2 702 -1987 702 -1987 0 net=5975
rlabel metal2 940 -1987 940 -1987 0 net=6611
rlabel metal2 1038 -1987 1038 -1987 0 net=7319
rlabel metal2 1087 -1987 1087 -1987 0 net=7651
rlabel metal2 1192 -1987 1192 -1987 0 net=8949
rlabel metal2 1388 -1987 1388 -1987 0 net=10021
rlabel metal2 1409 -1987 1409 -1987 0 net=10231
rlabel metal2 1584 -1987 1584 -1987 0 net=11665
rlabel metal2 233 -1989 233 -1989 0 net=3677
rlabel metal2 702 -1989 702 -1989 0 net=6663
rlabel metal2 1017 -1989 1017 -1989 0 net=6911
rlabel metal2 1213 -1989 1213 -1989 0 net=9611
rlabel metal2 1402 -1989 1402 -1989 0 net=11055
rlabel metal2 240 -1991 240 -1991 0 net=2605
rlabel metal2 408 -1991 408 -1991 0 net=5999
rlabel metal2 688 -1991 688 -1991 0 net=6603
rlabel metal2 1017 -1991 1017 -1991 0 net=9000
rlabel metal2 1409 -1991 1409 -1991 0 net=10373
rlabel metal2 1542 -1991 1542 -1991 0 net=12225
rlabel metal2 247 -1993 247 -1993 0 net=3011
rlabel metal2 324 -1993 324 -1993 0 net=5069
rlabel metal2 772 -1993 772 -1993 0 net=5707
rlabel metal2 975 -1993 975 -1993 0 net=6733
rlabel metal2 1129 -1993 1129 -1993 0 net=8217
rlabel metal2 1430 -1993 1430 -1993 0 net=8847
rlabel metal2 1598 -1993 1598 -1993 0 net=10215
rlabel metal2 107 -1995 107 -1995 0 net=4731
rlabel metal2 789 -1995 789 -1995 0 net=6689
rlabel metal2 1052 -1995 1052 -1995 0 net=7865
rlabel metal2 1276 -1995 1276 -1995 0 net=9185
rlabel metal2 1332 -1995 1332 -1995 0 net=9527
rlabel metal2 1556 -1995 1556 -1995 0 net=11117
rlabel metal2 243 -1997 243 -1997 0 net=1681
rlabel metal2 250 -1997 250 -1997 0 net=8430
rlabel metal2 1332 -1997 1332 -1997 0 net=9731
rlabel metal2 1556 -1997 1556 -1997 0 net=11355
rlabel metal2 254 -1999 254 -1999 0 net=2813
rlabel metal2 450 -1999 450 -1999 0 net=3287
rlabel metal2 667 -1999 667 -1999 0 net=7063
rlabel metal2 1255 -1999 1255 -1999 0 net=10399
rlabel metal2 1577 -1999 1577 -1999 0 net=12555
rlabel metal2 254 -2001 254 -2001 0 net=2191
rlabel metal2 303 -2001 303 -2001 0 net=1885
rlabel metal2 387 -2001 387 -2001 0 net=3985
rlabel metal2 576 -2001 576 -2001 0 net=3935
rlabel metal2 667 -2001 667 -2001 0 net=9657
rlabel metal2 1346 -2001 1346 -2001 0 net=10775
rlabel metal2 1521 -2001 1521 -2001 0 net=10989
rlabel metal2 268 -2003 268 -2003 0 net=3224
rlabel metal2 800 -2003 800 -2003 0 net=5426
rlabel metal2 1003 -2003 1003 -2003 0 net=6767
rlabel metal2 1262 -2003 1262 -2003 0 net=10095
rlabel metal2 198 -2005 198 -2005 0 net=2939
rlabel metal2 275 -2005 275 -2005 0 net=4354
rlabel metal2 548 -2005 548 -2005 0 net=4097
rlabel metal2 800 -2005 800 -2005 0 net=6031
rlabel metal2 1010 -2005 1010 -2005 0 net=6797
rlabel metal2 1311 -2005 1311 -2005 0 net=9305
rlabel metal2 110 -2007 110 -2007 0 net=1561
rlabel metal2 282 -2007 282 -2007 0 net=1610
rlabel metal2 457 -2007 457 -2007 0 net=3083
rlabel metal2 590 -2007 590 -2007 0 net=11653
rlabel metal2 114 -2009 114 -2009 0 net=2421
rlabel metal2 229 -2009 229 -2009 0 net=9435
rlabel metal2 114 -2011 114 -2011 0 net=9161
rlabel metal2 282 -2013 282 -2013 0 net=5103
rlabel metal2 807 -2013 807 -2013 0 net=6487
rlabel metal2 1045 -2013 1045 -2013 0 net=8053
rlabel metal2 289 -2015 289 -2015 0 net=2641
rlabel metal2 457 -2015 457 -2015 0 net=4503
rlabel metal2 793 -2015 793 -2015 0 net=5409
rlabel metal2 810 -2015 810 -2015 0 net=11301
rlabel metal2 303 -2017 303 -2017 0 net=1731
rlabel metal2 404 -2017 404 -2017 0 net=6967
rlabel metal2 1164 -2017 1164 -2017 0 net=8245
rlabel metal2 331 -2019 331 -2019 0 net=3239
rlabel metal2 429 -2019 429 -2019 0 net=4295
rlabel metal2 625 -2019 625 -2019 0 net=3149
rlabel metal2 485 -2021 485 -2021 0 net=4327
rlabel metal2 814 -2021 814 -2021 0 net=5509
rlabel metal2 863 -2021 863 -2021 0 net=5837
rlabel metal2 443 -2023 443 -2023 0 net=4587
rlabel metal2 499 -2023 499 -2023 0 net=8195
rlabel metal2 422 -2025 422 -2025 0 net=2383
rlabel metal2 478 -2025 478 -2025 0 net=3373
rlabel metal2 530 -2025 530 -2025 0 net=6387
rlabel metal2 562 -2025 562 -2025 0 net=5261
rlabel metal2 814 -2025 814 -2025 0 net=9318
rlabel metal2 44 -2027 44 -2027 0 net=4977
rlabel metal2 562 -2027 562 -2027 0 net=6503
rlabel metal2 1125 -2027 1125 -2027 0 net=10791
rlabel metal2 44 -2029 44 -2029 0 net=3571
rlabel metal2 212 -2029 212 -2029 0 net=5809
rlabel metal2 590 -2029 590 -2029 0 net=5132
rlabel metal2 891 -2029 891 -2029 0 net=6339
rlabel metal2 961 -2029 961 -2029 0 net=6989
rlabel metal2 128 -2031 128 -2031 0 net=7156
rlabel metal2 212 -2031 212 -2031 0 net=2869
rlabel metal2 737 -2031 737 -2031 0 net=4990
rlabel metal2 121 -2033 121 -2033 0 net=4963
rlabel metal2 758 -2033 758 -2033 0 net=5023
rlabel metal2 828 -2033 828 -2033 0 net=6875
rlabel metal2 121 -2035 121 -2035 0 net=4785
rlabel metal2 173 -2037 173 -2037 0 net=7363
rlabel metal2 191 -2039 191 -2039 0 net=2735
rlabel metal2 786 -2039 786 -2039 0 net=5933
rlabel metal2 261 -2041 261 -2041 0 net=2987
rlabel metal2 751 -2041 751 -2041 0 net=5859
rlabel metal2 296 -2043 296 -2043 0 net=3171
rlabel metal2 520 -2043 520 -2043 0 net=4657
rlabel metal2 751 -2043 751 -2043 0 net=10481
rlabel metal2 464 -2045 464 -2045 0 net=4275
rlabel metal2 86 -2047 86 -2047 0 net=4441
rlabel metal2 40 -2058 40 -2058 0 net=9766
rlabel metal2 1626 -2058 1626 -2058 0 net=11845
rlabel metal2 1661 -2058 1661 -2058 0 net=12159
rlabel metal2 1661 -2058 1661 -2058 0 net=12159
rlabel metal2 1675 -2058 1675 -2058 0 net=12283
rlabel metal2 1675 -2058 1675 -2058 0 net=12283
rlabel metal2 1738 -2058 1738 -2058 0 net=12715
rlabel metal2 1738 -2058 1738 -2058 0 net=12715
rlabel metal2 1759 -2058 1759 -2058 0 net=7537
rlabel metal2 44 -2060 44 -2060 0 net=3572
rlabel metal2 163 -2060 163 -2060 0 net=6504
rlabel metal2 611 -2060 611 -2060 0 net=4329
rlabel metal2 611 -2060 611 -2060 0 net=4329
rlabel metal2 632 -2060 632 -2060 0 net=9306
rlabel metal2 1626 -2060 1626 -2060 0 net=12111
rlabel metal2 1766 -2060 1766 -2060 0 net=8895
rlabel metal2 23 -2062 23 -2062 0 net=6805
rlabel metal2 663 -2062 663 -2062 0 net=5180
rlabel metal2 726 -2062 726 -2062 0 net=584
rlabel metal2 1066 -2062 1066 -2062 0 net=7175
rlabel metal2 1066 -2062 1066 -2062 0 net=7175
rlabel metal2 1080 -2062 1080 -2062 0 net=7343
rlabel metal2 1080 -2062 1080 -2062 0 net=7343
rlabel metal2 1090 -2062 1090 -2062 0 net=10468
rlabel metal2 1346 -2062 1346 -2062 0 net=10777
rlabel metal2 47 -2064 47 -2064 0 net=4742
rlabel metal2 688 -2064 688 -2064 0 net=4964
rlabel metal2 782 -2064 782 -2064 0 net=11136
rlabel metal2 1206 -2064 1206 -2064 0 net=8196
rlabel metal2 68 -2066 68 -2066 0 net=1569
rlabel metal2 142 -2066 142 -2066 0 net=1568
rlabel metal2 803 -2066 803 -2066 0 net=10928
rlabel metal2 100 -2068 100 -2068 0 net=1776
rlabel metal2 786 -2068 786 -2068 0 net=5861
rlabel metal2 835 -2068 835 -2068 0 net=5957
rlabel metal2 835 -2068 835 -2068 0 net=5957
rlabel metal2 873 -2068 873 -2068 0 net=1084
rlabel metal2 100 -2070 100 -2070 0 net=8625
rlabel metal2 919 -2070 919 -2070 0 net=6489
rlabel metal2 926 -2070 926 -2070 0 net=7900
rlabel metal2 1451 -2070 1451 -2070 0 net=11118
rlabel metal2 107 -2072 107 -2072 0 net=81
rlabel metal2 716 -2072 716 -2072 0 net=5223
rlabel metal2 758 -2072 758 -2072 0 net=5025
rlabel metal2 856 -2072 856 -2072 0 net=6033
rlabel metal2 912 -2072 912 -2072 0 net=6465
rlabel metal2 936 -2072 936 -2072 0 net=12170
rlabel metal2 107 -2074 107 -2074 0 net=3301
rlabel metal2 436 -2074 436 -2074 0 net=3382
rlabel metal2 779 -2074 779 -2074 0 net=5977
rlabel metal2 877 -2074 877 -2074 0 net=6509
rlabel metal2 985 -2074 985 -2074 0 net=11123
rlabel metal2 1703 -2074 1703 -2074 0 net=12493
rlabel metal2 114 -2076 114 -2076 0 net=3172
rlabel metal2 352 -2076 352 -2076 0 net=4625
rlabel metal2 453 -2076 453 -2076 0 net=3374
rlabel metal2 506 -2076 506 -2076 0 net=4845
rlabel metal2 744 -2076 744 -2076 0 net=11092
rlabel metal2 1696 -2076 1696 -2076 0 net=12427
rlabel metal2 54 -2078 54 -2078 0 net=2957
rlabel metal2 128 -2078 128 -2078 0 net=10232
rlabel metal2 1570 -2078 1570 -2078 0 net=11491
rlabel metal2 1682 -2078 1682 -2078 0 net=12375
rlabel metal2 128 -2080 128 -2080 0 net=1562
rlabel metal2 289 -2080 289 -2080 0 net=2643
rlabel metal2 359 -2080 359 -2080 0 net=1716
rlabel metal2 667 -2080 667 -2080 0 net=5410
rlabel metal2 898 -2080 898 -2080 0 net=6397
rlabel metal2 919 -2080 919 -2080 0 net=6613
rlabel metal2 947 -2080 947 -2080 0 net=8218
rlabel metal2 1395 -2080 1395 -2080 0 net=10107
rlabel metal2 1451 -2080 1451 -2080 0 net=11357
rlabel metal2 1605 -2080 1605 -2080 0 net=10217
rlabel metal2 121 -2082 121 -2082 0 net=4787
rlabel metal2 674 -2082 674 -2082 0 net=4732
rlabel metal2 758 -2082 758 -2082 0 net=8054
rlabel metal2 1269 -2082 1269 -2082 0 net=10321
rlabel metal2 1528 -2082 1528 -2082 0 net=11145
rlabel metal2 1605 -2082 1605 -2082 0 net=11667
rlabel metal2 1629 -2082 1629 -2082 0 net=1
rlabel metal2 121 -2084 121 -2084 0 net=2341
rlabel metal2 163 -2084 163 -2084 0 net=5879
rlabel metal2 884 -2084 884 -2084 0 net=6105
rlabel metal2 989 -2084 989 -2084 0 net=6386
rlabel metal2 1104 -2084 1104 -2084 0 net=10752
rlabel metal2 173 -2086 173 -2086 0 net=9856
rlabel metal2 1500 -2086 1500 -2086 0 net=10957
rlabel metal2 1535 -2086 1535 -2086 0 net=11303
rlabel metal2 1612 -2086 1612 -2086 0 net=11883
rlabel metal2 177 -2088 177 -2088 0 net=4210
rlabel metal2 821 -2088 821 -2088 0 net=5511
rlabel metal2 936 -2088 936 -2088 0 net=9787
rlabel metal2 1311 -2088 1311 -2088 0 net=9437
rlabel metal2 1353 -2088 1353 -2088 0 net=9773
rlabel metal2 1402 -2088 1402 -2088 0 net=11057
rlabel metal2 1619 -2088 1619 -2088 0 net=11699
rlabel metal2 177 -2090 177 -2090 0 net=5071
rlabel metal2 331 -2090 331 -2090 0 net=3241
rlabel metal2 534 -2090 534 -2090 0 net=1998
rlabel metal2 989 -2090 989 -2090 0 net=6913
rlabel metal2 1157 -2090 1157 -2090 0 net=8225
rlabel metal2 1199 -2090 1199 -2090 0 net=8611
rlabel metal2 1227 -2090 1227 -2090 0 net=8685
rlabel metal2 1325 -2090 1325 -2090 0 net=9659
rlabel metal2 1402 -2090 1402 -2090 0 net=10431
rlabel metal2 1584 -2090 1584 -2090 0 net=11655
rlabel metal2 51 -2092 51 -2092 0 net=5139
rlabel metal2 555 -2092 555 -2092 0 net=6389
rlabel metal2 1010 -2092 1010 -2092 0 net=6799
rlabel metal2 1073 -2092 1073 -2092 0 net=7321
rlabel metal2 1255 -2092 1255 -2092 0 net=11527
rlabel metal2 184 -2094 184 -2094 0 net=5435
rlabel metal2 950 -2094 950 -2094 0 net=8527
rlabel metal2 1258 -2094 1258 -2094 0 net=10990
rlabel metal2 184 -2096 184 -2096 0 net=5279
rlabel metal2 408 -2096 408 -2096 0 net=6001
rlabel metal2 1017 -2096 1017 -2096 0 net=6877
rlabel metal2 1073 -2096 1073 -2096 0 net=8657
rlabel metal2 1339 -2096 1339 -2096 0 net=10271
rlabel metal2 1423 -2096 1423 -2096 0 net=11999
rlabel metal2 1717 -2096 1717 -2096 0 net=12605
rlabel metal2 191 -2098 191 -2098 0 net=2736
rlabel metal2 674 -2098 674 -2098 0 net=3851
rlabel metal2 817 -2098 817 -2098 0 net=12543
rlabel metal2 142 -2100 142 -2100 0 net=2255
rlabel metal2 1031 -2100 1031 -2100 0 net=6969
rlabel metal2 1118 -2100 1118 -2100 0 net=9449
rlabel metal2 1444 -2100 1444 -2100 0 net=9415
rlabel metal2 191 -2102 191 -2102 0 net=2989
rlabel metal2 289 -2102 289 -2102 0 net=1719
rlabel metal2 1045 -2102 1045 -2102 0 net=7065
rlabel metal2 1129 -2102 1129 -2102 0 net=7867
rlabel metal2 1542 -2102 1542 -2102 0 net=12227
rlabel metal2 205 -2104 205 -2104 0 net=9532
rlabel metal2 1584 -2104 1584 -2104 0 net=12191
rlabel metal2 96 -2106 96 -2106 0 net=12245
rlabel metal2 205 -2108 205 -2108 0 net=2941
rlabel metal2 296 -2108 296 -2108 0 net=1733
rlabel metal2 310 -2108 310 -2108 0 net=3013
rlabel metal2 345 -2108 345 -2108 0 net=3720
rlabel metal2 366 -2108 366 -2108 0 net=9039
rlabel metal2 1374 -2108 1374 -2108 0 net=10709
rlabel metal2 208 -2110 208 -2110 0 net=4647
rlabel metal2 691 -2110 691 -2110 0 net=7479
rlabel metal2 1052 -2110 1052 -2110 0 net=7607
rlabel metal2 1115 -2110 1115 -2110 0 net=7653
rlabel metal2 1157 -2110 1157 -2110 0 net=9613
rlabel metal2 1220 -2110 1220 -2110 0 net=8715
rlabel metal2 1332 -2110 1332 -2110 0 net=9733
rlabel metal2 1507 -2110 1507 -2110 0 net=10097
rlabel metal2 212 -2112 212 -2112 0 net=2871
rlabel metal2 310 -2112 310 -2112 0 net=1887
rlabel metal2 324 -2112 324 -2112 0 net=6179
rlabel metal2 1101 -2112 1101 -2112 0 net=7551
rlabel metal2 1115 -2112 1115 -2112 0 net=10665
rlabel metal2 79 -2114 79 -2114 0 net=1925
rlabel metal2 338 -2114 338 -2114 0 net=2083
rlabel metal2 373 -2114 373 -2114 0 net=3807
rlabel metal2 408 -2114 408 -2114 0 net=4098
rlabel metal2 555 -2114 555 -2114 0 net=4047
rlabel metal2 576 -2114 576 -2114 0 net=3085
rlabel metal2 1171 -2114 1171 -2114 0 net=8373
rlabel metal2 1472 -2114 1472 -2114 0 net=10681
rlabel metal2 79 -2116 79 -2116 0 net=2051
rlabel metal2 156 -2118 156 -2118 0 net=6051
rlabel metal2 422 -2118 422 -2118 0 net=4979
rlabel metal2 1192 -2118 1192 -2118 0 net=8555
rlabel metal2 1234 -2118 1234 -2118 0 net=8971
rlabel metal2 1437 -2118 1437 -2118 0 net=10401
rlabel metal2 1724 -2118 1724 -2118 0 net=12621
rlabel metal2 131 -2120 131 -2120 0 net=2319
rlabel metal2 166 -2120 166 -2120 0 net=4157
rlabel metal2 593 -2120 593 -2120 0 net=9581
rlabel metal2 1409 -2120 1409 -2120 0 net=10375
rlabel metal2 1577 -2120 1577 -2120 0 net=12557
rlabel metal2 212 -2122 212 -2122 0 net=2041
rlabel metal2 905 -2122 905 -2122 0 net=11431
rlabel metal2 233 -2124 233 -2124 0 net=3679
rlabel metal2 541 -2124 541 -2124 0 net=3157
rlabel metal2 569 -2124 569 -2124 0 net=5709
rlabel metal2 1192 -2124 1192 -2124 0 net=9163
rlabel metal2 1388 -2124 1388 -2124 0 net=10023
rlabel metal2 233 -2126 233 -2126 0 net=2193
rlabel metal2 338 -2126 338 -2126 0 net=2815
rlabel metal2 429 -2126 429 -2126 0 net=4297
rlabel metal2 530 -2126 530 -2126 0 net=4763
rlabel metal2 607 -2126 607 -2126 0 net=11025
rlabel metal2 86 -2128 86 -2128 0 net=4443
rlabel metal2 345 -2128 345 -2128 0 net=2141
rlabel metal2 765 -2128 765 -2128 0 net=7495
rlabel metal2 1276 -2128 1276 -2128 0 net=11949
rlabel metal2 37 -2130 37 -2130 0 net=5587
rlabel metal2 772 -2130 772 -2130 0 net=6852
rlabel metal2 86 -2132 86 -2132 0 net=5810
rlabel metal2 485 -2132 485 -2132 0 net=4589
rlabel metal2 618 -2132 618 -2132 0 net=6359
rlabel metal2 1381 -2132 1381 -2132 0 net=9879
rlabel metal2 1479 -2132 1479 -2132 0 net=8849
rlabel metal2 30 -2134 30 -2134 0 net=3601
rlabel metal2 621 -2134 621 -2134 0 net=4728
rlabel metal2 660 -2134 660 -2134 0 net=8833
rlabel metal2 1360 -2134 1360 -2134 0 net=9815
rlabel metal2 1458 -2134 1458 -2134 0 net=10483
rlabel metal2 1486 -2134 1486 -2134 0 net=10793
rlabel metal2 51 -2136 51 -2136 0 net=3587
rlabel metal2 485 -2136 485 -2136 0 net=4821
rlabel metal2 1059 -2136 1059 -2136 0 net=10617
rlabel metal2 240 -2138 240 -2138 0 net=2607
rlabel metal2 387 -2138 387 -2138 0 net=3987
rlabel metal2 429 -2138 429 -2138 0 net=6657
rlabel metal2 1059 -2138 1059 -2138 0 net=7119
rlabel metal2 1318 -2138 1318 -2138 0 net=9489
rlabel metal2 170 -2140 170 -2140 0 net=2221
rlabel metal2 247 -2140 247 -2140 0 net=1683
rlabel metal2 387 -2140 387 -2140 0 net=2385
rlabel metal2 457 -2140 457 -2140 0 net=4505
rlabel metal2 968 -2140 968 -2140 0 net=6769
rlabel metal2 1087 -2140 1087 -2140 0 net=7365
rlabel metal2 1304 -2140 1304 -2140 0 net=9255
rlabel metal2 93 -2142 93 -2142 0 net=5609
rlabel metal2 464 -2142 464 -2142 0 net=4277
rlabel metal2 653 -2142 653 -2142 0 net=3936
rlabel metal2 814 -2142 814 -2142 0 net=7003
rlabel metal2 1094 -2142 1094 -2142 0 net=8067
rlabel metal2 1297 -2142 1297 -2142 0 net=9237
rlabel metal2 93 -2144 93 -2144 0 net=6604
rlabel metal2 1122 -2144 1122 -2144 0 net=7811
rlabel metal2 1283 -2144 1283 -2144 0 net=9187
rlabel metal2 58 -2146 58 -2146 0 net=4108
rlabel metal2 1241 -2146 1241 -2146 0 net=8951
rlabel metal2 58 -2148 58 -2148 0 net=3151
rlabel metal2 670 -2148 670 -2148 0 net=10393
rlabel metal2 170 -2150 170 -2150 0 net=12335
rlabel metal2 219 -2152 219 -2152 0 net=4749
rlabel metal2 471 -2152 471 -2152 0 net=3724
rlabel metal2 1185 -2152 1185 -2152 0 net=8785
rlabel metal2 198 -2154 198 -2154 0 net=2423
rlabel metal2 226 -2154 226 -2154 0 net=1509
rlabel metal2 362 -2154 362 -2154 0 net=3125
rlabel metal2 492 -2154 492 -2154 0 net=3065
rlabel metal2 492 -2154 492 -2154 0 net=3065
rlabel metal2 520 -2154 520 -2154 0 net=4659
rlabel metal2 751 -2154 751 -2154 0 net=7057
rlabel metal2 1164 -2154 1164 -2154 0 net=8247
rlabel metal2 198 -2156 198 -2156 0 net=1751
rlabel metal2 226 -2158 226 -2158 0 net=9528
rlabel metal2 229 -2160 229 -2160 0 net=3855
rlabel metal2 513 -2160 513 -2160 0 net=3438
rlabel metal2 583 -2160 583 -2160 0 net=4095
rlabel metal2 751 -2160 751 -2160 0 net=5935
rlabel metal2 1150 -2160 1150 -2160 0 net=8117
rlabel metal2 65 -2162 65 -2162 0 net=4807
rlabel metal2 583 -2162 583 -2162 0 net=4759
rlabel metal2 1136 -2162 1136 -2162 0 net=7871
rlabel metal2 65 -2164 65 -2164 0 net=6690
rlabel metal2 415 -2166 415 -2166 0 net=5903
rlabel metal2 982 -2166 982 -2166 0 net=7741
rlabel metal2 600 -2168 600 -2168 0 net=10169
rlabel metal2 625 -2170 625 -2170 0 net=6341
rlabel metal2 961 -2170 961 -2170 0 net=6991
rlabel metal2 695 -2172 695 -2172 0 net=4815
rlabel metal2 849 -2172 849 -2172 0 net=5787
rlabel metal2 975 -2172 975 -2172 0 net=6735
rlabel metal2 282 -2174 282 -2174 0 net=5105
rlabel metal2 849 -2174 849 -2174 0 net=5839
rlabel metal2 282 -2176 282 -2176 0 net=2649
rlabel metal2 639 -2176 639 -2176 0 net=6151
rlabel metal2 72 -2178 72 -2178 0 net=6425
rlabel metal2 702 -2178 702 -2178 0 net=6665
rlabel metal2 72 -2180 72 -2180 0 net=6623
rlabel metal2 380 -2182 380 -2182 0 net=2453
rlabel metal2 702 -2182 702 -2182 0 net=5262
rlabel metal2 933 -2182 933 -2182 0 net=9133
rlabel metal2 380 -2184 380 -2184 0 net=3289
rlabel metal2 450 -2186 450 -2186 0 net=6277
rlabel metal2 30 -2197 30 -2197 0 net=3602
rlabel metal2 453 -2197 453 -2197 0 net=4096
rlabel metal2 688 -2197 688 -2197 0 net=3086
rlabel metal2 796 -2197 796 -2197 0 net=9774
rlabel metal2 1437 -2197 1437 -2197 0 net=10377
rlabel metal2 1437 -2197 1437 -2197 0 net=10377
rlabel metal2 1500 -2197 1500 -2197 0 net=10667
rlabel metal2 1500 -2197 1500 -2197 0 net=10667
rlabel metal2 1535 -2197 1535 -2197 0 net=11027
rlabel metal2 1535 -2197 1535 -2197 0 net=11027
rlabel metal2 1570 -2197 1570 -2197 0 net=11305
rlabel metal2 1570 -2197 1570 -2197 0 net=11305
rlabel metal2 1640 -2197 1640 -2197 0 net=10794
rlabel metal2 1752 -2197 1752 -2197 0 net=8896
rlabel metal2 44 -2199 44 -2199 0 net=741
rlabel metal2 873 -2199 873 -2199 0 net=10322
rlabel metal2 1640 -2199 1640 -2199 0 net=12377
rlabel metal2 51 -2201 51 -2201 0 net=6624
rlabel metal2 89 -2201 89 -2201 0 net=1877
rlabel metal2 117 -2201 117 -2201 0 net=9416
rlabel metal2 1465 -2201 1465 -2201 0 net=10711
rlabel metal2 1647 -2201 1647 -2201 0 net=12229
rlabel metal2 1647 -2201 1647 -2201 0 net=12229
rlabel metal2 1682 -2201 1682 -2201 0 net=10218
rlabel metal2 51 -2203 51 -2203 0 net=6053
rlabel metal2 408 -2203 408 -2203 0 net=5979
rlabel metal2 786 -2203 786 -2203 0 net=5026
rlabel metal2 828 -2203 828 -2203 0 net=7868
rlabel metal2 1514 -2203 1514 -2203 0 net=11125
rlabel metal2 1682 -2203 1682 -2203 0 net=12545
rlabel metal2 58 -2205 58 -2205 0 net=3152
rlabel metal2 978 -2205 978 -2205 0 net=12000
rlabel metal2 1549 -2205 1549 -2205 0 net=11493
rlabel metal2 1696 -2205 1696 -2205 0 net=12717
rlabel metal2 58 -2207 58 -2207 0 net=6427
rlabel metal2 691 -2207 691 -2207 0 net=5224
rlabel metal2 723 -2207 723 -2207 0 net=9438
rlabel metal2 1423 -2207 1423 -2207 0 net=10403
rlabel metal2 1738 -2207 1738 -2207 0 net=7539
rlabel metal2 65 -2209 65 -2209 0 net=4569
rlabel metal2 607 -2209 607 -2209 0 net=4980
rlabel metal2 814 -2209 814 -2209 0 net=5513
rlabel metal2 828 -2209 828 -2209 0 net=6003
rlabel metal2 852 -2209 852 -2209 0 net=6970
rlabel metal2 1118 -2209 1118 -2209 0 net=12160
rlabel metal2 68 -2211 68 -2211 0 net=6806
rlabel metal2 590 -2211 590 -2211 0 net=4279
rlabel metal2 590 -2211 590 -2211 0 net=4279
rlabel metal2 611 -2211 611 -2211 0 net=4330
rlabel metal2 758 -2211 758 -2211 0 net=7655
rlabel metal2 1146 -2211 1146 -2211 0 net=12606
rlabel metal2 72 -2213 72 -2213 0 net=2343
rlabel metal2 131 -2213 131 -2213 0 net=6878
rlabel metal2 1031 -2213 1031 -2213 0 net=7543
rlabel metal2 1129 -2213 1129 -2213 0 net=8613
rlabel metal2 1227 -2213 1227 -2213 0 net=7323
rlabel metal2 89 -2215 89 -2215 0 net=5072
rlabel metal2 184 -2215 184 -2215 0 net=5281
rlabel metal2 618 -2215 618 -2215 0 net=10041
rlabel metal2 1507 -2215 1507 -2215 0 net=10683
rlabel metal2 93 -2217 93 -2217 0 net=4506
rlabel metal2 891 -2217 891 -2217 0 net=5788
rlabel metal2 999 -2217 999 -2217 0 net=11950
rlabel metal2 1335 -2217 1335 -2217 0 net=11846
rlabel metal2 96 -2219 96 -2219 0 net=7058
rlabel metal2 1192 -2219 1192 -2219 0 net=9165
rlabel metal2 96 -2221 96 -2221 0 net=4237
rlabel metal2 226 -2221 226 -2221 0 net=5905
rlabel metal2 450 -2221 450 -2221 0 net=4661
rlabel metal2 695 -2221 695 -2221 0 net=4816
rlabel metal2 733 -2221 733 -2221 0 net=12494
rlabel metal2 121 -2223 121 -2223 0 net=2195
rlabel metal2 236 -2223 236 -2223 0 net=8399
rlabel metal2 807 -2223 807 -2223 0 net=5959
rlabel metal2 842 -2223 842 -2223 0 net=6511
rlabel metal2 884 -2223 884 -2223 0 net=7177
rlabel metal2 1122 -2223 1122 -2223 0 net=12622
rlabel metal2 142 -2225 142 -2225 0 net=2257
rlabel metal2 152 -2225 152 -2225 0 net=10445
rlabel metal2 142 -2227 142 -2227 0 net=6343
rlabel metal2 639 -2227 639 -2227 0 net=6800
rlabel metal2 1066 -2227 1066 -2227 0 net=6957
rlabel metal2 170 -2229 170 -2229 0 net=1926
rlabel metal2 362 -2229 362 -2229 0 net=660
rlabel metal2 877 -2229 877 -2229 0 net=6361
rlabel metal2 933 -2229 933 -2229 0 net=8952
rlabel metal2 1346 -2229 1346 -2229 0 net=10433
rlabel metal2 170 -2231 170 -2231 0 net=127
rlabel metal2 569 -2231 569 -2231 0 net=5711
rlabel metal2 702 -2231 702 -2231 0 net=11700
rlabel metal2 177 -2233 177 -2233 0 net=2943
rlabel metal2 229 -2233 229 -2233 0 net=6390
rlabel metal2 999 -2233 999 -2233 0 net=7707
rlabel metal2 205 -2235 205 -2235 0 net=2143
rlabel metal2 464 -2235 464 -2235 0 net=3127
rlabel metal2 618 -2235 618 -2235 0 net=3853
rlabel metal2 702 -2235 702 -2235 0 net=8556
rlabel metal2 1227 -2235 1227 -2235 0 net=9189
rlabel metal2 1339 -2235 1339 -2235 0 net=10273
rlabel metal2 1626 -2235 1626 -2235 0 net=12113
rlabel metal2 100 -2237 100 -2237 0 net=8627
rlabel metal2 716 -2237 716 -2237 0 net=5937
rlabel metal2 772 -2237 772 -2237 0 net=11155
rlabel metal2 1612 -2237 1612 -2237 0 net=11885
rlabel metal2 44 -2239 44 -2239 0 net=8339
rlabel metal2 786 -2239 786 -2239 0 net=5863
rlabel metal2 821 -2239 821 -2239 0 net=5841
rlabel metal2 891 -2239 891 -2239 0 net=7067
rlabel metal2 1206 -2239 1206 -2239 0 net=9257
rlabel metal2 1339 -2239 1339 -2239 0 net=9881
rlabel metal2 1542 -2239 1542 -2239 0 net=10099
rlabel metal2 100 -2241 100 -2241 0 net=1571
rlabel metal2 191 -2241 191 -2241 0 net=2991
rlabel metal2 422 -2241 422 -2241 0 net=3989
rlabel metal2 471 -2241 471 -2241 0 net=3857
rlabel metal2 569 -2241 569 -2241 0 net=7121
rlabel metal2 1213 -2241 1213 -2241 0 net=9041
rlabel metal2 1276 -2241 1276 -2241 0 net=10619
rlabel metal2 1542 -2241 1542 -2241 0 net=11433
rlabel metal2 135 -2243 135 -2243 0 net=11656
rlabel metal2 191 -2245 191 -2245 0 net=2223
rlabel metal2 268 -2245 268 -2245 0 net=4049
rlabel metal2 586 -2245 586 -2245 0 net=8489
rlabel metal2 1237 -2245 1237 -2245 0 net=12284
rlabel metal2 107 -2247 107 -2247 0 net=3303
rlabel metal2 271 -2247 271 -2247 0 net=4764
rlabel metal2 548 -2247 548 -2247 0 net=3159
rlabel metal2 646 -2247 646 -2247 0 net=6279
rlabel metal2 730 -2247 730 -2247 0 net=10875
rlabel metal2 1486 -2247 1486 -2247 0 net=10779
rlabel metal2 1577 -2247 1577 -2247 0 net=11887
rlabel metal2 107 -2249 107 -2249 0 net=5881
rlabel metal2 233 -2249 233 -2249 0 net=1684
rlabel metal2 282 -2249 282 -2249 0 net=2650
rlabel metal2 800 -2249 800 -2249 0 net=6467
rlabel metal2 933 -2249 933 -2249 0 net=6771
rlabel metal2 1003 -2249 1003 -2249 0 net=7005
rlabel metal2 1255 -2249 1255 -2249 0 net=10171
rlabel metal2 1521 -2249 1521 -2249 0 net=12559
rlabel metal2 114 -2251 114 -2251 0 net=2959
rlabel metal2 282 -2251 282 -2251 0 net=4627
rlabel metal2 506 -2251 506 -2251 0 net=3242
rlabel metal2 737 -2251 737 -2251 0 net=5437
rlabel metal2 835 -2251 835 -2251 0 net=6667
rlabel metal2 1003 -2251 1003 -2251 0 net=7873
rlabel metal2 1283 -2251 1283 -2251 0 net=10109
rlabel metal2 163 -2253 163 -2253 0 net=4649
rlabel metal2 656 -2253 656 -2253 0 net=6445
rlabel metal2 747 -2253 747 -2253 0 net=12641
rlabel metal2 215 -2255 215 -2255 0 net=5911
rlabel metal2 751 -2255 751 -2255 0 net=6035
rlabel metal2 898 -2255 898 -2255 0 net=7481
rlabel metal2 1010 -2255 1010 -2255 0 net=9490
rlabel metal2 1388 -2255 1388 -2255 0 net=11529
rlabel metal2 156 -2257 156 -2257 0 net=2320
rlabel metal2 905 -2257 905 -2257 0 net=6615
rlabel metal2 926 -2257 926 -2257 0 net=6993
rlabel metal2 1038 -2257 1038 -2257 0 net=8529
rlabel metal2 1290 -2257 1290 -2257 0 net=8687
rlabel metal2 156 -2259 156 -2259 0 net=5141
rlabel metal2 541 -2259 541 -2259 0 net=6737
rlabel metal2 1010 -2259 1010 -2259 0 net=7553
rlabel metal2 1199 -2259 1199 -2259 0 net=8973
rlabel metal2 1290 -2259 1290 -2259 0 net=9735
rlabel metal2 1584 -2259 1584 -2259 0 net=12193
rlabel metal2 128 -2261 128 -2261 0 net=11815
rlabel metal2 40 -2263 40 -2263 0 net=3337
rlabel metal2 289 -2263 289 -2263 0 net=1721
rlabel metal2 761 -2263 761 -2263 0 net=7433
rlabel metal2 982 -2263 982 -2263 0 net=7743
rlabel metal2 1297 -2263 1297 -2263 0 net=9817
rlabel metal2 173 -2265 173 -2265 0 net=10083
rlabel metal2 173 -2267 173 -2267 0 net=1225
rlabel metal2 1013 -2267 1013 -2267 0 net=8409
rlabel metal2 1045 -2267 1045 -2267 0 net=8069
rlabel metal2 1108 -2267 1108 -2267 0 net=12247
rlabel metal2 289 -2269 289 -2269 0 net=3291
rlabel metal2 436 -2269 436 -2269 0 net=4809
rlabel metal2 520 -2269 520 -2269 0 net=10449
rlabel metal2 1668 -2269 1668 -2269 0 net=12429
rlabel metal2 114 -2271 114 -2271 0 net=9621
rlabel metal2 548 -2271 548 -2271 0 net=4847
rlabel metal2 849 -2271 849 -2271 0 net=12431
rlabel metal2 149 -2273 149 -2273 0 net=3757
rlabel metal2 681 -2273 681 -2273 0 net=4247
rlabel metal2 1017 -2273 1017 -2273 0 net=7609
rlabel metal2 1059 -2273 1059 -2273 0 net=8249
rlabel metal2 1318 -2273 1318 -2273 0 net=10395
rlabel metal2 1591 -2273 1591 -2273 0 net=12177
rlabel metal2 149 -2275 149 -2275 0 net=4445
rlabel metal2 296 -2275 296 -2275 0 net=1734
rlabel metal2 478 -2275 478 -2275 0 net=3589
rlabel metal2 1052 -2275 1052 -2275 0 net=7345
rlabel metal2 1094 -2275 1094 -2275 0 net=11058
rlabel metal2 219 -2277 219 -2277 0 net=2425
rlabel metal2 478 -2277 478 -2277 0 net=4591
rlabel metal2 1073 -2277 1073 -2277 0 net=8659
rlabel metal2 1185 -2277 1185 -2277 0 net=8835
rlabel metal2 1332 -2277 1332 -2277 0 net=9583
rlabel metal2 1458 -2277 1458 -2277 0 net=10485
rlabel metal2 1556 -2277 1556 -2277 0 net=11147
rlabel metal2 247 -2279 247 -2279 0 net=1511
rlabel metal2 296 -2279 296 -2279 0 net=5107
rlabel metal2 1073 -2279 1073 -2279 0 net=8119
rlabel metal2 1353 -2279 1353 -2279 0 net=9661
rlabel metal2 1479 -2279 1479 -2279 0 net=10959
rlabel metal2 1556 -2279 1556 -2279 0 net=11669
rlabel metal2 79 -2281 79 -2281 0 net=2053
rlabel metal2 303 -2281 303 -2281 0 net=2873
rlabel metal2 457 -2281 457 -2281 0 net=5611
rlabel metal2 968 -2281 968 -2281 0 net=9913
rlabel metal2 1360 -2281 1360 -2281 0 net=10025
rlabel metal2 1493 -2281 1493 -2281 0 net=8851
rlabel metal2 79 -2283 79 -2283 0 net=1753
rlabel metal2 310 -2283 310 -2283 0 net=1888
rlabel metal2 1136 -2283 1136 -2283 0 net=9789
rlabel metal2 1304 -2283 1304 -2283 0 net=9239
rlabel metal2 86 -2285 86 -2285 0 net=3647
rlabel metal2 492 -2285 492 -2285 0 net=3066
rlabel metal2 723 -2285 723 -2285 0 net=5333
rlabel metal2 1374 -2285 1374 -2285 0 net=11359
rlabel metal2 1493 -2285 1493 -2285 0 net=12337
rlabel metal2 138 -2287 138 -2287 0 net=5551
rlabel metal2 310 -2287 310 -2287 0 net=4823
rlabel metal2 499 -2287 499 -2287 0 net=4299
rlabel metal2 653 -2287 653 -2287 0 net=12593
rlabel metal2 198 -2289 198 -2289 0 net=4765
rlabel metal2 1157 -2289 1157 -2289 0 net=9615
rlabel metal2 1269 -2289 1269 -2289 0 net=9135
rlabel metal2 317 -2291 317 -2291 0 net=2063
rlabel metal2 744 -2291 744 -2291 0 net=10335
rlabel metal2 324 -2293 324 -2293 0 net=6181
rlabel metal2 975 -2293 975 -2293 0 net=6915
rlabel metal2 1083 -2293 1083 -2293 0 net=9639
rlabel metal2 324 -2295 324 -2295 0 net=2085
rlabel metal2 373 -2295 373 -2295 0 net=3809
rlabel metal2 499 -2295 499 -2295 0 net=6153
rlabel metal2 989 -2295 989 -2295 0 net=8375
rlabel metal2 275 -2297 275 -2297 0 net=2609
rlabel metal2 429 -2297 429 -2297 0 net=6659
rlabel metal2 744 -2297 744 -2297 0 net=6106
rlabel metal2 954 -2297 954 -2297 0 net=8167
rlabel metal2 212 -2299 212 -2299 0 net=2043
rlabel metal2 331 -2299 331 -2299 0 net=3015
rlabel metal2 429 -2299 429 -2299 0 net=2919
rlabel metal2 863 -2299 863 -2299 0 net=7813
rlabel metal2 1157 -2299 1157 -2299 0 net=8717
rlabel metal2 331 -2301 331 -2301 0 net=2091
rlabel metal2 1164 -2301 1164 -2301 0 net=8787
rlabel metal2 338 -2303 338 -2303 0 net=2817
rlabel metal2 415 -2303 415 -2303 0 net=2833
rlabel metal2 912 -2303 912 -2303 0 net=6399
rlabel metal2 1171 -2303 1171 -2303 0 net=7497
rlabel metal2 1241 -2303 1241 -2303 0 net=9451
rlabel metal2 338 -2305 338 -2305 0 net=2455
rlabel metal2 912 -2305 912 -2305 0 net=6491
rlabel metal2 947 -2305 947 -2305 0 net=5211
rlabel metal2 352 -2307 352 -2307 0 net=2645
rlabel metal2 940 -2307 940 -2307 0 net=7367
rlabel metal2 1143 -2307 1143 -2307 0 net=9821
rlabel metal2 352 -2309 352 -2309 0 net=4159
rlabel metal2 1087 -2309 1087 -2309 0 net=8227
rlabel metal2 359 -2311 359 -2311 0 net=2387
rlabel metal2 576 -2311 576 -2311 0 net=4789
rlabel metal2 996 -2311 996 -2311 0 net=8793
rlabel metal2 387 -2313 387 -2313 0 net=3681
rlabel metal2 667 -2313 667 -2313 0 net=5589
rlabel metal2 996 -2313 996 -2313 0 net=9667
rlabel metal2 443 -2315 443 -2315 0 net=4751
rlabel metal2 443 -2317 443 -2317 0 net=4761
rlabel metal2 471 -2319 471 -2319 0 net=4139
rlabel metal2 527 -2321 527 -2321 0 net=7701
rlabel metal2 51 -2332 51 -2332 0 net=6054
rlabel metal2 215 -2332 215 -2332 0 net=6916
rlabel metal2 982 -2332 982 -2332 0 net=7744
rlabel metal2 999 -2332 999 -2332 0 net=10780
rlabel metal2 1514 -2332 1514 -2332 0 net=11126
rlabel metal2 1605 -2332 1605 -2332 0 net=8852
rlabel metal2 51 -2334 51 -2334 0 net=5907
rlabel metal2 443 -2334 443 -2334 0 net=4762
rlabel metal2 856 -2334 856 -2334 0 net=6182
rlabel metal2 982 -2334 982 -2334 0 net=8071
rlabel metal2 1076 -2334 1076 -2334 0 net=10378
rlabel metal2 1493 -2334 1493 -2334 0 net=12339
rlabel metal2 1605 -2334 1605 -2334 0 net=12643
rlabel metal2 79 -2336 79 -2336 0 net=1754
rlabel metal2 733 -2336 733 -2336 0 net=278
rlabel metal2 1171 -2336 1171 -2336 0 net=9136
rlabel metal2 1612 -2336 1612 -2336 0 net=10101
rlabel metal2 79 -2338 79 -2338 0 net=9359
rlabel metal2 100 -2338 100 -2338 0 net=1572
rlabel metal2 1171 -2338 1171 -2338 0 net=8795
rlabel metal2 1244 -2338 1244 -2338 0 net=12430
rlabel metal2 86 -2340 86 -2340 0 net=12594
rlabel metal2 86 -2342 86 -2342 0 net=3339
rlabel metal2 135 -2342 135 -2342 0 net=2426
rlabel metal2 415 -2342 415 -2342 0 net=2835
rlabel metal2 450 -2342 450 -2342 0 net=4662
rlabel metal2 597 -2342 597 -2342 0 net=1878
rlabel metal2 660 -2342 660 -2342 0 net=6446
rlabel metal2 684 -2342 684 -2342 0 net=11816
rlabel metal2 93 -2344 93 -2344 0 net=3017
rlabel metal2 464 -2344 464 -2344 0 net=3991
rlabel metal2 492 -2344 492 -2344 0 net=6660
rlabel metal2 775 -2344 775 -2344 0 net=9166
rlabel metal2 1437 -2344 1437 -2344 0 net=10877
rlabel metal2 100 -2346 100 -2346 0 net=2961
rlabel metal2 345 -2346 345 -2346 0 net=2993
rlabel metal2 457 -2346 457 -2346 0 net=3649
rlabel metal2 502 -2346 502 -2346 0 net=828
rlabel metal2 548 -2346 548 -2346 0 net=4849
rlabel metal2 597 -2346 597 -2346 0 net=5091
rlabel metal2 691 -2346 691 -2346 0 net=11148
rlabel metal2 65 -2348 65 -2348 0 net=4571
rlabel metal2 464 -2348 464 -2348 0 net=3811
rlabel metal2 527 -2348 527 -2348 0 net=7703
rlabel metal2 1080 -2348 1080 -2348 0 net=9240
rlabel metal2 1556 -2348 1556 -2348 0 net=11671
rlabel metal2 65 -2350 65 -2350 0 net=4447
rlabel metal2 163 -2350 163 -2350 0 net=4650
rlabel metal2 240 -2350 240 -2350 0 net=3305
rlabel metal2 422 -2350 422 -2350 0 net=2903
rlabel metal2 733 -2350 733 -2350 0 net=11365
rlabel metal2 1521 -2350 1521 -2350 0 net=12561
rlabel metal2 96 -2352 96 -2352 0 net=12623
rlabel metal2 107 -2354 107 -2354 0 net=5883
rlabel metal2 548 -2354 548 -2354 0 net=3859
rlabel metal2 569 -2354 569 -2354 0 net=7122
rlabel metal2 800 -2354 800 -2354 0 net=6468
rlabel metal2 1248 -2354 1248 -2354 0 net=9617
rlabel metal2 1248 -2354 1248 -2354 0 net=9617
rlabel metal2 1304 -2354 1304 -2354 0 net=11886
rlabel metal2 107 -2356 107 -2356 0 net=9493
rlabel metal2 149 -2356 149 -2356 0 net=2145
rlabel metal2 212 -2356 212 -2356 0 net=2777
rlabel metal2 530 -2356 530 -2356 0 net=7415
rlabel metal2 989 -2356 989 -2356 0 net=8377
rlabel metal2 58 -2358 58 -2358 0 net=6429
rlabel metal2 212 -2358 212 -2358 0 net=8490
rlabel metal2 1304 -2358 1304 -2358 0 net=9915
rlabel metal2 1384 -2358 1384 -2358 0 net=11306
rlabel metal2 114 -2360 114 -2360 0 net=6154
rlabel metal2 576 -2360 576 -2360 0 net=4791
rlabel metal2 779 -2360 779 -2360 0 net=5439
rlabel metal2 856 -2360 856 -2360 0 net=12114
rlabel metal2 44 -2362 44 -2362 0 net=8341
rlabel metal2 618 -2362 618 -2362 0 net=3854
rlabel metal2 695 -2362 695 -2362 0 net=5713
rlabel metal2 863 -2362 863 -2362 0 net=7814
rlabel metal2 1178 -2362 1178 -2362 0 net=9137
rlabel metal2 1314 -2362 1314 -2362 0 net=12718
rlabel metal2 114 -2364 114 -2364 0 net=2389
rlabel metal2 432 -2364 432 -2364 0 net=6321
rlabel metal2 625 -2364 625 -2364 0 net=1723
rlabel metal2 1521 -2364 1521 -2364 0 net=12433
rlabel metal2 117 -2366 117 -2366 0 net=2019
rlabel metal2 240 -2366 240 -2366 0 net=3683
rlabel metal2 471 -2366 471 -2366 0 net=4141
rlabel metal2 590 -2366 590 -2366 0 net=4281
rlabel metal2 632 -2366 632 -2366 0 net=3590
rlabel metal2 863 -2366 863 -2366 0 net=9275
rlabel metal2 1283 -2366 1283 -2366 0 net=10111
rlabel metal2 1388 -2366 1388 -2366 0 net=11531
rlabel metal2 1570 -2366 1570 -2366 0 net=12195
rlabel metal2 128 -2368 128 -2368 0 net=5143
rlabel metal2 163 -2368 163 -2368 0 net=6669
rlabel metal2 870 -2368 870 -2368 0 net=6363
rlabel metal2 898 -2368 898 -2368 0 net=12546
rlabel metal2 135 -2370 135 -2370 0 net=5283
rlabel metal2 632 -2370 632 -2370 0 net=5213
rlabel metal2 954 -2370 954 -2370 0 net=10684
rlabel metal2 142 -2372 142 -2372 0 net=6345
rlabel metal2 898 -2372 898 -2372 0 net=8168
rlabel metal2 1332 -2372 1332 -2372 0 net=12230
rlabel metal2 142 -2374 142 -2374 0 net=4593
rlabel metal2 499 -2374 499 -2374 0 net=1389
rlabel metal2 1097 -2374 1097 -2374 0 net=10172
rlabel metal2 1388 -2374 1388 -2374 0 net=10337
rlabel metal2 1451 -2374 1451 -2374 0 net=11495
rlabel metal2 1598 -2374 1598 -2374 0 net=7711
rlabel metal2 170 -2376 170 -2376 0 net=3758
rlabel metal2 541 -2376 541 -2376 0 net=6738
rlabel metal2 828 -2376 828 -2376 0 net=6005
rlabel metal2 873 -2376 873 -2376 0 net=10668
rlabel metal2 170 -2378 170 -2378 0 net=4767
rlabel metal2 215 -2378 215 -2378 0 net=8628
rlabel metal2 688 -2378 688 -2378 0 net=5335
rlabel metal2 828 -2378 828 -2378 0 net=6959
rlabel metal2 1080 -2378 1080 -2378 0 net=7007
rlabel metal2 1108 -2378 1108 -2378 0 net=12249
rlabel metal2 156 -2380 156 -2380 0 net=7401
rlabel metal2 695 -2380 695 -2380 0 net=5613
rlabel metal2 723 -2380 723 -2380 0 net=5515
rlabel metal2 905 -2380 905 -2380 0 net=6617
rlabel metal2 905 -2380 905 -2380 0 net=6617
rlabel metal2 919 -2380 919 -2380 0 net=7435
rlabel metal2 996 -2380 996 -2380 0 net=7545
rlabel metal2 1066 -2380 1066 -2380 0 net=8661
rlabel metal2 1192 -2380 1192 -2380 0 net=9841
rlabel metal2 1395 -2380 1395 -2380 0 net=10405
rlabel metal2 198 -2382 198 -2382 0 net=5109
rlabel metal2 345 -2382 345 -2382 0 net=2819
rlabel metal2 387 -2382 387 -2382 0 net=2397
rlabel metal2 478 -2382 478 -2382 0 net=4249
rlabel metal2 709 -2382 709 -2382 0 net=5939
rlabel metal2 793 -2382 793 -2382 0 net=8401
rlabel metal2 1122 -2382 1122 -2382 0 net=8615
rlabel metal2 1143 -2382 1143 -2382 0 net=8975
rlabel metal2 1255 -2382 1255 -2382 0 net=9883
rlabel metal2 1374 -2382 1374 -2382 0 net=11361
rlabel metal2 226 -2384 226 -2384 0 net=2055
rlabel metal2 254 -2384 254 -2384 0 net=1513
rlabel metal2 268 -2384 268 -2384 0 net=4051
rlabel metal2 590 -2384 590 -2384 0 net=3129
rlabel metal2 639 -2384 639 -2384 0 net=10450
rlabel metal2 184 -2386 184 -2386 0 net=4239
rlabel metal2 254 -2386 254 -2386 0 net=2646
rlabel metal2 471 -2386 471 -2386 0 net=4752
rlabel metal2 786 -2386 786 -2386 0 net=5865
rlabel metal2 919 -2386 919 -2386 0 net=9043
rlabel metal2 1339 -2386 1339 -2386 0 net=10027
rlabel metal2 1374 -2386 1374 -2386 0 net=10447
rlabel metal2 184 -2388 184 -2388 0 net=3089
rlabel metal2 901 -2388 901 -2388 0 net=11019
rlabel metal2 268 -2390 268 -2390 0 net=2921
rlabel metal2 513 -2390 513 -2390 0 net=9623
rlabel metal2 1185 -2390 1185 -2390 0 net=8837
rlabel metal2 1360 -2390 1360 -2390 0 net=10275
rlabel metal2 1409 -2390 1409 -2390 0 net=10961
rlabel metal2 282 -2392 282 -2392 0 net=4629
rlabel metal2 520 -2392 520 -2392 0 net=3659
rlabel metal2 786 -2392 786 -2392 0 net=5843
rlabel metal2 901 -2392 901 -2392 0 net=9662
rlabel metal2 1479 -2392 1479 -2392 0 net=11889
rlabel metal2 282 -2394 282 -2394 0 net=3293
rlabel metal2 296 -2394 296 -2394 0 net=4331
rlabel metal2 814 -2394 814 -2394 0 net=6917
rlabel metal2 926 -2394 926 -2394 0 net=6995
rlabel metal2 957 -2394 957 -2394 0 net=10003
rlabel metal2 1346 -2394 1346 -2394 0 net=10435
rlabel metal2 1430 -2394 1430 -2394 0 net=12179
rlabel metal2 173 -2396 173 -2396 0 net=3783
rlabel metal2 303 -2396 303 -2396 0 net=5553
rlabel metal2 555 -2396 555 -2396 0 net=3160
rlabel metal2 646 -2396 646 -2396 0 net=6281
rlabel metal2 772 -2396 772 -2396 0 net=7263
rlabel metal2 884 -2396 884 -2396 0 net=7179
rlabel metal2 933 -2396 933 -2396 0 net=6773
rlabel metal2 971 -2396 971 -2396 0 net=10486
rlabel metal2 1577 -2396 1577 -2396 0 net=7540
rlabel metal2 177 -2398 177 -2398 0 net=2945
rlabel metal2 310 -2398 310 -2398 0 net=4825
rlabel metal2 604 -2398 604 -2398 0 net=6037
rlabel metal2 821 -2398 821 -2398 0 net=7324
rlabel metal2 58 -2400 58 -2400 0 net=4595
rlabel metal2 338 -2400 338 -2400 0 net=2457
rlabel metal2 653 -2400 653 -2400 0 net=5591
rlabel metal2 716 -2400 716 -2400 0 net=5913
rlabel metal2 744 -2400 744 -2400 0 net=6492
rlabel metal2 1024 -2400 1024 -2400 0 net=8411
rlabel metal2 1115 -2400 1115 -2400 0 net=6401
rlabel metal2 177 -2402 177 -2402 0 net=4810
rlabel metal2 667 -2402 667 -2402 0 net=5961
rlabel metal2 842 -2402 842 -2402 0 net=6513
rlabel metal2 891 -2402 891 -2402 0 net=7069
rlabel metal2 1017 -2402 1017 -2402 0 net=7611
rlabel metal2 1031 -2402 1031 -2402 0 net=9191
rlabel metal2 1318 -2402 1318 -2402 0 net=10397
rlabel metal2 1458 -2402 1458 -2402 0 net=11435
rlabel metal2 191 -2404 191 -2404 0 net=2225
rlabel metal2 352 -2404 352 -2404 0 net=4161
rlabel metal2 737 -2404 737 -2404 0 net=3737
rlabel metal2 842 -2404 842 -2404 0 net=7874
rlabel metal2 1038 -2404 1038 -2404 0 net=8531
rlabel metal2 1136 -2404 1136 -2404 0 net=9791
rlabel metal2 1535 -2404 1535 -2404 0 net=11029
rlabel metal2 191 -2406 191 -2406 0 net=2093
rlabel metal2 359 -2406 359 -2406 0 net=2611
rlabel metal2 436 -2406 436 -2406 0 net=4301
rlabel metal2 751 -2406 751 -2406 0 net=5547
rlabel metal2 1003 -2406 1003 -2406 0 net=9737
rlabel metal2 219 -2408 219 -2408 0 net=2259
rlabel metal2 506 -2408 506 -2408 0 net=3609
rlabel metal2 758 -2408 758 -2408 0 net=7657
rlabel metal2 1038 -2408 1038 -2408 0 net=8251
rlabel metal2 1115 -2408 1115 -2408 0 net=8719
rlabel metal2 1185 -2408 1185 -2408 0 net=9823
rlabel metal2 219 -2410 219 -2410 0 net=2065
rlabel metal2 324 -2410 324 -2410 0 net=2087
rlabel metal2 758 -2410 758 -2410 0 net=9107
rlabel metal2 1290 -2410 1290 -2410 0 net=10085
rlabel metal2 121 -2412 121 -2412 0 net=2197
rlabel metal2 324 -2412 324 -2412 0 net=3531
rlabel metal2 891 -2412 891 -2412 0 net=7554
rlabel metal2 1059 -2412 1059 -2412 0 net=8229
rlabel metal2 1136 -2412 1136 -2412 0 net=7709
rlabel metal2 72 -2414 72 -2414 0 net=2345
rlabel metal2 331 -2414 331 -2414 0 net=2175
rlabel metal2 961 -2414 961 -2414 0 net=7483
rlabel metal2 1073 -2414 1073 -2414 0 net=8121
rlabel metal2 1157 -2414 1157 -2414 0 net=8789
rlabel metal2 1199 -2414 1199 -2414 0 net=9259
rlabel metal2 1220 -2414 1220 -2414 0 net=7499
rlabel metal2 1325 -2414 1325 -2414 0 net=9497
rlabel metal2 1381 -2414 1381 -2414 0 net=9584
rlabel metal2 72 -2416 72 -2416 0 net=4211
rlabel metal2 1164 -2416 1164 -2416 0 net=8689
rlabel metal2 537 -2418 537 -2418 0 net=9329
rlabel metal2 1234 -2418 1234 -2418 0 net=9453
rlabel metal2 1276 -2418 1276 -2418 0 net=10621
rlabel metal2 933 -2420 933 -2420 0 net=6525
rlabel metal2 1206 -2420 1206 -2420 0 net=9818
rlabel metal2 940 -2422 940 -2422 0 net=7369
rlabel metal2 1241 -2422 1241 -2422 0 net=12351
rlabel metal2 940 -2424 940 -2424 0 net=7303
rlabel metal2 961 -2426 961 -2426 0 net=7347
rlabel metal2 1262 -2426 1262 -2426 0 net=9641
rlabel metal2 705 -2428 705 -2428 0 net=8101
rlabel metal2 1262 -2428 1262 -2428 0 net=9669
rlabel metal2 408 -2430 408 -2430 0 net=5980
rlabel metal2 1269 -2430 1269 -2430 0 net=10043
rlabel metal2 275 -2432 275 -2432 0 net=2045
rlabel metal2 1367 -2432 1367 -2432 0 net=10713
rlabel metal2 275 -2434 275 -2434 0 net=2875
rlabel metal2 1465 -2434 1465 -2434 0 net=11157
rlabel metal2 394 -2436 394 -2436 0 net=7325
rlabel metal2 1507 -2436 1507 -2436 0 net=12379
rlabel metal2 44 -2447 44 -2447 0 net=6671
rlabel metal2 184 -2447 184 -2447 0 net=3090
rlabel metal2 681 -2447 681 -2447 0 net=152
rlabel metal2 754 -2447 754 -2447 0 net=5714
rlabel metal2 786 -2447 786 -2447 0 net=5844
rlabel metal2 912 -2447 912 -2447 0 net=7071
rlabel metal2 86 -2449 86 -2449 0 net=3341
rlabel metal2 212 -2449 212 -2449 0 net=2965
rlabel metal2 212 -2449 212 -2449 0 net=2965
rlabel metal2 233 -2449 233 -2449 0 net=2021
rlabel metal2 233 -2449 233 -2449 0 net=2021
rlabel metal2 240 -2449 240 -2449 0 net=3684
rlabel metal2 870 -2449 870 -2449 0 net=6365
rlabel metal2 947 -2449 947 -2449 0 net=6775
rlabel metal2 947 -2449 947 -2449 0 net=6775
rlabel metal2 957 -2449 957 -2449 0 net=7546
rlabel metal2 1062 -2449 1062 -2449 0 net=11405
rlabel metal2 1675 -2449 1675 -2449 0 net=10103
rlabel metal2 86 -2451 86 -2451 0 net=5093
rlabel metal2 611 -2451 611 -2451 0 net=12434
rlabel metal2 1528 -2451 1528 -2451 0 net=12624
rlabel metal2 100 -2453 100 -2453 0 net=2963
rlabel metal2 257 -2453 257 -2453 0 net=4479
rlabel metal2 688 -2453 688 -2453 0 net=5336
rlabel metal2 779 -2453 779 -2453 0 net=5441
rlabel metal2 807 -2453 807 -2453 0 net=6996
rlabel metal2 971 -2453 971 -2453 0 net=8378
rlabel metal2 1605 -2453 1605 -2453 0 net=12645
rlabel metal2 107 -2455 107 -2455 0 net=9494
rlabel metal2 891 -2455 891 -2455 0 net=6939
rlabel metal2 1076 -2455 1076 -2455 0 net=10398
rlabel metal2 1367 -2455 1367 -2455 0 net=10715
rlabel metal2 1538 -2455 1538 -2455 0 net=11672
rlabel metal2 1577 -2455 1577 -2455 0 net=10781
rlabel metal2 72 -2457 72 -2457 0 net=4213
rlabel metal2 142 -2457 142 -2457 0 net=4594
rlabel metal2 180 -2457 180 -2457 0 net=10495
rlabel metal2 821 -2457 821 -2457 0 net=11387
rlabel metal2 142 -2459 142 -2459 0 net=1973
rlabel metal2 642 -2459 642 -2459 0 net=39
rlabel metal2 1227 -2459 1227 -2459 0 net=9793
rlabel metal2 1381 -2459 1381 -2459 0 net=11890
rlabel metal2 1500 -2459 1500 -2459 0 net=12251
rlabel metal2 152 -2461 152 -2461 0 net=10086
rlabel metal2 1300 -2461 1300 -2461 0 net=12180
rlabel metal2 1458 -2461 1458 -2461 0 net=11437
rlabel metal2 282 -2463 282 -2463 0 net=3294
rlabel metal2 562 -2463 562 -2463 0 net=4143
rlabel metal2 702 -2463 702 -2463 0 net=6961
rlabel metal2 842 -2463 842 -2463 0 net=5153
rlabel metal2 1115 -2463 1115 -2463 0 net=8721
rlabel metal2 1244 -2463 1244 -2463 0 net=9916
rlabel metal2 1311 -2463 1311 -2463 0 net=10795
rlabel metal2 1556 -2463 1556 -2463 0 net=12563
rlabel metal2 261 -2465 261 -2465 0 net=1515
rlabel metal2 296 -2465 296 -2465 0 net=4333
rlabel metal2 492 -2465 492 -2465 0 net=3651
rlabel metal2 593 -2465 593 -2465 0 net=7710
rlabel metal2 1157 -2465 1157 -2465 0 net=8791
rlabel metal2 226 -2467 226 -2467 0 net=2057
rlabel metal2 296 -2467 296 -2467 0 net=2261
rlabel metal2 411 -2467 411 -2467 0 net=3812
rlabel metal2 502 -2467 502 -2467 0 net=11915
rlabel metal2 93 -2469 93 -2469 0 net=3019
rlabel metal2 422 -2469 422 -2469 0 net=2905
rlabel metal2 506 -2469 506 -2469 0 net=3611
rlabel metal2 716 -2469 716 -2469 0 net=5915
rlabel metal2 845 -2469 845 -2469 0 net=10044
rlabel metal2 1276 -2469 1276 -2469 0 net=9643
rlabel metal2 1395 -2469 1395 -2469 0 net=10407
rlabel metal2 65 -2471 65 -2471 0 net=4449
rlabel metal2 226 -2471 226 -2471 0 net=2199
rlabel metal2 324 -2471 324 -2471 0 net=3532
rlabel metal2 506 -2471 506 -2471 0 net=3555
rlabel metal2 730 -2471 730 -2471 0 net=7370
rlabel metal2 1129 -2471 1129 -2471 0 net=8533
rlabel metal2 1199 -2471 1199 -2471 0 net=9261
rlabel metal2 1314 -2471 1314 -2471 0 net=1724
rlabel metal2 1507 -2471 1507 -2471 0 net=12381
rlabel metal2 65 -2473 65 -2473 0 net=9360
rlabel metal2 100 -2473 100 -2473 0 net=7351
rlabel metal2 324 -2473 324 -2473 0 net=2047
rlabel metal2 422 -2473 422 -2473 0 net=3993
rlabel metal2 513 -2473 513 -2473 0 net=4630
rlabel metal2 583 -2473 583 -2473 0 net=4851
rlabel metal2 751 -2473 751 -2473 0 net=5549
rlabel metal2 1465 -2473 1465 -2473 0 net=11159
rlabel metal2 58 -2475 58 -2475 0 net=4597
rlabel metal2 513 -2475 513 -2475 0 net=3131
rlabel metal2 597 -2475 597 -2475 0 net=5593
rlabel metal2 751 -2475 751 -2475 0 net=11005
rlabel metal2 58 -2477 58 -2477 0 net=5215
rlabel metal2 765 -2477 765 -2477 0 net=6283
rlabel metal2 919 -2477 919 -2477 0 net=9045
rlabel metal2 1276 -2477 1276 -2477 0 net=11497
rlabel metal2 1507 -2477 1507 -2477 0 net=12197
rlabel metal2 79 -2479 79 -2479 0 net=2821
rlabel metal2 401 -2479 401 -2479 0 net=5555
rlabel metal2 793 -2479 793 -2479 0 net=5867
rlabel metal2 852 -2479 852 -2479 0 net=8616
rlabel metal2 1129 -2479 1129 -2479 0 net=7713
rlabel metal2 121 -2481 121 -2481 0 net=2347
rlabel metal2 408 -2481 408 -2481 0 net=1075
rlabel metal2 929 -2481 929 -2481 0 net=10511
rlabel metal2 1514 -2481 1514 -2481 0 net=12341
rlabel metal2 121 -2483 121 -2483 0 net=5145
rlabel metal2 215 -2483 215 -2483 0 net=10873
rlabel metal2 128 -2485 128 -2485 0 net=2147
rlabel metal2 303 -2485 303 -2485 0 net=2946
rlabel metal2 436 -2485 436 -2485 0 net=4303
rlabel metal2 520 -2485 520 -2485 0 net=3660
rlabel metal2 677 -2485 677 -2485 0 net=11739
rlabel metal2 75 -2487 75 -2487 0 net=5989
rlabel metal2 450 -2487 450 -2487 0 net=2995
rlabel metal2 674 -2487 674 -2487 0 net=4409
rlabel metal2 877 -2487 877 -2487 0 net=6347
rlabel metal2 1024 -2487 1024 -2487 0 net=7613
rlabel metal2 1167 -2487 1167 -2487 0 net=10962
rlabel metal2 1416 -2487 1416 -2487 0 net=10623
rlabel metal2 149 -2489 149 -2489 0 net=3225
rlabel metal2 303 -2489 303 -2489 0 net=2399
rlabel metal2 429 -2489 429 -2489 0 net=11457
rlabel metal2 310 -2491 310 -2491 0 net=2459
rlabel metal2 387 -2491 387 -2491 0 net=4573
rlabel metal2 474 -2491 474 -2491 0 net=3111
rlabel metal2 520 -2491 520 -2491 0 net=7349
rlabel metal2 982 -2491 982 -2491 0 net=8073
rlabel metal2 1031 -2491 1031 -2491 0 net=9193
rlabel metal2 1332 -2491 1332 -2491 0 net=10005
rlabel metal2 1472 -2491 1472 -2491 0 net=11367
rlabel metal2 103 -2493 103 -2493 0 net=1927
rlabel metal2 432 -2493 432 -2493 0 net=12577
rlabel metal2 313 -2495 313 -2495 0 net=2612
rlabel metal2 443 -2495 443 -2495 0 net=2837
rlabel metal2 527 -2495 527 -2495 0 net=4052
rlabel metal2 576 -2495 576 -2495 0 net=8343
rlabel metal2 247 -2497 247 -2497 0 net=4241
rlabel metal2 366 -2497 366 -2497 0 net=2089
rlabel metal2 541 -2497 541 -2497 0 net=5517
rlabel metal2 877 -2497 877 -2497 0 net=6083
rlabel metal2 933 -2497 933 -2497 0 net=6527
rlabel metal2 1031 -2497 1031 -2497 0 net=7371
rlabel metal2 1199 -2497 1199 -2497 0 net=9885
rlabel metal2 1290 -2497 1290 -2497 0 net=10339
rlabel metal2 1395 -2497 1395 -2497 0 net=12353
rlabel metal2 219 -2499 219 -2499 0 net=2067
rlabel metal2 275 -2499 275 -2499 0 net=2877
rlabel metal2 415 -2499 415 -2499 0 net=2778
rlabel metal2 534 -2499 534 -2499 0 net=5885
rlabel metal2 810 -2499 810 -2499 0 net=9831
rlabel metal2 1542 -2499 1542 -2499 0 net=11031
rlabel metal2 198 -2501 198 -2501 0 net=5111
rlabel metal2 275 -2501 275 -2501 0 net=1655
rlabel metal2 884 -2501 884 -2501 0 net=6515
rlabel metal2 933 -2501 933 -2501 0 net=6317
rlabel metal2 1325 -2501 1325 -2501 0 net=9499
rlabel metal2 1339 -2501 1339 -2501 0 net=10029
rlabel metal2 173 -2503 173 -2503 0 net=4059
rlabel metal2 331 -2503 331 -2503 0 net=2177
rlabel metal2 534 -2503 534 -2503 0 net=4911
rlabel metal2 1038 -2503 1038 -2503 0 net=8253
rlabel metal2 1178 -2503 1178 -2503 0 net=9139
rlabel metal2 1339 -2503 1339 -2503 0 net=9511
rlabel metal2 51 -2505 51 -2505 0 net=5909
rlabel metal2 1003 -2505 1003 -2505 0 net=9739
rlabel metal2 1052 -2505 1052 -2505 0 net=8103
rlabel metal2 1185 -2505 1185 -2505 0 net=9825
rlabel metal2 1444 -2505 1444 -2505 0 net=11021
rlabel metal2 51 -2507 51 -2507 0 net=4769
rlabel metal2 268 -2507 268 -2507 0 net=2923
rlabel metal2 338 -2507 338 -2507 0 net=2227
rlabel metal2 415 -2507 415 -2507 0 net=4313
rlabel metal2 548 -2507 548 -2507 0 net=3861
rlabel metal2 590 -2507 590 -2507 0 net=6275
rlabel metal2 663 -2507 663 -2507 0 net=8523
rlabel metal2 1185 -2507 1185 -2507 0 net=11362
rlabel metal2 268 -2509 268 -2509 0 net=3785
rlabel metal2 338 -2509 338 -2509 0 net=3307
rlabel metal2 548 -2509 548 -2509 0 net=7729
rlabel metal2 1206 -2509 1206 -2509 0 net=11643
rlabel metal2 163 -2511 163 -2511 0 net=8617
rlabel metal2 1209 -2511 1209 -2511 0 net=10293
rlabel metal2 289 -2513 289 -2513 0 net=1867
rlabel metal2 569 -2513 569 -2513 0 net=6039
rlabel metal2 625 -2513 625 -2513 0 net=4283
rlabel metal2 695 -2513 695 -2513 0 net=5615
rlabel metal2 821 -2513 821 -2513 0 net=10143
rlabel metal2 156 -2515 156 -2515 0 net=7402
rlabel metal2 733 -2515 733 -2515 0 net=1460
rlabel metal2 156 -2517 156 -2517 0 net=2305
rlabel metal2 835 -2517 835 -2517 0 net=6007
rlabel metal2 926 -2517 926 -2517 0 net=7181
rlabel metal2 1010 -2517 1010 -2517 0 net=7485
rlabel metal2 1059 -2517 1059 -2517 0 net=8231
rlabel metal2 1083 -2517 1083 -2517 0 net=3699
rlabel metal2 1213 -2517 1213 -2517 0 net=8839
rlabel metal2 555 -2519 555 -2519 0 net=4827
rlabel metal2 709 -2519 709 -2519 0 net=5941
rlabel metal2 926 -2519 926 -2519 0 net=8431
rlabel metal2 1059 -2519 1059 -2519 0 net=9624
rlabel metal2 1213 -2519 1213 -2519 0 net=7501
rlabel metal2 1360 -2519 1360 -2519 0 net=10277
rlabel metal2 576 -2521 576 -2521 0 net=3739
rlabel metal2 863 -2521 863 -2521 0 net=9277
rlabel metal2 135 -2523 135 -2523 0 net=5284
rlabel metal2 863 -2523 863 -2523 0 net=6619
rlabel metal2 975 -2523 975 -2523 0 net=7417
rlabel metal2 1066 -2523 1066 -2523 0 net=8663
rlabel metal2 135 -2525 135 -2525 0 net=2095
rlabel metal2 394 -2525 394 -2525 0 net=7327
rlabel metal2 1087 -2525 1087 -2525 0 net=8123
rlabel metal2 1220 -2525 1220 -2525 0 net=9331
rlabel metal2 114 -2527 114 -2527 0 net=2391
rlabel metal2 394 -2527 394 -2527 0 net=5963
rlabel metal2 705 -2527 705 -2527 0 net=6521
rlabel metal2 1087 -2527 1087 -2527 0 net=11743
rlabel metal2 114 -2529 114 -2529 0 net=6323
rlabel metal2 660 -2529 660 -2529 0 net=4792
rlabel metal2 814 -2529 814 -2529 0 net=6919
rlabel metal2 1090 -2529 1090 -2529 0 net=11105
rlabel metal2 68 -2531 68 -2531 0 net=7361
rlabel metal2 660 -2531 660 -2531 0 net=10448
rlabel metal2 604 -2533 604 -2533 0 net=7305
rlabel metal2 1220 -2533 1220 -2533 0 net=6403
rlabel metal2 478 -2535 478 -2535 0 net=4251
rlabel metal2 1248 -2535 1248 -2535 0 net=9619
rlabel metal2 205 -2537 205 -2537 0 net=6431
rlabel metal2 667 -2537 667 -2537 0 net=1817
rlabel metal2 1143 -2537 1143 -2537 0 net=8977
rlabel metal2 1255 -2537 1255 -2537 0 net=10113
rlabel metal2 1374 -2537 1374 -2537 0 net=11533
rlabel metal2 1535 -2537 1535 -2537 0 net=11173
rlabel metal2 205 -2539 205 -2539 0 net=2461
rlabel metal2 1045 -2539 1045 -2539 0 net=7705
rlabel metal2 1234 -2539 1234 -2539 0 net=9455
rlabel metal2 1402 -2539 1402 -2539 0 net=10437
rlabel metal2 709 -2541 709 -2541 0 net=2131
rlabel metal2 814 -2541 814 -2541 0 net=5563
rlabel metal2 856 -2541 856 -2541 0 net=6531
rlabel metal2 989 -2541 989 -2541 0 net=7437
rlabel metal2 1171 -2541 1171 -2541 0 net=8797
rlabel metal2 1262 -2541 1262 -2541 0 net=9671
rlabel metal2 1437 -2541 1437 -2541 0 net=10879
rlabel metal2 555 -2543 555 -2543 0 net=5543
rlabel metal2 856 -2543 856 -2543 0 net=2799
rlabel metal2 989 -2543 989 -2543 0 net=8413
rlabel metal2 1164 -2543 1164 -2543 0 net=8691
rlabel metal2 1283 -2543 1283 -2543 0 net=9843
rlabel metal2 758 -2545 758 -2545 0 net=9109
rlabel metal2 730 -2547 730 -2547 0 net=3645
rlabel metal2 1017 -2547 1017 -2547 0 net=7659
rlabel metal2 1164 -2547 1164 -2547 0 net=10357
rlabel metal2 772 -2549 772 -2549 0 net=7265
rlabel metal2 1101 -2549 1101 -2549 0 net=8403
rlabel metal2 1195 -2549 1195 -2549 0 net=10255
rlabel metal2 646 -2551 646 -2551 0 net=4163
rlabel metal2 1080 -2551 1080 -2551 0 net=7009
rlabel metal2 345 -2553 345 -2553 0 net=4381
rlabel metal2 1080 -2553 1080 -2553 0 net=8563
rlabel metal2 72 -2564 72 -2564 0 net=6432
rlabel metal2 513 -2564 513 -2564 0 net=3132
rlabel metal2 789 -2564 789 -2564 0 net=8664
rlabel metal2 1678 -2564 1678 -2564 0 net=10104
rlabel metal2 75 -2566 75 -2566 0 net=11006
rlabel metal2 1703 -2566 1703 -2566 0 net=10782
rlabel metal2 79 -2568 79 -2568 0 net=2822
rlabel metal2 460 -2568 460 -2568 0 net=7306
rlabel metal2 618 -2568 618 -2568 0 net=7362
rlabel metal2 1192 -2568 1192 -2568 0 net=8535
rlabel metal2 1192 -2568 1192 -2568 0 net=8535
rlabel metal2 1346 -2568 1346 -2568 0 net=9645
rlabel metal2 1346 -2568 1346 -2568 0 net=9645
rlabel metal2 1430 -2568 1430 -2568 0 net=10513
rlabel metal2 1563 -2568 1563 -2568 0 net=11459
rlabel metal2 1703 -2568 1703 -2568 0 net=12579
rlabel metal2 93 -2570 93 -2570 0 net=4451
rlabel metal2 93 -2570 93 -2570 0 net=4451
rlabel metal2 100 -2570 100 -2570 0 net=5910
rlabel metal2 873 -2570 873 -2570 0 net=8564
rlabel metal2 1500 -2570 1500 -2570 0 net=11161
rlabel metal2 1626 -2570 1626 -2570 0 net=11917
rlabel metal2 100 -2572 100 -2572 0 net=2097
rlabel metal2 149 -2572 149 -2572 0 net=7328
rlabel metal2 1080 -2572 1080 -2572 0 net=7715
rlabel metal2 1178 -2572 1178 -2572 0 net=8525
rlabel metal2 1374 -2572 1374 -2572 0 net=11535
rlabel metal2 128 -2574 128 -2574 0 net=2149
rlabel metal2 170 -2574 170 -2574 0 net=2348
rlabel metal2 429 -2574 429 -2574 0 net=2800
rlabel metal2 873 -2574 873 -2574 0 net=8692
rlabel metal2 1374 -2574 1374 -2574 0 net=10145
rlabel metal2 58 -2576 58 -2576 0 net=5217
rlabel metal2 432 -2576 432 -2576 0 net=2090
rlabel metal2 548 -2576 548 -2576 0 net=5550
rlabel metal2 58 -2578 58 -2578 0 net=2049
rlabel metal2 373 -2578 373 -2578 0 net=1929
rlabel metal2 436 -2578 436 -2578 0 net=5991
rlabel metal2 555 -2578 555 -2578 0 net=5545
rlabel metal2 793 -2578 793 -2578 0 net=5617
rlabel metal2 793 -2578 793 -2578 0 net=5617
rlabel metal2 800 -2578 800 -2578 0 net=10497
rlabel metal2 1458 -2578 1458 -2578 0 net=12383
rlabel metal2 44 -2580 44 -2580 0 net=6673
rlabel metal2 576 -2580 576 -2580 0 net=3740
rlabel metal2 845 -2580 845 -2580 0 net=10030
rlabel metal2 44 -2582 44 -2582 0 net=8867
rlabel metal2 121 -2582 121 -2582 0 net=5147
rlabel metal2 201 -2582 201 -2582 0 net=8344
rlabel metal2 1542 -2582 1542 -2582 0 net=11023
rlabel metal2 128 -2584 128 -2584 0 net=5965
rlabel metal2 436 -2584 436 -2584 0 net=3419
rlabel metal2 506 -2584 506 -2584 0 net=3557
rlabel metal2 856 -2584 856 -2584 0 net=6285
rlabel metal2 898 -2584 898 -2584 0 net=6349
rlabel metal2 898 -2584 898 -2584 0 net=6349
rlabel metal2 926 -2584 926 -2584 0 net=9620
rlabel metal2 135 -2586 135 -2586 0 net=2769
rlabel metal2 670 -2586 670 -2586 0 net=10408
rlabel metal2 152 -2588 152 -2588 0 net=12541
rlabel metal2 240 -2590 240 -2590 0 net=2964
rlabel metal2 593 -2590 593 -2590 0 net=4144
rlabel metal2 625 -2590 625 -2590 0 net=7072
rlabel metal2 240 -2592 240 -2592 0 net=2059
rlabel metal2 268 -2592 268 -2592 0 net=3787
rlabel metal2 600 -2592 600 -2592 0 net=7706
rlabel metal2 1178 -2592 1178 -2592 0 net=8723
rlabel metal2 1262 -2592 1262 -2592 0 net=9195
rlabel metal2 1395 -2592 1395 -2592 0 net=12355
rlabel metal2 1696 -2592 1696 -2592 0 net=12647
rlabel metal2 226 -2594 226 -2594 0 net=2201
rlabel metal2 303 -2594 303 -2594 0 net=2401
rlabel metal2 401 -2594 401 -2594 0 net=5181
rlabel metal2 905 -2594 905 -2594 0 net=6523
rlabel metal2 954 -2594 954 -2594 0 net=10294
rlabel metal2 212 -2596 212 -2596 0 net=2967
rlabel metal2 233 -2596 233 -2596 0 net=2023
rlabel metal2 324 -2596 324 -2596 0 net=2229
rlabel metal2 506 -2596 506 -2596 0 net=6055
rlabel metal2 604 -2596 604 -2596 0 net=4411
rlabel metal2 681 -2596 681 -2596 0 net=4481
rlabel metal2 681 -2596 681 -2596 0 net=4481
rlabel metal2 730 -2596 730 -2596 0 net=4252
rlabel metal2 975 -2596 975 -2596 0 net=6921
rlabel metal2 975 -2596 975 -2596 0 net=6921
rlabel metal2 1034 -2596 1034 -2596 0 net=8153
rlabel metal2 1213 -2596 1213 -2596 0 net=7503
rlabel metal2 1395 -2596 1395 -2596 0 net=10257
rlabel metal2 1451 -2596 1451 -2596 0 net=10717
rlabel metal2 117 -2598 117 -2598 0 net=6577
rlabel metal2 1038 -2598 1038 -2598 0 net=9740
rlabel metal2 1087 -2598 1087 -2598 0 net=9111
rlabel metal2 1416 -2598 1416 -2598 0 net=10439
rlabel metal2 163 -2600 163 -2600 0 net=4541
rlabel metal2 611 -2600 611 -2600 0 net=4829
rlabel metal2 733 -2600 733 -2600 0 net=12459
rlabel metal2 163 -2602 163 -2602 0 net=457
rlabel metal2 632 -2602 632 -2602 0 net=4284
rlabel metal2 649 -2602 649 -2602 0 net=9456
rlabel metal2 1437 -2602 1437 -2602 0 net=10625
rlabel metal2 68 -2604 68 -2604 0 net=9921
rlabel metal2 1493 -2604 1493 -2604 0 net=11033
rlabel metal2 166 -2606 166 -2606 0 net=550
rlabel metal2 695 -2606 695 -2606 0 net=5327
rlabel metal2 884 -2606 884 -2606 0 net=6008
rlabel metal2 1010 -2606 1010 -2606 0 net=7419
rlabel metal2 1052 -2606 1052 -2606 0 net=7487
rlabel metal2 1052 -2606 1052 -2606 0 net=7487
rlabel metal2 1059 -2606 1059 -2606 0 net=8792
rlabel metal2 166 -2608 166 -2608 0 net=11740
rlabel metal2 198 -2610 198 -2610 0 net=4061
rlabel metal2 254 -2610 254 -2610 0 net=1516
rlabel metal2 296 -2610 296 -2610 0 net=2263
rlabel metal2 1003 -2610 1003 -2610 0 net=7183
rlabel metal2 1059 -2610 1059 -2610 0 net=7011
rlabel metal2 1122 -2610 1122 -2610 0 net=3700
rlabel metal2 1227 -2610 1227 -2610 0 net=8979
rlabel metal2 1276 -2610 1276 -2610 0 net=11499
rlabel metal2 65 -2612 65 -2612 0 net=7073
rlabel metal2 1066 -2612 1066 -2612 0 net=9513
rlabel metal2 1507 -2612 1507 -2612 0 net=12199
rlabel metal2 156 -2614 156 -2614 0 net=2307
rlabel metal2 373 -2614 373 -2614 0 net=3995
rlabel metal2 520 -2614 520 -2614 0 net=7350
rlabel metal2 1094 -2614 1094 -2614 0 net=7615
rlabel metal2 1276 -2614 1276 -2614 0 net=9333
rlabel metal2 1507 -2614 1507 -2614 0 net=12565
rlabel metal2 156 -2616 156 -2616 0 net=4383
rlabel metal2 520 -2616 520 -2616 0 net=3653
rlabel metal2 632 -2616 632 -2616 0 net=4853
rlabel metal2 733 -2616 733 -2616 0 net=3646
rlabel metal2 772 -2616 772 -2616 0 net=4164
rlabel metal2 957 -2616 957 -2616 0 net=12131
rlabel metal2 1283 -2616 1283 -2616 0 net=9279
rlabel metal2 1325 -2616 1325 -2616 0 net=9827
rlabel metal2 1514 -2616 1514 -2616 0 net=11175
rlabel metal2 212 -2618 212 -2618 0 net=4243
rlabel metal2 380 -2618 380 -2618 0 net=4575
rlabel metal2 464 -2618 464 -2618 0 net=2907
rlabel metal2 772 -2618 772 -2618 0 net=5869
rlabel metal2 821 -2618 821 -2618 0 net=6404
rlabel metal2 1255 -2618 1255 -2618 0 net=10115
rlabel metal2 1549 -2618 1549 -2618 0 net=11407
rlabel metal2 191 -2620 191 -2620 0 net=2393
rlabel metal2 492 -2620 492 -2620 0 net=4305
rlabel metal2 639 -2620 639 -2620 0 net=6276
rlabel metal2 716 -2620 716 -2620 0 net=7661
rlabel metal2 1122 -2620 1122 -2620 0 net=8125
rlabel metal2 1157 -2620 1157 -2620 0 net=8255
rlabel metal2 1255 -2620 1255 -2620 0 net=9141
rlabel metal2 1318 -2620 1318 -2620 0 net=9673
rlabel metal2 1612 -2620 1612 -2620 0 net=11745
rlabel metal2 184 -2622 184 -2622 0 net=3227
rlabel metal2 254 -2622 254 -2622 0 net=1701
rlabel metal2 261 -2622 261 -2622 0 net=1657
rlabel metal2 282 -2622 282 -2622 0 net=3113
rlabel metal2 646 -2622 646 -2622 0 net=6469
rlabel metal2 1199 -2622 1199 -2622 0 net=9887
rlabel metal2 142 -2624 142 -2624 0 net=1975
rlabel metal2 275 -2624 275 -2624 0 net=4459
rlabel metal2 418 -2624 418 -2624 0 net=5411
rlabel metal2 660 -2624 660 -2624 0 net=5564
rlabel metal2 821 -2624 821 -2624 0 net=5917
rlabel metal2 884 -2624 884 -2624 0 net=6319
rlabel metal2 957 -2624 957 -2624 0 net=11409
rlabel metal2 107 -2626 107 -2626 0 net=4214
rlabel metal2 457 -2626 457 -2626 0 net=2179
rlabel metal2 569 -2626 569 -2626 0 net=6041
rlabel metal2 894 -2626 894 -2626 0 net=11225
rlabel metal2 107 -2628 107 -2628 0 net=2463
rlabel metal2 310 -2628 310 -2628 0 net=2460
rlabel metal2 471 -2628 471 -2628 0 net=4335
rlabel metal2 744 -2628 744 -2628 0 net=5557
rlabel metal2 779 -2628 779 -2628 0 net=5443
rlabel metal2 933 -2628 933 -2628 0 net=6529
rlabel metal2 989 -2628 989 -2628 0 net=8415
rlabel metal2 1199 -2628 1199 -2628 0 net=8619
rlabel metal2 1269 -2628 1269 -2628 0 net=9047
rlabel metal2 72 -2630 72 -2630 0 net=4777
rlabel metal2 803 -2630 803 -2630 0 net=1242
rlabel metal2 1024 -2630 1024 -2630 0 net=8075
rlabel metal2 1150 -2630 1150 -2630 0 net=5797
rlabel metal2 142 -2632 142 -2632 0 net=1819
rlabel metal2 747 -2632 747 -2632 0 net=12297
rlabel metal2 177 -2634 177 -2634 0 net=3343
rlabel metal2 485 -2634 485 -2634 0 net=4599
rlabel metal2 653 -2634 653 -2634 0 net=2996
rlabel metal2 751 -2634 751 -2634 0 net=10874
rlabel metal2 1556 -2634 1556 -2634 0 net=11107
rlabel metal2 51 -2636 51 -2636 0 net=4771
rlabel metal2 205 -2636 205 -2636 0 net=1869
rlabel metal2 317 -2636 317 -2636 0 net=7353
rlabel metal2 751 -2636 751 -2636 0 net=8345
rlabel metal2 1157 -2636 1157 -2636 0 net=8405
rlabel metal2 1206 -2636 1206 -2636 0 net=8799
rlabel metal2 1269 -2636 1269 -2636 0 net=9263
rlabel metal2 1486 -2636 1486 -2636 0 net=12343
rlabel metal2 51 -2638 51 -2638 0 net=5519
rlabel metal2 597 -2638 597 -2638 0 net=5595
rlabel metal2 807 -2638 807 -2638 0 net=5943
rlabel metal2 947 -2638 947 -2638 0 net=6777
rlabel metal2 982 -2638 982 -2638 0 net=8433
rlabel metal2 1297 -2638 1297 -2638 0 net=9845
rlabel metal2 1556 -2638 1556 -2638 0 net=11439
rlabel metal2 121 -2640 121 -2640 0 net=6157
rlabel metal2 625 -2640 625 -2640 0 net=11801
rlabel metal2 247 -2642 247 -2642 0 net=2069
rlabel metal2 317 -2642 317 -2642 0 net=2839
rlabel metal2 534 -2642 534 -2642 0 net=4913
rlabel metal2 702 -2642 702 -2642 0 net=6963
rlabel metal2 1017 -2642 1017 -2642 0 net=7267
rlabel metal2 1062 -2642 1062 -2642 0 net=11611
rlabel metal2 86 -2644 86 -2644 0 net=5095
rlabel metal2 737 -2644 737 -2644 0 net=10669
rlabel metal2 86 -2646 86 -2646 0 net=12252
rlabel metal2 289 -2648 289 -2648 0 net=3613
rlabel metal2 534 -2648 534 -2648 0 net=3823
rlabel metal2 1017 -2648 1017 -2648 0 net=7373
rlabel metal2 1094 -2648 1094 -2648 0 net=8987
rlabel metal2 1290 -2648 1290 -2648 0 net=10341
rlabel metal2 338 -2650 338 -2650 0 net=3309
rlabel metal2 411 -2650 411 -2650 0 net=3465
rlabel metal2 541 -2650 541 -2650 0 net=6621
rlabel metal2 1031 -2650 1031 -2650 0 net=9985
rlabel metal2 219 -2652 219 -2652 0 net=5113
rlabel metal2 345 -2652 345 -2652 0 net=2133
rlabel metal2 737 -2652 737 -2652 0 net=6085
rlabel metal2 1097 -2652 1097 -2652 0 net=8840
rlabel metal2 82 -2654 82 -2654 0 net=4885
rlabel metal2 450 -2654 450 -2654 0 net=8905
rlabel metal2 1290 -2654 1290 -2654 0 net=9501
rlabel metal2 1472 -2654 1472 -2654 0 net=10881
rlabel metal2 628 -2656 628 -2656 0 net=6643
rlabel metal2 1101 -2656 1101 -2656 0 net=7731
rlabel metal2 1311 -2656 1311 -2656 0 net=9795
rlabel metal2 1535 -2656 1535 -2656 0 net=11389
rlabel metal2 443 -2658 443 -2658 0 net=11719
rlabel metal2 331 -2660 331 -2660 0 net=2925
rlabel metal2 709 -2660 709 -2660 0 net=5887
rlabel metal2 754 -2660 754 -2660 0 net=11605
rlabel metal2 331 -2662 331 -2662 0 net=3021
rlabel metal2 723 -2662 723 -2662 0 net=5155
rlabel metal2 863 -2662 863 -2662 0 net=7439
rlabel metal2 1115 -2662 1115 -2662 0 net=8105
rlabel metal2 1332 -2662 1332 -2662 0 net=9833
rlabel metal2 114 -2664 114 -2664 0 net=6325
rlabel metal2 366 -2664 366 -2664 0 net=2879
rlabel metal2 1073 -2664 1073 -2664 0 net=8233
rlabel metal2 1367 -2664 1367 -2664 0 net=10007
rlabel metal2 366 -2666 366 -2666 0 net=3863
rlabel metal2 768 -2666 768 -2666 0 net=7585
rlabel metal2 1388 -2666 1388 -2666 0 net=10279
rlabel metal2 415 -2668 415 -2668 0 net=4315
rlabel metal2 877 -2668 877 -2668 0 net=6367
rlabel metal2 1409 -2668 1409 -2668 0 net=10359
rlabel metal2 513 -2670 513 -2670 0 net=3883
rlabel metal2 912 -2670 912 -2670 0 net=6517
rlabel metal2 1465 -2670 1465 -2670 0 net=10797
rlabel metal2 740 -2672 740 -2672 0 net=11037
rlabel metal2 1528 -2672 1528 -2672 0 net=11369
rlabel metal2 919 -2674 919 -2674 0 net=6533
rlabel metal2 1444 -2674 1444 -2674 0 net=11645
rlabel metal2 870 -2676 870 -2676 0 net=10649
rlabel metal2 688 -2678 688 -2678 0 net=3612
rlabel metal2 968 -2678 968 -2678 0 net=6941
rlabel metal2 618 -2680 618 -2680 0 net=4453
rlabel metal2 677 -2682 677 -2682 0 net=7451
rlabel metal2 37 -2693 37 -2693 0 net=4337
rlabel metal2 579 -2693 579 -2693 0 net=5618
rlabel metal2 803 -2693 803 -2693 0 net=10258
rlabel metal2 51 -2695 51 -2695 0 net=5520
rlabel metal2 926 -2695 926 -2695 0 net=6524
rlabel metal2 1395 -2695 1395 -2695 0 net=12345
rlabel metal2 51 -2697 51 -2697 0 net=4245
rlabel metal2 250 -2697 250 -2697 0 net=5096
rlabel metal2 733 -2697 733 -2697 0 net=9514
rlabel metal2 1094 -2697 1094 -2697 0 net=12580
rlabel metal2 58 -2699 58 -2699 0 net=2050
rlabel metal2 649 -2699 649 -2699 0 net=3558
rlabel metal2 954 -2699 954 -2699 0 net=7616
rlabel metal2 1486 -2699 1486 -2699 0 net=12649
rlabel metal2 58 -2701 58 -2701 0 net=2061
rlabel metal2 250 -2701 250 -2701 0 net=4854
rlabel metal2 660 -2701 660 -2701 0 net=7355
rlabel metal2 758 -2701 758 -2701 0 net=2908
rlabel metal2 1066 -2701 1066 -2701 0 net=8127
rlabel metal2 1241 -2701 1241 -2701 0 net=9503
rlabel metal2 65 -2703 65 -2703 0 net=4914
rlabel metal2 660 -2703 660 -2703 0 net=6075
rlabel metal2 674 -2703 674 -2703 0 net=9846
rlabel metal2 65 -2705 65 -2705 0 net=5661
rlabel metal2 954 -2705 954 -2705 0 net=7733
rlabel metal2 1290 -2705 1290 -2705 0 net=10515
rlabel metal2 68 -2707 68 -2707 0 net=2880
rlabel metal2 1094 -2707 1094 -2707 0 net=10670
rlabel metal2 72 -2709 72 -2709 0 net=4778
rlabel metal2 453 -2709 453 -2709 0 net=3654
rlabel metal2 523 -2709 523 -2709 0 net=8526
rlabel metal2 1297 -2709 1297 -2709 0 net=10441
rlabel metal2 1430 -2709 1430 -2709 0 net=11441
rlabel metal2 82 -2711 82 -2711 0 net=5546
rlabel metal2 793 -2711 793 -2711 0 net=6645
rlabel metal2 957 -2711 957 -2711 0 net=11408
rlabel metal2 1556 -2711 1556 -2711 0 net=11607
rlabel metal2 110 -2713 110 -2713 0 net=9280
rlabel metal2 1416 -2713 1416 -2713 0 net=11803
rlabel metal2 114 -2715 114 -2715 0 net=6674
rlabel metal2 583 -2715 583 -2715 0 net=4316
rlabel metal2 1549 -2715 1549 -2715 0 net=11647
rlabel metal2 114 -2717 114 -2717 0 net=4601
rlabel metal2 653 -2717 653 -2717 0 net=10763
rlabel metal2 1283 -2717 1283 -2717 0 net=10499
rlabel metal2 117 -2719 117 -2719 0 net=4454
rlabel metal2 625 -2719 625 -2719 0 net=6320
rlabel metal2 947 -2719 947 -2719 0 net=5799
rlabel metal2 1423 -2719 1423 -2719 0 net=11919
rlabel metal2 121 -2721 121 -2721 0 net=6158
rlabel metal2 814 -2721 814 -2721 0 net=5444
rlabel metal2 849 -2721 849 -2721 0 net=7075
rlabel metal2 1034 -2721 1034 -2721 0 net=10116
rlabel metal2 121 -2723 121 -2723 0 net=3087
rlabel metal2 275 -2723 275 -2723 0 net=4461
rlabel metal2 289 -2723 289 -2723 0 net=3615
rlabel metal2 481 -2723 481 -2723 0 net=4306
rlabel metal2 583 -2723 583 -2723 0 net=6965
rlabel metal2 989 -2723 989 -2723 0 net=11024
rlabel metal2 107 -2725 107 -2725 0 net=2465
rlabel metal2 331 -2725 331 -2725 0 net=3022
rlabel metal2 786 -2725 786 -2725 0 net=6579
rlabel metal2 989 -2725 989 -2725 0 net=8981
rlabel metal2 1381 -2725 1381 -2725 0 net=11747
rlabel metal2 86 -2727 86 -2727 0 net=623
rlabel metal2 128 -2727 128 -2727 0 net=5966
rlabel metal2 758 -2727 758 -2727 0 net=6530
rlabel metal2 940 -2727 940 -2727 0 net=8155
rlabel metal2 1150 -2727 1150 -2727 0 net=9335
rlabel metal2 86 -2729 86 -2729 0 net=11108
rlabel metal2 93 -2731 93 -2731 0 net=4452
rlabel metal2 142 -2731 142 -2731 0 net=1820
rlabel metal2 688 -2731 688 -2731 0 net=8620
rlabel metal2 1227 -2731 1227 -2731 0 net=10361
rlabel metal2 72 -2733 72 -2733 0 net=6455
rlabel metal2 149 -2733 149 -2733 0 net=2151
rlabel metal2 166 -2733 166 -2733 0 net=6823
rlabel metal2 352 -2733 352 -2733 0 net=6327
rlabel metal2 667 -2733 667 -2733 0 net=4482
rlabel metal2 765 -2733 765 -2733 0 net=8536
rlabel metal2 1199 -2733 1199 -2733 0 net=9829
rlabel metal2 89 -2735 89 -2735 0 net=6675
rlabel metal2 149 -2735 149 -2735 0 net=9575
rlabel metal2 201 -2735 201 -2735 0 net=732
rlabel metal2 814 -2735 814 -2735 0 net=7441
rlabel metal2 873 -2735 873 -2735 0 net=10915
rlabel metal2 1192 -2735 1192 -2735 0 net=9889
rlabel metal2 89 -2737 89 -2737 0 net=5114
rlabel metal2 373 -2737 373 -2737 0 net=3996
rlabel metal2 429 -2737 429 -2737 0 net=5218
rlabel metal2 835 -2737 835 -2737 0 net=6350
rlabel metal2 933 -2737 933 -2737 0 net=7587
rlabel metal2 1101 -2737 1101 -2737 0 net=9797
rlabel metal2 1325 -2737 1325 -2737 0 net=11163
rlabel metal2 166 -2739 166 -2739 0 net=4663
rlabel metal2 593 -2739 593 -2739 0 net=266
rlabel metal2 1311 -2739 1311 -2739 0 net=11721
rlabel metal2 180 -2741 180 -2741 0 net=9048
rlabel metal2 184 -2743 184 -2743 0 net=1977
rlabel metal2 205 -2743 205 -2743 0 net=1871
rlabel metal2 359 -2743 359 -2743 0 net=2395
rlabel metal2 380 -2743 380 -2743 0 net=4576
rlabel metal2 380 -2743 380 -2743 0 net=4576
rlabel metal2 387 -2743 387 -2743 0 net=3311
rlabel metal2 387 -2743 387 -2743 0 net=3311
rlabel metal2 401 -2743 401 -2743 0 net=5183
rlabel metal2 597 -2743 597 -2743 0 net=12542
rlabel metal2 156 -2745 156 -2745 0 net=4385
rlabel metal2 212 -2745 212 -2745 0 net=2969
rlabel metal2 240 -2745 240 -2745 0 net=1659
rlabel metal2 268 -2745 268 -2745 0 net=2203
rlabel metal2 359 -2745 359 -2745 0 net=3467
rlabel metal2 506 -2745 506 -2745 0 net=6057
rlabel metal2 667 -2745 667 -2745 0 net=7375
rlabel metal2 1045 -2745 1045 -2745 0 net=11536
rlabel metal2 44 -2747 44 -2747 0 net=8868
rlabel metal2 254 -2747 254 -2747 0 net=1703
rlabel metal2 268 -2747 268 -2747 0 net=1597
rlabel metal2 485 -2747 485 -2747 0 net=5157
rlabel metal2 730 -2747 730 -2747 0 net=6287
rlabel metal2 863 -2747 863 -2747 0 net=6853
rlabel metal2 1339 -2747 1339 -2747 0 net=11411
rlabel metal2 44 -2749 44 -2749 0 net=2099
rlabel metal2 131 -2749 131 -2749 0 net=10487
rlabel metal2 835 -2749 835 -2749 0 net=7453
rlabel metal2 1003 -2749 1003 -2749 0 net=8235
rlabel metal2 1374 -2749 1374 -2749 0 net=10147
rlabel metal2 96 -2751 96 -2751 0 net=5489
rlabel metal2 184 -2751 184 -2751 0 net=3229
rlabel metal2 254 -2751 254 -2751 0 net=2537
rlabel metal2 401 -2751 401 -2751 0 net=3421
rlabel metal2 450 -2751 450 -2751 0 net=806
rlabel metal2 1017 -2751 1017 -2751 0 net=8435
rlabel metal2 1374 -2751 1374 -2751 0 net=10627
rlabel metal2 1458 -2751 1458 -2751 0 net=12385
rlabel metal2 100 -2753 100 -2753 0 net=3115
rlabel metal2 345 -2753 345 -2753 0 net=2134
rlabel metal2 1073 -2753 1073 -2753 0 net=9143
rlabel metal2 1437 -2753 1437 -2753 0 net=11461
rlabel metal2 275 -2755 275 -2755 0 net=2231
rlabel metal2 345 -2755 345 -2755 0 net=2181
rlabel metal2 520 -2755 520 -2755 0 net=7283
rlabel metal2 716 -2755 716 -2755 0 net=7663
rlabel metal2 884 -2755 884 -2755 0 net=11727
rlabel metal2 1458 -2755 1458 -2755 0 net=12357
rlabel metal2 233 -2757 233 -2757 0 net=4063
rlabel metal2 534 -2757 534 -2757 0 net=3824
rlabel metal2 1136 -2757 1136 -2757 0 net=9265
rlabel metal2 177 -2759 177 -2759 0 net=4773
rlabel metal2 282 -2759 282 -2759 0 net=3243
rlabel metal2 457 -2759 457 -2759 0 net=7329
rlabel metal2 229 -2761 229 -2761 0 net=9627
rlabel metal2 534 -2761 534 -2761 0 net=6923
rlabel metal2 1031 -2761 1031 -2761 0 net=9113
rlabel metal2 1171 -2761 1171 -2761 0 net=9987
rlabel metal2 317 -2763 317 -2763 0 net=2841
rlabel metal2 366 -2763 366 -2763 0 net=3865
rlabel metal2 541 -2763 541 -2763 0 net=6622
rlabel metal2 898 -2763 898 -2763 0 net=9077
rlabel metal2 975 -2763 975 -2763 0 net=7489
rlabel metal2 1269 -2763 1269 -2763 0 net=10719
rlabel metal2 296 -2765 296 -2765 0 net=2309
rlabel metal2 408 -2765 408 -2765 0 net=6543
rlabel metal2 1360 -2765 1360 -2765 0 net=11613
rlabel metal2 296 -2767 296 -2767 0 net=1931
rlabel metal2 429 -2767 429 -2767 0 net=4831
rlabel metal2 618 -2767 618 -2767 0 net=8077
rlabel metal2 1451 -2767 1451 -2767 0 net=12201
rlabel metal2 317 -2769 317 -2769 0 net=2927
rlabel metal2 499 -2769 499 -2769 0 net=5413
rlabel metal2 625 -2769 625 -2769 0 net=5889
rlabel metal2 716 -2769 716 -2769 0 net=9099
rlabel metal2 870 -2769 870 -2769 0 net=10963
rlabel metal2 1108 -2769 1108 -2769 0 net=9197
rlabel metal2 278 -2771 278 -2771 0 net=1
rlabel metal2 499 -2771 499 -2771 0 net=5559
rlabel metal2 751 -2771 751 -2771 0 net=5871
rlabel metal2 870 -2771 870 -2771 0 net=8417
rlabel metal2 1262 -2771 1262 -2771 0 net=10883
rlabel metal2 411 -2773 411 -2773 0 net=3788
rlabel metal2 541 -2773 541 -2773 0 net=4543
rlabel metal2 597 -2773 597 -2773 0 net=6535
rlabel metal2 1052 -2773 1052 -2773 0 net=9835
rlabel metal2 1472 -2773 1472 -2773 0 net=12567
rlabel metal2 415 -2775 415 -2775 0 net=2855
rlabel metal2 709 -2775 709 -2775 0 net=6369
rlabel metal2 894 -2775 894 -2775 0 net=12460
rlabel metal2 247 -2777 247 -2777 0 net=12285
rlabel metal2 919 -2777 919 -2777 0 net=8907
rlabel metal2 1332 -2777 1332 -2777 0 net=11391
rlabel metal2 422 -2779 422 -2779 0 net=8203
rlabel metal2 1164 -2779 1164 -2779 0 net=10009
rlabel metal2 1493 -2779 1493 -2779 0 net=11034
rlabel metal2 436 -2781 436 -2781 0 net=5993
rlabel metal2 555 -2781 555 -2781 0 net=5945
rlabel metal2 1213 -2781 1213 -2781 0 net=10651
rlabel metal2 1493 -2781 1493 -2781 0 net=12299
rlabel metal2 219 -2783 219 -2783 0 net=4887
rlabel metal2 562 -2783 562 -2783 0 net=5597
rlabel metal2 807 -2783 807 -2783 0 net=6779
rlabel metal2 1248 -2783 1248 -2783 0 net=12133
rlabel metal2 170 -2785 170 -2785 0 net=5149
rlabel metal2 527 -2785 527 -2785 0 net=4539
rlabel metal2 1206 -2785 1206 -2785 0 net=8801
rlabel metal2 1346 -2785 1346 -2785 0 net=9647
rlabel metal2 170 -2787 170 -2787 0 net=4165
rlabel metal2 842 -2787 842 -2787 0 net=11067
rlabel metal2 1346 -2787 1346 -2787 0 net=11177
rlabel metal2 79 -2789 79 -2789 0 net=446
rlabel metal2 79 -2791 79 -2791 0 net=2403
rlabel metal2 590 -2791 590 -2791 0 net=5918
rlabel metal2 842 -2791 842 -2791 0 net=6519
rlabel metal2 961 -2791 961 -2791 0 net=8107
rlabel metal2 1367 -2791 1367 -2791 0 net=10281
rlabel metal2 394 -2793 394 -2793 0 net=3345
rlabel metal2 600 -2793 600 -2793 0 net=6086
rlabel metal2 744 -2793 744 -2793 0 net=6043
rlabel metal2 912 -2793 912 -2793 0 net=6943
rlabel metal2 1115 -2793 1115 -2793 0 net=11753
rlabel metal2 135 -2795 135 -2795 0 net=2771
rlabel metal2 674 -2795 674 -2795 0 net=7717
rlabel metal2 135 -2797 135 -2797 0 net=6471
rlabel metal2 681 -2797 681 -2797 0 net=9674
rlabel metal2 464 -2799 464 -2799 0 net=7877
rlabel metal2 761 -2799 761 -2799 0 net=8753
rlabel metal2 821 -2799 821 -2799 0 net=7185
rlabel metal2 1318 -2799 1318 -2799 0 net=11039
rlabel metal2 163 -2801 163 -2801 0 net=11383
rlabel metal2 163 -2803 163 -2803 0 net=2264
rlabel metal2 999 -2803 999 -2803 0 net=9975
rlabel metal2 310 -2805 310 -2805 0 net=2071
rlabel metal2 765 -2805 765 -2805 0 net=10607
rlabel metal2 303 -2807 303 -2807 0 net=2025
rlabel metal2 768 -2807 768 -2807 0 net=7268
rlabel metal2 303 -2809 303 -2809 0 net=3885
rlabel metal2 772 -2809 772 -2809 0 net=9205
rlabel metal2 838 -2809 838 -2809 0 net=9367
rlabel metal2 1024 -2809 1024 -2809 0 net=8407
rlabel metal2 513 -2811 513 -2811 0 net=4413
rlabel metal2 891 -2811 891 -2811 0 net=8861
rlabel metal2 1157 -2811 1157 -2811 0 net=8725
rlabel metal2 604 -2813 604 -2813 0 net=5329
rlabel metal2 1178 -2813 1178 -2813 0 net=8257
rlabel metal2 695 -2815 695 -2815 0 net=7421
rlabel metal2 1220 -2815 1220 -2815 0 net=10799
rlabel metal2 1038 -2817 1038 -2817 0 net=7013
rlabel metal2 1465 -2817 1465 -2817 0 net=11227
rlabel metal2 1059 -2819 1059 -2819 0 net=9923
rlabel metal2 1304 -2821 1304 -2821 0 net=7505
rlabel metal2 1234 -2823 1234 -2823 0 net=8989
rlabel metal2 1353 -2823 1353 -2823 0 net=11501
rlabel metal2 1234 -2825 1234 -2825 0 net=10343
rlabel metal2 1402 -2827 1402 -2827 0 net=11371
rlabel metal2 1143 -2829 1143 -2829 0 net=8347
rlabel metal2 1143 -2831 1143 -2831 0 net=9319
rlabel metal2 30 -2842 30 -2842 0 net=9629
rlabel metal2 506 -2842 506 -2842 0 net=3866
rlabel metal2 765 -2842 765 -2842 0 net=6520
rlabel metal2 887 -2842 887 -2842 0 net=443
rlabel metal2 982 -2842 982 -2842 0 net=11372
rlabel metal2 1514 -2842 1514 -2842 0 net=11608
rlabel metal2 37 -2844 37 -2844 0 net=4338
rlabel metal2 583 -2844 583 -2844 0 net=6966
rlabel metal2 702 -2844 702 -2844 0 net=7357
rlabel metal2 898 -2844 898 -2844 0 net=10628
rlabel metal2 1395 -2844 1395 -2844 0 net=12347
rlabel metal2 37 -2846 37 -2846 0 net=5561
rlabel metal2 569 -2846 569 -2846 0 net=5185
rlabel metal2 593 -2846 593 -2846 0 net=6646
rlabel metal2 803 -2846 803 -2846 0 net=8108
rlabel metal2 996 -2846 996 -2846 0 net=9890
rlabel metal2 1202 -2846 1202 -2846 0 net=10282
rlabel metal2 44 -2848 44 -2848 0 net=2100
rlabel metal2 121 -2848 121 -2848 0 net=3088
rlabel metal2 607 -2848 607 -2848 0 net=6547
rlabel metal2 751 -2848 751 -2848 0 net=5873
rlabel metal2 775 -2848 775 -2848 0 net=9830
rlabel metal2 1276 -2848 1276 -2848 0 net=11393
rlabel metal2 1367 -2848 1367 -2848 0 net=11755
rlabel metal2 51 -2850 51 -2850 0 net=4246
rlabel metal2 250 -2850 250 -2850 0 net=11797
rlabel metal2 1388 -2850 1388 -2850 0 net=12135
rlabel metal2 51 -2852 51 -2852 0 net=5891
rlabel metal2 653 -2852 653 -2852 0 net=9207
rlabel metal2 877 -2852 877 -2852 0 net=12287
rlabel metal2 72 -2854 72 -2854 0 net=6456
rlabel metal2 1118 -2854 1118 -2854 0 net=12386
rlabel metal2 75 -2856 75 -2856 0 net=4540
rlabel metal2 618 -2856 618 -2856 0 net=8078
rlabel metal2 898 -2856 898 -2856 0 net=5297
rlabel metal2 86 -2858 86 -2858 0 net=3887
rlabel metal2 345 -2858 345 -2858 0 net=2182
rlabel metal2 751 -2858 751 -2858 0 net=6581
rlabel metal2 807 -2858 807 -2858 0 net=6780
rlabel metal2 947 -2858 947 -2858 0 net=5801
rlabel metal2 996 -2858 996 -2858 0 net=8128
rlabel metal2 1097 -2858 1097 -2858 0 net=11462
rlabel metal2 1500 -2858 1500 -2858 0 net=11649
rlabel metal2 93 -2860 93 -2860 0 net=1466
rlabel metal2 121 -2860 121 -2860 0 net=4377
rlabel metal2 268 -2860 268 -2860 0 net=1598
rlabel metal2 821 -2860 821 -2860 0 net=7187
rlabel metal2 821 -2860 821 -2860 0 net=7187
rlabel metal2 828 -2860 828 -2860 0 net=9115
rlabel metal2 1038 -2860 1038 -2860 0 net=7015
rlabel metal2 1164 -2860 1164 -2860 0 net=10010
rlabel metal2 1188 -2860 1188 -2860 0 net=11442
rlabel metal2 93 -2862 93 -2862 0 net=5331
rlabel metal2 618 -2862 618 -2862 0 net=9101
rlabel metal2 779 -2862 779 -2862 0 net=8755
rlabel metal2 1048 -2862 1048 -2862 0 net=9266
rlabel metal2 1185 -2862 1185 -2862 0 net=11069
rlabel metal2 1279 -2862 1279 -2862 0 net=12202
rlabel metal2 96 -2864 96 -2864 0 net=6924
rlabel metal2 625 -2864 625 -2864 0 net=7285
rlabel metal2 695 -2864 695 -2864 0 net=7423
rlabel metal2 856 -2864 856 -2864 0 net=7665
rlabel metal2 905 -2864 905 -2864 0 net=9369
rlabel metal2 1192 -2864 1192 -2864 0 net=10653
rlabel metal2 1248 -2864 1248 -2864 0 net=8803
rlabel metal2 100 -2866 100 -2866 0 net=3116
rlabel metal2 226 -2866 226 -2866 0 net=1705
rlabel metal2 268 -2866 268 -2866 0 net=3347
rlabel metal2 411 -2866 411 -2866 0 net=10727
rlabel metal2 1213 -2866 1213 -2866 0 net=10501
rlabel metal2 1318 -2866 1318 -2866 0 net=11041
rlabel metal2 1430 -2866 1430 -2866 0 net=12359
rlabel metal2 100 -2868 100 -2868 0 net=5395
rlabel metal2 275 -2868 275 -2868 0 net=2233
rlabel metal2 345 -2868 345 -2868 0 net=3313
rlabel metal2 429 -2868 429 -2868 0 net=4833
rlabel metal2 576 -2868 576 -2868 0 net=4665
rlabel metal2 709 -2868 709 -2868 0 net=6371
rlabel metal2 800 -2868 800 -2868 0 net=9997
rlabel metal2 1283 -2868 1283 -2868 0 net=4483
rlabel metal2 107 -2870 107 -2870 0 net=4545
rlabel metal2 646 -2870 646 -2870 0 net=12681
rlabel metal2 1458 -2870 1458 -2870 0 net=9649
rlabel metal2 128 -2872 128 -2872 0 net=7053
rlabel metal2 800 -2872 800 -2872 0 net=7077
rlabel metal2 866 -2872 866 -2872 0 net=7431
rlabel metal2 905 -2872 905 -2872 0 net=7589
rlabel metal2 940 -2872 940 -2872 0 net=8157
rlabel metal2 1129 -2872 1129 -2872 0 net=10917
rlabel metal2 1311 -2872 1311 -2872 0 net=11723
rlabel metal2 128 -2874 128 -2874 0 net=1661
rlabel metal2 275 -2874 275 -2874 0 net=2027
rlabel metal2 359 -2874 359 -2874 0 net=3469
rlabel metal2 450 -2874 450 -2874 0 net=7330
rlabel metal2 135 -2876 135 -2876 0 net=6473
rlabel metal2 541 -2876 541 -2876 0 net=6329
rlabel metal2 646 -2876 646 -2876 0 net=8983
rlabel metal2 1003 -2876 1003 -2876 0 net=8237
rlabel metal2 1311 -2876 1311 -2876 0 net=11615
rlabel metal2 1409 -2876 1409 -2876 0 net=11921
rlabel metal2 135 -2878 135 -2878 0 net=6311
rlabel metal2 191 -2878 191 -2878 0 net=2153
rlabel metal2 331 -2878 331 -2878 0 net=6825
rlabel metal2 457 -2878 457 -2878 0 net=5481
rlabel metal2 660 -2878 660 -2878 0 net=6077
rlabel metal2 716 -2878 716 -2878 0 net=6257
rlabel metal2 779 -2878 779 -2878 0 net=6855
rlabel metal2 912 -2878 912 -2878 0 net=6944
rlabel metal2 1080 -2878 1080 -2878 0 net=9977
rlabel metal2 1360 -2878 1360 -2878 0 net=11749
rlabel metal2 1423 -2878 1423 -2878 0 net=12651
rlabel metal2 142 -2880 142 -2880 0 net=6677
rlabel metal2 863 -2880 863 -2880 0 net=9336
rlabel metal2 1381 -2880 1381 -2880 0 net=11805
rlabel metal2 1486 -2880 1486 -2880 0 net=7507
rlabel metal2 142 -2882 142 -2882 0 net=2971
rlabel metal2 219 -2882 219 -2882 0 net=5151
rlabel metal2 474 -2882 474 -2882 0 net=9723
rlabel metal2 1150 -2882 1150 -2882 0 net=10363
rlabel metal2 1416 -2882 1416 -2882 0 net=12403
rlabel metal2 72 -2884 72 -2884 0 net=3457
rlabel metal2 219 -2884 219 -2884 0 net=3133
rlabel metal2 1003 -2884 1003 -2884 0 net=9145
rlabel metal2 1080 -2884 1080 -2884 0 net=9505
rlabel metal2 170 -2886 170 -2886 0 net=4166
rlabel metal2 523 -2886 523 -2886 0 net=7927
rlabel metal2 961 -2886 961 -2886 0 net=7491
rlabel metal2 1010 -2886 1010 -2886 0 net=8863
rlabel metal2 1122 -2886 1122 -2886 0 net=10765
rlabel metal2 1241 -2886 1241 -2886 0 net=10885
rlabel metal2 170 -2888 170 -2888 0 net=2947
rlabel metal2 177 -2890 177 -2890 0 net=1617
rlabel metal2 282 -2890 282 -2890 0 net=3245
rlabel metal2 660 -2890 660 -2890 0 net=6045
rlabel metal2 870 -2890 870 -2890 0 net=8419
rlabel metal2 1087 -2890 1087 -2890 0 net=10965
rlabel metal2 163 -2892 163 -2892 0 net=9903
rlabel metal2 331 -2892 331 -2892 0 net=2311
rlabel metal2 373 -2892 373 -2892 0 net=2396
rlabel metal2 527 -2892 527 -2892 0 net=4889
rlabel metal2 555 -2892 555 -2892 0 net=5947
rlabel metal2 667 -2892 667 -2892 0 net=7377
rlabel metal2 912 -2892 912 -2892 0 net=12300
rlabel metal2 114 -2894 114 -2894 0 net=4603
rlabel metal2 548 -2894 548 -2894 0 net=5415
rlabel metal2 667 -2894 667 -2894 0 net=8035
rlabel metal2 926 -2894 926 -2894 0 net=9079
rlabel metal2 1010 -2894 1010 -2894 0 net=8259
rlabel metal2 1493 -2894 1493 -2894 0 net=8349
rlabel metal2 163 -2896 163 -2896 0 net=3007
rlabel metal2 250 -2896 250 -2896 0 net=7449
rlabel metal2 926 -2896 926 -2896 0 net=8990
rlabel metal2 191 -2898 191 -2898 0 net=4387
rlabel metal2 359 -2898 359 -2898 0 net=6199
rlabel metal2 975 -2898 975 -2898 0 net=8727
rlabel metal2 1178 -2898 1178 -2898 0 net=10517
rlabel metal2 1304 -2898 1304 -2898 0 net=11503
rlabel metal2 205 -2900 205 -2900 0 net=2539
rlabel metal2 366 -2900 366 -2900 0 net=2823
rlabel metal2 674 -2900 674 -2900 0 net=7718
rlabel metal2 737 -2900 737 -2900 0 net=7879
rlabel metal2 968 -2900 968 -2900 0 net=10609
rlabel metal2 254 -2902 254 -2902 0 net=1872
rlabel metal2 380 -2902 380 -2902 0 net=4729
rlabel metal2 485 -2902 485 -2902 0 net=5159
rlabel metal2 597 -2902 597 -2902 0 net=6537
rlabel metal2 761 -2902 761 -2902 0 net=9491
rlabel metal2 1027 -2902 1027 -2902 0 net=11384
rlabel metal2 289 -2904 289 -2904 0 net=2467
rlabel metal2 380 -2904 380 -2904 0 net=3617
rlabel metal2 485 -2904 485 -2904 0 net=5599
rlabel metal2 611 -2904 611 -2904 0 net=7443
rlabel metal2 1052 -2904 1052 -2904 0 net=9837
rlabel metal2 1157 -2904 1157 -2904 0 net=11413
rlabel metal2 1479 -2904 1479 -2904 0 net=10149
rlabel metal2 44 -2906 44 -2906 0 net=4753
rlabel metal2 761 -2906 761 -2906 0 net=7987
rlabel metal2 1052 -2906 1052 -2906 0 net=9799
rlabel metal2 1255 -2906 1255 -2906 0 net=11729
rlabel metal2 65 -2908 65 -2908 0 net=5663
rlabel metal2 408 -2908 408 -2908 0 net=6545
rlabel metal2 814 -2908 814 -2908 0 net=7455
rlabel metal2 1059 -2908 1059 -2908 0 net=9925
rlabel metal2 1101 -2908 1101 -2908 0 net=9321
rlabel metal2 1255 -2908 1255 -2908 0 net=10443
rlabel metal2 65 -2910 65 -2910 0 net=2857
rlabel metal2 436 -2910 436 -2910 0 net=5995
rlabel metal2 733 -2910 733 -2910 0 net=11401
rlabel metal2 110 -2912 110 -2912 0 net=7225
rlabel metal2 1059 -2912 1059 -2912 0 net=9199
rlabel metal2 1143 -2912 1143 -2912 0 net=9989
rlabel metal2 1290 -2912 1290 -2912 0 net=11179
rlabel metal2 401 -2914 401 -2914 0 net=3423
rlabel metal2 436 -2914 436 -2914 0 net=4065
rlabel metal2 555 -2914 555 -2914 0 net=8909
rlabel metal2 1171 -2914 1171 -2914 0 net=10345
rlabel metal2 58 -2916 58 -2916 0 net=2062
rlabel metal2 408 -2916 408 -2916 0 net=2072
rlabel metal2 478 -2916 478 -2916 0 net=245
rlabel metal2 919 -2916 919 -2916 0 net=7735
rlabel metal2 1220 -2916 1220 -2916 0 net=10801
rlabel metal2 58 -2918 58 -2918 0 net=6059
rlabel metal2 723 -2918 723 -2918 0 net=10489
rlabel metal2 1220 -2918 1220 -2918 0 net=10721
rlabel metal2 114 -2920 114 -2920 0 net=1054
rlabel metal2 723 -2920 723 -2920 0 net=6289
rlabel metal2 891 -2920 891 -2920 0 net=12729
rlabel metal2 149 -2922 149 -2922 0 net=9577
rlabel metal2 954 -2922 954 -2922 0 net=8437
rlabel metal2 1269 -2922 1269 -2922 0 net=11165
rlabel metal2 149 -2924 149 -2924 0 net=3231
rlabel metal2 317 -2924 317 -2924 0 net=2929
rlabel metal2 471 -2924 471 -2924 0 net=2772
rlabel metal2 1017 -2924 1017 -2924 0 net=8408
rlabel metal2 184 -2926 184 -2926 0 net=1979
rlabel metal2 257 -2926 257 -2926 0 net=5225
rlabel metal2 404 -2926 404 -2926 0 net=9605
rlabel metal2 198 -2928 198 -2928 0 net=1933
rlabel metal2 422 -2928 422 -2928 0 net=8205
rlabel metal2 1024 -2928 1024 -2928 0 net=11228
rlabel metal2 79 -2930 79 -2930 0 net=2405
rlabel metal2 422 -2930 422 -2930 0 net=2705
rlabel metal2 1465 -2930 1465 -2930 0 net=12569
rlabel metal2 79 -2932 79 -2932 0 net=2843
rlabel metal2 471 -2932 471 -2932 0 net=7571
rlabel metal2 233 -2934 233 -2934 0 net=4775
rlabel metal2 233 -2936 233 -2936 0 net=2205
rlabel metal2 352 -2938 352 -2938 0 net=4415
rlabel metal2 443 -2940 443 -2940 0 net=4463
rlabel metal2 156 -2942 156 -2942 0 net=5491
rlabel metal2 30 -2953 30 -2953 0 net=9631
rlabel metal2 79 -2953 79 -2953 0 net=2844
rlabel metal2 523 -2953 523 -2953 0 net=716
rlabel metal2 635 -2953 635 -2953 0 net=9492
rlabel metal2 982 -2953 982 -2953 0 net=5802
rlabel metal2 1038 -2953 1038 -2953 0 net=8757
rlabel metal2 1062 -2953 1062 -2953 0 net=12360
rlabel metal2 1444 -2953 1444 -2953 0 net=7508
rlabel metal2 37 -2955 37 -2955 0 net=5562
rlabel metal2 100 -2955 100 -2955 0 net=5396
rlabel metal2 758 -2955 758 -2955 0 net=5874
rlabel metal2 821 -2955 821 -2955 0 net=7189
rlabel metal2 821 -2955 821 -2955 0 net=7189
rlabel metal2 828 -2955 828 -2955 0 net=9116
rlabel metal2 870 -2955 870 -2955 0 net=7450
rlabel metal2 1020 -2955 1020 -2955 0 net=10364
rlabel metal2 1199 -2955 1199 -2955 0 net=11395
rlabel metal2 1447 -2955 1447 -2955 0 net=11650
rlabel metal2 37 -2957 37 -2957 0 net=4379
rlabel metal2 124 -2957 124 -2957 0 net=2154
rlabel metal2 366 -2957 366 -2957 0 net=2824
rlabel metal2 870 -2957 870 -2957 0 net=12682
rlabel metal2 1472 -2957 1472 -2957 0 net=8351
rlabel metal2 44 -2959 44 -2959 0 net=4754
rlabel metal2 254 -2959 254 -2959 0 net=4776
rlabel metal2 373 -2959 373 -2959 0 net=6826
rlabel metal2 464 -2959 464 -2959 0 net=2930
rlabel metal2 684 -2959 684 -2959 0 net=4484
rlabel metal2 44 -2961 44 -2961 0 net=3233
rlabel metal2 156 -2961 156 -2961 0 net=3619
rlabel metal2 387 -2961 387 -2961 0 net=3471
rlabel metal2 387 -2961 387 -2961 0 net=3471
rlabel metal2 429 -2961 429 -2961 0 net=4730
rlabel metal2 534 -2961 534 -2961 0 net=6474
rlabel metal2 646 -2961 646 -2961 0 net=8984
rlabel metal2 936 -2961 936 -2961 0 net=7541
rlabel metal2 996 -2961 996 -2961 0 net=11070
rlabel metal2 1255 -2961 1255 -2961 0 net=10444
rlabel metal2 51 -2963 51 -2963 0 net=5892
rlabel metal2 611 -2963 611 -2963 0 net=7444
rlabel metal2 758 -2963 758 -2963 0 net=7227
rlabel metal2 877 -2963 877 -2963 0 net=7667
rlabel metal2 1038 -2963 1038 -2963 0 net=9839
rlabel metal2 1143 -2963 1143 -2963 0 net=9991
rlabel metal2 1255 -2963 1255 -2963 0 net=12289
rlabel metal2 51 -2965 51 -2965 0 net=10253
rlabel metal2 429 -2965 429 -2965 0 net=1755
rlabel metal2 828 -2965 828 -2965 0 net=11799
rlabel metal2 65 -2967 65 -2967 0 net=2859
rlabel metal2 93 -2967 93 -2967 0 net=5332
rlabel metal2 625 -2967 625 -2967 0 net=7287
rlabel metal2 793 -2967 793 -2967 0 net=7055
rlabel metal2 905 -2967 905 -2967 0 net=7591
rlabel metal2 905 -2967 905 -2967 0 net=7591
rlabel metal2 922 -2967 922 -2967 0 net=9800
rlabel metal2 1073 -2967 1073 -2967 0 net=8421
rlabel metal2 1143 -2967 1143 -2967 0 net=10887
rlabel metal2 1276 -2967 1276 -2967 0 net=11725
rlabel metal2 1374 -2967 1374 -2967 0 net=9651
rlabel metal2 65 -2969 65 -2969 0 net=10323
rlabel metal2 254 -2969 254 -2969 0 net=2029
rlabel metal2 289 -2969 289 -2969 0 net=5665
rlabel metal2 373 -2969 373 -2969 0 net=5997
rlabel metal2 632 -2969 632 -2969 0 net=6291
rlabel metal2 933 -2969 933 -2969 0 net=9081
rlabel metal2 996 -2969 996 -2969 0 net=11042
rlabel metal2 1458 -2969 1458 -2969 0 net=12571
rlabel metal2 100 -2971 100 -2971 0 net=6331
rlabel metal2 555 -2971 555 -2971 0 net=8911
rlabel metal2 954 -2971 954 -2971 0 net=8439
rlabel metal2 1090 -2971 1090 -2971 0 net=11922
rlabel metal2 1465 -2971 1465 -2971 0 net=10151
rlabel metal2 114 -2973 114 -2973 0 net=2127
rlabel metal2 159 -2973 159 -2973 0 net=4604
rlabel metal2 527 -2973 527 -2973 0 net=4891
rlabel metal2 555 -2973 555 -2973 0 net=5073
rlabel metal2 954 -2973 954 -2973 0 net=9147
rlabel metal2 1052 -2973 1052 -2973 0 net=9979
rlabel metal2 1136 -2973 1136 -2973 0 net=8239
rlabel metal2 1332 -2973 1332 -2973 0 net=8805
rlabel metal2 114 -2975 114 -2975 0 net=6313
rlabel metal2 177 -2975 177 -2975 0 net=3753
rlabel metal2 352 -2975 352 -2975 0 net=4416
rlabel metal2 646 -2975 646 -2975 0 net=4667
rlabel metal2 723 -2975 723 -2975 0 net=9011
rlabel metal2 1003 -2975 1003 -2975 0 net=9201
rlabel metal2 1129 -2975 1129 -2975 0 net=10347
rlabel metal2 121 -2977 121 -2977 0 net=4191
rlabel metal2 177 -2977 177 -2977 0 net=9606
rlabel metal2 180 -2979 180 -2979 0 net=5152
rlabel metal2 408 -2979 408 -2979 0 net=4939
rlabel metal2 534 -2979 534 -2979 0 net=8037
rlabel metal2 912 -2979 912 -2979 0 net=8729
rlabel metal2 1080 -2979 1080 -2979 0 net=9507
rlabel metal2 198 -2981 198 -2981 0 net=1934
rlabel metal2 653 -2981 653 -2981 0 net=9209
rlabel metal2 1080 -2981 1080 -2981 0 net=10491
rlabel metal2 1136 -2981 1136 -2981 0 net=10767
rlabel metal2 201 -2983 201 -2983 0 net=4464
rlabel metal2 562 -2983 562 -2983 0 net=7079
rlabel metal2 1108 -2983 1108 -2983 0 net=11167
rlabel metal2 219 -2985 219 -2985 0 net=3135
rlabel metal2 394 -2985 394 -2985 0 net=2997
rlabel metal2 1150 -2985 1150 -2985 0 net=10967
rlabel metal2 226 -2987 226 -2987 0 net=1707
rlabel metal2 352 -2987 352 -2987 0 net=3424
rlabel metal2 422 -2987 422 -2987 0 net=2707
rlabel metal2 565 -2987 565 -2987 0 net=6546
rlabel metal2 800 -2987 800 -2987 0 net=7457
rlabel metal2 1094 -2987 1094 -2987 0 net=7017
rlabel metal2 170 -2989 170 -2989 0 net=2949
rlabel metal2 233 -2989 233 -2989 0 net=2207
rlabel metal2 355 -2989 355 -2989 0 net=9167
rlabel metal2 506 -2989 506 -2989 0 net=7573
rlabel metal2 1094 -2989 1094 -2989 0 net=10655
rlabel metal2 1213 -2989 1213 -2989 0 net=10503
rlabel metal2 128 -2991 128 -2991 0 net=1663
rlabel metal2 243 -2991 243 -2991 0 net=927
rlabel metal2 1157 -2991 1157 -2991 0 net=11415
rlabel metal2 1227 -2991 1227 -2991 0 net=11505
rlabel metal2 58 -2993 58 -2993 0 net=6061
rlabel metal2 170 -2993 170 -2993 0 net=2541
rlabel metal2 257 -2993 257 -2993 0 net=5047
rlabel metal2 443 -2993 443 -2993 0 net=5493
rlabel metal2 506 -2993 506 -2993 0 net=6259
rlabel metal2 1031 -2993 1031 -2993 0 net=8159
rlabel metal2 58 -2995 58 -2995 0 net=3009
rlabel metal2 205 -2995 205 -2995 0 net=3519
rlabel metal2 569 -2995 569 -2995 0 net=4834
rlabel metal2 691 -2995 691 -2995 0 net=9926
rlabel metal2 1157 -2995 1157 -2995 0 net=10519
rlabel metal2 1192 -2995 1192 -2995 0 net=10803
rlabel metal2 86 -2997 86 -2997 0 net=3889
rlabel metal2 450 -2997 450 -2997 0 net=5417
rlabel metal2 569 -2997 569 -2997 0 net=5187
rlabel metal2 590 -2997 590 -2997 0 net=5160
rlabel metal2 1031 -2997 1031 -2997 0 net=9371
rlabel metal2 1087 -2997 1087 -2997 0 net=8515
rlabel metal2 86 -2999 86 -2999 0 net=5675
rlabel metal2 401 -2999 401 -2999 0 net=7301
rlabel metal2 1066 -2999 1066 -2999 0 net=9323
rlabel metal2 1178 -2999 1178 -2999 0 net=11807
rlabel metal2 163 -3001 163 -3001 0 net=9103
rlabel metal2 639 -3001 639 -3001 0 net=5949
rlabel metal2 667 -3001 667 -3001 0 net=10610
rlabel metal2 1381 -3001 1381 -3001 0 net=12405
rlabel metal2 261 -3003 261 -3003 0 net=5001
rlabel metal2 590 -3003 590 -3003 0 net=5299
rlabel metal2 926 -3003 926 -3003 0 net=9551
rlabel metal2 1234 -3003 1234 -3003 0 net=11731
rlabel metal2 1416 -3003 1416 -3003 0 net=12653
rlabel metal2 142 -3005 142 -3005 0 net=2972
rlabel metal2 264 -3005 264 -3005 0 net=3348
rlabel metal2 275 -3005 275 -3005 0 net=5483
rlabel metal2 502 -3005 502 -3005 0 net=5643
rlabel metal2 597 -3005 597 -3005 0 net=7379
rlabel metal2 898 -3005 898 -3005 0 net=10011
rlabel metal2 1311 -3005 1311 -3005 0 net=11617
rlabel metal2 107 -3007 107 -3007 0 net=4547
rlabel metal2 604 -3007 604 -3007 0 net=9578
rlabel metal2 1311 -3007 1311 -3007 0 net=12137
rlabel metal2 107 -3009 107 -3009 0 net=8207
rlabel metal2 611 -3009 611 -3009 0 net=3701
rlabel metal2 142 -3011 142 -3011 0 net=1981
rlabel metal2 264 -3011 264 -3011 0 net=6678
rlabel metal2 891 -3011 891 -3011 0 net=7737
rlabel metal2 184 -3013 184 -3013 0 net=4389
rlabel metal2 268 -3013 268 -3013 0 net=2469
rlabel metal2 359 -3013 359 -3013 0 net=6201
rlabel metal2 639 -3013 639 -3013 0 net=12730
rlabel metal2 191 -3015 191 -3015 0 net=5601
rlabel metal2 492 -3015 492 -3015 0 net=6047
rlabel metal2 667 -3015 667 -3015 0 net=7929
rlabel metal2 1346 -3015 1346 -3015 0 net=12349
rlabel metal2 282 -3017 282 -3017 0 net=9905
rlabel metal2 940 -3017 940 -3017 0 net=7493
rlabel metal2 282 -3019 282 -3019 0 net=2313
rlabel metal2 338 -3019 338 -3019 0 net=3315
rlabel metal2 401 -3019 401 -3019 0 net=3427
rlabel metal2 485 -3019 485 -3019 0 net=3685
rlabel metal2 807 -3019 807 -3019 0 net=7424
rlabel metal2 296 -3021 296 -3021 0 net=2407
rlabel metal2 404 -3021 404 -3021 0 net=6155
rlabel metal2 576 -3021 576 -3021 0 net=3246
rlabel metal2 296 -3023 296 -3023 0 net=10659
rlabel metal2 317 -3025 317 -3025 0 net=5227
rlabel metal2 618 -3025 618 -3025 0 net=2887
rlabel metal2 303 -3027 303 -3027 0 net=2235
rlabel metal2 331 -3027 331 -3027 0 net=2881
rlabel metal2 660 -3027 660 -3027 0 net=6079
rlabel metal2 716 -3027 716 -3027 0 net=6857
rlabel metal2 303 -3029 303 -3029 0 net=5685
rlabel metal2 345 -3031 345 -3031 0 net=4067
rlabel metal2 471 -3031 471 -3031 0 net=4073
rlabel metal2 779 -3031 779 -3031 0 net=6373
rlabel metal2 212 -3033 212 -3033 0 net=3459
rlabel metal2 674 -3033 674 -3033 0 net=6539
rlabel metal2 786 -3033 786 -3033 0 net=8583
rlabel metal2 212 -3035 212 -3035 0 net=1619
rlabel metal2 247 -3035 247 -3035 0 net=10935
rlabel metal2 681 -3035 681 -3035 0 net=6549
rlabel metal2 411 -3037 411 -3037 0 net=6979
rlabel metal2 681 -3037 681 -3037 0 net=7432
rlabel metal2 688 -3039 688 -3039 0 net=7359
rlabel metal2 856 -3039 856 -3039 0 net=7881
rlabel metal2 695 -3041 695 -3041 0 net=6583
rlabel metal2 842 -3041 842 -3041 0 net=7989
rlabel metal2 702 -3043 702 -3043 0 net=7623
rlabel metal2 856 -3043 856 -3043 0 net=9155
rlabel metal2 705 -3045 705 -3045 0 net=11923
rlabel metal2 751 -3047 751 -3047 0 net=6925
rlabel metal2 947 -3047 947 -3047 0 net=8261
rlabel metal2 1017 -3047 1017 -3047 0 net=9725
rlabel metal2 1010 -3049 1010 -3049 0 net=8865
rlabel metal2 1115 -3049 1115 -3049 0 net=10729
rlabel metal2 1045 -3051 1045 -3051 0 net=9999
rlabel metal2 1206 -3051 1206 -3051 0 net=11757
rlabel metal2 1164 -3053 1164 -3053 0 net=10723
rlabel metal2 1220 -3055 1220 -3055 0 net=10918
rlabel metal2 1248 -3057 1248 -3057 0 net=11403
rlabel metal2 1290 -3059 1290 -3059 0 net=11181
rlabel metal2 1290 -3061 1290 -3061 0 net=11751
rlabel metal2 37 -3072 37 -3072 0 net=4380
rlabel metal2 100 -3072 100 -3072 0 net=6332
rlabel metal2 590 -3072 590 -3072 0 net=5301
rlabel metal2 590 -3072 590 -3072 0 net=5301
rlabel metal2 621 -3072 621 -3072 0 net=7302
rlabel metal2 775 -3072 775 -3072 0 net=11404
rlabel metal2 1262 -3072 1262 -3072 0 net=7018
rlabel metal2 1293 -3072 1293 -3072 0 net=11182
rlabel metal2 1339 -3072 1339 -3072 0 net=11619
rlabel metal2 1367 -3072 1367 -3072 0 net=12407
rlabel metal2 1409 -3072 1409 -3072 0 net=12655
rlabel metal2 1451 -3072 1451 -3072 0 net=12573
rlabel metal2 44 -3074 44 -3074 0 net=3234
rlabel metal2 240 -3074 240 -3074 0 net=7542
rlabel metal2 1010 -3074 1010 -3074 0 net=8866
rlabel metal2 1090 -3074 1090 -3074 0 net=10504
rlabel metal2 1283 -3074 1283 -3074 0 net=12350
rlabel metal2 1458 -3074 1458 -3074 0 net=10153
rlabel metal2 51 -3076 51 -3076 0 net=10254
rlabel metal2 226 -3076 226 -3076 0 net=2951
rlabel metal2 243 -3076 243 -3076 0 net=3316
rlabel metal2 373 -3076 373 -3076 0 net=5998
rlabel metal2 639 -3076 639 -3076 0 net=7625
rlabel metal2 849 -3076 849 -3076 0 net=8440
rlabel metal2 982 -3076 982 -3076 0 net=10731
rlabel metal2 1143 -3076 1143 -3076 0 net=10889
rlabel metal2 1143 -3076 1143 -3076 0 net=10889
rlabel metal2 1171 -3076 1171 -3076 0 net=9509
rlabel metal2 1171 -3076 1171 -3076 0 net=9509
rlabel metal2 1220 -3076 1220 -3076 0 net=11752
rlabel metal2 1346 -3076 1346 -3076 0 net=9653
rlabel metal2 1465 -3076 1465 -3076 0 net=8353
rlabel metal2 58 -3078 58 -3078 0 net=3010
rlabel metal2 191 -3078 191 -3078 0 net=5602
rlabel metal2 254 -3078 254 -3078 0 net=2031
rlabel metal2 254 -3078 254 -3078 0 net=2031
rlabel metal2 289 -3078 289 -3078 0 net=3754
rlabel metal2 653 -3078 653 -3078 0 net=5950
rlabel metal2 740 -3078 740 -3078 0 net=10907
rlabel metal2 1010 -3078 1010 -3078 0 net=9981
rlabel metal2 1059 -3078 1059 -3078 0 net=11925
rlabel metal2 1262 -3078 1262 -3078 0 net=8807
rlabel metal2 72 -3080 72 -3080 0 net=9632
rlabel metal2 191 -3080 191 -3080 0 net=2471
rlabel metal2 299 -3080 299 -3080 0 net=1708
rlabel metal2 338 -3080 338 -3080 0 net=4941
rlabel metal2 513 -3080 513 -3080 0 net=6156
rlabel metal2 744 -3080 744 -3080 0 net=7459
rlabel metal2 807 -3080 807 -3080 0 net=9157
rlabel metal2 870 -3080 870 -3080 0 net=8262
rlabel metal2 961 -3080 961 -3080 0 net=10768
rlabel metal2 1164 -3080 1164 -3080 0 net=10725
rlabel metal2 1230 -3080 1230 -3080 0 net=12138
rlabel metal2 79 -3082 79 -3082 0 net=2860
rlabel metal2 436 -3082 436 -3082 0 net=3460
rlabel metal2 1066 -3082 1066 -3082 0 net=9325
rlabel metal2 1136 -3082 1136 -3082 0 net=11733
rlabel metal2 79 -3084 79 -3084 0 net=11741
rlabel metal2 100 -3084 100 -3084 0 net=6315
rlabel metal2 121 -3084 121 -3084 0 net=7123
rlabel metal2 782 -3084 782 -3084 0 net=9840
rlabel metal2 1052 -3084 1052 -3084 0 net=12291
rlabel metal2 86 -3086 86 -3086 0 net=5676
rlabel metal2 373 -3086 373 -3086 0 net=4075
rlabel metal2 478 -3086 478 -3086 0 net=9169
rlabel metal2 873 -3086 873 -3086 0 net=7592
rlabel metal2 929 -3086 929 -3086 0 net=11726
rlabel metal2 65 -3088 65 -3088 0 net=10325
rlabel metal2 93 -3088 93 -3088 0 net=9105
rlabel metal2 177 -3088 177 -3088 0 net=6980
rlabel metal2 436 -3088 436 -3088 0 net=10629
rlabel metal2 523 -3088 523 -3088 0 net=7056
rlabel metal2 884 -3088 884 -3088 0 net=7882
rlabel metal2 933 -3088 933 -3088 0 net=9083
rlabel metal2 964 -3088 964 -3088 0 net=9992
rlabel metal2 1276 -3088 1276 -3088 0 net=8517
rlabel metal2 107 -3090 107 -3090 0 net=8209
rlabel metal2 107 -3090 107 -3090 0 net=8209
rlabel metal2 114 -3090 114 -3090 0 net=6063
rlabel metal2 142 -3090 142 -3090 0 net=1982
rlabel metal2 226 -3090 226 -3090 0 net=7049
rlabel metal2 656 -3090 656 -3090 0 net=11800
rlabel metal2 884 -3090 884 -3090 0 net=7739
rlabel metal2 905 -3090 905 -3090 0 net=6635
rlabel metal2 996 -3090 996 -3090 0 net=12607
rlabel metal2 1066 -3090 1066 -3090 0 net=10657
rlabel metal2 1101 -3090 1101 -3090 0 net=9552
rlabel metal2 121 -3092 121 -3092 0 net=3621
rlabel metal2 163 -3092 163 -3092 0 net=3521
rlabel metal2 247 -3092 247 -3092 0 net=10
rlabel metal2 366 -3092 366 -3092 0 net=5667
rlabel metal2 520 -3092 520 -3092 0 net=3703
rlabel metal2 618 -3092 618 -3092 0 net=1378
rlabel metal2 912 -3092 912 -3092 0 net=8731
rlabel metal2 940 -3092 940 -3092 0 net=7494
rlabel metal2 975 -3092 975 -3092 0 net=2889
rlabel metal2 1101 -3092 1101 -3092 0 net=11397
rlabel metal2 142 -3094 142 -3094 0 net=2543
rlabel metal2 177 -3094 177 -3094 0 net=4391
rlabel metal2 198 -3094 198 -3094 0 net=7360
rlabel metal2 702 -3094 702 -3094 0 net=8758
rlabel metal2 1129 -3094 1129 -3094 0 net=10349
rlabel metal2 149 -3096 149 -3096 0 net=2129
rlabel metal2 149 -3096 149 -3096 0 net=2129
rlabel metal2 156 -3096 156 -3096 0 net=9567
rlabel metal2 303 -3096 303 -3096 0 net=5687
rlabel metal2 527 -3096 527 -3096 0 net=2709
rlabel metal2 940 -3096 940 -3096 0 net=9149
rlabel metal2 1017 -3096 1017 -3096 0 net=9727
rlabel metal2 1017 -3096 1017 -3096 0 net=9727
rlabel metal2 1073 -3096 1073 -3096 0 net=11759
rlabel metal2 128 -3098 128 -3098 0 net=2915
rlabel metal2 366 -3098 366 -3098 0 net=2773
rlabel metal2 898 -3098 898 -3098 0 net=10013
rlabel metal2 1164 -3098 1164 -3098 0 net=2845
rlabel metal2 170 -3100 170 -3100 0 net=5485
rlabel metal2 296 -3100 296 -3100 0 net=3473
rlabel metal2 394 -3100 394 -3100 0 net=2999
rlabel metal2 464 -3100 464 -3100 0 net=4525
rlabel metal2 674 -3100 674 -3100 0 net=10937
rlabel metal2 898 -3100 898 -3100 0 net=9373
rlabel metal2 1206 -3100 1206 -3100 0 net=8161
rlabel metal2 198 -3102 198 -3102 0 net=2315
rlabel metal2 352 -3102 352 -3102 0 net=5967
rlabel metal2 684 -3102 684 -3102 0 net=9906
rlabel metal2 786 -3102 786 -3102 0 net=8585
rlabel metal2 912 -3102 912 -3102 0 net=10493
rlabel metal2 201 -3104 201 -3104 0 net=3997
rlabel metal2 352 -3104 352 -3104 0 net=1757
rlabel metal2 471 -3104 471 -3104 0 net=7381
rlabel metal2 765 -3104 765 -3104 0 net=7289
rlabel metal2 793 -3104 793 -3104 0 net=7668
rlabel metal2 1031 -3104 1031 -3104 0 net=11169
rlabel metal2 233 -3106 233 -3106 0 net=1665
rlabel metal2 261 -3106 261 -3106 0 net=6027
rlabel metal2 401 -3106 401 -3106 0 net=3428
rlabel metal2 1024 -3106 1024 -3106 0 net=8423
rlabel metal2 212 -3108 212 -3108 0 net=1621
rlabel metal2 268 -3108 268 -3108 0 net=2209
rlabel metal2 380 -3108 380 -3108 0 net=3137
rlabel metal2 387 -3108 387 -3108 0 net=7109
rlabel metal2 723 -3108 723 -3108 0 net=9013
rlabel metal2 796 -3108 796 -3108 0 net=479
rlabel metal2 1080 -3108 1080 -3108 0 net=11507
rlabel metal2 222 -3110 222 -3110 0 net=4679
rlabel metal2 408 -3110 408 -3110 0 net=3687
rlabel metal2 506 -3110 506 -3110 0 net=6261
rlabel metal2 681 -3110 681 -3110 0 net=6585
rlabel metal2 723 -3110 723 -3110 0 net=7229
rlabel metal2 835 -3110 835 -3110 0 net=10661
rlabel metal2 1108 -3110 1108 -3110 0 net=10969
rlabel metal2 233 -3112 233 -3112 0 net=2883
rlabel metal2 380 -3112 380 -3112 0 net=7557
rlabel metal2 695 -3112 695 -3112 0 net=6551
rlabel metal2 758 -3112 758 -3112 0 net=7991
rlabel metal2 1122 -3112 1122 -3112 0 net=11809
rlabel metal2 275 -3114 275 -3114 0 net=4069
rlabel metal2 485 -3114 485 -3114 0 net=1521
rlabel metal2 709 -3114 709 -3114 0 net=6541
rlabel metal2 828 -3114 828 -3114 0 net=10697
rlabel metal2 1129 -3114 1129 -3114 0 net=11637
rlabel metal2 282 -3116 282 -3116 0 net=5075
rlabel metal2 576 -3116 576 -3116 0 net=5229
rlabel metal2 835 -3116 835 -3116 0 net=8953
rlabel metal2 1150 -3116 1150 -3116 0 net=7795
rlabel metal2 289 -3118 289 -3118 0 net=3375
rlabel metal2 814 -3118 814 -3118 0 net=7575
rlabel metal2 1178 -3118 1178 -3118 0 net=10805
rlabel metal2 310 -3120 310 -3120 0 net=4549
rlabel metal2 506 -3120 506 -3120 0 net=6293
rlabel metal2 814 -3120 814 -3120 0 net=7191
rlabel metal2 1192 -3120 1192 -3120 0 net=8241
rlabel metal2 317 -3122 317 -3122 0 net=2237
rlabel metal2 345 -3122 345 -3122 0 net=2409
rlabel metal2 457 -3122 457 -3122 0 net=2159
rlabel metal2 821 -3122 821 -3122 0 net=10001
rlabel metal2 135 -3124 135 -3124 0 net=4193
rlabel metal2 527 -3124 527 -3124 0 net=6203
rlabel metal2 1045 -3124 1045 -3124 0 net=11417
rlabel metal2 205 -3126 205 -3126 0 net=9917
rlabel metal2 534 -3126 534 -3126 0 net=8038
rlabel metal2 1157 -3126 1157 -3126 0 net=10521
rlabel metal2 450 -3128 450 -3128 0 net=5419
rlabel metal2 541 -3128 541 -3128 0 net=4893
rlabel metal2 583 -3128 583 -3128 0 net=5645
rlabel metal2 1157 -3128 1157 -3128 0 net=3767
rlabel metal2 450 -3130 450 -3130 0 net=5003
rlabel metal2 604 -3130 604 -3130 0 net=8912
rlabel metal2 422 -3132 422 -3132 0 net=5049
rlabel metal2 625 -3132 625 -3132 0 net=6859
rlabel metal2 863 -3132 863 -3132 0 net=9211
rlabel metal2 422 -3134 422 -3134 0 net=4633
rlabel metal2 716 -3134 716 -3134 0 net=6375
rlabel metal2 989 -3134 989 -3134 0 net=9203
rlabel metal2 492 -3136 492 -3136 0 net=6049
rlabel metal2 443 -3138 443 -3138 0 net=3891
rlabel metal2 499 -3138 499 -3138 0 net=5495
rlabel metal2 779 -3138 779 -3138 0 net=12311
rlabel metal2 499 -3140 499 -3140 0 net=5189
rlabel metal2 541 -3142 541 -3142 0 net=4669
rlabel metal2 562 -3144 562 -3144 0 net=7081
rlabel metal2 562 -3146 562 -3146 0 net=6927
rlabel metal2 569 -3148 569 -3148 0 net=6081
rlabel metal2 667 -3148 667 -3148 0 net=7931
rlabel metal2 135 -3150 135 -3150 0 net=11601
rlabel metal2 667 -3150 667 -3150 0 net=1519
rlabel metal2 58 -3161 58 -3161 0 net=2317
rlabel metal2 219 -3161 219 -3161 0 net=1759
rlabel metal2 373 -3161 373 -3161 0 net=4077
rlabel metal2 432 -3161 432 -3161 0 net=4894
rlabel metal2 569 -3161 569 -3161 0 net=6082
rlabel metal2 611 -3161 611 -3161 0 net=5230
rlabel metal2 667 -3161 667 -3161 0 net=1520
rlabel metal2 793 -3161 793 -3161 0 net=5647
rlabel metal2 845 -3161 845 -3161 0 net=9728
rlabel metal2 1080 -3161 1080 -3161 0 net=11509
rlabel metal2 1094 -3161 1094 -3161 0 net=2891
rlabel metal2 1101 -3161 1101 -3161 0 net=11399
rlabel metal2 1101 -3161 1101 -3161 0 net=11399
rlabel metal2 1188 -3161 1188 -3161 0 net=8808
rlabel metal2 1332 -3161 1332 -3161 0 net=9655
rlabel metal2 1353 -3161 1353 -3161 0 net=11621
rlabel metal2 1367 -3161 1367 -3161 0 net=12409
rlabel metal2 1367 -3161 1367 -3161 0 net=12409
rlabel metal2 1409 -3161 1409 -3161 0 net=12657
rlabel metal2 1409 -3161 1409 -3161 0 net=12657
rlabel metal2 1451 -3161 1451 -3161 0 net=12575
rlabel metal2 1451 -3161 1451 -3161 0 net=12575
rlabel metal2 1458 -3161 1458 -3161 0 net=10155
rlabel metal2 1458 -3161 1458 -3161 0 net=10155
rlabel metal2 1465 -3161 1465 -3161 0 net=8355
rlabel metal2 1465 -3161 1465 -3161 0 net=8355
rlabel metal2 65 -3163 65 -3163 0 net=11603
rlabel metal2 145 -3163 145 -3163 0 net=1291
rlabel metal2 306 -3163 306 -3163 0 net=4942
rlabel metal2 352 -3163 352 -3163 0 net=7111
rlabel metal2 415 -3163 415 -3163 0 net=3001
rlabel metal2 471 -3163 471 -3163 0 net=7382
rlabel metal2 653 -3163 653 -3163 0 net=7125
rlabel metal2 751 -3163 751 -3163 0 net=7933
rlabel metal2 856 -3163 856 -3163 0 net=12292
rlabel metal2 1080 -3163 1080 -3163 0 net=10971
rlabel metal2 1199 -3163 1199 -3163 0 net=10351
rlabel metal2 1199 -3163 1199 -3163 0 net=10351
rlabel metal2 1213 -3163 1213 -3163 0 net=10523
rlabel metal2 1213 -3163 1213 -3163 0 net=10523
rlabel metal2 1220 -3163 1220 -3163 0 net=10726
rlabel metal2 72 -3165 72 -3165 0 net=9919
rlabel metal2 296 -3165 296 -3165 0 net=3475
rlabel metal2 373 -3165 373 -3165 0 net=5191
rlabel metal2 513 -3165 513 -3165 0 net=5689
rlabel metal2 618 -3165 618 -3165 0 net=6542
rlabel metal2 716 -3165 716 -3165 0 net=6377
rlabel metal2 761 -3165 761 -3165 0 net=963
rlabel metal2 775 -3165 775 -3165 0 net=8954
rlabel metal2 856 -3165 856 -3165 0 net=10939
rlabel metal2 877 -3165 877 -3165 0 net=10909
rlabel metal2 975 -3165 975 -3165 0 net=12313
rlabel metal2 975 -3165 975 -3165 0 net=12313
rlabel metal2 985 -3165 985 -3165 0 net=11810
rlabel metal2 1227 -3165 1227 -3165 0 net=10505
rlabel metal2 1237 -3165 1237 -3165 0 net=8518
rlabel metal2 79 -3167 79 -3167 0 net=11742
rlabel metal2 250 -3167 250 -3167 0 net=7143
rlabel metal2 723 -3167 723 -3167 0 net=7231
rlabel metal2 723 -3167 723 -3167 0 net=7231
rlabel metal2 733 -3167 733 -3167 0 net=10494
rlabel metal2 919 -3167 919 -3167 0 net=2711
rlabel metal2 1094 -3167 1094 -3167 0 net=11639
rlabel metal2 79 -3169 79 -3169 0 net=9569
rlabel metal2 180 -3169 180 -3169 0 net=9891
rlabel metal2 688 -3169 688 -3169 0 net=10662
rlabel metal2 912 -3169 912 -3169 0 net=9085
rlabel metal2 964 -3169 964 -3169 0 net=9204
rlabel metal2 999 -3169 999 -3169 0 net=12608
rlabel metal2 1122 -3169 1122 -3169 0 net=8243
rlabel metal2 93 -3171 93 -3171 0 net=9106
rlabel metal2 327 -3171 327 -3171 0 net=313
rlabel metal2 387 -3171 387 -3171 0 net=2517
rlabel metal2 660 -3171 660 -3171 0 net=10002
rlabel metal2 835 -3171 835 -3171 0 net=10015
rlabel metal2 968 -3171 968 -3171 0 net=11927
rlabel metal2 1129 -3171 1129 -3171 0 net=11735
rlabel metal2 1192 -3171 1192 -3171 0 net=2437
rlabel metal2 93 -3173 93 -3173 0 net=5487
rlabel metal2 201 -3173 201 -3173 0 net=3741
rlabel metal2 401 -3173 401 -3173 0 net=4681
rlabel metal2 492 -3173 492 -3173 0 net=3893
rlabel metal2 534 -3173 534 -3173 0 net=5421
rlabel metal2 541 -3173 541 -3173 0 net=4670
rlabel metal2 870 -3173 870 -3173 0 net=9375
rlabel metal2 933 -3173 933 -3173 0 net=8733
rlabel metal2 989 -3173 989 -3173 0 net=11419
rlabel metal2 100 -3175 100 -3175 0 net=6316
rlabel metal2 156 -3175 156 -3175 0 net=2473
rlabel metal2 324 -3175 324 -3175 0 net=3999
rlabel metal2 415 -3175 415 -3175 0 net=4527
rlabel metal2 534 -3175 534 -3175 0 net=5051
rlabel metal2 569 -3175 569 -3175 0 net=9159
rlabel metal2 863 -3175 863 -3175 0 net=9213
rlabel metal2 933 -3175 933 -3175 0 net=11171
rlabel metal2 1045 -3175 1045 -3175 0 net=11761
rlabel metal2 100 -3177 100 -3177 0 net=3509
rlabel metal2 268 -3177 268 -3177 0 net=2210
rlabel metal2 422 -3177 422 -3177 0 net=4635
rlabel metal2 541 -3177 541 -3177 0 net=7083
rlabel metal2 660 -3177 660 -3177 0 net=8424
rlabel metal2 1031 -3177 1031 -3177 0 net=7593
rlabel metal2 114 -3179 114 -3179 0 net=6064
rlabel metal2 247 -3179 247 -3179 0 net=1667
rlabel metal2 422 -3179 422 -3179 0 net=3139
rlabel metal2 464 -3179 464 -3179 0 net=1523
rlabel metal2 492 -3179 492 -3179 0 net=5399
rlabel metal2 880 -3179 880 -3179 0 net=9049
rlabel metal2 940 -3179 940 -3179 0 net=9151
rlabel metal2 1006 -3179 1006 -3179 0 net=10658
rlabel metal2 1073 -3179 1073 -3179 0 net=7797
rlabel metal2 121 -3181 121 -3181 0 net=3622
rlabel metal2 436 -3181 436 -3181 0 net=10631
rlabel metal2 779 -3181 779 -3181 0 net=7577
rlabel metal2 1010 -3181 1010 -3181 0 net=9983
rlabel metal2 1115 -3181 1115 -3181 0 net=9327
rlabel metal2 121 -3183 121 -3183 0 net=7051
rlabel metal2 282 -3183 282 -3183 0 net=5077
rlabel metal2 443 -3183 443 -3183 0 net=2613
rlabel metal2 705 -3183 705 -3183 0 net=4915
rlabel metal2 1024 -3183 1024 -3183 0 net=3769
rlabel metal2 128 -3185 128 -3185 0 net=2916
rlabel metal2 128 -3185 128 -3185 0 net=2916
rlabel metal2 131 -3185 131 -3185 0 net=8129
rlabel metal2 282 -3185 282 -3185 0 net=2411
rlabel metal2 485 -3185 485 -3185 0 net=3705
rlabel metal2 548 -3185 548 -3185 0 net=5969
rlabel metal2 681 -3185 681 -3185 0 net=6587
rlabel metal2 695 -3185 695 -3185 0 net=6553
rlabel metal2 765 -3185 765 -3185 0 net=9015
rlabel metal2 884 -3185 884 -3185 0 net=7740
rlabel metal2 1115 -3185 1115 -3185 0 net=9215
rlabel metal2 135 -3187 135 -3187 0 net=2161
rlabel metal2 506 -3187 506 -3187 0 net=6295
rlabel metal2 800 -3187 800 -3187 0 net=9171
rlabel metal2 905 -3187 905 -3187 0 net=6637
rlabel metal2 1097 -3187 1097 -3187 0 net=1
rlabel metal2 1143 -3187 1143 -3187 0 net=10891
rlabel metal2 142 -3189 142 -3189 0 net=2544
rlabel metal2 331 -3189 331 -3189 0 net=2239
rlabel metal2 359 -3189 359 -3189 0 net=1501
rlabel metal2 1143 -3189 1143 -3189 0 net=2847
rlabel metal2 86 -3191 86 -3191 0 net=10326
rlabel metal2 149 -3191 149 -3191 0 net=2130
rlabel metal2 359 -3191 359 -3191 0 net=6029
rlabel metal2 408 -3191 408 -3191 0 net=3689
rlabel metal2 506 -3191 506 -3191 0 net=5497
rlabel metal2 597 -3191 597 -3191 0 net=6263
rlabel metal2 625 -3191 625 -3191 0 net=6861
rlabel metal2 786 -3191 786 -3191 0 net=7291
rlabel metal2 807 -3191 807 -3191 0 net=7193
rlabel metal2 884 -3191 884 -3191 0 net=8441
rlabel metal2 1157 -3191 1157 -3191 0 net=9510
rlabel metal2 86 -3193 86 -3193 0 net=8211
rlabel metal2 163 -3193 163 -3193 0 net=3523
rlabel metal2 380 -3193 380 -3193 0 net=7559
rlabel metal2 478 -3193 478 -3193 0 net=5669
rlabel metal2 607 -3193 607 -3193 0 net=2321
rlabel metal2 1164 -3193 1164 -3193 0 net=10806
rlabel metal2 107 -3195 107 -3195 0 net=2885
rlabel metal2 303 -3195 303 -3195 0 net=1695
rlabel metal2 632 -3195 632 -3195 0 net=6050
rlabel metal2 1171 -3195 1171 -3195 0 net=8163
rlabel metal2 163 -3197 163 -3197 0 net=2033
rlabel metal2 317 -3197 317 -3197 0 net=4195
rlabel metal2 562 -3197 562 -3197 0 net=6929
rlabel metal2 730 -3197 730 -3197 0 net=11913
rlabel metal2 814 -3197 814 -3197 0 net=8587
rlabel metal2 905 -3197 905 -3197 0 net=3725
rlabel metal2 1167 -3197 1167 -3197 0 net=7649
rlabel metal2 173 -3199 173 -3199 0 net=1573
rlabel metal2 254 -3199 254 -3199 0 net=1623
rlabel metal2 366 -3199 366 -3199 0 net=2775
rlabel metal2 527 -3199 527 -3199 0 net=6205
rlabel metal2 583 -3199 583 -3199 0 net=5303
rlabel metal2 639 -3199 639 -3199 0 net=7627
rlabel metal2 828 -3199 828 -3199 0 net=10699
rlabel metal2 926 -3199 926 -3199 0 net=10733
rlabel metal2 212 -3201 212 -3201 0 net=3117
rlabel metal2 366 -3201 366 -3201 0 net=9741
rlabel metal2 632 -3201 632 -3201 0 net=5293
rlabel metal2 646 -3201 646 -3201 0 net=1999
rlabel metal2 828 -3201 828 -3201 0 net=8537
rlabel metal2 177 -3203 177 -3203 0 net=4393
rlabel metal2 222 -3203 222 -3203 0 net=3247
rlabel metal2 310 -3203 310 -3203 0 net=4550
rlabel metal2 730 -3203 730 -3203 0 net=7461
rlabel metal2 961 -3203 961 -3203 0 net=11907
rlabel metal2 240 -3205 240 -3205 0 net=2953
rlabel metal2 450 -3205 450 -3205 0 net=5005
rlabel metal2 555 -3205 555 -3205 0 net=8933
rlabel metal2 744 -3205 744 -3205 0 net=7993
rlabel metal2 240 -3207 240 -3207 0 net=4071
rlabel metal2 289 -3207 289 -3207 0 net=3377
rlabel metal2 478 -3207 478 -3207 0 net=1895
rlabel metal2 247 -3209 247 -3209 0 net=6945
rlabel metal2 758 -3209 758 -3209 0 net=7827
rlabel metal2 261 -3211 261 -3211 0 net=4307
rlabel metal2 58 -3222 58 -3222 0 net=2318
rlabel metal2 250 -3222 250 -3222 0 net=243
rlabel metal2 250 -3222 250 -3222 0 net=243
rlabel metal2 317 -3222 317 -3222 0 net=3119
rlabel metal2 317 -3222 317 -3222 0 net=3119
rlabel metal2 338 -3222 338 -3222 0 net=3477
rlabel metal2 359 -3222 359 -3222 0 net=6030
rlabel metal2 380 -3222 380 -3222 0 net=2776
rlabel metal2 408 -3222 408 -3222 0 net=4196
rlabel metal2 702 -3222 702 -3222 0 net=6930
rlabel metal2 782 -3222 782 -3222 0 net=7594
rlabel metal2 1038 -3222 1038 -3222 0 net=9984
rlabel metal2 1066 -3222 1066 -3222 0 net=10973
rlabel metal2 1094 -3222 1094 -3222 0 net=11641
rlabel metal2 1094 -3222 1094 -3222 0 net=11641
rlabel metal2 1101 -3222 1101 -3222 0 net=11400
rlabel metal2 1129 -3222 1129 -3222 0 net=11737
rlabel metal2 1129 -3222 1129 -3222 0 net=11737
rlabel metal2 1136 -3222 1136 -3222 0 net=2892
rlabel metal2 1206 -3222 1206 -3222 0 net=7650
rlabel metal2 1290 -3222 1290 -3222 0 net=5987
rlabel metal2 1328 -3222 1328 -3222 0 net=9656
rlabel metal2 1360 -3222 1360 -3222 0 net=11623
rlabel metal2 1360 -3222 1360 -3222 0 net=11623
rlabel metal2 1367 -3222 1367 -3222 0 net=12411
rlabel metal2 1367 -3222 1367 -3222 0 net=12411
rlabel metal2 1409 -3222 1409 -3222 0 net=12659
rlabel metal2 1409 -3222 1409 -3222 0 net=12659
rlabel metal2 1451 -3222 1451 -3222 0 net=12576
rlabel metal2 1465 -3222 1465 -3222 0 net=8357
rlabel metal2 1465 -3222 1465 -3222 0 net=8357
rlabel metal2 65 -3224 65 -3224 0 net=11604
rlabel metal2 338 -3224 338 -3224 0 net=2241
rlabel metal2 359 -3224 359 -3224 0 net=2615
rlabel metal2 464 -3224 464 -3224 0 net=1524
rlabel metal2 604 -3224 604 -3224 0 net=9214
rlabel metal2 982 -3224 982 -3224 0 net=491
rlabel metal2 1234 -3224 1234 -3224 0 net=10506
rlabel metal2 1234 -3224 1234 -3224 0 net=10506
rlabel metal2 1451 -3224 1451 -3224 0 net=10157
rlabel metal2 72 -3226 72 -3226 0 net=9920
rlabel metal2 121 -3226 121 -3226 0 net=7052
rlabel metal2 380 -3226 380 -3226 0 net=4529
rlabel metal2 429 -3226 429 -3226 0 net=4078
rlabel metal2 499 -3226 499 -3226 0 net=3895
rlabel metal2 499 -3226 499 -3226 0 net=3895
rlabel metal2 520 -3226 520 -3226 0 net=3003
rlabel metal2 520 -3226 520 -3226 0 net=3003
rlabel metal2 534 -3226 534 -3226 0 net=5053
rlabel metal2 548 -3226 548 -3226 0 net=5970
rlabel metal2 737 -3226 737 -3226 0 net=6378
rlabel metal2 866 -3226 866 -3226 0 net=11172
rlabel metal2 982 -3226 982 -3226 0 net=11421
rlabel metal2 992 -3226 992 -3226 0 net=11762
rlabel metal2 1052 -3226 1052 -3226 0 net=2713
rlabel metal2 1125 -3226 1125 -3226 0 net=10769
rlabel metal2 1143 -3226 1143 -3226 0 net=2849
rlabel metal2 1143 -3226 1143 -3226 0 net=2849
rlabel metal2 1150 -3226 1150 -3226 0 net=9328
rlabel metal2 1213 -3226 1213 -3226 0 net=10525
rlabel metal2 79 -3228 79 -3228 0 net=9570
rlabel metal2 177 -3228 177 -3228 0 net=2135
rlabel metal2 201 -3228 201 -3228 0 net=2518
rlabel metal2 422 -3228 422 -3228 0 net=3141
rlabel metal2 443 -3228 443 -3228 0 net=3691
rlabel metal2 534 -3228 534 -3228 0 net=2001
rlabel metal2 730 -3228 730 -3228 0 net=7463
rlabel metal2 758 -3228 758 -3228 0 net=7829
rlabel metal2 786 -3228 786 -3228 0 net=11914
rlabel metal2 1017 -3228 1017 -3228 0 net=4916
rlabel metal2 1185 -3228 1185 -3228 0 net=10893
rlabel metal2 86 -3230 86 -3230 0 net=8212
rlabel metal2 131 -3230 131 -3230 0 net=2637
rlabel metal2 352 -3230 352 -3230 0 net=7113
rlabel metal2 450 -3230 450 -3230 0 net=3379
rlabel metal2 541 -3230 541 -3230 0 net=7085
rlabel metal2 733 -3230 733 -3230 0 net=9539
rlabel metal2 849 -3230 849 -3230 0 net=10700
rlabel metal2 996 -3230 996 -3230 0 net=1502
rlabel metal2 1150 -3230 1150 -3230 0 net=8165
rlabel metal2 1185 -3230 1185 -3230 0 net=10352
rlabel metal2 93 -3232 93 -3232 0 net=5488
rlabel metal2 187 -3232 187 -3232 0 net=9742
rlabel metal2 387 -3232 387 -3232 0 net=4001
rlabel metal2 450 -3232 450 -3232 0 net=4683
rlabel metal2 548 -3232 548 -3232 0 net=5671
rlabel metal2 604 -3232 604 -3232 0 net=2691
rlabel metal2 639 -3232 639 -3232 0 net=5295
rlabel metal2 765 -3232 765 -3232 0 net=8539
rlabel metal2 880 -3232 880 -3232 0 net=10734
rlabel metal2 933 -3232 933 -3232 0 net=11929
rlabel metal2 996 -3232 996 -3232 0 net=5285
rlabel metal2 100 -3234 100 -3234 0 net=3510
rlabel metal2 247 -3234 247 -3234 0 net=4308
rlabel metal2 282 -3234 282 -3234 0 net=2413
rlabel metal2 366 -3234 366 -3234 0 net=3425
rlabel metal2 474 -3234 474 -3234 0 net=7757
rlabel metal2 611 -3234 611 -3234 0 net=5691
rlabel metal2 807 -3234 807 -3234 0 net=7195
rlabel metal2 898 -3234 898 -3234 0 net=9051
rlabel metal2 940 -3234 940 -3234 0 net=6639
rlabel metal2 1059 -3234 1059 -3234 0 net=8244
rlabel metal2 1160 -3234 1160 -3234 0 net=3027
rlabel metal2 114 -3236 114 -3236 0 net=5400
rlabel metal2 555 -3236 555 -3236 0 net=9172
rlabel metal2 898 -3236 898 -3236 0 net=9087
rlabel metal2 919 -3236 919 -3236 0 net=9665
rlabel metal2 1164 -3236 1164 -3236 0 net=2439
rlabel metal2 135 -3238 135 -3238 0 net=2163
rlabel metal2 191 -3238 191 -3238 0 net=3661
rlabel metal2 555 -3238 555 -3238 0 net=6207
rlabel metal2 569 -3238 569 -3238 0 net=9160
rlabel metal2 611 -3238 611 -3238 0 net=7127
rlabel metal2 800 -3238 800 -3238 0 net=7293
rlabel metal2 856 -3238 856 -3238 0 net=10941
rlabel metal2 940 -3238 940 -3238 0 net=9153
rlabel metal2 1073 -3238 1073 -3238 0 net=7799
rlabel metal2 1073 -3238 1073 -3238 0 net=7799
rlabel metal2 1080 -3238 1080 -3238 0 net=9217
rlabel metal2 149 -3240 149 -3240 0 net=5201
rlabel metal2 527 -3240 527 -3240 0 net=5007
rlabel metal2 618 -3240 618 -3240 0 net=6265
rlabel metal2 628 -3240 628 -3240 0 net=7994
rlabel metal2 793 -3240 793 -3240 0 net=7935
rlabel metal2 884 -3240 884 -3240 0 net=8443
rlabel metal2 947 -3240 947 -3240 0 net=8735
rlabel metal2 1087 -3240 1087 -3240 0 net=11511
rlabel metal2 152 -3242 152 -3242 0 net=9573
rlabel metal2 618 -3242 618 -3242 0 net=5209
rlabel metal2 653 -3242 653 -3242 0 net=6589
rlabel metal2 744 -3242 744 -3242 0 net=7629
rlabel metal2 793 -3242 793 -3242 0 net=9017
rlabel metal2 842 -3242 842 -3242 0 net=5649
rlabel metal2 226 -3244 226 -3244 0 net=1575
rlabel metal2 264 -3244 264 -3244 0 net=9457
rlabel metal2 296 -3244 296 -3244 0 net=3743
rlabel metal2 513 -3244 513 -3244 0 net=4637
rlabel metal2 558 -3244 558 -3244 0 net=5422
rlabel metal2 751 -3244 751 -3244 0 net=7579
rlabel metal2 821 -3244 821 -3244 0 net=11909
rlabel metal2 107 -3246 107 -3246 0 net=2886
rlabel metal2 268 -3246 268 -3246 0 net=1669
rlabel metal2 296 -3246 296 -3246 0 net=1697
rlabel metal2 394 -3246 394 -3246 0 net=7560
rlabel metal2 635 -3246 635 -3246 0 net=10632
rlabel metal2 842 -3246 842 -3246 0 net=9377
rlabel metal2 884 -3246 884 -3246 0 net=3727
rlabel metal2 961 -3246 961 -3246 0 net=3771
rlabel metal2 156 -3248 156 -3248 0 net=2474
rlabel metal2 506 -3248 506 -3248 0 net=5499
rlabel metal2 562 -3248 562 -3248 0 net=5305
rlabel metal2 660 -3248 660 -3248 0 net=7645
rlabel metal2 772 -3248 772 -3248 0 net=8589
rlabel metal2 870 -3248 870 -3248 0 net=10911
rlabel metal2 905 -3248 905 -3248 0 net=12315
rlabel metal2 156 -3250 156 -3250 0 net=9385
rlabel metal2 268 -3250 268 -3250 0 net=6947
rlabel metal2 436 -3250 436 -3250 0 net=5079
rlabel metal2 660 -3250 660 -3250 0 net=6863
rlabel metal2 877 -3250 877 -3250 0 net=2322
rlabel metal2 198 -3252 198 -3252 0 net=1911
rlabel metal2 373 -3252 373 -3252 0 net=5193
rlabel metal2 506 -3252 506 -3252 0 net=3189
rlabel metal2 667 -3252 667 -3252 0 net=9893
rlabel metal2 184 -3254 184 -3254 0 net=8131
rlabel metal2 219 -3254 219 -3254 0 net=1761
rlabel metal2 331 -3254 331 -3254 0 net=3525
rlabel metal2 590 -3254 590 -3254 0 net=8935
rlabel metal2 212 -3256 212 -3256 0 net=4395
rlabel metal2 226 -3256 226 -3256 0 net=1625
rlabel metal2 310 -3256 310 -3256 0 net=2955
rlabel metal2 667 -3256 667 -3256 0 net=7145
rlabel metal2 212 -3258 212 -3258 0 net=3249
rlabel metal2 310 -3258 310 -3258 0 net=1897
rlabel metal2 674 -3258 674 -3258 0 net=6297
rlabel metal2 709 -3258 709 -3258 0 net=6555
rlabel metal2 1454 -3258 1454 -3258 0 net=1
rlabel metal2 163 -3260 163 -3260 0 net=2035
rlabel metal2 478 -3260 478 -3260 0 net=3707
rlabel metal2 681 -3260 681 -3260 0 net=7233
rlabel metal2 163 -3262 163 -3262 0 net=5235
rlabel metal2 408 -3262 408 -3262 0 net=5097
rlabel metal2 709 -3262 709 -3262 0 net=10017
rlabel metal2 208 -3264 208 -3264 0 net=4072
rlabel metal2 240 -3266 240 -3266 0 net=1687
rlabel metal2 163 -3277 163 -3277 0 net=5236
rlabel metal2 243 -3277 243 -3277 0 net=2002
rlabel metal2 593 -3277 593 -3277 0 net=7086
rlabel metal2 670 -3277 670 -3277 0 net=6298
rlabel metal2 684 -3277 684 -3277 0 net=5296
rlabel metal2 723 -3277 723 -3277 0 net=9666
rlabel metal2 936 -3277 936 -3277 0 net=9154
rlabel metal2 947 -3277 947 -3277 0 net=5651
rlabel metal2 982 -3277 982 -3277 0 net=11423
rlabel metal2 1003 -3277 1003 -3277 0 net=6640
rlabel metal2 1066 -3277 1066 -3277 0 net=10975
rlabel metal2 1066 -3277 1066 -3277 0 net=10975
rlabel metal2 1073 -3277 1073 -3277 0 net=7801
rlabel metal2 1094 -3277 1094 -3277 0 net=11642
rlabel metal2 1094 -3277 1094 -3277 0 net=11642
rlabel metal2 1108 -3277 1108 -3277 0 net=11513
rlabel metal2 1122 -3277 1122 -3277 0 net=11738
rlabel metal2 1136 -3277 1136 -3277 0 net=10770
rlabel metal2 1171 -3277 1171 -3277 0 net=3028
rlabel metal2 1206 -3277 1206 -3277 0 net=10895
rlabel metal2 1216 -3277 1216 -3277 0 net=10526
rlabel metal2 1251 -3277 1251 -3277 0 net=5988
rlabel metal2 1360 -3277 1360 -3277 0 net=11625
rlabel metal2 1360 -3277 1360 -3277 0 net=11625
rlabel metal2 1367 -3277 1367 -3277 0 net=12413
rlabel metal2 1367 -3277 1367 -3277 0 net=12413
rlabel metal2 1409 -3277 1409 -3277 0 net=12661
rlabel metal2 1409 -3277 1409 -3277 0 net=12661
rlabel metal2 1451 -3277 1451 -3277 0 net=10158
rlabel metal2 177 -3279 177 -3279 0 net=2137
rlabel metal2 208 -3279 208 -3279 0 net=2441
rlabel metal2 289 -3279 289 -3279 0 net=1912
rlabel metal2 415 -3279 415 -3279 0 net=7115
rlabel metal2 688 -3279 688 -3279 0 net=7647
rlabel metal2 730 -3279 730 -3279 0 net=7580
rlabel metal2 779 -3279 779 -3279 0 net=7936
rlabel metal2 807 -3279 807 -3279 0 net=7294
rlabel metal2 838 -3279 838 -3279 0 net=5286
rlabel metal2 1073 -3279 1073 -3279 0 net=9219
rlabel metal2 1097 -3279 1097 -3279 0 net=8491
rlabel metal2 1458 -3279 1458 -3279 0 net=8358
rlabel metal2 177 -3281 177 -3281 0 net=6949
rlabel metal2 282 -3281 282 -3281 0 net=1671
rlabel metal2 331 -3281 331 -3281 0 net=2956
rlabel metal2 394 -3281 394 -3281 0 net=5210
rlabel metal2 639 -3281 639 -3281 0 net=5693
rlabel metal2 681 -3281 681 -3281 0 net=7235
rlabel metal2 751 -3281 751 -3281 0 net=7831
rlabel metal2 779 -3281 779 -3281 0 net=9541
rlabel metal2 793 -3281 793 -3281 0 net=9019
rlabel metal2 814 -3281 814 -3281 0 net=9895
rlabel metal2 856 -3281 856 -3281 0 net=3383
rlabel metal2 912 -3281 912 -3281 0 net=8445
rlabel metal2 940 -3281 940 -3281 0 net=8737
rlabel metal2 1101 -3281 1101 -3281 0 net=2715
rlabel metal2 1125 -3281 1125 -3281 0 net=2440
rlabel metal2 184 -3283 184 -3283 0 net=3662
rlabel metal2 212 -3283 212 -3283 0 net=3251
rlabel metal2 212 -3283 212 -3283 0 net=3251
rlabel metal2 226 -3283 226 -3283 0 net=1627
rlabel metal2 282 -3283 282 -3283 0 net=1699
rlabel metal2 324 -3283 324 -3283 0 net=2639
rlabel metal2 415 -3283 415 -3283 0 net=3143
rlabel metal2 457 -3283 457 -3283 0 net=3380
rlabel metal2 593 -3283 593 -3283 0 net=10018
rlabel metal2 712 -3283 712 -3283 0 net=9953
rlabel metal2 828 -3283 828 -3283 0 net=7197
rlabel metal2 828 -3283 828 -3283 0 net=7197
rlabel metal2 863 -3283 863 -3283 0 net=3729
rlabel metal2 912 -3283 912 -3283 0 net=11931
rlabel metal2 954 -3283 954 -3283 0 net=3773
rlabel metal2 1136 -3283 1136 -3283 0 net=8166
rlabel metal2 156 -3285 156 -3285 0 net=9387
rlabel metal2 226 -3285 226 -3285 0 net=186
rlabel metal2 639 -3285 639 -3285 0 net=6865
rlabel metal2 681 -3285 681 -3285 0 net=9591
rlabel metal2 870 -3285 870 -3285 0 net=10913
rlabel metal2 926 -3285 926 -3285 0 net=9053
rlabel metal2 1143 -3285 1143 -3285 0 net=2851
rlabel metal2 1143 -3285 1143 -3285 0 net=2851
rlabel metal2 184 -3287 184 -3287 0 net=8133
rlabel metal2 296 -3287 296 -3287 0 net=7581
rlabel metal2 576 -3287 576 -3287 0 net=9574
rlabel metal2 187 -3289 187 -3289 0 net=1563
rlabel metal2 331 -3289 331 -3289 0 net=3479
rlabel metal2 359 -3289 359 -3289 0 net=2617
rlabel metal2 359 -3289 359 -3289 0 net=2617
rlabel metal2 366 -3289 366 -3289 0 net=3426
rlabel metal2 597 -3289 597 -3289 0 net=7759
rlabel metal2 744 -3289 744 -3289 0 net=7631
rlabel metal2 793 -3289 793 -3289 0 net=11911
rlabel metal2 877 -3289 877 -3289 0 net=9089
rlabel metal2 198 -3291 198 -3291 0 net=4397
rlabel metal2 338 -3291 338 -3291 0 net=2243
rlabel metal2 366 -3291 366 -3291 0 net=4003
rlabel metal2 422 -3291 422 -3291 0 net=3745
rlabel metal2 471 -3291 471 -3291 0 net=3709
rlabel metal2 488 -3291 488 -3291 0 net=5080
rlabel metal2 611 -3291 611 -3291 0 net=7129
rlabel metal2 611 -3291 611 -3291 0 net=7129
rlabel metal2 635 -3291 635 -3291 0 net=5133
rlabel metal2 891 -3291 891 -3291 0 net=10943
rlabel metal2 170 -3293 170 -3293 0 net=2165
rlabel metal2 373 -3293 373 -3293 0 net=3527
rlabel metal2 446 -3293 446 -3293 0 net=11035
rlabel metal2 758 -3293 758 -3293 0 net=8541
rlabel metal2 821 -3293 821 -3293 0 net=9379
rlabel metal2 898 -3293 898 -3293 0 net=12317
rlabel metal2 219 -3295 219 -3295 0 net=2037
rlabel metal2 275 -3295 275 -3295 0 net=9459
rlabel metal2 422 -3295 422 -3295 0 net=3191
rlabel metal2 534 -3295 534 -3295 0 net=5055
rlabel metal2 555 -3295 555 -3295 0 net=6209
rlabel metal2 660 -3295 660 -3295 0 net=6557
rlabel metal2 765 -3295 765 -3295 0 net=8591
rlabel metal2 842 -3295 842 -3295 0 net=1068
rlabel metal2 880 -3295 880 -3295 0 net=7035
rlabel metal2 233 -3297 233 -3297 0 net=5099
rlabel metal2 464 -3297 464 -3297 0 net=5203
rlabel metal2 576 -3297 576 -3297 0 net=3937
rlabel metal2 716 -3297 716 -3297 0 net=7465
rlabel metal2 254 -3299 254 -3299 0 net=1577
rlabel metal2 317 -3299 317 -3299 0 net=3121
rlabel metal2 464 -3299 464 -3299 0 net=2692
rlabel metal2 695 -3299 695 -3299 0 net=8937
rlabel metal2 254 -3301 254 -3301 0 net=2415
rlabel metal2 401 -3301 401 -3301 0 net=7695
rlabel metal2 737 -3301 737 -3301 0 net=6299
rlabel metal2 310 -3303 310 -3303 0 net=1899
rlabel metal2 352 -3303 352 -3303 0 net=2427
rlabel metal2 492 -3303 492 -3303 0 net=1688
rlabel metal2 583 -3303 583 -3303 0 net=5569
rlabel metal2 303 -3305 303 -3305 0 net=1763
rlabel metal2 380 -3305 380 -3305 0 net=4531
rlabel metal2 604 -3305 604 -3305 0 net=6563
rlabel metal2 303 -3307 303 -3307 0 net=1709
rlabel metal2 380 -3309 380 -3309 0 net=7959
rlabel metal2 401 -3311 401 -3311 0 net=4685
rlabel metal2 467 -3311 467 -3311 0 net=9461
rlabel metal2 436 -3313 436 -3313 0 net=5195
rlabel metal2 436 -3315 436 -3315 0 net=3693
rlabel metal2 450 -3315 450 -3315 0 net=6267
rlabel metal2 324 -3317 324 -3317 0 net=3023
rlabel metal2 474 -3317 474 -3317 0 net=5500
rlabel metal2 625 -3317 625 -3317 0 net=6591
rlabel metal2 478 -3319 478 -3319 0 net=3897
rlabel metal2 513 -3319 513 -3319 0 net=7147
rlabel metal2 499 -3321 499 -3321 0 net=3005
rlabel metal2 548 -3321 548 -3321 0 net=5673
rlabel metal2 506 -3323 506 -3323 0 net=11325
rlabel metal2 520 -3325 520 -3325 0 net=4639
rlabel metal2 548 -3325 548 -3325 0 net=5307
rlabel metal2 408 -3327 408 -3327 0 net=11679
rlabel metal2 527 -3329 527 -3329 0 net=5009
rlabel metal2 184 -3340 184 -3340 0 net=8135
rlabel metal2 184 -3340 184 -3340 0 net=8135
rlabel metal2 191 -3340 191 -3340 0 net=9389
rlabel metal2 261 -3340 261 -3340 0 net=1197
rlabel metal2 621 -3340 621 -3340 0 net=7632
rlabel metal2 807 -3340 807 -3340 0 net=9592
rlabel metal2 870 -3340 870 -3340 0 net=5134
rlabel metal2 1115 -3340 1115 -3340 0 net=11515
rlabel metal2 1139 -3340 1139 -3340 0 net=2852
rlabel metal2 1213 -3340 1213 -3340 0 net=10897
rlabel metal2 1213 -3340 1213 -3340 0 net=10897
rlabel metal2 1353 -3340 1353 -3340 0 net=12415
rlabel metal2 1409 -3340 1409 -3340 0 net=12663
rlabel metal2 1409 -3340 1409 -3340 0 net=12663
rlabel metal2 191 -3342 191 -3342 0 net=5101
rlabel metal2 240 -3342 240 -3342 0 net=2443
rlabel metal2 264 -3342 264 -3342 0 net=1578
rlabel metal2 282 -3342 282 -3342 0 net=1700
rlabel metal2 429 -3342 429 -3342 0 net=3529
rlabel metal2 429 -3342 429 -3342 0 net=3529
rlabel metal2 471 -3342 471 -3342 0 net=3710
rlabel metal2 576 -3342 576 -3342 0 net=3939
rlabel metal2 604 -3342 604 -3342 0 net=6565
rlabel metal2 695 -3342 695 -3342 0 net=7697
rlabel metal2 695 -3342 695 -3342 0 net=7697
rlabel metal2 702 -3342 702 -3342 0 net=7648
rlabel metal2 702 -3342 702 -3342 0 net=7648
rlabel metal2 709 -3342 709 -3342 0 net=1170
rlabel metal2 779 -3342 779 -3342 0 net=9543
rlabel metal2 779 -3342 779 -3342 0 net=9543
rlabel metal2 821 -3342 821 -3342 0 net=9381
rlabel metal2 842 -3342 842 -3342 0 net=10914
rlabel metal2 894 -3342 894 -3342 0 net=10944
rlabel metal2 940 -3342 940 -3342 0 net=8739
rlabel metal2 940 -3342 940 -3342 0 net=8739
rlabel metal2 947 -3342 947 -3342 0 net=9054
rlabel metal2 975 -3342 975 -3342 0 net=5653
rlabel metal2 1059 -3342 1059 -3342 0 net=9220
rlabel metal2 1108 -3342 1108 -3342 0 net=2717
rlabel metal2 1290 -3342 1290 -3342 0 net=8493
rlabel metal2 198 -3344 198 -3344 0 net=4399
rlabel metal2 254 -3344 254 -3344 0 net=2417
rlabel metal2 282 -3344 282 -3344 0 net=1673
rlabel metal2 303 -3344 303 -3344 0 net=1711
rlabel metal2 338 -3344 338 -3344 0 net=2166
rlabel metal2 471 -3344 471 -3344 0 net=4641
rlabel metal2 541 -3344 541 -3344 0 net=667
rlabel metal2 989 -3344 989 -3344 0 net=11425
rlabel metal2 989 -3344 989 -3344 0 net=11425
rlabel metal2 1062 -3344 1062 -3344 0 net=10976
rlabel metal2 1073 -3344 1073 -3344 0 net=7803
rlabel metal2 1360 -3344 1360 -3344 0 net=11627
rlabel metal2 1360 -3344 1360 -3344 0 net=11627
rlabel metal2 198 -3346 198 -3346 0 net=2429
rlabel metal2 355 -3346 355 -3346 0 net=11326
rlabel metal2 513 -3346 513 -3346 0 net=7149
rlabel metal2 513 -3346 513 -3346 0 net=7149
rlabel metal2 520 -3346 520 -3346 0 net=5011
rlabel metal2 558 -3346 558 -3346 0 net=12689
rlabel metal2 604 -3346 604 -3346 0 net=7117
rlabel metal2 660 -3346 660 -3346 0 net=6559
rlabel metal2 712 -3346 712 -3346 0 net=11912
rlabel metal2 828 -3346 828 -3346 0 net=7198
rlabel metal2 849 -3346 849 -3346 0 net=9897
rlabel metal2 849 -3346 849 -3346 0 net=9897
rlabel metal2 856 -3346 856 -3346 0 net=3385
rlabel metal2 856 -3346 856 -3346 0 net=3385
rlabel metal2 870 -3346 870 -3346 0 net=7037
rlabel metal2 919 -3346 919 -3346 0 net=8447
rlabel metal2 919 -3346 919 -3346 0 net=8447
rlabel metal2 926 -3346 926 -3346 0 net=3775
rlabel metal2 226 -3348 226 -3348 0 net=9269
rlabel metal2 737 -3348 737 -3348 0 net=9020
rlabel metal2 884 -3348 884 -3348 0 net=6301
rlabel metal2 905 -3348 905 -3348 0 net=11933
rlabel metal2 247 -3350 247 -3350 0 net=1629
rlabel metal2 268 -3350 268 -3350 0 net=1564
rlabel metal2 492 -3350 492 -3350 0 net=5196
rlabel metal2 555 -3350 555 -3350 0 net=5205
rlabel metal2 737 -3350 737 -3350 0 net=8543
rlabel metal2 775 -3350 775 -3350 0 net=11817
rlabel metal2 877 -3350 877 -3350 0 net=9091
rlabel metal2 212 -3352 212 -3352 0 net=3253
rlabel metal2 289 -3352 289 -3352 0 net=1901
rlabel metal2 366 -3352 366 -3352 0 net=4004
rlabel metal2 383 -3352 383 -3352 0 net=9460
rlabel metal2 394 -3352 394 -3352 0 net=2640
rlabel metal2 495 -3352 495 -3352 0 net=12017
rlabel metal2 744 -3352 744 -3352 0 net=11036
rlabel metal2 863 -3352 863 -3352 0 net=3731
rlabel metal2 177 -3354 177 -3354 0 net=6950
rlabel metal2 397 -3354 397 -3354 0 net=357
rlabel metal2 744 -3354 744 -3354 0 net=8939
rlabel metal2 863 -3354 863 -3354 0 net=12318
rlabel metal2 177 -3356 177 -3356 0 net=11609
rlabel metal2 296 -3356 296 -3356 0 net=7583
rlabel metal2 373 -3356 373 -3356 0 net=3123
rlabel metal2 443 -3356 443 -3356 0 net=9439
rlabel metal2 576 -3356 576 -3356 0 net=10529
rlabel metal2 758 -3356 758 -3356 0 net=8593
rlabel metal2 205 -3358 205 -3358 0 net=2139
rlabel metal2 219 -3358 219 -3358 0 net=2039
rlabel metal2 296 -3358 296 -3358 0 net=2619
rlabel metal2 373 -3358 373 -3358 0 net=3747
rlabel metal2 499 -3358 499 -3358 0 net=3006
rlabel metal2 751 -3358 751 -3358 0 net=7833
rlabel metal2 205 -3360 205 -3360 0 net=3025
rlabel metal2 359 -3360 359 -3360 0 net=1821
rlabel metal2 499 -3360 499 -3360 0 net=11681
rlabel metal2 730 -3360 730 -3360 0 net=7961
rlabel metal2 219 -3362 219 -3362 0 net=3481
rlabel metal2 415 -3362 415 -3362 0 net=3145
rlabel metal2 716 -3362 716 -3362 0 net=7467
rlabel metal2 303 -3364 303 -3364 0 net=1765
rlabel metal2 317 -3364 317 -3364 0 net=12243
rlabel metal2 450 -3364 450 -3364 0 net=6269
rlabel metal2 639 -3364 639 -3364 0 net=6867
rlabel metal2 310 -3366 310 -3366 0 net=3193
rlabel metal2 450 -3366 450 -3366 0 net=3899
rlabel metal2 639 -3366 639 -3366 0 net=5695
rlabel metal2 306 -3368 306 -3368 0 net=1
rlabel metal2 478 -3368 478 -3368 0 net=5057
rlabel metal2 667 -3368 667 -3368 0 net=9395
rlabel metal2 324 -3370 324 -3370 0 net=2245
rlabel metal2 352 -3370 352 -3370 0 net=9579
rlabel metal2 625 -3370 625 -3370 0 net=6593
rlabel metal2 331 -3372 331 -3372 0 net=3695
rlabel metal2 611 -3372 611 -3372 0 net=7131
rlabel metal2 345 -3374 345 -3374 0 net=2785
rlabel metal2 611 -3374 611 -3374 0 net=7761
rlabel metal2 401 -3376 401 -3376 0 net=4687
rlabel metal2 723 -3376 723 -3376 0 net=12293
rlabel metal2 401 -3378 401 -3378 0 net=3873
rlabel metal2 814 -3378 814 -3378 0 net=9954
rlabel metal2 408 -3380 408 -3380 0 net=4533
rlabel metal2 814 -3380 814 -3380 0 net=1865
rlabel metal2 485 -3382 485 -3382 0 net=5674
rlabel metal2 653 -3384 653 -3384 0 net=7237
rlabel metal2 583 -3386 583 -3386 0 net=5571
rlabel metal2 583 -3388 583 -3388 0 net=9463
rlabel metal2 548 -3390 548 -3390 0 net=5309
rlabel metal2 548 -3392 548 -3392 0 net=6211
rlabel metal2 446 -3394 446 -3394 0 net=11293
rlabel metal2 177 -3405 177 -3405 0 net=11610
rlabel metal2 247 -3405 247 -3405 0 net=2040
rlabel metal2 366 -3405 366 -3405 0 net=7584
rlabel metal2 443 -3405 443 -3405 0 net=9441
rlabel metal2 443 -3405 443 -3405 0 net=9441
rlabel metal2 457 -3405 457 -3405 0 net=3146
rlabel metal2 499 -3405 499 -3405 0 net=11682
rlabel metal2 513 -3405 513 -3405 0 net=7150
rlabel metal2 632 -3405 632 -3405 0 net=5311
rlabel metal2 674 -3405 674 -3405 0 net=9397
rlabel metal2 674 -3405 674 -3405 0 net=9397
rlabel metal2 695 -3405 695 -3405 0 net=7699
rlabel metal2 709 -3405 709 -3405 0 net=6561
rlabel metal2 709 -3405 709 -3405 0 net=6561
rlabel metal2 719 -3405 719 -3405 0 net=8544
rlabel metal2 744 -3405 744 -3405 0 net=8941
rlabel metal2 744 -3405 744 -3405 0 net=8941
rlabel metal2 751 -3405 751 -3405 0 net=7963
rlabel metal2 751 -3405 751 -3405 0 net=7963
rlabel metal2 765 -3405 765 -3405 0 net=7834
rlabel metal2 782 -3405 782 -3405 0 net=4779
rlabel metal2 989 -3405 989 -3405 0 net=11427
rlabel metal2 989 -3405 989 -3405 0 net=11427
rlabel metal2 996 -3405 996 -3405 0 net=5655
rlabel metal2 996 -3405 996 -3405 0 net=5655
rlabel metal2 1073 -3405 1073 -3405 0 net=7805
rlabel metal2 1073 -3405 1073 -3405 0 net=7805
rlabel metal2 1115 -3405 1115 -3405 0 net=2719
rlabel metal2 1115 -3405 1115 -3405 0 net=2719
rlabel metal2 1122 -3405 1122 -3405 0 net=11517
rlabel metal2 1122 -3405 1122 -3405 0 net=11517
rlabel metal2 1213 -3405 1213 -3405 0 net=10899
rlabel metal2 1213 -3405 1213 -3405 0 net=10899
rlabel metal2 1353 -3405 1353 -3405 0 net=12417
rlabel metal2 1353 -3405 1353 -3405 0 net=12417
rlabel metal2 1360 -3405 1360 -3405 0 net=11629
rlabel metal2 1360 -3405 1360 -3405 0 net=11629
rlabel metal2 1367 -3405 1367 -3405 0 net=8495
rlabel metal2 1409 -3405 1409 -3405 0 net=12665
rlabel metal2 1409 -3405 1409 -3405 0 net=12665
rlabel metal2 184 -3407 184 -3407 0 net=8136
rlabel metal2 264 -3407 264 -3407 0 net=3254
rlabel metal2 275 -3407 275 -3407 0 net=2418
rlabel metal2 467 -3407 467 -3407 0 net=7118
rlabel metal2 632 -3407 632 -3407 0 net=7239
rlabel metal2 681 -3407 681 -3407 0 net=10531
rlabel metal2 772 -3407 772 -3407 0 net=9544
rlabel metal2 831 -3407 831 -3407 0 net=3386
rlabel metal2 891 -3407 891 -3407 0 net=3776
rlabel metal2 940 -3407 940 -3407 0 net=8741
rlabel metal2 940 -3407 940 -3407 0 net=8741
rlabel metal2 947 -3407 947 -3407 0 net=8545
rlabel metal2 968 -3407 968 -3407 0 net=7477
rlabel metal2 212 -3409 212 -3409 0 net=2140
rlabel metal2 233 -3409 233 -3409 0 net=9391
rlabel metal2 282 -3409 282 -3409 0 net=1675
rlabel metal2 282 -3409 282 -3409 0 net=1675
rlabel metal2 310 -3409 310 -3409 0 net=3195
rlabel metal2 471 -3409 471 -3409 0 net=4643
rlabel metal2 499 -3409 499 -3409 0 net=8747
rlabel metal2 558 -3409 558 -3409 0 net=7132
rlabel metal2 653 -3409 653 -3409 0 net=6595
rlabel metal2 688 -3409 688 -3409 0 net=5572
rlabel metal2 842 -3409 842 -3409 0 net=7038
rlabel metal2 912 -3409 912 -3409 0 net=9093
rlabel metal2 954 -3409 954 -3409 0 net=9607
rlabel metal2 254 -3411 254 -3411 0 net=1631
rlabel metal2 317 -3411 317 -3411 0 net=12244
rlabel metal2 341 -3411 341 -3411 0 net=3124
rlabel metal2 408 -3411 408 -3411 0 net=4535
rlabel metal2 478 -3411 478 -3411 0 net=5059
rlabel metal2 520 -3411 520 -3411 0 net=5012
rlabel metal2 569 -3411 569 -3411 0 net=12691
rlabel metal2 625 -3411 625 -3411 0 net=5697
rlabel metal2 660 -3411 660 -3411 0 net=5207
rlabel metal2 688 -3411 688 -3411 0 net=12295
rlabel metal2 730 -3411 730 -3411 0 net=7469
rlabel metal2 842 -3411 842 -3411 0 net=11657
rlabel metal2 849 -3411 849 -3411 0 net=9899
rlabel metal2 849 -3411 849 -3411 0 net=9899
rlabel metal2 856 -3411 856 -3411 0 net=6303
rlabel metal2 905 -3411 905 -3411 0 net=11935
rlabel metal2 919 -3411 919 -3411 0 net=8449
rlabel metal2 919 -3411 919 -3411 0 net=8449
rlabel metal2 961 -3411 961 -3411 0 net=3789
rlabel metal2 191 -3413 191 -3413 0 net=5102
rlabel metal2 352 -3413 352 -3413 0 net=3875
rlabel metal2 534 -3413 534 -3413 0 net=6212
rlabel metal2 569 -3413 569 -3413 0 net=3940
rlabel metal2 597 -3413 597 -3413 0 net=11295
rlabel metal2 695 -3413 695 -3413 0 net=6869
rlabel metal2 723 -3413 723 -3413 0 net=1866
rlabel metal2 863 -3413 863 -3413 0 net=8693
rlabel metal2 877 -3413 877 -3413 0 net=3733
rlabel metal2 240 -3415 240 -3415 0 net=4401
rlabel metal2 261 -3415 261 -3415 0 net=2445
rlabel metal2 289 -3415 289 -3415 0 net=1903
rlabel metal2 327 -3415 327 -3415 0 net=9580
rlabel metal2 488 -3415 488 -3415 0 net=9857
rlabel metal2 541 -3415 541 -3415 0 net=3259
rlabel metal2 730 -3415 730 -3415 0 net=8595
rlabel metal2 821 -3415 821 -3415 0 net=11819
rlabel metal2 198 -3417 198 -3417 0 net=2431
rlabel metal2 331 -3417 331 -3417 0 net=3697
rlabel metal2 527 -3417 527 -3417 0 net=12019
rlabel metal2 562 -3417 562 -3417 0 net=6271
rlabel metal2 639 -3417 639 -3417 0 net=950
rlabel metal2 821 -3417 821 -3417 0 net=9383
rlabel metal2 359 -3419 359 -3419 0 net=1823
rlabel metal2 562 -3419 562 -3419 0 net=9465
rlabel metal2 646 -3419 646 -3419 0 net=9271
rlabel metal2 296 -3421 296 -3421 0 net=2621
rlabel metal2 373 -3421 373 -3421 0 net=3749
rlabel metal2 583 -3421 583 -3421 0 net=7763
rlabel metal2 618 -3421 618 -3421 0 net=6567
rlabel metal2 733 -3421 733 -3421 0 net=1
rlabel metal2 219 -3423 219 -3423 0 net=3483
rlabel metal2 303 -3423 303 -3423 0 net=1767
rlabel metal2 303 -3425 303 -3425 0 net=3530
rlabel metal2 429 -3427 429 -3427 0 net=4689
rlabel metal2 436 -3429 436 -3429 0 net=3901
rlabel metal2 422 -3431 422 -3431 0 net=1713
rlabel metal2 345 -3433 345 -3433 0 net=2787
rlabel metal2 324 -3435 324 -3435 0 net=2247
rlabel metal2 205 -3437 205 -3437 0 net=3026
rlabel metal2 222 -3448 222 -3448 0 net=536
rlabel metal2 338 -3448 338 -3448 0 net=3877
rlabel metal2 359 -3448 359 -3448 0 net=2623
rlabel metal2 401 -3448 401 -3448 0 net=3698
rlabel metal2 478 -3448 478 -3448 0 net=4645
rlabel metal2 492 -3448 492 -3448 0 net=5061
rlabel metal2 492 -3448 492 -3448 0 net=5061
rlabel metal2 506 -3448 506 -3448 0 net=3261
rlabel metal2 548 -3448 548 -3448 0 net=12021
rlabel metal2 548 -3448 548 -3448 0 net=12021
rlabel metal2 597 -3448 597 -3448 0 net=6273
rlabel metal2 614 -3448 614 -3448 0 net=5698
rlabel metal2 642 -3448 642 -3448 0 net=12296
rlabel metal2 698 -3448 698 -3448 0 net=7700
rlabel metal2 709 -3448 709 -3448 0 net=6562
rlabel metal2 740 -3448 740 -3448 0 net=7470
rlabel metal2 765 -3448 765 -3448 0 net=10532
rlabel metal2 782 -3448 782 -3448 0 net=394
rlabel metal2 982 -3448 982 -3448 0 net=4781
rlabel metal2 1073 -3448 1073 -3448 0 net=7806
rlabel metal2 1094 -3448 1094 -3448 0 net=3790
rlabel metal2 1223 -3448 1223 -3448 0 net=4507
rlabel metal2 1353 -3448 1353 -3448 0 net=12419
rlabel metal2 1353 -3448 1353 -3448 0 net=12419
rlabel metal2 1360 -3448 1360 -3448 0 net=11631
rlabel metal2 1360 -3448 1360 -3448 0 net=11631
rlabel metal2 1409 -3448 1409 -3448 0 net=12667
rlabel metal2 254 -3450 254 -3450 0 net=4403
rlabel metal2 264 -3450 264 -3450 0 net=1091
rlabel metal2 471 -3450 471 -3450 0 net=4537
rlabel metal2 520 -3450 520 -3450 0 net=2689
rlabel metal2 621 -3450 621 -3450 0 net=1438
rlabel metal2 737 -3450 737 -3450 0 net=7965
rlabel metal2 821 -3450 821 -3450 0 net=9384
rlabel metal2 831 -3450 831 -3450 0 net=9900
rlabel metal2 856 -3450 856 -3450 0 net=6305
rlabel metal2 856 -3450 856 -3450 0 net=6305
rlabel metal2 884 -3450 884 -3450 0 net=3735
rlabel metal2 884 -3450 884 -3450 0 net=3735
rlabel metal2 912 -3450 912 -3450 0 net=11937
rlabel metal2 912 -3450 912 -3450 0 net=11937
rlabel metal2 919 -3450 919 -3450 0 net=8451
rlabel metal2 919 -3450 919 -3450 0 net=8451
rlabel metal2 926 -3450 926 -3450 0 net=9095
rlabel metal2 926 -3450 926 -3450 0 net=9095
rlabel metal2 933 -3450 933 -3450 0 net=10551
rlabel metal2 957 -3450 957 -3450 0 net=7478
rlabel metal2 989 -3450 989 -3450 0 net=11429
rlabel metal2 989 -3450 989 -3450 0 net=11429
rlabel metal2 996 -3450 996 -3450 0 net=5657
rlabel metal2 996 -3450 996 -3450 0 net=5657
rlabel metal2 1010 -3450 1010 -3450 0 net=9608
rlabel metal2 1115 -3450 1115 -3450 0 net=2721
rlabel metal2 1115 -3450 1115 -3450 0 net=2721
rlabel metal2 1122 -3450 1122 -3450 0 net=11519
rlabel metal2 1122 -3450 1122 -3450 0 net=11519
rlabel metal2 1213 -3450 1213 -3450 0 net=10901
rlabel metal2 1213 -3450 1213 -3450 0 net=10901
rlabel metal2 1395 -3450 1395 -3450 0 net=8497
rlabel metal2 240 -3452 240 -3452 0 net=2433
rlabel metal2 268 -3452 268 -3452 0 net=2446
rlabel metal2 292 -3452 292 -3452 0 net=2073
rlabel metal2 373 -3452 373 -3452 0 net=1769
rlabel metal2 408 -3452 408 -3452 0 net=3751
rlabel metal2 422 -3452 422 -3452 0 net=2788
rlabel metal2 541 -3452 541 -3452 0 net=11549
rlabel metal2 625 -3452 625 -3452 0 net=7241
rlabel metal2 646 -3452 646 -3452 0 net=6569
rlabel metal2 646 -3452 646 -3452 0 net=6569
rlabel metal2 653 -3452 653 -3452 0 net=6597
rlabel metal2 653 -3452 653 -3452 0 net=6597
rlabel metal2 674 -3452 674 -3452 0 net=9398
rlabel metal2 695 -3452 695 -3452 0 net=6871
rlabel metal2 719 -3452 719 -3452 0 net=8596
rlabel metal2 824 -3452 824 -3452 0 net=400
rlabel metal2 275 -3454 275 -3454 0 net=9392
rlabel metal2 317 -3454 317 -3454 0 net=1904
rlabel metal2 345 -3454 345 -3454 0 net=2249
rlabel metal2 394 -3454 394 -3454 0 net=3196
rlabel metal2 569 -3454 569 -3454 0 net=7765
rlabel metal2 667 -3454 667 -3454 0 net=5313
rlabel metal2 681 -3454 681 -3454 0 net=5208
rlabel metal2 835 -3454 835 -3454 0 net=9273
rlabel metal2 940 -3454 940 -3454 0 net=8743
rlabel metal2 940 -3454 940 -3454 0 net=8743
rlabel metal2 947 -3454 947 -3454 0 net=8546
rlabel metal2 282 -3456 282 -3456 0 net=1677
rlabel metal2 310 -3456 310 -3456 0 net=1633
rlabel metal2 387 -3456 387 -3456 0 net=1825
rlabel metal2 422 -3456 422 -3456 0 net=4690
rlabel metal2 443 -3456 443 -3456 0 net=9443
rlabel metal2 443 -3456 443 -3456 0 net=9443
rlabel metal2 450 -3456 450 -3456 0 net=1714
rlabel metal2 576 -3456 576 -3456 0 net=12693
rlabel metal2 660 -3456 660 -3456 0 net=11297
rlabel metal2 688 -3456 688 -3456 0 net=8942
rlabel metal2 821 -3456 821 -3456 0 net=3791
rlabel metal2 842 -3456 842 -3456 0 net=11659
rlabel metal2 842 -3456 842 -3456 0 net=11659
rlabel metal2 849 -3456 849 -3456 0 net=8694
rlabel metal2 296 -3458 296 -3458 0 net=3485
rlabel metal2 425 -3458 425 -3458 0 net=1140
rlabel metal2 660 -3458 660 -3458 0 net=9819
rlabel metal2 863 -3458 863 -3458 0 net=11821
rlabel metal2 429 -3460 429 -3460 0 net=3903
rlabel metal2 555 -3460 555 -3460 0 net=8749
rlabel metal2 695 -3460 695 -3460 0 net=6901
rlabel metal2 555 -3462 555 -3462 0 net=9467
rlabel metal2 534 -3464 534 -3464 0 net=9859
rlabel metal2 261 -3475 261 -3475 0 net=4405
rlabel metal2 303 -3475 303 -3475 0 net=1679
rlabel metal2 317 -3475 317 -3475 0 net=1634
rlabel metal2 331 -3475 331 -3475 0 net=3487
rlabel metal2 331 -3475 331 -3475 0 net=3487
rlabel metal2 338 -3475 338 -3475 0 net=3879
rlabel metal2 338 -3475 338 -3475 0 net=3879
rlabel metal2 352 -3475 352 -3475 0 net=2251
rlabel metal2 352 -3475 352 -3475 0 net=2251
rlabel metal2 380 -3475 380 -3475 0 net=2624
rlabel metal2 415 -3475 415 -3475 0 net=3752
rlabel metal2 467 -3475 467 -3475 0 net=2690
rlabel metal2 541 -3475 541 -3475 0 net=11551
rlabel metal2 541 -3475 541 -3475 0 net=11551
rlabel metal2 548 -3475 548 -3475 0 net=12023
rlabel metal2 569 -3475 569 -3475 0 net=7767
rlabel metal2 569 -3475 569 -3475 0 net=7767
rlabel metal2 583 -3475 583 -3475 0 net=12695
rlabel metal2 597 -3475 597 -3475 0 net=9820
rlabel metal2 681 -3475 681 -3475 0 net=11299
rlabel metal2 695 -3475 695 -3475 0 net=5377
rlabel metal2 835 -3475 835 -3475 0 net=3793
rlabel metal2 835 -3475 835 -3475 0 net=3793
rlabel metal2 842 -3475 842 -3475 0 net=11661
rlabel metal2 852 -3475 852 -3475 0 net=6306
rlabel metal2 870 -3475 870 -3475 0 net=11822
rlabel metal2 891 -3475 891 -3475 0 net=9274
rlabel metal2 989 -3475 989 -3475 0 net=11430
rlabel metal2 996 -3475 996 -3475 0 net=5659
rlabel metal2 996 -3475 996 -3475 0 net=5659
rlabel metal2 1066 -3475 1066 -3475 0 net=4783
rlabel metal2 1115 -3475 1115 -3475 0 net=2723
rlabel metal2 1213 -3475 1213 -3475 0 net=10902
rlabel metal2 1353 -3475 1353 -3475 0 net=12421
rlabel metal2 1353 -3475 1353 -3475 0 net=12421
rlabel metal2 1360 -3475 1360 -3475 0 net=11633
rlabel metal2 1360 -3475 1360 -3475 0 net=11633
rlabel metal2 1409 -3475 1409 -3475 0 net=8499
rlabel metal2 254 -3477 254 -3477 0 net=2435
rlabel metal2 394 -3477 394 -3477 0 net=1826
rlabel metal2 418 -3477 418 -3477 0 net=1400
rlabel metal2 709 -3477 709 -3477 0 net=6873
rlabel metal2 726 -3477 726 -3477 0 net=7966
rlabel metal2 758 -3477 758 -3477 0 net=6902
rlabel metal2 877 -3477 877 -3477 0 net=11341
rlabel metal2 905 -3477 905 -3477 0 net=10553
rlabel metal2 940 -3477 940 -3477 0 net=8745
rlabel metal2 940 -3477 940 -3477 0 net=8745
rlabel metal2 1115 -3477 1115 -3477 0 net=11520
rlabel metal2 1220 -3477 1220 -3477 0 net=4508
rlabel metal2 1409 -3477 1409 -3477 0 net=12668
rlabel metal2 401 -3479 401 -3479 0 net=1771
rlabel metal2 429 -3479 429 -3479 0 net=3904
rlabel metal2 471 -3479 471 -3479 0 net=3262
rlabel metal2 548 -3479 548 -3479 0 net=9469
rlabel metal2 576 -3479 576 -3479 0 net=8751
rlabel metal2 604 -3479 604 -3479 0 net=6274
rlabel metal2 646 -3479 646 -3479 0 net=6571
rlabel metal2 674 -3479 674 -3479 0 net=5315
rlabel metal2 884 -3479 884 -3479 0 net=3736
rlabel metal2 884 -3479 884 -3479 0 net=3736
rlabel metal2 912 -3479 912 -3479 0 net=11939
rlabel metal2 912 -3479 912 -3479 0 net=11939
rlabel metal2 919 -3479 919 -3479 0 net=8453
rlabel metal2 919 -3479 919 -3479 0 net=8453
rlabel metal2 926 -3479 926 -3479 0 net=9097
rlabel metal2 926 -3479 926 -3479 0 net=9097
rlabel metal2 359 -3481 359 -3481 0 net=2074
rlabel metal2 436 -3481 436 -3481 0 net=9445
rlabel metal2 478 -3481 478 -3481 0 net=4646
rlabel metal2 513 -3481 513 -3481 0 net=217
rlabel metal2 653 -3481 653 -3481 0 net=6599
rlabel metal2 653 -3481 653 -3481 0 net=6599
rlabel metal2 1412 -3481 1412 -3481 0 net=1
rlabel metal2 478 -3483 478 -3483 0 net=5351
rlabel metal2 485 -3485 485 -3485 0 net=4538
rlabel metal2 562 -3485 562 -3485 0 net=9861
rlabel metal2 611 -3485 611 -3485 0 net=7242
rlabel metal2 492 -3487 492 -3487 0 net=5062
rlabel metal2 261 -3498 261 -3498 0 net=2436
rlabel metal2 310 -3498 310 -3498 0 net=1680
rlabel metal2 331 -3498 331 -3498 0 net=3488
rlabel metal2 352 -3498 352 -3498 0 net=2253
rlabel metal2 408 -3498 408 -3498 0 net=1772
rlabel metal2 429 -3498 429 -3498 0 net=9446
rlabel metal2 541 -3498 541 -3498 0 net=11552
rlabel metal2 555 -3498 555 -3498 0 net=12024
rlabel metal2 569 -3498 569 -3498 0 net=7769
rlabel metal2 569 -3498 569 -3498 0 net=7769
rlabel metal2 583 -3498 583 -3498 0 net=8752
rlabel metal2 646 -3498 646 -3498 0 net=6600
rlabel metal2 660 -3498 660 -3498 0 net=6573
rlabel metal2 681 -3498 681 -3498 0 net=5316
rlabel metal2 716 -3498 716 -3498 0 net=6874
rlabel metal2 828 -3498 828 -3498 0 net=5379
rlabel metal2 877 -3498 877 -3498 0 net=11343
rlabel metal2 877 -3498 877 -3498 0 net=11343
rlabel metal2 898 -3498 898 -3498 0 net=10554
rlabel metal2 912 -3498 912 -3498 0 net=11940
rlabel metal2 912 -3498 912 -3498 0 net=11940
rlabel metal2 919 -3498 919 -3498 0 net=8454
rlabel metal2 919 -3498 919 -3498 0 net=8454
rlabel metal2 922 -3498 922 -3498 0 net=9098
rlabel metal2 940 -3498 940 -3498 0 net=8746
rlabel metal2 989 -3498 989 -3498 0 net=5660
rlabel metal2 1094 -3498 1094 -3498 0 net=4784
rlabel metal2 1118 -3498 1118 -3498 0 net=2724
rlabel metal2 1353 -3498 1353 -3498 0 net=12423
rlabel metal2 1353 -3498 1353 -3498 0 net=12423
rlabel metal2 1360 -3498 1360 -3498 0 net=11635
rlabel metal2 1412 -3498 1412 -3498 0 net=8500
rlabel metal2 268 -3500 268 -3500 0 net=4407
rlabel metal2 331 -3500 331 -3500 0 net=3881
rlabel metal2 355 -3500 355 -3500 0 net=5352
rlabel metal2 541 -3500 541 -3500 0 net=9471
rlabel metal2 576 -3500 576 -3500 0 net=9863
rlabel metal2 688 -3500 688 -3500 0 net=11300
rlabel metal2 688 -3500 688 -3500 0 net=11300
rlabel metal2 835 -3500 835 -3500 0 net=3794
rlabel metal2 576 -3502 576 -3502 0 net=12696
rlabel metal2 842 -3502 842 -3502 0 net=11662
rlabel metal2 271 -3513 271 -3513 0 net=4408
rlabel metal2 327 -3513 327 -3513 0 net=3882
rlabel metal2 355 -3513 355 -3513 0 net=2254
rlabel metal2 541 -3513 541 -3513 0 net=9472
rlabel metal2 565 -3513 565 -3513 0 net=7770
rlabel metal2 579 -3513 579 -3513 0 net=9864
rlabel metal2 660 -3513 660 -3513 0 net=6574
rlabel metal2 856 -3513 856 -3513 0 net=11344
rlabel metal2 1353 -3513 1353 -3513 0 net=12424
rlabel metal2 1363 -3513 1363 -3513 0 net=11636
rlabel metal2 870 -3515 870 -3515 0 net=5380
<< end >>
