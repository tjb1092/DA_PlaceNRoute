magic
tech scmos
timestamp 1555071785 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 36 -10 42 -4
rect 43 -10 49 -4
rect 50 -10 56 -4
rect 57 -10 63 -4
rect 64 -10 70 -4
rect 134 -10 140 -4
rect 141 -10 147 -4
rect 148 -10 151 -4
rect 176 -10 179 -4
rect 183 -10 189 -4
rect 190 -10 196 -4
rect 197 -10 200 -4
rect 204 -10 210 -4
rect 211 -10 217 -4
rect 218 -10 221 -4
rect 225 -10 231 -4
rect 232 -10 238 -4
rect 239 -10 242 -4
rect 1 -29 7 -23
rect 8 -29 14 -23
rect 15 -29 21 -23
rect 22 -29 28 -23
rect 29 -29 35 -23
rect 36 -29 42 -23
rect 43 -29 49 -23
rect 50 -29 56 -23
rect 57 -29 63 -23
rect 64 -29 70 -23
rect 127 -29 133 -23
rect 134 -29 137 -23
rect 141 -29 144 -23
rect 148 -29 154 -23
rect 155 -29 161 -23
rect 162 -29 165 -23
rect 169 -29 175 -23
rect 176 -29 179 -23
rect 183 -29 189 -23
rect 190 -29 196 -23
rect 197 -29 200 -23
rect 204 -29 207 -23
rect 211 -29 217 -23
rect 218 -29 224 -23
rect 225 -29 231 -23
rect 232 -29 235 -23
rect 239 -29 242 -23
rect 246 -29 252 -23
rect 253 -29 259 -23
rect 295 -29 301 -23
rect 323 -29 329 -23
rect 330 -29 333 -23
rect 1 -56 7 -50
rect 8 -56 14 -50
rect 15 -56 21 -50
rect 22 -56 28 -50
rect 29 -56 35 -50
rect 36 -56 42 -50
rect 43 -56 49 -50
rect 50 -56 56 -50
rect 57 -56 63 -50
rect 64 -56 70 -50
rect 71 -56 77 -50
rect 134 -56 137 -50
rect 141 -56 147 -50
rect 148 -56 154 -50
rect 155 -56 161 -50
rect 162 -56 168 -50
rect 169 -56 175 -50
rect 176 -56 182 -50
rect 183 -56 186 -50
rect 190 -56 193 -50
rect 197 -56 203 -50
rect 204 -56 210 -50
rect 211 -56 214 -50
rect 218 -56 224 -50
rect 225 -56 231 -50
rect 232 -56 235 -50
rect 239 -56 242 -50
rect 246 -56 249 -50
rect 253 -56 259 -50
rect 260 -56 263 -50
rect 267 -56 273 -50
rect 274 -56 280 -50
rect 281 -56 284 -50
rect 288 -56 291 -50
rect 295 -56 301 -50
rect 302 -56 305 -50
rect 323 -56 326 -50
rect 330 -56 333 -50
rect 1 -79 7 -73
rect 8 -79 14 -73
rect 15 -79 21 -73
rect 22 -79 28 -73
rect 29 -79 35 -73
rect 36 -79 42 -73
rect 43 -79 49 -73
rect 50 -79 56 -73
rect 85 -79 91 -73
rect 99 -79 105 -73
rect 106 -79 109 -73
rect 113 -79 119 -73
rect 120 -79 123 -73
rect 127 -79 130 -73
rect 134 -79 140 -73
rect 141 -79 147 -73
rect 148 -79 151 -73
rect 155 -79 161 -73
rect 162 -79 168 -73
rect 169 -79 172 -73
rect 176 -79 179 -73
rect 183 -79 189 -73
rect 190 -79 193 -73
rect 197 -79 203 -73
rect 204 -79 207 -73
rect 211 -79 217 -73
rect 218 -79 224 -73
rect 225 -79 231 -73
rect 232 -79 238 -73
rect 239 -79 242 -73
rect 246 -79 252 -73
rect 253 -79 256 -73
rect 260 -79 263 -73
rect 267 -79 273 -73
rect 274 -79 277 -73
rect 281 -79 284 -73
rect 288 -79 294 -73
rect 295 -79 298 -73
rect 302 -79 308 -73
rect 309 -79 315 -73
rect 316 -79 322 -73
rect 323 -79 326 -73
rect 330 -79 333 -73
rect 1 -104 7 -98
rect 8 -104 14 -98
rect 15 -104 21 -98
rect 22 -104 28 -98
rect 29 -104 35 -98
rect 36 -104 42 -98
rect 43 -104 49 -98
rect 50 -104 56 -98
rect 85 -104 91 -98
rect 99 -104 105 -98
rect 106 -104 109 -98
rect 113 -104 116 -98
rect 120 -104 126 -98
rect 127 -104 133 -98
rect 134 -104 137 -98
rect 141 -104 147 -98
rect 148 -104 151 -98
rect 155 -104 161 -98
rect 162 -104 168 -98
rect 169 -104 175 -98
rect 176 -104 182 -98
rect 183 -104 186 -98
rect 190 -104 196 -98
rect 197 -104 200 -98
rect 204 -104 210 -98
rect 211 -104 217 -98
rect 218 -104 224 -98
rect 225 -104 231 -98
rect 232 -104 235 -98
rect 239 -104 245 -98
rect 246 -104 249 -98
rect 253 -104 256 -98
rect 260 -104 263 -98
rect 267 -104 273 -98
rect 274 -104 277 -98
rect 281 -104 287 -98
rect 288 -104 294 -98
rect 295 -104 298 -98
rect 302 -104 305 -98
rect 309 -104 312 -98
rect 316 -104 319 -98
rect 323 -104 329 -98
rect 379 -104 385 -98
rect 1 -129 7 -123
rect 8 -129 14 -123
rect 15 -129 21 -123
rect 22 -129 28 -123
rect 29 -129 35 -123
rect 36 -129 42 -123
rect 43 -129 49 -123
rect 78 -129 84 -123
rect 85 -129 91 -123
rect 99 -129 105 -123
rect 106 -129 109 -123
rect 113 -129 119 -123
rect 120 -129 126 -123
rect 127 -129 133 -123
rect 134 -129 137 -123
rect 141 -129 147 -123
rect 148 -129 154 -123
rect 155 -129 158 -123
rect 162 -129 165 -123
rect 169 -129 175 -123
rect 176 -129 182 -123
rect 183 -129 186 -123
rect 190 -129 196 -123
rect 197 -129 200 -123
rect 204 -129 207 -123
rect 211 -129 217 -123
rect 218 -129 221 -123
rect 225 -129 231 -123
rect 232 -129 238 -123
rect 239 -129 242 -123
rect 253 -129 256 -123
rect 260 -129 263 -123
rect 267 -129 270 -123
rect 295 -129 301 -123
rect 302 -129 305 -123
rect 309 -129 315 -123
rect 316 -129 319 -123
rect 379 -129 382 -123
rect 1 -154 7 -148
rect 8 -154 14 -148
rect 15 -154 21 -148
rect 22 -154 28 -148
rect 29 -154 35 -148
rect 36 -154 42 -148
rect 43 -154 49 -148
rect 78 -154 84 -148
rect 106 -154 109 -148
rect 113 -154 116 -148
rect 120 -154 123 -148
rect 127 -154 133 -148
rect 134 -154 140 -148
rect 141 -154 147 -148
rect 148 -154 154 -148
rect 155 -154 161 -148
rect 162 -154 165 -148
rect 169 -154 175 -148
rect 176 -154 179 -148
rect 183 -154 189 -148
rect 190 -154 193 -148
rect 197 -154 203 -148
rect 204 -154 210 -148
rect 211 -154 217 -148
rect 218 -154 221 -148
rect 225 -154 228 -148
rect 232 -154 235 -148
rect 239 -154 245 -148
rect 253 -154 259 -148
rect 260 -154 263 -148
rect 267 -154 273 -148
rect 274 -154 277 -148
rect 309 -154 315 -148
rect 316 -154 322 -148
rect 323 -154 326 -148
rect 379 -154 385 -148
rect 386 -154 389 -148
rect 1 -177 7 -171
rect 8 -177 14 -171
rect 15 -177 21 -171
rect 22 -177 28 -171
rect 29 -177 35 -171
rect 78 -177 84 -171
rect 113 -177 119 -171
rect 120 -177 126 -171
rect 127 -177 133 -171
rect 134 -177 137 -171
rect 141 -177 147 -171
rect 148 -177 154 -171
rect 155 -177 161 -171
rect 162 -177 165 -171
rect 169 -177 172 -171
rect 176 -177 179 -171
rect 183 -177 189 -171
rect 190 -177 196 -171
rect 197 -177 200 -171
rect 204 -177 207 -171
rect 211 -177 217 -171
rect 218 -177 221 -171
rect 225 -177 231 -171
rect 232 -177 238 -171
rect 239 -177 242 -171
rect 246 -177 249 -171
rect 253 -177 256 -171
rect 260 -177 263 -171
rect 267 -177 273 -171
rect 274 -177 280 -171
rect 281 -177 287 -171
rect 288 -177 291 -171
rect 295 -177 298 -171
rect 302 -177 305 -171
rect 309 -177 315 -171
rect 316 -177 319 -171
rect 323 -177 326 -171
rect 330 -177 333 -171
rect 337 -177 343 -171
rect 344 -177 347 -171
rect 351 -177 357 -171
rect 358 -177 364 -171
rect 365 -177 368 -171
rect 372 -177 375 -171
rect 379 -177 385 -171
rect 386 -177 389 -171
rect 393 -177 396 -171
rect 407 -177 413 -171
rect 414 -177 417 -171
rect 435 -177 441 -171
rect 442 -177 445 -171
rect 1 -204 7 -198
rect 8 -204 14 -198
rect 15 -204 21 -198
rect 22 -204 28 -198
rect 71 -204 77 -198
rect 78 -204 81 -198
rect 85 -204 91 -198
rect 92 -204 98 -198
rect 99 -204 105 -198
rect 106 -204 109 -198
rect 113 -204 119 -198
rect 120 -204 123 -198
rect 127 -204 133 -198
rect 134 -204 140 -198
rect 141 -204 147 -198
rect 148 -204 151 -198
rect 155 -204 158 -198
rect 162 -204 165 -198
rect 169 -204 172 -198
rect 176 -204 179 -198
rect 183 -204 186 -198
rect 190 -204 193 -198
rect 197 -204 203 -198
rect 204 -204 210 -198
rect 211 -204 217 -198
rect 218 -204 224 -198
rect 225 -204 231 -198
rect 232 -204 235 -198
rect 239 -204 242 -198
rect 246 -204 252 -198
rect 253 -204 256 -198
rect 260 -204 266 -198
rect 267 -204 270 -198
rect 274 -204 277 -198
rect 281 -204 287 -198
rect 288 -204 291 -198
rect 295 -204 298 -198
rect 302 -204 308 -198
rect 309 -204 312 -198
rect 316 -204 319 -198
rect 323 -204 326 -198
rect 330 -204 333 -198
rect 337 -204 340 -198
rect 344 -204 347 -198
rect 351 -204 354 -198
rect 358 -204 361 -198
rect 365 -204 371 -198
rect 372 -204 375 -198
rect 379 -204 385 -198
rect 393 -204 396 -198
rect 400 -204 406 -198
rect 407 -204 410 -198
rect 414 -204 417 -198
rect 421 -204 427 -198
rect 428 -204 434 -198
rect 435 -204 438 -198
rect 442 -204 448 -198
rect 1 -237 7 -231
rect 8 -237 14 -231
rect 15 -237 21 -231
rect 22 -237 28 -231
rect 29 -237 35 -231
rect 64 -237 70 -231
rect 71 -237 77 -231
rect 78 -237 81 -231
rect 85 -237 88 -231
rect 92 -237 95 -231
rect 99 -237 102 -231
rect 106 -237 109 -231
rect 113 -237 116 -231
rect 120 -237 123 -231
rect 127 -237 130 -231
rect 134 -237 140 -231
rect 141 -237 144 -231
rect 148 -237 154 -231
rect 155 -237 161 -231
rect 162 -237 168 -231
rect 169 -237 172 -231
rect 176 -237 182 -231
rect 183 -237 189 -231
rect 190 -237 193 -231
rect 197 -237 203 -231
rect 204 -237 210 -231
rect 211 -237 214 -231
rect 218 -237 224 -231
rect 225 -237 231 -231
rect 232 -237 238 -231
rect 239 -237 245 -231
rect 246 -237 252 -231
rect 253 -237 259 -231
rect 260 -237 266 -231
rect 267 -237 270 -231
rect 274 -237 277 -231
rect 281 -237 284 -231
rect 288 -237 291 -231
rect 295 -237 298 -231
rect 302 -237 305 -231
rect 309 -237 312 -231
rect 316 -237 319 -231
rect 323 -237 329 -231
rect 330 -237 333 -231
rect 337 -237 340 -231
rect 344 -237 347 -231
rect 351 -237 354 -231
rect 358 -237 361 -231
rect 365 -237 371 -231
rect 372 -237 375 -231
rect 379 -237 385 -231
rect 386 -237 389 -231
rect 414 -237 420 -231
rect 421 -237 424 -231
rect 435 -237 441 -231
rect 1 -280 7 -274
rect 8 -280 14 -274
rect 15 -280 21 -274
rect 22 -280 28 -274
rect 29 -280 35 -274
rect 36 -280 42 -274
rect 50 -280 56 -274
rect 71 -280 77 -274
rect 78 -280 81 -274
rect 85 -280 91 -274
rect 92 -280 95 -274
rect 99 -280 105 -274
rect 106 -280 109 -274
rect 113 -280 116 -274
rect 120 -280 126 -274
rect 127 -280 133 -274
rect 134 -280 140 -274
rect 141 -280 147 -274
rect 148 -280 154 -274
rect 155 -280 158 -274
rect 162 -280 165 -274
rect 169 -280 172 -274
rect 176 -280 179 -274
rect 183 -280 189 -274
rect 190 -280 196 -274
rect 197 -280 200 -274
rect 204 -280 210 -274
rect 211 -280 217 -274
rect 218 -280 224 -274
rect 225 -280 231 -274
rect 232 -280 235 -274
rect 239 -280 242 -274
rect 246 -280 249 -274
rect 253 -280 259 -274
rect 260 -280 263 -274
rect 267 -280 273 -274
rect 274 -280 277 -274
rect 281 -280 284 -274
rect 288 -280 294 -274
rect 295 -280 301 -274
rect 302 -280 308 -274
rect 309 -280 312 -274
rect 316 -280 319 -274
rect 323 -280 326 -274
rect 330 -280 333 -274
rect 337 -280 340 -274
rect 344 -280 347 -274
rect 351 -280 354 -274
rect 358 -280 361 -274
rect 365 -280 368 -274
rect 372 -280 375 -274
rect 379 -280 382 -274
rect 386 -280 389 -274
rect 393 -280 396 -274
rect 400 -280 403 -274
rect 407 -280 410 -274
rect 414 -280 420 -274
rect 421 -280 424 -274
rect 428 -280 431 -274
rect 435 -280 441 -274
rect 442 -280 445 -274
rect 449 -280 455 -274
rect 456 -280 459 -274
rect 526 -280 532 -274
rect 533 -280 536 -274
rect 1 -321 7 -315
rect 8 -321 14 -315
rect 15 -321 21 -315
rect 29 -321 35 -315
rect 43 -321 49 -315
rect 50 -321 56 -315
rect 57 -321 60 -315
rect 64 -321 70 -315
rect 71 -321 77 -315
rect 78 -321 84 -315
rect 85 -321 88 -315
rect 92 -321 95 -315
rect 99 -321 102 -315
rect 106 -321 112 -315
rect 113 -321 116 -315
rect 120 -321 123 -315
rect 127 -321 130 -315
rect 134 -321 137 -315
rect 141 -321 147 -315
rect 148 -321 154 -315
rect 155 -321 161 -315
rect 162 -321 165 -315
rect 169 -321 175 -315
rect 176 -321 179 -315
rect 183 -321 186 -315
rect 190 -321 196 -315
rect 197 -321 200 -315
rect 204 -321 210 -315
rect 211 -321 214 -315
rect 218 -321 221 -315
rect 225 -321 231 -315
rect 232 -321 235 -315
rect 239 -321 245 -315
rect 246 -321 252 -315
rect 253 -321 259 -315
rect 260 -321 266 -315
rect 267 -321 270 -315
rect 274 -321 277 -315
rect 281 -321 287 -315
rect 288 -321 291 -315
rect 295 -321 301 -315
rect 302 -321 305 -315
rect 309 -321 312 -315
rect 316 -321 319 -315
rect 323 -321 329 -315
rect 330 -321 333 -315
rect 337 -321 340 -315
rect 344 -321 347 -315
rect 351 -321 354 -315
rect 358 -321 361 -315
rect 365 -321 368 -315
rect 372 -321 378 -315
rect 379 -321 382 -315
rect 386 -321 389 -315
rect 393 -321 396 -315
rect 400 -321 403 -315
rect 407 -321 410 -315
rect 414 -321 420 -315
rect 421 -321 424 -315
rect 428 -321 434 -315
rect 435 -321 438 -315
rect 449 -321 455 -315
rect 519 -321 525 -315
rect 526 -321 529 -315
rect 1 -368 7 -362
rect 8 -368 14 -362
rect 15 -368 21 -362
rect 22 -368 28 -362
rect 29 -368 35 -362
rect 36 -368 39 -362
rect 43 -368 46 -362
rect 50 -368 53 -362
rect 57 -368 60 -362
rect 64 -368 67 -362
rect 71 -368 74 -362
rect 78 -368 84 -362
rect 85 -368 91 -362
rect 92 -368 98 -362
rect 99 -368 102 -362
rect 106 -368 112 -362
rect 113 -368 119 -362
rect 120 -368 126 -362
rect 127 -368 133 -362
rect 134 -368 140 -362
rect 141 -368 147 -362
rect 148 -368 151 -362
rect 155 -368 158 -362
rect 162 -368 168 -362
rect 169 -368 175 -362
rect 176 -368 179 -362
rect 183 -368 186 -362
rect 190 -368 196 -362
rect 197 -368 203 -362
rect 204 -368 207 -362
rect 211 -368 217 -362
rect 218 -368 221 -362
rect 225 -368 228 -362
rect 232 -368 235 -362
rect 239 -368 245 -362
rect 246 -368 252 -362
rect 253 -368 259 -362
rect 260 -368 266 -362
rect 267 -368 273 -362
rect 274 -368 280 -362
rect 281 -368 287 -362
rect 288 -368 291 -362
rect 295 -368 298 -362
rect 302 -368 308 -362
rect 309 -368 312 -362
rect 316 -368 322 -362
rect 323 -368 329 -362
rect 330 -368 333 -362
rect 337 -368 340 -362
rect 344 -368 347 -362
rect 351 -368 354 -362
rect 358 -368 361 -362
rect 365 -368 368 -362
rect 372 -368 375 -362
rect 379 -368 382 -362
rect 386 -368 392 -362
rect 393 -368 396 -362
rect 400 -368 403 -362
rect 407 -368 410 -362
rect 414 -368 417 -362
rect 421 -368 424 -362
rect 428 -368 431 -362
rect 435 -368 438 -362
rect 442 -368 445 -362
rect 449 -368 452 -362
rect 456 -368 459 -362
rect 463 -368 469 -362
rect 470 -368 473 -362
rect 512 -368 515 -362
rect 1 -419 7 -413
rect 15 -419 21 -413
rect 22 -419 25 -413
rect 29 -419 32 -413
rect 36 -419 42 -413
rect 43 -419 49 -413
rect 50 -419 56 -413
rect 57 -419 63 -413
rect 64 -419 70 -413
rect 71 -419 74 -413
rect 78 -419 81 -413
rect 85 -419 88 -413
rect 92 -419 95 -413
rect 99 -419 105 -413
rect 106 -419 112 -413
rect 113 -419 116 -413
rect 120 -419 123 -413
rect 127 -419 130 -413
rect 134 -419 140 -413
rect 141 -419 147 -413
rect 148 -419 154 -413
rect 155 -419 161 -413
rect 162 -419 168 -413
rect 169 -419 172 -413
rect 176 -419 179 -413
rect 183 -419 186 -413
rect 190 -419 196 -413
rect 197 -419 200 -413
rect 204 -419 210 -413
rect 211 -419 217 -413
rect 218 -419 221 -413
rect 225 -419 231 -413
rect 232 -419 235 -413
rect 239 -419 242 -413
rect 246 -419 249 -413
rect 253 -419 256 -413
rect 260 -419 266 -413
rect 267 -419 273 -413
rect 274 -419 277 -413
rect 281 -419 287 -413
rect 288 -419 291 -413
rect 295 -419 298 -413
rect 302 -419 305 -413
rect 309 -419 315 -413
rect 316 -419 322 -413
rect 323 -419 329 -413
rect 330 -419 333 -413
rect 337 -419 343 -413
rect 344 -419 350 -413
rect 351 -419 354 -413
rect 358 -419 361 -413
rect 365 -419 368 -413
rect 372 -419 375 -413
rect 379 -419 382 -413
rect 386 -419 389 -413
rect 393 -419 396 -413
rect 400 -419 403 -413
rect 407 -419 410 -413
rect 414 -419 420 -413
rect 421 -419 424 -413
rect 428 -419 431 -413
rect 435 -419 438 -413
rect 442 -419 445 -413
rect 449 -419 452 -413
rect 456 -419 459 -413
rect 463 -419 466 -413
rect 470 -419 473 -413
rect 477 -419 483 -413
rect 484 -419 490 -413
rect 491 -419 494 -413
rect 498 -419 501 -413
rect 505 -419 511 -413
rect 512 -419 515 -413
rect 519 -419 522 -413
rect 526 -419 529 -413
rect 1 -470 4 -464
rect 8 -470 11 -464
rect 15 -470 18 -464
rect 22 -470 28 -464
rect 29 -470 35 -464
rect 36 -470 39 -464
rect 43 -470 46 -464
rect 50 -470 56 -464
rect 57 -470 60 -464
rect 64 -470 67 -464
rect 71 -470 74 -464
rect 78 -470 81 -464
rect 85 -470 88 -464
rect 92 -470 98 -464
rect 99 -470 102 -464
rect 106 -470 109 -464
rect 113 -470 119 -464
rect 120 -470 126 -464
rect 127 -470 133 -464
rect 134 -470 137 -464
rect 141 -470 144 -464
rect 148 -470 154 -464
rect 155 -470 161 -464
rect 162 -470 168 -464
rect 169 -470 175 -464
rect 176 -470 179 -464
rect 183 -470 186 -464
rect 190 -470 196 -464
rect 197 -470 203 -464
rect 204 -470 207 -464
rect 211 -470 214 -464
rect 218 -470 224 -464
rect 225 -470 231 -464
rect 232 -470 235 -464
rect 239 -470 245 -464
rect 246 -470 249 -464
rect 253 -470 259 -464
rect 260 -470 266 -464
rect 267 -470 270 -464
rect 274 -470 280 -464
rect 281 -470 287 -464
rect 288 -470 291 -464
rect 295 -470 298 -464
rect 302 -470 305 -464
rect 309 -470 315 -464
rect 316 -470 322 -464
rect 323 -470 326 -464
rect 330 -470 333 -464
rect 337 -470 340 -464
rect 344 -470 350 -464
rect 351 -470 357 -464
rect 358 -470 364 -464
rect 365 -470 371 -464
rect 372 -470 378 -464
rect 379 -470 382 -464
rect 386 -470 389 -464
rect 393 -470 396 -464
rect 400 -470 403 -464
rect 407 -470 410 -464
rect 414 -470 417 -464
rect 421 -470 424 -464
rect 428 -470 431 -464
rect 435 -470 438 -464
rect 442 -470 445 -464
rect 449 -470 452 -464
rect 456 -470 459 -464
rect 463 -470 466 -464
rect 470 -470 473 -464
rect 477 -470 480 -464
rect 484 -470 487 -464
rect 491 -470 494 -464
rect 498 -470 501 -464
rect 505 -470 508 -464
rect 512 -470 515 -464
rect 519 -470 522 -464
rect 526 -470 529 -464
rect 533 -470 536 -464
rect 540 -470 543 -464
rect 547 -470 550 -464
rect 554 -470 560 -464
rect 561 -470 564 -464
rect 568 -470 574 -464
rect 575 -470 578 -464
rect 15 -527 18 -521
rect 22 -527 25 -521
rect 29 -527 32 -521
rect 36 -527 39 -521
rect 43 -527 46 -521
rect 50 -527 53 -521
rect 57 -527 60 -521
rect 64 -527 70 -521
rect 71 -527 77 -521
rect 78 -527 84 -521
rect 85 -527 91 -521
rect 92 -527 95 -521
rect 99 -527 102 -521
rect 106 -527 109 -521
rect 113 -527 119 -521
rect 120 -527 126 -521
rect 127 -527 133 -521
rect 134 -527 140 -521
rect 141 -527 147 -521
rect 148 -527 151 -521
rect 155 -527 161 -521
rect 162 -527 165 -521
rect 169 -527 172 -521
rect 176 -527 179 -521
rect 183 -527 189 -521
rect 190 -527 193 -521
rect 197 -527 203 -521
rect 204 -527 207 -521
rect 211 -527 214 -521
rect 218 -527 224 -521
rect 225 -527 231 -521
rect 232 -527 235 -521
rect 239 -527 245 -521
rect 246 -527 249 -521
rect 253 -527 256 -521
rect 260 -527 266 -521
rect 267 -527 270 -521
rect 274 -527 280 -521
rect 281 -527 287 -521
rect 288 -527 294 -521
rect 295 -527 301 -521
rect 302 -527 305 -521
rect 309 -527 315 -521
rect 316 -527 319 -521
rect 323 -527 329 -521
rect 330 -527 333 -521
rect 337 -527 340 -521
rect 344 -527 350 -521
rect 351 -527 357 -521
rect 358 -527 361 -521
rect 365 -527 371 -521
rect 372 -527 378 -521
rect 379 -527 382 -521
rect 386 -527 392 -521
rect 393 -527 396 -521
rect 400 -527 403 -521
rect 407 -527 410 -521
rect 414 -527 417 -521
rect 421 -527 427 -521
rect 428 -527 431 -521
rect 435 -527 438 -521
rect 442 -527 445 -521
rect 449 -527 452 -521
rect 456 -527 459 -521
rect 463 -527 466 -521
rect 470 -527 473 -521
rect 477 -527 480 -521
rect 484 -527 487 -521
rect 491 -527 494 -521
rect 498 -527 501 -521
rect 505 -527 511 -521
rect 512 -527 518 -521
rect 519 -527 522 -521
rect 540 -527 543 -521
rect 561 -527 564 -521
rect 8 -576 11 -570
rect 15 -576 21 -570
rect 22 -576 28 -570
rect 29 -576 32 -570
rect 36 -576 42 -570
rect 43 -576 49 -570
rect 50 -576 53 -570
rect 57 -576 63 -570
rect 64 -576 70 -570
rect 71 -576 74 -570
rect 78 -576 81 -570
rect 85 -576 91 -570
rect 92 -576 95 -570
rect 99 -576 105 -570
rect 106 -576 112 -570
rect 113 -576 119 -570
rect 120 -576 123 -570
rect 127 -576 130 -570
rect 134 -576 137 -570
rect 141 -576 144 -570
rect 148 -576 151 -570
rect 155 -576 158 -570
rect 162 -576 165 -570
rect 169 -576 175 -570
rect 176 -576 179 -570
rect 183 -576 189 -570
rect 190 -576 193 -570
rect 197 -576 200 -570
rect 204 -576 210 -570
rect 211 -576 217 -570
rect 218 -576 224 -570
rect 225 -576 231 -570
rect 232 -576 238 -570
rect 239 -576 245 -570
rect 246 -576 249 -570
rect 253 -576 259 -570
rect 260 -576 263 -570
rect 267 -576 273 -570
rect 274 -576 277 -570
rect 281 -576 287 -570
rect 288 -576 291 -570
rect 295 -576 298 -570
rect 302 -576 308 -570
rect 309 -576 315 -570
rect 316 -576 319 -570
rect 323 -576 326 -570
rect 330 -576 333 -570
rect 337 -576 343 -570
rect 344 -576 347 -570
rect 351 -576 354 -570
rect 358 -576 364 -570
rect 365 -576 371 -570
rect 372 -576 375 -570
rect 379 -576 382 -570
rect 386 -576 389 -570
rect 393 -576 396 -570
rect 400 -576 403 -570
rect 407 -576 410 -570
rect 414 -576 417 -570
rect 421 -576 424 -570
rect 428 -576 434 -570
rect 435 -576 438 -570
rect 442 -576 445 -570
rect 449 -576 452 -570
rect 456 -576 459 -570
rect 463 -576 466 -570
rect 470 -576 473 -570
rect 477 -576 480 -570
rect 484 -576 487 -570
rect 491 -576 494 -570
rect 498 -576 504 -570
rect 505 -576 508 -570
rect 512 -576 518 -570
rect 519 -576 522 -570
rect 526 -576 532 -570
rect 533 -576 536 -570
rect 540 -576 543 -570
rect 547 -576 553 -570
rect 554 -576 557 -570
rect 561 -576 564 -570
rect 8 -619 11 -613
rect 15 -619 18 -613
rect 22 -619 25 -613
rect 29 -619 32 -613
rect 36 -619 39 -613
rect 43 -619 49 -613
rect 50 -619 56 -613
rect 57 -619 60 -613
rect 64 -619 70 -613
rect 71 -619 74 -613
rect 78 -619 84 -613
rect 85 -619 91 -613
rect 92 -619 95 -613
rect 99 -619 105 -613
rect 106 -619 109 -613
rect 113 -619 119 -613
rect 120 -619 123 -613
rect 127 -619 133 -613
rect 134 -619 140 -613
rect 141 -619 147 -613
rect 148 -619 151 -613
rect 155 -619 158 -613
rect 162 -619 165 -613
rect 169 -619 172 -613
rect 176 -619 182 -613
rect 183 -619 189 -613
rect 190 -619 193 -613
rect 197 -619 200 -613
rect 204 -619 207 -613
rect 211 -619 217 -613
rect 218 -619 224 -613
rect 225 -619 231 -613
rect 232 -619 235 -613
rect 239 -619 242 -613
rect 246 -619 249 -613
rect 253 -619 256 -613
rect 260 -619 263 -613
rect 267 -619 270 -613
rect 274 -619 277 -613
rect 281 -619 284 -613
rect 288 -619 294 -613
rect 295 -619 301 -613
rect 302 -619 305 -613
rect 309 -619 315 -613
rect 316 -619 319 -613
rect 323 -619 329 -613
rect 330 -619 333 -613
rect 337 -619 343 -613
rect 344 -619 347 -613
rect 351 -619 357 -613
rect 358 -619 361 -613
rect 365 -619 368 -613
rect 372 -619 375 -613
rect 379 -619 382 -613
rect 386 -619 389 -613
rect 393 -619 399 -613
rect 400 -619 403 -613
rect 407 -619 410 -613
rect 414 -619 420 -613
rect 421 -619 424 -613
rect 428 -619 431 -613
rect 435 -619 438 -613
rect 442 -619 445 -613
rect 449 -619 452 -613
rect 456 -619 459 -613
rect 463 -619 466 -613
rect 470 -619 473 -613
rect 477 -619 483 -613
rect 484 -619 487 -613
rect 491 -619 494 -613
rect 498 -619 501 -613
rect 505 -619 511 -613
rect 512 -619 518 -613
rect 519 -619 525 -613
rect 526 -619 529 -613
rect 533 -619 536 -613
rect 540 -619 543 -613
rect 547 -619 550 -613
rect 554 -619 557 -613
rect 561 -619 567 -613
rect 36 -666 42 -660
rect 43 -666 46 -660
rect 50 -666 53 -660
rect 57 -666 63 -660
rect 64 -666 67 -660
rect 71 -666 77 -660
rect 78 -666 81 -660
rect 85 -666 88 -660
rect 92 -666 98 -660
rect 99 -666 105 -660
rect 106 -666 109 -660
rect 113 -666 119 -660
rect 120 -666 123 -660
rect 127 -666 133 -660
rect 134 -666 137 -660
rect 141 -666 147 -660
rect 148 -666 151 -660
rect 155 -666 158 -660
rect 162 -666 165 -660
rect 169 -666 175 -660
rect 176 -666 179 -660
rect 183 -666 186 -660
rect 190 -666 193 -660
rect 197 -666 203 -660
rect 204 -666 210 -660
rect 211 -666 214 -660
rect 218 -666 221 -660
rect 225 -666 228 -660
rect 232 -666 235 -660
rect 239 -666 245 -660
rect 246 -666 252 -660
rect 253 -666 256 -660
rect 260 -666 263 -660
rect 267 -666 273 -660
rect 274 -666 277 -660
rect 281 -666 284 -660
rect 288 -666 291 -660
rect 295 -666 298 -660
rect 302 -666 305 -660
rect 309 -666 312 -660
rect 316 -666 322 -660
rect 323 -666 326 -660
rect 330 -666 336 -660
rect 337 -666 343 -660
rect 344 -666 350 -660
rect 351 -666 357 -660
rect 358 -666 361 -660
rect 365 -666 368 -660
rect 372 -666 378 -660
rect 379 -666 382 -660
rect 386 -666 389 -660
rect 393 -666 399 -660
rect 400 -666 406 -660
rect 407 -666 410 -660
rect 414 -666 417 -660
rect 421 -666 424 -660
rect 428 -666 431 -660
rect 435 -666 438 -660
rect 442 -666 445 -660
rect 449 -666 452 -660
rect 456 -666 459 -660
rect 463 -666 466 -660
rect 470 -666 476 -660
rect 477 -666 480 -660
rect 484 -666 490 -660
rect 491 -666 494 -660
rect 498 -666 501 -660
rect 505 -666 508 -660
rect 512 -666 518 -660
rect 519 -666 522 -660
rect 526 -666 532 -660
rect 533 -666 536 -660
rect 540 -666 546 -660
rect 547 -666 550 -660
rect 554 -666 557 -660
rect 561 -666 567 -660
rect 582 -666 585 -660
rect 15 -715 18 -709
rect 22 -715 25 -709
rect 29 -715 35 -709
rect 36 -715 39 -709
rect 43 -715 46 -709
rect 50 -715 53 -709
rect 57 -715 63 -709
rect 64 -715 70 -709
rect 71 -715 77 -709
rect 78 -715 81 -709
rect 85 -715 88 -709
rect 92 -715 95 -709
rect 99 -715 105 -709
rect 106 -715 112 -709
rect 113 -715 116 -709
rect 120 -715 123 -709
rect 127 -715 130 -709
rect 134 -715 140 -709
rect 141 -715 144 -709
rect 148 -715 154 -709
rect 155 -715 158 -709
rect 162 -715 168 -709
rect 169 -715 172 -709
rect 176 -715 179 -709
rect 183 -715 189 -709
rect 190 -715 196 -709
rect 197 -715 203 -709
rect 204 -715 207 -709
rect 211 -715 214 -709
rect 218 -715 224 -709
rect 225 -715 228 -709
rect 232 -715 235 -709
rect 239 -715 242 -709
rect 246 -715 249 -709
rect 253 -715 256 -709
rect 260 -715 263 -709
rect 267 -715 270 -709
rect 274 -715 277 -709
rect 281 -715 287 -709
rect 288 -715 291 -709
rect 295 -715 301 -709
rect 302 -715 305 -709
rect 309 -715 315 -709
rect 316 -715 319 -709
rect 323 -715 326 -709
rect 330 -715 336 -709
rect 337 -715 343 -709
rect 344 -715 350 -709
rect 351 -715 354 -709
rect 358 -715 361 -709
rect 365 -715 368 -709
rect 372 -715 375 -709
rect 379 -715 385 -709
rect 386 -715 392 -709
rect 393 -715 399 -709
rect 400 -715 403 -709
rect 407 -715 410 -709
rect 414 -715 417 -709
rect 421 -715 427 -709
rect 428 -715 431 -709
rect 435 -715 438 -709
rect 442 -715 445 -709
rect 449 -715 452 -709
rect 456 -715 459 -709
rect 463 -715 466 -709
rect 470 -715 473 -709
rect 477 -715 480 -709
rect 484 -715 487 -709
rect 491 -715 497 -709
rect 498 -715 501 -709
rect 505 -715 508 -709
rect 512 -715 515 -709
rect 519 -715 522 -709
rect 526 -715 529 -709
rect 533 -715 536 -709
rect 540 -715 543 -709
rect 547 -715 550 -709
rect 554 -715 557 -709
rect 561 -715 564 -709
rect 568 -715 574 -709
rect 575 -715 578 -709
rect 582 -715 585 -709
rect 589 -715 595 -709
rect 596 -715 602 -709
rect 603 -715 606 -709
rect 610 -715 616 -709
rect 617 -715 620 -709
rect 624 -715 630 -709
rect 631 -715 634 -709
rect 638 -715 641 -709
rect 645 -715 648 -709
rect 29 -766 35 -760
rect 36 -766 42 -760
rect 43 -766 46 -760
rect 50 -766 53 -760
rect 57 -766 60 -760
rect 64 -766 67 -760
rect 71 -766 74 -760
rect 78 -766 81 -760
rect 85 -766 88 -760
rect 92 -766 95 -760
rect 99 -766 105 -760
rect 106 -766 109 -760
rect 113 -766 119 -760
rect 120 -766 123 -760
rect 127 -766 130 -760
rect 134 -766 140 -760
rect 141 -766 147 -760
rect 148 -766 154 -760
rect 155 -766 158 -760
rect 162 -766 165 -760
rect 169 -766 172 -760
rect 176 -766 179 -760
rect 183 -766 186 -760
rect 190 -766 196 -760
rect 197 -766 200 -760
rect 204 -766 210 -760
rect 211 -766 217 -760
rect 218 -766 224 -760
rect 225 -766 231 -760
rect 232 -766 235 -760
rect 239 -766 242 -760
rect 246 -766 252 -760
rect 253 -766 259 -760
rect 260 -766 263 -760
rect 267 -766 270 -760
rect 274 -766 280 -760
rect 281 -766 287 -760
rect 288 -766 294 -760
rect 295 -766 298 -760
rect 302 -766 308 -760
rect 309 -766 312 -760
rect 316 -766 319 -760
rect 323 -766 326 -760
rect 330 -766 336 -760
rect 337 -766 343 -760
rect 344 -766 350 -760
rect 351 -766 354 -760
rect 358 -766 364 -760
rect 365 -766 368 -760
rect 372 -766 378 -760
rect 379 -766 382 -760
rect 386 -766 389 -760
rect 393 -766 399 -760
rect 400 -766 403 -760
rect 407 -766 410 -760
rect 414 -766 417 -760
rect 421 -766 424 -760
rect 428 -766 431 -760
rect 435 -766 438 -760
rect 442 -766 448 -760
rect 449 -766 452 -760
rect 456 -766 459 -760
rect 463 -766 466 -760
rect 470 -766 476 -760
rect 477 -766 480 -760
rect 484 -766 490 -760
rect 491 -766 494 -760
rect 498 -766 501 -760
rect 505 -766 508 -760
rect 512 -766 515 -760
rect 519 -766 522 -760
rect 526 -766 532 -760
rect 533 -766 536 -760
rect 540 -766 543 -760
rect 554 -766 557 -760
rect 610 -766 616 -760
rect 22 -823 28 -817
rect 29 -823 35 -817
rect 36 -823 39 -817
rect 43 -823 46 -817
rect 50 -823 53 -817
rect 57 -823 63 -817
rect 64 -823 67 -817
rect 71 -823 77 -817
rect 78 -823 81 -817
rect 85 -823 88 -817
rect 92 -823 95 -817
rect 99 -823 105 -817
rect 106 -823 112 -817
rect 113 -823 119 -817
rect 120 -823 126 -817
rect 127 -823 130 -817
rect 134 -823 137 -817
rect 141 -823 147 -817
rect 148 -823 154 -817
rect 155 -823 161 -817
rect 162 -823 168 -817
rect 169 -823 172 -817
rect 176 -823 179 -817
rect 183 -823 189 -817
rect 190 -823 193 -817
rect 197 -823 203 -817
rect 204 -823 207 -817
rect 211 -823 217 -817
rect 218 -823 221 -817
rect 225 -823 228 -817
rect 232 -823 238 -817
rect 239 -823 242 -817
rect 246 -823 252 -817
rect 253 -823 259 -817
rect 260 -823 266 -817
rect 267 -823 270 -817
rect 274 -823 277 -817
rect 281 -823 284 -817
rect 288 -823 291 -817
rect 295 -823 301 -817
rect 302 -823 305 -817
rect 309 -823 315 -817
rect 316 -823 322 -817
rect 323 -823 326 -817
rect 330 -823 336 -817
rect 337 -823 340 -817
rect 344 -823 350 -817
rect 351 -823 357 -817
rect 358 -823 361 -817
rect 365 -823 368 -817
rect 372 -823 378 -817
rect 379 -823 382 -817
rect 386 -823 389 -817
rect 393 -823 396 -817
rect 400 -823 406 -817
rect 407 -823 410 -817
rect 414 -823 417 -817
rect 421 -823 424 -817
rect 428 -823 431 -817
rect 435 -823 438 -817
rect 442 -823 445 -817
rect 449 -823 452 -817
rect 456 -823 462 -817
rect 463 -823 466 -817
rect 470 -823 473 -817
rect 477 -823 480 -817
rect 484 -823 487 -817
rect 491 -823 494 -817
rect 498 -823 501 -817
rect 505 -823 508 -817
rect 512 -823 515 -817
rect 519 -823 522 -817
rect 526 -823 529 -817
rect 533 -823 536 -817
rect 540 -823 543 -817
rect 547 -823 550 -817
rect 554 -823 560 -817
rect 22 -886 28 -880
rect 29 -886 35 -880
rect 36 -886 42 -880
rect 43 -886 49 -880
rect 50 -886 53 -880
rect 57 -886 60 -880
rect 64 -886 67 -880
rect 71 -886 77 -880
rect 78 -886 81 -880
rect 85 -886 88 -880
rect 92 -886 95 -880
rect 99 -886 102 -880
rect 106 -886 109 -880
rect 113 -886 119 -880
rect 120 -886 126 -880
rect 127 -886 133 -880
rect 134 -886 140 -880
rect 141 -886 144 -880
rect 148 -886 151 -880
rect 155 -886 161 -880
rect 162 -886 168 -880
rect 169 -886 175 -880
rect 176 -886 182 -880
rect 183 -886 186 -880
rect 190 -886 196 -880
rect 197 -886 203 -880
rect 204 -886 210 -880
rect 211 -886 214 -880
rect 218 -886 221 -880
rect 225 -886 228 -880
rect 232 -886 235 -880
rect 239 -886 242 -880
rect 246 -886 249 -880
rect 253 -886 256 -880
rect 260 -886 263 -880
rect 267 -886 270 -880
rect 274 -886 277 -880
rect 281 -886 287 -880
rect 288 -886 291 -880
rect 295 -886 301 -880
rect 302 -886 308 -880
rect 309 -886 315 -880
rect 316 -886 319 -880
rect 323 -886 326 -880
rect 330 -886 336 -880
rect 337 -886 340 -880
rect 344 -886 350 -880
rect 351 -886 357 -880
rect 358 -886 361 -880
rect 365 -886 368 -880
rect 372 -886 378 -880
rect 379 -886 385 -880
rect 386 -886 389 -880
rect 393 -886 396 -880
rect 400 -886 403 -880
rect 407 -886 410 -880
rect 414 -886 417 -880
rect 421 -886 424 -880
rect 428 -886 431 -880
rect 435 -886 438 -880
rect 442 -886 445 -880
rect 449 -886 452 -880
rect 456 -886 459 -880
rect 463 -886 469 -880
rect 470 -886 476 -880
rect 477 -886 480 -880
rect 484 -886 487 -880
rect 491 -886 494 -880
rect 498 -886 501 -880
rect 505 -886 508 -880
rect 512 -886 515 -880
rect 519 -886 525 -880
rect 526 -886 529 -880
rect 533 -886 536 -880
rect 8 -941 11 -935
rect 15 -941 18 -935
rect 22 -941 25 -935
rect 29 -941 35 -935
rect 36 -941 39 -935
rect 43 -941 49 -935
rect 50 -941 53 -935
rect 57 -941 60 -935
rect 64 -941 67 -935
rect 71 -941 77 -935
rect 78 -941 84 -935
rect 85 -941 91 -935
rect 92 -941 95 -935
rect 99 -941 105 -935
rect 106 -941 109 -935
rect 113 -941 116 -935
rect 120 -941 123 -935
rect 127 -941 130 -935
rect 134 -941 140 -935
rect 141 -941 144 -935
rect 148 -941 154 -935
rect 155 -941 161 -935
rect 162 -941 168 -935
rect 169 -941 172 -935
rect 176 -941 179 -935
rect 183 -941 186 -935
rect 190 -941 196 -935
rect 197 -941 203 -935
rect 204 -941 210 -935
rect 211 -941 217 -935
rect 218 -941 224 -935
rect 225 -941 231 -935
rect 232 -941 235 -935
rect 239 -941 242 -935
rect 246 -941 249 -935
rect 253 -941 256 -935
rect 260 -941 266 -935
rect 267 -941 270 -935
rect 274 -941 277 -935
rect 281 -941 284 -935
rect 288 -941 294 -935
rect 295 -941 298 -935
rect 302 -941 308 -935
rect 309 -941 312 -935
rect 316 -941 319 -935
rect 323 -941 329 -935
rect 330 -941 336 -935
rect 337 -941 340 -935
rect 344 -941 347 -935
rect 351 -941 357 -935
rect 358 -941 361 -935
rect 365 -941 368 -935
rect 372 -941 375 -935
rect 379 -941 385 -935
rect 386 -941 389 -935
rect 393 -941 399 -935
rect 400 -941 403 -935
rect 407 -941 413 -935
rect 414 -941 417 -935
rect 421 -941 424 -935
rect 428 -941 431 -935
rect 435 -941 438 -935
rect 442 -941 448 -935
rect 449 -941 452 -935
rect 456 -941 459 -935
rect 463 -941 469 -935
rect 470 -941 473 -935
rect 477 -941 480 -935
rect 484 -941 487 -935
rect 491 -941 494 -935
rect 498 -941 501 -935
rect 505 -941 508 -935
rect 512 -941 515 -935
rect 519 -941 522 -935
rect 1 -990 4 -984
rect 8 -990 11 -984
rect 15 -990 21 -984
rect 22 -990 28 -984
rect 29 -990 35 -984
rect 36 -990 42 -984
rect 43 -990 46 -984
rect 50 -990 53 -984
rect 57 -990 63 -984
rect 64 -990 67 -984
rect 71 -990 77 -984
rect 78 -990 84 -984
rect 85 -990 88 -984
rect 92 -990 98 -984
rect 99 -990 105 -984
rect 106 -990 109 -984
rect 113 -990 116 -984
rect 120 -990 123 -984
rect 127 -990 133 -984
rect 134 -990 140 -984
rect 141 -990 144 -984
rect 148 -990 151 -984
rect 155 -990 161 -984
rect 162 -990 168 -984
rect 169 -990 172 -984
rect 176 -990 182 -984
rect 183 -990 189 -984
rect 190 -990 196 -984
rect 197 -990 203 -984
rect 204 -990 207 -984
rect 211 -990 214 -984
rect 218 -990 224 -984
rect 225 -990 231 -984
rect 232 -990 238 -984
rect 239 -990 245 -984
rect 246 -990 249 -984
rect 253 -990 259 -984
rect 260 -990 266 -984
rect 267 -990 270 -984
rect 274 -990 277 -984
rect 281 -990 284 -984
rect 288 -990 294 -984
rect 295 -990 301 -984
rect 302 -990 305 -984
rect 309 -990 312 -984
rect 316 -990 319 -984
rect 323 -990 326 -984
rect 330 -990 336 -984
rect 337 -990 343 -984
rect 344 -990 347 -984
rect 351 -990 357 -984
rect 358 -990 361 -984
rect 365 -990 368 -984
rect 372 -990 375 -984
rect 379 -990 382 -984
rect 386 -990 389 -984
rect 393 -990 396 -984
rect 400 -990 403 -984
rect 407 -990 410 -984
rect 414 -990 417 -984
rect 421 -990 424 -984
rect 428 -990 431 -984
rect 435 -990 438 -984
rect 442 -990 445 -984
rect 449 -990 452 -984
rect 456 -990 459 -984
rect 463 -990 469 -984
rect 470 -990 476 -984
rect 477 -990 480 -984
rect 491 -990 494 -984
rect 505 -990 508 -984
rect 15 -1037 21 -1031
rect 22 -1037 25 -1031
rect 29 -1037 35 -1031
rect 36 -1037 39 -1031
rect 43 -1037 49 -1031
rect 57 -1037 60 -1031
rect 78 -1037 84 -1031
rect 85 -1037 88 -1031
rect 92 -1037 98 -1031
rect 99 -1037 105 -1031
rect 106 -1037 109 -1031
rect 113 -1037 116 -1031
rect 120 -1037 123 -1031
rect 127 -1037 130 -1031
rect 134 -1037 140 -1031
rect 141 -1037 144 -1031
rect 148 -1037 154 -1031
rect 155 -1037 161 -1031
rect 162 -1037 168 -1031
rect 169 -1037 172 -1031
rect 176 -1037 179 -1031
rect 183 -1037 189 -1031
rect 190 -1037 193 -1031
rect 197 -1037 200 -1031
rect 204 -1037 207 -1031
rect 211 -1037 217 -1031
rect 218 -1037 224 -1031
rect 225 -1037 231 -1031
rect 232 -1037 235 -1031
rect 239 -1037 242 -1031
rect 246 -1037 249 -1031
rect 253 -1037 256 -1031
rect 260 -1037 263 -1031
rect 267 -1037 270 -1031
rect 274 -1037 280 -1031
rect 281 -1037 287 -1031
rect 288 -1037 291 -1031
rect 295 -1037 301 -1031
rect 302 -1037 308 -1031
rect 309 -1037 312 -1031
rect 316 -1037 319 -1031
rect 323 -1037 329 -1031
rect 330 -1037 336 -1031
rect 337 -1037 343 -1031
rect 344 -1037 347 -1031
rect 351 -1037 354 -1031
rect 358 -1037 361 -1031
rect 365 -1037 368 -1031
rect 372 -1037 375 -1031
rect 379 -1037 382 -1031
rect 386 -1037 389 -1031
rect 393 -1037 396 -1031
rect 400 -1037 403 -1031
rect 407 -1037 410 -1031
rect 414 -1037 420 -1031
rect 421 -1037 427 -1031
rect 428 -1037 431 -1031
rect 435 -1037 441 -1031
rect 442 -1037 448 -1031
rect 449 -1037 452 -1031
rect 456 -1037 462 -1031
rect 463 -1037 469 -1031
rect 470 -1037 473 -1031
rect 477 -1037 480 -1031
rect 484 -1037 490 -1031
rect 29 -1082 32 -1076
rect 36 -1082 39 -1076
rect 43 -1082 49 -1076
rect 50 -1082 53 -1076
rect 57 -1082 63 -1076
rect 64 -1082 70 -1076
rect 71 -1082 74 -1076
rect 78 -1082 81 -1076
rect 85 -1082 88 -1076
rect 92 -1082 98 -1076
rect 99 -1082 102 -1076
rect 106 -1082 112 -1076
rect 113 -1082 119 -1076
rect 120 -1082 123 -1076
rect 127 -1082 130 -1076
rect 134 -1082 137 -1076
rect 141 -1082 147 -1076
rect 148 -1082 154 -1076
rect 155 -1082 161 -1076
rect 162 -1082 168 -1076
rect 169 -1082 175 -1076
rect 176 -1082 179 -1076
rect 183 -1082 186 -1076
rect 190 -1082 196 -1076
rect 197 -1082 203 -1076
rect 204 -1082 207 -1076
rect 211 -1082 217 -1076
rect 218 -1082 224 -1076
rect 225 -1082 231 -1076
rect 232 -1082 238 -1076
rect 239 -1082 242 -1076
rect 246 -1082 249 -1076
rect 253 -1082 256 -1076
rect 260 -1082 263 -1076
rect 267 -1082 273 -1076
rect 274 -1082 280 -1076
rect 281 -1082 287 -1076
rect 288 -1082 294 -1076
rect 295 -1082 298 -1076
rect 302 -1082 308 -1076
rect 309 -1082 312 -1076
rect 316 -1082 319 -1076
rect 323 -1082 326 -1076
rect 330 -1082 333 -1076
rect 337 -1082 343 -1076
rect 344 -1082 350 -1076
rect 351 -1082 354 -1076
rect 358 -1082 361 -1076
rect 365 -1082 368 -1076
rect 372 -1082 375 -1076
rect 379 -1082 382 -1076
rect 386 -1082 389 -1076
rect 393 -1082 396 -1076
rect 400 -1082 403 -1076
rect 407 -1082 410 -1076
rect 414 -1082 417 -1076
rect 421 -1082 424 -1076
rect 428 -1082 431 -1076
rect 435 -1082 438 -1076
rect 442 -1082 445 -1076
rect 449 -1082 452 -1076
rect 456 -1082 459 -1076
rect 463 -1082 466 -1076
rect 470 -1082 476 -1076
rect 477 -1082 483 -1076
rect 484 -1082 487 -1076
rect 491 -1082 497 -1076
rect 498 -1082 501 -1076
rect 43 -1115 49 -1109
rect 64 -1115 67 -1109
rect 71 -1115 74 -1109
rect 78 -1115 84 -1109
rect 85 -1115 91 -1109
rect 92 -1115 98 -1109
rect 99 -1115 102 -1109
rect 106 -1115 112 -1109
rect 113 -1115 116 -1109
rect 120 -1115 126 -1109
rect 127 -1115 130 -1109
rect 134 -1115 137 -1109
rect 141 -1115 147 -1109
rect 148 -1115 151 -1109
rect 155 -1115 158 -1109
rect 162 -1115 168 -1109
rect 169 -1115 172 -1109
rect 176 -1115 179 -1109
rect 183 -1115 186 -1109
rect 190 -1115 196 -1109
rect 197 -1115 203 -1109
rect 204 -1115 210 -1109
rect 211 -1115 217 -1109
rect 218 -1115 224 -1109
rect 225 -1115 231 -1109
rect 232 -1115 238 -1109
rect 239 -1115 242 -1109
rect 246 -1115 252 -1109
rect 253 -1115 256 -1109
rect 260 -1115 263 -1109
rect 267 -1115 273 -1109
rect 274 -1115 277 -1109
rect 281 -1115 287 -1109
rect 288 -1115 291 -1109
rect 295 -1115 298 -1109
rect 302 -1115 305 -1109
rect 309 -1115 315 -1109
rect 316 -1115 319 -1109
rect 323 -1115 326 -1109
rect 330 -1115 336 -1109
rect 337 -1115 340 -1109
rect 344 -1115 347 -1109
rect 351 -1115 357 -1109
rect 358 -1115 361 -1109
rect 365 -1115 371 -1109
rect 372 -1115 375 -1109
rect 379 -1115 382 -1109
rect 386 -1115 389 -1109
rect 393 -1115 399 -1109
rect 400 -1115 403 -1109
rect 407 -1115 413 -1109
rect 414 -1115 417 -1109
rect 421 -1115 424 -1109
rect 428 -1115 434 -1109
rect 435 -1115 438 -1109
rect 442 -1115 445 -1109
rect 449 -1115 455 -1109
rect 456 -1115 459 -1109
rect 43 -1148 49 -1142
rect 50 -1148 53 -1142
rect 57 -1148 63 -1142
rect 64 -1148 67 -1142
rect 71 -1148 77 -1142
rect 78 -1148 84 -1142
rect 85 -1148 91 -1142
rect 92 -1148 98 -1142
rect 99 -1148 102 -1142
rect 106 -1148 112 -1142
rect 113 -1148 116 -1142
rect 120 -1148 123 -1142
rect 127 -1148 133 -1142
rect 134 -1148 140 -1142
rect 141 -1148 144 -1142
rect 148 -1148 151 -1142
rect 155 -1148 158 -1142
rect 162 -1148 165 -1142
rect 169 -1148 172 -1142
rect 176 -1148 179 -1142
rect 183 -1148 189 -1142
rect 190 -1148 196 -1142
rect 197 -1148 200 -1142
rect 204 -1148 210 -1142
rect 211 -1148 217 -1142
rect 218 -1148 224 -1142
rect 225 -1148 231 -1142
rect 232 -1148 235 -1142
rect 239 -1148 245 -1142
rect 246 -1148 252 -1142
rect 253 -1148 259 -1142
rect 260 -1148 263 -1142
rect 267 -1148 273 -1142
rect 274 -1148 277 -1142
rect 281 -1148 284 -1142
rect 288 -1148 291 -1142
rect 295 -1148 298 -1142
rect 302 -1148 308 -1142
rect 309 -1148 315 -1142
rect 316 -1148 319 -1142
rect 323 -1148 326 -1142
rect 330 -1148 333 -1142
rect 337 -1148 340 -1142
rect 344 -1148 347 -1142
rect 351 -1148 354 -1142
rect 358 -1148 361 -1142
rect 365 -1148 368 -1142
rect 372 -1148 375 -1142
rect 379 -1148 385 -1142
rect 386 -1148 392 -1142
rect 393 -1148 396 -1142
rect 400 -1148 406 -1142
rect 407 -1148 410 -1142
rect 414 -1148 417 -1142
rect 421 -1148 424 -1142
rect 442 -1148 448 -1142
rect 449 -1148 452 -1142
rect 43 -1185 49 -1179
rect 50 -1185 53 -1179
rect 57 -1185 63 -1179
rect 64 -1185 70 -1179
rect 71 -1185 77 -1179
rect 78 -1185 84 -1179
rect 85 -1185 91 -1179
rect 92 -1185 98 -1179
rect 99 -1185 102 -1179
rect 106 -1185 109 -1179
rect 113 -1185 119 -1179
rect 120 -1185 123 -1179
rect 127 -1185 130 -1179
rect 134 -1185 137 -1179
rect 141 -1185 147 -1179
rect 148 -1185 154 -1179
rect 155 -1185 158 -1179
rect 162 -1185 168 -1179
rect 169 -1185 175 -1179
rect 176 -1185 182 -1179
rect 183 -1185 186 -1179
rect 190 -1185 196 -1179
rect 197 -1185 203 -1179
rect 204 -1185 207 -1179
rect 211 -1185 214 -1179
rect 218 -1185 224 -1179
rect 225 -1185 231 -1179
rect 232 -1185 238 -1179
rect 239 -1185 245 -1179
rect 246 -1185 252 -1179
rect 253 -1185 259 -1179
rect 260 -1185 263 -1179
rect 267 -1185 270 -1179
rect 274 -1185 277 -1179
rect 281 -1185 284 -1179
rect 288 -1185 294 -1179
rect 295 -1185 301 -1179
rect 302 -1185 308 -1179
rect 309 -1185 312 -1179
rect 316 -1185 319 -1179
rect 323 -1185 326 -1179
rect 330 -1185 333 -1179
rect 337 -1185 340 -1179
rect 344 -1185 350 -1179
rect 351 -1185 354 -1179
rect 358 -1185 361 -1179
rect 365 -1185 368 -1179
rect 372 -1185 375 -1179
rect 379 -1185 382 -1179
rect 386 -1185 389 -1179
rect 393 -1185 396 -1179
rect 400 -1185 403 -1179
rect 414 -1185 420 -1179
rect 421 -1185 424 -1179
rect 428 -1185 431 -1179
rect 43 -1212 49 -1206
rect 64 -1212 70 -1206
rect 71 -1212 74 -1206
rect 78 -1212 84 -1206
rect 85 -1212 91 -1206
rect 92 -1212 98 -1206
rect 99 -1212 102 -1206
rect 106 -1212 109 -1206
rect 113 -1212 119 -1206
rect 120 -1212 123 -1206
rect 127 -1212 130 -1206
rect 134 -1212 140 -1206
rect 141 -1212 147 -1206
rect 148 -1212 154 -1206
rect 155 -1212 161 -1206
rect 162 -1212 168 -1206
rect 169 -1212 172 -1206
rect 176 -1212 179 -1206
rect 183 -1212 189 -1206
rect 190 -1212 196 -1206
rect 197 -1212 200 -1206
rect 204 -1212 207 -1206
rect 211 -1212 214 -1206
rect 218 -1212 224 -1206
rect 225 -1212 231 -1206
rect 232 -1212 235 -1206
rect 239 -1212 245 -1206
rect 246 -1212 249 -1206
rect 253 -1212 256 -1206
rect 281 -1212 284 -1206
rect 288 -1212 294 -1206
rect 295 -1212 298 -1206
rect 302 -1212 308 -1206
rect 309 -1212 315 -1206
rect 316 -1212 319 -1206
rect 323 -1212 326 -1206
rect 330 -1212 333 -1206
rect 337 -1212 343 -1206
rect 344 -1212 347 -1206
rect 351 -1212 357 -1206
rect 358 -1212 361 -1206
rect 365 -1212 368 -1206
rect 372 -1212 378 -1206
rect 379 -1212 382 -1206
rect 407 -1212 410 -1206
rect 421 -1212 427 -1206
rect 428 -1212 431 -1206
rect 22 -1235 28 -1229
rect 29 -1235 35 -1229
rect 36 -1235 39 -1229
rect 43 -1235 49 -1229
rect 50 -1235 53 -1229
rect 57 -1235 60 -1229
rect 64 -1235 70 -1229
rect 71 -1235 77 -1229
rect 78 -1235 81 -1229
rect 92 -1235 95 -1229
rect 99 -1235 102 -1229
rect 106 -1235 112 -1229
rect 113 -1235 119 -1229
rect 120 -1235 126 -1229
rect 127 -1235 133 -1229
rect 134 -1235 140 -1229
rect 141 -1235 144 -1229
rect 148 -1235 151 -1229
rect 155 -1235 161 -1229
rect 162 -1235 165 -1229
rect 169 -1235 175 -1229
rect 176 -1235 182 -1229
rect 183 -1235 186 -1229
rect 190 -1235 193 -1229
rect 197 -1235 203 -1229
rect 204 -1235 210 -1229
rect 211 -1235 217 -1229
rect 218 -1235 224 -1229
rect 225 -1235 231 -1229
rect 232 -1235 235 -1229
rect 239 -1235 242 -1229
rect 246 -1235 252 -1229
rect 253 -1235 256 -1229
rect 260 -1235 266 -1229
rect 267 -1235 270 -1229
rect 274 -1235 277 -1229
rect 281 -1235 284 -1229
rect 288 -1235 294 -1229
rect 295 -1235 301 -1229
rect 302 -1235 305 -1229
rect 309 -1235 312 -1229
rect 316 -1235 322 -1229
rect 323 -1235 329 -1229
rect 337 -1235 340 -1229
rect 344 -1235 350 -1229
rect 351 -1235 354 -1229
rect 358 -1235 361 -1229
rect 365 -1235 371 -1229
rect 372 -1235 375 -1229
rect 400 -1235 403 -1229
rect 407 -1235 413 -1229
rect 414 -1235 420 -1229
rect 421 -1235 424 -1229
rect 428 -1235 434 -1229
rect 22 -1260 28 -1254
rect 29 -1260 32 -1254
rect 36 -1260 42 -1254
rect 43 -1260 49 -1254
rect 57 -1260 60 -1254
rect 64 -1260 70 -1254
rect 71 -1260 77 -1254
rect 78 -1260 81 -1254
rect 99 -1260 105 -1254
rect 106 -1260 112 -1254
rect 113 -1260 116 -1254
rect 120 -1260 123 -1254
rect 127 -1260 130 -1254
rect 134 -1260 140 -1254
rect 141 -1260 147 -1254
rect 148 -1260 154 -1254
rect 155 -1260 161 -1254
rect 162 -1260 168 -1254
rect 169 -1260 172 -1254
rect 176 -1260 179 -1254
rect 183 -1260 189 -1254
rect 190 -1260 196 -1254
rect 197 -1260 203 -1254
rect 204 -1260 210 -1254
rect 211 -1260 214 -1254
rect 218 -1260 224 -1254
rect 225 -1260 231 -1254
rect 232 -1260 235 -1254
rect 239 -1260 245 -1254
rect 246 -1260 252 -1254
rect 253 -1260 259 -1254
rect 260 -1260 263 -1254
rect 267 -1260 270 -1254
rect 274 -1260 280 -1254
rect 281 -1260 287 -1254
rect 288 -1260 291 -1254
rect 295 -1260 301 -1254
rect 302 -1260 305 -1254
rect 316 -1260 322 -1254
rect 323 -1260 326 -1254
rect 330 -1260 336 -1254
rect 337 -1260 340 -1254
rect 344 -1260 350 -1254
rect 351 -1260 357 -1254
rect 358 -1260 361 -1254
rect 365 -1260 371 -1254
<< polysilicon >>
rect 138 -5 139 -3
rect 142 -11 143 -9
rect 145 -11 146 -9
rect 149 -5 150 -3
rect 149 -11 150 -9
rect 177 -5 178 -3
rect 177 -11 178 -9
rect 187 -5 188 -3
rect 184 -11 185 -9
rect 187 -11 188 -9
rect 191 -5 192 -3
rect 198 -5 199 -3
rect 198 -11 199 -9
rect 205 -5 206 -3
rect 208 -11 209 -9
rect 212 -5 213 -3
rect 215 -5 216 -3
rect 219 -5 220 -3
rect 219 -11 220 -9
rect 226 -5 227 -3
rect 229 -11 230 -9
rect 236 -11 237 -9
rect 240 -5 241 -3
rect 240 -11 241 -9
rect 128 -30 129 -28
rect 135 -24 136 -22
rect 135 -30 136 -28
rect 142 -24 143 -22
rect 142 -30 143 -28
rect 152 -30 153 -28
rect 156 -24 157 -22
rect 159 -30 160 -28
rect 163 -24 164 -22
rect 163 -30 164 -28
rect 170 -24 171 -22
rect 177 -24 178 -22
rect 177 -30 178 -28
rect 184 -24 185 -22
rect 191 -24 192 -22
rect 198 -24 199 -22
rect 198 -30 199 -28
rect 205 -24 206 -22
rect 205 -30 206 -28
rect 215 -24 216 -22
rect 219 -24 220 -22
rect 226 -24 227 -22
rect 229 -24 230 -22
rect 226 -30 227 -28
rect 229 -30 230 -28
rect 233 -24 234 -22
rect 233 -30 234 -28
rect 240 -24 241 -22
rect 240 -30 241 -28
rect 247 -24 248 -22
rect 254 -24 255 -22
rect 296 -30 297 -28
rect 324 -24 325 -22
rect 327 -30 328 -28
rect 331 -24 332 -22
rect 331 -30 332 -28
rect 135 -51 136 -49
rect 135 -57 136 -55
rect 145 -51 146 -49
rect 142 -57 143 -55
rect 152 -51 153 -49
rect 159 -51 160 -49
rect 163 -51 164 -49
rect 173 -51 174 -49
rect 170 -57 171 -55
rect 177 -51 178 -49
rect 184 -51 185 -49
rect 184 -57 185 -55
rect 191 -51 192 -49
rect 191 -57 192 -55
rect 198 -51 199 -49
rect 201 -51 202 -49
rect 205 -51 206 -49
rect 208 -51 209 -49
rect 212 -51 213 -49
rect 212 -57 213 -55
rect 219 -51 220 -49
rect 222 -51 223 -49
rect 219 -57 220 -55
rect 226 -51 227 -49
rect 229 -51 230 -49
rect 229 -57 230 -55
rect 233 -51 234 -49
rect 233 -57 234 -55
rect 240 -51 241 -49
rect 240 -57 241 -55
rect 247 -51 248 -49
rect 247 -57 248 -55
rect 254 -57 255 -55
rect 261 -51 262 -49
rect 261 -57 262 -55
rect 268 -51 269 -49
rect 268 -57 269 -55
rect 278 -57 279 -55
rect 282 -51 283 -49
rect 282 -57 283 -55
rect 289 -51 290 -49
rect 289 -57 290 -55
rect 296 -57 297 -55
rect 299 -57 300 -55
rect 303 -51 304 -49
rect 303 -57 304 -55
rect 324 -51 325 -49
rect 324 -57 325 -55
rect 331 -51 332 -49
rect 331 -57 332 -55
rect 89 -80 90 -78
rect 103 -74 104 -72
rect 107 -74 108 -72
rect 107 -80 108 -78
rect 117 -80 118 -78
rect 121 -74 122 -72
rect 121 -80 122 -78
rect 128 -74 129 -72
rect 128 -80 129 -78
rect 138 -80 139 -78
rect 142 -74 143 -72
rect 142 -80 143 -78
rect 145 -80 146 -78
rect 149 -74 150 -72
rect 149 -80 150 -78
rect 159 -74 160 -72
rect 163 -74 164 -72
rect 166 -74 167 -72
rect 170 -74 171 -72
rect 170 -80 171 -78
rect 177 -74 178 -72
rect 177 -80 178 -78
rect 184 -74 185 -72
rect 191 -74 192 -72
rect 191 -80 192 -78
rect 201 -74 202 -72
rect 198 -80 199 -78
rect 205 -74 206 -72
rect 205 -80 206 -78
rect 215 -80 216 -78
rect 219 -74 220 -72
rect 222 -80 223 -78
rect 226 -74 227 -72
rect 229 -80 230 -78
rect 236 -80 237 -78
rect 240 -74 241 -72
rect 240 -80 241 -78
rect 247 -80 248 -78
rect 254 -74 255 -72
rect 254 -80 255 -78
rect 261 -74 262 -72
rect 261 -80 262 -78
rect 271 -80 272 -78
rect 275 -74 276 -72
rect 275 -80 276 -78
rect 282 -74 283 -72
rect 282 -80 283 -78
rect 292 -74 293 -72
rect 292 -80 293 -78
rect 296 -74 297 -72
rect 296 -80 297 -78
rect 306 -74 307 -72
rect 313 -74 314 -72
rect 317 -80 318 -78
rect 320 -80 321 -78
rect 324 -74 325 -72
rect 324 -80 325 -78
rect 331 -74 332 -72
rect 331 -80 332 -78
rect 89 -99 90 -97
rect 100 -99 101 -97
rect 103 -105 104 -103
rect 107 -99 108 -97
rect 107 -105 108 -103
rect 114 -99 115 -97
rect 114 -105 115 -103
rect 121 -99 122 -97
rect 124 -105 125 -103
rect 128 -99 129 -97
rect 131 -99 132 -97
rect 128 -105 129 -103
rect 135 -99 136 -97
rect 135 -105 136 -103
rect 145 -99 146 -97
rect 149 -99 150 -97
rect 149 -105 150 -103
rect 159 -99 160 -97
rect 163 -99 164 -97
rect 166 -99 167 -97
rect 163 -105 164 -103
rect 170 -105 171 -103
rect 177 -105 178 -103
rect 180 -105 181 -103
rect 184 -99 185 -97
rect 184 -105 185 -103
rect 194 -99 195 -97
rect 198 -99 199 -97
rect 198 -105 199 -103
rect 205 -105 206 -103
rect 208 -105 209 -103
rect 212 -99 213 -97
rect 212 -105 213 -103
rect 215 -105 216 -103
rect 219 -99 220 -97
rect 222 -99 223 -97
rect 219 -105 220 -103
rect 226 -99 227 -97
rect 229 -99 230 -97
rect 229 -105 230 -103
rect 233 -99 234 -97
rect 233 -105 234 -103
rect 240 -105 241 -103
rect 243 -105 244 -103
rect 247 -99 248 -97
rect 247 -105 248 -103
rect 254 -99 255 -97
rect 254 -105 255 -103
rect 261 -99 262 -97
rect 261 -105 262 -103
rect 268 -105 269 -103
rect 271 -105 272 -103
rect 275 -99 276 -97
rect 275 -105 276 -103
rect 282 -105 283 -103
rect 289 -105 290 -103
rect 296 -99 297 -97
rect 296 -105 297 -103
rect 303 -99 304 -97
rect 303 -105 304 -103
rect 310 -99 311 -97
rect 310 -105 311 -103
rect 317 -99 318 -97
rect 317 -105 318 -103
rect 324 -99 325 -97
rect 324 -105 325 -103
rect 383 -105 384 -103
rect 79 -130 80 -128
rect 86 -124 87 -122
rect 86 -130 87 -128
rect 103 -124 104 -122
rect 107 -124 108 -122
rect 107 -130 108 -128
rect 114 -124 115 -122
rect 117 -130 118 -128
rect 124 -124 125 -122
rect 121 -130 122 -128
rect 128 -130 129 -128
rect 131 -130 132 -128
rect 135 -124 136 -122
rect 135 -130 136 -128
rect 145 -124 146 -122
rect 152 -130 153 -128
rect 156 -124 157 -122
rect 156 -130 157 -128
rect 163 -124 164 -122
rect 163 -130 164 -128
rect 173 -130 174 -128
rect 180 -124 181 -122
rect 177 -130 178 -128
rect 184 -124 185 -122
rect 184 -130 185 -128
rect 191 -124 192 -122
rect 194 -130 195 -128
rect 198 -124 199 -122
rect 198 -130 199 -128
rect 205 -124 206 -122
rect 205 -130 206 -128
rect 212 -124 213 -122
rect 215 -124 216 -122
rect 215 -130 216 -128
rect 219 -124 220 -122
rect 219 -130 220 -128
rect 226 -124 227 -122
rect 229 -130 230 -128
rect 236 -124 237 -122
rect 240 -124 241 -122
rect 240 -130 241 -128
rect 254 -124 255 -122
rect 254 -130 255 -128
rect 261 -124 262 -122
rect 261 -130 262 -128
rect 268 -124 269 -122
rect 268 -130 269 -128
rect 299 -124 300 -122
rect 296 -130 297 -128
rect 299 -130 300 -128
rect 303 -124 304 -122
rect 303 -130 304 -128
rect 310 -124 311 -122
rect 317 -124 318 -122
rect 317 -130 318 -128
rect 380 -124 381 -122
rect 380 -130 381 -128
rect 79 -149 80 -147
rect 82 -149 83 -147
rect 82 -155 83 -153
rect 107 -149 108 -147
rect 107 -155 108 -153
rect 114 -149 115 -147
rect 114 -155 115 -153
rect 121 -149 122 -147
rect 121 -155 122 -153
rect 128 -149 129 -147
rect 131 -149 132 -147
rect 138 -149 139 -147
rect 135 -155 136 -153
rect 138 -155 139 -153
rect 142 -149 143 -147
rect 145 -149 146 -147
rect 152 -149 153 -147
rect 152 -155 153 -153
rect 156 -149 157 -147
rect 159 -149 160 -147
rect 163 -149 164 -147
rect 163 -155 164 -153
rect 170 -149 171 -147
rect 173 -149 174 -147
rect 173 -155 174 -153
rect 177 -149 178 -147
rect 177 -155 178 -153
rect 184 -155 185 -153
rect 187 -155 188 -153
rect 191 -149 192 -147
rect 191 -155 192 -153
rect 198 -149 199 -147
rect 201 -155 202 -153
rect 205 -149 206 -147
rect 208 -149 209 -147
rect 205 -155 206 -153
rect 215 -149 216 -147
rect 212 -155 213 -153
rect 215 -155 216 -153
rect 219 -149 220 -147
rect 219 -155 220 -153
rect 226 -149 227 -147
rect 226 -155 227 -153
rect 233 -149 234 -147
rect 233 -155 234 -153
rect 243 -155 244 -153
rect 254 -149 255 -147
rect 257 -149 258 -147
rect 254 -155 255 -153
rect 261 -149 262 -147
rect 261 -155 262 -153
rect 268 -149 269 -147
rect 271 -149 272 -147
rect 268 -155 269 -153
rect 271 -155 272 -153
rect 275 -149 276 -147
rect 275 -155 276 -153
rect 310 -149 311 -147
rect 313 -155 314 -153
rect 317 -149 318 -147
rect 317 -155 318 -153
rect 320 -155 321 -153
rect 324 -149 325 -147
rect 324 -155 325 -153
rect 383 -155 384 -153
rect 387 -149 388 -147
rect 387 -155 388 -153
rect 82 -172 83 -170
rect 117 -172 118 -170
rect 124 -172 125 -170
rect 121 -178 122 -176
rect 131 -178 132 -176
rect 135 -172 136 -170
rect 135 -178 136 -176
rect 145 -172 146 -170
rect 152 -172 153 -170
rect 156 -172 157 -170
rect 159 -178 160 -176
rect 163 -172 164 -170
rect 163 -178 164 -176
rect 170 -172 171 -170
rect 170 -178 171 -176
rect 177 -172 178 -170
rect 177 -178 178 -176
rect 184 -178 185 -176
rect 191 -172 192 -170
rect 198 -172 199 -170
rect 198 -178 199 -176
rect 205 -172 206 -170
rect 205 -178 206 -176
rect 212 -172 213 -170
rect 215 -172 216 -170
rect 219 -172 220 -170
rect 219 -178 220 -176
rect 226 -172 227 -170
rect 229 -172 230 -170
rect 229 -178 230 -176
rect 233 -172 234 -170
rect 233 -178 234 -176
rect 240 -172 241 -170
rect 240 -178 241 -176
rect 247 -172 248 -170
rect 247 -178 248 -176
rect 254 -172 255 -170
rect 254 -178 255 -176
rect 261 -172 262 -170
rect 261 -178 262 -176
rect 271 -178 272 -176
rect 278 -172 279 -170
rect 275 -178 276 -176
rect 282 -172 283 -170
rect 285 -178 286 -176
rect 289 -172 290 -170
rect 289 -178 290 -176
rect 296 -172 297 -170
rect 296 -178 297 -176
rect 303 -172 304 -170
rect 303 -178 304 -176
rect 313 -178 314 -176
rect 317 -172 318 -170
rect 317 -178 318 -176
rect 324 -172 325 -170
rect 324 -178 325 -176
rect 331 -172 332 -170
rect 331 -178 332 -176
rect 341 -172 342 -170
rect 345 -172 346 -170
rect 345 -178 346 -176
rect 352 -172 353 -170
rect 355 -178 356 -176
rect 359 -172 360 -170
rect 362 -172 363 -170
rect 366 -172 367 -170
rect 366 -178 367 -176
rect 373 -172 374 -170
rect 373 -178 374 -176
rect 380 -172 381 -170
rect 383 -172 384 -170
rect 387 -172 388 -170
rect 387 -178 388 -176
rect 394 -172 395 -170
rect 394 -178 395 -176
rect 408 -172 409 -170
rect 408 -178 409 -176
rect 415 -172 416 -170
rect 415 -178 416 -176
rect 436 -172 437 -170
rect 443 -172 444 -170
rect 443 -178 444 -176
rect 75 -199 76 -197
rect 79 -199 80 -197
rect 79 -205 80 -203
rect 86 -199 87 -197
rect 89 -199 90 -197
rect 86 -205 87 -203
rect 93 -199 94 -197
rect 96 -205 97 -203
rect 103 -205 104 -203
rect 107 -199 108 -197
rect 107 -205 108 -203
rect 114 -205 115 -203
rect 121 -199 122 -197
rect 121 -205 122 -203
rect 128 -199 129 -197
rect 131 -199 132 -197
rect 131 -205 132 -203
rect 135 -199 136 -197
rect 142 -199 143 -197
rect 145 -205 146 -203
rect 149 -199 150 -197
rect 149 -205 150 -203
rect 156 -199 157 -197
rect 156 -205 157 -203
rect 163 -199 164 -197
rect 163 -205 164 -203
rect 170 -199 171 -197
rect 170 -205 171 -203
rect 177 -199 178 -197
rect 177 -205 178 -203
rect 184 -199 185 -197
rect 184 -205 185 -203
rect 191 -199 192 -197
rect 191 -205 192 -203
rect 201 -199 202 -197
rect 205 -199 206 -197
rect 205 -205 206 -203
rect 212 -199 213 -197
rect 215 -199 216 -197
rect 212 -205 213 -203
rect 219 -199 220 -197
rect 219 -205 220 -203
rect 229 -199 230 -197
rect 229 -205 230 -203
rect 233 -199 234 -197
rect 233 -205 234 -203
rect 240 -199 241 -197
rect 240 -205 241 -203
rect 250 -199 251 -197
rect 247 -205 248 -203
rect 254 -199 255 -197
rect 254 -205 255 -203
rect 261 -199 262 -197
rect 264 -205 265 -203
rect 268 -199 269 -197
rect 268 -205 269 -203
rect 275 -199 276 -197
rect 275 -205 276 -203
rect 282 -199 283 -197
rect 285 -199 286 -197
rect 289 -199 290 -197
rect 289 -205 290 -203
rect 296 -199 297 -197
rect 296 -205 297 -203
rect 303 -199 304 -197
rect 306 -205 307 -203
rect 310 -199 311 -197
rect 310 -205 311 -203
rect 317 -199 318 -197
rect 317 -205 318 -203
rect 324 -199 325 -197
rect 324 -205 325 -203
rect 331 -199 332 -197
rect 331 -205 332 -203
rect 338 -199 339 -197
rect 338 -205 339 -203
rect 345 -199 346 -197
rect 345 -205 346 -203
rect 352 -199 353 -197
rect 352 -205 353 -203
rect 359 -199 360 -197
rect 359 -205 360 -203
rect 369 -199 370 -197
rect 369 -205 370 -203
rect 373 -199 374 -197
rect 373 -205 374 -203
rect 380 -199 381 -197
rect 383 -199 384 -197
rect 380 -205 381 -203
rect 383 -205 384 -203
rect 394 -199 395 -197
rect 394 -205 395 -203
rect 401 -199 402 -197
rect 401 -205 402 -203
rect 404 -205 405 -203
rect 408 -199 409 -197
rect 408 -205 409 -203
rect 415 -199 416 -197
rect 415 -205 416 -203
rect 422 -199 423 -197
rect 432 -199 433 -197
rect 436 -199 437 -197
rect 436 -205 437 -203
rect 443 -199 444 -197
rect 68 -238 69 -236
rect 72 -232 73 -230
rect 79 -232 80 -230
rect 79 -238 80 -236
rect 86 -232 87 -230
rect 86 -238 87 -236
rect 93 -232 94 -230
rect 93 -238 94 -236
rect 100 -232 101 -230
rect 100 -238 101 -236
rect 107 -232 108 -230
rect 107 -238 108 -236
rect 114 -232 115 -230
rect 114 -238 115 -236
rect 121 -232 122 -230
rect 121 -238 122 -236
rect 128 -232 129 -230
rect 128 -238 129 -236
rect 135 -238 136 -236
rect 138 -238 139 -236
rect 142 -232 143 -230
rect 142 -238 143 -236
rect 149 -232 150 -230
rect 149 -238 150 -236
rect 152 -238 153 -236
rect 159 -232 160 -230
rect 156 -238 157 -236
rect 159 -238 160 -236
rect 166 -238 167 -236
rect 170 -232 171 -230
rect 170 -238 171 -236
rect 177 -232 178 -230
rect 180 -232 181 -230
rect 180 -238 181 -236
rect 187 -232 188 -230
rect 187 -238 188 -236
rect 191 -232 192 -230
rect 191 -238 192 -236
rect 198 -232 199 -230
rect 201 -232 202 -230
rect 205 -232 206 -230
rect 205 -238 206 -236
rect 212 -232 213 -230
rect 212 -238 213 -236
rect 219 -232 220 -230
rect 222 -232 223 -230
rect 219 -238 220 -236
rect 226 -232 227 -230
rect 229 -232 230 -230
rect 226 -238 227 -236
rect 233 -232 234 -230
rect 236 -232 237 -230
rect 240 -232 241 -230
rect 240 -238 241 -236
rect 243 -238 244 -236
rect 247 -232 248 -230
rect 250 -238 251 -236
rect 257 -232 258 -230
rect 254 -238 255 -236
rect 261 -232 262 -230
rect 261 -238 262 -236
rect 264 -238 265 -236
rect 268 -232 269 -230
rect 268 -238 269 -236
rect 275 -232 276 -230
rect 275 -238 276 -236
rect 282 -232 283 -230
rect 282 -238 283 -236
rect 289 -232 290 -230
rect 289 -238 290 -236
rect 296 -232 297 -230
rect 296 -238 297 -236
rect 303 -232 304 -230
rect 303 -238 304 -236
rect 310 -232 311 -230
rect 310 -238 311 -236
rect 317 -232 318 -230
rect 317 -238 318 -236
rect 324 -232 325 -230
rect 331 -232 332 -230
rect 331 -238 332 -236
rect 338 -232 339 -230
rect 338 -238 339 -236
rect 345 -232 346 -230
rect 345 -238 346 -236
rect 352 -232 353 -230
rect 352 -238 353 -236
rect 359 -232 360 -230
rect 359 -238 360 -236
rect 366 -238 367 -236
rect 369 -238 370 -236
rect 373 -232 374 -230
rect 373 -238 374 -236
rect 380 -232 381 -230
rect 387 -232 388 -230
rect 387 -238 388 -236
rect 418 -238 419 -236
rect 422 -232 423 -230
rect 422 -238 423 -236
rect 439 -232 440 -230
rect 30 -281 31 -279
rect 33 -281 34 -279
rect 37 -281 38 -279
rect 54 -281 55 -279
rect 72 -275 73 -273
rect 79 -275 80 -273
rect 79 -281 80 -279
rect 86 -275 87 -273
rect 93 -275 94 -273
rect 93 -281 94 -279
rect 103 -281 104 -279
rect 107 -275 108 -273
rect 107 -281 108 -279
rect 114 -275 115 -273
rect 114 -281 115 -279
rect 121 -275 122 -273
rect 121 -281 122 -279
rect 131 -275 132 -273
rect 131 -281 132 -279
rect 135 -275 136 -273
rect 145 -275 146 -273
rect 149 -275 150 -273
rect 152 -275 153 -273
rect 149 -281 150 -279
rect 152 -281 153 -279
rect 156 -275 157 -273
rect 156 -281 157 -279
rect 163 -275 164 -273
rect 163 -281 164 -279
rect 170 -275 171 -273
rect 170 -281 171 -279
rect 177 -275 178 -273
rect 177 -281 178 -279
rect 184 -275 185 -273
rect 187 -275 188 -273
rect 184 -281 185 -279
rect 187 -281 188 -279
rect 194 -275 195 -273
rect 194 -281 195 -279
rect 198 -275 199 -273
rect 198 -281 199 -279
rect 205 -275 206 -273
rect 208 -275 209 -273
rect 212 -275 213 -273
rect 215 -275 216 -273
rect 219 -281 220 -279
rect 222 -281 223 -279
rect 226 -275 227 -273
rect 229 -275 230 -273
rect 226 -281 227 -279
rect 233 -275 234 -273
rect 233 -281 234 -279
rect 240 -275 241 -273
rect 240 -281 241 -279
rect 247 -275 248 -273
rect 247 -281 248 -279
rect 254 -275 255 -273
rect 257 -275 258 -273
rect 254 -281 255 -279
rect 261 -275 262 -273
rect 261 -281 262 -279
rect 268 -275 269 -273
rect 271 -275 272 -273
rect 268 -281 269 -279
rect 275 -275 276 -273
rect 275 -281 276 -279
rect 282 -275 283 -273
rect 282 -281 283 -279
rect 292 -275 293 -273
rect 292 -281 293 -279
rect 296 -275 297 -273
rect 299 -275 300 -273
rect 296 -281 297 -279
rect 303 -275 304 -273
rect 306 -281 307 -279
rect 310 -275 311 -273
rect 310 -281 311 -279
rect 317 -275 318 -273
rect 317 -281 318 -279
rect 324 -275 325 -273
rect 324 -281 325 -279
rect 331 -275 332 -273
rect 331 -281 332 -279
rect 338 -275 339 -273
rect 338 -281 339 -279
rect 345 -275 346 -273
rect 345 -281 346 -279
rect 352 -275 353 -273
rect 352 -281 353 -279
rect 359 -275 360 -273
rect 359 -281 360 -279
rect 366 -275 367 -273
rect 366 -281 367 -279
rect 373 -275 374 -273
rect 373 -281 374 -279
rect 380 -275 381 -273
rect 380 -281 381 -279
rect 387 -275 388 -273
rect 387 -281 388 -279
rect 394 -275 395 -273
rect 394 -281 395 -279
rect 401 -275 402 -273
rect 401 -281 402 -279
rect 408 -275 409 -273
rect 408 -281 409 -279
rect 415 -275 416 -273
rect 418 -275 419 -273
rect 415 -281 416 -279
rect 422 -275 423 -273
rect 422 -281 423 -279
rect 429 -275 430 -273
rect 429 -281 430 -279
rect 439 -275 440 -273
rect 443 -275 444 -273
rect 443 -281 444 -279
rect 450 -275 451 -273
rect 453 -275 454 -273
rect 450 -281 451 -279
rect 457 -275 458 -273
rect 457 -281 458 -279
rect 530 -275 531 -273
rect 534 -275 535 -273
rect 534 -281 535 -279
rect 30 -316 31 -314
rect 47 -316 48 -314
rect 51 -316 52 -314
rect 58 -316 59 -314
rect 58 -322 59 -320
rect 68 -316 69 -314
rect 75 -316 76 -314
rect 82 -316 83 -314
rect 82 -322 83 -320
rect 86 -316 87 -314
rect 86 -322 87 -320
rect 93 -316 94 -314
rect 93 -322 94 -320
rect 100 -316 101 -314
rect 100 -322 101 -320
rect 107 -322 108 -320
rect 110 -322 111 -320
rect 114 -316 115 -314
rect 114 -322 115 -320
rect 121 -316 122 -314
rect 121 -322 122 -320
rect 128 -316 129 -314
rect 128 -322 129 -320
rect 135 -316 136 -314
rect 135 -322 136 -320
rect 142 -316 143 -314
rect 145 -316 146 -314
rect 142 -322 143 -320
rect 149 -316 150 -314
rect 149 -322 150 -320
rect 152 -322 153 -320
rect 159 -322 160 -320
rect 163 -316 164 -314
rect 163 -322 164 -320
rect 170 -316 171 -314
rect 170 -322 171 -320
rect 177 -316 178 -314
rect 177 -322 178 -320
rect 184 -316 185 -314
rect 184 -322 185 -320
rect 191 -316 192 -314
rect 194 -322 195 -320
rect 198 -316 199 -314
rect 198 -322 199 -320
rect 205 -316 206 -314
rect 208 -316 209 -314
rect 212 -316 213 -314
rect 212 -322 213 -320
rect 219 -316 220 -314
rect 219 -322 220 -320
rect 226 -316 227 -314
rect 229 -316 230 -314
rect 229 -322 230 -320
rect 233 -316 234 -314
rect 233 -322 234 -320
rect 243 -316 244 -314
rect 240 -322 241 -320
rect 243 -322 244 -320
rect 247 -316 248 -314
rect 247 -322 248 -320
rect 250 -322 251 -320
rect 254 -322 255 -320
rect 261 -316 262 -314
rect 264 -322 265 -320
rect 268 -316 269 -314
rect 268 -322 269 -320
rect 275 -316 276 -314
rect 275 -322 276 -320
rect 282 -316 283 -314
rect 282 -322 283 -320
rect 285 -322 286 -320
rect 289 -316 290 -314
rect 289 -322 290 -320
rect 296 -316 297 -314
rect 299 -316 300 -314
rect 299 -322 300 -320
rect 303 -316 304 -314
rect 303 -322 304 -320
rect 310 -316 311 -314
rect 310 -322 311 -320
rect 317 -316 318 -314
rect 317 -322 318 -320
rect 324 -322 325 -320
rect 331 -316 332 -314
rect 331 -322 332 -320
rect 338 -316 339 -314
rect 338 -322 339 -320
rect 345 -316 346 -314
rect 345 -322 346 -320
rect 352 -316 353 -314
rect 352 -322 353 -320
rect 359 -316 360 -314
rect 359 -322 360 -320
rect 366 -316 367 -314
rect 366 -322 367 -320
rect 376 -316 377 -314
rect 373 -322 374 -320
rect 380 -316 381 -314
rect 380 -322 381 -320
rect 387 -316 388 -314
rect 387 -322 388 -320
rect 394 -316 395 -314
rect 394 -322 395 -320
rect 401 -316 402 -314
rect 401 -322 402 -320
rect 408 -316 409 -314
rect 408 -322 409 -320
rect 418 -316 419 -314
rect 422 -316 423 -314
rect 422 -322 423 -320
rect 429 -322 430 -320
rect 436 -316 437 -314
rect 436 -322 437 -320
rect 453 -316 454 -314
rect 520 -322 521 -320
rect 523 -322 524 -320
rect 527 -316 528 -314
rect 527 -322 528 -320
rect 19 -363 20 -361
rect 16 -369 17 -367
rect 23 -363 24 -361
rect 30 -369 31 -367
rect 37 -363 38 -361
rect 37 -369 38 -367
rect 44 -363 45 -361
rect 44 -369 45 -367
rect 51 -363 52 -361
rect 51 -369 52 -367
rect 58 -363 59 -361
rect 58 -369 59 -367
rect 65 -363 66 -361
rect 65 -369 66 -367
rect 72 -363 73 -361
rect 72 -369 73 -367
rect 82 -363 83 -361
rect 82 -369 83 -367
rect 86 -363 87 -361
rect 89 -369 90 -367
rect 96 -363 97 -361
rect 93 -369 94 -367
rect 100 -363 101 -361
rect 100 -369 101 -367
rect 107 -363 108 -361
rect 110 -363 111 -361
rect 107 -369 108 -367
rect 110 -369 111 -367
rect 114 -363 115 -361
rect 117 -363 118 -361
rect 114 -369 115 -367
rect 117 -369 118 -367
rect 124 -363 125 -361
rect 124 -369 125 -367
rect 131 -363 132 -361
rect 131 -369 132 -367
rect 135 -363 136 -361
rect 138 -363 139 -361
rect 135 -369 136 -367
rect 145 -363 146 -361
rect 142 -369 143 -367
rect 149 -363 150 -361
rect 149 -369 150 -367
rect 156 -363 157 -361
rect 156 -369 157 -367
rect 166 -363 167 -361
rect 166 -369 167 -367
rect 170 -363 171 -361
rect 173 -369 174 -367
rect 177 -363 178 -361
rect 177 -369 178 -367
rect 184 -363 185 -361
rect 184 -369 185 -367
rect 194 -363 195 -361
rect 191 -369 192 -367
rect 198 -363 199 -361
rect 201 -363 202 -361
rect 205 -363 206 -361
rect 205 -369 206 -367
rect 212 -363 213 -361
rect 215 -363 216 -361
rect 212 -369 213 -367
rect 219 -363 220 -361
rect 219 -369 220 -367
rect 226 -363 227 -361
rect 226 -369 227 -367
rect 233 -363 234 -361
rect 233 -369 234 -367
rect 240 -363 241 -361
rect 243 -363 244 -361
rect 240 -369 241 -367
rect 243 -369 244 -367
rect 250 -363 251 -361
rect 247 -369 248 -367
rect 250 -369 251 -367
rect 254 -369 255 -367
rect 261 -363 262 -361
rect 264 -363 265 -361
rect 261 -369 262 -367
rect 271 -363 272 -361
rect 268 -369 269 -367
rect 271 -369 272 -367
rect 275 -369 276 -367
rect 278 -369 279 -367
rect 285 -363 286 -361
rect 282 -369 283 -367
rect 289 -363 290 -361
rect 289 -369 290 -367
rect 296 -363 297 -361
rect 296 -369 297 -367
rect 306 -363 307 -361
rect 310 -363 311 -361
rect 310 -369 311 -367
rect 317 -369 318 -367
rect 320 -369 321 -367
rect 324 -363 325 -361
rect 327 -363 328 -361
rect 324 -369 325 -367
rect 331 -363 332 -361
rect 331 -369 332 -367
rect 338 -363 339 -361
rect 338 -369 339 -367
rect 345 -363 346 -361
rect 345 -369 346 -367
rect 352 -363 353 -361
rect 352 -369 353 -367
rect 359 -363 360 -361
rect 359 -369 360 -367
rect 366 -363 367 -361
rect 366 -369 367 -367
rect 373 -363 374 -361
rect 373 -369 374 -367
rect 380 -363 381 -361
rect 380 -369 381 -367
rect 390 -363 391 -361
rect 387 -369 388 -367
rect 390 -369 391 -367
rect 394 -363 395 -361
rect 394 -369 395 -367
rect 401 -363 402 -361
rect 401 -369 402 -367
rect 408 -363 409 -361
rect 408 -369 409 -367
rect 415 -363 416 -361
rect 415 -369 416 -367
rect 422 -363 423 -361
rect 422 -369 423 -367
rect 429 -363 430 -361
rect 429 -369 430 -367
rect 436 -363 437 -361
rect 436 -369 437 -367
rect 443 -363 444 -361
rect 443 -369 444 -367
rect 450 -363 451 -361
rect 450 -369 451 -367
rect 457 -363 458 -361
rect 457 -369 458 -367
rect 467 -363 468 -361
rect 471 -363 472 -361
rect 471 -369 472 -367
rect 513 -363 514 -361
rect 513 -369 514 -367
rect 16 -414 17 -412
rect 23 -414 24 -412
rect 23 -420 24 -418
rect 30 -414 31 -412
rect 30 -420 31 -418
rect 37 -414 38 -412
rect 44 -414 45 -412
rect 51 -420 52 -418
rect 58 -414 59 -412
rect 65 -414 66 -412
rect 72 -414 73 -412
rect 72 -420 73 -418
rect 79 -414 80 -412
rect 79 -420 80 -418
rect 86 -414 87 -412
rect 86 -420 87 -418
rect 93 -414 94 -412
rect 93 -420 94 -418
rect 100 -414 101 -412
rect 103 -414 104 -412
rect 107 -414 108 -412
rect 110 -414 111 -412
rect 110 -420 111 -418
rect 114 -414 115 -412
rect 114 -420 115 -418
rect 121 -414 122 -412
rect 121 -420 122 -418
rect 128 -414 129 -412
rect 128 -420 129 -418
rect 138 -414 139 -412
rect 142 -420 143 -418
rect 145 -420 146 -418
rect 152 -414 153 -412
rect 156 -414 157 -412
rect 159 -414 160 -412
rect 166 -414 167 -412
rect 170 -414 171 -412
rect 170 -420 171 -418
rect 177 -414 178 -412
rect 177 -420 178 -418
rect 184 -414 185 -412
rect 191 -414 192 -412
rect 194 -414 195 -412
rect 198 -414 199 -412
rect 198 -420 199 -418
rect 208 -414 209 -412
rect 212 -414 213 -412
rect 215 -414 216 -412
rect 215 -420 216 -418
rect 219 -414 220 -412
rect 219 -420 220 -418
rect 226 -414 227 -412
rect 229 -414 230 -412
rect 226 -420 227 -418
rect 229 -420 230 -418
rect 233 -414 234 -412
rect 233 -420 234 -418
rect 240 -414 241 -412
rect 240 -420 241 -418
rect 247 -414 248 -412
rect 247 -420 248 -418
rect 254 -414 255 -412
rect 254 -420 255 -418
rect 261 -414 262 -412
rect 261 -420 262 -418
rect 264 -420 265 -418
rect 268 -414 269 -412
rect 275 -414 276 -412
rect 275 -420 276 -418
rect 282 -414 283 -412
rect 285 -420 286 -418
rect 289 -414 290 -412
rect 289 -420 290 -418
rect 296 -414 297 -412
rect 296 -420 297 -418
rect 303 -414 304 -412
rect 303 -420 304 -418
rect 310 -414 311 -412
rect 313 -414 314 -412
rect 317 -414 318 -412
rect 320 -420 321 -418
rect 324 -414 325 -412
rect 327 -414 328 -412
rect 324 -420 325 -418
rect 327 -420 328 -418
rect 331 -414 332 -412
rect 331 -420 332 -418
rect 341 -420 342 -418
rect 348 -414 349 -412
rect 352 -414 353 -412
rect 352 -420 353 -418
rect 359 -414 360 -412
rect 359 -420 360 -418
rect 366 -414 367 -412
rect 366 -420 367 -418
rect 373 -414 374 -412
rect 373 -420 374 -418
rect 380 -414 381 -412
rect 380 -420 381 -418
rect 387 -414 388 -412
rect 387 -420 388 -418
rect 394 -414 395 -412
rect 394 -420 395 -418
rect 397 -420 398 -418
rect 401 -414 402 -412
rect 401 -420 402 -418
rect 408 -414 409 -412
rect 408 -420 409 -418
rect 415 -414 416 -412
rect 418 -414 419 -412
rect 415 -420 416 -418
rect 422 -414 423 -412
rect 422 -420 423 -418
rect 429 -414 430 -412
rect 429 -420 430 -418
rect 436 -414 437 -412
rect 436 -420 437 -418
rect 443 -414 444 -412
rect 443 -420 444 -418
rect 450 -414 451 -412
rect 450 -420 451 -418
rect 457 -414 458 -412
rect 457 -420 458 -418
rect 464 -414 465 -412
rect 464 -420 465 -418
rect 471 -414 472 -412
rect 471 -420 472 -418
rect 481 -414 482 -412
rect 485 -420 486 -418
rect 492 -414 493 -412
rect 492 -420 493 -418
rect 499 -414 500 -412
rect 499 -420 500 -418
rect 506 -414 507 -412
rect 506 -420 507 -418
rect 513 -414 514 -412
rect 513 -420 514 -418
rect 520 -414 521 -412
rect 520 -420 521 -418
rect 527 -414 528 -412
rect 527 -420 528 -418
rect 2 -465 3 -463
rect 2 -471 3 -469
rect 9 -465 10 -463
rect 9 -471 10 -469
rect 16 -465 17 -463
rect 16 -471 17 -469
rect 23 -471 24 -469
rect 30 -465 31 -463
rect 37 -465 38 -463
rect 37 -471 38 -469
rect 44 -465 45 -463
rect 44 -471 45 -469
rect 54 -465 55 -463
rect 54 -471 55 -469
rect 58 -465 59 -463
rect 58 -471 59 -469
rect 65 -465 66 -463
rect 65 -471 66 -469
rect 72 -465 73 -463
rect 72 -471 73 -469
rect 79 -465 80 -463
rect 79 -471 80 -469
rect 86 -465 87 -463
rect 86 -471 87 -469
rect 96 -465 97 -463
rect 93 -471 94 -469
rect 96 -471 97 -469
rect 100 -465 101 -463
rect 100 -471 101 -469
rect 107 -465 108 -463
rect 107 -471 108 -469
rect 114 -471 115 -469
rect 121 -465 122 -463
rect 121 -471 122 -469
rect 124 -471 125 -469
rect 128 -471 129 -469
rect 131 -471 132 -469
rect 135 -465 136 -463
rect 135 -471 136 -469
rect 142 -465 143 -463
rect 142 -471 143 -469
rect 149 -471 150 -469
rect 152 -471 153 -469
rect 159 -465 160 -463
rect 156 -471 157 -469
rect 166 -465 167 -463
rect 163 -471 164 -469
rect 170 -465 171 -463
rect 173 -465 174 -463
rect 170 -471 171 -469
rect 177 -465 178 -463
rect 177 -471 178 -469
rect 184 -471 185 -469
rect 191 -465 192 -463
rect 191 -471 192 -469
rect 198 -465 199 -463
rect 201 -465 202 -463
rect 201 -471 202 -469
rect 205 -465 206 -463
rect 205 -471 206 -469
rect 212 -465 213 -463
rect 212 -471 213 -469
rect 219 -465 220 -463
rect 222 -465 223 -463
rect 219 -471 220 -469
rect 229 -465 230 -463
rect 229 -471 230 -469
rect 233 -465 234 -463
rect 233 -471 234 -469
rect 240 -465 241 -463
rect 243 -465 244 -463
rect 240 -471 241 -469
rect 247 -465 248 -463
rect 247 -471 248 -469
rect 254 -465 255 -463
rect 261 -471 262 -469
rect 264 -471 265 -469
rect 268 -465 269 -463
rect 268 -471 269 -469
rect 275 -465 276 -463
rect 278 -465 279 -463
rect 278 -471 279 -469
rect 282 -465 283 -463
rect 285 -465 286 -463
rect 282 -471 283 -469
rect 285 -471 286 -469
rect 289 -465 290 -463
rect 289 -471 290 -469
rect 296 -465 297 -463
rect 296 -471 297 -469
rect 303 -465 304 -463
rect 303 -471 304 -469
rect 313 -465 314 -463
rect 310 -471 311 -469
rect 313 -471 314 -469
rect 317 -471 318 -469
rect 320 -471 321 -469
rect 324 -465 325 -463
rect 324 -471 325 -469
rect 331 -465 332 -463
rect 331 -471 332 -469
rect 338 -465 339 -463
rect 338 -471 339 -469
rect 345 -465 346 -463
rect 348 -465 349 -463
rect 352 -465 353 -463
rect 359 -465 360 -463
rect 359 -471 360 -469
rect 366 -471 367 -469
rect 373 -471 374 -469
rect 380 -465 381 -463
rect 380 -471 381 -469
rect 387 -465 388 -463
rect 387 -471 388 -469
rect 394 -465 395 -463
rect 397 -465 398 -463
rect 394 -471 395 -469
rect 401 -465 402 -463
rect 401 -471 402 -469
rect 408 -465 409 -463
rect 408 -471 409 -469
rect 415 -465 416 -463
rect 415 -471 416 -469
rect 422 -465 423 -463
rect 422 -471 423 -469
rect 429 -465 430 -463
rect 429 -471 430 -469
rect 436 -465 437 -463
rect 436 -471 437 -469
rect 443 -465 444 -463
rect 443 -471 444 -469
rect 450 -465 451 -463
rect 450 -471 451 -469
rect 457 -465 458 -463
rect 457 -471 458 -469
rect 464 -465 465 -463
rect 464 -471 465 -469
rect 471 -465 472 -463
rect 471 -471 472 -469
rect 478 -465 479 -463
rect 478 -471 479 -469
rect 485 -465 486 -463
rect 485 -471 486 -469
rect 492 -465 493 -463
rect 492 -471 493 -469
rect 499 -465 500 -463
rect 499 -471 500 -469
rect 506 -465 507 -463
rect 506 -471 507 -469
rect 513 -465 514 -463
rect 513 -471 514 -469
rect 520 -465 521 -463
rect 520 -471 521 -469
rect 527 -465 528 -463
rect 527 -471 528 -469
rect 534 -465 535 -463
rect 534 -471 535 -469
rect 541 -465 542 -463
rect 541 -471 542 -469
rect 548 -465 549 -463
rect 548 -471 549 -469
rect 555 -471 556 -469
rect 558 -471 559 -469
rect 562 -465 563 -463
rect 562 -471 563 -469
rect 572 -471 573 -469
rect 576 -465 577 -463
rect 576 -471 577 -469
rect 16 -522 17 -520
rect 16 -528 17 -526
rect 23 -522 24 -520
rect 23 -528 24 -526
rect 30 -522 31 -520
rect 30 -528 31 -526
rect 37 -522 38 -520
rect 37 -528 38 -526
rect 44 -522 45 -520
rect 44 -528 45 -526
rect 51 -522 52 -520
rect 51 -528 52 -526
rect 58 -522 59 -520
rect 58 -528 59 -526
rect 65 -522 66 -520
rect 68 -528 69 -526
rect 75 -522 76 -520
rect 75 -528 76 -526
rect 79 -522 80 -520
rect 82 -522 83 -520
rect 86 -522 87 -520
rect 89 -522 90 -520
rect 89 -528 90 -526
rect 93 -522 94 -520
rect 93 -528 94 -526
rect 100 -522 101 -520
rect 100 -528 101 -526
rect 107 -522 108 -520
rect 107 -528 108 -526
rect 117 -522 118 -520
rect 114 -528 115 -526
rect 124 -522 125 -520
rect 121 -528 122 -526
rect 124 -528 125 -526
rect 128 -528 129 -526
rect 131 -528 132 -526
rect 138 -528 139 -526
rect 145 -528 146 -526
rect 149 -522 150 -520
rect 149 -528 150 -526
rect 159 -522 160 -520
rect 156 -528 157 -526
rect 159 -528 160 -526
rect 163 -522 164 -520
rect 163 -528 164 -526
rect 170 -522 171 -520
rect 170 -528 171 -526
rect 177 -522 178 -520
rect 177 -528 178 -526
rect 184 -522 185 -520
rect 187 -528 188 -526
rect 191 -522 192 -520
rect 191 -528 192 -526
rect 201 -522 202 -520
rect 201 -528 202 -526
rect 205 -522 206 -520
rect 205 -528 206 -526
rect 212 -522 213 -520
rect 212 -528 213 -526
rect 219 -522 220 -520
rect 222 -522 223 -520
rect 219 -528 220 -526
rect 226 -522 227 -520
rect 229 -522 230 -520
rect 226 -528 227 -526
rect 233 -522 234 -520
rect 233 -528 234 -526
rect 240 -522 241 -520
rect 243 -522 244 -520
rect 240 -528 241 -526
rect 247 -522 248 -520
rect 247 -528 248 -526
rect 254 -522 255 -520
rect 254 -528 255 -526
rect 261 -522 262 -520
rect 264 -522 265 -520
rect 261 -528 262 -526
rect 264 -528 265 -526
rect 268 -522 269 -520
rect 268 -528 269 -526
rect 275 -522 276 -520
rect 278 -528 279 -526
rect 282 -522 283 -520
rect 285 -522 286 -520
rect 285 -528 286 -526
rect 289 -522 290 -520
rect 292 -522 293 -520
rect 292 -528 293 -526
rect 296 -522 297 -520
rect 299 -522 300 -520
rect 299 -528 300 -526
rect 303 -522 304 -520
rect 303 -528 304 -526
rect 310 -522 311 -520
rect 310 -528 311 -526
rect 313 -528 314 -526
rect 317 -522 318 -520
rect 317 -528 318 -526
rect 324 -528 325 -526
rect 331 -522 332 -520
rect 331 -528 332 -526
rect 338 -522 339 -520
rect 338 -528 339 -526
rect 345 -522 346 -520
rect 348 -528 349 -526
rect 355 -522 356 -520
rect 352 -528 353 -526
rect 359 -522 360 -520
rect 359 -528 360 -526
rect 366 -522 367 -520
rect 369 -522 370 -520
rect 373 -528 374 -526
rect 376 -528 377 -526
rect 380 -522 381 -520
rect 380 -528 381 -526
rect 390 -522 391 -520
rect 394 -522 395 -520
rect 394 -528 395 -526
rect 401 -522 402 -520
rect 401 -528 402 -526
rect 408 -522 409 -520
rect 408 -528 409 -526
rect 415 -522 416 -520
rect 415 -528 416 -526
rect 425 -522 426 -520
rect 429 -522 430 -520
rect 429 -528 430 -526
rect 436 -522 437 -520
rect 436 -528 437 -526
rect 443 -522 444 -520
rect 443 -528 444 -526
rect 450 -522 451 -520
rect 450 -528 451 -526
rect 457 -522 458 -520
rect 457 -528 458 -526
rect 464 -522 465 -520
rect 464 -528 465 -526
rect 471 -522 472 -520
rect 471 -528 472 -526
rect 478 -522 479 -520
rect 478 -528 479 -526
rect 485 -522 486 -520
rect 485 -528 486 -526
rect 492 -522 493 -520
rect 492 -528 493 -526
rect 499 -522 500 -520
rect 499 -528 500 -526
rect 509 -522 510 -520
rect 506 -528 507 -526
rect 509 -528 510 -526
rect 513 -522 514 -520
rect 513 -528 514 -526
rect 520 -522 521 -520
rect 520 -528 521 -526
rect 541 -522 542 -520
rect 541 -528 542 -526
rect 562 -522 563 -520
rect 562 -528 563 -526
rect 9 -571 10 -569
rect 9 -577 10 -575
rect 16 -571 17 -569
rect 23 -577 24 -575
rect 30 -571 31 -569
rect 30 -577 31 -575
rect 40 -571 41 -569
rect 44 -577 45 -575
rect 51 -571 52 -569
rect 51 -577 52 -575
rect 58 -571 59 -569
rect 58 -577 59 -575
rect 68 -571 69 -569
rect 65 -577 66 -575
rect 72 -571 73 -569
rect 72 -577 73 -575
rect 79 -571 80 -569
rect 79 -577 80 -575
rect 86 -577 87 -575
rect 89 -577 90 -575
rect 93 -571 94 -569
rect 93 -577 94 -575
rect 103 -571 104 -569
rect 100 -577 101 -575
rect 107 -571 108 -569
rect 110 -577 111 -575
rect 117 -571 118 -569
rect 114 -577 115 -575
rect 117 -577 118 -575
rect 121 -571 122 -569
rect 121 -577 122 -575
rect 128 -571 129 -569
rect 128 -577 129 -575
rect 135 -571 136 -569
rect 135 -577 136 -575
rect 142 -571 143 -569
rect 142 -577 143 -575
rect 149 -571 150 -569
rect 149 -577 150 -575
rect 156 -571 157 -569
rect 156 -577 157 -575
rect 163 -571 164 -569
rect 163 -577 164 -575
rect 170 -571 171 -569
rect 173 -577 174 -575
rect 177 -571 178 -569
rect 177 -577 178 -575
rect 184 -571 185 -569
rect 187 -577 188 -575
rect 191 -571 192 -569
rect 191 -577 192 -575
rect 198 -571 199 -569
rect 198 -577 199 -575
rect 205 -571 206 -569
rect 208 -571 209 -569
rect 205 -577 206 -575
rect 208 -577 209 -575
rect 215 -571 216 -569
rect 219 -571 220 -569
rect 222 -571 223 -569
rect 219 -577 220 -575
rect 229 -571 230 -569
rect 229 -577 230 -575
rect 236 -571 237 -569
rect 233 -577 234 -575
rect 236 -577 237 -575
rect 240 -571 241 -569
rect 247 -571 248 -569
rect 247 -577 248 -575
rect 254 -571 255 -569
rect 257 -571 258 -569
rect 261 -571 262 -569
rect 261 -577 262 -575
rect 268 -571 269 -569
rect 271 -571 272 -569
rect 268 -577 269 -575
rect 271 -577 272 -575
rect 275 -571 276 -569
rect 275 -577 276 -575
rect 282 -571 283 -569
rect 285 -577 286 -575
rect 289 -571 290 -569
rect 289 -577 290 -575
rect 296 -571 297 -569
rect 296 -577 297 -575
rect 306 -571 307 -569
rect 306 -577 307 -575
rect 313 -571 314 -569
rect 313 -577 314 -575
rect 317 -571 318 -569
rect 317 -577 318 -575
rect 324 -571 325 -569
rect 324 -577 325 -575
rect 331 -571 332 -569
rect 331 -577 332 -575
rect 338 -571 339 -569
rect 341 -571 342 -569
rect 338 -577 339 -575
rect 345 -571 346 -569
rect 345 -577 346 -575
rect 352 -571 353 -569
rect 352 -577 353 -575
rect 359 -571 360 -569
rect 362 -571 363 -569
rect 359 -577 360 -575
rect 362 -577 363 -575
rect 366 -571 367 -569
rect 369 -571 370 -569
rect 373 -571 374 -569
rect 373 -577 374 -575
rect 380 -571 381 -569
rect 380 -577 381 -575
rect 387 -571 388 -569
rect 387 -577 388 -575
rect 394 -571 395 -569
rect 394 -577 395 -575
rect 401 -571 402 -569
rect 401 -577 402 -575
rect 408 -571 409 -569
rect 408 -577 409 -575
rect 415 -571 416 -569
rect 415 -577 416 -575
rect 422 -571 423 -569
rect 422 -577 423 -575
rect 429 -571 430 -569
rect 432 -577 433 -575
rect 436 -571 437 -569
rect 436 -577 437 -575
rect 443 -571 444 -569
rect 443 -577 444 -575
rect 450 -571 451 -569
rect 450 -577 451 -575
rect 457 -571 458 -569
rect 457 -577 458 -575
rect 464 -571 465 -569
rect 464 -577 465 -575
rect 471 -571 472 -569
rect 471 -577 472 -575
rect 478 -571 479 -569
rect 478 -577 479 -575
rect 485 -571 486 -569
rect 485 -577 486 -575
rect 492 -571 493 -569
rect 492 -577 493 -575
rect 499 -577 500 -575
rect 506 -571 507 -569
rect 506 -577 507 -575
rect 513 -577 514 -575
rect 520 -571 521 -569
rect 520 -577 521 -575
rect 527 -571 528 -569
rect 530 -571 531 -569
rect 527 -577 528 -575
rect 530 -577 531 -575
rect 534 -571 535 -569
rect 534 -577 535 -575
rect 541 -571 542 -569
rect 541 -577 542 -575
rect 548 -577 549 -575
rect 555 -571 556 -569
rect 555 -577 556 -575
rect 562 -571 563 -569
rect 562 -577 563 -575
rect 9 -614 10 -612
rect 9 -620 10 -618
rect 16 -614 17 -612
rect 16 -620 17 -618
rect 23 -614 24 -612
rect 23 -620 24 -618
rect 30 -614 31 -612
rect 30 -620 31 -618
rect 37 -614 38 -612
rect 37 -620 38 -618
rect 44 -620 45 -618
rect 47 -620 48 -618
rect 51 -614 52 -612
rect 54 -614 55 -612
rect 58 -614 59 -612
rect 58 -620 59 -618
rect 65 -614 66 -612
rect 68 -620 69 -618
rect 72 -614 73 -612
rect 72 -620 73 -618
rect 79 -614 80 -612
rect 82 -614 83 -612
rect 86 -620 87 -618
rect 89 -620 90 -618
rect 93 -614 94 -612
rect 93 -620 94 -618
rect 103 -614 104 -612
rect 103 -620 104 -618
rect 107 -614 108 -612
rect 107 -620 108 -618
rect 114 -620 115 -618
rect 121 -614 122 -612
rect 121 -620 122 -618
rect 131 -614 132 -612
rect 131 -620 132 -618
rect 135 -614 136 -612
rect 138 -614 139 -612
rect 142 -614 143 -612
rect 145 -614 146 -612
rect 142 -620 143 -618
rect 149 -614 150 -612
rect 149 -620 150 -618
rect 156 -614 157 -612
rect 156 -620 157 -618
rect 163 -614 164 -612
rect 163 -620 164 -618
rect 170 -614 171 -612
rect 170 -620 171 -618
rect 177 -620 178 -618
rect 180 -620 181 -618
rect 187 -620 188 -618
rect 191 -614 192 -612
rect 191 -620 192 -618
rect 198 -614 199 -612
rect 198 -620 199 -618
rect 205 -614 206 -612
rect 205 -620 206 -618
rect 212 -614 213 -612
rect 212 -620 213 -618
rect 219 -614 220 -612
rect 222 -614 223 -612
rect 219 -620 220 -618
rect 222 -620 223 -618
rect 226 -614 227 -612
rect 229 -614 230 -612
rect 226 -620 227 -618
rect 233 -614 234 -612
rect 233 -620 234 -618
rect 240 -614 241 -612
rect 240 -620 241 -618
rect 247 -614 248 -612
rect 247 -620 248 -618
rect 254 -614 255 -612
rect 254 -620 255 -618
rect 261 -614 262 -612
rect 261 -620 262 -618
rect 268 -614 269 -612
rect 268 -620 269 -618
rect 275 -614 276 -612
rect 275 -620 276 -618
rect 282 -614 283 -612
rect 282 -620 283 -618
rect 289 -614 290 -612
rect 289 -620 290 -618
rect 292 -620 293 -618
rect 299 -614 300 -612
rect 296 -620 297 -618
rect 299 -620 300 -618
rect 303 -614 304 -612
rect 303 -620 304 -618
rect 310 -614 311 -612
rect 310 -620 311 -618
rect 317 -614 318 -612
rect 317 -620 318 -618
rect 327 -614 328 -612
rect 324 -620 325 -618
rect 327 -620 328 -618
rect 331 -614 332 -612
rect 331 -620 332 -618
rect 338 -614 339 -612
rect 341 -614 342 -612
rect 341 -620 342 -618
rect 345 -614 346 -612
rect 345 -620 346 -618
rect 352 -614 353 -612
rect 352 -620 353 -618
rect 355 -620 356 -618
rect 359 -614 360 -612
rect 359 -620 360 -618
rect 366 -614 367 -612
rect 366 -620 367 -618
rect 373 -614 374 -612
rect 373 -620 374 -618
rect 380 -614 381 -612
rect 380 -620 381 -618
rect 387 -614 388 -612
rect 387 -620 388 -618
rect 394 -614 395 -612
rect 394 -620 395 -618
rect 397 -620 398 -618
rect 401 -614 402 -612
rect 401 -620 402 -618
rect 408 -614 409 -612
rect 408 -620 409 -618
rect 418 -620 419 -618
rect 422 -614 423 -612
rect 422 -620 423 -618
rect 429 -614 430 -612
rect 429 -620 430 -618
rect 436 -614 437 -612
rect 436 -620 437 -618
rect 443 -614 444 -612
rect 443 -620 444 -618
rect 450 -614 451 -612
rect 450 -620 451 -618
rect 457 -614 458 -612
rect 457 -620 458 -618
rect 464 -614 465 -612
rect 464 -620 465 -618
rect 471 -614 472 -612
rect 471 -620 472 -618
rect 481 -614 482 -612
rect 481 -620 482 -618
rect 485 -614 486 -612
rect 485 -620 486 -618
rect 492 -614 493 -612
rect 492 -620 493 -618
rect 499 -614 500 -612
rect 499 -620 500 -618
rect 509 -614 510 -612
rect 513 -614 514 -612
rect 516 -614 517 -612
rect 516 -620 517 -618
rect 520 -614 521 -612
rect 523 -614 524 -612
rect 527 -614 528 -612
rect 527 -620 528 -618
rect 534 -614 535 -612
rect 534 -620 535 -618
rect 541 -614 542 -612
rect 541 -620 542 -618
rect 548 -614 549 -612
rect 548 -620 549 -618
rect 555 -614 556 -612
rect 555 -620 556 -618
rect 562 -614 563 -612
rect 40 -661 41 -659
rect 44 -661 45 -659
rect 44 -667 45 -665
rect 51 -661 52 -659
rect 51 -667 52 -665
rect 61 -661 62 -659
rect 58 -667 59 -665
rect 65 -661 66 -659
rect 65 -667 66 -665
rect 72 -661 73 -659
rect 75 -661 76 -659
rect 79 -661 80 -659
rect 79 -667 80 -665
rect 86 -661 87 -659
rect 86 -667 87 -665
rect 96 -661 97 -659
rect 100 -661 101 -659
rect 100 -667 101 -665
rect 103 -667 104 -665
rect 107 -661 108 -659
rect 107 -667 108 -665
rect 114 -661 115 -659
rect 117 -661 118 -659
rect 114 -667 115 -665
rect 121 -661 122 -659
rect 121 -667 122 -665
rect 128 -661 129 -659
rect 131 -661 132 -659
rect 135 -661 136 -659
rect 135 -667 136 -665
rect 142 -667 143 -665
rect 149 -661 150 -659
rect 149 -667 150 -665
rect 156 -661 157 -659
rect 156 -667 157 -665
rect 163 -661 164 -659
rect 163 -667 164 -665
rect 170 -661 171 -659
rect 170 -667 171 -665
rect 177 -661 178 -659
rect 177 -667 178 -665
rect 184 -661 185 -659
rect 184 -667 185 -665
rect 191 -661 192 -659
rect 191 -667 192 -665
rect 201 -667 202 -665
rect 208 -661 209 -659
rect 205 -667 206 -665
rect 212 -661 213 -659
rect 212 -667 213 -665
rect 219 -661 220 -659
rect 219 -667 220 -665
rect 226 -661 227 -659
rect 226 -667 227 -665
rect 233 -661 234 -659
rect 233 -667 234 -665
rect 243 -667 244 -665
rect 247 -661 248 -659
rect 250 -661 251 -659
rect 247 -667 248 -665
rect 250 -667 251 -665
rect 254 -661 255 -659
rect 254 -667 255 -665
rect 261 -661 262 -659
rect 261 -667 262 -665
rect 268 -667 269 -665
rect 271 -667 272 -665
rect 275 -661 276 -659
rect 275 -667 276 -665
rect 282 -661 283 -659
rect 282 -667 283 -665
rect 289 -661 290 -659
rect 289 -667 290 -665
rect 296 -661 297 -659
rect 296 -667 297 -665
rect 303 -661 304 -659
rect 303 -667 304 -665
rect 310 -661 311 -659
rect 310 -667 311 -665
rect 320 -661 321 -659
rect 320 -667 321 -665
rect 324 -661 325 -659
rect 324 -667 325 -665
rect 331 -661 332 -659
rect 334 -661 335 -659
rect 338 -661 339 -659
rect 341 -661 342 -659
rect 338 -667 339 -665
rect 345 -661 346 -659
rect 348 -661 349 -659
rect 345 -667 346 -665
rect 348 -667 349 -665
rect 352 -661 353 -659
rect 359 -661 360 -659
rect 359 -667 360 -665
rect 366 -661 367 -659
rect 366 -667 367 -665
rect 373 -667 374 -665
rect 376 -667 377 -665
rect 380 -661 381 -659
rect 380 -667 381 -665
rect 387 -661 388 -659
rect 387 -667 388 -665
rect 397 -661 398 -659
rect 394 -667 395 -665
rect 397 -667 398 -665
rect 401 -661 402 -659
rect 401 -667 402 -665
rect 404 -667 405 -665
rect 408 -661 409 -659
rect 408 -667 409 -665
rect 415 -661 416 -659
rect 415 -667 416 -665
rect 422 -661 423 -659
rect 422 -667 423 -665
rect 429 -661 430 -659
rect 429 -667 430 -665
rect 436 -661 437 -659
rect 436 -667 437 -665
rect 443 -661 444 -659
rect 443 -667 444 -665
rect 450 -661 451 -659
rect 450 -667 451 -665
rect 457 -661 458 -659
rect 457 -667 458 -665
rect 464 -661 465 -659
rect 464 -667 465 -665
rect 471 -661 472 -659
rect 474 -661 475 -659
rect 471 -667 472 -665
rect 474 -667 475 -665
rect 478 -661 479 -659
rect 478 -667 479 -665
rect 488 -661 489 -659
rect 488 -667 489 -665
rect 492 -661 493 -659
rect 492 -667 493 -665
rect 499 -661 500 -659
rect 499 -667 500 -665
rect 506 -661 507 -659
rect 506 -667 507 -665
rect 513 -661 514 -659
rect 516 -661 517 -659
rect 516 -667 517 -665
rect 520 -661 521 -659
rect 520 -667 521 -665
rect 530 -661 531 -659
rect 530 -667 531 -665
rect 534 -661 535 -659
rect 534 -667 535 -665
rect 544 -661 545 -659
rect 544 -667 545 -665
rect 548 -661 549 -659
rect 548 -667 549 -665
rect 555 -661 556 -659
rect 555 -667 556 -665
rect 562 -661 563 -659
rect 583 -661 584 -659
rect 583 -667 584 -665
rect 16 -710 17 -708
rect 16 -716 17 -714
rect 23 -710 24 -708
rect 23 -716 24 -714
rect 30 -710 31 -708
rect 37 -710 38 -708
rect 37 -716 38 -714
rect 44 -710 45 -708
rect 44 -716 45 -714
rect 51 -710 52 -708
rect 51 -716 52 -714
rect 58 -716 59 -714
rect 65 -710 66 -708
rect 65 -716 66 -714
rect 72 -710 73 -708
rect 72 -716 73 -714
rect 75 -716 76 -714
rect 79 -710 80 -708
rect 79 -716 80 -714
rect 86 -710 87 -708
rect 86 -716 87 -714
rect 93 -710 94 -708
rect 93 -716 94 -714
rect 103 -710 104 -708
rect 103 -716 104 -714
rect 110 -710 111 -708
rect 107 -716 108 -714
rect 114 -710 115 -708
rect 114 -716 115 -714
rect 121 -710 122 -708
rect 121 -716 122 -714
rect 128 -710 129 -708
rect 128 -716 129 -714
rect 135 -710 136 -708
rect 142 -710 143 -708
rect 142 -716 143 -714
rect 149 -710 150 -708
rect 149 -716 150 -714
rect 152 -716 153 -714
rect 156 -710 157 -708
rect 156 -716 157 -714
rect 163 -710 164 -708
rect 166 -710 167 -708
rect 163 -716 164 -714
rect 170 -710 171 -708
rect 170 -716 171 -714
rect 177 -710 178 -708
rect 177 -716 178 -714
rect 184 -710 185 -708
rect 184 -716 185 -714
rect 187 -716 188 -714
rect 194 -710 195 -708
rect 191 -716 192 -714
rect 194 -716 195 -714
rect 198 -710 199 -708
rect 201 -710 202 -708
rect 198 -716 199 -714
rect 201 -716 202 -714
rect 205 -710 206 -708
rect 205 -716 206 -714
rect 212 -710 213 -708
rect 212 -716 213 -714
rect 219 -710 220 -708
rect 219 -716 220 -714
rect 222 -716 223 -714
rect 226 -710 227 -708
rect 226 -716 227 -714
rect 233 -710 234 -708
rect 233 -716 234 -714
rect 240 -710 241 -708
rect 240 -716 241 -714
rect 247 -710 248 -708
rect 247 -716 248 -714
rect 254 -710 255 -708
rect 254 -716 255 -714
rect 261 -710 262 -708
rect 261 -716 262 -714
rect 268 -710 269 -708
rect 268 -716 269 -714
rect 275 -710 276 -708
rect 275 -716 276 -714
rect 282 -716 283 -714
rect 289 -710 290 -708
rect 289 -716 290 -714
rect 296 -710 297 -708
rect 299 -710 300 -708
rect 296 -716 297 -714
rect 303 -710 304 -708
rect 303 -716 304 -714
rect 310 -710 311 -708
rect 310 -716 311 -714
rect 317 -710 318 -708
rect 317 -716 318 -714
rect 324 -710 325 -708
rect 324 -716 325 -714
rect 331 -710 332 -708
rect 334 -710 335 -708
rect 331 -716 332 -714
rect 334 -716 335 -714
rect 338 -710 339 -708
rect 338 -716 339 -714
rect 345 -710 346 -708
rect 345 -716 346 -714
rect 348 -716 349 -714
rect 352 -710 353 -708
rect 352 -716 353 -714
rect 359 -710 360 -708
rect 359 -716 360 -714
rect 366 -710 367 -708
rect 366 -716 367 -714
rect 373 -710 374 -708
rect 373 -716 374 -714
rect 380 -710 381 -708
rect 380 -716 381 -714
rect 383 -716 384 -714
rect 387 -710 388 -708
rect 387 -716 388 -714
rect 394 -716 395 -714
rect 397 -716 398 -714
rect 401 -710 402 -708
rect 401 -716 402 -714
rect 408 -710 409 -708
rect 408 -716 409 -714
rect 415 -710 416 -708
rect 415 -716 416 -714
rect 422 -710 423 -708
rect 425 -716 426 -714
rect 429 -710 430 -708
rect 429 -716 430 -714
rect 436 -710 437 -708
rect 436 -716 437 -714
rect 443 -710 444 -708
rect 443 -716 444 -714
rect 450 -710 451 -708
rect 450 -716 451 -714
rect 457 -710 458 -708
rect 457 -716 458 -714
rect 464 -710 465 -708
rect 464 -716 465 -714
rect 471 -710 472 -708
rect 471 -716 472 -714
rect 478 -710 479 -708
rect 478 -716 479 -714
rect 485 -710 486 -708
rect 485 -716 486 -714
rect 495 -716 496 -714
rect 499 -710 500 -708
rect 499 -716 500 -714
rect 506 -710 507 -708
rect 506 -716 507 -714
rect 513 -710 514 -708
rect 513 -716 514 -714
rect 520 -710 521 -708
rect 520 -716 521 -714
rect 527 -710 528 -708
rect 527 -716 528 -714
rect 534 -710 535 -708
rect 534 -716 535 -714
rect 541 -710 542 -708
rect 541 -716 542 -714
rect 548 -710 549 -708
rect 548 -716 549 -714
rect 555 -710 556 -708
rect 555 -716 556 -714
rect 562 -710 563 -708
rect 562 -716 563 -714
rect 572 -710 573 -708
rect 569 -716 570 -714
rect 572 -716 573 -714
rect 576 -710 577 -708
rect 576 -716 577 -714
rect 583 -710 584 -708
rect 583 -716 584 -714
rect 593 -710 594 -708
rect 593 -716 594 -714
rect 597 -716 598 -714
rect 600 -716 601 -714
rect 604 -710 605 -708
rect 604 -716 605 -714
rect 611 -710 612 -708
rect 614 -716 615 -714
rect 618 -710 619 -708
rect 618 -716 619 -714
rect 628 -710 629 -708
rect 632 -710 633 -708
rect 632 -716 633 -714
rect 639 -710 640 -708
rect 639 -716 640 -714
rect 646 -710 647 -708
rect 646 -716 647 -714
rect 33 -761 34 -759
rect 33 -767 34 -765
rect 40 -767 41 -765
rect 44 -761 45 -759
rect 44 -767 45 -765
rect 51 -761 52 -759
rect 51 -767 52 -765
rect 58 -761 59 -759
rect 58 -767 59 -765
rect 65 -761 66 -759
rect 65 -767 66 -765
rect 72 -761 73 -759
rect 72 -767 73 -765
rect 79 -761 80 -759
rect 79 -767 80 -765
rect 86 -761 87 -759
rect 86 -767 87 -765
rect 93 -761 94 -759
rect 93 -767 94 -765
rect 103 -761 104 -759
rect 107 -761 108 -759
rect 107 -767 108 -765
rect 114 -761 115 -759
rect 117 -767 118 -765
rect 121 -761 122 -759
rect 121 -767 122 -765
rect 128 -761 129 -759
rect 128 -767 129 -765
rect 135 -761 136 -759
rect 135 -767 136 -765
rect 142 -761 143 -759
rect 145 -767 146 -765
rect 149 -761 150 -759
rect 152 -761 153 -759
rect 149 -767 150 -765
rect 152 -767 153 -765
rect 156 -761 157 -759
rect 156 -767 157 -765
rect 163 -761 164 -759
rect 163 -767 164 -765
rect 170 -761 171 -759
rect 170 -767 171 -765
rect 177 -761 178 -759
rect 177 -767 178 -765
rect 184 -761 185 -759
rect 184 -767 185 -765
rect 194 -761 195 -759
rect 191 -767 192 -765
rect 194 -767 195 -765
rect 198 -761 199 -759
rect 198 -767 199 -765
rect 205 -761 206 -759
rect 205 -767 206 -765
rect 215 -761 216 -759
rect 212 -767 213 -765
rect 215 -767 216 -765
rect 222 -761 223 -759
rect 219 -767 220 -765
rect 222 -767 223 -765
rect 229 -761 230 -759
rect 226 -767 227 -765
rect 229 -767 230 -765
rect 233 -761 234 -759
rect 233 -767 234 -765
rect 240 -761 241 -759
rect 240 -767 241 -765
rect 250 -761 251 -759
rect 247 -767 248 -765
rect 254 -761 255 -759
rect 257 -761 258 -759
rect 257 -767 258 -765
rect 261 -761 262 -759
rect 261 -767 262 -765
rect 268 -761 269 -759
rect 268 -767 269 -765
rect 278 -761 279 -759
rect 275 -767 276 -765
rect 285 -761 286 -759
rect 285 -767 286 -765
rect 292 -761 293 -759
rect 292 -767 293 -765
rect 296 -761 297 -759
rect 296 -767 297 -765
rect 303 -761 304 -759
rect 303 -767 304 -765
rect 306 -767 307 -765
rect 310 -761 311 -759
rect 310 -767 311 -765
rect 317 -761 318 -759
rect 317 -767 318 -765
rect 324 -761 325 -759
rect 324 -767 325 -765
rect 331 -761 332 -759
rect 334 -761 335 -759
rect 331 -767 332 -765
rect 338 -761 339 -759
rect 338 -767 339 -765
rect 341 -767 342 -765
rect 348 -761 349 -759
rect 352 -761 353 -759
rect 352 -767 353 -765
rect 359 -761 360 -759
rect 362 -761 363 -759
rect 359 -767 360 -765
rect 366 -761 367 -759
rect 366 -767 367 -765
rect 373 -767 374 -765
rect 376 -767 377 -765
rect 380 -761 381 -759
rect 380 -767 381 -765
rect 387 -761 388 -759
rect 387 -767 388 -765
rect 394 -761 395 -759
rect 397 -767 398 -765
rect 401 -761 402 -759
rect 401 -767 402 -765
rect 408 -761 409 -759
rect 408 -767 409 -765
rect 415 -761 416 -759
rect 415 -767 416 -765
rect 422 -761 423 -759
rect 422 -767 423 -765
rect 429 -761 430 -759
rect 429 -767 430 -765
rect 436 -761 437 -759
rect 436 -767 437 -765
rect 443 -767 444 -765
rect 446 -767 447 -765
rect 450 -761 451 -759
rect 450 -767 451 -765
rect 457 -761 458 -759
rect 457 -767 458 -765
rect 464 -761 465 -759
rect 464 -767 465 -765
rect 471 -761 472 -759
rect 474 -761 475 -759
rect 471 -767 472 -765
rect 478 -761 479 -759
rect 478 -767 479 -765
rect 485 -761 486 -759
rect 488 -761 489 -759
rect 492 -761 493 -759
rect 492 -767 493 -765
rect 499 -761 500 -759
rect 499 -767 500 -765
rect 506 -761 507 -759
rect 506 -767 507 -765
rect 513 -761 514 -759
rect 513 -767 514 -765
rect 520 -761 521 -759
rect 520 -767 521 -765
rect 527 -761 528 -759
rect 530 -761 531 -759
rect 530 -767 531 -765
rect 534 -761 535 -759
rect 534 -767 535 -765
rect 541 -761 542 -759
rect 541 -767 542 -765
rect 555 -761 556 -759
rect 555 -767 556 -765
rect 611 -761 612 -759
rect 26 -818 27 -816
rect 30 -818 31 -816
rect 37 -818 38 -816
rect 37 -824 38 -822
rect 44 -818 45 -816
rect 44 -824 45 -822
rect 51 -818 52 -816
rect 51 -824 52 -822
rect 58 -818 59 -816
rect 65 -818 66 -816
rect 65 -824 66 -822
rect 72 -818 73 -816
rect 79 -818 80 -816
rect 79 -824 80 -822
rect 86 -818 87 -816
rect 86 -824 87 -822
rect 93 -818 94 -816
rect 93 -824 94 -822
rect 103 -818 104 -816
rect 107 -818 108 -816
rect 110 -824 111 -822
rect 114 -818 115 -816
rect 121 -818 122 -816
rect 124 -824 125 -822
rect 128 -818 129 -816
rect 128 -824 129 -822
rect 135 -818 136 -816
rect 135 -824 136 -822
rect 142 -818 143 -816
rect 145 -818 146 -816
rect 145 -824 146 -822
rect 152 -818 153 -816
rect 149 -824 150 -822
rect 152 -824 153 -822
rect 156 -818 157 -816
rect 159 -824 160 -822
rect 163 -818 164 -816
rect 166 -818 167 -816
rect 163 -824 164 -822
rect 170 -818 171 -816
rect 170 -824 171 -822
rect 177 -818 178 -816
rect 177 -824 178 -822
rect 187 -818 188 -816
rect 187 -824 188 -822
rect 191 -818 192 -816
rect 191 -824 192 -822
rect 198 -824 199 -822
rect 201 -824 202 -822
rect 205 -818 206 -816
rect 205 -824 206 -822
rect 212 -818 213 -816
rect 215 -818 216 -816
rect 219 -818 220 -816
rect 219 -824 220 -822
rect 226 -818 227 -816
rect 226 -824 227 -822
rect 236 -818 237 -816
rect 233 -824 234 -822
rect 236 -824 237 -822
rect 240 -818 241 -816
rect 240 -824 241 -822
rect 247 -818 248 -816
rect 247 -824 248 -822
rect 254 -818 255 -816
rect 257 -818 258 -816
rect 257 -824 258 -822
rect 261 -818 262 -816
rect 261 -824 262 -822
rect 268 -818 269 -816
rect 268 -824 269 -822
rect 275 -818 276 -816
rect 275 -824 276 -822
rect 282 -818 283 -816
rect 282 -824 283 -822
rect 289 -818 290 -816
rect 289 -824 290 -822
rect 296 -818 297 -816
rect 296 -824 297 -822
rect 303 -818 304 -816
rect 303 -824 304 -822
rect 313 -818 314 -816
rect 310 -824 311 -822
rect 313 -824 314 -822
rect 317 -818 318 -816
rect 317 -824 318 -822
rect 320 -824 321 -822
rect 324 -818 325 -816
rect 324 -824 325 -822
rect 331 -818 332 -816
rect 334 -818 335 -816
rect 338 -818 339 -816
rect 338 -824 339 -822
rect 348 -824 349 -822
rect 352 -818 353 -816
rect 355 -824 356 -822
rect 359 -818 360 -816
rect 359 -824 360 -822
rect 366 -818 367 -816
rect 366 -824 367 -822
rect 376 -818 377 -816
rect 373 -824 374 -822
rect 376 -824 377 -822
rect 380 -818 381 -816
rect 380 -824 381 -822
rect 387 -818 388 -816
rect 387 -824 388 -822
rect 394 -818 395 -816
rect 394 -824 395 -822
rect 404 -818 405 -816
rect 401 -824 402 -822
rect 404 -824 405 -822
rect 408 -818 409 -816
rect 408 -824 409 -822
rect 415 -818 416 -816
rect 415 -824 416 -822
rect 422 -818 423 -816
rect 422 -824 423 -822
rect 429 -818 430 -816
rect 429 -824 430 -822
rect 436 -818 437 -816
rect 436 -824 437 -822
rect 443 -818 444 -816
rect 443 -824 444 -822
rect 450 -818 451 -816
rect 450 -824 451 -822
rect 460 -818 461 -816
rect 464 -818 465 -816
rect 464 -824 465 -822
rect 471 -818 472 -816
rect 471 -824 472 -822
rect 478 -818 479 -816
rect 478 -824 479 -822
rect 485 -818 486 -816
rect 485 -824 486 -822
rect 492 -818 493 -816
rect 492 -824 493 -822
rect 499 -818 500 -816
rect 499 -824 500 -822
rect 506 -818 507 -816
rect 506 -824 507 -822
rect 513 -818 514 -816
rect 513 -824 514 -822
rect 520 -818 521 -816
rect 520 -824 521 -822
rect 527 -818 528 -816
rect 527 -824 528 -822
rect 534 -818 535 -816
rect 534 -824 535 -822
rect 541 -818 542 -816
rect 541 -824 542 -822
rect 548 -818 549 -816
rect 548 -824 549 -822
rect 555 -818 556 -816
rect 558 -818 559 -816
rect 558 -824 559 -822
rect 26 -881 27 -879
rect 30 -881 31 -879
rect 37 -881 38 -879
rect 40 -881 41 -879
rect 44 -881 45 -879
rect 44 -887 45 -885
rect 51 -881 52 -879
rect 51 -887 52 -885
rect 58 -881 59 -879
rect 58 -887 59 -885
rect 65 -881 66 -879
rect 65 -887 66 -885
rect 72 -881 73 -879
rect 75 -881 76 -879
rect 79 -881 80 -879
rect 79 -887 80 -885
rect 86 -881 87 -879
rect 86 -887 87 -885
rect 93 -881 94 -879
rect 93 -887 94 -885
rect 100 -881 101 -879
rect 100 -887 101 -885
rect 107 -881 108 -879
rect 107 -887 108 -885
rect 114 -881 115 -879
rect 117 -881 118 -879
rect 121 -881 122 -879
rect 124 -887 125 -885
rect 128 -881 129 -879
rect 128 -887 129 -885
rect 138 -887 139 -885
rect 142 -881 143 -879
rect 142 -887 143 -885
rect 149 -881 150 -879
rect 149 -887 150 -885
rect 156 -881 157 -879
rect 156 -887 157 -885
rect 159 -887 160 -885
rect 163 -881 164 -879
rect 163 -887 164 -885
rect 166 -887 167 -885
rect 173 -881 174 -879
rect 170 -887 171 -885
rect 180 -881 181 -879
rect 180 -887 181 -885
rect 184 -881 185 -879
rect 184 -887 185 -885
rect 194 -881 195 -879
rect 191 -887 192 -885
rect 194 -887 195 -885
rect 201 -881 202 -879
rect 201 -887 202 -885
rect 205 -887 206 -885
rect 208 -887 209 -885
rect 212 -881 213 -879
rect 212 -887 213 -885
rect 219 -881 220 -879
rect 219 -887 220 -885
rect 226 -881 227 -879
rect 226 -887 227 -885
rect 233 -881 234 -879
rect 233 -887 234 -885
rect 240 -881 241 -879
rect 240 -887 241 -885
rect 247 -881 248 -879
rect 247 -887 248 -885
rect 254 -881 255 -879
rect 254 -887 255 -885
rect 261 -881 262 -879
rect 261 -887 262 -885
rect 268 -881 269 -879
rect 268 -887 269 -885
rect 275 -881 276 -879
rect 275 -887 276 -885
rect 285 -881 286 -879
rect 282 -887 283 -885
rect 285 -887 286 -885
rect 289 -881 290 -879
rect 289 -887 290 -885
rect 296 -881 297 -879
rect 296 -887 297 -885
rect 306 -881 307 -879
rect 306 -887 307 -885
rect 310 -881 311 -879
rect 313 -881 314 -879
rect 310 -887 311 -885
rect 313 -887 314 -885
rect 317 -881 318 -879
rect 317 -887 318 -885
rect 324 -881 325 -879
rect 324 -887 325 -885
rect 331 -881 332 -879
rect 334 -881 335 -879
rect 334 -887 335 -885
rect 338 -881 339 -879
rect 338 -887 339 -885
rect 348 -881 349 -879
rect 345 -887 346 -885
rect 348 -887 349 -885
rect 352 -881 353 -879
rect 355 -881 356 -879
rect 352 -887 353 -885
rect 355 -887 356 -885
rect 359 -881 360 -879
rect 359 -887 360 -885
rect 366 -881 367 -879
rect 366 -887 367 -885
rect 373 -881 374 -879
rect 373 -887 374 -885
rect 380 -887 381 -885
rect 383 -887 384 -885
rect 387 -881 388 -879
rect 387 -887 388 -885
rect 394 -881 395 -879
rect 394 -887 395 -885
rect 401 -881 402 -879
rect 401 -887 402 -885
rect 408 -881 409 -879
rect 408 -887 409 -885
rect 415 -881 416 -879
rect 415 -887 416 -885
rect 422 -881 423 -879
rect 422 -887 423 -885
rect 429 -881 430 -879
rect 429 -887 430 -885
rect 436 -881 437 -879
rect 436 -887 437 -885
rect 443 -881 444 -879
rect 443 -887 444 -885
rect 450 -881 451 -879
rect 450 -887 451 -885
rect 457 -881 458 -879
rect 457 -887 458 -885
rect 464 -881 465 -879
rect 467 -881 468 -879
rect 474 -881 475 -879
rect 474 -887 475 -885
rect 478 -881 479 -879
rect 478 -887 479 -885
rect 485 -881 486 -879
rect 485 -887 486 -885
rect 492 -881 493 -879
rect 492 -887 493 -885
rect 499 -881 500 -879
rect 499 -887 500 -885
rect 506 -881 507 -879
rect 506 -887 507 -885
rect 513 -881 514 -879
rect 513 -887 514 -885
rect 520 -887 521 -885
rect 523 -887 524 -885
rect 527 -881 528 -879
rect 527 -887 528 -885
rect 534 -881 535 -879
rect 534 -887 535 -885
rect 9 -936 10 -934
rect 9 -942 10 -940
rect 16 -936 17 -934
rect 16 -942 17 -940
rect 23 -936 24 -934
rect 23 -942 24 -940
rect 30 -942 31 -940
rect 37 -936 38 -934
rect 37 -942 38 -940
rect 44 -936 45 -934
rect 51 -936 52 -934
rect 51 -942 52 -940
rect 58 -936 59 -934
rect 58 -942 59 -940
rect 65 -936 66 -934
rect 65 -942 66 -940
rect 72 -936 73 -934
rect 82 -942 83 -940
rect 86 -942 87 -940
rect 93 -936 94 -934
rect 93 -942 94 -940
rect 100 -942 101 -940
rect 103 -942 104 -940
rect 107 -936 108 -934
rect 107 -942 108 -940
rect 114 -936 115 -934
rect 114 -942 115 -940
rect 121 -936 122 -934
rect 121 -942 122 -940
rect 128 -936 129 -934
rect 128 -942 129 -940
rect 135 -936 136 -934
rect 142 -936 143 -934
rect 142 -942 143 -940
rect 149 -936 150 -934
rect 152 -936 153 -934
rect 159 -936 160 -934
rect 156 -942 157 -940
rect 159 -942 160 -940
rect 166 -936 167 -934
rect 163 -942 164 -940
rect 166 -942 167 -940
rect 170 -936 171 -934
rect 170 -942 171 -940
rect 177 -936 178 -934
rect 177 -942 178 -940
rect 184 -936 185 -934
rect 184 -942 185 -940
rect 194 -936 195 -934
rect 191 -942 192 -940
rect 201 -936 202 -934
rect 198 -942 199 -940
rect 201 -942 202 -940
rect 205 -936 206 -934
rect 208 -936 209 -934
rect 205 -942 206 -940
rect 212 -936 213 -934
rect 212 -942 213 -940
rect 219 -936 220 -934
rect 222 -936 223 -934
rect 219 -942 220 -940
rect 226 -936 227 -934
rect 229 -936 230 -934
rect 226 -942 227 -940
rect 229 -942 230 -940
rect 233 -936 234 -934
rect 233 -942 234 -940
rect 240 -936 241 -934
rect 240 -942 241 -940
rect 247 -936 248 -934
rect 247 -942 248 -940
rect 254 -936 255 -934
rect 254 -942 255 -940
rect 264 -936 265 -934
rect 264 -942 265 -940
rect 268 -936 269 -934
rect 268 -942 269 -940
rect 275 -936 276 -934
rect 275 -942 276 -940
rect 282 -936 283 -934
rect 282 -942 283 -940
rect 292 -936 293 -934
rect 289 -942 290 -940
rect 296 -936 297 -934
rect 296 -942 297 -940
rect 306 -936 307 -934
rect 306 -942 307 -940
rect 310 -936 311 -934
rect 310 -942 311 -940
rect 317 -936 318 -934
rect 317 -942 318 -940
rect 324 -936 325 -934
rect 324 -942 325 -940
rect 327 -942 328 -940
rect 331 -936 332 -934
rect 334 -936 335 -934
rect 334 -942 335 -940
rect 338 -936 339 -934
rect 338 -942 339 -940
rect 345 -936 346 -934
rect 345 -942 346 -940
rect 352 -942 353 -940
rect 359 -936 360 -934
rect 359 -942 360 -940
rect 366 -936 367 -934
rect 366 -942 367 -940
rect 373 -936 374 -934
rect 373 -942 374 -940
rect 380 -936 381 -934
rect 387 -936 388 -934
rect 387 -942 388 -940
rect 397 -936 398 -934
rect 394 -942 395 -940
rect 401 -936 402 -934
rect 401 -942 402 -940
rect 408 -936 409 -934
rect 415 -936 416 -934
rect 415 -942 416 -940
rect 422 -936 423 -934
rect 422 -942 423 -940
rect 429 -936 430 -934
rect 429 -942 430 -940
rect 436 -936 437 -934
rect 436 -942 437 -940
rect 443 -942 444 -940
rect 450 -936 451 -934
rect 450 -942 451 -940
rect 457 -936 458 -934
rect 457 -942 458 -940
rect 464 -942 465 -940
rect 471 -936 472 -934
rect 471 -942 472 -940
rect 478 -936 479 -934
rect 478 -942 479 -940
rect 485 -936 486 -934
rect 485 -942 486 -940
rect 492 -936 493 -934
rect 492 -942 493 -940
rect 499 -936 500 -934
rect 499 -942 500 -940
rect 506 -936 507 -934
rect 506 -942 507 -940
rect 513 -936 514 -934
rect 513 -942 514 -940
rect 520 -936 521 -934
rect 520 -942 521 -940
rect 2 -985 3 -983
rect 2 -991 3 -989
rect 9 -985 10 -983
rect 9 -991 10 -989
rect 16 -985 17 -983
rect 16 -991 17 -989
rect 23 -985 24 -983
rect 30 -985 31 -983
rect 33 -991 34 -989
rect 37 -991 38 -989
rect 40 -991 41 -989
rect 44 -985 45 -983
rect 44 -991 45 -989
rect 51 -985 52 -983
rect 51 -991 52 -989
rect 58 -991 59 -989
rect 61 -991 62 -989
rect 65 -985 66 -983
rect 65 -991 66 -989
rect 75 -985 76 -983
rect 79 -991 80 -989
rect 82 -991 83 -989
rect 86 -985 87 -983
rect 86 -991 87 -989
rect 96 -985 97 -983
rect 93 -991 94 -989
rect 96 -991 97 -989
rect 103 -985 104 -983
rect 103 -991 104 -989
rect 107 -985 108 -983
rect 107 -991 108 -989
rect 114 -985 115 -983
rect 114 -991 115 -989
rect 121 -985 122 -983
rect 121 -991 122 -989
rect 128 -991 129 -989
rect 131 -991 132 -989
rect 135 -985 136 -983
rect 138 -985 139 -983
rect 142 -985 143 -983
rect 142 -991 143 -989
rect 149 -985 150 -983
rect 149 -991 150 -989
rect 159 -985 160 -983
rect 159 -991 160 -989
rect 163 -985 164 -983
rect 166 -985 167 -983
rect 163 -991 164 -989
rect 170 -985 171 -983
rect 170 -991 171 -989
rect 177 -985 178 -983
rect 177 -991 178 -989
rect 184 -985 185 -983
rect 187 -985 188 -983
rect 184 -991 185 -989
rect 187 -991 188 -989
rect 191 -985 192 -983
rect 194 -985 195 -983
rect 191 -991 192 -989
rect 194 -991 195 -989
rect 198 -985 199 -983
rect 201 -985 202 -983
rect 198 -991 199 -989
rect 205 -985 206 -983
rect 205 -991 206 -989
rect 212 -985 213 -983
rect 212 -991 213 -989
rect 219 -985 220 -983
rect 222 -985 223 -983
rect 219 -991 220 -989
rect 222 -991 223 -989
rect 226 -991 227 -989
rect 229 -991 230 -989
rect 233 -985 234 -983
rect 243 -991 244 -989
rect 247 -985 248 -983
rect 247 -991 248 -989
rect 257 -985 258 -983
rect 254 -991 255 -989
rect 261 -985 262 -983
rect 264 -985 265 -983
rect 261 -991 262 -989
rect 268 -985 269 -983
rect 268 -991 269 -989
rect 275 -985 276 -983
rect 275 -991 276 -989
rect 282 -985 283 -983
rect 282 -991 283 -989
rect 292 -985 293 -983
rect 289 -991 290 -989
rect 292 -991 293 -989
rect 296 -985 297 -983
rect 299 -985 300 -983
rect 303 -985 304 -983
rect 303 -991 304 -989
rect 310 -985 311 -983
rect 310 -991 311 -989
rect 317 -985 318 -983
rect 317 -991 318 -989
rect 324 -985 325 -983
rect 324 -991 325 -989
rect 331 -985 332 -983
rect 334 -985 335 -983
rect 338 -985 339 -983
rect 338 -991 339 -989
rect 341 -991 342 -989
rect 345 -985 346 -983
rect 345 -991 346 -989
rect 355 -985 356 -983
rect 352 -991 353 -989
rect 359 -985 360 -983
rect 359 -991 360 -989
rect 366 -985 367 -983
rect 366 -991 367 -989
rect 373 -985 374 -983
rect 373 -991 374 -989
rect 380 -985 381 -983
rect 380 -991 381 -989
rect 387 -985 388 -983
rect 387 -991 388 -989
rect 394 -985 395 -983
rect 394 -991 395 -989
rect 401 -985 402 -983
rect 401 -991 402 -989
rect 408 -985 409 -983
rect 408 -991 409 -989
rect 415 -985 416 -983
rect 415 -991 416 -989
rect 422 -985 423 -983
rect 422 -991 423 -989
rect 429 -985 430 -983
rect 429 -991 430 -989
rect 436 -985 437 -983
rect 436 -991 437 -989
rect 443 -985 444 -983
rect 443 -991 444 -989
rect 450 -985 451 -983
rect 450 -991 451 -989
rect 457 -985 458 -983
rect 457 -991 458 -989
rect 467 -985 468 -983
rect 464 -991 465 -989
rect 471 -985 472 -983
rect 474 -991 475 -989
rect 478 -985 479 -983
rect 478 -991 479 -989
rect 492 -985 493 -983
rect 492 -991 493 -989
rect 506 -985 507 -983
rect 506 -991 507 -989
rect 16 -1032 17 -1030
rect 23 -1032 24 -1030
rect 23 -1038 24 -1036
rect 33 -1038 34 -1036
rect 37 -1032 38 -1030
rect 37 -1038 38 -1036
rect 47 -1032 48 -1030
rect 58 -1032 59 -1030
rect 58 -1038 59 -1036
rect 82 -1032 83 -1030
rect 79 -1038 80 -1036
rect 86 -1032 87 -1030
rect 86 -1038 87 -1036
rect 93 -1032 94 -1030
rect 96 -1038 97 -1036
rect 100 -1038 101 -1036
rect 107 -1032 108 -1030
rect 107 -1038 108 -1036
rect 114 -1032 115 -1030
rect 114 -1038 115 -1036
rect 121 -1032 122 -1030
rect 121 -1038 122 -1036
rect 128 -1032 129 -1030
rect 128 -1038 129 -1036
rect 135 -1038 136 -1036
rect 138 -1038 139 -1036
rect 142 -1032 143 -1030
rect 142 -1038 143 -1036
rect 149 -1032 150 -1030
rect 149 -1038 150 -1036
rect 156 -1032 157 -1030
rect 156 -1038 157 -1036
rect 166 -1032 167 -1030
rect 170 -1032 171 -1030
rect 170 -1038 171 -1036
rect 177 -1032 178 -1030
rect 177 -1038 178 -1036
rect 184 -1038 185 -1036
rect 191 -1032 192 -1030
rect 191 -1038 192 -1036
rect 198 -1032 199 -1030
rect 198 -1038 199 -1036
rect 205 -1032 206 -1030
rect 205 -1038 206 -1036
rect 212 -1032 213 -1030
rect 215 -1032 216 -1030
rect 222 -1032 223 -1030
rect 219 -1038 220 -1036
rect 229 -1032 230 -1030
rect 226 -1038 227 -1036
rect 229 -1038 230 -1036
rect 233 -1032 234 -1030
rect 233 -1038 234 -1036
rect 240 -1032 241 -1030
rect 240 -1038 241 -1036
rect 247 -1032 248 -1030
rect 247 -1038 248 -1036
rect 254 -1032 255 -1030
rect 254 -1038 255 -1036
rect 261 -1032 262 -1030
rect 261 -1038 262 -1036
rect 268 -1032 269 -1030
rect 268 -1038 269 -1036
rect 278 -1032 279 -1030
rect 278 -1038 279 -1036
rect 285 -1032 286 -1030
rect 285 -1038 286 -1036
rect 289 -1032 290 -1030
rect 289 -1038 290 -1036
rect 299 -1038 300 -1036
rect 303 -1038 304 -1036
rect 310 -1032 311 -1030
rect 310 -1038 311 -1036
rect 317 -1032 318 -1030
rect 317 -1038 318 -1036
rect 327 -1032 328 -1030
rect 324 -1038 325 -1036
rect 327 -1038 328 -1036
rect 334 -1032 335 -1030
rect 338 -1032 339 -1030
rect 338 -1038 339 -1036
rect 345 -1032 346 -1030
rect 345 -1038 346 -1036
rect 352 -1032 353 -1030
rect 352 -1038 353 -1036
rect 359 -1032 360 -1030
rect 359 -1038 360 -1036
rect 366 -1032 367 -1030
rect 366 -1038 367 -1036
rect 373 -1032 374 -1030
rect 373 -1038 374 -1036
rect 380 -1032 381 -1030
rect 380 -1038 381 -1036
rect 387 -1032 388 -1030
rect 387 -1038 388 -1036
rect 394 -1032 395 -1030
rect 394 -1038 395 -1036
rect 401 -1032 402 -1030
rect 401 -1038 402 -1036
rect 408 -1032 409 -1030
rect 408 -1038 409 -1036
rect 415 -1032 416 -1030
rect 418 -1032 419 -1030
rect 418 -1038 419 -1036
rect 422 -1038 423 -1036
rect 429 -1032 430 -1030
rect 429 -1038 430 -1036
rect 439 -1032 440 -1030
rect 436 -1038 437 -1036
rect 446 -1032 447 -1030
rect 443 -1038 444 -1036
rect 450 -1032 451 -1030
rect 450 -1038 451 -1036
rect 460 -1032 461 -1030
rect 457 -1038 458 -1036
rect 460 -1038 461 -1036
rect 467 -1032 468 -1030
rect 467 -1038 468 -1036
rect 471 -1032 472 -1030
rect 471 -1038 472 -1036
rect 478 -1032 479 -1030
rect 478 -1038 479 -1036
rect 488 -1032 489 -1030
rect 485 -1038 486 -1036
rect 488 -1038 489 -1036
rect 30 -1077 31 -1075
rect 30 -1083 31 -1081
rect 37 -1077 38 -1075
rect 37 -1083 38 -1081
rect 44 -1083 45 -1081
rect 47 -1083 48 -1081
rect 51 -1077 52 -1075
rect 51 -1083 52 -1081
rect 58 -1083 59 -1081
rect 61 -1083 62 -1081
rect 68 -1077 69 -1075
rect 65 -1083 66 -1081
rect 72 -1077 73 -1075
rect 72 -1083 73 -1081
rect 79 -1077 80 -1075
rect 79 -1083 80 -1081
rect 86 -1077 87 -1075
rect 86 -1083 87 -1081
rect 96 -1077 97 -1075
rect 96 -1083 97 -1081
rect 100 -1077 101 -1075
rect 100 -1083 101 -1081
rect 110 -1077 111 -1075
rect 110 -1083 111 -1081
rect 114 -1077 115 -1075
rect 117 -1077 118 -1075
rect 121 -1077 122 -1075
rect 121 -1083 122 -1081
rect 128 -1077 129 -1075
rect 128 -1083 129 -1081
rect 135 -1077 136 -1075
rect 135 -1083 136 -1081
rect 142 -1077 143 -1075
rect 145 -1083 146 -1081
rect 149 -1077 150 -1075
rect 149 -1083 150 -1081
rect 156 -1077 157 -1075
rect 159 -1077 160 -1075
rect 156 -1083 157 -1081
rect 159 -1083 160 -1081
rect 163 -1077 164 -1075
rect 163 -1083 164 -1081
rect 173 -1077 174 -1075
rect 170 -1083 171 -1081
rect 173 -1083 174 -1081
rect 177 -1077 178 -1075
rect 177 -1083 178 -1081
rect 184 -1077 185 -1075
rect 184 -1083 185 -1081
rect 191 -1077 192 -1075
rect 191 -1083 192 -1081
rect 194 -1083 195 -1081
rect 198 -1077 199 -1075
rect 201 -1083 202 -1081
rect 205 -1077 206 -1075
rect 205 -1083 206 -1081
rect 215 -1077 216 -1075
rect 212 -1083 213 -1081
rect 215 -1083 216 -1081
rect 222 -1077 223 -1075
rect 222 -1083 223 -1081
rect 226 -1083 227 -1081
rect 229 -1083 230 -1081
rect 233 -1077 234 -1075
rect 236 -1083 237 -1081
rect 240 -1077 241 -1075
rect 240 -1083 241 -1081
rect 247 -1077 248 -1075
rect 247 -1083 248 -1081
rect 254 -1077 255 -1075
rect 254 -1083 255 -1081
rect 261 -1077 262 -1075
rect 261 -1083 262 -1081
rect 268 -1077 269 -1075
rect 271 -1083 272 -1081
rect 275 -1077 276 -1075
rect 278 -1077 279 -1075
rect 278 -1083 279 -1081
rect 282 -1077 283 -1075
rect 289 -1077 290 -1075
rect 296 -1077 297 -1075
rect 296 -1083 297 -1081
rect 303 -1077 304 -1075
rect 306 -1077 307 -1075
rect 303 -1083 304 -1081
rect 310 -1077 311 -1075
rect 310 -1083 311 -1081
rect 317 -1077 318 -1075
rect 317 -1083 318 -1081
rect 324 -1077 325 -1075
rect 324 -1083 325 -1081
rect 331 -1077 332 -1075
rect 331 -1083 332 -1081
rect 338 -1077 339 -1075
rect 341 -1077 342 -1075
rect 338 -1083 339 -1081
rect 341 -1083 342 -1081
rect 345 -1077 346 -1075
rect 348 -1077 349 -1075
rect 348 -1083 349 -1081
rect 352 -1077 353 -1075
rect 352 -1083 353 -1081
rect 359 -1077 360 -1075
rect 359 -1083 360 -1081
rect 366 -1077 367 -1075
rect 366 -1083 367 -1081
rect 373 -1077 374 -1075
rect 373 -1083 374 -1081
rect 380 -1077 381 -1075
rect 380 -1083 381 -1081
rect 387 -1077 388 -1075
rect 387 -1083 388 -1081
rect 394 -1077 395 -1075
rect 394 -1083 395 -1081
rect 401 -1077 402 -1075
rect 401 -1083 402 -1081
rect 408 -1077 409 -1075
rect 408 -1083 409 -1081
rect 415 -1077 416 -1075
rect 415 -1083 416 -1081
rect 422 -1077 423 -1075
rect 422 -1083 423 -1081
rect 429 -1077 430 -1075
rect 429 -1083 430 -1081
rect 436 -1077 437 -1075
rect 436 -1083 437 -1081
rect 443 -1077 444 -1075
rect 443 -1083 444 -1081
rect 450 -1077 451 -1075
rect 450 -1083 451 -1081
rect 457 -1077 458 -1075
rect 457 -1083 458 -1081
rect 464 -1077 465 -1075
rect 464 -1083 465 -1081
rect 471 -1083 472 -1081
rect 478 -1083 479 -1081
rect 481 -1083 482 -1081
rect 485 -1077 486 -1075
rect 485 -1083 486 -1081
rect 495 -1077 496 -1075
rect 495 -1083 496 -1081
rect 499 -1077 500 -1075
rect 499 -1083 500 -1081
rect 47 -1116 48 -1114
rect 65 -1110 66 -1108
rect 65 -1116 66 -1114
rect 72 -1110 73 -1108
rect 72 -1116 73 -1114
rect 79 -1110 80 -1108
rect 82 -1110 83 -1108
rect 86 -1110 87 -1108
rect 89 -1110 90 -1108
rect 93 -1116 94 -1114
rect 100 -1110 101 -1108
rect 100 -1116 101 -1114
rect 107 -1110 108 -1108
rect 114 -1110 115 -1108
rect 114 -1116 115 -1114
rect 121 -1110 122 -1108
rect 124 -1110 125 -1108
rect 124 -1116 125 -1114
rect 128 -1110 129 -1108
rect 128 -1116 129 -1114
rect 135 -1110 136 -1108
rect 135 -1116 136 -1114
rect 142 -1116 143 -1114
rect 149 -1110 150 -1108
rect 149 -1116 150 -1114
rect 156 -1110 157 -1108
rect 156 -1116 157 -1114
rect 163 -1110 164 -1108
rect 170 -1110 171 -1108
rect 170 -1116 171 -1114
rect 177 -1110 178 -1108
rect 177 -1116 178 -1114
rect 184 -1110 185 -1108
rect 184 -1116 185 -1114
rect 191 -1116 192 -1114
rect 194 -1116 195 -1114
rect 201 -1116 202 -1114
rect 208 -1110 209 -1108
rect 208 -1116 209 -1114
rect 212 -1110 213 -1108
rect 215 -1110 216 -1108
rect 212 -1116 213 -1114
rect 222 -1110 223 -1108
rect 226 -1110 227 -1108
rect 226 -1116 227 -1114
rect 229 -1116 230 -1114
rect 233 -1110 234 -1108
rect 236 -1110 237 -1108
rect 233 -1116 234 -1114
rect 240 -1110 241 -1108
rect 240 -1116 241 -1114
rect 247 -1110 248 -1108
rect 250 -1116 251 -1114
rect 254 -1110 255 -1108
rect 254 -1116 255 -1114
rect 261 -1110 262 -1108
rect 261 -1116 262 -1114
rect 268 -1110 269 -1108
rect 271 -1110 272 -1108
rect 268 -1116 269 -1114
rect 271 -1116 272 -1114
rect 275 -1110 276 -1108
rect 275 -1116 276 -1114
rect 285 -1116 286 -1114
rect 289 -1110 290 -1108
rect 289 -1116 290 -1114
rect 296 -1110 297 -1108
rect 296 -1116 297 -1114
rect 303 -1110 304 -1108
rect 303 -1116 304 -1114
rect 310 -1110 311 -1108
rect 310 -1116 311 -1114
rect 313 -1116 314 -1114
rect 317 -1110 318 -1108
rect 317 -1116 318 -1114
rect 324 -1110 325 -1108
rect 324 -1116 325 -1114
rect 331 -1110 332 -1108
rect 331 -1116 332 -1114
rect 334 -1116 335 -1114
rect 338 -1110 339 -1108
rect 338 -1116 339 -1114
rect 345 -1110 346 -1108
rect 345 -1116 346 -1114
rect 352 -1116 353 -1114
rect 359 -1110 360 -1108
rect 359 -1116 360 -1114
rect 366 -1110 367 -1108
rect 369 -1110 370 -1108
rect 369 -1116 370 -1114
rect 373 -1110 374 -1108
rect 373 -1116 374 -1114
rect 380 -1110 381 -1108
rect 380 -1116 381 -1114
rect 387 -1110 388 -1108
rect 387 -1116 388 -1114
rect 394 -1110 395 -1108
rect 397 -1116 398 -1114
rect 401 -1110 402 -1108
rect 401 -1116 402 -1114
rect 408 -1116 409 -1114
rect 415 -1110 416 -1108
rect 415 -1116 416 -1114
rect 422 -1110 423 -1108
rect 422 -1116 423 -1114
rect 432 -1110 433 -1108
rect 432 -1116 433 -1114
rect 436 -1110 437 -1108
rect 436 -1116 437 -1114
rect 443 -1110 444 -1108
rect 443 -1116 444 -1114
rect 450 -1116 451 -1114
rect 457 -1110 458 -1108
rect 457 -1116 458 -1114
rect 47 -1149 48 -1147
rect 51 -1143 52 -1141
rect 51 -1149 52 -1147
rect 58 -1149 59 -1147
rect 65 -1143 66 -1141
rect 65 -1149 66 -1147
rect 72 -1143 73 -1141
rect 75 -1143 76 -1141
rect 82 -1143 83 -1141
rect 82 -1149 83 -1147
rect 86 -1149 87 -1147
rect 89 -1149 90 -1147
rect 93 -1143 94 -1141
rect 100 -1143 101 -1141
rect 100 -1149 101 -1147
rect 110 -1143 111 -1141
rect 107 -1149 108 -1147
rect 114 -1143 115 -1141
rect 114 -1149 115 -1147
rect 121 -1143 122 -1141
rect 121 -1149 122 -1147
rect 128 -1149 129 -1147
rect 135 -1149 136 -1147
rect 142 -1143 143 -1141
rect 142 -1149 143 -1147
rect 149 -1143 150 -1141
rect 149 -1149 150 -1147
rect 156 -1143 157 -1141
rect 156 -1149 157 -1147
rect 163 -1143 164 -1141
rect 163 -1149 164 -1147
rect 170 -1143 171 -1141
rect 170 -1149 171 -1147
rect 177 -1143 178 -1141
rect 177 -1149 178 -1147
rect 184 -1149 185 -1147
rect 187 -1149 188 -1147
rect 191 -1143 192 -1141
rect 194 -1143 195 -1141
rect 198 -1143 199 -1141
rect 198 -1149 199 -1147
rect 205 -1143 206 -1141
rect 208 -1149 209 -1147
rect 212 -1149 213 -1147
rect 215 -1149 216 -1147
rect 222 -1143 223 -1141
rect 222 -1149 223 -1147
rect 226 -1143 227 -1141
rect 229 -1143 230 -1141
rect 226 -1149 227 -1147
rect 229 -1149 230 -1147
rect 233 -1143 234 -1141
rect 233 -1149 234 -1147
rect 240 -1143 241 -1141
rect 243 -1143 244 -1141
rect 240 -1149 241 -1147
rect 243 -1149 244 -1147
rect 247 -1143 248 -1141
rect 247 -1149 248 -1147
rect 254 -1143 255 -1141
rect 257 -1143 258 -1141
rect 257 -1149 258 -1147
rect 261 -1143 262 -1141
rect 261 -1149 262 -1147
rect 268 -1143 269 -1141
rect 268 -1149 269 -1147
rect 271 -1149 272 -1147
rect 275 -1143 276 -1141
rect 275 -1149 276 -1147
rect 282 -1143 283 -1141
rect 282 -1149 283 -1147
rect 289 -1143 290 -1141
rect 289 -1149 290 -1147
rect 296 -1143 297 -1141
rect 296 -1149 297 -1147
rect 303 -1143 304 -1141
rect 306 -1143 307 -1141
rect 306 -1149 307 -1147
rect 310 -1143 311 -1141
rect 310 -1149 311 -1147
rect 313 -1149 314 -1147
rect 317 -1143 318 -1141
rect 317 -1149 318 -1147
rect 324 -1143 325 -1141
rect 324 -1149 325 -1147
rect 331 -1143 332 -1141
rect 331 -1149 332 -1147
rect 338 -1143 339 -1141
rect 338 -1149 339 -1147
rect 345 -1143 346 -1141
rect 345 -1149 346 -1147
rect 352 -1143 353 -1141
rect 352 -1149 353 -1147
rect 359 -1143 360 -1141
rect 359 -1149 360 -1147
rect 366 -1143 367 -1141
rect 366 -1149 367 -1147
rect 373 -1143 374 -1141
rect 373 -1149 374 -1147
rect 383 -1143 384 -1141
rect 387 -1143 388 -1141
rect 394 -1143 395 -1141
rect 394 -1149 395 -1147
rect 401 -1143 402 -1141
rect 404 -1143 405 -1141
rect 401 -1149 402 -1147
rect 404 -1149 405 -1147
rect 408 -1143 409 -1141
rect 408 -1149 409 -1147
rect 415 -1143 416 -1141
rect 415 -1149 416 -1147
rect 422 -1143 423 -1141
rect 422 -1149 423 -1147
rect 446 -1149 447 -1147
rect 450 -1143 451 -1141
rect 450 -1149 451 -1147
rect 47 -1186 48 -1184
rect 51 -1180 52 -1178
rect 51 -1186 52 -1184
rect 61 -1180 62 -1178
rect 65 -1180 66 -1178
rect 75 -1186 76 -1184
rect 79 -1186 80 -1184
rect 89 -1186 90 -1184
rect 93 -1186 94 -1184
rect 100 -1180 101 -1178
rect 100 -1186 101 -1184
rect 107 -1180 108 -1178
rect 107 -1186 108 -1184
rect 117 -1180 118 -1178
rect 121 -1180 122 -1178
rect 121 -1186 122 -1184
rect 128 -1180 129 -1178
rect 128 -1186 129 -1184
rect 135 -1180 136 -1178
rect 135 -1186 136 -1184
rect 145 -1180 146 -1178
rect 142 -1186 143 -1184
rect 149 -1186 150 -1184
rect 152 -1186 153 -1184
rect 156 -1180 157 -1178
rect 156 -1186 157 -1184
rect 166 -1186 167 -1184
rect 173 -1186 174 -1184
rect 177 -1186 178 -1184
rect 184 -1180 185 -1178
rect 184 -1186 185 -1184
rect 191 -1180 192 -1178
rect 194 -1180 195 -1178
rect 191 -1186 192 -1184
rect 201 -1186 202 -1184
rect 205 -1180 206 -1178
rect 205 -1186 206 -1184
rect 212 -1180 213 -1178
rect 212 -1186 213 -1184
rect 222 -1186 223 -1184
rect 226 -1180 227 -1178
rect 226 -1186 227 -1184
rect 229 -1186 230 -1184
rect 233 -1180 234 -1178
rect 236 -1180 237 -1178
rect 236 -1186 237 -1184
rect 243 -1180 244 -1178
rect 240 -1186 241 -1184
rect 247 -1180 248 -1178
rect 254 -1180 255 -1178
rect 261 -1180 262 -1178
rect 261 -1186 262 -1184
rect 268 -1180 269 -1178
rect 268 -1186 269 -1184
rect 275 -1180 276 -1178
rect 275 -1186 276 -1184
rect 282 -1180 283 -1178
rect 282 -1186 283 -1184
rect 289 -1186 290 -1184
rect 292 -1186 293 -1184
rect 296 -1180 297 -1178
rect 299 -1180 300 -1178
rect 303 -1180 304 -1178
rect 303 -1186 304 -1184
rect 310 -1180 311 -1178
rect 310 -1186 311 -1184
rect 317 -1180 318 -1178
rect 317 -1186 318 -1184
rect 324 -1180 325 -1178
rect 324 -1186 325 -1184
rect 331 -1180 332 -1178
rect 331 -1186 332 -1184
rect 338 -1180 339 -1178
rect 338 -1186 339 -1184
rect 345 -1186 346 -1184
rect 348 -1186 349 -1184
rect 352 -1180 353 -1178
rect 352 -1186 353 -1184
rect 359 -1180 360 -1178
rect 359 -1186 360 -1184
rect 366 -1180 367 -1178
rect 366 -1186 367 -1184
rect 373 -1180 374 -1178
rect 373 -1186 374 -1184
rect 380 -1180 381 -1178
rect 380 -1186 381 -1184
rect 387 -1180 388 -1178
rect 387 -1186 388 -1184
rect 394 -1180 395 -1178
rect 394 -1186 395 -1184
rect 401 -1180 402 -1178
rect 401 -1186 402 -1184
rect 415 -1180 416 -1178
rect 418 -1180 419 -1178
rect 415 -1186 416 -1184
rect 422 -1180 423 -1178
rect 422 -1186 423 -1184
rect 429 -1180 430 -1178
rect 429 -1186 430 -1184
rect 47 -1207 48 -1205
rect 65 -1207 66 -1205
rect 68 -1207 69 -1205
rect 72 -1207 73 -1205
rect 72 -1213 73 -1211
rect 79 -1207 80 -1205
rect 82 -1207 83 -1205
rect 79 -1213 80 -1211
rect 89 -1213 90 -1211
rect 96 -1207 97 -1205
rect 100 -1207 101 -1205
rect 100 -1213 101 -1211
rect 107 -1207 108 -1205
rect 107 -1213 108 -1211
rect 114 -1207 115 -1205
rect 114 -1213 115 -1211
rect 121 -1207 122 -1205
rect 121 -1213 122 -1211
rect 128 -1207 129 -1205
rect 128 -1213 129 -1211
rect 135 -1207 136 -1205
rect 138 -1207 139 -1205
rect 135 -1213 136 -1211
rect 138 -1213 139 -1211
rect 145 -1207 146 -1205
rect 142 -1213 143 -1211
rect 149 -1207 150 -1205
rect 152 -1213 153 -1211
rect 156 -1207 157 -1205
rect 159 -1207 160 -1205
rect 156 -1213 157 -1211
rect 159 -1213 160 -1211
rect 166 -1207 167 -1205
rect 163 -1213 164 -1211
rect 170 -1207 171 -1205
rect 170 -1213 171 -1211
rect 177 -1207 178 -1205
rect 177 -1213 178 -1211
rect 184 -1207 185 -1205
rect 187 -1213 188 -1211
rect 194 -1213 195 -1211
rect 198 -1207 199 -1205
rect 198 -1213 199 -1211
rect 205 -1207 206 -1205
rect 205 -1213 206 -1211
rect 212 -1207 213 -1205
rect 212 -1213 213 -1211
rect 219 -1207 220 -1205
rect 222 -1207 223 -1205
rect 222 -1213 223 -1211
rect 226 -1207 227 -1205
rect 229 -1207 230 -1205
rect 229 -1213 230 -1211
rect 233 -1207 234 -1205
rect 233 -1213 234 -1211
rect 240 -1207 241 -1205
rect 243 -1213 244 -1211
rect 247 -1207 248 -1205
rect 247 -1213 248 -1211
rect 254 -1207 255 -1205
rect 254 -1213 255 -1211
rect 282 -1207 283 -1205
rect 282 -1213 283 -1211
rect 289 -1207 290 -1205
rect 292 -1207 293 -1205
rect 292 -1213 293 -1211
rect 296 -1207 297 -1205
rect 296 -1213 297 -1211
rect 303 -1207 304 -1205
rect 303 -1213 304 -1211
rect 306 -1213 307 -1211
rect 310 -1213 311 -1211
rect 313 -1213 314 -1211
rect 317 -1207 318 -1205
rect 317 -1213 318 -1211
rect 324 -1207 325 -1205
rect 324 -1213 325 -1211
rect 331 -1207 332 -1205
rect 331 -1213 332 -1211
rect 341 -1207 342 -1205
rect 341 -1213 342 -1211
rect 345 -1207 346 -1205
rect 345 -1213 346 -1211
rect 352 -1213 353 -1211
rect 359 -1207 360 -1205
rect 359 -1213 360 -1211
rect 366 -1207 367 -1205
rect 366 -1213 367 -1211
rect 373 -1213 374 -1211
rect 380 -1207 381 -1205
rect 380 -1213 381 -1211
rect 408 -1207 409 -1205
rect 408 -1213 409 -1211
rect 422 -1207 423 -1205
rect 425 -1213 426 -1211
rect 429 -1207 430 -1205
rect 429 -1213 430 -1211
rect 23 -1236 24 -1234
rect 33 -1230 34 -1228
rect 37 -1230 38 -1228
rect 37 -1236 38 -1234
rect 44 -1230 45 -1228
rect 51 -1230 52 -1228
rect 51 -1236 52 -1234
rect 58 -1230 59 -1228
rect 58 -1236 59 -1234
rect 65 -1230 66 -1228
rect 65 -1236 66 -1234
rect 72 -1230 73 -1228
rect 79 -1230 80 -1228
rect 79 -1236 80 -1234
rect 93 -1230 94 -1228
rect 93 -1236 94 -1234
rect 100 -1230 101 -1228
rect 100 -1236 101 -1234
rect 110 -1236 111 -1234
rect 114 -1236 115 -1234
rect 117 -1236 118 -1234
rect 121 -1230 122 -1228
rect 124 -1230 125 -1228
rect 128 -1230 129 -1228
rect 128 -1236 129 -1234
rect 138 -1236 139 -1234
rect 142 -1230 143 -1228
rect 142 -1236 143 -1234
rect 149 -1230 150 -1228
rect 149 -1236 150 -1234
rect 159 -1236 160 -1234
rect 163 -1230 164 -1228
rect 163 -1236 164 -1234
rect 173 -1230 174 -1228
rect 170 -1236 171 -1234
rect 180 -1230 181 -1228
rect 184 -1230 185 -1228
rect 184 -1236 185 -1234
rect 191 -1230 192 -1228
rect 191 -1236 192 -1234
rect 201 -1230 202 -1228
rect 205 -1236 206 -1234
rect 208 -1236 209 -1234
rect 212 -1230 213 -1228
rect 215 -1230 216 -1228
rect 215 -1236 216 -1234
rect 219 -1230 220 -1228
rect 222 -1230 223 -1228
rect 222 -1236 223 -1234
rect 229 -1230 230 -1228
rect 233 -1230 234 -1228
rect 233 -1236 234 -1234
rect 240 -1230 241 -1228
rect 240 -1236 241 -1234
rect 250 -1236 251 -1234
rect 254 -1230 255 -1228
rect 254 -1236 255 -1234
rect 261 -1236 262 -1234
rect 268 -1230 269 -1228
rect 268 -1236 269 -1234
rect 275 -1230 276 -1228
rect 275 -1236 276 -1234
rect 282 -1230 283 -1228
rect 282 -1236 283 -1234
rect 292 -1230 293 -1228
rect 299 -1236 300 -1234
rect 303 -1230 304 -1228
rect 303 -1236 304 -1234
rect 310 -1230 311 -1228
rect 310 -1236 311 -1234
rect 317 -1230 318 -1228
rect 320 -1230 321 -1228
rect 327 -1236 328 -1234
rect 338 -1230 339 -1228
rect 338 -1236 339 -1234
rect 345 -1230 346 -1228
rect 352 -1230 353 -1228
rect 352 -1236 353 -1234
rect 359 -1230 360 -1228
rect 359 -1236 360 -1234
rect 366 -1230 367 -1228
rect 373 -1230 374 -1228
rect 373 -1236 374 -1234
rect 401 -1230 402 -1228
rect 401 -1236 402 -1234
rect 408 -1236 409 -1234
rect 415 -1236 416 -1234
rect 422 -1230 423 -1228
rect 422 -1236 423 -1234
rect 432 -1230 433 -1228
rect 23 -1255 24 -1253
rect 30 -1255 31 -1253
rect 30 -1261 31 -1259
rect 37 -1261 38 -1259
rect 44 -1255 45 -1253
rect 58 -1255 59 -1253
rect 58 -1261 59 -1259
rect 68 -1261 69 -1259
rect 75 -1255 76 -1253
rect 72 -1261 73 -1259
rect 79 -1255 80 -1253
rect 79 -1261 80 -1259
rect 103 -1255 104 -1253
rect 107 -1261 108 -1259
rect 114 -1255 115 -1253
rect 114 -1261 115 -1259
rect 121 -1255 122 -1253
rect 121 -1261 122 -1259
rect 128 -1255 129 -1253
rect 128 -1261 129 -1259
rect 138 -1261 139 -1259
rect 145 -1255 146 -1253
rect 142 -1261 143 -1259
rect 152 -1255 153 -1253
rect 152 -1261 153 -1259
rect 159 -1255 160 -1253
rect 163 -1261 164 -1259
rect 170 -1255 171 -1253
rect 170 -1261 171 -1259
rect 177 -1255 178 -1253
rect 177 -1261 178 -1259
rect 187 -1261 188 -1259
rect 194 -1255 195 -1253
rect 198 -1261 199 -1259
rect 208 -1255 209 -1253
rect 205 -1261 206 -1259
rect 208 -1261 209 -1259
rect 212 -1255 213 -1253
rect 212 -1261 213 -1259
rect 219 -1255 220 -1253
rect 222 -1255 223 -1253
rect 226 -1255 227 -1253
rect 226 -1261 227 -1259
rect 233 -1255 234 -1253
rect 233 -1261 234 -1259
rect 240 -1255 241 -1253
rect 250 -1261 251 -1259
rect 257 -1255 258 -1253
rect 261 -1255 262 -1253
rect 261 -1261 262 -1259
rect 268 -1255 269 -1253
rect 268 -1261 269 -1259
rect 278 -1255 279 -1253
rect 285 -1261 286 -1259
rect 289 -1255 290 -1253
rect 289 -1261 290 -1259
rect 296 -1261 297 -1259
rect 303 -1255 304 -1253
rect 303 -1261 304 -1259
rect 317 -1261 318 -1259
rect 324 -1255 325 -1253
rect 324 -1261 325 -1259
rect 334 -1255 335 -1253
rect 338 -1255 339 -1253
rect 338 -1261 339 -1259
rect 348 -1261 349 -1259
rect 355 -1261 356 -1259
rect 359 -1255 360 -1253
rect 359 -1261 360 -1259
rect 369 -1255 370 -1253
<< metal1 >>
rect 138 0 150 1
rect 177 0 192 1
rect 198 0 216 1
rect 226 0 241 1
rect 187 -2 206 -1
rect 212 -2 220 -1
rect 135 -13 185 -12
rect 187 -13 230 -12
rect 240 -13 248 -12
rect 324 -13 332 -12
rect 145 -15 150 -14
rect 163 -15 171 -14
rect 177 -15 185 -14
rect 191 -15 234 -14
rect 156 -17 178 -16
rect 198 -17 206 -16
rect 208 -17 220 -16
rect 226 -17 255 -16
rect 198 -19 216 -18
rect 219 -19 241 -18
rect 229 -21 237 -20
rect 128 -32 146 -31
rect 198 -32 220 -31
rect 222 -32 262 -31
rect 268 -32 290 -31
rect 296 -32 304 -31
rect 324 -32 332 -31
rect 135 -34 153 -33
rect 198 -34 248 -33
rect 327 -34 332 -33
rect 135 -36 153 -35
rect 201 -36 234 -35
rect 142 -38 160 -37
rect 173 -38 234 -37
rect 159 -40 178 -39
rect 205 -40 227 -39
rect 163 -42 178 -41
rect 205 -42 241 -41
rect 163 -44 185 -43
rect 208 -44 213 -43
rect 226 -44 283 -43
rect 229 -46 241 -45
rect 191 -48 230 -47
rect 103 -59 108 -58
rect 121 -59 136 -58
rect 142 -59 164 -58
rect 205 -59 213 -58
rect 226 -59 248 -58
rect 261 -59 314 -58
rect 128 -61 160 -60
rect 191 -61 262 -60
rect 268 -61 283 -60
rect 289 -61 307 -60
rect 142 -63 150 -62
rect 184 -63 192 -62
rect 229 -63 234 -62
rect 240 -63 255 -62
rect 275 -63 279 -62
rect 282 -63 300 -62
rect 177 -65 185 -64
rect 201 -65 241 -64
rect 296 -65 304 -64
rect 219 -67 255 -66
rect 292 -67 297 -66
rect 170 -69 220 -68
rect 166 -71 171 -70
rect 100 -82 108 -81
rect 114 -82 132 -81
rect 138 -82 150 -81
rect 159 -82 164 -81
rect 166 -82 178 -81
rect 184 -82 195 -81
rect 205 -82 213 -81
rect 229 -82 255 -81
rect 275 -82 304 -81
rect 317 -82 325 -81
rect 107 -84 129 -83
rect 149 -84 171 -83
rect 191 -84 199 -83
rect 222 -84 230 -83
rect 233 -84 248 -83
rect 282 -84 293 -83
rect 296 -84 311 -83
rect 317 -84 321 -83
rect 324 -84 332 -83
rect 121 -86 146 -85
rect 198 -86 216 -85
rect 219 -86 248 -85
rect 117 -88 122 -87
rect 128 -88 136 -87
rect 142 -88 146 -87
rect 222 -88 297 -87
rect 226 -90 255 -89
rect 236 -92 262 -91
rect 240 -94 276 -93
rect 261 -96 272 -95
rect 86 -107 104 -106
rect 107 -107 129 -106
rect 135 -107 146 -106
rect 149 -107 181 -106
rect 198 -107 220 -106
rect 229 -107 276 -106
rect 282 -107 297 -106
rect 380 -107 384 -106
rect 114 -109 125 -108
rect 135 -109 164 -108
rect 198 -109 213 -108
rect 215 -109 234 -108
rect 243 -109 304 -108
rect 103 -111 115 -110
rect 156 -111 185 -110
rect 205 -111 237 -110
rect 247 -111 272 -110
rect 289 -111 311 -110
rect 107 -113 125 -112
rect 163 -113 171 -112
rect 177 -113 216 -112
rect 268 -113 318 -112
rect 180 -115 206 -114
rect 208 -115 220 -114
rect 261 -115 269 -114
rect 303 -115 325 -114
rect 184 -117 192 -116
rect 212 -117 300 -116
rect 310 -117 318 -116
rect 254 -119 262 -118
rect 226 -121 255 -120
rect 79 -132 83 -131
rect 107 -132 143 -131
rect 156 -132 195 -131
rect 219 -132 234 -131
rect 257 -132 262 -131
rect 268 -132 272 -131
rect 296 -132 304 -131
rect 310 -132 318 -131
rect 380 -132 388 -131
rect 79 -134 87 -133
rect 107 -134 118 -133
rect 131 -134 139 -133
rect 159 -134 216 -133
rect 226 -134 269 -133
rect 275 -134 318 -133
rect 114 -136 122 -135
rect 128 -136 132 -135
rect 135 -136 153 -135
rect 163 -136 178 -135
rect 184 -136 230 -135
rect 254 -136 262 -135
rect 299 -136 325 -135
rect 128 -138 157 -137
rect 170 -138 255 -137
rect 145 -140 164 -139
rect 173 -140 178 -139
rect 191 -140 216 -139
rect 121 -142 174 -141
rect 205 -142 220 -141
rect 152 -144 209 -143
rect 205 -146 241 -145
rect 107 -157 153 -156
rect 156 -157 164 -156
rect 173 -157 178 -156
rect 187 -157 192 -156
rect 198 -157 227 -156
rect 233 -157 248 -156
rect 254 -157 304 -156
rect 317 -157 342 -156
rect 359 -157 374 -156
rect 387 -157 395 -156
rect 408 -157 416 -156
rect 436 -157 444 -156
rect 114 -159 118 -158
rect 121 -159 136 -158
rect 152 -159 185 -158
rect 212 -159 255 -158
rect 261 -159 272 -158
rect 296 -159 314 -158
rect 317 -159 325 -158
rect 331 -159 353 -158
rect 362 -159 381 -158
rect 383 -159 388 -158
rect 124 -161 139 -160
rect 163 -161 202 -160
rect 205 -161 213 -160
rect 215 -161 220 -160
rect 226 -161 367 -160
rect 135 -163 146 -162
rect 170 -163 192 -162
rect 205 -163 216 -162
rect 219 -163 230 -162
rect 233 -163 290 -162
rect 320 -163 346 -162
rect 177 -165 244 -164
rect 261 -165 276 -164
rect 278 -165 325 -164
rect 240 -167 283 -166
rect 268 -169 384 -168
rect 75 -180 80 -179
rect 86 -180 122 -179
rect 135 -180 143 -179
rect 149 -180 199 -179
rect 229 -180 248 -179
rect 250 -180 360 -179
rect 369 -180 388 -179
rect 415 -180 423 -179
rect 432 -180 444 -179
rect 89 -182 94 -181
rect 107 -182 129 -181
rect 156 -182 160 -181
rect 163 -182 269 -181
rect 271 -182 325 -181
rect 338 -182 374 -181
rect 383 -182 395 -181
rect 401 -182 416 -181
rect 436 -182 444 -181
rect 121 -184 136 -183
rect 170 -184 213 -183
rect 233 -184 262 -183
rect 296 -184 314 -183
rect 317 -184 356 -183
rect 380 -184 395 -183
rect 170 -186 220 -185
rect 229 -186 234 -185
rect 254 -186 276 -185
rect 303 -186 311 -185
rect 317 -186 332 -185
rect 345 -186 374 -185
rect 177 -188 216 -187
rect 219 -188 276 -187
rect 285 -188 346 -187
rect 177 -190 185 -189
rect 191 -190 206 -189
rect 254 -190 283 -189
rect 285 -190 353 -189
rect 163 -192 206 -191
rect 261 -192 325 -191
rect 331 -192 367 -191
rect 184 -194 241 -193
rect 296 -194 304 -193
rect 201 -196 241 -195
rect 72 -207 97 -206
rect 100 -207 122 -206
rect 128 -207 227 -206
rect 261 -207 332 -206
rect 345 -207 388 -206
rect 394 -207 402 -206
rect 404 -207 409 -206
rect 415 -207 423 -206
rect 436 -207 440 -206
rect 79 -209 87 -208
rect 103 -209 108 -208
rect 121 -209 248 -208
rect 268 -209 304 -208
rect 306 -209 318 -208
rect 373 -209 384 -208
rect 79 -211 146 -210
rect 149 -211 230 -210
rect 236 -211 346 -210
rect 373 -211 381 -210
rect 86 -213 188 -212
rect 191 -213 220 -212
rect 222 -213 241 -212
rect 257 -213 269 -212
rect 275 -213 318 -212
rect 359 -213 381 -212
rect 93 -215 150 -214
rect 156 -215 181 -214
rect 198 -215 248 -214
rect 310 -215 332 -214
rect 107 -217 220 -216
rect 229 -217 339 -216
rect 142 -219 164 -218
rect 170 -219 265 -218
rect 296 -219 311 -218
rect 324 -219 339 -218
rect 159 -221 192 -220
rect 201 -221 276 -220
rect 324 -221 353 -220
rect 170 -223 178 -222
rect 205 -223 255 -222
rect 352 -223 370 -222
rect 131 -225 178 -224
rect 184 -225 206 -224
rect 212 -225 297 -224
rect 212 -227 234 -226
rect 240 -227 360 -226
rect 233 -229 283 -228
rect 68 -240 157 -239
rect 170 -240 188 -239
rect 229 -240 318 -239
rect 359 -240 444 -239
rect 450 -240 458 -239
rect 530 -240 535 -239
rect 86 -242 160 -241
rect 170 -242 206 -241
rect 240 -242 276 -241
rect 292 -242 360 -241
rect 366 -242 454 -241
rect 79 -244 206 -243
rect 243 -244 304 -243
rect 331 -244 367 -243
rect 369 -244 388 -243
rect 394 -244 440 -243
rect 72 -246 80 -245
rect 93 -246 185 -245
rect 194 -246 241 -245
rect 250 -246 346 -245
rect 418 -246 423 -245
rect 93 -248 213 -247
rect 254 -248 265 -247
rect 271 -248 339 -247
rect 345 -248 353 -247
rect 373 -248 423 -247
rect 100 -250 136 -249
rect 138 -250 188 -249
rect 208 -250 374 -249
rect 408 -250 419 -249
rect 107 -252 167 -251
rect 177 -252 192 -251
rect 212 -252 248 -251
rect 254 -252 381 -251
rect 107 -254 115 -253
rect 121 -254 227 -253
rect 257 -254 318 -253
rect 338 -254 416 -253
rect 114 -256 146 -255
rect 180 -256 234 -255
rect 261 -256 325 -255
rect 121 -258 150 -257
rect 198 -258 227 -257
rect 261 -258 269 -257
rect 275 -258 300 -257
rect 303 -258 388 -257
rect 128 -260 164 -259
rect 268 -260 332 -259
rect 131 -262 216 -261
rect 296 -262 430 -261
rect 135 -264 157 -263
rect 296 -264 402 -263
rect 142 -266 153 -265
rect 310 -266 353 -265
rect 86 -268 153 -267
rect 219 -268 311 -267
rect 149 -270 283 -269
rect 282 -272 290 -271
rect 30 -283 38 -282
rect 47 -283 150 -282
rect 177 -283 213 -282
rect 222 -283 262 -282
rect 268 -283 402 -282
rect 415 -283 437 -282
rect 453 -283 458 -282
rect 527 -283 535 -282
rect 30 -285 34 -284
rect 51 -285 55 -284
rect 58 -285 132 -284
rect 135 -285 164 -284
rect 184 -285 220 -284
rect 243 -285 451 -284
rect 68 -287 185 -286
rect 194 -287 395 -286
rect 401 -287 423 -286
rect 75 -289 80 -288
rect 82 -289 192 -288
rect 205 -289 220 -288
rect 247 -289 290 -288
rect 292 -289 367 -288
rect 387 -289 423 -288
rect 86 -291 104 -290
rect 107 -291 122 -290
rect 149 -291 171 -290
rect 208 -291 241 -290
rect 254 -291 353 -290
rect 380 -291 388 -290
rect 394 -291 409 -290
rect 93 -293 262 -292
rect 268 -293 276 -292
rect 282 -293 304 -292
rect 306 -293 311 -292
rect 338 -293 367 -292
rect 408 -293 419 -292
rect 93 -295 115 -294
rect 121 -295 146 -294
rect 156 -295 178 -294
rect 226 -295 276 -294
rect 296 -295 430 -294
rect 100 -297 153 -296
rect 163 -297 325 -296
rect 352 -297 377 -296
rect 114 -299 199 -298
rect 226 -299 248 -298
rect 299 -299 444 -298
rect 128 -301 283 -300
rect 310 -301 318 -300
rect 142 -303 297 -302
rect 317 -303 346 -302
rect 170 -305 339 -304
rect 198 -307 234 -306
rect 331 -307 346 -306
rect 187 -309 234 -308
rect 331 -309 360 -308
rect 229 -311 381 -310
rect 359 -313 374 -312
rect 19 -324 24 -323
rect 37 -324 94 -323
rect 96 -324 167 -323
rect 194 -324 276 -323
rect 282 -324 367 -323
rect 373 -324 472 -323
rect 513 -324 521 -323
rect 523 -324 528 -323
rect 51 -326 202 -325
rect 219 -326 297 -325
rect 327 -326 332 -325
rect 408 -326 416 -325
rect 422 -326 458 -325
rect 58 -328 108 -327
rect 110 -328 139 -327
rect 145 -328 157 -327
rect 159 -328 178 -327
rect 198 -328 244 -327
rect 247 -328 318 -327
rect 331 -328 381 -327
rect 390 -328 409 -327
rect 436 -328 468 -327
rect 58 -330 87 -329
rect 100 -330 150 -329
rect 177 -330 185 -329
rect 198 -330 381 -329
rect 387 -330 437 -329
rect 65 -332 136 -331
rect 149 -332 171 -331
rect 184 -332 251 -331
rect 254 -332 367 -331
rect 401 -332 423 -331
rect 82 -334 143 -333
rect 212 -334 220 -333
rect 243 -334 339 -333
rect 72 -336 83 -335
rect 86 -336 122 -335
rect 124 -336 216 -335
rect 250 -336 304 -335
rect 100 -338 108 -337
rect 110 -338 153 -337
rect 163 -338 213 -337
rect 261 -338 311 -337
rect 114 -340 227 -339
rect 264 -340 374 -339
rect 44 -342 115 -341
rect 117 -342 206 -341
rect 264 -342 444 -341
rect 128 -344 230 -343
rect 268 -344 272 -343
rect 285 -344 290 -343
rect 299 -344 402 -343
rect 131 -346 136 -345
rect 194 -346 339 -345
rect 233 -348 286 -347
rect 289 -348 307 -347
rect 310 -348 360 -347
rect 170 -350 234 -349
rect 352 -350 360 -349
rect 345 -352 353 -351
rect 345 -354 430 -353
rect 394 -356 430 -355
rect 240 -358 395 -357
rect 240 -360 451 -359
rect 23 -371 101 -370
rect 121 -371 153 -370
rect 198 -371 272 -370
rect 275 -371 437 -370
rect 443 -371 528 -370
rect 30 -373 118 -372
rect 135 -373 167 -372
rect 226 -373 304 -372
rect 317 -373 367 -372
rect 387 -373 458 -372
rect 481 -373 500 -372
rect 30 -375 174 -374
rect 226 -375 311 -374
rect 331 -375 458 -374
rect 37 -377 115 -376
rect 128 -377 167 -376
rect 233 -377 279 -376
rect 282 -377 465 -376
rect 44 -379 125 -378
rect 138 -379 171 -378
rect 233 -379 314 -378
rect 338 -379 388 -378
rect 390 -379 416 -378
rect 418 -379 521 -378
rect 44 -381 104 -380
rect 149 -381 216 -380
rect 240 -381 297 -380
rect 310 -381 402 -380
rect 415 -381 444 -380
rect 450 -381 493 -380
rect 51 -383 101 -382
rect 243 -383 346 -382
rect 348 -383 367 -382
rect 394 -383 507 -382
rect 58 -385 111 -384
rect 254 -385 283 -384
rect 296 -385 321 -384
rect 352 -385 402 -384
rect 408 -385 451 -384
rect 58 -387 160 -386
rect 254 -387 290 -386
rect 352 -387 472 -386
rect 65 -389 192 -388
rect 250 -389 472 -388
rect 65 -391 83 -390
rect 86 -391 209 -390
rect 261 -391 381 -390
rect 408 -391 423 -390
rect 72 -393 94 -392
rect 110 -393 248 -392
rect 261 -393 395 -392
rect 72 -395 213 -394
rect 268 -395 430 -394
rect 79 -397 108 -396
rect 131 -397 290 -396
rect 324 -397 423 -396
rect 37 -399 108 -398
rect 114 -399 325 -398
rect 359 -399 381 -398
rect 89 -401 143 -400
rect 156 -401 192 -400
rect 212 -401 332 -400
rect 373 -401 430 -400
rect 93 -403 185 -402
rect 229 -403 360 -402
rect 156 -405 437 -404
rect 177 -407 248 -406
rect 275 -407 328 -406
rect 177 -409 195 -408
rect 240 -409 269 -408
rect 317 -409 374 -408
rect 184 -411 206 -410
rect 16 -422 80 -421
rect 86 -422 90 -421
rect 93 -422 216 -421
rect 247 -422 265 -421
rect 268 -422 283 -421
rect 289 -422 293 -421
rect 324 -422 500 -421
rect 520 -422 549 -421
rect 30 -424 146 -423
rect 159 -424 458 -423
rect 464 -424 542 -423
rect 30 -426 111 -425
rect 114 -426 213 -425
rect 219 -426 248 -425
rect 254 -426 325 -425
rect 327 -426 409 -425
rect 415 -426 577 -425
rect 44 -428 223 -427
rect 240 -428 255 -427
rect 261 -428 493 -427
rect 527 -428 563 -427
rect 2 -430 241 -429
rect 278 -430 297 -429
rect 338 -430 486 -429
rect 51 -432 55 -431
rect 58 -432 122 -431
rect 128 -432 202 -431
rect 219 -432 500 -431
rect 37 -434 122 -433
rect 135 -434 167 -433
rect 173 -434 465 -433
rect 471 -434 479 -433
rect 65 -436 199 -435
rect 226 -436 528 -435
rect 72 -438 321 -437
rect 341 -438 402 -437
rect 429 -438 521 -437
rect 72 -440 171 -439
rect 191 -440 276 -439
rect 285 -440 472 -439
rect 9 -442 171 -441
rect 177 -442 286 -441
rect 289 -442 304 -441
rect 348 -442 486 -441
rect 79 -444 346 -443
rect 352 -444 409 -443
rect 436 -444 535 -443
rect 86 -446 185 -445
rect 198 -446 230 -445
rect 296 -446 314 -445
rect 359 -446 458 -445
rect 96 -448 101 -447
rect 107 -448 143 -447
rect 177 -448 244 -447
rect 366 -448 402 -447
rect 436 -448 444 -447
rect 142 -450 360 -449
rect 380 -450 430 -449
rect 443 -450 507 -449
rect 23 -452 507 -451
rect 205 -454 353 -453
rect 373 -454 381 -453
rect 387 -454 493 -453
rect 229 -456 416 -455
rect 275 -458 388 -457
rect 394 -458 398 -457
rect 394 -460 423 -459
rect 397 -462 423 -461
rect 9 -473 122 -472
rect 131 -473 192 -472
rect 219 -473 248 -472
rect 275 -473 472 -472
rect 555 -473 563 -472
rect 16 -475 118 -474
rect 152 -475 178 -474
rect 184 -475 314 -474
rect 355 -475 535 -474
rect 558 -475 563 -474
rect 16 -477 94 -476
rect 107 -477 279 -476
rect 282 -477 472 -476
rect 23 -479 150 -478
rect 159 -479 423 -478
rect 425 -479 486 -478
rect 30 -481 55 -480
rect 58 -481 97 -480
rect 107 -481 234 -480
rect 240 -481 339 -480
rect 359 -481 542 -480
rect 37 -483 241 -482
rect 285 -483 409 -482
rect 464 -483 573 -482
rect 2 -485 286 -484
rect 299 -485 360 -484
rect 373 -485 458 -484
rect 541 -485 549 -484
rect 37 -487 115 -486
rect 142 -487 150 -486
rect 163 -487 507 -486
rect 44 -489 125 -488
rect 135 -489 164 -488
rect 170 -489 178 -488
rect 184 -489 269 -488
rect 303 -489 318 -488
rect 331 -489 339 -488
rect 394 -489 486 -488
rect 51 -491 346 -490
rect 380 -491 395 -490
rect 408 -491 416 -490
rect 436 -491 465 -490
rect 72 -493 230 -492
rect 233 -493 370 -492
rect 380 -493 402 -492
rect 457 -493 500 -492
rect 44 -495 230 -494
rect 289 -495 304 -494
rect 310 -495 528 -494
rect 75 -497 94 -496
rect 124 -497 220 -496
rect 222 -497 577 -496
rect 86 -499 265 -498
rect 289 -499 297 -498
rect 310 -499 325 -498
rect 331 -499 451 -498
rect 82 -501 87 -500
rect 89 -501 129 -500
rect 156 -501 416 -500
rect 429 -501 451 -500
rect 170 -503 244 -502
rect 264 -503 269 -502
rect 296 -503 493 -502
rect 191 -505 262 -504
rect 320 -505 402 -504
rect 429 -505 444 -504
rect 478 -505 493 -504
rect 65 -507 262 -506
rect 282 -507 479 -506
rect 58 -509 66 -508
rect 201 -509 248 -508
rect 292 -509 444 -508
rect 201 -511 510 -510
rect 212 -513 318 -512
rect 366 -513 437 -512
rect 205 -515 213 -514
rect 226 -515 255 -514
rect 366 -515 521 -514
rect 79 -517 206 -516
rect 387 -517 521 -516
rect 23 -519 80 -518
rect 390 -519 500 -518
rect 9 -530 17 -529
rect 23 -530 129 -529
rect 131 -530 171 -529
rect 177 -530 188 -529
rect 198 -530 213 -529
rect 215 -530 220 -529
rect 226 -530 500 -529
rect 509 -530 556 -529
rect 16 -532 258 -531
rect 268 -532 272 -531
rect 275 -532 370 -531
rect 373 -532 528 -531
rect 30 -534 69 -533
rect 79 -534 101 -533
rect 107 -534 178 -533
rect 205 -534 293 -533
rect 296 -534 318 -533
rect 331 -534 367 -533
rect 373 -534 521 -533
rect 30 -536 69 -535
rect 103 -536 206 -535
rect 219 -536 514 -535
rect 37 -538 202 -537
rect 254 -538 300 -537
rect 306 -538 409 -537
rect 478 -538 535 -537
rect 40 -540 90 -539
rect 107 -540 164 -539
rect 254 -540 388 -539
rect 464 -540 479 -539
rect 485 -540 507 -539
rect 44 -542 139 -541
rect 156 -542 286 -541
rect 289 -542 377 -541
rect 492 -542 521 -541
rect 51 -544 185 -543
rect 208 -544 507 -543
rect 51 -546 76 -545
rect 114 -546 262 -545
rect 268 -546 304 -545
rect 313 -546 423 -545
rect 492 -546 531 -545
rect 58 -548 122 -547
rect 124 -548 146 -547
rect 149 -548 157 -547
rect 163 -548 279 -547
rect 282 -548 472 -547
rect 58 -550 73 -549
rect 117 -550 311 -549
rect 313 -550 444 -549
rect 121 -552 223 -551
rect 317 -552 325 -551
rect 331 -552 342 -551
rect 345 -552 451 -551
rect 128 -554 171 -553
rect 229 -554 325 -553
rect 348 -554 437 -553
rect 443 -554 458 -553
rect 135 -556 234 -555
rect 240 -556 437 -555
rect 149 -558 192 -557
rect 240 -558 262 -557
rect 352 -558 472 -557
rect 159 -560 192 -559
rect 338 -560 353 -559
rect 359 -560 409 -559
rect 415 -560 451 -559
rect 142 -562 360 -561
rect 362 -562 465 -561
rect 236 -564 339 -563
rect 394 -564 416 -563
rect 429 -564 458 -563
rect 394 -566 402 -565
rect 429 -566 486 -565
rect 264 -568 402 -567
rect 9 -579 90 -578
rect 121 -579 283 -578
rect 289 -579 304 -578
rect 338 -579 395 -578
rect 429 -579 451 -578
rect 464 -579 528 -578
rect 530 -579 542 -578
rect 9 -581 111 -580
rect 121 -581 132 -580
rect 135 -581 213 -580
rect 222 -581 332 -580
rect 338 -581 346 -580
rect 359 -581 416 -580
rect 432 -581 521 -580
rect 534 -581 549 -580
rect 23 -583 59 -582
rect 72 -583 83 -582
rect 86 -583 227 -582
rect 233 -583 248 -582
rect 254 -583 276 -582
rect 324 -583 332 -582
rect 341 -583 346 -582
rect 352 -583 360 -582
rect 366 -583 381 -582
rect 436 -583 500 -582
rect 520 -583 542 -582
rect 23 -585 101 -584
rect 135 -585 363 -584
rect 380 -585 388 -584
rect 436 -585 510 -584
rect 523 -585 535 -584
rect 30 -587 115 -586
rect 138 -587 164 -586
rect 170 -587 188 -586
rect 191 -587 220 -586
rect 236 -587 517 -586
rect 30 -589 52 -588
rect 54 -589 66 -588
rect 72 -589 129 -588
rect 145 -589 157 -588
rect 191 -589 286 -588
rect 352 -589 549 -588
rect 16 -591 52 -590
rect 58 -591 66 -590
rect 79 -591 118 -590
rect 142 -591 157 -590
rect 198 -591 230 -590
rect 240 -591 395 -590
rect 443 -591 465 -590
rect 471 -591 528 -590
rect 37 -593 45 -592
rect 79 -593 108 -592
rect 149 -593 174 -592
rect 198 -593 272 -592
rect 275 -593 318 -592
rect 387 -593 423 -592
rect 443 -593 458 -592
rect 481 -593 507 -592
rect 103 -595 164 -594
rect 205 -595 297 -594
rect 373 -595 458 -594
rect 485 -595 514 -594
rect 142 -597 374 -596
rect 401 -597 472 -596
rect 485 -597 493 -596
rect 499 -597 514 -596
rect 149 -599 311 -598
rect 450 -599 479 -598
rect 205 -601 328 -600
rect 208 -603 234 -602
rect 247 -603 262 -602
rect 268 -603 493 -602
rect 177 -605 269 -604
rect 289 -605 423 -604
rect 219 -607 300 -606
rect 306 -607 402 -606
rect 229 -609 318 -608
rect 261 -611 314 -610
rect 9 -622 69 -621
rect 72 -622 132 -621
rect 142 -622 227 -621
rect 233 -622 293 -621
rect 296 -622 381 -621
rect 394 -622 437 -621
rect 443 -622 475 -621
rect 499 -622 507 -621
rect 513 -622 584 -621
rect 16 -624 62 -623
rect 65 -624 118 -623
rect 163 -624 178 -623
rect 184 -624 199 -623
rect 219 -624 248 -623
rect 261 -624 419 -623
rect 422 -624 437 -623
rect 450 -624 489 -623
rect 516 -624 535 -623
rect 544 -624 556 -623
rect 23 -626 90 -625
rect 93 -626 101 -625
rect 103 -626 300 -625
rect 310 -626 360 -625
rect 401 -626 444 -625
rect 520 -626 542 -625
rect 555 -626 563 -625
rect 30 -628 48 -627
rect 51 -628 59 -627
rect 72 -628 80 -627
rect 96 -628 209 -627
rect 222 -628 262 -627
rect 275 -628 311 -627
rect 317 -628 451 -627
rect 527 -628 535 -627
rect 37 -630 45 -629
rect 107 -630 136 -629
rect 149 -630 178 -629
rect 226 -630 304 -629
rect 327 -630 430 -629
rect 44 -632 321 -631
rect 334 -632 388 -631
rect 397 -632 430 -631
rect 86 -634 108 -633
rect 114 -634 220 -633
rect 233 -634 251 -633
rect 275 -634 349 -633
rect 352 -634 458 -633
rect 75 -636 87 -635
rect 114 -636 248 -635
rect 296 -636 374 -635
rect 380 -636 398 -635
rect 408 -636 416 -635
rect 422 -636 472 -635
rect 131 -638 360 -637
rect 366 -638 472 -637
rect 149 -640 157 -639
rect 163 -640 213 -639
rect 240 -640 290 -639
rect 324 -640 458 -639
rect 128 -642 157 -641
rect 170 -642 188 -641
rect 191 -642 304 -641
rect 324 -642 531 -641
rect 40 -644 171 -643
rect 180 -644 192 -643
rect 205 -644 213 -643
rect 254 -644 290 -643
rect 331 -644 367 -643
rect 401 -644 409 -643
rect 254 -646 549 -645
rect 331 -648 388 -647
rect 481 -648 549 -647
rect 338 -650 479 -649
rect 341 -652 500 -651
rect 268 -654 342 -653
rect 345 -654 353 -653
rect 355 -654 493 -653
rect 345 -656 465 -655
rect 485 -656 493 -655
rect 464 -658 517 -657
rect 16 -669 66 -668
rect 107 -669 111 -668
rect 114 -669 136 -668
rect 156 -669 272 -668
rect 296 -669 318 -668
rect 320 -669 430 -668
rect 471 -669 619 -668
rect 628 -669 640 -668
rect 23 -671 104 -670
rect 156 -671 178 -670
rect 205 -671 213 -670
rect 240 -671 290 -670
rect 303 -671 405 -670
rect 471 -671 479 -670
rect 485 -671 489 -670
rect 499 -671 514 -670
rect 516 -671 521 -670
rect 527 -671 612 -670
rect 30 -673 38 -672
rect 44 -673 101 -672
rect 163 -673 167 -672
rect 170 -673 234 -672
rect 247 -673 304 -672
rect 345 -673 577 -672
rect 583 -673 647 -672
rect 44 -675 52 -674
rect 58 -675 80 -674
rect 93 -675 104 -674
rect 114 -675 164 -674
rect 170 -675 227 -674
rect 247 -675 300 -674
rect 348 -675 367 -674
rect 376 -675 416 -674
rect 478 -675 493 -674
rect 499 -675 556 -674
rect 593 -675 633 -674
rect 51 -677 335 -676
rect 352 -677 374 -676
rect 380 -677 402 -676
rect 415 -677 458 -676
rect 506 -677 521 -676
rect 530 -677 535 -676
rect 548 -677 563 -676
rect 65 -679 87 -678
rect 191 -679 227 -678
rect 250 -679 465 -678
rect 72 -681 80 -680
rect 86 -681 122 -680
rect 201 -681 206 -680
rect 212 -681 276 -680
rect 296 -681 556 -680
rect 121 -683 199 -682
rect 219 -683 276 -682
rect 324 -683 374 -682
rect 380 -683 605 -682
rect 177 -685 202 -684
rect 219 -685 244 -684
rect 254 -685 325 -684
rect 331 -685 535 -684
rect 184 -687 255 -686
rect 261 -687 290 -686
rect 338 -687 507 -686
rect 135 -689 262 -688
rect 268 -689 549 -688
rect 149 -691 185 -690
rect 194 -691 269 -690
rect 310 -691 339 -690
rect 359 -691 402 -690
rect 443 -691 458 -690
rect 128 -693 150 -692
rect 233 -693 311 -692
rect 366 -693 409 -692
rect 443 -693 545 -692
rect 282 -695 360 -694
rect 387 -695 584 -694
rect 387 -697 437 -696
rect 450 -697 465 -696
rect 345 -699 437 -698
rect 450 -699 573 -698
rect 394 -701 430 -700
rect 397 -703 423 -702
rect 408 -705 475 -704
rect 422 -707 542 -706
rect 16 -718 59 -717
rect 86 -718 136 -717
rect 142 -718 150 -717
rect 152 -718 188 -717
rect 194 -718 206 -717
rect 219 -718 255 -717
rect 261 -718 346 -717
rect 348 -718 416 -717
rect 422 -718 489 -717
rect 495 -718 535 -717
rect 541 -718 615 -717
rect 23 -720 66 -719
rect 79 -720 150 -719
rect 156 -720 262 -719
rect 268 -720 332 -719
rect 334 -720 472 -719
rect 474 -720 535 -719
rect 562 -720 601 -719
rect 611 -720 633 -719
rect 33 -722 38 -721
rect 44 -722 76 -721
rect 79 -722 115 -721
rect 156 -722 286 -721
rect 296 -722 325 -721
rect 338 -722 465 -721
rect 499 -722 573 -721
rect 593 -722 647 -721
rect 44 -724 122 -723
rect 163 -724 178 -723
rect 194 -724 304 -723
rect 310 -724 507 -723
rect 527 -724 531 -723
rect 569 -724 605 -723
rect 51 -726 258 -725
rect 268 -726 290 -725
rect 310 -726 360 -725
rect 366 -726 528 -725
rect 597 -726 640 -725
rect 51 -728 129 -727
rect 163 -728 230 -727
rect 240 -728 304 -727
rect 317 -728 325 -727
rect 352 -728 542 -727
rect 65 -730 73 -729
rect 86 -730 94 -729
rect 103 -730 458 -729
rect 464 -730 556 -729
rect 58 -732 104 -731
rect 114 -732 129 -731
rect 170 -732 202 -731
rect 205 -732 297 -731
rect 317 -732 332 -731
rect 352 -732 360 -731
rect 366 -732 514 -731
rect 555 -732 619 -731
rect 72 -734 108 -733
rect 121 -734 216 -733
rect 226 -734 241 -733
rect 247 -734 384 -733
rect 397 -734 521 -733
rect 93 -736 153 -735
rect 170 -736 213 -735
rect 250 -736 388 -735
rect 408 -736 521 -735
rect 107 -738 199 -737
rect 222 -738 388 -737
rect 408 -738 444 -737
rect 450 -738 458 -737
rect 506 -738 577 -737
rect 177 -740 192 -739
rect 222 -740 363 -739
rect 373 -740 493 -739
rect 184 -742 199 -741
rect 254 -742 349 -741
rect 380 -742 479 -741
rect 142 -744 185 -743
rect 275 -744 279 -743
rect 282 -744 402 -743
rect 415 -744 472 -743
rect 478 -744 549 -743
rect 292 -746 402 -745
rect 425 -746 584 -745
rect 334 -748 514 -747
rect 338 -750 451 -749
rect 380 -752 437 -751
rect 429 -754 500 -753
rect 394 -756 430 -755
rect 394 -758 437 -757
rect 26 -769 34 -768
rect 40 -769 150 -768
rect 152 -769 374 -768
rect 387 -769 395 -768
rect 397 -769 458 -768
rect 471 -769 521 -768
rect 534 -769 559 -768
rect 30 -771 38 -770
rect 44 -771 115 -770
rect 128 -771 167 -770
rect 170 -771 192 -770
rect 212 -771 269 -770
rect 275 -771 437 -770
rect 446 -771 479 -770
rect 492 -771 528 -770
rect 44 -773 94 -772
rect 128 -773 188 -772
rect 212 -773 311 -772
rect 324 -773 339 -772
rect 352 -773 461 -772
rect 513 -773 549 -772
rect 51 -775 146 -774
rect 156 -775 195 -774
rect 219 -775 262 -774
rect 285 -775 318 -774
rect 334 -775 486 -774
rect 499 -775 514 -774
rect 520 -775 556 -774
rect 51 -777 122 -776
rect 156 -777 192 -776
rect 222 -777 290 -776
rect 292 -777 377 -776
rect 401 -777 500 -776
rect 58 -779 143 -778
rect 163 -779 332 -778
rect 338 -779 444 -778
rect 492 -779 556 -778
rect 58 -781 66 -780
rect 72 -781 153 -780
rect 163 -781 283 -780
rect 303 -781 388 -780
rect 429 -781 535 -780
rect 65 -783 332 -782
rect 359 -783 465 -782
rect 72 -785 146 -784
rect 170 -785 258 -784
rect 261 -785 423 -784
rect 443 -785 531 -784
rect 86 -787 118 -786
rect 121 -787 437 -786
rect 464 -787 507 -786
rect 86 -789 206 -788
rect 226 -789 276 -788
rect 303 -789 353 -788
rect 359 -789 381 -788
rect 404 -789 430 -788
rect 93 -791 258 -790
rect 306 -791 479 -790
rect 177 -793 325 -792
rect 103 -795 178 -794
rect 184 -795 227 -794
rect 229 -795 367 -794
rect 205 -797 216 -796
rect 233 -797 269 -796
rect 313 -797 507 -796
rect 215 -799 220 -798
rect 236 -799 342 -798
rect 366 -799 409 -798
rect 247 -801 297 -800
rect 317 -801 472 -800
rect 247 -803 423 -802
rect 254 -805 542 -804
rect 296 -807 381 -806
rect 450 -807 542 -806
rect 376 -809 409 -808
rect 415 -809 451 -808
rect 107 -811 416 -810
rect 79 -813 108 -812
rect 79 -815 199 -814
rect 26 -826 41 -825
rect 44 -826 237 -825
rect 240 -826 248 -825
rect 254 -826 286 -825
rect 306 -826 486 -825
rect 30 -828 38 -827
rect 44 -828 73 -827
rect 75 -828 111 -827
rect 114 -828 143 -827
rect 145 -828 318 -827
rect 320 -828 388 -827
rect 401 -828 465 -827
rect 467 -828 542 -827
rect 51 -830 160 -829
rect 173 -830 195 -829
rect 201 -830 405 -829
rect 450 -830 486 -829
rect 37 -832 52 -831
rect 58 -832 181 -831
rect 187 -832 311 -831
rect 313 -832 549 -831
rect 79 -834 164 -833
rect 212 -834 220 -833
rect 240 -834 276 -833
rect 296 -834 451 -833
rect 457 -834 465 -833
rect 79 -836 171 -835
rect 177 -836 220 -835
rect 261 -836 325 -835
rect 331 -836 367 -835
rect 373 -836 514 -835
rect 86 -838 202 -837
rect 205 -838 262 -837
rect 310 -838 318 -837
rect 324 -838 360 -837
rect 366 -838 430 -837
rect 86 -840 136 -839
rect 149 -840 559 -839
rect 100 -842 227 -841
rect 257 -842 514 -841
rect 107 -844 192 -843
rect 226 -844 283 -843
rect 313 -844 472 -843
rect 117 -846 430 -845
rect 121 -848 304 -847
rect 348 -848 500 -847
rect 124 -850 129 -849
rect 149 -850 335 -849
rect 338 -850 500 -849
rect 93 -852 129 -851
rect 156 -852 276 -851
rect 289 -852 339 -851
rect 355 -852 535 -851
rect 65 -854 94 -853
rect 163 -854 185 -853
rect 247 -854 356 -853
rect 359 -854 409 -853
rect 520 -854 535 -853
rect 65 -856 199 -855
rect 268 -856 290 -855
rect 373 -856 507 -855
rect 268 -858 381 -857
rect 387 -858 475 -857
rect 492 -858 507 -857
rect 376 -860 528 -859
rect 348 -862 528 -861
rect 401 -864 437 -863
rect 408 -866 423 -865
rect 436 -866 479 -865
rect 352 -868 479 -867
rect 415 -870 493 -869
rect 394 -872 416 -871
rect 422 -872 444 -871
rect 152 -874 444 -873
rect 233 -876 395 -875
rect 233 -878 297 -877
rect 9 -889 136 -888
rect 142 -889 157 -888
rect 159 -889 493 -888
rect 520 -889 535 -888
rect 16 -891 209 -890
rect 240 -891 265 -890
rect 268 -891 335 -890
rect 348 -891 486 -890
rect 520 -891 524 -890
rect 23 -893 45 -892
rect 58 -893 346 -892
rect 355 -893 437 -892
rect 457 -893 493 -892
rect 44 -895 52 -894
rect 58 -895 73 -894
rect 79 -895 171 -894
rect 177 -895 213 -894
rect 240 -895 335 -894
rect 359 -895 363 -894
rect 380 -895 514 -894
rect 37 -897 213 -896
rect 233 -897 381 -896
rect 383 -897 514 -896
rect 51 -899 286 -898
rect 313 -899 409 -898
rect 422 -899 475 -898
rect 478 -899 486 -898
rect 65 -901 139 -900
rect 142 -901 255 -900
rect 282 -901 325 -900
rect 331 -901 500 -900
rect 65 -903 192 -902
rect 194 -903 262 -902
rect 282 -903 325 -902
rect 352 -903 500 -902
rect 86 -905 230 -904
rect 296 -905 423 -904
rect 436 -905 444 -904
rect 478 -905 507 -904
rect 93 -907 164 -906
rect 201 -907 293 -906
rect 317 -907 346 -906
rect 359 -907 402 -906
rect 506 -907 528 -906
rect 93 -909 129 -908
rect 149 -909 269 -908
rect 317 -909 339 -908
rect 394 -909 409 -908
rect 100 -911 181 -910
rect 205 -911 290 -910
rect 397 -911 472 -910
rect 107 -913 307 -912
rect 401 -913 416 -912
rect 107 -915 248 -914
rect 275 -915 339 -914
rect 415 -915 430 -914
rect 114 -917 150 -916
rect 152 -917 171 -916
rect 201 -917 248 -916
rect 306 -917 367 -916
rect 429 -917 451 -916
rect 121 -919 185 -918
rect 208 -919 297 -918
rect 387 -919 451 -918
rect 124 -921 167 -920
rect 184 -921 223 -920
rect 226 -921 234 -920
rect 362 -921 388 -920
rect 128 -923 195 -922
rect 219 -923 276 -922
rect 159 -925 311 -924
rect 166 -927 255 -926
rect 205 -929 311 -928
rect 219 -931 367 -930
rect 226 -933 458 -932
rect 2 -944 164 -943
rect 201 -944 423 -943
rect 443 -944 500 -943
rect 16 -946 104 -945
rect 107 -946 111 -945
rect 114 -946 139 -945
rect 142 -946 192 -945
rect 212 -946 241 -945
rect 257 -946 297 -945
rect 299 -946 416 -945
rect 429 -946 444 -945
rect 464 -946 486 -945
rect 9 -948 192 -947
rect 222 -948 262 -947
rect 268 -948 304 -947
rect 310 -948 409 -947
rect 467 -948 493 -947
rect 23 -950 31 -949
rect 37 -950 199 -949
rect 254 -950 311 -949
rect 324 -950 402 -949
rect 492 -950 514 -949
rect 9 -952 31 -951
rect 44 -952 185 -951
rect 187 -952 213 -951
rect 268 -952 276 -951
rect 296 -952 325 -951
rect 327 -952 416 -951
rect 16 -954 24 -953
rect 51 -954 167 -953
rect 198 -954 430 -953
rect 51 -956 59 -955
rect 65 -956 202 -955
rect 247 -956 276 -955
rect 338 -956 381 -955
rect 394 -956 479 -955
rect 65 -958 206 -957
rect 306 -958 395 -957
rect 478 -958 507 -957
rect 75 -960 101 -959
rect 107 -960 171 -959
rect 177 -960 206 -959
rect 331 -960 339 -959
rect 345 -960 402 -959
rect 506 -960 521 -959
rect 86 -962 157 -961
rect 163 -962 283 -961
rect 289 -962 346 -961
rect 352 -962 451 -961
rect 86 -964 293 -963
rect 373 -964 423 -963
rect 93 -966 104 -965
rect 110 -966 171 -965
rect 177 -966 265 -965
rect 373 -966 388 -965
rect 96 -968 472 -967
rect 114 -970 167 -969
rect 194 -970 248 -969
rect 264 -970 437 -969
rect 457 -970 472 -969
rect 121 -972 220 -971
rect 226 -972 458 -971
rect 128 -974 185 -973
rect 233 -974 283 -973
rect 359 -974 388 -973
rect 82 -976 234 -975
rect 355 -976 360 -975
rect 366 -976 437 -975
rect 135 -978 143 -977
rect 149 -978 230 -977
rect 334 -978 367 -977
rect 159 -980 220 -979
rect 334 -980 451 -979
rect 121 -982 160 -981
rect 9 -993 38 -992
rect 44 -993 220 -992
rect 229 -993 241 -992
rect 278 -993 381 -992
rect 418 -993 437 -992
rect 439 -993 479 -992
rect 488 -993 507 -992
rect 23 -995 34 -994
rect 37 -995 48 -994
rect 51 -995 59 -994
rect 65 -995 94 -994
rect 107 -995 185 -994
rect 187 -995 276 -994
rect 289 -995 318 -994
rect 341 -995 444 -994
rect 446 -995 479 -994
rect 40 -997 94 -996
rect 107 -997 195 -996
rect 215 -997 230 -996
rect 233 -997 346 -996
rect 352 -997 451 -996
rect 467 -997 472 -996
rect 474 -997 493 -996
rect 58 -999 62 -998
rect 79 -999 115 -998
rect 131 -999 325 -998
rect 327 -999 346 -998
rect 380 -999 388 -998
rect 415 -999 451 -998
rect 82 -1001 458 -1000
rect 2 -1003 83 -1002
rect 86 -1003 244 -1002
rect 285 -1003 290 -1002
rect 303 -1003 318 -1002
rect 334 -1003 353 -1002
rect 366 -1003 388 -1002
rect 422 -1003 465 -1002
rect 86 -1005 104 -1004
rect 149 -1005 160 -1004
rect 163 -1005 167 -1004
rect 170 -1005 227 -1004
rect 310 -1005 367 -1004
rect 96 -1007 115 -1006
rect 149 -1007 430 -1006
rect 156 -1009 171 -1008
rect 191 -1009 283 -1008
rect 415 -1009 430 -1008
rect 191 -1011 213 -1010
rect 222 -1011 311 -1010
rect 212 -1013 269 -1012
rect 128 -1015 269 -1014
rect 128 -1017 178 -1016
rect 222 -1017 409 -1016
rect 177 -1019 199 -1018
rect 394 -1019 409 -1018
rect 198 -1021 262 -1020
rect 373 -1021 395 -1020
rect 254 -1023 262 -1022
rect 373 -1023 461 -1022
rect 254 -1025 339 -1024
rect 338 -1027 402 -1026
rect 292 -1029 402 -1028
rect 23 -1040 34 -1039
rect 51 -1040 59 -1039
rect 72 -1040 80 -1039
rect 86 -1040 101 -1039
rect 117 -1040 122 -1039
rect 128 -1040 157 -1039
rect 159 -1040 297 -1039
rect 299 -1040 360 -1039
rect 408 -1040 423 -1039
rect 443 -1040 451 -1039
rect 460 -1040 468 -1039
rect 488 -1040 500 -1039
rect 30 -1042 38 -1041
rect 68 -1042 80 -1041
rect 100 -1042 115 -1041
rect 121 -1042 139 -1041
rect 149 -1042 171 -1041
rect 177 -1042 185 -1041
rect 205 -1042 227 -1041
rect 233 -1042 276 -1041
rect 285 -1042 318 -1041
rect 324 -1042 388 -1041
rect 401 -1042 423 -1041
rect 429 -1042 451 -1041
rect 464 -1042 472 -1041
rect 37 -1044 97 -1043
rect 110 -1044 157 -1043
rect 163 -1044 255 -1043
rect 261 -1044 307 -1043
rect 331 -1044 339 -1043
rect 345 -1044 360 -1043
rect 394 -1044 402 -1043
rect 408 -1044 496 -1043
rect 86 -1046 115 -1045
rect 128 -1046 486 -1045
rect 135 -1048 143 -1047
rect 177 -1048 220 -1047
rect 222 -1048 279 -1047
rect 303 -1048 367 -1047
rect 418 -1048 458 -1047
rect 478 -1048 486 -1047
rect 107 -1050 143 -1049
rect 184 -1050 192 -1049
rect 198 -1050 206 -1049
rect 215 -1050 388 -1049
rect 96 -1052 192 -1051
rect 198 -1052 416 -1051
rect 135 -1054 174 -1053
rect 233 -1054 262 -1053
rect 268 -1054 325 -1053
rect 338 -1054 430 -1053
rect 240 -1056 283 -1055
rect 303 -1056 444 -1055
rect 240 -1058 328 -1057
rect 341 -1058 458 -1057
rect 247 -1060 255 -1059
rect 268 -1060 367 -1059
rect 149 -1062 248 -1061
rect 278 -1062 318 -1061
rect 348 -1062 381 -1061
rect 310 -1064 395 -1063
rect 289 -1066 311 -1065
rect 373 -1066 381 -1065
rect 229 -1068 374 -1067
rect 289 -1070 353 -1069
rect 352 -1072 437 -1071
rect 345 -1074 437 -1073
rect 30 -1085 45 -1084
rect 47 -1085 62 -1084
rect 86 -1085 90 -1084
rect 96 -1085 178 -1084
rect 191 -1085 209 -1084
rect 212 -1085 325 -1084
rect 338 -1085 402 -1084
rect 432 -1085 465 -1084
rect 471 -1085 479 -1084
rect 481 -1085 486 -1084
rect 495 -1085 500 -1084
rect 37 -1087 202 -1086
rect 212 -1087 342 -1086
rect 345 -1087 388 -1086
rect 401 -1087 458 -1086
rect 51 -1089 66 -1088
rect 100 -1089 160 -1088
rect 170 -1089 248 -1088
rect 271 -1089 311 -1088
rect 338 -1089 374 -1088
rect 450 -1089 458 -1088
rect 58 -1091 111 -1090
rect 114 -1091 136 -1090
rect 149 -1091 241 -1090
rect 271 -1091 332 -1090
rect 348 -1091 381 -1090
rect 65 -1093 73 -1092
rect 100 -1093 122 -1092
rect 124 -1093 136 -1092
rect 149 -1093 227 -1092
rect 229 -1093 318 -1092
rect 352 -1093 388 -1092
rect 72 -1095 87 -1094
rect 163 -1095 171 -1094
rect 173 -1095 237 -1094
rect 240 -1095 248 -1094
rect 268 -1095 318 -1094
rect 366 -1095 377 -1094
rect 380 -1095 416 -1094
rect 82 -1097 122 -1096
rect 156 -1097 164 -1096
rect 177 -1097 223 -1096
rect 226 -1097 332 -1096
rect 366 -1097 444 -1096
rect 156 -1099 279 -1098
rect 289 -1099 360 -1098
rect 369 -1099 430 -1098
rect 194 -1101 216 -1100
rect 236 -1101 255 -1100
rect 275 -1101 297 -1100
rect 310 -1101 325 -1100
rect 359 -1101 395 -1100
rect 422 -1101 444 -1100
rect 107 -1103 216 -1102
rect 233 -1103 255 -1102
rect 261 -1103 297 -1102
rect 373 -1103 409 -1102
rect 145 -1105 262 -1104
rect 376 -1105 423 -1104
rect 205 -1107 223 -1106
rect 394 -1107 416 -1106
rect 47 -1118 52 -1117
rect 72 -1118 83 -1117
rect 100 -1118 125 -1117
rect 149 -1118 209 -1117
rect 212 -1118 223 -1117
rect 229 -1118 314 -1117
rect 334 -1118 388 -1117
rect 394 -1118 402 -1117
rect 408 -1118 444 -1117
rect 65 -1120 73 -1119
rect 100 -1120 269 -1119
rect 285 -1120 297 -1119
rect 306 -1120 332 -1119
rect 338 -1120 398 -1119
rect 408 -1120 416 -1119
rect 422 -1120 451 -1119
rect 65 -1122 76 -1121
rect 110 -1122 122 -1121
rect 149 -1122 227 -1121
rect 233 -1122 258 -1121
rect 275 -1122 297 -1121
rect 317 -1122 339 -1121
rect 352 -1122 360 -1121
rect 366 -1122 402 -1121
rect 415 -1122 433 -1121
rect 450 -1122 458 -1121
rect 114 -1124 143 -1123
rect 170 -1124 283 -1123
rect 289 -1124 311 -1123
rect 317 -1124 381 -1123
rect 387 -1124 405 -1123
rect 422 -1124 437 -1123
rect 114 -1126 129 -1125
rect 135 -1126 143 -1125
rect 170 -1126 230 -1125
rect 240 -1126 272 -1125
rect 310 -1126 346 -1125
rect 177 -1128 202 -1127
rect 205 -1128 234 -1127
rect 243 -1128 353 -1127
rect 184 -1130 192 -1129
rect 198 -1130 241 -1129
rect 247 -1130 304 -1129
rect 331 -1130 374 -1129
rect 163 -1132 192 -1131
rect 226 -1132 384 -1131
rect 254 -1134 276 -1133
rect 303 -1134 360 -1133
rect 156 -1136 255 -1135
rect 268 -1136 290 -1135
rect 324 -1136 374 -1135
rect 156 -1138 195 -1137
rect 250 -1138 325 -1137
rect 345 -1138 370 -1137
rect 177 -1140 195 -1139
rect 47 -1151 52 -1150
rect 58 -1151 83 -1150
rect 89 -1151 108 -1150
rect 114 -1151 185 -1150
rect 191 -1151 206 -1150
rect 212 -1151 297 -1150
rect 299 -1151 388 -1150
rect 394 -1151 405 -1150
rect 408 -1151 419 -1150
rect 446 -1151 451 -1150
rect 51 -1153 62 -1152
rect 65 -1153 87 -1152
rect 107 -1153 129 -1152
rect 135 -1153 150 -1152
rect 170 -1153 185 -1152
rect 194 -1153 283 -1152
rect 303 -1153 374 -1152
rect 65 -1155 188 -1154
rect 212 -1155 237 -1154
rect 240 -1155 339 -1154
rect 100 -1157 136 -1156
rect 142 -1157 146 -1156
rect 177 -1157 209 -1156
rect 222 -1157 234 -1156
rect 243 -1157 262 -1156
rect 271 -1157 318 -1156
rect 324 -1157 328 -1156
rect 338 -1157 367 -1156
rect 100 -1159 216 -1158
rect 226 -1159 346 -1158
rect 359 -1159 367 -1158
rect 117 -1161 122 -1160
rect 128 -1161 244 -1160
rect 247 -1161 360 -1160
rect 121 -1163 157 -1162
rect 226 -1163 283 -1162
rect 306 -1163 374 -1162
rect 156 -1165 164 -1164
rect 229 -1165 269 -1164
rect 310 -1165 381 -1164
rect 198 -1167 269 -1166
rect 296 -1167 311 -1166
rect 313 -1167 416 -1166
rect 233 -1169 290 -1168
rect 317 -1169 402 -1168
rect 415 -1169 430 -1168
rect 254 -1171 262 -1170
rect 324 -1171 332 -1170
rect 352 -1171 402 -1170
rect 247 -1173 353 -1172
rect 257 -1175 395 -1174
rect 327 -1177 332 -1176
rect 51 -1188 69 -1187
rect 72 -1188 76 -1187
rect 89 -1188 97 -1187
rect 100 -1188 143 -1187
rect 156 -1188 223 -1187
rect 229 -1188 276 -1187
rect 289 -1188 325 -1187
rect 338 -1188 349 -1187
rect 408 -1188 416 -1187
rect 422 -1188 426 -1187
rect 65 -1190 83 -1189
rect 93 -1190 101 -1189
rect 107 -1190 150 -1189
rect 166 -1190 199 -1189
rect 219 -1190 311 -1189
rect 324 -1190 353 -1189
rect 422 -1190 430 -1189
rect 79 -1192 167 -1191
rect 170 -1192 178 -1191
rect 184 -1192 202 -1191
rect 229 -1192 255 -1191
rect 268 -1192 293 -1191
rect 303 -1192 332 -1191
rect 345 -1192 388 -1191
rect 425 -1192 430 -1191
rect 79 -1194 115 -1193
rect 121 -1194 153 -1193
rect 159 -1194 178 -1193
rect 240 -1194 318 -1193
rect 331 -1194 342 -1193
rect 345 -1194 402 -1193
rect 107 -1196 146 -1195
rect 149 -1196 192 -1195
rect 233 -1196 241 -1195
rect 247 -1196 262 -1195
rect 282 -1196 304 -1195
rect 317 -1196 374 -1195
rect 128 -1198 227 -1197
rect 236 -1198 283 -1197
rect 289 -1198 360 -1197
rect 128 -1200 157 -1199
rect 184 -1200 227 -1199
rect 292 -1200 297 -1199
rect 359 -1200 367 -1199
rect 135 -1202 174 -1201
rect 366 -1202 395 -1201
rect 121 -1204 136 -1203
rect 138 -1204 223 -1203
rect 33 -1215 38 -1214
rect 44 -1215 52 -1214
rect 58 -1215 66 -1214
rect 72 -1215 80 -1214
rect 89 -1215 101 -1214
rect 107 -1215 174 -1214
rect 180 -1215 206 -1214
rect 229 -1215 248 -1214
rect 254 -1215 269 -1214
rect 303 -1215 342 -1214
rect 373 -1215 381 -1214
rect 401 -1215 409 -1214
rect 422 -1215 430 -1214
rect 72 -1217 80 -1216
rect 93 -1217 139 -1216
rect 152 -1217 160 -1216
rect 163 -1217 213 -1216
rect 229 -1217 241 -1216
rect 243 -1217 293 -1216
rect 296 -1217 304 -1216
rect 306 -1217 325 -1216
rect 331 -1217 353 -1216
rect 425 -1217 433 -1216
rect 114 -1219 122 -1218
rect 128 -1219 143 -1218
rect 163 -1219 178 -1218
rect 184 -1219 202 -1218
rect 212 -1219 255 -1218
rect 275 -1219 293 -1218
rect 310 -1219 346 -1218
rect 352 -1219 367 -1218
rect 100 -1221 129 -1220
rect 135 -1221 157 -1220
rect 170 -1221 188 -1220
rect 191 -1221 223 -1220
rect 282 -1221 311 -1220
rect 317 -1221 321 -1220
rect 338 -1221 346 -1220
rect 366 -1221 374 -1220
rect 121 -1223 150 -1222
rect 194 -1223 199 -1222
rect 215 -1223 318 -1222
rect 124 -1225 143 -1224
rect 222 -1225 234 -1224
rect 282 -1225 314 -1224
rect 219 -1227 234 -1226
rect 30 -1238 38 -1237
rect 44 -1238 52 -1237
rect 65 -1238 76 -1237
rect 93 -1238 118 -1237
rect 128 -1238 150 -1237
rect 152 -1238 209 -1237
rect 222 -1238 269 -1237
rect 275 -1238 290 -1237
rect 299 -1238 311 -1237
rect 324 -1238 328 -1237
rect 334 -1238 339 -1237
rect 369 -1238 374 -1237
rect 401 -1238 409 -1237
rect 415 -1238 423 -1237
rect 100 -1240 115 -1239
rect 128 -1240 139 -1239
rect 142 -1240 146 -1239
rect 163 -1240 216 -1239
rect 226 -1240 279 -1239
rect 338 -1240 353 -1239
rect 103 -1242 122 -1241
rect 177 -1242 192 -1241
rect 194 -1242 241 -1241
rect 250 -1242 269 -1241
rect 110 -1244 115 -1243
rect 205 -1244 283 -1243
rect 208 -1246 255 -1245
rect 212 -1248 223 -1247
rect 233 -1248 258 -1247
rect 170 -1250 234 -1249
rect 170 -1252 185 -1251
rect 219 -1252 241 -1251
rect 30 -1263 38 -1262
rect 58 -1263 69 -1262
rect 72 -1263 80 -1262
rect 107 -1263 115 -1262
rect 121 -1263 153 -1262
rect 170 -1263 206 -1262
rect 208 -1263 213 -1262
rect 226 -1263 269 -1262
rect 285 -1263 290 -1262
rect 296 -1263 304 -1262
rect 317 -1263 325 -1262
rect 338 -1263 349 -1262
rect 355 -1263 360 -1262
rect 128 -1265 139 -1264
rect 142 -1265 164 -1264
rect 177 -1265 188 -1264
rect 198 -1265 234 -1264
rect 250 -1265 262 -1264
<< m2contact >>
rect 138 0 139 1
rect 149 0 150 1
rect 177 0 178 1
rect 191 0 192 1
rect 198 0 199 1
rect 215 0 216 1
rect 226 0 227 1
rect 240 0 241 1
rect 187 -2 188 -1
rect 205 -2 206 -1
rect 212 -2 213 -1
rect 219 -2 220 -1
rect 135 -13 136 -12
rect 184 -13 185 -12
rect 187 -13 188 -12
rect 229 -13 230 -12
rect 240 -13 241 -12
rect 247 -13 248 -12
rect 324 -13 325 -12
rect 331 -13 332 -12
rect 145 -15 146 -14
rect 149 -15 150 -14
rect 163 -15 164 -14
rect 170 -15 171 -14
rect 177 -15 178 -14
rect 184 -15 185 -14
rect 191 -15 192 -14
rect 233 -15 234 -14
rect 156 -17 157 -16
rect 177 -17 178 -16
rect 198 -17 199 -16
rect 205 -17 206 -16
rect 208 -17 209 -16
rect 219 -17 220 -16
rect 226 -17 227 -16
rect 254 -17 255 -16
rect 198 -19 199 -18
rect 215 -19 216 -18
rect 219 -19 220 -18
rect 240 -19 241 -18
rect 229 -21 230 -20
rect 236 -21 237 -20
rect 128 -32 129 -31
rect 145 -32 146 -31
rect 198 -32 199 -31
rect 219 -32 220 -31
rect 222 -32 223 -31
rect 261 -32 262 -31
rect 268 -32 269 -31
rect 289 -32 290 -31
rect 296 -32 297 -31
rect 303 -32 304 -31
rect 324 -32 325 -31
rect 331 -32 332 -31
rect 135 -34 136 -33
rect 152 -34 153 -33
rect 198 -34 199 -33
rect 247 -34 248 -33
rect 327 -34 328 -33
rect 331 -34 332 -33
rect 135 -36 136 -35
rect 152 -36 153 -35
rect 201 -36 202 -35
rect 233 -36 234 -35
rect 142 -38 143 -37
rect 159 -38 160 -37
rect 173 -38 174 -37
rect 233 -38 234 -37
rect 159 -40 160 -39
rect 177 -40 178 -39
rect 205 -40 206 -39
rect 226 -40 227 -39
rect 163 -42 164 -41
rect 177 -42 178 -41
rect 205 -42 206 -41
rect 240 -42 241 -41
rect 163 -44 164 -43
rect 184 -44 185 -43
rect 208 -44 209 -43
rect 212 -44 213 -43
rect 226 -44 227 -43
rect 282 -44 283 -43
rect 229 -46 230 -45
rect 240 -46 241 -45
rect 191 -48 192 -47
rect 229 -48 230 -47
rect 103 -59 104 -58
rect 107 -59 108 -58
rect 121 -59 122 -58
rect 135 -59 136 -58
rect 142 -59 143 -58
rect 163 -59 164 -58
rect 205 -59 206 -58
rect 212 -59 213 -58
rect 226 -59 227 -58
rect 247 -59 248 -58
rect 261 -59 262 -58
rect 313 -59 314 -58
rect 128 -61 129 -60
rect 159 -61 160 -60
rect 191 -61 192 -60
rect 261 -61 262 -60
rect 268 -61 269 -60
rect 282 -61 283 -60
rect 289 -61 290 -60
rect 306 -61 307 -60
rect 142 -63 143 -62
rect 149 -63 150 -62
rect 184 -63 185 -62
rect 191 -63 192 -62
rect 229 -63 230 -62
rect 233 -63 234 -62
rect 240 -63 241 -62
rect 254 -63 255 -62
rect 275 -63 276 -62
rect 278 -63 279 -62
rect 282 -63 283 -62
rect 299 -63 300 -62
rect 177 -65 178 -64
rect 184 -65 185 -64
rect 201 -65 202 -64
rect 240 -65 241 -64
rect 296 -65 297 -64
rect 303 -65 304 -64
rect 219 -67 220 -66
rect 254 -67 255 -66
rect 292 -67 293 -66
rect 296 -67 297 -66
rect 170 -69 171 -68
rect 219 -69 220 -68
rect 166 -71 167 -70
rect 170 -71 171 -70
rect 100 -82 101 -81
rect 107 -82 108 -81
rect 114 -82 115 -81
rect 131 -82 132 -81
rect 138 -82 139 -81
rect 149 -82 150 -81
rect 159 -82 160 -81
rect 163 -82 164 -81
rect 166 -82 167 -81
rect 177 -82 178 -81
rect 184 -82 185 -81
rect 194 -82 195 -81
rect 205 -82 206 -81
rect 212 -82 213 -81
rect 229 -82 230 -81
rect 254 -82 255 -81
rect 275 -82 276 -81
rect 303 -82 304 -81
rect 317 -82 318 -81
rect 324 -82 325 -81
rect 107 -84 108 -83
rect 128 -84 129 -83
rect 149 -84 150 -83
rect 170 -84 171 -83
rect 191 -84 192 -83
rect 198 -84 199 -83
rect 222 -84 223 -83
rect 229 -84 230 -83
rect 233 -84 234 -83
rect 247 -84 248 -83
rect 282 -84 283 -83
rect 292 -84 293 -83
rect 296 -84 297 -83
rect 310 -84 311 -83
rect 317 -84 318 -83
rect 320 -84 321 -83
rect 324 -84 325 -83
rect 331 -84 332 -83
rect 121 -86 122 -85
rect 145 -86 146 -85
rect 198 -86 199 -85
rect 215 -86 216 -85
rect 219 -86 220 -85
rect 247 -86 248 -85
rect 117 -88 118 -87
rect 121 -88 122 -87
rect 128 -88 129 -87
rect 135 -88 136 -87
rect 142 -88 143 -87
rect 145 -88 146 -87
rect 222 -88 223 -87
rect 296 -88 297 -87
rect 226 -90 227 -89
rect 254 -90 255 -89
rect 236 -92 237 -91
rect 261 -92 262 -91
rect 240 -94 241 -93
rect 275 -94 276 -93
rect 261 -96 262 -95
rect 271 -96 272 -95
rect 86 -107 87 -106
rect 103 -107 104 -106
rect 107 -107 108 -106
rect 128 -107 129 -106
rect 135 -107 136 -106
rect 145 -107 146 -106
rect 149 -107 150 -106
rect 180 -107 181 -106
rect 198 -107 199 -106
rect 219 -107 220 -106
rect 229 -107 230 -106
rect 275 -107 276 -106
rect 282 -107 283 -106
rect 296 -107 297 -106
rect 380 -107 381 -106
rect 383 -107 384 -106
rect 114 -109 115 -108
rect 124 -109 125 -108
rect 135 -109 136 -108
rect 163 -109 164 -108
rect 198 -109 199 -108
rect 212 -109 213 -108
rect 215 -109 216 -108
rect 233 -109 234 -108
rect 243 -109 244 -108
rect 303 -109 304 -108
rect 103 -111 104 -110
rect 114 -111 115 -110
rect 156 -111 157 -110
rect 184 -111 185 -110
rect 205 -111 206 -110
rect 236 -111 237 -110
rect 247 -111 248 -110
rect 271 -111 272 -110
rect 289 -111 290 -110
rect 310 -111 311 -110
rect 107 -113 108 -112
rect 124 -113 125 -112
rect 163 -113 164 -112
rect 170 -113 171 -112
rect 177 -113 178 -112
rect 215 -113 216 -112
rect 268 -113 269 -112
rect 317 -113 318 -112
rect 180 -115 181 -114
rect 205 -115 206 -114
rect 208 -115 209 -114
rect 219 -115 220 -114
rect 261 -115 262 -114
rect 268 -115 269 -114
rect 303 -115 304 -114
rect 324 -115 325 -114
rect 184 -117 185 -116
rect 191 -117 192 -116
rect 212 -117 213 -116
rect 299 -117 300 -116
rect 310 -117 311 -116
rect 317 -117 318 -116
rect 254 -119 255 -118
rect 261 -119 262 -118
rect 226 -121 227 -120
rect 254 -121 255 -120
rect 79 -132 80 -131
rect 82 -132 83 -131
rect 107 -132 108 -131
rect 142 -132 143 -131
rect 156 -132 157 -131
rect 194 -132 195 -131
rect 219 -132 220 -131
rect 233 -132 234 -131
rect 257 -132 258 -131
rect 261 -132 262 -131
rect 268 -132 269 -131
rect 271 -132 272 -131
rect 296 -132 297 -131
rect 303 -132 304 -131
rect 310 -132 311 -131
rect 317 -132 318 -131
rect 380 -132 381 -131
rect 387 -132 388 -131
rect 79 -134 80 -133
rect 86 -134 87 -133
rect 107 -134 108 -133
rect 117 -134 118 -133
rect 131 -134 132 -133
rect 138 -134 139 -133
rect 159 -134 160 -133
rect 215 -134 216 -133
rect 226 -134 227 -133
rect 268 -134 269 -133
rect 275 -134 276 -133
rect 317 -134 318 -133
rect 114 -136 115 -135
rect 121 -136 122 -135
rect 128 -136 129 -135
rect 131 -136 132 -135
rect 135 -136 136 -135
rect 152 -136 153 -135
rect 163 -136 164 -135
rect 177 -136 178 -135
rect 184 -136 185 -135
rect 229 -136 230 -135
rect 254 -136 255 -135
rect 261 -136 262 -135
rect 299 -136 300 -135
rect 324 -136 325 -135
rect 128 -138 129 -137
rect 156 -138 157 -137
rect 170 -138 171 -137
rect 254 -138 255 -137
rect 145 -140 146 -139
rect 163 -140 164 -139
rect 173 -140 174 -139
rect 177 -140 178 -139
rect 191 -140 192 -139
rect 215 -140 216 -139
rect 121 -142 122 -141
rect 173 -142 174 -141
rect 205 -142 206 -141
rect 219 -142 220 -141
rect 152 -144 153 -143
rect 208 -144 209 -143
rect 205 -146 206 -145
rect 240 -146 241 -145
rect 107 -157 108 -156
rect 152 -157 153 -156
rect 156 -157 157 -156
rect 163 -157 164 -156
rect 173 -157 174 -156
rect 177 -157 178 -156
rect 187 -157 188 -156
rect 191 -157 192 -156
rect 198 -157 199 -156
rect 226 -157 227 -156
rect 233 -157 234 -156
rect 247 -157 248 -156
rect 254 -157 255 -156
rect 303 -157 304 -156
rect 317 -157 318 -156
rect 341 -157 342 -156
rect 359 -157 360 -156
rect 373 -157 374 -156
rect 387 -157 388 -156
rect 394 -157 395 -156
rect 408 -157 409 -156
rect 415 -157 416 -156
rect 436 -157 437 -156
rect 443 -157 444 -156
rect 114 -159 115 -158
rect 117 -159 118 -158
rect 121 -159 122 -158
rect 135 -159 136 -158
rect 152 -159 153 -158
rect 184 -159 185 -158
rect 212 -159 213 -158
rect 254 -159 255 -158
rect 261 -159 262 -158
rect 271 -159 272 -158
rect 296 -159 297 -158
rect 313 -159 314 -158
rect 317 -159 318 -158
rect 324 -159 325 -158
rect 331 -159 332 -158
rect 352 -159 353 -158
rect 362 -159 363 -158
rect 380 -159 381 -158
rect 383 -159 384 -158
rect 387 -159 388 -158
rect 124 -161 125 -160
rect 138 -161 139 -160
rect 163 -161 164 -160
rect 201 -161 202 -160
rect 205 -161 206 -160
rect 212 -161 213 -160
rect 215 -161 216 -160
rect 219 -161 220 -160
rect 226 -161 227 -160
rect 366 -161 367 -160
rect 135 -163 136 -162
rect 145 -163 146 -162
rect 170 -163 171 -162
rect 191 -163 192 -162
rect 205 -163 206 -162
rect 215 -163 216 -162
rect 219 -163 220 -162
rect 229 -163 230 -162
rect 233 -163 234 -162
rect 289 -163 290 -162
rect 320 -163 321 -162
rect 345 -163 346 -162
rect 177 -165 178 -164
rect 243 -165 244 -164
rect 261 -165 262 -164
rect 275 -165 276 -164
rect 278 -165 279 -164
rect 324 -165 325 -164
rect 240 -167 241 -166
rect 282 -167 283 -166
rect 268 -169 269 -168
rect 383 -169 384 -168
rect 75 -180 76 -179
rect 79 -180 80 -179
rect 86 -180 87 -179
rect 121 -180 122 -179
rect 135 -180 136 -179
rect 142 -180 143 -179
rect 149 -180 150 -179
rect 198 -180 199 -179
rect 229 -180 230 -179
rect 247 -180 248 -179
rect 250 -180 251 -179
rect 359 -180 360 -179
rect 369 -180 370 -179
rect 387 -180 388 -179
rect 415 -180 416 -179
rect 422 -180 423 -179
rect 432 -180 433 -179
rect 443 -180 444 -179
rect 89 -182 90 -181
rect 93 -182 94 -181
rect 107 -182 108 -181
rect 128 -182 129 -181
rect 156 -182 157 -181
rect 159 -182 160 -181
rect 163 -182 164 -181
rect 268 -182 269 -181
rect 271 -182 272 -181
rect 324 -182 325 -181
rect 338 -182 339 -181
rect 373 -182 374 -181
rect 383 -182 384 -181
rect 394 -182 395 -181
rect 401 -182 402 -181
rect 415 -182 416 -181
rect 436 -182 437 -181
rect 443 -182 444 -181
rect 121 -184 122 -183
rect 135 -184 136 -183
rect 170 -184 171 -183
rect 212 -184 213 -183
rect 233 -184 234 -183
rect 261 -184 262 -183
rect 296 -184 297 -183
rect 313 -184 314 -183
rect 317 -184 318 -183
rect 355 -184 356 -183
rect 380 -184 381 -183
rect 394 -184 395 -183
rect 170 -186 171 -185
rect 219 -186 220 -185
rect 229 -186 230 -185
rect 233 -186 234 -185
rect 254 -186 255 -185
rect 275 -186 276 -185
rect 303 -186 304 -185
rect 310 -186 311 -185
rect 317 -186 318 -185
rect 331 -186 332 -185
rect 345 -186 346 -185
rect 373 -186 374 -185
rect 177 -188 178 -187
rect 215 -188 216 -187
rect 219 -188 220 -187
rect 275 -188 276 -187
rect 285 -188 286 -187
rect 345 -188 346 -187
rect 177 -190 178 -189
rect 184 -190 185 -189
rect 191 -190 192 -189
rect 205 -190 206 -189
rect 254 -190 255 -189
rect 282 -190 283 -189
rect 285 -190 286 -189
rect 352 -190 353 -189
rect 163 -192 164 -191
rect 205 -192 206 -191
rect 261 -192 262 -191
rect 324 -192 325 -191
rect 331 -192 332 -191
rect 366 -192 367 -191
rect 184 -194 185 -193
rect 240 -194 241 -193
rect 296 -194 297 -193
rect 303 -194 304 -193
rect 201 -196 202 -195
rect 240 -196 241 -195
rect 72 -207 73 -206
rect 96 -207 97 -206
rect 100 -207 101 -206
rect 121 -207 122 -206
rect 128 -207 129 -206
rect 226 -207 227 -206
rect 261 -207 262 -206
rect 331 -207 332 -206
rect 345 -207 346 -206
rect 387 -207 388 -206
rect 394 -207 395 -206
rect 401 -207 402 -206
rect 404 -207 405 -206
rect 408 -207 409 -206
rect 415 -207 416 -206
rect 422 -207 423 -206
rect 436 -207 437 -206
rect 439 -207 440 -206
rect 79 -209 80 -208
rect 86 -209 87 -208
rect 103 -209 104 -208
rect 107 -209 108 -208
rect 121 -209 122 -208
rect 247 -209 248 -208
rect 268 -209 269 -208
rect 303 -209 304 -208
rect 306 -209 307 -208
rect 317 -209 318 -208
rect 373 -209 374 -208
rect 383 -209 384 -208
rect 79 -211 80 -210
rect 145 -211 146 -210
rect 149 -211 150 -210
rect 229 -211 230 -210
rect 236 -211 237 -210
rect 345 -211 346 -210
rect 373 -211 374 -210
rect 380 -211 381 -210
rect 86 -213 87 -212
rect 187 -213 188 -212
rect 191 -213 192 -212
rect 219 -213 220 -212
rect 222 -213 223 -212
rect 240 -213 241 -212
rect 257 -213 258 -212
rect 268 -213 269 -212
rect 275 -213 276 -212
rect 317 -213 318 -212
rect 359 -213 360 -212
rect 380 -213 381 -212
rect 93 -215 94 -214
rect 149 -215 150 -214
rect 156 -215 157 -214
rect 180 -215 181 -214
rect 198 -215 199 -214
rect 247 -215 248 -214
rect 310 -215 311 -214
rect 331 -215 332 -214
rect 107 -217 108 -216
rect 219 -217 220 -216
rect 229 -217 230 -216
rect 338 -217 339 -216
rect 142 -219 143 -218
rect 163 -219 164 -218
rect 170 -219 171 -218
rect 264 -219 265 -218
rect 296 -219 297 -218
rect 310 -219 311 -218
rect 324 -219 325 -218
rect 338 -219 339 -218
rect 159 -221 160 -220
rect 191 -221 192 -220
rect 201 -221 202 -220
rect 275 -221 276 -220
rect 324 -221 325 -220
rect 352 -221 353 -220
rect 170 -223 171 -222
rect 177 -223 178 -222
rect 205 -223 206 -222
rect 254 -223 255 -222
rect 352 -223 353 -222
rect 369 -223 370 -222
rect 131 -225 132 -224
rect 177 -225 178 -224
rect 184 -225 185 -224
rect 205 -225 206 -224
rect 212 -225 213 -224
rect 296 -225 297 -224
rect 212 -227 213 -226
rect 233 -227 234 -226
rect 240 -227 241 -226
rect 359 -227 360 -226
rect 233 -229 234 -228
rect 282 -229 283 -228
rect 68 -240 69 -239
rect 156 -240 157 -239
rect 170 -240 171 -239
rect 187 -240 188 -239
rect 229 -240 230 -239
rect 317 -240 318 -239
rect 359 -240 360 -239
rect 443 -240 444 -239
rect 450 -240 451 -239
rect 457 -240 458 -239
rect 530 -240 531 -239
rect 534 -240 535 -239
rect 86 -242 87 -241
rect 159 -242 160 -241
rect 170 -242 171 -241
rect 205 -242 206 -241
rect 240 -242 241 -241
rect 275 -242 276 -241
rect 292 -242 293 -241
rect 359 -242 360 -241
rect 366 -242 367 -241
rect 453 -242 454 -241
rect 79 -244 80 -243
rect 205 -244 206 -243
rect 243 -244 244 -243
rect 303 -244 304 -243
rect 331 -244 332 -243
rect 366 -244 367 -243
rect 369 -244 370 -243
rect 387 -244 388 -243
rect 394 -244 395 -243
rect 439 -244 440 -243
rect 72 -246 73 -245
rect 79 -246 80 -245
rect 93 -246 94 -245
rect 184 -246 185 -245
rect 194 -246 195 -245
rect 240 -246 241 -245
rect 250 -246 251 -245
rect 345 -246 346 -245
rect 418 -246 419 -245
rect 422 -246 423 -245
rect 93 -248 94 -247
rect 212 -248 213 -247
rect 254 -248 255 -247
rect 264 -248 265 -247
rect 271 -248 272 -247
rect 338 -248 339 -247
rect 345 -248 346 -247
rect 352 -248 353 -247
rect 373 -248 374 -247
rect 422 -248 423 -247
rect 100 -250 101 -249
rect 135 -250 136 -249
rect 138 -250 139 -249
rect 187 -250 188 -249
rect 208 -250 209 -249
rect 373 -250 374 -249
rect 408 -250 409 -249
rect 418 -250 419 -249
rect 107 -252 108 -251
rect 166 -252 167 -251
rect 177 -252 178 -251
rect 191 -252 192 -251
rect 212 -252 213 -251
rect 247 -252 248 -251
rect 254 -252 255 -251
rect 380 -252 381 -251
rect 107 -254 108 -253
rect 114 -254 115 -253
rect 121 -254 122 -253
rect 226 -254 227 -253
rect 257 -254 258 -253
rect 317 -254 318 -253
rect 338 -254 339 -253
rect 415 -254 416 -253
rect 114 -256 115 -255
rect 145 -256 146 -255
rect 180 -256 181 -255
rect 233 -256 234 -255
rect 261 -256 262 -255
rect 324 -256 325 -255
rect 121 -258 122 -257
rect 149 -258 150 -257
rect 198 -258 199 -257
rect 226 -258 227 -257
rect 261 -258 262 -257
rect 268 -258 269 -257
rect 275 -258 276 -257
rect 299 -258 300 -257
rect 303 -258 304 -257
rect 387 -258 388 -257
rect 128 -260 129 -259
rect 163 -260 164 -259
rect 268 -260 269 -259
rect 331 -260 332 -259
rect 131 -262 132 -261
rect 215 -262 216 -261
rect 296 -262 297 -261
rect 429 -262 430 -261
rect 135 -264 136 -263
rect 156 -264 157 -263
rect 296 -264 297 -263
rect 401 -264 402 -263
rect 142 -266 143 -265
rect 152 -266 153 -265
rect 310 -266 311 -265
rect 352 -266 353 -265
rect 86 -268 87 -267
rect 152 -268 153 -267
rect 219 -268 220 -267
rect 310 -268 311 -267
rect 149 -270 150 -269
rect 282 -270 283 -269
rect 282 -272 283 -271
rect 289 -272 290 -271
rect 30 -283 31 -282
rect 37 -283 38 -282
rect 47 -283 48 -282
rect 149 -283 150 -282
rect 177 -283 178 -282
rect 212 -283 213 -282
rect 222 -283 223 -282
rect 261 -283 262 -282
rect 268 -283 269 -282
rect 401 -283 402 -282
rect 415 -283 416 -282
rect 436 -283 437 -282
rect 453 -283 454 -282
rect 457 -283 458 -282
rect 527 -283 528 -282
rect 534 -283 535 -282
rect 30 -285 31 -284
rect 33 -285 34 -284
rect 51 -285 52 -284
rect 54 -285 55 -284
rect 58 -285 59 -284
rect 131 -285 132 -284
rect 135 -285 136 -284
rect 163 -285 164 -284
rect 184 -285 185 -284
rect 219 -285 220 -284
rect 243 -285 244 -284
rect 450 -285 451 -284
rect 68 -287 69 -286
rect 184 -287 185 -286
rect 194 -287 195 -286
rect 394 -287 395 -286
rect 401 -287 402 -286
rect 422 -287 423 -286
rect 75 -289 76 -288
rect 79 -289 80 -288
rect 82 -289 83 -288
rect 191 -289 192 -288
rect 205 -289 206 -288
rect 219 -289 220 -288
rect 247 -289 248 -288
rect 289 -289 290 -288
rect 292 -289 293 -288
rect 366 -289 367 -288
rect 387 -289 388 -288
rect 422 -289 423 -288
rect 86 -291 87 -290
rect 103 -291 104 -290
rect 107 -291 108 -290
rect 121 -291 122 -290
rect 149 -291 150 -290
rect 170 -291 171 -290
rect 208 -291 209 -290
rect 240 -291 241 -290
rect 254 -291 255 -290
rect 352 -291 353 -290
rect 380 -291 381 -290
rect 387 -291 388 -290
rect 394 -291 395 -290
rect 408 -291 409 -290
rect 93 -293 94 -292
rect 261 -293 262 -292
rect 268 -293 269 -292
rect 275 -293 276 -292
rect 282 -293 283 -292
rect 303 -293 304 -292
rect 306 -293 307 -292
rect 310 -293 311 -292
rect 338 -293 339 -292
rect 366 -293 367 -292
rect 408 -293 409 -292
rect 418 -293 419 -292
rect 93 -295 94 -294
rect 114 -295 115 -294
rect 121 -295 122 -294
rect 145 -295 146 -294
rect 156 -295 157 -294
rect 177 -295 178 -294
rect 226 -295 227 -294
rect 275 -295 276 -294
rect 296 -295 297 -294
rect 429 -295 430 -294
rect 100 -297 101 -296
rect 152 -297 153 -296
rect 163 -297 164 -296
rect 324 -297 325 -296
rect 352 -297 353 -296
rect 376 -297 377 -296
rect 114 -299 115 -298
rect 198 -299 199 -298
rect 226 -299 227 -298
rect 247 -299 248 -298
rect 299 -299 300 -298
rect 443 -299 444 -298
rect 128 -301 129 -300
rect 282 -301 283 -300
rect 310 -301 311 -300
rect 317 -301 318 -300
rect 142 -303 143 -302
rect 296 -303 297 -302
rect 317 -303 318 -302
rect 345 -303 346 -302
rect 170 -305 171 -304
rect 338 -305 339 -304
rect 198 -307 199 -306
rect 233 -307 234 -306
rect 331 -307 332 -306
rect 345 -307 346 -306
rect 187 -309 188 -308
rect 233 -309 234 -308
rect 331 -309 332 -308
rect 359 -309 360 -308
rect 229 -311 230 -310
rect 380 -311 381 -310
rect 359 -313 360 -312
rect 373 -313 374 -312
rect 19 -324 20 -323
rect 23 -324 24 -323
rect 37 -324 38 -323
rect 93 -324 94 -323
rect 96 -324 97 -323
rect 166 -324 167 -323
rect 194 -324 195 -323
rect 275 -324 276 -323
rect 282 -324 283 -323
rect 366 -324 367 -323
rect 373 -324 374 -323
rect 471 -324 472 -323
rect 513 -324 514 -323
rect 520 -324 521 -323
rect 523 -324 524 -323
rect 527 -324 528 -323
rect 51 -326 52 -325
rect 201 -326 202 -325
rect 219 -326 220 -325
rect 296 -326 297 -325
rect 327 -326 328 -325
rect 331 -326 332 -325
rect 408 -326 409 -325
rect 415 -326 416 -325
rect 422 -326 423 -325
rect 457 -326 458 -325
rect 58 -328 59 -327
rect 107 -328 108 -327
rect 110 -328 111 -327
rect 138 -328 139 -327
rect 145 -328 146 -327
rect 156 -328 157 -327
rect 159 -328 160 -327
rect 177 -328 178 -327
rect 198 -328 199 -327
rect 243 -328 244 -327
rect 247 -328 248 -327
rect 317 -328 318 -327
rect 331 -328 332 -327
rect 380 -328 381 -327
rect 390 -328 391 -327
rect 408 -328 409 -327
rect 436 -328 437 -327
rect 467 -328 468 -327
rect 58 -330 59 -329
rect 86 -330 87 -329
rect 100 -330 101 -329
rect 149 -330 150 -329
rect 177 -330 178 -329
rect 184 -330 185 -329
rect 198 -330 199 -329
rect 380 -330 381 -329
rect 387 -330 388 -329
rect 436 -330 437 -329
rect 65 -332 66 -331
rect 135 -332 136 -331
rect 149 -332 150 -331
rect 170 -332 171 -331
rect 184 -332 185 -331
rect 250 -332 251 -331
rect 254 -332 255 -331
rect 366 -332 367 -331
rect 401 -332 402 -331
rect 422 -332 423 -331
rect 82 -334 83 -333
rect 142 -334 143 -333
rect 212 -334 213 -333
rect 219 -334 220 -333
rect 243 -334 244 -333
rect 338 -334 339 -333
rect 72 -336 73 -335
rect 82 -336 83 -335
rect 86 -336 87 -335
rect 121 -336 122 -335
rect 124 -336 125 -335
rect 215 -336 216 -335
rect 250 -336 251 -335
rect 303 -336 304 -335
rect 100 -338 101 -337
rect 107 -338 108 -337
rect 110 -338 111 -337
rect 152 -338 153 -337
rect 163 -338 164 -337
rect 212 -338 213 -337
rect 261 -338 262 -337
rect 310 -338 311 -337
rect 114 -340 115 -339
rect 226 -340 227 -339
rect 264 -340 265 -339
rect 373 -340 374 -339
rect 44 -342 45 -341
rect 114 -342 115 -341
rect 117 -342 118 -341
rect 205 -342 206 -341
rect 264 -342 265 -341
rect 443 -342 444 -341
rect 128 -344 129 -343
rect 229 -344 230 -343
rect 268 -344 269 -343
rect 271 -344 272 -343
rect 285 -344 286 -343
rect 289 -344 290 -343
rect 299 -344 300 -343
rect 401 -344 402 -343
rect 131 -346 132 -345
rect 135 -346 136 -345
rect 194 -346 195 -345
rect 338 -346 339 -345
rect 233 -348 234 -347
rect 285 -348 286 -347
rect 289 -348 290 -347
rect 306 -348 307 -347
rect 310 -348 311 -347
rect 359 -348 360 -347
rect 170 -350 171 -349
rect 233 -350 234 -349
rect 352 -350 353 -349
rect 359 -350 360 -349
rect 345 -352 346 -351
rect 352 -352 353 -351
rect 345 -354 346 -353
rect 429 -354 430 -353
rect 394 -356 395 -355
rect 429 -356 430 -355
rect 240 -358 241 -357
rect 394 -358 395 -357
rect 240 -360 241 -359
rect 450 -360 451 -359
rect 23 -371 24 -370
rect 100 -371 101 -370
rect 121 -371 122 -370
rect 152 -371 153 -370
rect 198 -371 199 -370
rect 271 -371 272 -370
rect 275 -371 276 -370
rect 436 -371 437 -370
rect 443 -371 444 -370
rect 527 -371 528 -370
rect 30 -373 31 -372
rect 117 -373 118 -372
rect 135 -373 136 -372
rect 166 -373 167 -372
rect 226 -373 227 -372
rect 303 -373 304 -372
rect 317 -373 318 -372
rect 366 -373 367 -372
rect 387 -373 388 -372
rect 457 -373 458 -372
rect 481 -373 482 -372
rect 499 -373 500 -372
rect 30 -375 31 -374
rect 173 -375 174 -374
rect 226 -375 227 -374
rect 310 -375 311 -374
rect 331 -375 332 -374
rect 457 -375 458 -374
rect 37 -377 38 -376
rect 114 -377 115 -376
rect 128 -377 129 -376
rect 166 -377 167 -376
rect 233 -377 234 -376
rect 278 -377 279 -376
rect 282 -377 283 -376
rect 464 -377 465 -376
rect 44 -379 45 -378
rect 124 -379 125 -378
rect 138 -379 139 -378
rect 170 -379 171 -378
rect 233 -379 234 -378
rect 313 -379 314 -378
rect 338 -379 339 -378
rect 387 -379 388 -378
rect 390 -379 391 -378
rect 415 -379 416 -378
rect 418 -379 419 -378
rect 520 -379 521 -378
rect 44 -381 45 -380
rect 103 -381 104 -380
rect 149 -381 150 -380
rect 215 -381 216 -380
rect 240 -381 241 -380
rect 296 -381 297 -380
rect 310 -381 311 -380
rect 401 -381 402 -380
rect 415 -381 416 -380
rect 443 -381 444 -380
rect 450 -381 451 -380
rect 492 -381 493 -380
rect 51 -383 52 -382
rect 100 -383 101 -382
rect 243 -383 244 -382
rect 345 -383 346 -382
rect 348 -383 349 -382
rect 366 -383 367 -382
rect 394 -383 395 -382
rect 506 -383 507 -382
rect 58 -385 59 -384
rect 110 -385 111 -384
rect 254 -385 255 -384
rect 282 -385 283 -384
rect 296 -385 297 -384
rect 320 -385 321 -384
rect 352 -385 353 -384
rect 401 -385 402 -384
rect 408 -385 409 -384
rect 450 -385 451 -384
rect 58 -387 59 -386
rect 159 -387 160 -386
rect 254 -387 255 -386
rect 289 -387 290 -386
rect 352 -387 353 -386
rect 471 -387 472 -386
rect 65 -389 66 -388
rect 191 -389 192 -388
rect 250 -389 251 -388
rect 471 -389 472 -388
rect 65 -391 66 -390
rect 82 -391 83 -390
rect 86 -391 87 -390
rect 208 -391 209 -390
rect 261 -391 262 -390
rect 380 -391 381 -390
rect 408 -391 409 -390
rect 422 -391 423 -390
rect 72 -393 73 -392
rect 93 -393 94 -392
rect 110 -393 111 -392
rect 247 -393 248 -392
rect 261 -393 262 -392
rect 394 -393 395 -392
rect 72 -395 73 -394
rect 212 -395 213 -394
rect 268 -395 269 -394
rect 429 -395 430 -394
rect 79 -397 80 -396
rect 107 -397 108 -396
rect 131 -397 132 -396
rect 289 -397 290 -396
rect 324 -397 325 -396
rect 422 -397 423 -396
rect 37 -399 38 -398
rect 107 -399 108 -398
rect 114 -399 115 -398
rect 324 -399 325 -398
rect 359 -399 360 -398
rect 380 -399 381 -398
rect 89 -401 90 -400
rect 142 -401 143 -400
rect 156 -401 157 -400
rect 191 -401 192 -400
rect 212 -401 213 -400
rect 331 -401 332 -400
rect 373 -401 374 -400
rect 429 -401 430 -400
rect 93 -403 94 -402
rect 184 -403 185 -402
rect 229 -403 230 -402
rect 359 -403 360 -402
rect 156 -405 157 -404
rect 436 -405 437 -404
rect 177 -407 178 -406
rect 247 -407 248 -406
rect 275 -407 276 -406
rect 327 -407 328 -406
rect 177 -409 178 -408
rect 194 -409 195 -408
rect 240 -409 241 -408
rect 268 -409 269 -408
rect 317 -409 318 -408
rect 373 -409 374 -408
rect 184 -411 185 -410
rect 205 -411 206 -410
rect 16 -422 17 -421
rect 79 -422 80 -421
rect 86 -422 87 -421
rect 89 -422 90 -421
rect 93 -422 94 -421
rect 215 -422 216 -421
rect 247 -422 248 -421
rect 264 -422 265 -421
rect 268 -422 269 -421
rect 282 -422 283 -421
rect 289 -422 290 -421
rect 292 -422 293 -421
rect 324 -422 325 -421
rect 499 -422 500 -421
rect 520 -422 521 -421
rect 548 -422 549 -421
rect 30 -424 31 -423
rect 145 -424 146 -423
rect 159 -424 160 -423
rect 457 -424 458 -423
rect 464 -424 465 -423
rect 541 -424 542 -423
rect 30 -426 31 -425
rect 110 -426 111 -425
rect 114 -426 115 -425
rect 212 -426 213 -425
rect 219 -426 220 -425
rect 247 -426 248 -425
rect 254 -426 255 -425
rect 324 -426 325 -425
rect 327 -426 328 -425
rect 408 -426 409 -425
rect 415 -426 416 -425
rect 576 -426 577 -425
rect 44 -428 45 -427
rect 222 -428 223 -427
rect 240 -428 241 -427
rect 254 -428 255 -427
rect 261 -428 262 -427
rect 492 -428 493 -427
rect 527 -428 528 -427
rect 562 -428 563 -427
rect 2 -430 3 -429
rect 240 -430 241 -429
rect 278 -430 279 -429
rect 296 -430 297 -429
rect 338 -430 339 -429
rect 485 -430 486 -429
rect 51 -432 52 -431
rect 54 -432 55 -431
rect 58 -432 59 -431
rect 121 -432 122 -431
rect 128 -432 129 -431
rect 201 -432 202 -431
rect 219 -432 220 -431
rect 499 -432 500 -431
rect 37 -434 38 -433
rect 121 -434 122 -433
rect 135 -434 136 -433
rect 166 -434 167 -433
rect 173 -434 174 -433
rect 464 -434 465 -433
rect 471 -434 472 -433
rect 478 -434 479 -433
rect 65 -436 66 -435
rect 198 -436 199 -435
rect 226 -436 227 -435
rect 527 -436 528 -435
rect 72 -438 73 -437
rect 320 -438 321 -437
rect 341 -438 342 -437
rect 401 -438 402 -437
rect 429 -438 430 -437
rect 520 -438 521 -437
rect 72 -440 73 -439
rect 170 -440 171 -439
rect 191 -440 192 -439
rect 275 -440 276 -439
rect 285 -440 286 -439
rect 471 -440 472 -439
rect 9 -442 10 -441
rect 170 -442 171 -441
rect 177 -442 178 -441
rect 285 -442 286 -441
rect 289 -442 290 -441
rect 303 -442 304 -441
rect 348 -442 349 -441
rect 485 -442 486 -441
rect 79 -444 80 -443
rect 345 -444 346 -443
rect 352 -444 353 -443
rect 408 -444 409 -443
rect 436 -444 437 -443
rect 534 -444 535 -443
rect 86 -446 87 -445
rect 184 -446 185 -445
rect 198 -446 199 -445
rect 229 -446 230 -445
rect 296 -446 297 -445
rect 313 -446 314 -445
rect 359 -446 360 -445
rect 457 -446 458 -445
rect 96 -448 97 -447
rect 100 -448 101 -447
rect 107 -448 108 -447
rect 142 -448 143 -447
rect 177 -448 178 -447
rect 243 -448 244 -447
rect 366 -448 367 -447
rect 401 -448 402 -447
rect 436 -448 437 -447
rect 443 -448 444 -447
rect 142 -450 143 -449
rect 359 -450 360 -449
rect 380 -450 381 -449
rect 429 -450 430 -449
rect 443 -450 444 -449
rect 506 -450 507 -449
rect 23 -452 24 -451
rect 506 -452 507 -451
rect 205 -454 206 -453
rect 352 -454 353 -453
rect 373 -454 374 -453
rect 380 -454 381 -453
rect 387 -454 388 -453
rect 492 -454 493 -453
rect 229 -456 230 -455
rect 415 -456 416 -455
rect 275 -458 276 -457
rect 387 -458 388 -457
rect 394 -458 395 -457
rect 397 -458 398 -457
rect 394 -460 395 -459
rect 422 -460 423 -459
rect 397 -462 398 -461
rect 422 -462 423 -461
rect 9 -473 10 -472
rect 121 -473 122 -472
rect 131 -473 132 -472
rect 191 -473 192 -472
rect 219 -473 220 -472
rect 247 -473 248 -472
rect 275 -473 276 -472
rect 471 -473 472 -472
rect 555 -473 556 -472
rect 562 -473 563 -472
rect 16 -475 17 -474
rect 117 -475 118 -474
rect 152 -475 153 -474
rect 177 -475 178 -474
rect 184 -475 185 -474
rect 313 -475 314 -474
rect 355 -475 356 -474
rect 534 -475 535 -474
rect 558 -475 559 -474
rect 562 -475 563 -474
rect 16 -477 17 -476
rect 93 -477 94 -476
rect 107 -477 108 -476
rect 278 -477 279 -476
rect 282 -477 283 -476
rect 471 -477 472 -476
rect 23 -479 24 -478
rect 149 -479 150 -478
rect 159 -479 160 -478
rect 422 -479 423 -478
rect 425 -479 426 -478
rect 485 -479 486 -478
rect 30 -481 31 -480
rect 54 -481 55 -480
rect 58 -481 59 -480
rect 96 -481 97 -480
rect 107 -481 108 -480
rect 233 -481 234 -480
rect 240 -481 241 -480
rect 338 -481 339 -480
rect 359 -481 360 -480
rect 541 -481 542 -480
rect 37 -483 38 -482
rect 240 -483 241 -482
rect 285 -483 286 -482
rect 408 -483 409 -482
rect 464 -483 465 -482
rect 572 -483 573 -482
rect 2 -485 3 -484
rect 285 -485 286 -484
rect 299 -485 300 -484
rect 359 -485 360 -484
rect 373 -485 374 -484
rect 457 -485 458 -484
rect 541 -485 542 -484
rect 548 -485 549 -484
rect 37 -487 38 -486
rect 114 -487 115 -486
rect 142 -487 143 -486
rect 149 -487 150 -486
rect 163 -487 164 -486
rect 506 -487 507 -486
rect 44 -489 45 -488
rect 124 -489 125 -488
rect 135 -489 136 -488
rect 163 -489 164 -488
rect 170 -489 171 -488
rect 177 -489 178 -488
rect 184 -489 185 -488
rect 268 -489 269 -488
rect 303 -489 304 -488
rect 317 -489 318 -488
rect 331 -489 332 -488
rect 338 -489 339 -488
rect 394 -489 395 -488
rect 485 -489 486 -488
rect 51 -491 52 -490
rect 345 -491 346 -490
rect 380 -491 381 -490
rect 394 -491 395 -490
rect 408 -491 409 -490
rect 415 -491 416 -490
rect 436 -491 437 -490
rect 464 -491 465 -490
rect 72 -493 73 -492
rect 229 -493 230 -492
rect 233 -493 234 -492
rect 369 -493 370 -492
rect 380 -493 381 -492
rect 401 -493 402 -492
rect 457 -493 458 -492
rect 499 -493 500 -492
rect 44 -495 45 -494
rect 229 -495 230 -494
rect 289 -495 290 -494
rect 303 -495 304 -494
rect 310 -495 311 -494
rect 527 -495 528 -494
rect 75 -497 76 -496
rect 93 -497 94 -496
rect 124 -497 125 -496
rect 219 -497 220 -496
rect 222 -497 223 -496
rect 576 -497 577 -496
rect 86 -499 87 -498
rect 264 -499 265 -498
rect 289 -499 290 -498
rect 296 -499 297 -498
rect 310 -499 311 -498
rect 324 -499 325 -498
rect 331 -499 332 -498
rect 450 -499 451 -498
rect 82 -501 83 -500
rect 86 -501 87 -500
rect 89 -501 90 -500
rect 128 -501 129 -500
rect 156 -501 157 -500
rect 415 -501 416 -500
rect 429 -501 430 -500
rect 450 -501 451 -500
rect 170 -503 171 -502
rect 243 -503 244 -502
rect 264 -503 265 -502
rect 268 -503 269 -502
rect 296 -503 297 -502
rect 492 -503 493 -502
rect 191 -505 192 -504
rect 261 -505 262 -504
rect 320 -505 321 -504
rect 401 -505 402 -504
rect 429 -505 430 -504
rect 443 -505 444 -504
rect 478 -505 479 -504
rect 492 -505 493 -504
rect 65 -507 66 -506
rect 261 -507 262 -506
rect 282 -507 283 -506
rect 478 -507 479 -506
rect 58 -509 59 -508
rect 65 -509 66 -508
rect 201 -509 202 -508
rect 247 -509 248 -508
rect 292 -509 293 -508
rect 443 -509 444 -508
rect 201 -511 202 -510
rect 509 -511 510 -510
rect 212 -513 213 -512
rect 317 -513 318 -512
rect 366 -513 367 -512
rect 436 -513 437 -512
rect 205 -515 206 -514
rect 212 -515 213 -514
rect 226 -515 227 -514
rect 254 -515 255 -514
rect 366 -515 367 -514
rect 520 -515 521 -514
rect 79 -517 80 -516
rect 205 -517 206 -516
rect 387 -517 388 -516
rect 520 -517 521 -516
rect 23 -519 24 -518
rect 79 -519 80 -518
rect 390 -519 391 -518
rect 499 -519 500 -518
rect 9 -530 10 -529
rect 16 -530 17 -529
rect 23 -530 24 -529
rect 128 -530 129 -529
rect 131 -530 132 -529
rect 170 -530 171 -529
rect 177 -530 178 -529
rect 187 -530 188 -529
rect 198 -530 199 -529
rect 212 -530 213 -529
rect 215 -530 216 -529
rect 219 -530 220 -529
rect 226 -530 227 -529
rect 499 -530 500 -529
rect 509 -530 510 -529
rect 555 -530 556 -529
rect 16 -532 17 -531
rect 257 -532 258 -531
rect 268 -532 269 -531
rect 271 -532 272 -531
rect 275 -532 276 -531
rect 369 -532 370 -531
rect 373 -532 374 -531
rect 527 -532 528 -531
rect 30 -534 31 -533
rect 68 -534 69 -533
rect 79 -534 80 -533
rect 100 -534 101 -533
rect 107 -534 108 -533
rect 177 -534 178 -533
rect 205 -534 206 -533
rect 292 -534 293 -533
rect 296 -534 297 -533
rect 317 -534 318 -533
rect 331 -534 332 -533
rect 366 -534 367 -533
rect 373 -534 374 -533
rect 520 -534 521 -533
rect 30 -536 31 -535
rect 68 -536 69 -535
rect 103 -536 104 -535
rect 205 -536 206 -535
rect 219 -536 220 -535
rect 513 -536 514 -535
rect 37 -538 38 -537
rect 201 -538 202 -537
rect 254 -538 255 -537
rect 299 -538 300 -537
rect 306 -538 307 -537
rect 408 -538 409 -537
rect 478 -538 479 -537
rect 534 -538 535 -537
rect 40 -540 41 -539
rect 89 -540 90 -539
rect 107 -540 108 -539
rect 163 -540 164 -539
rect 254 -540 255 -539
rect 387 -540 388 -539
rect 464 -540 465 -539
rect 478 -540 479 -539
rect 485 -540 486 -539
rect 506 -540 507 -539
rect 44 -542 45 -541
rect 138 -542 139 -541
rect 156 -542 157 -541
rect 285 -542 286 -541
rect 289 -542 290 -541
rect 376 -542 377 -541
rect 492 -542 493 -541
rect 520 -542 521 -541
rect 51 -544 52 -543
rect 184 -544 185 -543
rect 208 -544 209 -543
rect 506 -544 507 -543
rect 51 -546 52 -545
rect 75 -546 76 -545
rect 114 -546 115 -545
rect 261 -546 262 -545
rect 268 -546 269 -545
rect 303 -546 304 -545
rect 313 -546 314 -545
rect 422 -546 423 -545
rect 492 -546 493 -545
rect 530 -546 531 -545
rect 58 -548 59 -547
rect 121 -548 122 -547
rect 124 -548 125 -547
rect 145 -548 146 -547
rect 149 -548 150 -547
rect 156 -548 157 -547
rect 163 -548 164 -547
rect 278 -548 279 -547
rect 282 -548 283 -547
rect 471 -548 472 -547
rect 58 -550 59 -549
rect 72 -550 73 -549
rect 117 -550 118 -549
rect 310 -550 311 -549
rect 313 -550 314 -549
rect 443 -550 444 -549
rect 121 -552 122 -551
rect 222 -552 223 -551
rect 317 -552 318 -551
rect 324 -552 325 -551
rect 331 -552 332 -551
rect 341 -552 342 -551
rect 345 -552 346 -551
rect 450 -552 451 -551
rect 128 -554 129 -553
rect 170 -554 171 -553
rect 229 -554 230 -553
rect 324 -554 325 -553
rect 348 -554 349 -553
rect 436 -554 437 -553
rect 443 -554 444 -553
rect 457 -554 458 -553
rect 135 -556 136 -555
rect 233 -556 234 -555
rect 240 -556 241 -555
rect 436 -556 437 -555
rect 149 -558 150 -557
rect 191 -558 192 -557
rect 240 -558 241 -557
rect 261 -558 262 -557
rect 352 -558 353 -557
rect 471 -558 472 -557
rect 159 -560 160 -559
rect 191 -560 192 -559
rect 338 -560 339 -559
rect 352 -560 353 -559
rect 359 -560 360 -559
rect 408 -560 409 -559
rect 415 -560 416 -559
rect 450 -560 451 -559
rect 142 -562 143 -561
rect 359 -562 360 -561
rect 362 -562 363 -561
rect 464 -562 465 -561
rect 236 -564 237 -563
rect 338 -564 339 -563
rect 394 -564 395 -563
rect 415 -564 416 -563
rect 429 -564 430 -563
rect 457 -564 458 -563
rect 394 -566 395 -565
rect 401 -566 402 -565
rect 429 -566 430 -565
rect 485 -566 486 -565
rect 264 -568 265 -567
rect 401 -568 402 -567
rect 9 -579 10 -578
rect 89 -579 90 -578
rect 121 -579 122 -578
rect 282 -579 283 -578
rect 289 -579 290 -578
rect 303 -579 304 -578
rect 338 -579 339 -578
rect 394 -579 395 -578
rect 429 -579 430 -578
rect 450 -579 451 -578
rect 464 -579 465 -578
rect 527 -579 528 -578
rect 530 -579 531 -578
rect 541 -579 542 -578
rect 9 -581 10 -580
rect 110 -581 111 -580
rect 121 -581 122 -580
rect 131 -581 132 -580
rect 135 -581 136 -580
rect 212 -581 213 -580
rect 222 -581 223 -580
rect 331 -581 332 -580
rect 338 -581 339 -580
rect 345 -581 346 -580
rect 359 -581 360 -580
rect 415 -581 416 -580
rect 432 -581 433 -580
rect 520 -581 521 -580
rect 534 -581 535 -580
rect 548 -581 549 -580
rect 23 -583 24 -582
rect 58 -583 59 -582
rect 72 -583 73 -582
rect 82 -583 83 -582
rect 86 -583 87 -582
rect 226 -583 227 -582
rect 233 -583 234 -582
rect 247 -583 248 -582
rect 254 -583 255 -582
rect 275 -583 276 -582
rect 324 -583 325 -582
rect 331 -583 332 -582
rect 341 -583 342 -582
rect 345 -583 346 -582
rect 352 -583 353 -582
rect 359 -583 360 -582
rect 366 -583 367 -582
rect 380 -583 381 -582
rect 436 -583 437 -582
rect 499 -583 500 -582
rect 520 -583 521 -582
rect 541 -583 542 -582
rect 23 -585 24 -584
rect 100 -585 101 -584
rect 135 -585 136 -584
rect 362 -585 363 -584
rect 380 -585 381 -584
rect 387 -585 388 -584
rect 436 -585 437 -584
rect 509 -585 510 -584
rect 523 -585 524 -584
rect 534 -585 535 -584
rect 30 -587 31 -586
rect 114 -587 115 -586
rect 138 -587 139 -586
rect 163 -587 164 -586
rect 170 -587 171 -586
rect 187 -587 188 -586
rect 191 -587 192 -586
rect 219 -587 220 -586
rect 236 -587 237 -586
rect 516 -587 517 -586
rect 30 -589 31 -588
rect 51 -589 52 -588
rect 54 -589 55 -588
rect 65 -589 66 -588
rect 72 -589 73 -588
rect 128 -589 129 -588
rect 145 -589 146 -588
rect 156 -589 157 -588
rect 191 -589 192 -588
rect 285 -589 286 -588
rect 352 -589 353 -588
rect 548 -589 549 -588
rect 16 -591 17 -590
rect 51 -591 52 -590
rect 58 -591 59 -590
rect 65 -591 66 -590
rect 79 -591 80 -590
rect 117 -591 118 -590
rect 142 -591 143 -590
rect 156 -591 157 -590
rect 198 -591 199 -590
rect 229 -591 230 -590
rect 240 -591 241 -590
rect 394 -591 395 -590
rect 443 -591 444 -590
rect 464 -591 465 -590
rect 471 -591 472 -590
rect 527 -591 528 -590
rect 37 -593 38 -592
rect 44 -593 45 -592
rect 79 -593 80 -592
rect 107 -593 108 -592
rect 149 -593 150 -592
rect 173 -593 174 -592
rect 198 -593 199 -592
rect 271 -593 272 -592
rect 275 -593 276 -592
rect 317 -593 318 -592
rect 387 -593 388 -592
rect 422 -593 423 -592
rect 443 -593 444 -592
rect 457 -593 458 -592
rect 481 -593 482 -592
rect 506 -593 507 -592
rect 103 -595 104 -594
rect 163 -595 164 -594
rect 205 -595 206 -594
rect 296 -595 297 -594
rect 373 -595 374 -594
rect 457 -595 458 -594
rect 485 -595 486 -594
rect 513 -595 514 -594
rect 142 -597 143 -596
rect 373 -597 374 -596
rect 401 -597 402 -596
rect 471 -597 472 -596
rect 485 -597 486 -596
rect 492 -597 493 -596
rect 499 -597 500 -596
rect 513 -597 514 -596
rect 149 -599 150 -598
rect 310 -599 311 -598
rect 450 -599 451 -598
rect 478 -599 479 -598
rect 205 -601 206 -600
rect 327 -601 328 -600
rect 208 -603 209 -602
rect 233 -603 234 -602
rect 247 -603 248 -602
rect 261 -603 262 -602
rect 268 -603 269 -602
rect 492 -603 493 -602
rect 177 -605 178 -604
rect 268 -605 269 -604
rect 289 -605 290 -604
rect 422 -605 423 -604
rect 219 -607 220 -606
rect 299 -607 300 -606
rect 306 -607 307 -606
rect 401 -607 402 -606
rect 229 -609 230 -608
rect 317 -609 318 -608
rect 261 -611 262 -610
rect 313 -611 314 -610
rect 9 -622 10 -621
rect 68 -622 69 -621
rect 72 -622 73 -621
rect 131 -622 132 -621
rect 142 -622 143 -621
rect 226 -622 227 -621
rect 233 -622 234 -621
rect 292 -622 293 -621
rect 296 -622 297 -621
rect 380 -622 381 -621
rect 394 -622 395 -621
rect 436 -622 437 -621
rect 443 -622 444 -621
rect 474 -622 475 -621
rect 499 -622 500 -621
rect 506 -622 507 -621
rect 513 -622 514 -621
rect 583 -622 584 -621
rect 16 -624 17 -623
rect 61 -624 62 -623
rect 65 -624 66 -623
rect 117 -624 118 -623
rect 163 -624 164 -623
rect 177 -624 178 -623
rect 184 -624 185 -623
rect 198 -624 199 -623
rect 219 -624 220 -623
rect 247 -624 248 -623
rect 261 -624 262 -623
rect 418 -624 419 -623
rect 422 -624 423 -623
rect 436 -624 437 -623
rect 450 -624 451 -623
rect 488 -624 489 -623
rect 516 -624 517 -623
rect 534 -624 535 -623
rect 544 -624 545 -623
rect 555 -624 556 -623
rect 23 -626 24 -625
rect 89 -626 90 -625
rect 93 -626 94 -625
rect 100 -626 101 -625
rect 103 -626 104 -625
rect 299 -626 300 -625
rect 310 -626 311 -625
rect 359 -626 360 -625
rect 401 -626 402 -625
rect 443 -626 444 -625
rect 520 -626 521 -625
rect 541 -626 542 -625
rect 555 -626 556 -625
rect 562 -626 563 -625
rect 30 -628 31 -627
rect 47 -628 48 -627
rect 51 -628 52 -627
rect 58 -628 59 -627
rect 72 -628 73 -627
rect 79 -628 80 -627
rect 96 -628 97 -627
rect 208 -628 209 -627
rect 222 -628 223 -627
rect 261 -628 262 -627
rect 275 -628 276 -627
rect 310 -628 311 -627
rect 317 -628 318 -627
rect 450 -628 451 -627
rect 527 -628 528 -627
rect 534 -628 535 -627
rect 37 -630 38 -629
rect 44 -630 45 -629
rect 107 -630 108 -629
rect 135 -630 136 -629
rect 149 -630 150 -629
rect 177 -630 178 -629
rect 226 -630 227 -629
rect 303 -630 304 -629
rect 327 -630 328 -629
rect 429 -630 430 -629
rect 44 -632 45 -631
rect 320 -632 321 -631
rect 334 -632 335 -631
rect 387 -632 388 -631
rect 397 -632 398 -631
rect 429 -632 430 -631
rect 86 -634 87 -633
rect 107 -634 108 -633
rect 114 -634 115 -633
rect 219 -634 220 -633
rect 233 -634 234 -633
rect 250 -634 251 -633
rect 275 -634 276 -633
rect 348 -634 349 -633
rect 352 -634 353 -633
rect 457 -634 458 -633
rect 75 -636 76 -635
rect 86 -636 87 -635
rect 114 -636 115 -635
rect 247 -636 248 -635
rect 296 -636 297 -635
rect 373 -636 374 -635
rect 380 -636 381 -635
rect 397 -636 398 -635
rect 408 -636 409 -635
rect 415 -636 416 -635
rect 422 -636 423 -635
rect 471 -636 472 -635
rect 131 -638 132 -637
rect 359 -638 360 -637
rect 366 -638 367 -637
rect 471 -638 472 -637
rect 149 -640 150 -639
rect 156 -640 157 -639
rect 163 -640 164 -639
rect 212 -640 213 -639
rect 240 -640 241 -639
rect 289 -640 290 -639
rect 324 -640 325 -639
rect 457 -640 458 -639
rect 128 -642 129 -641
rect 156 -642 157 -641
rect 170 -642 171 -641
rect 187 -642 188 -641
rect 191 -642 192 -641
rect 303 -642 304 -641
rect 324 -642 325 -641
rect 530 -642 531 -641
rect 40 -644 41 -643
rect 170 -644 171 -643
rect 180 -644 181 -643
rect 191 -644 192 -643
rect 205 -644 206 -643
rect 212 -644 213 -643
rect 254 -644 255 -643
rect 289 -644 290 -643
rect 331 -644 332 -643
rect 366 -644 367 -643
rect 401 -644 402 -643
rect 408 -644 409 -643
rect 254 -646 255 -645
rect 548 -646 549 -645
rect 331 -648 332 -647
rect 387 -648 388 -647
rect 481 -648 482 -647
rect 548 -648 549 -647
rect 338 -650 339 -649
rect 478 -650 479 -649
rect 341 -652 342 -651
rect 499 -652 500 -651
rect 268 -654 269 -653
rect 341 -654 342 -653
rect 345 -654 346 -653
rect 352 -654 353 -653
rect 355 -654 356 -653
rect 492 -654 493 -653
rect 345 -656 346 -655
rect 464 -656 465 -655
rect 485 -656 486 -655
rect 492 -656 493 -655
rect 464 -658 465 -657
rect 516 -658 517 -657
rect 16 -669 17 -668
rect 65 -669 66 -668
rect 107 -669 108 -668
rect 110 -669 111 -668
rect 114 -669 115 -668
rect 135 -669 136 -668
rect 156 -669 157 -668
rect 271 -669 272 -668
rect 296 -669 297 -668
rect 317 -669 318 -668
rect 320 -669 321 -668
rect 429 -669 430 -668
rect 471 -669 472 -668
rect 618 -669 619 -668
rect 628 -669 629 -668
rect 639 -669 640 -668
rect 23 -671 24 -670
rect 103 -671 104 -670
rect 156 -671 157 -670
rect 177 -671 178 -670
rect 205 -671 206 -670
rect 212 -671 213 -670
rect 240 -671 241 -670
rect 289 -671 290 -670
rect 303 -671 304 -670
rect 404 -671 405 -670
rect 471 -671 472 -670
rect 478 -671 479 -670
rect 485 -671 486 -670
rect 488 -671 489 -670
rect 499 -671 500 -670
rect 513 -671 514 -670
rect 516 -671 517 -670
rect 520 -671 521 -670
rect 527 -671 528 -670
rect 611 -671 612 -670
rect 30 -673 31 -672
rect 37 -673 38 -672
rect 44 -673 45 -672
rect 100 -673 101 -672
rect 163 -673 164 -672
rect 166 -673 167 -672
rect 170 -673 171 -672
rect 233 -673 234 -672
rect 247 -673 248 -672
rect 303 -673 304 -672
rect 345 -673 346 -672
rect 576 -673 577 -672
rect 583 -673 584 -672
rect 646 -673 647 -672
rect 44 -675 45 -674
rect 51 -675 52 -674
rect 58 -675 59 -674
rect 79 -675 80 -674
rect 93 -675 94 -674
rect 103 -675 104 -674
rect 114 -675 115 -674
rect 163 -675 164 -674
rect 170 -675 171 -674
rect 226 -675 227 -674
rect 247 -675 248 -674
rect 299 -675 300 -674
rect 348 -675 349 -674
rect 366 -675 367 -674
rect 376 -675 377 -674
rect 415 -675 416 -674
rect 478 -675 479 -674
rect 492 -675 493 -674
rect 499 -675 500 -674
rect 555 -675 556 -674
rect 593 -675 594 -674
rect 632 -675 633 -674
rect 51 -677 52 -676
rect 334 -677 335 -676
rect 352 -677 353 -676
rect 373 -677 374 -676
rect 380 -677 381 -676
rect 401 -677 402 -676
rect 415 -677 416 -676
rect 457 -677 458 -676
rect 506 -677 507 -676
rect 520 -677 521 -676
rect 530 -677 531 -676
rect 534 -677 535 -676
rect 548 -677 549 -676
rect 562 -677 563 -676
rect 65 -679 66 -678
rect 86 -679 87 -678
rect 191 -679 192 -678
rect 226 -679 227 -678
rect 250 -679 251 -678
rect 464 -679 465 -678
rect 72 -681 73 -680
rect 79 -681 80 -680
rect 86 -681 87 -680
rect 121 -681 122 -680
rect 201 -681 202 -680
rect 205 -681 206 -680
rect 212 -681 213 -680
rect 275 -681 276 -680
rect 296 -681 297 -680
rect 555 -681 556 -680
rect 121 -683 122 -682
rect 198 -683 199 -682
rect 219 -683 220 -682
rect 275 -683 276 -682
rect 324 -683 325 -682
rect 373 -683 374 -682
rect 380 -683 381 -682
rect 604 -683 605 -682
rect 177 -685 178 -684
rect 201 -685 202 -684
rect 219 -685 220 -684
rect 243 -685 244 -684
rect 254 -685 255 -684
rect 324 -685 325 -684
rect 331 -685 332 -684
rect 534 -685 535 -684
rect 184 -687 185 -686
rect 254 -687 255 -686
rect 261 -687 262 -686
rect 289 -687 290 -686
rect 338 -687 339 -686
rect 506 -687 507 -686
rect 135 -689 136 -688
rect 261 -689 262 -688
rect 268 -689 269 -688
rect 548 -689 549 -688
rect 149 -691 150 -690
rect 184 -691 185 -690
rect 194 -691 195 -690
rect 268 -691 269 -690
rect 310 -691 311 -690
rect 338 -691 339 -690
rect 359 -691 360 -690
rect 401 -691 402 -690
rect 443 -691 444 -690
rect 457 -691 458 -690
rect 128 -693 129 -692
rect 149 -693 150 -692
rect 233 -693 234 -692
rect 310 -693 311 -692
rect 366 -693 367 -692
rect 408 -693 409 -692
rect 443 -693 444 -692
rect 544 -693 545 -692
rect 282 -695 283 -694
rect 359 -695 360 -694
rect 387 -695 388 -694
rect 583 -695 584 -694
rect 387 -697 388 -696
rect 436 -697 437 -696
rect 450 -697 451 -696
rect 464 -697 465 -696
rect 345 -699 346 -698
rect 436 -699 437 -698
rect 450 -699 451 -698
rect 572 -699 573 -698
rect 394 -701 395 -700
rect 429 -701 430 -700
rect 397 -703 398 -702
rect 422 -703 423 -702
rect 408 -705 409 -704
rect 474 -705 475 -704
rect 422 -707 423 -706
rect 541 -707 542 -706
rect 16 -718 17 -717
rect 58 -718 59 -717
rect 86 -718 87 -717
rect 135 -718 136 -717
rect 142 -718 143 -717
rect 149 -718 150 -717
rect 152 -718 153 -717
rect 187 -718 188 -717
rect 194 -718 195 -717
rect 205 -718 206 -717
rect 219 -718 220 -717
rect 254 -718 255 -717
rect 261 -718 262 -717
rect 345 -718 346 -717
rect 348 -718 349 -717
rect 415 -718 416 -717
rect 422 -718 423 -717
rect 488 -718 489 -717
rect 495 -718 496 -717
rect 534 -718 535 -717
rect 541 -718 542 -717
rect 614 -718 615 -717
rect 23 -720 24 -719
rect 65 -720 66 -719
rect 79 -720 80 -719
rect 149 -720 150 -719
rect 156 -720 157 -719
rect 261 -720 262 -719
rect 268 -720 269 -719
rect 331 -720 332 -719
rect 334 -720 335 -719
rect 471 -720 472 -719
rect 474 -720 475 -719
rect 534 -720 535 -719
rect 562 -720 563 -719
rect 600 -720 601 -719
rect 611 -720 612 -719
rect 632 -720 633 -719
rect 33 -722 34 -721
rect 37 -722 38 -721
rect 44 -722 45 -721
rect 75 -722 76 -721
rect 79 -722 80 -721
rect 114 -722 115 -721
rect 156 -722 157 -721
rect 285 -722 286 -721
rect 296 -722 297 -721
rect 324 -722 325 -721
rect 338 -722 339 -721
rect 464 -722 465 -721
rect 499 -722 500 -721
rect 572 -722 573 -721
rect 593 -722 594 -721
rect 646 -722 647 -721
rect 44 -724 45 -723
rect 121 -724 122 -723
rect 163 -724 164 -723
rect 177 -724 178 -723
rect 194 -724 195 -723
rect 303 -724 304 -723
rect 310 -724 311 -723
rect 506 -724 507 -723
rect 527 -724 528 -723
rect 530 -724 531 -723
rect 569 -724 570 -723
rect 604 -724 605 -723
rect 51 -726 52 -725
rect 257 -726 258 -725
rect 268 -726 269 -725
rect 289 -726 290 -725
rect 310 -726 311 -725
rect 359 -726 360 -725
rect 366 -726 367 -725
rect 527 -726 528 -725
rect 597 -726 598 -725
rect 639 -726 640 -725
rect 51 -728 52 -727
rect 128 -728 129 -727
rect 163 -728 164 -727
rect 229 -728 230 -727
rect 240 -728 241 -727
rect 303 -728 304 -727
rect 317 -728 318 -727
rect 324 -728 325 -727
rect 352 -728 353 -727
rect 541 -728 542 -727
rect 65 -730 66 -729
rect 72 -730 73 -729
rect 86 -730 87 -729
rect 93 -730 94 -729
rect 103 -730 104 -729
rect 457 -730 458 -729
rect 464 -730 465 -729
rect 555 -730 556 -729
rect 58 -732 59 -731
rect 103 -732 104 -731
rect 114 -732 115 -731
rect 128 -732 129 -731
rect 170 -732 171 -731
rect 201 -732 202 -731
rect 205 -732 206 -731
rect 296 -732 297 -731
rect 317 -732 318 -731
rect 331 -732 332 -731
rect 352 -732 353 -731
rect 359 -732 360 -731
rect 366 -732 367 -731
rect 513 -732 514 -731
rect 555 -732 556 -731
rect 618 -732 619 -731
rect 72 -734 73 -733
rect 107 -734 108 -733
rect 121 -734 122 -733
rect 215 -734 216 -733
rect 226 -734 227 -733
rect 240 -734 241 -733
rect 247 -734 248 -733
rect 383 -734 384 -733
rect 397 -734 398 -733
rect 520 -734 521 -733
rect 93 -736 94 -735
rect 152 -736 153 -735
rect 170 -736 171 -735
rect 212 -736 213 -735
rect 250 -736 251 -735
rect 387 -736 388 -735
rect 408 -736 409 -735
rect 520 -736 521 -735
rect 107 -738 108 -737
rect 198 -738 199 -737
rect 222 -738 223 -737
rect 387 -738 388 -737
rect 408 -738 409 -737
rect 443 -738 444 -737
rect 450 -738 451 -737
rect 457 -738 458 -737
rect 506 -738 507 -737
rect 576 -738 577 -737
rect 177 -740 178 -739
rect 191 -740 192 -739
rect 222 -740 223 -739
rect 362 -740 363 -739
rect 373 -740 374 -739
rect 492 -740 493 -739
rect 184 -742 185 -741
rect 198 -742 199 -741
rect 254 -742 255 -741
rect 348 -742 349 -741
rect 380 -742 381 -741
rect 478 -742 479 -741
rect 142 -744 143 -743
rect 184 -744 185 -743
rect 275 -744 276 -743
rect 278 -744 279 -743
rect 282 -744 283 -743
rect 401 -744 402 -743
rect 415 -744 416 -743
rect 471 -744 472 -743
rect 478 -744 479 -743
rect 548 -744 549 -743
rect 292 -746 293 -745
rect 401 -746 402 -745
rect 425 -746 426 -745
rect 583 -746 584 -745
rect 334 -748 335 -747
rect 513 -748 514 -747
rect 338 -750 339 -749
rect 450 -750 451 -749
rect 380 -752 381 -751
rect 436 -752 437 -751
rect 429 -754 430 -753
rect 499 -754 500 -753
rect 394 -756 395 -755
rect 429 -756 430 -755
rect 394 -758 395 -757
rect 436 -758 437 -757
rect 26 -769 27 -768
rect 33 -769 34 -768
rect 40 -769 41 -768
rect 149 -769 150 -768
rect 152 -769 153 -768
rect 373 -769 374 -768
rect 387 -769 388 -768
rect 394 -769 395 -768
rect 397 -769 398 -768
rect 457 -769 458 -768
rect 471 -769 472 -768
rect 520 -769 521 -768
rect 534 -769 535 -768
rect 558 -769 559 -768
rect 30 -771 31 -770
rect 37 -771 38 -770
rect 44 -771 45 -770
rect 114 -771 115 -770
rect 128 -771 129 -770
rect 166 -771 167 -770
rect 170 -771 171 -770
rect 191 -771 192 -770
rect 212 -771 213 -770
rect 268 -771 269 -770
rect 275 -771 276 -770
rect 436 -771 437 -770
rect 446 -771 447 -770
rect 478 -771 479 -770
rect 492 -771 493 -770
rect 527 -771 528 -770
rect 44 -773 45 -772
rect 93 -773 94 -772
rect 128 -773 129 -772
rect 187 -773 188 -772
rect 212 -773 213 -772
rect 310 -773 311 -772
rect 324 -773 325 -772
rect 338 -773 339 -772
rect 352 -773 353 -772
rect 460 -773 461 -772
rect 513 -773 514 -772
rect 548 -773 549 -772
rect 51 -775 52 -774
rect 145 -775 146 -774
rect 156 -775 157 -774
rect 194 -775 195 -774
rect 219 -775 220 -774
rect 261 -775 262 -774
rect 285 -775 286 -774
rect 317 -775 318 -774
rect 334 -775 335 -774
rect 485 -775 486 -774
rect 499 -775 500 -774
rect 513 -775 514 -774
rect 520 -775 521 -774
rect 555 -775 556 -774
rect 51 -777 52 -776
rect 121 -777 122 -776
rect 156 -777 157 -776
rect 191 -777 192 -776
rect 222 -777 223 -776
rect 289 -777 290 -776
rect 292 -777 293 -776
rect 376 -777 377 -776
rect 401 -777 402 -776
rect 499 -777 500 -776
rect 58 -779 59 -778
rect 142 -779 143 -778
rect 163 -779 164 -778
rect 331 -779 332 -778
rect 338 -779 339 -778
rect 443 -779 444 -778
rect 492 -779 493 -778
rect 555 -779 556 -778
rect 58 -781 59 -780
rect 65 -781 66 -780
rect 72 -781 73 -780
rect 152 -781 153 -780
rect 163 -781 164 -780
rect 282 -781 283 -780
rect 303 -781 304 -780
rect 387 -781 388 -780
rect 429 -781 430 -780
rect 534 -781 535 -780
rect 65 -783 66 -782
rect 331 -783 332 -782
rect 359 -783 360 -782
rect 464 -783 465 -782
rect 72 -785 73 -784
rect 145 -785 146 -784
rect 170 -785 171 -784
rect 257 -785 258 -784
rect 261 -785 262 -784
rect 422 -785 423 -784
rect 443 -785 444 -784
rect 530 -785 531 -784
rect 86 -787 87 -786
rect 117 -787 118 -786
rect 121 -787 122 -786
rect 436 -787 437 -786
rect 464 -787 465 -786
rect 506 -787 507 -786
rect 86 -789 87 -788
rect 205 -789 206 -788
rect 226 -789 227 -788
rect 275 -789 276 -788
rect 303 -789 304 -788
rect 352 -789 353 -788
rect 359 -789 360 -788
rect 380 -789 381 -788
rect 404 -789 405 -788
rect 429 -789 430 -788
rect 93 -791 94 -790
rect 257 -791 258 -790
rect 306 -791 307 -790
rect 478 -791 479 -790
rect 177 -793 178 -792
rect 324 -793 325 -792
rect 103 -795 104 -794
rect 177 -795 178 -794
rect 184 -795 185 -794
rect 226 -795 227 -794
rect 229 -795 230 -794
rect 366 -795 367 -794
rect 205 -797 206 -796
rect 215 -797 216 -796
rect 233 -797 234 -796
rect 268 -797 269 -796
rect 313 -797 314 -796
rect 506 -797 507 -796
rect 215 -799 216 -798
rect 219 -799 220 -798
rect 236 -799 237 -798
rect 341 -799 342 -798
rect 366 -799 367 -798
rect 408 -799 409 -798
rect 247 -801 248 -800
rect 296 -801 297 -800
rect 317 -801 318 -800
rect 471 -801 472 -800
rect 247 -803 248 -802
rect 422 -803 423 -802
rect 254 -805 255 -804
rect 541 -805 542 -804
rect 296 -807 297 -806
rect 380 -807 381 -806
rect 450 -807 451 -806
rect 541 -807 542 -806
rect 376 -809 377 -808
rect 408 -809 409 -808
rect 415 -809 416 -808
rect 450 -809 451 -808
rect 107 -811 108 -810
rect 415 -811 416 -810
rect 79 -813 80 -812
rect 107 -813 108 -812
rect 79 -815 80 -814
rect 198 -815 199 -814
rect 26 -826 27 -825
rect 40 -826 41 -825
rect 44 -826 45 -825
rect 236 -826 237 -825
rect 240 -826 241 -825
rect 247 -826 248 -825
rect 254 -826 255 -825
rect 285 -826 286 -825
rect 306 -826 307 -825
rect 485 -826 486 -825
rect 30 -828 31 -827
rect 37 -828 38 -827
rect 44 -828 45 -827
rect 72 -828 73 -827
rect 75 -828 76 -827
rect 110 -828 111 -827
rect 114 -828 115 -827
rect 142 -828 143 -827
rect 145 -828 146 -827
rect 317 -828 318 -827
rect 320 -828 321 -827
rect 387 -828 388 -827
rect 401 -828 402 -827
rect 464 -828 465 -827
rect 467 -828 468 -827
rect 541 -828 542 -827
rect 51 -830 52 -829
rect 159 -830 160 -829
rect 173 -830 174 -829
rect 194 -830 195 -829
rect 201 -830 202 -829
rect 404 -830 405 -829
rect 450 -830 451 -829
rect 485 -830 486 -829
rect 37 -832 38 -831
rect 51 -832 52 -831
rect 58 -832 59 -831
rect 180 -832 181 -831
rect 187 -832 188 -831
rect 310 -832 311 -831
rect 313 -832 314 -831
rect 548 -832 549 -831
rect 79 -834 80 -833
rect 163 -834 164 -833
rect 212 -834 213 -833
rect 219 -834 220 -833
rect 240 -834 241 -833
rect 275 -834 276 -833
rect 296 -834 297 -833
rect 450 -834 451 -833
rect 457 -834 458 -833
rect 464 -834 465 -833
rect 79 -836 80 -835
rect 170 -836 171 -835
rect 177 -836 178 -835
rect 219 -836 220 -835
rect 261 -836 262 -835
rect 324 -836 325 -835
rect 331 -836 332 -835
rect 366 -836 367 -835
rect 373 -836 374 -835
rect 513 -836 514 -835
rect 86 -838 87 -837
rect 201 -838 202 -837
rect 205 -838 206 -837
rect 261 -838 262 -837
rect 310 -838 311 -837
rect 317 -838 318 -837
rect 324 -838 325 -837
rect 359 -838 360 -837
rect 366 -838 367 -837
rect 429 -838 430 -837
rect 86 -840 87 -839
rect 135 -840 136 -839
rect 149 -840 150 -839
rect 558 -840 559 -839
rect 100 -842 101 -841
rect 226 -842 227 -841
rect 257 -842 258 -841
rect 513 -842 514 -841
rect 107 -844 108 -843
rect 191 -844 192 -843
rect 226 -844 227 -843
rect 282 -844 283 -843
rect 313 -844 314 -843
rect 471 -844 472 -843
rect 117 -846 118 -845
rect 429 -846 430 -845
rect 121 -848 122 -847
rect 303 -848 304 -847
rect 348 -848 349 -847
rect 499 -848 500 -847
rect 124 -850 125 -849
rect 128 -850 129 -849
rect 149 -850 150 -849
rect 334 -850 335 -849
rect 338 -850 339 -849
rect 499 -850 500 -849
rect 93 -852 94 -851
rect 128 -852 129 -851
rect 156 -852 157 -851
rect 275 -852 276 -851
rect 289 -852 290 -851
rect 338 -852 339 -851
rect 355 -852 356 -851
rect 534 -852 535 -851
rect 65 -854 66 -853
rect 93 -854 94 -853
rect 163 -854 164 -853
rect 184 -854 185 -853
rect 247 -854 248 -853
rect 355 -854 356 -853
rect 359 -854 360 -853
rect 408 -854 409 -853
rect 520 -854 521 -853
rect 534 -854 535 -853
rect 65 -856 66 -855
rect 198 -856 199 -855
rect 268 -856 269 -855
rect 289 -856 290 -855
rect 373 -856 374 -855
rect 506 -856 507 -855
rect 268 -858 269 -857
rect 380 -858 381 -857
rect 387 -858 388 -857
rect 474 -858 475 -857
rect 492 -858 493 -857
rect 506 -858 507 -857
rect 376 -860 377 -859
rect 527 -860 528 -859
rect 348 -862 349 -861
rect 527 -862 528 -861
rect 401 -864 402 -863
rect 436 -864 437 -863
rect 408 -866 409 -865
rect 422 -866 423 -865
rect 436 -866 437 -865
rect 478 -866 479 -865
rect 352 -868 353 -867
rect 478 -868 479 -867
rect 415 -870 416 -869
rect 492 -870 493 -869
rect 394 -872 395 -871
rect 415 -872 416 -871
rect 422 -872 423 -871
rect 443 -872 444 -871
rect 152 -874 153 -873
rect 443 -874 444 -873
rect 233 -876 234 -875
rect 394 -876 395 -875
rect 233 -878 234 -877
rect 296 -878 297 -877
rect 9 -889 10 -888
rect 135 -889 136 -888
rect 142 -889 143 -888
rect 156 -889 157 -888
rect 159 -889 160 -888
rect 492 -889 493 -888
rect 520 -889 521 -888
rect 534 -889 535 -888
rect 16 -891 17 -890
rect 208 -891 209 -890
rect 240 -891 241 -890
rect 264 -891 265 -890
rect 268 -891 269 -890
rect 334 -891 335 -890
rect 348 -891 349 -890
rect 485 -891 486 -890
rect 520 -891 521 -890
rect 523 -891 524 -890
rect 23 -893 24 -892
rect 44 -893 45 -892
rect 58 -893 59 -892
rect 345 -893 346 -892
rect 355 -893 356 -892
rect 436 -893 437 -892
rect 457 -893 458 -892
rect 492 -893 493 -892
rect 44 -895 45 -894
rect 51 -895 52 -894
rect 58 -895 59 -894
rect 72 -895 73 -894
rect 79 -895 80 -894
rect 170 -895 171 -894
rect 177 -895 178 -894
rect 212 -895 213 -894
rect 240 -895 241 -894
rect 334 -895 335 -894
rect 359 -895 360 -894
rect 362 -895 363 -894
rect 380 -895 381 -894
rect 513 -895 514 -894
rect 37 -897 38 -896
rect 212 -897 213 -896
rect 233 -897 234 -896
rect 380 -897 381 -896
rect 383 -897 384 -896
rect 513 -897 514 -896
rect 51 -899 52 -898
rect 285 -899 286 -898
rect 313 -899 314 -898
rect 408 -899 409 -898
rect 422 -899 423 -898
rect 474 -899 475 -898
rect 478 -899 479 -898
rect 485 -899 486 -898
rect 65 -901 66 -900
rect 138 -901 139 -900
rect 142 -901 143 -900
rect 254 -901 255 -900
rect 282 -901 283 -900
rect 324 -901 325 -900
rect 331 -901 332 -900
rect 499 -901 500 -900
rect 65 -903 66 -902
rect 191 -903 192 -902
rect 194 -903 195 -902
rect 261 -903 262 -902
rect 282 -903 283 -902
rect 324 -903 325 -902
rect 352 -903 353 -902
rect 499 -903 500 -902
rect 86 -905 87 -904
rect 229 -905 230 -904
rect 296 -905 297 -904
rect 422 -905 423 -904
rect 436 -905 437 -904
rect 443 -905 444 -904
rect 478 -905 479 -904
rect 506 -905 507 -904
rect 93 -907 94 -906
rect 163 -907 164 -906
rect 201 -907 202 -906
rect 292 -907 293 -906
rect 317 -907 318 -906
rect 345 -907 346 -906
rect 359 -907 360 -906
rect 401 -907 402 -906
rect 506 -907 507 -906
rect 527 -907 528 -906
rect 93 -909 94 -908
rect 128 -909 129 -908
rect 149 -909 150 -908
rect 268 -909 269 -908
rect 317 -909 318 -908
rect 338 -909 339 -908
rect 394 -909 395 -908
rect 408 -909 409 -908
rect 100 -911 101 -910
rect 180 -911 181 -910
rect 205 -911 206 -910
rect 289 -911 290 -910
rect 397 -911 398 -910
rect 471 -911 472 -910
rect 107 -913 108 -912
rect 306 -913 307 -912
rect 401 -913 402 -912
rect 415 -913 416 -912
rect 107 -915 108 -914
rect 247 -915 248 -914
rect 275 -915 276 -914
rect 338 -915 339 -914
rect 415 -915 416 -914
rect 429 -915 430 -914
rect 114 -917 115 -916
rect 149 -917 150 -916
rect 152 -917 153 -916
rect 170 -917 171 -916
rect 201 -917 202 -916
rect 247 -917 248 -916
rect 306 -917 307 -916
rect 366 -917 367 -916
rect 429 -917 430 -916
rect 450 -917 451 -916
rect 121 -919 122 -918
rect 184 -919 185 -918
rect 208 -919 209 -918
rect 296 -919 297 -918
rect 387 -919 388 -918
rect 450 -919 451 -918
rect 124 -921 125 -920
rect 166 -921 167 -920
rect 184 -921 185 -920
rect 222 -921 223 -920
rect 226 -921 227 -920
rect 233 -921 234 -920
rect 362 -921 363 -920
rect 387 -921 388 -920
rect 128 -923 129 -922
rect 194 -923 195 -922
rect 219 -923 220 -922
rect 275 -923 276 -922
rect 159 -925 160 -924
rect 310 -925 311 -924
rect 166 -927 167 -926
rect 254 -927 255 -926
rect 205 -929 206 -928
rect 310 -929 311 -928
rect 219 -931 220 -930
rect 366 -931 367 -930
rect 226 -933 227 -932
rect 457 -933 458 -932
rect 2 -944 3 -943
rect 163 -944 164 -943
rect 201 -944 202 -943
rect 422 -944 423 -943
rect 443 -944 444 -943
rect 499 -944 500 -943
rect 16 -946 17 -945
rect 103 -946 104 -945
rect 107 -946 108 -945
rect 110 -946 111 -945
rect 114 -946 115 -945
rect 138 -946 139 -945
rect 142 -946 143 -945
rect 191 -946 192 -945
rect 212 -946 213 -945
rect 240 -946 241 -945
rect 257 -946 258 -945
rect 296 -946 297 -945
rect 299 -946 300 -945
rect 415 -946 416 -945
rect 429 -946 430 -945
rect 443 -946 444 -945
rect 464 -946 465 -945
rect 485 -946 486 -945
rect 9 -948 10 -947
rect 191 -948 192 -947
rect 222 -948 223 -947
rect 261 -948 262 -947
rect 268 -948 269 -947
rect 303 -948 304 -947
rect 310 -948 311 -947
rect 408 -948 409 -947
rect 467 -948 468 -947
rect 492 -948 493 -947
rect 23 -950 24 -949
rect 30 -950 31 -949
rect 37 -950 38 -949
rect 198 -950 199 -949
rect 254 -950 255 -949
rect 310 -950 311 -949
rect 324 -950 325 -949
rect 401 -950 402 -949
rect 492 -950 493 -949
rect 513 -950 514 -949
rect 9 -952 10 -951
rect 30 -952 31 -951
rect 44 -952 45 -951
rect 184 -952 185 -951
rect 187 -952 188 -951
rect 212 -952 213 -951
rect 268 -952 269 -951
rect 275 -952 276 -951
rect 296 -952 297 -951
rect 324 -952 325 -951
rect 327 -952 328 -951
rect 415 -952 416 -951
rect 16 -954 17 -953
rect 23 -954 24 -953
rect 51 -954 52 -953
rect 166 -954 167 -953
rect 198 -954 199 -953
rect 429 -954 430 -953
rect 51 -956 52 -955
rect 58 -956 59 -955
rect 65 -956 66 -955
rect 201 -956 202 -955
rect 247 -956 248 -955
rect 275 -956 276 -955
rect 338 -956 339 -955
rect 380 -956 381 -955
rect 394 -956 395 -955
rect 478 -956 479 -955
rect 65 -958 66 -957
rect 205 -958 206 -957
rect 306 -958 307 -957
rect 394 -958 395 -957
rect 478 -958 479 -957
rect 506 -958 507 -957
rect 75 -960 76 -959
rect 100 -960 101 -959
rect 107 -960 108 -959
rect 170 -960 171 -959
rect 177 -960 178 -959
rect 205 -960 206 -959
rect 331 -960 332 -959
rect 338 -960 339 -959
rect 345 -960 346 -959
rect 401 -960 402 -959
rect 506 -960 507 -959
rect 520 -960 521 -959
rect 86 -962 87 -961
rect 156 -962 157 -961
rect 163 -962 164 -961
rect 282 -962 283 -961
rect 289 -962 290 -961
rect 345 -962 346 -961
rect 352 -962 353 -961
rect 450 -962 451 -961
rect 86 -964 87 -963
rect 292 -964 293 -963
rect 373 -964 374 -963
rect 422 -964 423 -963
rect 93 -966 94 -965
rect 103 -966 104 -965
rect 110 -966 111 -965
rect 170 -966 171 -965
rect 177 -966 178 -965
rect 264 -966 265 -965
rect 373 -966 374 -965
rect 387 -966 388 -965
rect 96 -968 97 -967
rect 471 -968 472 -967
rect 114 -970 115 -969
rect 166 -970 167 -969
rect 194 -970 195 -969
rect 247 -970 248 -969
rect 264 -970 265 -969
rect 436 -970 437 -969
rect 457 -970 458 -969
rect 471 -970 472 -969
rect 121 -972 122 -971
rect 219 -972 220 -971
rect 226 -972 227 -971
rect 457 -972 458 -971
rect 128 -974 129 -973
rect 184 -974 185 -973
rect 233 -974 234 -973
rect 282 -974 283 -973
rect 359 -974 360 -973
rect 387 -974 388 -973
rect 82 -976 83 -975
rect 233 -976 234 -975
rect 355 -976 356 -975
rect 359 -976 360 -975
rect 366 -976 367 -975
rect 436 -976 437 -975
rect 135 -978 136 -977
rect 142 -978 143 -977
rect 149 -978 150 -977
rect 229 -978 230 -977
rect 334 -978 335 -977
rect 366 -978 367 -977
rect 159 -980 160 -979
rect 219 -980 220 -979
rect 334 -980 335 -979
rect 450 -980 451 -979
rect 121 -982 122 -981
rect 159 -982 160 -981
rect 9 -993 10 -992
rect 37 -993 38 -992
rect 44 -993 45 -992
rect 219 -993 220 -992
rect 229 -993 230 -992
rect 240 -993 241 -992
rect 278 -993 279 -992
rect 380 -993 381 -992
rect 418 -993 419 -992
rect 436 -993 437 -992
rect 439 -993 440 -992
rect 478 -993 479 -992
rect 488 -993 489 -992
rect 506 -993 507 -992
rect 23 -995 24 -994
rect 33 -995 34 -994
rect 37 -995 38 -994
rect 47 -995 48 -994
rect 51 -995 52 -994
rect 58 -995 59 -994
rect 65 -995 66 -994
rect 93 -995 94 -994
rect 107 -995 108 -994
rect 184 -995 185 -994
rect 187 -995 188 -994
rect 275 -995 276 -994
rect 289 -995 290 -994
rect 317 -995 318 -994
rect 341 -995 342 -994
rect 443 -995 444 -994
rect 446 -995 447 -994
rect 478 -995 479 -994
rect 40 -997 41 -996
rect 93 -997 94 -996
rect 107 -997 108 -996
rect 194 -997 195 -996
rect 215 -997 216 -996
rect 229 -997 230 -996
rect 233 -997 234 -996
rect 345 -997 346 -996
rect 352 -997 353 -996
rect 450 -997 451 -996
rect 467 -997 468 -996
rect 471 -997 472 -996
rect 474 -997 475 -996
rect 492 -997 493 -996
rect 58 -999 59 -998
rect 61 -999 62 -998
rect 79 -999 80 -998
rect 114 -999 115 -998
rect 131 -999 132 -998
rect 324 -999 325 -998
rect 327 -999 328 -998
rect 345 -999 346 -998
rect 380 -999 381 -998
rect 387 -999 388 -998
rect 415 -999 416 -998
rect 450 -999 451 -998
rect 82 -1001 83 -1000
rect 457 -1001 458 -1000
rect 2 -1003 3 -1002
rect 82 -1003 83 -1002
rect 86 -1003 87 -1002
rect 243 -1003 244 -1002
rect 285 -1003 286 -1002
rect 289 -1003 290 -1002
rect 303 -1003 304 -1002
rect 317 -1003 318 -1002
rect 334 -1003 335 -1002
rect 352 -1003 353 -1002
rect 366 -1003 367 -1002
rect 387 -1003 388 -1002
rect 422 -1003 423 -1002
rect 464 -1003 465 -1002
rect 86 -1005 87 -1004
rect 103 -1005 104 -1004
rect 149 -1005 150 -1004
rect 159 -1005 160 -1004
rect 163 -1005 164 -1004
rect 166 -1005 167 -1004
rect 170 -1005 171 -1004
rect 226 -1005 227 -1004
rect 310 -1005 311 -1004
rect 366 -1005 367 -1004
rect 96 -1007 97 -1006
rect 114 -1007 115 -1006
rect 149 -1007 150 -1006
rect 429 -1007 430 -1006
rect 156 -1009 157 -1008
rect 170 -1009 171 -1008
rect 191 -1009 192 -1008
rect 282 -1009 283 -1008
rect 415 -1009 416 -1008
rect 429 -1009 430 -1008
rect 191 -1011 192 -1010
rect 212 -1011 213 -1010
rect 222 -1011 223 -1010
rect 310 -1011 311 -1010
rect 212 -1013 213 -1012
rect 268 -1013 269 -1012
rect 128 -1015 129 -1014
rect 268 -1015 269 -1014
rect 128 -1017 129 -1016
rect 177 -1017 178 -1016
rect 222 -1017 223 -1016
rect 408 -1017 409 -1016
rect 177 -1019 178 -1018
rect 198 -1019 199 -1018
rect 394 -1019 395 -1018
rect 408 -1019 409 -1018
rect 198 -1021 199 -1020
rect 261 -1021 262 -1020
rect 373 -1021 374 -1020
rect 394 -1021 395 -1020
rect 254 -1023 255 -1022
rect 261 -1023 262 -1022
rect 373 -1023 374 -1022
rect 460 -1023 461 -1022
rect 254 -1025 255 -1024
rect 338 -1025 339 -1024
rect 338 -1027 339 -1026
rect 401 -1027 402 -1026
rect 292 -1029 293 -1028
rect 401 -1029 402 -1028
rect 23 -1040 24 -1039
rect 33 -1040 34 -1039
rect 51 -1040 52 -1039
rect 58 -1040 59 -1039
rect 72 -1040 73 -1039
rect 79 -1040 80 -1039
rect 86 -1040 87 -1039
rect 100 -1040 101 -1039
rect 117 -1040 118 -1039
rect 121 -1040 122 -1039
rect 128 -1040 129 -1039
rect 156 -1040 157 -1039
rect 159 -1040 160 -1039
rect 296 -1040 297 -1039
rect 299 -1040 300 -1039
rect 359 -1040 360 -1039
rect 408 -1040 409 -1039
rect 422 -1040 423 -1039
rect 443 -1040 444 -1039
rect 450 -1040 451 -1039
rect 460 -1040 461 -1039
rect 467 -1040 468 -1039
rect 488 -1040 489 -1039
rect 499 -1040 500 -1039
rect 30 -1042 31 -1041
rect 37 -1042 38 -1041
rect 68 -1042 69 -1041
rect 79 -1042 80 -1041
rect 100 -1042 101 -1041
rect 114 -1042 115 -1041
rect 121 -1042 122 -1041
rect 138 -1042 139 -1041
rect 149 -1042 150 -1041
rect 170 -1042 171 -1041
rect 177 -1042 178 -1041
rect 184 -1042 185 -1041
rect 205 -1042 206 -1041
rect 226 -1042 227 -1041
rect 233 -1042 234 -1041
rect 275 -1042 276 -1041
rect 285 -1042 286 -1041
rect 317 -1042 318 -1041
rect 324 -1042 325 -1041
rect 387 -1042 388 -1041
rect 401 -1042 402 -1041
rect 422 -1042 423 -1041
rect 429 -1042 430 -1041
rect 450 -1042 451 -1041
rect 464 -1042 465 -1041
rect 471 -1042 472 -1041
rect 37 -1044 38 -1043
rect 96 -1044 97 -1043
rect 110 -1044 111 -1043
rect 156 -1044 157 -1043
rect 163 -1044 164 -1043
rect 254 -1044 255 -1043
rect 261 -1044 262 -1043
rect 306 -1044 307 -1043
rect 331 -1044 332 -1043
rect 338 -1044 339 -1043
rect 345 -1044 346 -1043
rect 359 -1044 360 -1043
rect 394 -1044 395 -1043
rect 401 -1044 402 -1043
rect 408 -1044 409 -1043
rect 495 -1044 496 -1043
rect 86 -1046 87 -1045
rect 114 -1046 115 -1045
rect 128 -1046 129 -1045
rect 485 -1046 486 -1045
rect 135 -1048 136 -1047
rect 142 -1048 143 -1047
rect 177 -1048 178 -1047
rect 219 -1048 220 -1047
rect 222 -1048 223 -1047
rect 278 -1048 279 -1047
rect 303 -1048 304 -1047
rect 366 -1048 367 -1047
rect 418 -1048 419 -1047
rect 457 -1048 458 -1047
rect 478 -1048 479 -1047
rect 485 -1048 486 -1047
rect 107 -1050 108 -1049
rect 142 -1050 143 -1049
rect 184 -1050 185 -1049
rect 191 -1050 192 -1049
rect 198 -1050 199 -1049
rect 205 -1050 206 -1049
rect 215 -1050 216 -1049
rect 387 -1050 388 -1049
rect 96 -1052 97 -1051
rect 191 -1052 192 -1051
rect 198 -1052 199 -1051
rect 415 -1052 416 -1051
rect 135 -1054 136 -1053
rect 173 -1054 174 -1053
rect 233 -1054 234 -1053
rect 261 -1054 262 -1053
rect 268 -1054 269 -1053
rect 324 -1054 325 -1053
rect 338 -1054 339 -1053
rect 429 -1054 430 -1053
rect 240 -1056 241 -1055
rect 282 -1056 283 -1055
rect 303 -1056 304 -1055
rect 443 -1056 444 -1055
rect 240 -1058 241 -1057
rect 327 -1058 328 -1057
rect 341 -1058 342 -1057
rect 457 -1058 458 -1057
rect 247 -1060 248 -1059
rect 254 -1060 255 -1059
rect 268 -1060 269 -1059
rect 366 -1060 367 -1059
rect 149 -1062 150 -1061
rect 247 -1062 248 -1061
rect 278 -1062 279 -1061
rect 317 -1062 318 -1061
rect 348 -1062 349 -1061
rect 380 -1062 381 -1061
rect 310 -1064 311 -1063
rect 394 -1064 395 -1063
rect 289 -1066 290 -1065
rect 310 -1066 311 -1065
rect 373 -1066 374 -1065
rect 380 -1066 381 -1065
rect 229 -1068 230 -1067
rect 373 -1068 374 -1067
rect 289 -1070 290 -1069
rect 352 -1070 353 -1069
rect 352 -1072 353 -1071
rect 436 -1072 437 -1071
rect 345 -1074 346 -1073
rect 436 -1074 437 -1073
rect 30 -1085 31 -1084
rect 44 -1085 45 -1084
rect 47 -1085 48 -1084
rect 61 -1085 62 -1084
rect 86 -1085 87 -1084
rect 89 -1085 90 -1084
rect 96 -1085 97 -1084
rect 177 -1085 178 -1084
rect 191 -1085 192 -1084
rect 208 -1085 209 -1084
rect 212 -1085 213 -1084
rect 324 -1085 325 -1084
rect 338 -1085 339 -1084
rect 401 -1085 402 -1084
rect 432 -1085 433 -1084
rect 464 -1085 465 -1084
rect 471 -1085 472 -1084
rect 478 -1085 479 -1084
rect 481 -1085 482 -1084
rect 485 -1085 486 -1084
rect 495 -1085 496 -1084
rect 499 -1085 500 -1084
rect 37 -1087 38 -1086
rect 201 -1087 202 -1086
rect 212 -1087 213 -1086
rect 341 -1087 342 -1086
rect 345 -1087 346 -1086
rect 387 -1087 388 -1086
rect 401 -1087 402 -1086
rect 457 -1087 458 -1086
rect 51 -1089 52 -1088
rect 65 -1089 66 -1088
rect 100 -1089 101 -1088
rect 159 -1089 160 -1088
rect 170 -1089 171 -1088
rect 247 -1089 248 -1088
rect 271 -1089 272 -1088
rect 310 -1089 311 -1088
rect 338 -1089 339 -1088
rect 373 -1089 374 -1088
rect 450 -1089 451 -1088
rect 457 -1089 458 -1088
rect 58 -1091 59 -1090
rect 110 -1091 111 -1090
rect 114 -1091 115 -1090
rect 135 -1091 136 -1090
rect 149 -1091 150 -1090
rect 240 -1091 241 -1090
rect 271 -1091 272 -1090
rect 331 -1091 332 -1090
rect 348 -1091 349 -1090
rect 380 -1091 381 -1090
rect 65 -1093 66 -1092
rect 72 -1093 73 -1092
rect 100 -1093 101 -1092
rect 121 -1093 122 -1092
rect 124 -1093 125 -1092
rect 135 -1093 136 -1092
rect 149 -1093 150 -1092
rect 226 -1093 227 -1092
rect 229 -1093 230 -1092
rect 317 -1093 318 -1092
rect 352 -1093 353 -1092
rect 387 -1093 388 -1092
rect 72 -1095 73 -1094
rect 86 -1095 87 -1094
rect 163 -1095 164 -1094
rect 170 -1095 171 -1094
rect 173 -1095 174 -1094
rect 236 -1095 237 -1094
rect 240 -1095 241 -1094
rect 247 -1095 248 -1094
rect 268 -1095 269 -1094
rect 317 -1095 318 -1094
rect 366 -1095 367 -1094
rect 376 -1095 377 -1094
rect 380 -1095 381 -1094
rect 415 -1095 416 -1094
rect 82 -1097 83 -1096
rect 121 -1097 122 -1096
rect 156 -1097 157 -1096
rect 163 -1097 164 -1096
rect 177 -1097 178 -1096
rect 222 -1097 223 -1096
rect 226 -1097 227 -1096
rect 331 -1097 332 -1096
rect 366 -1097 367 -1096
rect 443 -1097 444 -1096
rect 156 -1099 157 -1098
rect 278 -1099 279 -1098
rect 289 -1099 290 -1098
rect 359 -1099 360 -1098
rect 369 -1099 370 -1098
rect 429 -1099 430 -1098
rect 194 -1101 195 -1100
rect 215 -1101 216 -1100
rect 236 -1101 237 -1100
rect 254 -1101 255 -1100
rect 275 -1101 276 -1100
rect 296 -1101 297 -1100
rect 310 -1101 311 -1100
rect 324 -1101 325 -1100
rect 359 -1101 360 -1100
rect 394 -1101 395 -1100
rect 422 -1101 423 -1100
rect 443 -1101 444 -1100
rect 107 -1103 108 -1102
rect 215 -1103 216 -1102
rect 233 -1103 234 -1102
rect 254 -1103 255 -1102
rect 261 -1103 262 -1102
rect 296 -1103 297 -1102
rect 373 -1103 374 -1102
rect 408 -1103 409 -1102
rect 145 -1105 146 -1104
rect 261 -1105 262 -1104
rect 376 -1105 377 -1104
rect 422 -1105 423 -1104
rect 205 -1107 206 -1106
rect 222 -1107 223 -1106
rect 394 -1107 395 -1106
rect 415 -1107 416 -1106
rect 47 -1118 48 -1117
rect 51 -1118 52 -1117
rect 72 -1118 73 -1117
rect 82 -1118 83 -1117
rect 100 -1118 101 -1117
rect 124 -1118 125 -1117
rect 149 -1118 150 -1117
rect 208 -1118 209 -1117
rect 212 -1118 213 -1117
rect 222 -1118 223 -1117
rect 229 -1118 230 -1117
rect 313 -1118 314 -1117
rect 334 -1118 335 -1117
rect 387 -1118 388 -1117
rect 394 -1118 395 -1117
rect 401 -1118 402 -1117
rect 408 -1118 409 -1117
rect 443 -1118 444 -1117
rect 65 -1120 66 -1119
rect 72 -1120 73 -1119
rect 100 -1120 101 -1119
rect 268 -1120 269 -1119
rect 285 -1120 286 -1119
rect 296 -1120 297 -1119
rect 306 -1120 307 -1119
rect 331 -1120 332 -1119
rect 338 -1120 339 -1119
rect 397 -1120 398 -1119
rect 408 -1120 409 -1119
rect 415 -1120 416 -1119
rect 422 -1120 423 -1119
rect 450 -1120 451 -1119
rect 65 -1122 66 -1121
rect 75 -1122 76 -1121
rect 110 -1122 111 -1121
rect 121 -1122 122 -1121
rect 149 -1122 150 -1121
rect 226 -1122 227 -1121
rect 233 -1122 234 -1121
rect 257 -1122 258 -1121
rect 275 -1122 276 -1121
rect 296 -1122 297 -1121
rect 317 -1122 318 -1121
rect 338 -1122 339 -1121
rect 352 -1122 353 -1121
rect 359 -1122 360 -1121
rect 366 -1122 367 -1121
rect 401 -1122 402 -1121
rect 415 -1122 416 -1121
rect 432 -1122 433 -1121
rect 450 -1122 451 -1121
rect 457 -1122 458 -1121
rect 114 -1124 115 -1123
rect 142 -1124 143 -1123
rect 170 -1124 171 -1123
rect 282 -1124 283 -1123
rect 289 -1124 290 -1123
rect 310 -1124 311 -1123
rect 317 -1124 318 -1123
rect 380 -1124 381 -1123
rect 387 -1124 388 -1123
rect 404 -1124 405 -1123
rect 422 -1124 423 -1123
rect 436 -1124 437 -1123
rect 114 -1126 115 -1125
rect 128 -1126 129 -1125
rect 135 -1126 136 -1125
rect 142 -1126 143 -1125
rect 170 -1126 171 -1125
rect 229 -1126 230 -1125
rect 240 -1126 241 -1125
rect 271 -1126 272 -1125
rect 310 -1126 311 -1125
rect 345 -1126 346 -1125
rect 177 -1128 178 -1127
rect 201 -1128 202 -1127
rect 205 -1128 206 -1127
rect 233 -1128 234 -1127
rect 243 -1128 244 -1127
rect 352 -1128 353 -1127
rect 184 -1130 185 -1129
rect 191 -1130 192 -1129
rect 198 -1130 199 -1129
rect 240 -1130 241 -1129
rect 247 -1130 248 -1129
rect 303 -1130 304 -1129
rect 331 -1130 332 -1129
rect 373 -1130 374 -1129
rect 163 -1132 164 -1131
rect 191 -1132 192 -1131
rect 226 -1132 227 -1131
rect 383 -1132 384 -1131
rect 254 -1134 255 -1133
rect 275 -1134 276 -1133
rect 303 -1134 304 -1133
rect 359 -1134 360 -1133
rect 156 -1136 157 -1135
rect 254 -1136 255 -1135
rect 268 -1136 269 -1135
rect 289 -1136 290 -1135
rect 324 -1136 325 -1135
rect 373 -1136 374 -1135
rect 156 -1138 157 -1137
rect 194 -1138 195 -1137
rect 250 -1138 251 -1137
rect 324 -1138 325 -1137
rect 345 -1138 346 -1137
rect 369 -1138 370 -1137
rect 177 -1140 178 -1139
rect 194 -1140 195 -1139
rect 47 -1151 48 -1150
rect 51 -1151 52 -1150
rect 58 -1151 59 -1150
rect 82 -1151 83 -1150
rect 89 -1151 90 -1150
rect 107 -1151 108 -1150
rect 114 -1151 115 -1150
rect 184 -1151 185 -1150
rect 191 -1151 192 -1150
rect 205 -1151 206 -1150
rect 212 -1151 213 -1150
rect 296 -1151 297 -1150
rect 299 -1151 300 -1150
rect 387 -1151 388 -1150
rect 394 -1151 395 -1150
rect 404 -1151 405 -1150
rect 408 -1151 409 -1150
rect 418 -1151 419 -1150
rect 446 -1151 447 -1150
rect 450 -1151 451 -1150
rect 51 -1153 52 -1152
rect 61 -1153 62 -1152
rect 65 -1153 66 -1152
rect 86 -1153 87 -1152
rect 107 -1153 108 -1152
rect 128 -1153 129 -1152
rect 135 -1153 136 -1152
rect 149 -1153 150 -1152
rect 170 -1153 171 -1152
rect 184 -1153 185 -1152
rect 194 -1153 195 -1152
rect 282 -1153 283 -1152
rect 303 -1153 304 -1152
rect 373 -1153 374 -1152
rect 65 -1155 66 -1154
rect 187 -1155 188 -1154
rect 212 -1155 213 -1154
rect 236 -1155 237 -1154
rect 240 -1155 241 -1154
rect 338 -1155 339 -1154
rect 100 -1157 101 -1156
rect 135 -1157 136 -1156
rect 142 -1157 143 -1156
rect 145 -1157 146 -1156
rect 177 -1157 178 -1156
rect 208 -1157 209 -1156
rect 222 -1157 223 -1156
rect 233 -1157 234 -1156
rect 243 -1157 244 -1156
rect 261 -1157 262 -1156
rect 271 -1157 272 -1156
rect 317 -1157 318 -1156
rect 324 -1157 325 -1156
rect 327 -1157 328 -1156
rect 338 -1157 339 -1156
rect 366 -1157 367 -1156
rect 100 -1159 101 -1158
rect 215 -1159 216 -1158
rect 226 -1159 227 -1158
rect 345 -1159 346 -1158
rect 359 -1159 360 -1158
rect 366 -1159 367 -1158
rect 117 -1161 118 -1160
rect 121 -1161 122 -1160
rect 128 -1161 129 -1160
rect 243 -1161 244 -1160
rect 247 -1161 248 -1160
rect 359 -1161 360 -1160
rect 121 -1163 122 -1162
rect 156 -1163 157 -1162
rect 226 -1163 227 -1162
rect 282 -1163 283 -1162
rect 306 -1163 307 -1162
rect 373 -1163 374 -1162
rect 156 -1165 157 -1164
rect 163 -1165 164 -1164
rect 229 -1165 230 -1164
rect 268 -1165 269 -1164
rect 310 -1165 311 -1164
rect 380 -1165 381 -1164
rect 198 -1167 199 -1166
rect 268 -1167 269 -1166
rect 296 -1167 297 -1166
rect 310 -1167 311 -1166
rect 313 -1167 314 -1166
rect 415 -1167 416 -1166
rect 233 -1169 234 -1168
rect 289 -1169 290 -1168
rect 317 -1169 318 -1168
rect 401 -1169 402 -1168
rect 415 -1169 416 -1168
rect 429 -1169 430 -1168
rect 254 -1171 255 -1170
rect 261 -1171 262 -1170
rect 324 -1171 325 -1170
rect 331 -1171 332 -1170
rect 352 -1171 353 -1170
rect 401 -1171 402 -1170
rect 247 -1173 248 -1172
rect 352 -1173 353 -1172
rect 257 -1175 258 -1174
rect 394 -1175 395 -1174
rect 327 -1177 328 -1176
rect 331 -1177 332 -1176
rect 51 -1188 52 -1187
rect 68 -1188 69 -1187
rect 72 -1188 73 -1187
rect 75 -1188 76 -1187
rect 89 -1188 90 -1187
rect 96 -1188 97 -1187
rect 100 -1188 101 -1187
rect 142 -1188 143 -1187
rect 156 -1188 157 -1187
rect 222 -1188 223 -1187
rect 229 -1188 230 -1187
rect 275 -1188 276 -1187
rect 289 -1188 290 -1187
rect 324 -1188 325 -1187
rect 338 -1188 339 -1187
rect 348 -1188 349 -1187
rect 408 -1188 409 -1187
rect 415 -1188 416 -1187
rect 422 -1188 423 -1187
rect 425 -1188 426 -1187
rect 65 -1190 66 -1189
rect 82 -1190 83 -1189
rect 93 -1190 94 -1189
rect 100 -1190 101 -1189
rect 107 -1190 108 -1189
rect 149 -1190 150 -1189
rect 166 -1190 167 -1189
rect 198 -1190 199 -1189
rect 219 -1190 220 -1189
rect 310 -1190 311 -1189
rect 324 -1190 325 -1189
rect 352 -1190 353 -1189
rect 422 -1190 423 -1189
rect 429 -1190 430 -1189
rect 79 -1192 80 -1191
rect 166 -1192 167 -1191
rect 170 -1192 171 -1191
rect 177 -1192 178 -1191
rect 184 -1192 185 -1191
rect 201 -1192 202 -1191
rect 229 -1192 230 -1191
rect 254 -1192 255 -1191
rect 268 -1192 269 -1191
rect 292 -1192 293 -1191
rect 303 -1192 304 -1191
rect 331 -1192 332 -1191
rect 345 -1192 346 -1191
rect 387 -1192 388 -1191
rect 425 -1192 426 -1191
rect 429 -1192 430 -1191
rect 79 -1194 80 -1193
rect 114 -1194 115 -1193
rect 121 -1194 122 -1193
rect 152 -1194 153 -1193
rect 159 -1194 160 -1193
rect 177 -1194 178 -1193
rect 240 -1194 241 -1193
rect 317 -1194 318 -1193
rect 331 -1194 332 -1193
rect 341 -1194 342 -1193
rect 345 -1194 346 -1193
rect 401 -1194 402 -1193
rect 107 -1196 108 -1195
rect 145 -1196 146 -1195
rect 149 -1196 150 -1195
rect 191 -1196 192 -1195
rect 233 -1196 234 -1195
rect 240 -1196 241 -1195
rect 247 -1196 248 -1195
rect 261 -1196 262 -1195
rect 282 -1196 283 -1195
rect 303 -1196 304 -1195
rect 317 -1196 318 -1195
rect 373 -1196 374 -1195
rect 128 -1198 129 -1197
rect 226 -1198 227 -1197
rect 236 -1198 237 -1197
rect 282 -1198 283 -1197
rect 289 -1198 290 -1197
rect 359 -1198 360 -1197
rect 128 -1200 129 -1199
rect 156 -1200 157 -1199
rect 184 -1200 185 -1199
rect 226 -1200 227 -1199
rect 292 -1200 293 -1199
rect 296 -1200 297 -1199
rect 359 -1200 360 -1199
rect 366 -1200 367 -1199
rect 135 -1202 136 -1201
rect 173 -1202 174 -1201
rect 366 -1202 367 -1201
rect 394 -1202 395 -1201
rect 121 -1204 122 -1203
rect 135 -1204 136 -1203
rect 138 -1204 139 -1203
rect 222 -1204 223 -1203
rect 33 -1215 34 -1214
rect 37 -1215 38 -1214
rect 44 -1215 45 -1214
rect 51 -1215 52 -1214
rect 58 -1215 59 -1214
rect 65 -1215 66 -1214
rect 72 -1215 73 -1214
rect 79 -1215 80 -1214
rect 89 -1215 90 -1214
rect 100 -1215 101 -1214
rect 107 -1215 108 -1214
rect 173 -1215 174 -1214
rect 180 -1215 181 -1214
rect 205 -1215 206 -1214
rect 229 -1215 230 -1214
rect 247 -1215 248 -1214
rect 254 -1215 255 -1214
rect 268 -1215 269 -1214
rect 303 -1215 304 -1214
rect 341 -1215 342 -1214
rect 373 -1215 374 -1214
rect 380 -1215 381 -1214
rect 401 -1215 402 -1214
rect 408 -1215 409 -1214
rect 422 -1215 423 -1214
rect 429 -1215 430 -1214
rect 72 -1217 73 -1216
rect 79 -1217 80 -1216
rect 93 -1217 94 -1216
rect 138 -1217 139 -1216
rect 152 -1217 153 -1216
rect 159 -1217 160 -1216
rect 163 -1217 164 -1216
rect 212 -1217 213 -1216
rect 229 -1217 230 -1216
rect 240 -1217 241 -1216
rect 243 -1217 244 -1216
rect 292 -1217 293 -1216
rect 296 -1217 297 -1216
rect 303 -1217 304 -1216
rect 306 -1217 307 -1216
rect 324 -1217 325 -1216
rect 331 -1217 332 -1216
rect 352 -1217 353 -1216
rect 425 -1217 426 -1216
rect 432 -1217 433 -1216
rect 114 -1219 115 -1218
rect 121 -1219 122 -1218
rect 128 -1219 129 -1218
rect 142 -1219 143 -1218
rect 163 -1219 164 -1218
rect 177 -1219 178 -1218
rect 184 -1219 185 -1218
rect 201 -1219 202 -1218
rect 212 -1219 213 -1218
rect 254 -1219 255 -1218
rect 275 -1219 276 -1218
rect 292 -1219 293 -1218
rect 310 -1219 311 -1218
rect 345 -1219 346 -1218
rect 352 -1219 353 -1218
rect 366 -1219 367 -1218
rect 100 -1221 101 -1220
rect 128 -1221 129 -1220
rect 135 -1221 136 -1220
rect 156 -1221 157 -1220
rect 170 -1221 171 -1220
rect 187 -1221 188 -1220
rect 191 -1221 192 -1220
rect 222 -1221 223 -1220
rect 282 -1221 283 -1220
rect 310 -1221 311 -1220
rect 317 -1221 318 -1220
rect 320 -1221 321 -1220
rect 338 -1221 339 -1220
rect 345 -1221 346 -1220
rect 366 -1221 367 -1220
rect 373 -1221 374 -1220
rect 121 -1223 122 -1222
rect 149 -1223 150 -1222
rect 194 -1223 195 -1222
rect 198 -1223 199 -1222
rect 215 -1223 216 -1222
rect 317 -1223 318 -1222
rect 124 -1225 125 -1224
rect 142 -1225 143 -1224
rect 222 -1225 223 -1224
rect 233 -1225 234 -1224
rect 282 -1225 283 -1224
rect 313 -1225 314 -1224
rect 219 -1227 220 -1226
rect 233 -1227 234 -1226
rect 30 -1238 31 -1237
rect 37 -1238 38 -1237
rect 44 -1238 45 -1237
rect 51 -1238 52 -1237
rect 65 -1238 66 -1237
rect 75 -1238 76 -1237
rect 93 -1238 94 -1237
rect 117 -1238 118 -1237
rect 128 -1238 129 -1237
rect 149 -1238 150 -1237
rect 152 -1238 153 -1237
rect 208 -1238 209 -1237
rect 222 -1238 223 -1237
rect 268 -1238 269 -1237
rect 275 -1238 276 -1237
rect 289 -1238 290 -1237
rect 299 -1238 300 -1237
rect 310 -1238 311 -1237
rect 324 -1238 325 -1237
rect 327 -1238 328 -1237
rect 334 -1238 335 -1237
rect 338 -1238 339 -1237
rect 369 -1238 370 -1237
rect 373 -1238 374 -1237
rect 401 -1238 402 -1237
rect 408 -1238 409 -1237
rect 415 -1238 416 -1237
rect 422 -1238 423 -1237
rect 100 -1240 101 -1239
rect 114 -1240 115 -1239
rect 128 -1240 129 -1239
rect 138 -1240 139 -1239
rect 142 -1240 143 -1239
rect 145 -1240 146 -1239
rect 163 -1240 164 -1239
rect 215 -1240 216 -1239
rect 226 -1240 227 -1239
rect 278 -1240 279 -1239
rect 338 -1240 339 -1239
rect 352 -1240 353 -1239
rect 103 -1242 104 -1241
rect 121 -1242 122 -1241
rect 177 -1242 178 -1241
rect 191 -1242 192 -1241
rect 194 -1242 195 -1241
rect 240 -1242 241 -1241
rect 250 -1242 251 -1241
rect 268 -1242 269 -1241
rect 110 -1244 111 -1243
rect 114 -1244 115 -1243
rect 205 -1244 206 -1243
rect 282 -1244 283 -1243
rect 208 -1246 209 -1245
rect 254 -1246 255 -1245
rect 212 -1248 213 -1247
rect 222 -1248 223 -1247
rect 233 -1248 234 -1247
rect 257 -1248 258 -1247
rect 170 -1250 171 -1249
rect 233 -1250 234 -1249
rect 170 -1252 171 -1251
rect 184 -1252 185 -1251
rect 219 -1252 220 -1251
rect 240 -1252 241 -1251
rect 30 -1263 31 -1262
rect 37 -1263 38 -1262
rect 58 -1263 59 -1262
rect 68 -1263 69 -1262
rect 72 -1263 73 -1262
rect 79 -1263 80 -1262
rect 107 -1263 108 -1262
rect 114 -1263 115 -1262
rect 121 -1263 122 -1262
rect 152 -1263 153 -1262
rect 170 -1263 171 -1262
rect 205 -1263 206 -1262
rect 208 -1263 209 -1262
rect 212 -1263 213 -1262
rect 226 -1263 227 -1262
rect 268 -1263 269 -1262
rect 285 -1263 286 -1262
rect 289 -1263 290 -1262
rect 296 -1263 297 -1262
rect 303 -1263 304 -1262
rect 317 -1263 318 -1262
rect 324 -1263 325 -1262
rect 338 -1263 339 -1262
rect 348 -1263 349 -1262
rect 355 -1263 356 -1262
rect 359 -1263 360 -1262
rect 128 -1265 129 -1264
rect 138 -1265 139 -1264
rect 142 -1265 143 -1264
rect 163 -1265 164 -1264
rect 177 -1265 178 -1264
rect 187 -1265 188 -1264
rect 198 -1265 199 -1264
rect 233 -1265 234 -1264
rect 250 -1265 251 -1264
rect 261 -1265 262 -1264
<< metal2 >>
rect 138 -3 139 1
rect 149 -3 150 1
rect 177 -3 178 1
rect 191 -3 192 1
rect 198 -3 199 1
rect 215 -3 216 1
rect 226 -3 227 1
rect 240 -3 241 1
rect 187 -3 188 -1
rect 205 -3 206 -1
rect 212 -3 213 -1
rect 219 -3 220 -1
rect 135 -22 136 -12
rect 184 -13 185 -11
rect 187 -13 188 -11
rect 229 -13 230 -11
rect 240 -13 241 -11
rect 247 -22 248 -12
rect 324 -22 325 -12
rect 331 -22 332 -12
rect 142 -15 143 -11
rect 142 -22 143 -14
rect 142 -15 143 -11
rect 142 -22 143 -14
rect 145 -15 146 -11
rect 149 -15 150 -11
rect 163 -22 164 -14
rect 170 -22 171 -14
rect 177 -15 178 -11
rect 184 -22 185 -14
rect 191 -22 192 -14
rect 233 -22 234 -14
rect 156 -22 157 -16
rect 177 -22 178 -16
rect 198 -17 199 -11
rect 205 -22 206 -16
rect 208 -17 209 -11
rect 219 -17 220 -11
rect 226 -22 227 -16
rect 254 -22 255 -16
rect 198 -22 199 -18
rect 215 -22 216 -18
rect 219 -22 220 -18
rect 240 -22 241 -18
rect 229 -22 230 -20
rect 236 -21 237 -11
rect 128 -32 129 -30
rect 145 -49 146 -31
rect 198 -32 199 -30
rect 219 -49 220 -31
rect 222 -49 223 -31
rect 261 -49 262 -31
rect 268 -49 269 -31
rect 289 -49 290 -31
rect 296 -32 297 -30
rect 303 -49 304 -31
rect 324 -49 325 -31
rect 331 -32 332 -30
rect 135 -34 136 -30
rect 152 -34 153 -30
rect 198 -49 199 -33
rect 247 -49 248 -33
rect 327 -34 328 -30
rect 331 -49 332 -33
rect 135 -49 136 -35
rect 152 -49 153 -35
rect 201 -49 202 -35
rect 233 -36 234 -30
rect 142 -38 143 -30
rect 159 -38 160 -30
rect 173 -49 174 -37
rect 233 -49 234 -37
rect 159 -49 160 -39
rect 177 -40 178 -30
rect 205 -40 206 -30
rect 226 -40 227 -30
rect 163 -42 164 -30
rect 177 -49 178 -41
rect 205 -49 206 -41
rect 240 -42 241 -30
rect 163 -49 164 -43
rect 184 -49 185 -43
rect 208 -49 209 -43
rect 212 -49 213 -43
rect 226 -49 227 -43
rect 282 -49 283 -43
rect 229 -46 230 -30
rect 240 -49 241 -45
rect 191 -49 192 -47
rect 229 -49 230 -47
rect 103 -72 104 -58
rect 107 -72 108 -58
rect 121 -72 122 -58
rect 135 -59 136 -57
rect 142 -59 143 -57
rect 163 -72 164 -58
rect 205 -72 206 -58
rect 212 -59 213 -57
rect 226 -72 227 -58
rect 247 -59 248 -57
rect 261 -59 262 -57
rect 313 -72 314 -58
rect 324 -59 325 -57
rect 324 -72 325 -58
rect 324 -59 325 -57
rect 324 -72 325 -58
rect 331 -59 332 -57
rect 331 -72 332 -58
rect 331 -59 332 -57
rect 331 -72 332 -58
rect 128 -72 129 -60
rect 159 -72 160 -60
rect 191 -61 192 -57
rect 261 -72 262 -60
rect 268 -61 269 -57
rect 282 -61 283 -57
rect 289 -61 290 -57
rect 306 -72 307 -60
rect 142 -72 143 -62
rect 149 -72 150 -62
rect 184 -63 185 -57
rect 191 -72 192 -62
rect 229 -63 230 -57
rect 233 -63 234 -57
rect 240 -63 241 -57
rect 254 -63 255 -57
rect 275 -72 276 -62
rect 278 -63 279 -57
rect 282 -72 283 -62
rect 299 -63 300 -57
rect 177 -72 178 -64
rect 184 -72 185 -64
rect 201 -72 202 -64
rect 240 -72 241 -64
rect 296 -65 297 -57
rect 303 -65 304 -57
rect 219 -67 220 -57
rect 254 -72 255 -66
rect 292 -72 293 -66
rect 296 -72 297 -66
rect 170 -69 171 -57
rect 219 -72 220 -68
rect 166 -72 167 -70
rect 170 -72 171 -70
rect 89 -82 90 -80
rect 89 -97 90 -81
rect 89 -82 90 -80
rect 89 -97 90 -81
rect 100 -97 101 -81
rect 107 -82 108 -80
rect 114 -97 115 -81
rect 131 -97 132 -81
rect 138 -82 139 -80
rect 149 -82 150 -80
rect 159 -97 160 -81
rect 163 -97 164 -81
rect 166 -97 167 -81
rect 177 -82 178 -80
rect 184 -97 185 -81
rect 194 -97 195 -81
rect 205 -82 206 -80
rect 212 -97 213 -81
rect 229 -82 230 -80
rect 254 -82 255 -80
rect 275 -82 276 -80
rect 303 -97 304 -81
rect 317 -82 318 -80
rect 324 -82 325 -80
rect 107 -97 108 -83
rect 128 -84 129 -80
rect 149 -97 150 -83
rect 170 -84 171 -80
rect 191 -84 192 -80
rect 198 -84 199 -80
rect 222 -84 223 -80
rect 229 -97 230 -83
rect 233 -97 234 -83
rect 247 -84 248 -80
rect 282 -84 283 -80
rect 292 -84 293 -80
rect 296 -84 297 -80
rect 310 -97 311 -83
rect 317 -97 318 -83
rect 320 -84 321 -80
rect 324 -97 325 -83
rect 331 -84 332 -80
rect 121 -86 122 -80
rect 145 -86 146 -80
rect 198 -97 199 -85
rect 215 -86 216 -80
rect 219 -97 220 -85
rect 247 -97 248 -85
rect 117 -88 118 -80
rect 121 -97 122 -87
rect 128 -97 129 -87
rect 135 -97 136 -87
rect 142 -88 143 -80
rect 145 -97 146 -87
rect 222 -97 223 -87
rect 296 -97 297 -87
rect 226 -97 227 -89
rect 254 -97 255 -89
rect 236 -92 237 -80
rect 261 -92 262 -80
rect 240 -94 241 -80
rect 275 -97 276 -93
rect 261 -97 262 -95
rect 271 -96 272 -80
rect 86 -122 87 -106
rect 103 -107 104 -105
rect 107 -107 108 -105
rect 128 -107 129 -105
rect 135 -107 136 -105
rect 145 -122 146 -106
rect 149 -107 150 -105
rect 180 -107 181 -105
rect 198 -107 199 -105
rect 219 -107 220 -105
rect 229 -107 230 -105
rect 275 -107 276 -105
rect 282 -107 283 -105
rect 296 -107 297 -105
rect 380 -122 381 -106
rect 383 -107 384 -105
rect 114 -109 115 -105
rect 124 -109 125 -105
rect 135 -122 136 -108
rect 163 -109 164 -105
rect 198 -122 199 -108
rect 212 -109 213 -105
rect 215 -109 216 -105
rect 233 -109 234 -105
rect 240 -109 241 -105
rect 240 -122 241 -108
rect 240 -109 241 -105
rect 240 -122 241 -108
rect 243 -109 244 -105
rect 303 -109 304 -105
rect 103 -122 104 -110
rect 114 -122 115 -110
rect 156 -122 157 -110
rect 184 -111 185 -105
rect 205 -111 206 -105
rect 236 -122 237 -110
rect 247 -111 248 -105
rect 271 -111 272 -105
rect 289 -111 290 -105
rect 310 -111 311 -105
rect 107 -122 108 -112
rect 124 -122 125 -112
rect 163 -122 164 -112
rect 170 -113 171 -105
rect 177 -113 178 -105
rect 215 -122 216 -112
rect 268 -113 269 -105
rect 317 -113 318 -105
rect 180 -122 181 -114
rect 205 -122 206 -114
rect 208 -115 209 -105
rect 219 -122 220 -114
rect 261 -115 262 -105
rect 268 -122 269 -114
rect 303 -122 304 -114
rect 324 -115 325 -105
rect 184 -122 185 -116
rect 191 -122 192 -116
rect 212 -122 213 -116
rect 299 -122 300 -116
rect 310 -122 311 -116
rect 317 -122 318 -116
rect 254 -119 255 -105
rect 261 -122 262 -118
rect 226 -122 227 -120
rect 254 -122 255 -120
rect 79 -132 80 -130
rect 82 -147 83 -131
rect 107 -132 108 -130
rect 142 -147 143 -131
rect 156 -132 157 -130
rect 194 -132 195 -130
rect 198 -132 199 -130
rect 198 -147 199 -131
rect 198 -132 199 -130
rect 198 -147 199 -131
rect 219 -132 220 -130
rect 233 -147 234 -131
rect 257 -147 258 -131
rect 261 -132 262 -130
rect 268 -132 269 -130
rect 271 -147 272 -131
rect 296 -132 297 -130
rect 303 -132 304 -130
rect 310 -147 311 -131
rect 317 -132 318 -130
rect 380 -132 381 -130
rect 387 -147 388 -131
rect 79 -147 80 -133
rect 86 -134 87 -130
rect 107 -147 108 -133
rect 117 -134 118 -130
rect 131 -134 132 -130
rect 138 -147 139 -133
rect 159 -147 160 -133
rect 215 -134 216 -130
rect 226 -147 227 -133
rect 268 -147 269 -133
rect 275 -147 276 -133
rect 317 -147 318 -133
rect 114 -147 115 -135
rect 121 -136 122 -130
rect 128 -136 129 -130
rect 131 -147 132 -135
rect 135 -136 136 -130
rect 152 -136 153 -130
rect 163 -136 164 -130
rect 177 -136 178 -130
rect 184 -136 185 -130
rect 229 -136 230 -130
rect 254 -136 255 -130
rect 261 -147 262 -135
rect 299 -136 300 -130
rect 324 -147 325 -135
rect 128 -147 129 -137
rect 156 -147 157 -137
rect 170 -147 171 -137
rect 254 -147 255 -137
rect 145 -147 146 -139
rect 163 -147 164 -139
rect 173 -140 174 -130
rect 177 -147 178 -139
rect 191 -147 192 -139
rect 215 -147 216 -139
rect 121 -147 122 -141
rect 173 -147 174 -141
rect 205 -142 206 -130
rect 219 -147 220 -141
rect 152 -147 153 -143
rect 208 -147 209 -143
rect 205 -147 206 -145
rect 240 -146 241 -130
rect 82 -157 83 -155
rect 82 -170 83 -156
rect 82 -157 83 -155
rect 82 -170 83 -156
rect 107 -157 108 -155
rect 152 -157 153 -155
rect 156 -170 157 -156
rect 163 -157 164 -155
rect 173 -157 174 -155
rect 177 -157 178 -155
rect 187 -157 188 -155
rect 191 -157 192 -155
rect 198 -170 199 -156
rect 226 -157 227 -155
rect 233 -157 234 -155
rect 247 -170 248 -156
rect 254 -157 255 -155
rect 303 -170 304 -156
rect 317 -157 318 -155
rect 341 -170 342 -156
rect 359 -170 360 -156
rect 373 -170 374 -156
rect 387 -157 388 -155
rect 394 -170 395 -156
rect 408 -170 409 -156
rect 415 -170 416 -156
rect 436 -170 437 -156
rect 443 -170 444 -156
rect 114 -159 115 -155
rect 117 -170 118 -158
rect 121 -159 122 -155
rect 135 -159 136 -155
rect 152 -170 153 -158
rect 184 -159 185 -155
rect 212 -159 213 -155
rect 254 -170 255 -158
rect 261 -159 262 -155
rect 271 -159 272 -155
rect 296 -170 297 -158
rect 313 -159 314 -155
rect 317 -170 318 -158
rect 324 -159 325 -155
rect 331 -170 332 -158
rect 352 -170 353 -158
rect 362 -170 363 -158
rect 380 -170 381 -158
rect 383 -159 384 -155
rect 387 -170 388 -158
rect 124 -170 125 -160
rect 138 -161 139 -155
rect 163 -170 164 -160
rect 201 -161 202 -155
rect 205 -161 206 -155
rect 212 -170 213 -160
rect 215 -161 216 -155
rect 219 -161 220 -155
rect 226 -170 227 -160
rect 366 -170 367 -160
rect 135 -170 136 -162
rect 145 -170 146 -162
rect 170 -170 171 -162
rect 191 -170 192 -162
rect 205 -170 206 -162
rect 215 -170 216 -162
rect 219 -170 220 -162
rect 229 -170 230 -162
rect 233 -170 234 -162
rect 289 -170 290 -162
rect 320 -163 321 -155
rect 345 -170 346 -162
rect 177 -170 178 -164
rect 243 -165 244 -155
rect 261 -170 262 -164
rect 275 -165 276 -155
rect 278 -170 279 -164
rect 324 -170 325 -164
rect 240 -170 241 -166
rect 282 -170 283 -166
rect 268 -169 269 -155
rect 383 -170 384 -168
rect 75 -197 76 -179
rect 79 -197 80 -179
rect 86 -197 87 -179
rect 121 -180 122 -178
rect 131 -180 132 -178
rect 131 -197 132 -179
rect 131 -180 132 -178
rect 131 -197 132 -179
rect 135 -180 136 -178
rect 142 -197 143 -179
rect 149 -197 150 -179
rect 198 -180 199 -178
rect 229 -180 230 -178
rect 247 -180 248 -178
rect 250 -197 251 -179
rect 359 -197 360 -179
rect 369 -197 370 -179
rect 387 -180 388 -178
rect 408 -180 409 -178
rect 408 -197 409 -179
rect 408 -180 409 -178
rect 408 -197 409 -179
rect 415 -180 416 -178
rect 422 -197 423 -179
rect 432 -197 433 -179
rect 443 -180 444 -178
rect 89 -197 90 -181
rect 93 -197 94 -181
rect 107 -197 108 -181
rect 128 -197 129 -181
rect 156 -197 157 -181
rect 159 -182 160 -178
rect 163 -182 164 -178
rect 268 -197 269 -181
rect 271 -182 272 -178
rect 324 -182 325 -178
rect 338 -197 339 -181
rect 373 -182 374 -178
rect 383 -197 384 -181
rect 394 -182 395 -178
rect 401 -197 402 -181
rect 415 -197 416 -181
rect 436 -197 437 -181
rect 443 -197 444 -181
rect 121 -197 122 -183
rect 135 -197 136 -183
rect 170 -184 171 -178
rect 212 -197 213 -183
rect 233 -184 234 -178
rect 261 -184 262 -178
rect 289 -184 290 -178
rect 289 -197 290 -183
rect 289 -184 290 -178
rect 289 -197 290 -183
rect 296 -184 297 -178
rect 313 -184 314 -178
rect 317 -184 318 -178
rect 355 -184 356 -178
rect 380 -197 381 -183
rect 394 -197 395 -183
rect 170 -197 171 -185
rect 219 -186 220 -178
rect 229 -197 230 -185
rect 233 -197 234 -185
rect 254 -186 255 -178
rect 275 -186 276 -178
rect 303 -186 304 -178
rect 310 -197 311 -185
rect 317 -197 318 -185
rect 331 -186 332 -178
rect 345 -186 346 -178
rect 373 -197 374 -185
rect 177 -188 178 -178
rect 215 -197 216 -187
rect 219 -197 220 -187
rect 275 -197 276 -187
rect 285 -188 286 -178
rect 345 -197 346 -187
rect 177 -197 178 -189
rect 184 -190 185 -178
rect 191 -197 192 -189
rect 205 -190 206 -178
rect 254 -197 255 -189
rect 282 -197 283 -189
rect 285 -197 286 -189
rect 352 -197 353 -189
rect 163 -197 164 -191
rect 205 -197 206 -191
rect 261 -197 262 -191
rect 324 -197 325 -191
rect 331 -197 332 -191
rect 366 -192 367 -178
rect 184 -197 185 -193
rect 240 -194 241 -178
rect 296 -197 297 -193
rect 303 -197 304 -193
rect 201 -197 202 -195
rect 240 -197 241 -195
rect 72 -230 73 -206
rect 96 -207 97 -205
rect 100 -230 101 -206
rect 121 -207 122 -205
rect 128 -230 129 -206
rect 226 -230 227 -206
rect 261 -230 262 -206
rect 331 -207 332 -205
rect 345 -207 346 -205
rect 387 -230 388 -206
rect 394 -207 395 -205
rect 401 -207 402 -205
rect 404 -207 405 -205
rect 408 -207 409 -205
rect 415 -207 416 -205
rect 422 -230 423 -206
rect 436 -207 437 -205
rect 439 -230 440 -206
rect 79 -209 80 -205
rect 86 -209 87 -205
rect 103 -209 104 -205
rect 107 -209 108 -205
rect 114 -209 115 -205
rect 114 -230 115 -208
rect 114 -209 115 -205
rect 114 -230 115 -208
rect 121 -230 122 -208
rect 247 -209 248 -205
rect 268 -209 269 -205
rect 303 -230 304 -208
rect 306 -209 307 -205
rect 317 -209 318 -205
rect 373 -209 374 -205
rect 383 -209 384 -205
rect 79 -230 80 -210
rect 145 -211 146 -205
rect 149 -211 150 -205
rect 229 -211 230 -205
rect 236 -230 237 -210
rect 345 -230 346 -210
rect 373 -230 374 -210
rect 380 -211 381 -205
rect 86 -230 87 -212
rect 187 -230 188 -212
rect 191 -213 192 -205
rect 219 -213 220 -205
rect 222 -230 223 -212
rect 240 -213 241 -205
rect 257 -230 258 -212
rect 268 -230 269 -212
rect 275 -213 276 -205
rect 317 -230 318 -212
rect 359 -213 360 -205
rect 380 -230 381 -212
rect 93 -230 94 -214
rect 149 -230 150 -214
rect 156 -215 157 -205
rect 180 -230 181 -214
rect 198 -230 199 -214
rect 247 -230 248 -214
rect 289 -215 290 -205
rect 289 -230 290 -214
rect 289 -215 290 -205
rect 289 -230 290 -214
rect 310 -215 311 -205
rect 331 -230 332 -214
rect 107 -230 108 -216
rect 219 -230 220 -216
rect 229 -230 230 -216
rect 338 -217 339 -205
rect 142 -230 143 -218
rect 163 -219 164 -205
rect 170 -219 171 -205
rect 264 -219 265 -205
rect 296 -219 297 -205
rect 310 -230 311 -218
rect 324 -219 325 -205
rect 338 -230 339 -218
rect 159 -230 160 -220
rect 191 -230 192 -220
rect 201 -230 202 -220
rect 275 -230 276 -220
rect 324 -230 325 -220
rect 352 -221 353 -205
rect 170 -230 171 -222
rect 177 -223 178 -205
rect 205 -223 206 -205
rect 254 -223 255 -205
rect 352 -230 353 -222
rect 369 -223 370 -205
rect 131 -225 132 -205
rect 177 -230 178 -224
rect 184 -225 185 -205
rect 205 -230 206 -224
rect 212 -225 213 -205
rect 296 -230 297 -224
rect 212 -230 213 -226
rect 233 -227 234 -205
rect 240 -230 241 -226
rect 359 -230 360 -226
rect 233 -230 234 -228
rect 282 -230 283 -228
rect 68 -240 69 -238
rect 156 -240 157 -238
rect 170 -240 171 -238
rect 187 -240 188 -238
rect 229 -273 230 -239
rect 317 -240 318 -238
rect 359 -240 360 -238
rect 443 -273 444 -239
rect 450 -273 451 -239
rect 457 -273 458 -239
rect 530 -273 531 -239
rect 534 -273 535 -239
rect 86 -242 87 -238
rect 159 -242 160 -238
rect 170 -273 171 -241
rect 205 -242 206 -238
rect 240 -242 241 -238
rect 275 -242 276 -238
rect 292 -273 293 -241
rect 359 -273 360 -241
rect 366 -242 367 -238
rect 453 -273 454 -241
rect 79 -244 80 -238
rect 205 -273 206 -243
rect 243 -244 244 -238
rect 303 -244 304 -238
rect 331 -244 332 -238
rect 366 -273 367 -243
rect 369 -244 370 -238
rect 387 -244 388 -238
rect 394 -273 395 -243
rect 439 -273 440 -243
rect 72 -273 73 -245
rect 79 -273 80 -245
rect 93 -246 94 -238
rect 184 -273 185 -245
rect 194 -273 195 -245
rect 240 -273 241 -245
rect 250 -246 251 -238
rect 345 -246 346 -238
rect 418 -246 419 -238
rect 422 -246 423 -238
rect 93 -273 94 -247
rect 212 -248 213 -238
rect 254 -248 255 -238
rect 264 -248 265 -238
rect 271 -273 272 -247
rect 338 -248 339 -238
rect 345 -273 346 -247
rect 352 -248 353 -238
rect 373 -248 374 -238
rect 422 -273 423 -247
rect 100 -250 101 -238
rect 135 -250 136 -238
rect 138 -250 139 -238
rect 187 -273 188 -249
rect 208 -273 209 -249
rect 373 -273 374 -249
rect 408 -273 409 -249
rect 418 -273 419 -249
rect 107 -252 108 -238
rect 166 -252 167 -238
rect 177 -273 178 -251
rect 191 -252 192 -238
rect 212 -273 213 -251
rect 247 -273 248 -251
rect 254 -273 255 -251
rect 380 -273 381 -251
rect 107 -273 108 -253
rect 114 -254 115 -238
rect 121 -254 122 -238
rect 226 -254 227 -238
rect 257 -273 258 -253
rect 317 -273 318 -253
rect 338 -273 339 -253
rect 415 -273 416 -253
rect 114 -273 115 -255
rect 145 -273 146 -255
rect 180 -256 181 -238
rect 233 -273 234 -255
rect 261 -256 262 -238
rect 324 -273 325 -255
rect 121 -273 122 -257
rect 149 -258 150 -238
rect 198 -273 199 -257
rect 226 -273 227 -257
rect 261 -273 262 -257
rect 268 -258 269 -238
rect 275 -273 276 -257
rect 299 -273 300 -257
rect 303 -273 304 -257
rect 387 -273 388 -257
rect 128 -260 129 -238
rect 163 -273 164 -259
rect 268 -273 269 -259
rect 331 -273 332 -259
rect 131 -273 132 -261
rect 215 -273 216 -261
rect 296 -262 297 -238
rect 429 -273 430 -261
rect 135 -273 136 -263
rect 156 -273 157 -263
rect 296 -273 297 -263
rect 401 -273 402 -263
rect 142 -266 143 -238
rect 152 -266 153 -238
rect 310 -266 311 -238
rect 352 -273 353 -265
rect 86 -273 87 -267
rect 152 -273 153 -267
rect 219 -268 220 -238
rect 310 -273 311 -267
rect 149 -273 150 -269
rect 282 -270 283 -238
rect 282 -273 283 -271
rect 289 -272 290 -238
rect 30 -283 31 -281
rect 37 -283 38 -281
rect 47 -314 48 -282
rect 149 -283 150 -281
rect 177 -283 178 -281
rect 212 -314 213 -282
rect 222 -283 223 -281
rect 261 -283 262 -281
rect 268 -283 269 -281
rect 401 -283 402 -281
rect 415 -283 416 -281
rect 436 -314 437 -282
rect 453 -314 454 -282
rect 457 -283 458 -281
rect 527 -314 528 -282
rect 534 -283 535 -281
rect 30 -314 31 -284
rect 33 -285 34 -281
rect 51 -314 52 -284
rect 54 -285 55 -281
rect 58 -314 59 -284
rect 131 -285 132 -281
rect 135 -314 136 -284
rect 163 -285 164 -281
rect 184 -285 185 -281
rect 219 -285 220 -281
rect 243 -314 244 -284
rect 450 -285 451 -281
rect 68 -314 69 -286
rect 184 -314 185 -286
rect 194 -287 195 -281
rect 394 -287 395 -281
rect 401 -314 402 -286
rect 422 -287 423 -281
rect 75 -314 76 -288
rect 79 -289 80 -281
rect 82 -314 83 -288
rect 191 -314 192 -288
rect 205 -314 206 -288
rect 219 -314 220 -288
rect 247 -289 248 -281
rect 289 -314 290 -288
rect 292 -289 293 -281
rect 366 -289 367 -281
rect 387 -289 388 -281
rect 422 -314 423 -288
rect 86 -314 87 -290
rect 103 -291 104 -281
rect 107 -291 108 -281
rect 121 -291 122 -281
rect 149 -314 150 -290
rect 170 -291 171 -281
rect 208 -314 209 -290
rect 240 -291 241 -281
rect 254 -291 255 -281
rect 352 -291 353 -281
rect 380 -291 381 -281
rect 387 -314 388 -290
rect 394 -314 395 -290
rect 408 -291 409 -281
rect 93 -293 94 -281
rect 261 -314 262 -292
rect 268 -314 269 -292
rect 275 -293 276 -281
rect 282 -293 283 -281
rect 303 -314 304 -292
rect 306 -293 307 -281
rect 310 -293 311 -281
rect 338 -293 339 -281
rect 366 -314 367 -292
rect 408 -314 409 -292
rect 418 -314 419 -292
rect 93 -314 94 -294
rect 114 -295 115 -281
rect 121 -314 122 -294
rect 145 -314 146 -294
rect 156 -295 157 -281
rect 177 -314 178 -294
rect 226 -295 227 -281
rect 275 -314 276 -294
rect 296 -295 297 -281
rect 429 -295 430 -281
rect 100 -314 101 -296
rect 152 -297 153 -281
rect 163 -314 164 -296
rect 324 -297 325 -281
rect 352 -314 353 -296
rect 376 -314 377 -296
rect 114 -314 115 -298
rect 198 -299 199 -281
rect 226 -314 227 -298
rect 247 -314 248 -298
rect 299 -314 300 -298
rect 443 -299 444 -281
rect 128 -314 129 -300
rect 282 -314 283 -300
rect 310 -314 311 -300
rect 317 -301 318 -281
rect 142 -314 143 -302
rect 296 -314 297 -302
rect 317 -314 318 -302
rect 345 -303 346 -281
rect 170 -314 171 -304
rect 338 -314 339 -304
rect 198 -314 199 -306
rect 233 -307 234 -281
rect 331 -307 332 -281
rect 345 -314 346 -306
rect 187 -309 188 -281
rect 233 -314 234 -308
rect 331 -314 332 -308
rect 359 -309 360 -281
rect 229 -314 230 -310
rect 380 -314 381 -310
rect 359 -314 360 -312
rect 373 -313 374 -281
rect 19 -361 20 -323
rect 23 -361 24 -323
rect 37 -361 38 -323
rect 93 -324 94 -322
rect 96 -361 97 -323
rect 166 -361 167 -323
rect 194 -324 195 -322
rect 275 -324 276 -322
rect 282 -324 283 -322
rect 366 -324 367 -322
rect 373 -324 374 -322
rect 471 -361 472 -323
rect 513 -361 514 -323
rect 520 -324 521 -322
rect 523 -324 524 -322
rect 527 -324 528 -322
rect 51 -361 52 -325
rect 201 -361 202 -325
rect 219 -326 220 -322
rect 296 -361 297 -325
rect 324 -326 325 -322
rect 324 -361 325 -325
rect 324 -326 325 -322
rect 324 -361 325 -325
rect 327 -361 328 -325
rect 331 -326 332 -322
rect 408 -326 409 -322
rect 415 -361 416 -325
rect 422 -326 423 -322
rect 457 -361 458 -325
rect 58 -328 59 -322
rect 107 -328 108 -322
rect 110 -328 111 -322
rect 138 -361 139 -327
rect 145 -361 146 -327
rect 156 -361 157 -327
rect 159 -328 160 -322
rect 177 -328 178 -322
rect 198 -328 199 -322
rect 243 -328 244 -322
rect 247 -328 248 -322
rect 317 -328 318 -322
rect 331 -361 332 -327
rect 380 -328 381 -322
rect 390 -361 391 -327
rect 408 -361 409 -327
rect 436 -328 437 -322
rect 467 -361 468 -327
rect 58 -361 59 -329
rect 86 -330 87 -322
rect 100 -330 101 -322
rect 149 -330 150 -322
rect 177 -361 178 -329
rect 184 -330 185 -322
rect 198 -361 199 -329
rect 380 -361 381 -329
rect 387 -330 388 -322
rect 436 -361 437 -329
rect 65 -361 66 -331
rect 135 -332 136 -322
rect 149 -361 150 -331
rect 170 -332 171 -322
rect 184 -361 185 -331
rect 250 -332 251 -322
rect 254 -332 255 -322
rect 366 -361 367 -331
rect 401 -332 402 -322
rect 422 -361 423 -331
rect 82 -334 83 -322
rect 142 -334 143 -322
rect 212 -334 213 -322
rect 219 -361 220 -333
rect 243 -361 244 -333
rect 338 -334 339 -322
rect 72 -361 73 -335
rect 82 -361 83 -335
rect 86 -361 87 -335
rect 121 -336 122 -322
rect 124 -361 125 -335
rect 215 -361 216 -335
rect 250 -361 251 -335
rect 303 -336 304 -322
rect 100 -361 101 -337
rect 107 -361 108 -337
rect 110 -361 111 -337
rect 152 -338 153 -322
rect 163 -338 164 -322
rect 212 -361 213 -337
rect 261 -361 262 -337
rect 310 -338 311 -322
rect 114 -340 115 -322
rect 226 -361 227 -339
rect 264 -340 265 -322
rect 373 -361 374 -339
rect 44 -361 45 -341
rect 114 -361 115 -341
rect 117 -361 118 -341
rect 205 -361 206 -341
rect 264 -361 265 -341
rect 443 -361 444 -341
rect 128 -344 129 -322
rect 229 -344 230 -322
rect 268 -344 269 -322
rect 271 -361 272 -343
rect 285 -344 286 -322
rect 289 -344 290 -322
rect 299 -344 300 -322
rect 401 -361 402 -343
rect 131 -361 132 -345
rect 135 -361 136 -345
rect 194 -361 195 -345
rect 338 -361 339 -345
rect 233 -348 234 -322
rect 285 -361 286 -347
rect 289 -361 290 -347
rect 306 -361 307 -347
rect 310 -361 311 -347
rect 359 -348 360 -322
rect 170 -361 171 -349
rect 233 -361 234 -349
rect 352 -350 353 -322
rect 359 -361 360 -349
rect 345 -352 346 -322
rect 352 -361 353 -351
rect 345 -361 346 -353
rect 429 -354 430 -322
rect 394 -356 395 -322
rect 429 -361 430 -355
rect 240 -358 241 -322
rect 394 -361 395 -357
rect 240 -361 241 -359
rect 450 -361 451 -359
rect 16 -371 17 -369
rect 16 -412 17 -370
rect 16 -371 17 -369
rect 16 -412 17 -370
rect 23 -412 24 -370
rect 100 -371 101 -369
rect 121 -412 122 -370
rect 152 -412 153 -370
rect 198 -412 199 -370
rect 271 -371 272 -369
rect 275 -371 276 -369
rect 436 -371 437 -369
rect 443 -371 444 -369
rect 527 -412 528 -370
rect 30 -373 31 -369
rect 117 -373 118 -369
rect 135 -373 136 -369
rect 166 -373 167 -369
rect 219 -373 220 -369
rect 219 -412 220 -372
rect 219 -373 220 -369
rect 219 -412 220 -372
rect 226 -373 227 -369
rect 303 -412 304 -372
rect 317 -373 318 -369
rect 366 -373 367 -369
rect 387 -373 388 -369
rect 457 -373 458 -369
rect 481 -412 482 -372
rect 499 -412 500 -372
rect 513 -373 514 -369
rect 513 -412 514 -372
rect 513 -373 514 -369
rect 513 -412 514 -372
rect 30 -412 31 -374
rect 173 -375 174 -369
rect 226 -412 227 -374
rect 310 -375 311 -369
rect 331 -375 332 -369
rect 457 -412 458 -374
rect 37 -377 38 -369
rect 114 -377 115 -369
rect 128 -412 129 -376
rect 166 -412 167 -376
rect 233 -377 234 -369
rect 278 -377 279 -369
rect 282 -377 283 -369
rect 464 -412 465 -376
rect 44 -379 45 -369
rect 124 -379 125 -369
rect 138 -412 139 -378
rect 170 -412 171 -378
rect 233 -412 234 -378
rect 313 -412 314 -378
rect 338 -379 339 -369
rect 387 -412 388 -378
rect 390 -379 391 -369
rect 415 -379 416 -369
rect 418 -412 419 -378
rect 520 -412 521 -378
rect 44 -412 45 -380
rect 103 -412 104 -380
rect 149 -381 150 -369
rect 215 -412 216 -380
rect 240 -381 241 -369
rect 296 -381 297 -369
rect 310 -412 311 -380
rect 401 -381 402 -369
rect 415 -412 416 -380
rect 443 -412 444 -380
rect 450 -381 451 -369
rect 492 -412 493 -380
rect 51 -383 52 -369
rect 100 -412 101 -382
rect 243 -383 244 -369
rect 345 -383 346 -369
rect 348 -412 349 -382
rect 366 -412 367 -382
rect 394 -383 395 -369
rect 506 -412 507 -382
rect 58 -385 59 -369
rect 110 -385 111 -369
rect 254 -385 255 -369
rect 282 -412 283 -384
rect 296 -412 297 -384
rect 320 -385 321 -369
rect 352 -385 353 -369
rect 401 -412 402 -384
rect 408 -385 409 -369
rect 450 -412 451 -384
rect 58 -412 59 -386
rect 159 -412 160 -386
rect 254 -412 255 -386
rect 289 -387 290 -369
rect 352 -412 353 -386
rect 471 -387 472 -369
rect 65 -389 66 -369
rect 191 -389 192 -369
rect 250 -389 251 -369
rect 471 -412 472 -388
rect 65 -412 66 -390
rect 82 -391 83 -369
rect 86 -412 87 -390
rect 208 -412 209 -390
rect 261 -391 262 -369
rect 380 -391 381 -369
rect 408 -412 409 -390
rect 422 -391 423 -369
rect 72 -393 73 -369
rect 93 -393 94 -369
rect 110 -412 111 -392
rect 247 -393 248 -369
rect 261 -412 262 -392
rect 394 -412 395 -392
rect 72 -412 73 -394
rect 212 -395 213 -369
rect 268 -395 269 -369
rect 429 -395 430 -369
rect 79 -412 80 -396
rect 107 -397 108 -369
rect 131 -397 132 -369
rect 289 -412 290 -396
rect 324 -397 325 -369
rect 422 -412 423 -396
rect 37 -412 38 -398
rect 107 -412 108 -398
rect 114 -412 115 -398
rect 324 -412 325 -398
rect 359 -399 360 -369
rect 380 -412 381 -398
rect 89 -401 90 -369
rect 142 -401 143 -369
rect 156 -401 157 -369
rect 191 -412 192 -400
rect 212 -412 213 -400
rect 331 -412 332 -400
rect 373 -401 374 -369
rect 429 -412 430 -400
rect 93 -412 94 -402
rect 184 -403 185 -369
rect 229 -412 230 -402
rect 359 -412 360 -402
rect 156 -412 157 -404
rect 436 -412 437 -404
rect 177 -407 178 -369
rect 247 -412 248 -406
rect 275 -412 276 -406
rect 327 -412 328 -406
rect 177 -412 178 -408
rect 194 -412 195 -408
rect 240 -412 241 -408
rect 268 -412 269 -408
rect 317 -412 318 -408
rect 373 -412 374 -408
rect 184 -412 185 -410
rect 205 -411 206 -369
rect 16 -463 17 -421
rect 79 -422 80 -420
rect 86 -422 87 -420
rect 89 -462 90 -421
rect 93 -422 94 -420
rect 215 -422 216 -420
rect 233 -422 234 -420
rect 233 -463 234 -421
rect 233 -422 234 -420
rect 233 -463 234 -421
rect 247 -422 248 -420
rect 264 -422 265 -420
rect 268 -463 269 -421
rect 282 -463 283 -421
rect 289 -422 290 -420
rect 292 -462 293 -421
rect 324 -422 325 -420
rect 499 -422 500 -420
rect 513 -422 514 -420
rect 513 -463 514 -421
rect 513 -422 514 -420
rect 513 -463 514 -421
rect 520 -422 521 -420
rect 548 -463 549 -421
rect 30 -424 31 -420
rect 145 -424 146 -420
rect 159 -463 160 -423
rect 457 -424 458 -420
rect 464 -424 465 -420
rect 541 -463 542 -423
rect 30 -463 31 -425
rect 110 -426 111 -420
rect 114 -426 115 -420
rect 212 -463 213 -425
rect 219 -426 220 -420
rect 247 -463 248 -425
rect 254 -426 255 -420
rect 324 -463 325 -425
rect 327 -426 328 -420
rect 408 -426 409 -420
rect 415 -426 416 -420
rect 576 -463 577 -425
rect 44 -463 45 -427
rect 222 -463 223 -427
rect 240 -428 241 -420
rect 254 -463 255 -427
rect 261 -428 262 -420
rect 492 -428 493 -420
rect 527 -428 528 -420
rect 562 -463 563 -427
rect 2 -463 3 -429
rect 240 -463 241 -429
rect 278 -463 279 -429
rect 296 -430 297 -420
rect 331 -430 332 -420
rect 331 -463 332 -429
rect 331 -430 332 -420
rect 331 -463 332 -429
rect 338 -463 339 -429
rect 485 -430 486 -420
rect 51 -432 52 -420
rect 54 -463 55 -431
rect 58 -463 59 -431
rect 121 -432 122 -420
rect 128 -432 129 -420
rect 201 -463 202 -431
rect 219 -463 220 -431
rect 499 -463 500 -431
rect 37 -463 38 -433
rect 121 -463 122 -433
rect 135 -463 136 -433
rect 166 -463 167 -433
rect 173 -463 174 -433
rect 464 -463 465 -433
rect 471 -434 472 -420
rect 478 -463 479 -433
rect 65 -463 66 -435
rect 198 -436 199 -420
rect 226 -436 227 -420
rect 527 -463 528 -435
rect 72 -438 73 -420
rect 320 -438 321 -420
rect 341 -438 342 -420
rect 401 -438 402 -420
rect 429 -438 430 -420
rect 520 -463 521 -437
rect 72 -463 73 -439
rect 170 -440 171 -420
rect 191 -463 192 -439
rect 275 -440 276 -420
rect 285 -440 286 -420
rect 471 -463 472 -439
rect 9 -463 10 -441
rect 170 -463 171 -441
rect 177 -442 178 -420
rect 285 -463 286 -441
rect 289 -463 290 -441
rect 303 -442 304 -420
rect 348 -463 349 -441
rect 485 -463 486 -441
rect 79 -463 80 -443
rect 345 -463 346 -443
rect 352 -444 353 -420
rect 408 -463 409 -443
rect 436 -444 437 -420
rect 534 -463 535 -443
rect 86 -463 87 -445
rect 198 -463 199 -445
rect 229 -446 230 -420
rect 296 -463 297 -445
rect 313 -463 314 -445
rect 359 -446 360 -420
rect 457 -463 458 -445
rect 96 -463 97 -447
rect 100 -463 101 -447
rect 107 -463 108 -447
rect 142 -448 143 -420
rect 177 -463 178 -447
rect 243 -463 244 -447
rect 366 -448 367 -420
rect 401 -463 402 -447
rect 436 -463 437 -447
rect 443 -448 444 -420
rect 450 -448 451 -420
rect 450 -463 451 -447
rect 450 -448 451 -420
rect 450 -463 451 -447
rect 142 -463 143 -449
rect 359 -463 360 -449
rect 380 -450 381 -420
rect 429 -463 430 -449
rect 443 -463 444 -449
rect 506 -450 507 -420
rect 23 -452 24 -420
rect 506 -463 507 -451
rect 205 -463 206 -453
rect 352 -463 353 -453
rect 373 -454 374 -420
rect 380 -463 381 -453
rect 387 -454 388 -420
rect 492 -463 493 -453
rect 229 -463 230 -455
rect 415 -463 416 -455
rect 275 -463 276 -457
rect 387 -463 388 -457
rect 394 -458 395 -420
rect 397 -458 398 -420
rect 394 -463 395 -459
rect 422 -460 423 -420
rect 397 -463 398 -461
rect 422 -463 423 -461
rect 9 -473 10 -471
rect 121 -473 122 -471
rect 131 -473 132 -471
rect 191 -473 192 -471
rect 219 -473 220 -471
rect 247 -473 248 -471
rect 275 -520 276 -472
rect 471 -473 472 -471
rect 513 -473 514 -471
rect 513 -520 514 -472
rect 513 -473 514 -471
rect 513 -520 514 -472
rect 555 -473 556 -471
rect 562 -473 563 -471
rect 16 -475 17 -471
rect 117 -520 118 -474
rect 152 -475 153 -471
rect 177 -475 178 -471
rect 184 -475 185 -471
rect 313 -475 314 -471
rect 355 -520 356 -474
rect 534 -475 535 -471
rect 558 -475 559 -471
rect 562 -520 563 -474
rect 16 -520 17 -476
rect 93 -477 94 -471
rect 100 -477 101 -471
rect 100 -520 101 -476
rect 100 -477 101 -471
rect 100 -520 101 -476
rect 107 -477 108 -471
rect 278 -477 279 -471
rect 282 -477 283 -471
rect 471 -520 472 -476
rect 23 -479 24 -471
rect 149 -479 150 -471
rect 159 -520 160 -478
rect 422 -479 423 -471
rect 425 -520 426 -478
rect 485 -479 486 -471
rect 30 -520 31 -480
rect 54 -481 55 -471
rect 58 -481 59 -471
rect 96 -481 97 -471
rect 107 -520 108 -480
rect 233 -481 234 -471
rect 240 -481 241 -471
rect 338 -481 339 -471
rect 359 -481 360 -471
rect 541 -481 542 -471
rect 37 -483 38 -471
rect 240 -520 241 -482
rect 285 -483 286 -471
rect 408 -483 409 -471
rect 464 -483 465 -471
rect 572 -483 573 -471
rect 2 -485 3 -471
rect 285 -520 286 -484
rect 299 -520 300 -484
rect 359 -520 360 -484
rect 373 -485 374 -471
rect 457 -485 458 -471
rect 541 -520 542 -484
rect 548 -485 549 -471
rect 37 -520 38 -486
rect 114 -487 115 -471
rect 142 -487 143 -471
rect 149 -520 150 -486
rect 163 -487 164 -471
rect 506 -487 507 -471
rect 44 -489 45 -471
rect 124 -489 125 -471
rect 135 -489 136 -471
rect 163 -520 164 -488
rect 170 -489 171 -471
rect 177 -520 178 -488
rect 184 -520 185 -488
rect 268 -489 269 -471
rect 303 -489 304 -471
rect 317 -489 318 -471
rect 331 -489 332 -471
rect 338 -520 339 -488
rect 394 -489 395 -471
rect 485 -520 486 -488
rect 51 -520 52 -490
rect 345 -520 346 -490
rect 380 -491 381 -471
rect 394 -520 395 -490
rect 408 -520 409 -490
rect 415 -491 416 -471
rect 436 -491 437 -471
rect 464 -520 465 -490
rect 72 -493 73 -471
rect 229 -493 230 -471
rect 233 -520 234 -492
rect 369 -520 370 -492
rect 380 -520 381 -492
rect 401 -493 402 -471
rect 457 -520 458 -492
rect 499 -493 500 -471
rect 44 -520 45 -494
rect 229 -520 230 -494
rect 289 -495 290 -471
rect 303 -520 304 -494
rect 310 -495 311 -471
rect 527 -495 528 -471
rect 75 -520 76 -496
rect 93 -520 94 -496
rect 124 -520 125 -496
rect 219 -520 220 -496
rect 222 -520 223 -496
rect 576 -497 577 -471
rect 86 -499 87 -471
rect 264 -499 265 -471
rect 289 -520 290 -498
rect 296 -499 297 -471
rect 310 -520 311 -498
rect 324 -499 325 -471
rect 331 -520 332 -498
rect 450 -499 451 -471
rect 82 -520 83 -500
rect 86 -520 87 -500
rect 89 -520 90 -500
rect 128 -501 129 -471
rect 156 -501 157 -471
rect 415 -520 416 -500
rect 429 -501 430 -471
rect 450 -520 451 -500
rect 170 -520 171 -502
rect 243 -520 244 -502
rect 264 -520 265 -502
rect 268 -520 269 -502
rect 296 -520 297 -502
rect 492 -503 493 -471
rect 191 -520 192 -504
rect 261 -505 262 -471
rect 320 -505 321 -471
rect 401 -520 402 -504
rect 429 -520 430 -504
rect 443 -505 444 -471
rect 478 -505 479 -471
rect 492 -520 493 -504
rect 65 -507 66 -471
rect 261 -520 262 -506
rect 282 -520 283 -506
rect 478 -520 479 -506
rect 58 -520 59 -508
rect 65 -520 66 -508
rect 201 -509 202 -471
rect 247 -520 248 -508
rect 292 -520 293 -508
rect 443 -520 444 -508
rect 201 -520 202 -510
rect 509 -520 510 -510
rect 212 -513 213 -471
rect 317 -520 318 -512
rect 366 -513 367 -471
rect 436 -520 437 -512
rect 205 -515 206 -471
rect 212 -520 213 -514
rect 226 -520 227 -514
rect 254 -520 255 -514
rect 366 -520 367 -514
rect 520 -515 521 -471
rect 79 -517 80 -471
rect 205 -520 206 -516
rect 387 -517 388 -471
rect 520 -520 521 -516
rect 23 -520 24 -518
rect 79 -520 80 -518
rect 390 -520 391 -518
rect 499 -520 500 -518
rect 9 -569 10 -529
rect 16 -530 17 -528
rect 23 -530 24 -528
rect 128 -530 129 -528
rect 131 -530 132 -528
rect 170 -530 171 -528
rect 177 -530 178 -528
rect 187 -530 188 -528
rect 198 -569 199 -529
rect 212 -530 213 -528
rect 215 -569 216 -529
rect 219 -530 220 -528
rect 226 -530 227 -528
rect 499 -530 500 -528
rect 509 -530 510 -528
rect 555 -569 556 -529
rect 562 -530 563 -528
rect 562 -569 563 -529
rect 562 -530 563 -528
rect 562 -569 563 -529
rect 16 -569 17 -531
rect 257 -569 258 -531
rect 268 -532 269 -528
rect 271 -569 272 -531
rect 275 -569 276 -531
rect 369 -569 370 -531
rect 373 -532 374 -528
rect 527 -569 528 -531
rect 541 -532 542 -528
rect 541 -569 542 -531
rect 541 -532 542 -528
rect 541 -569 542 -531
rect 30 -534 31 -528
rect 68 -534 69 -528
rect 79 -569 80 -533
rect 100 -534 101 -528
rect 107 -534 108 -528
rect 177 -569 178 -533
rect 205 -534 206 -528
rect 292 -534 293 -528
rect 296 -569 297 -533
rect 317 -534 318 -528
rect 331 -534 332 -528
rect 366 -569 367 -533
rect 373 -569 374 -533
rect 520 -534 521 -528
rect 30 -569 31 -535
rect 68 -569 69 -535
rect 93 -536 94 -528
rect 93 -569 94 -535
rect 93 -536 94 -528
rect 93 -569 94 -535
rect 103 -569 104 -535
rect 205 -569 206 -535
rect 219 -569 220 -535
rect 513 -536 514 -528
rect 37 -538 38 -528
rect 201 -538 202 -528
rect 247 -538 248 -528
rect 247 -569 248 -537
rect 247 -538 248 -528
rect 247 -569 248 -537
rect 254 -538 255 -528
rect 299 -538 300 -528
rect 306 -569 307 -537
rect 408 -538 409 -528
rect 478 -538 479 -528
rect 534 -569 535 -537
rect 40 -569 41 -539
rect 89 -540 90 -528
rect 107 -569 108 -539
rect 163 -540 164 -528
rect 254 -569 255 -539
rect 387 -569 388 -539
rect 464 -540 465 -528
rect 478 -569 479 -539
rect 485 -540 486 -528
rect 506 -540 507 -528
rect 44 -542 45 -528
rect 138 -542 139 -528
rect 156 -542 157 -528
rect 285 -542 286 -528
rect 289 -569 290 -541
rect 376 -542 377 -528
rect 380 -542 381 -528
rect 380 -569 381 -541
rect 380 -542 381 -528
rect 380 -569 381 -541
rect 492 -542 493 -528
rect 520 -569 521 -541
rect 51 -544 52 -528
rect 184 -569 185 -543
rect 208 -569 209 -543
rect 506 -569 507 -543
rect 51 -569 52 -545
rect 75 -546 76 -528
rect 114 -546 115 -528
rect 261 -546 262 -528
rect 268 -569 269 -545
rect 303 -546 304 -528
rect 313 -546 314 -528
rect 422 -569 423 -545
rect 492 -569 493 -545
rect 530 -569 531 -545
rect 58 -548 59 -528
rect 121 -548 122 -528
rect 124 -548 125 -528
rect 145 -548 146 -528
rect 149 -548 150 -528
rect 156 -569 157 -547
rect 163 -569 164 -547
rect 278 -548 279 -528
rect 282 -569 283 -547
rect 471 -548 472 -528
rect 58 -569 59 -549
rect 72 -569 73 -549
rect 117 -569 118 -549
rect 310 -550 311 -528
rect 313 -569 314 -549
rect 443 -550 444 -528
rect 121 -569 122 -551
rect 222 -569 223 -551
rect 317 -569 318 -551
rect 324 -552 325 -528
rect 331 -569 332 -551
rect 341 -569 342 -551
rect 345 -569 346 -551
rect 450 -552 451 -528
rect 128 -569 129 -553
rect 170 -569 171 -553
rect 229 -569 230 -553
rect 324 -569 325 -553
rect 348 -554 349 -528
rect 436 -554 437 -528
rect 443 -569 444 -553
rect 457 -554 458 -528
rect 135 -569 136 -555
rect 233 -556 234 -528
rect 240 -556 241 -528
rect 436 -569 437 -555
rect 149 -569 150 -557
rect 191 -558 192 -528
rect 240 -569 241 -557
rect 261 -569 262 -557
rect 352 -558 353 -528
rect 471 -569 472 -557
rect 159 -560 160 -528
rect 191 -569 192 -559
rect 338 -560 339 -528
rect 352 -569 353 -559
rect 359 -560 360 -528
rect 408 -569 409 -559
rect 415 -560 416 -528
rect 450 -569 451 -559
rect 142 -569 143 -561
rect 359 -569 360 -561
rect 362 -569 363 -561
rect 464 -569 465 -561
rect 236 -569 237 -563
rect 338 -569 339 -563
rect 394 -564 395 -528
rect 415 -569 416 -563
rect 429 -564 430 -528
rect 457 -569 458 -563
rect 394 -569 395 -565
rect 401 -566 402 -528
rect 429 -569 430 -565
rect 485 -569 486 -565
rect 264 -568 265 -528
rect 401 -569 402 -567
rect 9 -579 10 -577
rect 89 -579 90 -577
rect 93 -579 94 -577
rect 93 -612 94 -578
rect 93 -579 94 -577
rect 93 -612 94 -578
rect 121 -579 122 -577
rect 282 -612 283 -578
rect 289 -579 290 -577
rect 303 -612 304 -578
rect 338 -579 339 -577
rect 394 -579 395 -577
rect 408 -579 409 -577
rect 408 -612 409 -578
rect 408 -579 409 -577
rect 408 -612 409 -578
rect 429 -612 430 -578
rect 450 -579 451 -577
rect 464 -579 465 -577
rect 527 -579 528 -577
rect 530 -579 531 -577
rect 541 -579 542 -577
rect 555 -579 556 -577
rect 555 -612 556 -578
rect 555 -579 556 -577
rect 555 -612 556 -578
rect 562 -579 563 -577
rect 562 -612 563 -578
rect 562 -579 563 -577
rect 562 -612 563 -578
rect 9 -612 10 -580
rect 110 -581 111 -577
rect 121 -612 122 -580
rect 131 -612 132 -580
rect 135 -581 136 -577
rect 212 -612 213 -580
rect 222 -612 223 -580
rect 331 -581 332 -577
rect 338 -612 339 -580
rect 345 -581 346 -577
rect 359 -581 360 -577
rect 415 -581 416 -577
rect 432 -581 433 -577
rect 520 -581 521 -577
rect 534 -581 535 -577
rect 548 -581 549 -577
rect 23 -583 24 -577
rect 58 -583 59 -577
rect 72 -583 73 -577
rect 82 -612 83 -582
rect 86 -583 87 -577
rect 226 -612 227 -582
rect 233 -583 234 -577
rect 247 -583 248 -577
rect 254 -612 255 -582
rect 275 -583 276 -577
rect 324 -583 325 -577
rect 331 -612 332 -582
rect 341 -612 342 -582
rect 345 -612 346 -582
rect 352 -583 353 -577
rect 359 -612 360 -582
rect 366 -612 367 -582
rect 380 -583 381 -577
rect 436 -583 437 -577
rect 499 -583 500 -577
rect 520 -612 521 -582
rect 541 -612 542 -582
rect 23 -612 24 -584
rect 100 -585 101 -577
rect 135 -612 136 -584
rect 362 -585 363 -577
rect 380 -612 381 -584
rect 387 -585 388 -577
rect 436 -612 437 -584
rect 509 -612 510 -584
rect 523 -612 524 -584
rect 534 -612 535 -584
rect 30 -587 31 -577
rect 114 -587 115 -577
rect 138 -612 139 -586
rect 163 -587 164 -577
rect 170 -612 171 -586
rect 187 -587 188 -577
rect 191 -587 192 -577
rect 219 -587 220 -577
rect 236 -587 237 -577
rect 516 -612 517 -586
rect 30 -612 31 -588
rect 51 -589 52 -577
rect 54 -612 55 -588
rect 65 -589 66 -577
rect 72 -612 73 -588
rect 128 -589 129 -577
rect 145 -612 146 -588
rect 156 -589 157 -577
rect 191 -612 192 -588
rect 285 -589 286 -577
rect 352 -612 353 -588
rect 548 -612 549 -588
rect 16 -612 17 -590
rect 51 -612 52 -590
rect 58 -612 59 -590
rect 65 -612 66 -590
rect 79 -591 80 -577
rect 117 -591 118 -577
rect 142 -591 143 -577
rect 156 -612 157 -590
rect 198 -591 199 -577
rect 229 -591 230 -577
rect 240 -612 241 -590
rect 394 -612 395 -590
rect 443 -591 444 -577
rect 464 -612 465 -590
rect 471 -591 472 -577
rect 527 -612 528 -590
rect 37 -612 38 -592
rect 44 -593 45 -577
rect 79 -612 80 -592
rect 107 -612 108 -592
rect 149 -593 150 -577
rect 173 -593 174 -577
rect 198 -612 199 -592
rect 271 -593 272 -577
rect 275 -612 276 -592
rect 317 -593 318 -577
rect 387 -612 388 -592
rect 422 -593 423 -577
rect 443 -612 444 -592
rect 457 -593 458 -577
rect 481 -612 482 -592
rect 506 -593 507 -577
rect 103 -612 104 -594
rect 163 -612 164 -594
rect 205 -595 206 -577
rect 296 -595 297 -577
rect 373 -595 374 -577
rect 457 -612 458 -594
rect 485 -595 486 -577
rect 513 -595 514 -577
rect 142 -612 143 -596
rect 373 -612 374 -596
rect 401 -597 402 -577
rect 471 -612 472 -596
rect 485 -612 486 -596
rect 492 -597 493 -577
rect 499 -612 500 -596
rect 513 -612 514 -596
rect 149 -612 150 -598
rect 310 -612 311 -598
rect 450 -612 451 -598
rect 478 -599 479 -577
rect 205 -612 206 -600
rect 327 -612 328 -600
rect 208 -603 209 -577
rect 233 -612 234 -602
rect 247 -612 248 -602
rect 261 -603 262 -577
rect 268 -603 269 -577
rect 492 -612 493 -602
rect 177 -605 178 -577
rect 268 -612 269 -604
rect 289 -612 290 -604
rect 422 -612 423 -604
rect 219 -612 220 -606
rect 299 -612 300 -606
rect 306 -607 307 -577
rect 401 -612 402 -606
rect 229 -612 230 -608
rect 317 -612 318 -608
rect 261 -612 262 -610
rect 313 -611 314 -577
rect 9 -622 10 -620
rect 68 -622 69 -620
rect 72 -622 73 -620
rect 131 -622 132 -620
rect 142 -622 143 -620
rect 226 -622 227 -620
rect 233 -622 234 -620
rect 292 -622 293 -620
rect 296 -622 297 -620
rect 380 -622 381 -620
rect 394 -622 395 -620
rect 436 -622 437 -620
rect 443 -622 444 -620
rect 474 -659 475 -621
rect 499 -622 500 -620
rect 506 -659 507 -621
rect 513 -659 514 -621
rect 583 -659 584 -621
rect 16 -624 17 -620
rect 61 -659 62 -623
rect 65 -659 66 -623
rect 117 -659 118 -623
rect 121 -624 122 -620
rect 121 -659 122 -623
rect 121 -624 122 -620
rect 121 -659 122 -623
rect 163 -624 164 -620
rect 177 -624 178 -620
rect 184 -659 185 -623
rect 198 -624 199 -620
rect 219 -624 220 -620
rect 247 -624 248 -620
rect 261 -624 262 -620
rect 418 -624 419 -620
rect 422 -624 423 -620
rect 436 -659 437 -623
rect 450 -624 451 -620
rect 488 -659 489 -623
rect 516 -624 517 -620
rect 534 -624 535 -620
rect 544 -659 545 -623
rect 555 -624 556 -620
rect 23 -626 24 -620
rect 89 -626 90 -620
rect 93 -626 94 -620
rect 100 -659 101 -625
rect 103 -626 104 -620
rect 299 -626 300 -620
rect 310 -626 311 -620
rect 359 -626 360 -620
rect 401 -626 402 -620
rect 443 -659 444 -625
rect 520 -659 521 -625
rect 541 -626 542 -620
rect 555 -659 556 -625
rect 562 -659 563 -625
rect 30 -628 31 -620
rect 47 -628 48 -620
rect 51 -659 52 -627
rect 58 -628 59 -620
rect 72 -659 73 -627
rect 79 -659 80 -627
rect 96 -659 97 -627
rect 208 -659 209 -627
rect 222 -628 223 -620
rect 261 -659 262 -627
rect 275 -628 276 -620
rect 310 -659 311 -627
rect 317 -628 318 -620
rect 450 -659 451 -627
rect 527 -628 528 -620
rect 534 -659 535 -627
rect 37 -630 38 -620
rect 44 -630 45 -620
rect 107 -630 108 -620
rect 135 -659 136 -629
rect 149 -630 150 -620
rect 177 -659 178 -629
rect 226 -659 227 -629
rect 303 -630 304 -620
rect 327 -630 328 -620
rect 429 -630 430 -620
rect 44 -659 45 -631
rect 320 -659 321 -631
rect 334 -659 335 -631
rect 387 -632 388 -620
rect 397 -632 398 -620
rect 429 -659 430 -631
rect 86 -634 87 -620
rect 107 -659 108 -633
rect 114 -634 115 -620
rect 219 -659 220 -633
rect 233 -659 234 -633
rect 250 -659 251 -633
rect 275 -659 276 -633
rect 348 -659 349 -633
rect 352 -634 353 -620
rect 457 -634 458 -620
rect 75 -659 76 -635
rect 86 -659 87 -635
rect 114 -659 115 -635
rect 247 -659 248 -635
rect 282 -636 283 -620
rect 282 -659 283 -635
rect 282 -636 283 -620
rect 282 -659 283 -635
rect 296 -659 297 -635
rect 373 -636 374 -620
rect 380 -659 381 -635
rect 397 -659 398 -635
rect 408 -636 409 -620
rect 415 -659 416 -635
rect 422 -659 423 -635
rect 471 -636 472 -620
rect 131 -659 132 -637
rect 359 -659 360 -637
rect 366 -638 367 -620
rect 471 -659 472 -637
rect 149 -659 150 -639
rect 156 -640 157 -620
rect 163 -659 164 -639
rect 212 -640 213 -620
rect 240 -640 241 -620
rect 289 -640 290 -620
rect 324 -640 325 -620
rect 457 -659 458 -639
rect 128 -659 129 -641
rect 156 -659 157 -641
rect 170 -642 171 -620
rect 187 -642 188 -620
rect 191 -642 192 -620
rect 303 -659 304 -641
rect 324 -659 325 -641
rect 530 -659 531 -641
rect 40 -659 41 -643
rect 170 -659 171 -643
rect 180 -644 181 -620
rect 191 -659 192 -643
rect 205 -644 206 -620
rect 212 -659 213 -643
rect 254 -644 255 -620
rect 289 -659 290 -643
rect 331 -644 332 -620
rect 366 -659 367 -643
rect 401 -659 402 -643
rect 408 -659 409 -643
rect 254 -659 255 -645
rect 548 -646 549 -620
rect 331 -659 332 -647
rect 387 -659 388 -647
rect 481 -648 482 -620
rect 548 -659 549 -647
rect 338 -659 339 -649
rect 478 -659 479 -649
rect 341 -652 342 -620
rect 499 -659 500 -651
rect 268 -654 269 -620
rect 341 -659 342 -653
rect 345 -654 346 -620
rect 352 -659 353 -653
rect 355 -654 356 -620
rect 492 -654 493 -620
rect 345 -659 346 -655
rect 464 -656 465 -620
rect 485 -656 486 -620
rect 492 -659 493 -655
rect 464 -659 465 -657
rect 516 -659 517 -657
rect 16 -708 17 -668
rect 65 -669 66 -667
rect 107 -669 108 -667
rect 110 -708 111 -668
rect 114 -669 115 -667
rect 135 -669 136 -667
rect 142 -669 143 -667
rect 142 -708 143 -668
rect 142 -669 143 -667
rect 142 -708 143 -668
rect 156 -669 157 -667
rect 271 -669 272 -667
rect 296 -669 297 -667
rect 317 -708 318 -668
rect 320 -669 321 -667
rect 429 -669 430 -667
rect 471 -669 472 -667
rect 618 -708 619 -668
rect 628 -708 629 -668
rect 639 -708 640 -668
rect 23 -708 24 -670
rect 103 -671 104 -667
rect 156 -708 157 -670
rect 177 -671 178 -667
rect 205 -671 206 -667
rect 212 -671 213 -667
rect 240 -708 241 -670
rect 289 -671 290 -667
rect 303 -671 304 -667
rect 404 -671 405 -667
rect 471 -708 472 -670
rect 478 -671 479 -667
rect 485 -708 486 -670
rect 488 -671 489 -667
rect 499 -671 500 -667
rect 513 -708 514 -670
rect 516 -671 517 -667
rect 520 -671 521 -667
rect 527 -708 528 -670
rect 611 -708 612 -670
rect 30 -708 31 -672
rect 37 -708 38 -672
rect 44 -673 45 -667
rect 100 -673 101 -667
rect 163 -673 164 -667
rect 166 -708 167 -672
rect 170 -673 171 -667
rect 233 -673 234 -667
rect 247 -673 248 -667
rect 303 -708 304 -672
rect 345 -673 346 -667
rect 576 -708 577 -672
rect 583 -673 584 -667
rect 646 -708 647 -672
rect 44 -708 45 -674
rect 51 -675 52 -667
rect 58 -675 59 -667
rect 79 -675 80 -667
rect 93 -708 94 -674
rect 103 -708 104 -674
rect 114 -708 115 -674
rect 163 -708 164 -674
rect 170 -708 171 -674
rect 226 -675 227 -667
rect 247 -708 248 -674
rect 299 -708 300 -674
rect 348 -675 349 -667
rect 366 -675 367 -667
rect 376 -675 377 -667
rect 415 -675 416 -667
rect 478 -708 479 -674
rect 492 -675 493 -667
rect 499 -708 500 -674
rect 555 -675 556 -667
rect 593 -708 594 -674
rect 632 -708 633 -674
rect 51 -708 52 -676
rect 334 -708 335 -676
rect 352 -708 353 -676
rect 373 -677 374 -667
rect 380 -677 381 -667
rect 401 -677 402 -667
rect 415 -708 416 -676
rect 457 -677 458 -667
rect 506 -677 507 -667
rect 520 -708 521 -676
rect 530 -677 531 -667
rect 534 -677 535 -667
rect 548 -677 549 -667
rect 562 -708 563 -676
rect 65 -708 66 -678
rect 86 -679 87 -667
rect 191 -679 192 -667
rect 226 -708 227 -678
rect 250 -679 251 -667
rect 464 -679 465 -667
rect 72 -708 73 -680
rect 79 -708 80 -680
rect 86 -708 87 -680
rect 121 -681 122 -667
rect 201 -681 202 -667
rect 205 -708 206 -680
rect 212 -708 213 -680
rect 275 -681 276 -667
rect 296 -708 297 -680
rect 555 -708 556 -680
rect 121 -708 122 -682
rect 198 -708 199 -682
rect 219 -683 220 -667
rect 275 -708 276 -682
rect 324 -683 325 -667
rect 373 -708 374 -682
rect 380 -708 381 -682
rect 604 -708 605 -682
rect 177 -708 178 -684
rect 201 -708 202 -684
rect 219 -708 220 -684
rect 243 -685 244 -667
rect 254 -685 255 -667
rect 324 -708 325 -684
rect 331 -708 332 -684
rect 534 -708 535 -684
rect 184 -687 185 -667
rect 254 -708 255 -686
rect 261 -687 262 -667
rect 289 -708 290 -686
rect 338 -687 339 -667
rect 506 -708 507 -686
rect 135 -708 136 -688
rect 261 -708 262 -688
rect 268 -689 269 -667
rect 548 -708 549 -688
rect 149 -691 150 -667
rect 184 -708 185 -690
rect 194 -708 195 -690
rect 268 -708 269 -690
rect 310 -691 311 -667
rect 338 -708 339 -690
rect 359 -691 360 -667
rect 401 -708 402 -690
rect 443 -691 444 -667
rect 457 -708 458 -690
rect 128 -708 129 -692
rect 149 -708 150 -692
rect 233 -708 234 -692
rect 310 -708 311 -692
rect 366 -708 367 -692
rect 408 -693 409 -667
rect 443 -708 444 -692
rect 544 -693 545 -667
rect 282 -695 283 -667
rect 359 -708 360 -694
rect 387 -695 388 -667
rect 583 -708 584 -694
rect 387 -708 388 -696
rect 436 -697 437 -667
rect 450 -697 451 -667
rect 464 -708 465 -696
rect 345 -708 346 -698
rect 436 -708 437 -698
rect 450 -708 451 -698
rect 572 -708 573 -698
rect 394 -701 395 -667
rect 429 -708 430 -700
rect 397 -703 398 -667
rect 422 -703 423 -667
rect 408 -708 409 -704
rect 474 -705 475 -667
rect 422 -708 423 -706
rect 541 -708 542 -706
rect 16 -718 17 -716
rect 58 -718 59 -716
rect 86 -718 87 -716
rect 135 -759 136 -717
rect 142 -718 143 -716
rect 149 -718 150 -716
rect 152 -718 153 -716
rect 187 -718 188 -716
rect 194 -718 195 -716
rect 205 -718 206 -716
rect 219 -718 220 -716
rect 254 -718 255 -716
rect 261 -718 262 -716
rect 345 -718 346 -716
rect 348 -718 349 -716
rect 415 -718 416 -716
rect 422 -759 423 -717
rect 488 -759 489 -717
rect 495 -718 496 -716
rect 534 -718 535 -716
rect 541 -718 542 -716
rect 614 -718 615 -716
rect 23 -720 24 -716
rect 65 -720 66 -716
rect 79 -720 80 -716
rect 149 -759 150 -719
rect 156 -720 157 -716
rect 261 -759 262 -719
rect 268 -720 269 -716
rect 331 -720 332 -716
rect 334 -720 335 -716
rect 471 -720 472 -716
rect 474 -759 475 -719
rect 534 -759 535 -719
rect 562 -720 563 -716
rect 600 -720 601 -716
rect 611 -759 612 -719
rect 632 -720 633 -716
rect 33 -759 34 -721
rect 37 -722 38 -716
rect 44 -722 45 -716
rect 75 -722 76 -716
rect 79 -759 80 -721
rect 114 -722 115 -716
rect 156 -759 157 -721
rect 285 -759 286 -721
rect 296 -722 297 -716
rect 324 -722 325 -716
rect 338 -722 339 -716
rect 464 -722 465 -716
rect 485 -722 486 -716
rect 485 -759 486 -721
rect 485 -722 486 -716
rect 485 -759 486 -721
rect 499 -722 500 -716
rect 572 -722 573 -716
rect 593 -722 594 -716
rect 646 -722 647 -716
rect 44 -759 45 -723
rect 121 -724 122 -716
rect 163 -724 164 -716
rect 177 -724 178 -716
rect 194 -759 195 -723
rect 303 -724 304 -716
rect 310 -724 311 -716
rect 506 -724 507 -716
rect 527 -724 528 -716
rect 530 -759 531 -723
rect 569 -724 570 -716
rect 604 -724 605 -716
rect 51 -726 52 -716
rect 257 -759 258 -725
rect 268 -759 269 -725
rect 289 -726 290 -716
rect 310 -759 311 -725
rect 359 -726 360 -716
rect 366 -726 367 -716
rect 527 -759 528 -725
rect 597 -726 598 -716
rect 639 -726 640 -716
rect 51 -759 52 -727
rect 128 -728 129 -716
rect 163 -759 164 -727
rect 229 -759 230 -727
rect 233 -728 234 -716
rect 233 -759 234 -727
rect 233 -728 234 -716
rect 233 -759 234 -727
rect 240 -728 241 -716
rect 303 -759 304 -727
rect 317 -728 318 -716
rect 324 -759 325 -727
rect 352 -728 353 -716
rect 541 -759 542 -727
rect 65 -759 66 -729
rect 72 -730 73 -716
rect 86 -759 87 -729
rect 93 -730 94 -716
rect 103 -730 104 -716
rect 457 -730 458 -716
rect 464 -759 465 -729
rect 555 -730 556 -716
rect 58 -759 59 -731
rect 103 -759 104 -731
rect 114 -759 115 -731
rect 128 -759 129 -731
rect 170 -732 171 -716
rect 201 -732 202 -716
rect 205 -759 206 -731
rect 296 -759 297 -731
rect 317 -759 318 -731
rect 331 -759 332 -731
rect 352 -759 353 -731
rect 359 -759 360 -731
rect 366 -759 367 -731
rect 513 -732 514 -716
rect 555 -759 556 -731
rect 618 -732 619 -716
rect 72 -759 73 -733
rect 107 -734 108 -716
rect 121 -759 122 -733
rect 215 -759 216 -733
rect 226 -734 227 -716
rect 240 -759 241 -733
rect 247 -734 248 -716
rect 383 -734 384 -716
rect 397 -734 398 -716
rect 520 -734 521 -716
rect 93 -759 94 -735
rect 152 -759 153 -735
rect 170 -759 171 -735
rect 212 -736 213 -716
rect 250 -759 251 -735
rect 387 -736 388 -716
rect 408 -736 409 -716
rect 520 -759 521 -735
rect 107 -759 108 -737
rect 198 -738 199 -716
rect 222 -738 223 -716
rect 387 -759 388 -737
rect 408 -759 409 -737
rect 443 -738 444 -716
rect 450 -738 451 -716
rect 457 -759 458 -737
rect 506 -759 507 -737
rect 576 -738 577 -716
rect 177 -759 178 -739
rect 191 -740 192 -716
rect 222 -759 223 -739
rect 362 -759 363 -739
rect 373 -740 374 -716
rect 492 -759 493 -739
rect 184 -742 185 -716
rect 198 -759 199 -741
rect 254 -759 255 -741
rect 348 -759 349 -741
rect 380 -742 381 -716
rect 478 -742 479 -716
rect 142 -759 143 -743
rect 184 -759 185 -743
rect 275 -744 276 -716
rect 278 -759 279 -743
rect 282 -744 283 -716
rect 401 -744 402 -716
rect 415 -759 416 -743
rect 471 -759 472 -743
rect 478 -759 479 -743
rect 548 -744 549 -716
rect 292 -759 293 -745
rect 401 -759 402 -745
rect 425 -746 426 -716
rect 583 -746 584 -716
rect 334 -759 335 -747
rect 513 -759 514 -747
rect 338 -759 339 -749
rect 450 -759 451 -749
rect 380 -759 381 -751
rect 436 -752 437 -716
rect 429 -754 430 -716
rect 499 -759 500 -753
rect 394 -756 395 -716
rect 429 -759 430 -755
rect 394 -759 395 -757
rect 436 -759 437 -757
rect 26 -816 27 -768
rect 33 -769 34 -767
rect 40 -769 41 -767
rect 149 -769 150 -767
rect 152 -769 153 -767
rect 373 -769 374 -767
rect 387 -769 388 -767
rect 394 -816 395 -768
rect 397 -769 398 -767
rect 457 -769 458 -767
rect 471 -769 472 -767
rect 520 -769 521 -767
rect 534 -769 535 -767
rect 558 -816 559 -768
rect 30 -816 31 -770
rect 37 -816 38 -770
rect 44 -771 45 -767
rect 114 -816 115 -770
rect 128 -771 129 -767
rect 166 -816 167 -770
rect 170 -771 171 -767
rect 191 -771 192 -767
rect 212 -771 213 -767
rect 268 -771 269 -767
rect 275 -771 276 -767
rect 436 -771 437 -767
rect 446 -771 447 -767
rect 478 -771 479 -767
rect 492 -771 493 -767
rect 527 -816 528 -770
rect 44 -816 45 -772
rect 93 -773 94 -767
rect 128 -816 129 -772
rect 187 -816 188 -772
rect 212 -816 213 -772
rect 310 -773 311 -767
rect 324 -773 325 -767
rect 338 -773 339 -767
rect 352 -773 353 -767
rect 460 -816 461 -772
rect 513 -773 514 -767
rect 548 -816 549 -772
rect 51 -775 52 -767
rect 145 -775 146 -767
rect 156 -775 157 -767
rect 194 -775 195 -767
rect 219 -775 220 -767
rect 261 -775 262 -767
rect 285 -775 286 -767
rect 317 -775 318 -767
rect 334 -816 335 -774
rect 485 -816 486 -774
rect 499 -775 500 -767
rect 513 -816 514 -774
rect 520 -816 521 -774
rect 555 -775 556 -767
rect 51 -816 52 -776
rect 121 -777 122 -767
rect 135 -777 136 -767
rect 135 -816 136 -776
rect 135 -777 136 -767
rect 135 -816 136 -776
rect 156 -816 157 -776
rect 191 -816 192 -776
rect 222 -777 223 -767
rect 289 -816 290 -776
rect 292 -777 293 -767
rect 376 -777 377 -767
rect 401 -777 402 -767
rect 499 -816 500 -776
rect 58 -779 59 -767
rect 142 -816 143 -778
rect 163 -779 164 -767
rect 331 -779 332 -767
rect 338 -816 339 -778
rect 443 -779 444 -767
rect 492 -816 493 -778
rect 555 -816 556 -778
rect 58 -816 59 -780
rect 65 -781 66 -767
rect 72 -781 73 -767
rect 152 -816 153 -780
rect 163 -816 164 -780
rect 282 -816 283 -780
rect 303 -781 304 -767
rect 387 -816 388 -780
rect 429 -781 430 -767
rect 534 -816 535 -780
rect 65 -816 66 -782
rect 331 -816 332 -782
rect 359 -783 360 -767
rect 464 -783 465 -767
rect 72 -816 73 -784
rect 145 -816 146 -784
rect 170 -816 171 -784
rect 257 -785 258 -767
rect 261 -816 262 -784
rect 422 -785 423 -767
rect 443 -816 444 -784
rect 530 -785 531 -767
rect 86 -787 87 -767
rect 117 -787 118 -767
rect 121 -816 122 -786
rect 436 -816 437 -786
rect 464 -816 465 -786
rect 506 -787 507 -767
rect 86 -816 87 -788
rect 205 -789 206 -767
rect 226 -789 227 -767
rect 275 -816 276 -788
rect 303 -816 304 -788
rect 352 -816 353 -788
rect 359 -816 360 -788
rect 380 -789 381 -767
rect 404 -816 405 -788
rect 429 -816 430 -788
rect 93 -816 94 -790
rect 257 -816 258 -790
rect 306 -791 307 -767
rect 478 -816 479 -790
rect 177 -793 178 -767
rect 324 -816 325 -792
rect 103 -816 104 -794
rect 177 -816 178 -794
rect 184 -795 185 -767
rect 226 -816 227 -794
rect 229 -795 230 -767
rect 366 -795 367 -767
rect 205 -816 206 -796
rect 215 -797 216 -767
rect 233 -797 234 -767
rect 268 -816 269 -796
rect 313 -816 314 -796
rect 506 -816 507 -796
rect 215 -816 216 -798
rect 219 -816 220 -798
rect 236 -816 237 -798
rect 341 -799 342 -767
rect 366 -816 367 -798
rect 408 -799 409 -767
rect 240 -801 241 -767
rect 240 -816 241 -800
rect 240 -801 241 -767
rect 240 -816 241 -800
rect 247 -801 248 -767
rect 296 -801 297 -767
rect 317 -816 318 -800
rect 471 -816 472 -800
rect 247 -816 248 -802
rect 422 -816 423 -802
rect 254 -816 255 -804
rect 541 -805 542 -767
rect 296 -816 297 -806
rect 380 -816 381 -806
rect 450 -807 451 -767
rect 541 -816 542 -806
rect 376 -816 377 -808
rect 408 -816 409 -808
rect 415 -809 416 -767
rect 450 -816 451 -808
rect 107 -811 108 -767
rect 415 -816 416 -810
rect 79 -813 80 -767
rect 107 -816 108 -812
rect 79 -816 80 -814
rect 198 -815 199 -767
rect 26 -879 27 -825
rect 40 -879 41 -825
rect 44 -826 45 -824
rect 236 -826 237 -824
rect 240 -826 241 -824
rect 247 -826 248 -824
rect 254 -879 255 -825
rect 285 -879 286 -825
rect 306 -879 307 -825
rect 485 -826 486 -824
rect 30 -879 31 -827
rect 37 -828 38 -824
rect 44 -879 45 -827
rect 72 -879 73 -827
rect 75 -879 76 -827
rect 110 -828 111 -824
rect 114 -879 115 -827
rect 142 -879 143 -827
rect 145 -828 146 -824
rect 317 -828 318 -824
rect 320 -828 321 -824
rect 387 -828 388 -824
rect 401 -828 402 -824
rect 464 -828 465 -824
rect 467 -879 468 -827
rect 541 -828 542 -824
rect 51 -830 52 -824
rect 159 -830 160 -824
rect 173 -879 174 -829
rect 194 -879 195 -829
rect 201 -830 202 -824
rect 404 -830 405 -824
rect 450 -830 451 -824
rect 485 -879 486 -829
rect 37 -879 38 -831
rect 51 -879 52 -831
rect 58 -879 59 -831
rect 180 -879 181 -831
rect 187 -832 188 -824
rect 310 -832 311 -824
rect 313 -832 314 -824
rect 548 -832 549 -824
rect 79 -834 80 -824
rect 163 -834 164 -824
rect 212 -879 213 -833
rect 219 -834 220 -824
rect 240 -879 241 -833
rect 275 -834 276 -824
rect 296 -834 297 -824
rect 450 -879 451 -833
rect 457 -879 458 -833
rect 464 -879 465 -833
rect 79 -879 80 -835
rect 170 -836 171 -824
rect 177 -836 178 -824
rect 219 -879 220 -835
rect 261 -836 262 -824
rect 324 -836 325 -824
rect 331 -879 332 -835
rect 366 -836 367 -824
rect 373 -836 374 -824
rect 513 -836 514 -824
rect 86 -838 87 -824
rect 201 -879 202 -837
rect 205 -838 206 -824
rect 261 -879 262 -837
rect 310 -879 311 -837
rect 317 -879 318 -837
rect 324 -879 325 -837
rect 359 -838 360 -824
rect 366 -879 367 -837
rect 429 -838 430 -824
rect 86 -879 87 -839
rect 135 -840 136 -824
rect 149 -840 150 -824
rect 558 -840 559 -824
rect 100 -879 101 -841
rect 226 -842 227 -824
rect 257 -842 258 -824
rect 513 -879 514 -841
rect 107 -879 108 -843
rect 191 -844 192 -824
rect 226 -879 227 -843
rect 282 -844 283 -824
rect 313 -879 314 -843
rect 471 -844 472 -824
rect 117 -879 118 -845
rect 429 -879 430 -845
rect 121 -879 122 -847
rect 303 -848 304 -824
rect 348 -848 349 -824
rect 499 -848 500 -824
rect 124 -850 125 -824
rect 128 -850 129 -824
rect 149 -879 150 -849
rect 334 -879 335 -849
rect 338 -850 339 -824
rect 499 -879 500 -849
rect 93 -852 94 -824
rect 128 -879 129 -851
rect 156 -879 157 -851
rect 275 -879 276 -851
rect 289 -852 290 -824
rect 338 -879 339 -851
rect 355 -852 356 -824
rect 534 -852 535 -824
rect 65 -854 66 -824
rect 93 -879 94 -853
rect 163 -879 164 -853
rect 184 -879 185 -853
rect 247 -879 248 -853
rect 355 -879 356 -853
rect 359 -879 360 -853
rect 408 -854 409 -824
rect 520 -854 521 -824
rect 534 -879 535 -853
rect 65 -879 66 -855
rect 198 -856 199 -824
rect 268 -856 269 -824
rect 289 -879 290 -855
rect 373 -879 374 -855
rect 506 -856 507 -824
rect 268 -879 269 -857
rect 380 -858 381 -824
rect 387 -879 388 -857
rect 474 -879 475 -857
rect 492 -858 493 -824
rect 506 -879 507 -857
rect 376 -860 377 -824
rect 527 -860 528 -824
rect 348 -879 349 -861
rect 527 -879 528 -861
rect 401 -879 402 -863
rect 436 -864 437 -824
rect 408 -879 409 -865
rect 422 -866 423 -824
rect 436 -879 437 -865
rect 478 -866 479 -824
rect 352 -879 353 -867
rect 478 -879 479 -867
rect 415 -870 416 -824
rect 492 -879 493 -869
rect 394 -872 395 -824
rect 415 -879 416 -871
rect 422 -879 423 -871
rect 443 -872 444 -824
rect 152 -874 153 -824
rect 443 -879 444 -873
rect 233 -876 234 -824
rect 394 -879 395 -875
rect 233 -879 234 -877
rect 296 -879 297 -877
rect 9 -934 10 -888
rect 135 -934 136 -888
rect 142 -889 143 -887
rect 156 -889 157 -887
rect 159 -889 160 -887
rect 492 -889 493 -887
rect 520 -889 521 -887
rect 534 -889 535 -887
rect 16 -934 17 -890
rect 208 -891 209 -887
rect 240 -891 241 -887
rect 264 -934 265 -890
rect 268 -891 269 -887
rect 334 -891 335 -887
rect 348 -891 349 -887
rect 485 -891 486 -887
rect 520 -934 521 -890
rect 523 -891 524 -887
rect 23 -934 24 -892
rect 44 -893 45 -887
rect 58 -893 59 -887
rect 345 -893 346 -887
rect 355 -893 356 -887
rect 436 -893 437 -887
rect 457 -893 458 -887
rect 492 -934 493 -892
rect 44 -934 45 -894
rect 51 -895 52 -887
rect 58 -934 59 -894
rect 72 -934 73 -894
rect 79 -895 80 -887
rect 170 -895 171 -887
rect 177 -934 178 -894
rect 212 -895 213 -887
rect 240 -934 241 -894
rect 334 -934 335 -894
rect 359 -895 360 -887
rect 362 -921 363 -894
rect 373 -895 374 -887
rect 373 -934 374 -894
rect 373 -895 374 -887
rect 373 -934 374 -894
rect 380 -895 381 -887
rect 513 -895 514 -887
rect 37 -934 38 -896
rect 212 -934 213 -896
rect 233 -897 234 -887
rect 380 -934 381 -896
rect 383 -897 384 -887
rect 513 -934 514 -896
rect 51 -934 52 -898
rect 285 -899 286 -887
rect 313 -899 314 -887
rect 408 -899 409 -887
rect 422 -899 423 -887
rect 474 -899 475 -887
rect 478 -899 479 -887
rect 485 -934 486 -898
rect 65 -901 66 -887
rect 138 -901 139 -887
rect 142 -934 143 -900
rect 254 -901 255 -887
rect 282 -901 283 -887
rect 324 -901 325 -887
rect 331 -934 332 -900
rect 499 -901 500 -887
rect 65 -934 66 -902
rect 191 -903 192 -887
rect 194 -903 195 -887
rect 261 -903 262 -887
rect 282 -934 283 -902
rect 324 -934 325 -902
rect 352 -903 353 -887
rect 499 -934 500 -902
rect 86 -905 87 -887
rect 229 -934 230 -904
rect 296 -905 297 -887
rect 422 -934 423 -904
rect 436 -934 437 -904
rect 443 -905 444 -887
rect 478 -934 479 -904
rect 506 -905 507 -887
rect 93 -907 94 -887
rect 163 -907 164 -887
rect 201 -907 202 -887
rect 292 -934 293 -906
rect 317 -907 318 -887
rect 345 -934 346 -906
rect 359 -934 360 -906
rect 401 -907 402 -887
rect 506 -934 507 -906
rect 527 -907 528 -887
rect 93 -934 94 -908
rect 128 -909 129 -887
rect 149 -909 150 -887
rect 268 -934 269 -908
rect 317 -934 318 -908
rect 338 -909 339 -887
rect 394 -909 395 -887
rect 408 -934 409 -908
rect 100 -911 101 -887
rect 180 -911 181 -887
rect 205 -911 206 -887
rect 289 -911 290 -887
rect 397 -934 398 -910
rect 471 -934 472 -910
rect 107 -913 108 -887
rect 306 -913 307 -887
rect 401 -934 402 -912
rect 415 -913 416 -887
rect 107 -934 108 -914
rect 247 -915 248 -887
rect 275 -915 276 -887
rect 338 -934 339 -914
rect 415 -934 416 -914
rect 429 -915 430 -887
rect 114 -934 115 -916
rect 149 -934 150 -916
rect 152 -934 153 -916
rect 170 -934 171 -916
rect 201 -934 202 -916
rect 247 -934 248 -916
rect 306 -934 307 -916
rect 366 -917 367 -887
rect 429 -934 430 -916
rect 450 -917 451 -887
rect 121 -934 122 -918
rect 184 -919 185 -887
rect 208 -934 209 -918
rect 296 -934 297 -918
rect 387 -919 388 -887
rect 450 -934 451 -918
rect 124 -921 125 -887
rect 166 -921 167 -887
rect 184 -934 185 -920
rect 222 -934 223 -920
rect 226 -921 227 -887
rect 233 -934 234 -920
rect 387 -934 388 -920
rect 128 -934 129 -922
rect 194 -934 195 -922
rect 219 -923 220 -887
rect 275 -934 276 -922
rect 159 -934 160 -924
rect 310 -925 311 -887
rect 166 -934 167 -926
rect 254 -934 255 -926
rect 205 -934 206 -928
rect 310 -934 311 -928
rect 219 -934 220 -930
rect 366 -934 367 -930
rect 226 -934 227 -932
rect 457 -934 458 -932
rect 2 -983 3 -943
rect 163 -944 164 -942
rect 201 -944 202 -942
rect 422 -944 423 -942
rect 443 -944 444 -942
rect 499 -944 500 -942
rect 16 -946 17 -942
rect 103 -946 104 -942
rect 107 -946 108 -942
rect 110 -966 111 -945
rect 114 -946 115 -942
rect 138 -983 139 -945
rect 142 -946 143 -942
rect 191 -946 192 -942
rect 212 -946 213 -942
rect 240 -946 241 -942
rect 257 -983 258 -945
rect 296 -946 297 -942
rect 299 -983 300 -945
rect 415 -946 416 -942
rect 429 -946 430 -942
rect 443 -983 444 -945
rect 464 -946 465 -942
rect 485 -946 486 -942
rect 9 -948 10 -942
rect 191 -983 192 -947
rect 222 -983 223 -947
rect 261 -983 262 -947
rect 268 -948 269 -942
rect 303 -983 304 -947
rect 310 -948 311 -942
rect 408 -983 409 -947
rect 467 -983 468 -947
rect 492 -948 493 -942
rect 23 -950 24 -942
rect 30 -950 31 -942
rect 37 -950 38 -942
rect 198 -950 199 -942
rect 254 -950 255 -942
rect 310 -983 311 -949
rect 317 -950 318 -942
rect 317 -983 318 -949
rect 317 -950 318 -942
rect 317 -983 318 -949
rect 324 -950 325 -942
rect 401 -950 402 -942
rect 492 -983 493 -949
rect 513 -950 514 -942
rect 9 -983 10 -951
rect 30 -983 31 -951
rect 44 -983 45 -951
rect 184 -952 185 -942
rect 187 -983 188 -951
rect 212 -983 213 -951
rect 268 -983 269 -951
rect 275 -952 276 -942
rect 296 -983 297 -951
rect 324 -983 325 -951
rect 327 -952 328 -942
rect 415 -983 416 -951
rect 16 -983 17 -953
rect 23 -983 24 -953
rect 51 -954 52 -942
rect 166 -954 167 -942
rect 198 -983 199 -953
rect 429 -983 430 -953
rect 51 -983 52 -955
rect 58 -956 59 -942
rect 65 -956 66 -942
rect 201 -983 202 -955
rect 247 -956 248 -942
rect 275 -983 276 -955
rect 338 -956 339 -942
rect 380 -983 381 -955
rect 394 -956 395 -942
rect 478 -956 479 -942
rect 65 -983 66 -957
rect 205 -958 206 -942
rect 306 -958 307 -942
rect 394 -983 395 -957
rect 478 -983 479 -957
rect 506 -958 507 -942
rect 75 -983 76 -959
rect 100 -960 101 -942
rect 107 -983 108 -959
rect 170 -960 171 -942
rect 177 -960 178 -942
rect 205 -983 206 -959
rect 331 -983 332 -959
rect 338 -983 339 -959
rect 345 -960 346 -942
rect 401 -983 402 -959
rect 506 -983 507 -959
rect 520 -960 521 -942
rect 86 -962 87 -942
rect 156 -962 157 -942
rect 163 -983 164 -961
rect 282 -962 283 -942
rect 289 -962 290 -942
rect 345 -983 346 -961
rect 352 -962 353 -942
rect 450 -962 451 -942
rect 86 -983 87 -963
rect 292 -983 293 -963
rect 373 -964 374 -942
rect 422 -983 423 -963
rect 93 -966 94 -942
rect 103 -983 104 -965
rect 170 -983 171 -965
rect 177 -983 178 -965
rect 264 -966 265 -942
rect 373 -983 374 -965
rect 387 -966 388 -942
rect 96 -983 97 -967
rect 471 -968 472 -942
rect 114 -983 115 -969
rect 166 -983 167 -969
rect 194 -983 195 -969
rect 247 -983 248 -969
rect 264 -983 265 -969
rect 436 -970 437 -942
rect 457 -970 458 -942
rect 471 -983 472 -969
rect 121 -972 122 -942
rect 219 -972 220 -942
rect 226 -972 227 -942
rect 457 -983 458 -971
rect 128 -974 129 -942
rect 184 -983 185 -973
rect 233 -974 234 -942
rect 282 -983 283 -973
rect 359 -974 360 -942
rect 387 -983 388 -973
rect 82 -976 83 -942
rect 233 -983 234 -975
rect 355 -983 356 -975
rect 359 -983 360 -975
rect 366 -976 367 -942
rect 436 -983 437 -975
rect 135 -983 136 -977
rect 142 -983 143 -977
rect 149 -983 150 -977
rect 229 -978 230 -942
rect 334 -978 335 -942
rect 366 -983 367 -977
rect 159 -980 160 -942
rect 219 -983 220 -979
rect 334 -983 335 -979
rect 450 -983 451 -979
rect 121 -983 122 -981
rect 159 -983 160 -981
rect 9 -993 10 -991
rect 37 -993 38 -991
rect 44 -993 45 -991
rect 219 -993 220 -991
rect 229 -993 230 -991
rect 240 -1030 241 -992
rect 247 -993 248 -991
rect 247 -1030 248 -992
rect 247 -993 248 -991
rect 247 -1030 248 -992
rect 278 -1030 279 -992
rect 380 -993 381 -991
rect 418 -1030 419 -992
rect 436 -993 437 -991
rect 439 -1030 440 -992
rect 478 -993 479 -991
rect 488 -1030 489 -992
rect 506 -993 507 -991
rect 16 -995 17 -991
rect 16 -1030 17 -994
rect 16 -995 17 -991
rect 16 -1030 17 -994
rect 23 -1030 24 -994
rect 33 -995 34 -991
rect 37 -1030 38 -994
rect 47 -1030 48 -994
rect 51 -995 52 -991
rect 58 -995 59 -991
rect 65 -995 66 -991
rect 93 -995 94 -991
rect 107 -995 108 -991
rect 184 -995 185 -991
rect 187 -995 188 -991
rect 275 -995 276 -991
rect 289 -995 290 -991
rect 317 -995 318 -991
rect 341 -995 342 -991
rect 443 -995 444 -991
rect 446 -1030 447 -994
rect 478 -1030 479 -994
rect 40 -997 41 -991
rect 93 -1030 94 -996
rect 107 -1030 108 -996
rect 194 -997 195 -991
rect 205 -997 206 -991
rect 205 -1030 206 -996
rect 205 -997 206 -991
rect 205 -1030 206 -996
rect 215 -1030 216 -996
rect 229 -1030 230 -996
rect 233 -1030 234 -996
rect 345 -997 346 -991
rect 352 -997 353 -991
rect 450 -997 451 -991
rect 467 -1030 468 -996
rect 471 -1030 472 -996
rect 474 -997 475 -991
rect 492 -997 493 -991
rect 58 -1030 59 -998
rect 61 -999 62 -991
rect 79 -999 80 -991
rect 114 -999 115 -991
rect 121 -999 122 -991
rect 121 -1030 122 -998
rect 121 -999 122 -991
rect 121 -1030 122 -998
rect 131 -999 132 -991
rect 324 -999 325 -991
rect 327 -1030 328 -998
rect 345 -1030 346 -998
rect 359 -999 360 -991
rect 359 -1030 360 -998
rect 359 -999 360 -991
rect 359 -1030 360 -998
rect 380 -1030 381 -998
rect 387 -999 388 -991
rect 415 -999 416 -991
rect 450 -1030 451 -998
rect 82 -1001 83 -991
rect 457 -1001 458 -991
rect 2 -1003 3 -991
rect 82 -1030 83 -1002
rect 86 -1003 87 -991
rect 243 -1003 244 -991
rect 285 -1030 286 -1002
rect 289 -1030 290 -1002
rect 303 -1003 304 -991
rect 317 -1030 318 -1002
rect 334 -1030 335 -1002
rect 352 -1030 353 -1002
rect 366 -1003 367 -991
rect 387 -1030 388 -1002
rect 422 -1003 423 -991
rect 464 -1003 465 -991
rect 86 -1030 87 -1004
rect 103 -1005 104 -991
rect 142 -1005 143 -991
rect 142 -1030 143 -1004
rect 142 -1005 143 -991
rect 142 -1030 143 -1004
rect 149 -1005 150 -991
rect 159 -1005 160 -991
rect 163 -1005 164 -991
rect 166 -1030 167 -1004
rect 170 -1005 171 -991
rect 226 -1005 227 -991
rect 310 -1005 311 -991
rect 366 -1030 367 -1004
rect 96 -1007 97 -991
rect 114 -1030 115 -1006
rect 149 -1030 150 -1006
rect 429 -1007 430 -991
rect 156 -1030 157 -1008
rect 170 -1030 171 -1008
rect 191 -1009 192 -991
rect 282 -1009 283 -991
rect 415 -1030 416 -1008
rect 429 -1030 430 -1008
rect 191 -1030 192 -1010
rect 212 -1011 213 -991
rect 222 -1011 223 -991
rect 310 -1030 311 -1010
rect 212 -1030 213 -1012
rect 268 -1013 269 -991
rect 128 -1015 129 -991
rect 268 -1030 269 -1014
rect 128 -1030 129 -1016
rect 177 -1017 178 -991
rect 222 -1030 223 -1016
rect 408 -1017 409 -991
rect 177 -1030 178 -1018
rect 198 -1019 199 -991
rect 394 -1019 395 -991
rect 408 -1030 409 -1018
rect 198 -1030 199 -1020
rect 261 -1021 262 -991
rect 373 -1021 374 -991
rect 394 -1030 395 -1020
rect 254 -1023 255 -991
rect 261 -1030 262 -1022
rect 373 -1030 374 -1022
rect 460 -1030 461 -1022
rect 254 -1030 255 -1024
rect 338 -1025 339 -991
rect 338 -1030 339 -1026
rect 401 -1027 402 -991
rect 292 -1029 293 -991
rect 401 -1030 402 -1028
rect 23 -1040 24 -1038
rect 33 -1040 34 -1038
rect 51 -1075 52 -1039
rect 58 -1040 59 -1038
rect 72 -1075 73 -1039
rect 79 -1040 80 -1038
rect 86 -1040 87 -1038
rect 100 -1040 101 -1038
rect 117 -1075 118 -1039
rect 121 -1040 122 -1038
rect 128 -1040 129 -1038
rect 156 -1040 157 -1038
rect 159 -1075 160 -1039
rect 296 -1075 297 -1039
rect 299 -1040 300 -1038
rect 359 -1040 360 -1038
rect 408 -1040 409 -1038
rect 422 -1040 423 -1038
rect 443 -1040 444 -1038
rect 450 -1040 451 -1038
rect 460 -1040 461 -1038
rect 467 -1040 468 -1038
rect 488 -1040 489 -1038
rect 499 -1075 500 -1039
rect 30 -1075 31 -1041
rect 37 -1042 38 -1038
rect 68 -1075 69 -1041
rect 79 -1075 80 -1041
rect 100 -1075 101 -1041
rect 114 -1042 115 -1038
rect 121 -1075 122 -1041
rect 138 -1042 139 -1038
rect 149 -1042 150 -1038
rect 170 -1042 171 -1038
rect 177 -1042 178 -1038
rect 184 -1042 185 -1038
rect 205 -1042 206 -1038
rect 226 -1042 227 -1038
rect 233 -1042 234 -1038
rect 275 -1075 276 -1041
rect 285 -1042 286 -1038
rect 317 -1042 318 -1038
rect 324 -1042 325 -1038
rect 387 -1042 388 -1038
rect 401 -1042 402 -1038
rect 422 -1075 423 -1041
rect 429 -1042 430 -1038
rect 450 -1075 451 -1041
rect 464 -1075 465 -1041
rect 471 -1042 472 -1038
rect 37 -1075 38 -1043
rect 96 -1044 97 -1038
rect 110 -1075 111 -1043
rect 156 -1075 157 -1043
rect 163 -1075 164 -1043
rect 254 -1044 255 -1038
rect 261 -1044 262 -1038
rect 306 -1075 307 -1043
rect 331 -1075 332 -1043
rect 338 -1044 339 -1038
rect 345 -1044 346 -1038
rect 359 -1075 360 -1043
rect 394 -1044 395 -1038
rect 401 -1075 402 -1043
rect 408 -1075 409 -1043
rect 495 -1075 496 -1043
rect 86 -1075 87 -1045
rect 114 -1075 115 -1045
rect 128 -1075 129 -1045
rect 485 -1046 486 -1038
rect 135 -1048 136 -1038
rect 142 -1048 143 -1038
rect 177 -1075 178 -1047
rect 219 -1048 220 -1038
rect 222 -1075 223 -1047
rect 278 -1048 279 -1038
rect 303 -1048 304 -1038
rect 366 -1048 367 -1038
rect 418 -1048 419 -1038
rect 457 -1048 458 -1038
rect 478 -1048 479 -1038
rect 485 -1075 486 -1047
rect 107 -1050 108 -1038
rect 142 -1075 143 -1049
rect 184 -1075 185 -1049
rect 191 -1050 192 -1038
rect 198 -1050 199 -1038
rect 205 -1075 206 -1049
rect 215 -1075 216 -1049
rect 387 -1075 388 -1049
rect 96 -1075 97 -1051
rect 191 -1075 192 -1051
rect 198 -1075 199 -1051
rect 415 -1075 416 -1051
rect 135 -1075 136 -1053
rect 173 -1075 174 -1053
rect 233 -1075 234 -1053
rect 261 -1075 262 -1053
rect 268 -1054 269 -1038
rect 324 -1075 325 -1053
rect 338 -1075 339 -1053
rect 429 -1075 430 -1053
rect 240 -1056 241 -1038
rect 282 -1075 283 -1055
rect 303 -1075 304 -1055
rect 443 -1075 444 -1055
rect 240 -1075 241 -1057
rect 327 -1058 328 -1038
rect 341 -1075 342 -1057
rect 457 -1075 458 -1057
rect 247 -1060 248 -1038
rect 254 -1075 255 -1059
rect 268 -1075 269 -1059
rect 366 -1075 367 -1059
rect 149 -1075 150 -1061
rect 247 -1075 248 -1061
rect 278 -1075 279 -1061
rect 317 -1075 318 -1061
rect 348 -1075 349 -1061
rect 380 -1062 381 -1038
rect 310 -1064 311 -1038
rect 394 -1075 395 -1063
rect 289 -1066 290 -1038
rect 310 -1075 311 -1065
rect 373 -1066 374 -1038
rect 380 -1075 381 -1065
rect 229 -1068 230 -1038
rect 373 -1075 374 -1067
rect 289 -1075 290 -1069
rect 352 -1070 353 -1038
rect 352 -1075 353 -1071
rect 436 -1072 437 -1038
rect 345 -1075 346 -1073
rect 436 -1075 437 -1073
rect 30 -1085 31 -1083
rect 44 -1085 45 -1083
rect 47 -1085 48 -1083
rect 61 -1085 62 -1083
rect 79 -1085 80 -1083
rect 79 -1108 80 -1084
rect 79 -1085 80 -1083
rect 79 -1108 80 -1084
rect 86 -1085 87 -1083
rect 89 -1108 90 -1084
rect 96 -1085 97 -1083
rect 177 -1085 178 -1083
rect 184 -1085 185 -1083
rect 184 -1108 185 -1084
rect 184 -1085 185 -1083
rect 184 -1108 185 -1084
rect 191 -1085 192 -1083
rect 208 -1108 209 -1084
rect 212 -1085 213 -1083
rect 324 -1085 325 -1083
rect 338 -1085 339 -1083
rect 401 -1085 402 -1083
rect 432 -1108 433 -1084
rect 464 -1085 465 -1083
rect 471 -1085 472 -1083
rect 478 -1085 479 -1083
rect 481 -1085 482 -1083
rect 485 -1085 486 -1083
rect 495 -1085 496 -1083
rect 499 -1085 500 -1083
rect 37 -1087 38 -1083
rect 201 -1087 202 -1083
rect 212 -1108 213 -1086
rect 341 -1087 342 -1083
rect 345 -1108 346 -1086
rect 387 -1087 388 -1083
rect 401 -1108 402 -1086
rect 457 -1087 458 -1083
rect 51 -1089 52 -1083
rect 65 -1089 66 -1083
rect 100 -1089 101 -1083
rect 159 -1089 160 -1083
rect 170 -1089 171 -1083
rect 247 -1089 248 -1083
rect 271 -1089 272 -1083
rect 310 -1089 311 -1083
rect 338 -1108 339 -1088
rect 373 -1089 374 -1083
rect 436 -1089 437 -1083
rect 436 -1108 437 -1088
rect 436 -1089 437 -1083
rect 436 -1108 437 -1088
rect 450 -1089 451 -1083
rect 457 -1108 458 -1088
rect 58 -1091 59 -1083
rect 110 -1091 111 -1083
rect 114 -1108 115 -1090
rect 135 -1091 136 -1083
rect 149 -1091 150 -1083
rect 240 -1091 241 -1083
rect 271 -1108 272 -1090
rect 331 -1091 332 -1083
rect 348 -1091 349 -1083
rect 380 -1091 381 -1083
rect 65 -1108 66 -1092
rect 72 -1093 73 -1083
rect 100 -1108 101 -1092
rect 121 -1093 122 -1083
rect 124 -1108 125 -1092
rect 135 -1108 136 -1092
rect 149 -1108 150 -1092
rect 226 -1093 227 -1083
rect 229 -1093 230 -1083
rect 317 -1093 318 -1083
rect 352 -1093 353 -1083
rect 387 -1108 388 -1092
rect 72 -1108 73 -1094
rect 86 -1108 87 -1094
rect 128 -1095 129 -1083
rect 128 -1108 129 -1094
rect 128 -1095 129 -1083
rect 128 -1108 129 -1094
rect 163 -1095 164 -1083
rect 170 -1108 171 -1094
rect 173 -1095 174 -1083
rect 236 -1095 237 -1083
rect 240 -1108 241 -1094
rect 247 -1108 248 -1094
rect 268 -1108 269 -1094
rect 317 -1108 318 -1094
rect 366 -1095 367 -1083
rect 376 -1105 377 -1094
rect 380 -1108 381 -1094
rect 415 -1095 416 -1083
rect 82 -1108 83 -1096
rect 121 -1108 122 -1096
rect 156 -1097 157 -1083
rect 163 -1108 164 -1096
rect 177 -1108 178 -1096
rect 222 -1097 223 -1083
rect 226 -1108 227 -1096
rect 331 -1108 332 -1096
rect 366 -1108 367 -1096
rect 443 -1097 444 -1083
rect 156 -1108 157 -1098
rect 278 -1099 279 -1083
rect 289 -1108 290 -1098
rect 359 -1099 360 -1083
rect 369 -1108 370 -1098
rect 429 -1099 430 -1083
rect 194 -1101 195 -1083
rect 215 -1101 216 -1083
rect 236 -1108 237 -1100
rect 254 -1101 255 -1083
rect 275 -1108 276 -1100
rect 296 -1101 297 -1083
rect 303 -1101 304 -1083
rect 303 -1108 304 -1100
rect 303 -1101 304 -1083
rect 303 -1108 304 -1100
rect 310 -1108 311 -1100
rect 324 -1108 325 -1100
rect 359 -1108 360 -1100
rect 394 -1101 395 -1083
rect 422 -1101 423 -1083
rect 443 -1108 444 -1100
rect 107 -1108 108 -1102
rect 215 -1108 216 -1102
rect 233 -1108 234 -1102
rect 254 -1108 255 -1102
rect 261 -1103 262 -1083
rect 296 -1108 297 -1102
rect 373 -1108 374 -1102
rect 408 -1103 409 -1083
rect 145 -1105 146 -1083
rect 261 -1108 262 -1104
rect 422 -1108 423 -1104
rect 205 -1107 206 -1083
rect 222 -1108 223 -1106
rect 394 -1108 395 -1106
rect 415 -1108 416 -1106
rect 47 -1118 48 -1116
rect 51 -1141 52 -1117
rect 72 -1118 73 -1116
rect 82 -1141 83 -1117
rect 93 -1118 94 -1116
rect 93 -1141 94 -1117
rect 93 -1118 94 -1116
rect 93 -1141 94 -1117
rect 100 -1118 101 -1116
rect 124 -1118 125 -1116
rect 149 -1118 150 -1116
rect 208 -1118 209 -1116
rect 212 -1118 213 -1116
rect 222 -1141 223 -1117
rect 229 -1118 230 -1116
rect 313 -1118 314 -1116
rect 334 -1118 335 -1116
rect 387 -1118 388 -1116
rect 394 -1141 395 -1117
rect 401 -1118 402 -1116
rect 408 -1118 409 -1116
rect 443 -1118 444 -1116
rect 65 -1120 66 -1116
rect 72 -1141 73 -1119
rect 100 -1141 101 -1119
rect 268 -1120 269 -1116
rect 285 -1120 286 -1116
rect 296 -1120 297 -1116
rect 306 -1141 307 -1119
rect 331 -1120 332 -1116
rect 338 -1120 339 -1116
rect 397 -1120 398 -1116
rect 408 -1141 409 -1119
rect 415 -1120 416 -1116
rect 422 -1120 423 -1116
rect 450 -1120 451 -1116
rect 65 -1141 66 -1121
rect 75 -1141 76 -1121
rect 110 -1141 111 -1121
rect 121 -1141 122 -1121
rect 149 -1141 150 -1121
rect 226 -1122 227 -1116
rect 233 -1122 234 -1116
rect 257 -1141 258 -1121
rect 261 -1122 262 -1116
rect 261 -1141 262 -1121
rect 261 -1122 262 -1116
rect 261 -1141 262 -1121
rect 275 -1122 276 -1116
rect 296 -1141 297 -1121
rect 317 -1122 318 -1116
rect 338 -1141 339 -1121
rect 352 -1122 353 -1116
rect 359 -1122 360 -1116
rect 366 -1141 367 -1121
rect 401 -1141 402 -1121
rect 415 -1141 416 -1121
rect 432 -1122 433 -1116
rect 450 -1141 451 -1121
rect 457 -1122 458 -1116
rect 114 -1124 115 -1116
rect 142 -1124 143 -1116
rect 170 -1124 171 -1116
rect 282 -1141 283 -1123
rect 289 -1124 290 -1116
rect 310 -1124 311 -1116
rect 317 -1141 318 -1123
rect 380 -1124 381 -1116
rect 387 -1141 388 -1123
rect 404 -1141 405 -1123
rect 422 -1141 423 -1123
rect 436 -1124 437 -1116
rect 114 -1141 115 -1125
rect 128 -1126 129 -1116
rect 135 -1126 136 -1116
rect 142 -1141 143 -1125
rect 170 -1141 171 -1125
rect 229 -1141 230 -1125
rect 240 -1126 241 -1116
rect 271 -1126 272 -1116
rect 310 -1141 311 -1125
rect 345 -1126 346 -1116
rect 177 -1128 178 -1116
rect 201 -1128 202 -1116
rect 205 -1141 206 -1127
rect 233 -1141 234 -1127
rect 243 -1141 244 -1127
rect 352 -1141 353 -1127
rect 184 -1130 185 -1116
rect 191 -1130 192 -1116
rect 198 -1141 199 -1129
rect 240 -1141 241 -1129
rect 247 -1141 248 -1129
rect 303 -1130 304 -1116
rect 331 -1141 332 -1129
rect 373 -1130 374 -1116
rect 163 -1141 164 -1131
rect 191 -1141 192 -1131
rect 226 -1141 227 -1131
rect 383 -1141 384 -1131
rect 254 -1134 255 -1116
rect 275 -1141 276 -1133
rect 303 -1141 304 -1133
rect 359 -1141 360 -1133
rect 156 -1136 157 -1116
rect 254 -1141 255 -1135
rect 268 -1141 269 -1135
rect 289 -1141 290 -1135
rect 324 -1136 325 -1116
rect 373 -1141 374 -1135
rect 156 -1141 157 -1137
rect 194 -1138 195 -1116
rect 250 -1138 251 -1116
rect 324 -1141 325 -1137
rect 345 -1141 346 -1137
rect 369 -1138 370 -1116
rect 177 -1141 178 -1139
rect 194 -1141 195 -1139
rect 47 -1151 48 -1149
rect 51 -1151 52 -1149
rect 58 -1151 59 -1149
rect 82 -1151 83 -1149
rect 89 -1151 90 -1149
rect 107 -1151 108 -1149
rect 114 -1151 115 -1149
rect 184 -1151 185 -1149
rect 191 -1178 192 -1150
rect 205 -1178 206 -1150
rect 212 -1151 213 -1149
rect 296 -1151 297 -1149
rect 299 -1178 300 -1150
rect 387 -1178 388 -1150
rect 394 -1151 395 -1149
rect 404 -1151 405 -1149
rect 408 -1151 409 -1149
rect 418 -1178 419 -1150
rect 422 -1151 423 -1149
rect 422 -1178 423 -1150
rect 422 -1151 423 -1149
rect 422 -1178 423 -1150
rect 446 -1151 447 -1149
rect 450 -1151 451 -1149
rect 51 -1178 52 -1152
rect 61 -1178 62 -1152
rect 65 -1153 66 -1149
rect 86 -1153 87 -1149
rect 107 -1178 108 -1152
rect 128 -1153 129 -1149
rect 135 -1153 136 -1149
rect 149 -1153 150 -1149
rect 170 -1153 171 -1149
rect 184 -1178 185 -1152
rect 194 -1178 195 -1152
rect 282 -1153 283 -1149
rect 303 -1178 304 -1152
rect 373 -1153 374 -1149
rect 65 -1178 66 -1154
rect 187 -1155 188 -1149
rect 212 -1178 213 -1154
rect 236 -1178 237 -1154
rect 240 -1155 241 -1149
rect 338 -1155 339 -1149
rect 100 -1157 101 -1149
rect 135 -1178 136 -1156
rect 142 -1157 143 -1149
rect 145 -1178 146 -1156
rect 177 -1157 178 -1149
rect 208 -1157 209 -1149
rect 222 -1157 223 -1149
rect 233 -1157 234 -1149
rect 243 -1157 244 -1149
rect 261 -1157 262 -1149
rect 271 -1157 272 -1149
rect 317 -1157 318 -1149
rect 324 -1157 325 -1149
rect 327 -1177 328 -1156
rect 338 -1178 339 -1156
rect 366 -1157 367 -1149
rect 100 -1178 101 -1158
rect 215 -1159 216 -1149
rect 226 -1159 227 -1149
rect 345 -1159 346 -1149
rect 359 -1159 360 -1149
rect 366 -1178 367 -1158
rect 117 -1178 118 -1160
rect 121 -1161 122 -1149
rect 128 -1178 129 -1160
rect 243 -1178 244 -1160
rect 247 -1161 248 -1149
rect 359 -1178 360 -1160
rect 121 -1178 122 -1162
rect 156 -1163 157 -1149
rect 226 -1178 227 -1162
rect 282 -1178 283 -1162
rect 306 -1163 307 -1149
rect 373 -1178 374 -1162
rect 156 -1178 157 -1164
rect 163 -1165 164 -1149
rect 229 -1165 230 -1149
rect 268 -1165 269 -1149
rect 275 -1165 276 -1149
rect 275 -1178 276 -1164
rect 275 -1165 276 -1149
rect 275 -1178 276 -1164
rect 310 -1165 311 -1149
rect 380 -1178 381 -1164
rect 198 -1167 199 -1149
rect 268 -1178 269 -1166
rect 296 -1178 297 -1166
rect 310 -1178 311 -1166
rect 313 -1167 314 -1149
rect 415 -1167 416 -1149
rect 233 -1178 234 -1168
rect 289 -1169 290 -1149
rect 317 -1178 318 -1168
rect 401 -1169 402 -1149
rect 415 -1178 416 -1168
rect 429 -1178 430 -1168
rect 254 -1178 255 -1170
rect 261 -1178 262 -1170
rect 324 -1178 325 -1170
rect 331 -1171 332 -1149
rect 352 -1171 353 -1149
rect 401 -1178 402 -1170
rect 247 -1178 248 -1172
rect 352 -1178 353 -1172
rect 257 -1175 258 -1149
rect 394 -1178 395 -1174
rect 331 -1178 332 -1176
rect 47 -1188 48 -1186
rect 47 -1205 48 -1187
rect 47 -1188 48 -1186
rect 47 -1205 48 -1187
rect 51 -1188 52 -1186
rect 68 -1205 69 -1187
rect 72 -1205 73 -1187
rect 75 -1188 76 -1186
rect 89 -1188 90 -1186
rect 96 -1205 97 -1187
rect 100 -1188 101 -1186
rect 142 -1188 143 -1186
rect 156 -1188 157 -1186
rect 222 -1188 223 -1186
rect 229 -1188 230 -1186
rect 275 -1188 276 -1186
rect 289 -1188 290 -1186
rect 324 -1188 325 -1186
rect 338 -1188 339 -1186
rect 348 -1188 349 -1186
rect 380 -1188 381 -1186
rect 380 -1205 381 -1187
rect 380 -1188 381 -1186
rect 380 -1205 381 -1187
rect 408 -1205 409 -1187
rect 415 -1188 416 -1186
rect 422 -1188 423 -1186
rect 425 -1192 426 -1187
rect 65 -1205 66 -1189
rect 82 -1205 83 -1189
rect 93 -1190 94 -1186
rect 100 -1205 101 -1189
rect 107 -1190 108 -1186
rect 149 -1190 150 -1186
rect 166 -1190 167 -1186
rect 198 -1205 199 -1189
rect 205 -1190 206 -1186
rect 205 -1205 206 -1189
rect 205 -1190 206 -1186
rect 205 -1205 206 -1189
rect 212 -1190 213 -1186
rect 212 -1205 213 -1189
rect 212 -1190 213 -1186
rect 212 -1205 213 -1189
rect 219 -1205 220 -1189
rect 310 -1190 311 -1186
rect 324 -1205 325 -1189
rect 352 -1190 353 -1186
rect 422 -1205 423 -1189
rect 429 -1190 430 -1186
rect 79 -1192 80 -1186
rect 166 -1205 167 -1191
rect 170 -1205 171 -1191
rect 177 -1192 178 -1186
rect 184 -1192 185 -1186
rect 201 -1192 202 -1186
rect 229 -1205 230 -1191
rect 254 -1205 255 -1191
rect 268 -1192 269 -1186
rect 292 -1192 293 -1186
rect 303 -1192 304 -1186
rect 331 -1192 332 -1186
rect 345 -1192 346 -1186
rect 387 -1192 388 -1186
rect 429 -1205 430 -1191
rect 79 -1205 80 -1193
rect 114 -1205 115 -1193
rect 121 -1194 122 -1186
rect 152 -1194 153 -1186
rect 159 -1205 160 -1193
rect 177 -1205 178 -1193
rect 240 -1194 241 -1186
rect 317 -1194 318 -1186
rect 331 -1205 332 -1193
rect 341 -1205 342 -1193
rect 345 -1205 346 -1193
rect 401 -1194 402 -1186
rect 107 -1205 108 -1195
rect 145 -1205 146 -1195
rect 149 -1205 150 -1195
rect 191 -1196 192 -1186
rect 233 -1205 234 -1195
rect 240 -1205 241 -1195
rect 247 -1205 248 -1195
rect 261 -1196 262 -1186
rect 282 -1196 283 -1186
rect 303 -1205 304 -1195
rect 317 -1205 318 -1195
rect 373 -1196 374 -1186
rect 128 -1198 129 -1186
rect 226 -1198 227 -1186
rect 236 -1198 237 -1186
rect 282 -1205 283 -1197
rect 289 -1205 290 -1197
rect 359 -1198 360 -1186
rect 128 -1205 129 -1199
rect 156 -1205 157 -1199
rect 184 -1205 185 -1199
rect 226 -1205 227 -1199
rect 292 -1205 293 -1199
rect 296 -1205 297 -1199
rect 359 -1205 360 -1199
rect 366 -1200 367 -1186
rect 135 -1202 136 -1186
rect 173 -1202 174 -1186
rect 366 -1205 367 -1201
rect 394 -1202 395 -1186
rect 121 -1205 122 -1203
rect 135 -1205 136 -1203
rect 138 -1205 139 -1203
rect 222 -1205 223 -1203
rect 33 -1228 34 -1214
rect 37 -1228 38 -1214
rect 44 -1228 45 -1214
rect 51 -1228 52 -1214
rect 58 -1228 59 -1214
rect 65 -1228 66 -1214
rect 72 -1215 73 -1213
rect 79 -1215 80 -1213
rect 89 -1215 90 -1213
rect 100 -1215 101 -1213
rect 107 -1215 108 -1213
rect 173 -1228 174 -1214
rect 180 -1228 181 -1214
rect 205 -1215 206 -1213
rect 229 -1215 230 -1213
rect 247 -1215 248 -1213
rect 254 -1215 255 -1213
rect 268 -1228 269 -1214
rect 303 -1215 304 -1213
rect 341 -1215 342 -1213
rect 359 -1215 360 -1213
rect 359 -1228 360 -1214
rect 359 -1215 360 -1213
rect 359 -1228 360 -1214
rect 373 -1215 374 -1213
rect 380 -1215 381 -1213
rect 401 -1228 402 -1214
rect 408 -1215 409 -1213
rect 422 -1228 423 -1214
rect 429 -1215 430 -1213
rect 72 -1228 73 -1216
rect 79 -1228 80 -1216
rect 93 -1228 94 -1216
rect 138 -1217 139 -1213
rect 152 -1217 153 -1213
rect 159 -1217 160 -1213
rect 163 -1217 164 -1213
rect 212 -1217 213 -1213
rect 229 -1228 230 -1216
rect 240 -1228 241 -1216
rect 243 -1217 244 -1213
rect 292 -1217 293 -1213
rect 296 -1217 297 -1213
rect 303 -1228 304 -1216
rect 306 -1217 307 -1213
rect 324 -1217 325 -1213
rect 331 -1217 332 -1213
rect 352 -1217 353 -1213
rect 425 -1217 426 -1213
rect 432 -1228 433 -1216
rect 114 -1219 115 -1213
rect 121 -1219 122 -1213
rect 128 -1219 129 -1213
rect 142 -1219 143 -1213
rect 163 -1228 164 -1218
rect 177 -1219 178 -1213
rect 184 -1228 185 -1218
rect 201 -1228 202 -1218
rect 212 -1228 213 -1218
rect 254 -1228 255 -1218
rect 275 -1228 276 -1218
rect 292 -1228 293 -1218
rect 310 -1219 311 -1213
rect 345 -1219 346 -1213
rect 352 -1228 353 -1218
rect 366 -1219 367 -1213
rect 100 -1228 101 -1220
rect 128 -1228 129 -1220
rect 135 -1221 136 -1213
rect 156 -1221 157 -1213
rect 170 -1221 171 -1213
rect 187 -1221 188 -1213
rect 191 -1228 192 -1220
rect 222 -1221 223 -1213
rect 282 -1221 283 -1213
rect 310 -1228 311 -1220
rect 317 -1221 318 -1213
rect 320 -1228 321 -1220
rect 338 -1228 339 -1220
rect 345 -1228 346 -1220
rect 366 -1228 367 -1220
rect 373 -1228 374 -1220
rect 121 -1228 122 -1222
rect 149 -1228 150 -1222
rect 194 -1223 195 -1213
rect 198 -1223 199 -1213
rect 215 -1228 216 -1222
rect 317 -1228 318 -1222
rect 124 -1228 125 -1224
rect 142 -1228 143 -1224
rect 222 -1228 223 -1224
rect 233 -1225 234 -1213
rect 282 -1228 283 -1224
rect 313 -1225 314 -1213
rect 219 -1228 220 -1226
rect 233 -1228 234 -1226
rect 23 -1238 24 -1236
rect 23 -1253 24 -1237
rect 23 -1238 24 -1236
rect 23 -1253 24 -1237
rect 30 -1253 31 -1237
rect 37 -1238 38 -1236
rect 44 -1253 45 -1237
rect 51 -1238 52 -1236
rect 58 -1238 59 -1236
rect 58 -1253 59 -1237
rect 58 -1238 59 -1236
rect 58 -1253 59 -1237
rect 65 -1238 66 -1236
rect 75 -1253 76 -1237
rect 79 -1238 80 -1236
rect 79 -1253 80 -1237
rect 79 -1238 80 -1236
rect 79 -1253 80 -1237
rect 93 -1238 94 -1236
rect 117 -1238 118 -1236
rect 128 -1238 129 -1236
rect 149 -1238 150 -1236
rect 152 -1253 153 -1237
rect 208 -1238 209 -1236
rect 222 -1238 223 -1236
rect 268 -1238 269 -1236
rect 275 -1238 276 -1236
rect 289 -1253 290 -1237
rect 299 -1238 300 -1236
rect 310 -1238 311 -1236
rect 324 -1253 325 -1237
rect 327 -1238 328 -1236
rect 334 -1253 335 -1237
rect 338 -1238 339 -1236
rect 359 -1238 360 -1236
rect 359 -1253 360 -1237
rect 359 -1238 360 -1236
rect 359 -1253 360 -1237
rect 369 -1253 370 -1237
rect 373 -1238 374 -1236
rect 401 -1238 402 -1236
rect 408 -1238 409 -1236
rect 415 -1238 416 -1236
rect 422 -1238 423 -1236
rect 100 -1240 101 -1236
rect 114 -1240 115 -1236
rect 128 -1253 129 -1239
rect 138 -1240 139 -1236
rect 142 -1240 143 -1236
rect 145 -1253 146 -1239
rect 159 -1240 160 -1236
rect 159 -1253 160 -1239
rect 159 -1240 160 -1236
rect 159 -1253 160 -1239
rect 163 -1240 164 -1236
rect 215 -1240 216 -1236
rect 226 -1253 227 -1239
rect 278 -1253 279 -1239
rect 303 -1240 304 -1236
rect 303 -1253 304 -1239
rect 303 -1240 304 -1236
rect 303 -1253 304 -1239
rect 338 -1253 339 -1239
rect 352 -1240 353 -1236
rect 103 -1253 104 -1241
rect 121 -1253 122 -1241
rect 177 -1253 178 -1241
rect 191 -1242 192 -1236
rect 194 -1253 195 -1241
rect 240 -1242 241 -1236
rect 250 -1242 251 -1236
rect 268 -1253 269 -1241
rect 110 -1244 111 -1236
rect 114 -1253 115 -1243
rect 205 -1244 206 -1236
rect 282 -1244 283 -1236
rect 208 -1253 209 -1245
rect 254 -1246 255 -1236
rect 261 -1246 262 -1236
rect 261 -1253 262 -1245
rect 261 -1246 262 -1236
rect 261 -1253 262 -1245
rect 212 -1253 213 -1247
rect 222 -1253 223 -1247
rect 233 -1248 234 -1236
rect 257 -1253 258 -1247
rect 170 -1250 171 -1236
rect 233 -1253 234 -1249
rect 170 -1253 171 -1251
rect 184 -1252 185 -1236
rect 219 -1253 220 -1251
rect 240 -1253 241 -1251
rect 30 -1263 31 -1261
rect 37 -1263 38 -1261
rect 58 -1263 59 -1261
rect 68 -1263 69 -1261
rect 72 -1263 73 -1261
rect 79 -1263 80 -1261
rect 107 -1263 108 -1261
rect 114 -1263 115 -1261
rect 121 -1263 122 -1261
rect 152 -1263 153 -1261
rect 170 -1263 171 -1261
rect 205 -1263 206 -1261
rect 208 -1263 209 -1261
rect 212 -1263 213 -1261
rect 226 -1263 227 -1261
rect 268 -1263 269 -1261
rect 285 -1263 286 -1261
rect 289 -1263 290 -1261
rect 296 -1263 297 -1261
rect 303 -1263 304 -1261
rect 317 -1263 318 -1261
rect 324 -1263 325 -1261
rect 338 -1263 339 -1261
rect 348 -1263 349 -1261
rect 355 -1263 356 -1261
rect 359 -1263 360 -1261
rect 128 -1265 129 -1261
rect 138 -1265 139 -1261
rect 142 -1265 143 -1261
rect 163 -1265 164 -1261
rect 177 -1265 178 -1261
rect 187 -1265 188 -1261
rect 198 -1265 199 -1261
rect 233 -1265 234 -1261
rect 250 -1265 251 -1261
rect 261 -1265 262 -1261
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=28
rlabel pdiffusion 10 -8 10 -8 0 cellNo=121
rlabel pdiffusion 17 -8 17 -8 0 cellNo=40
rlabel pdiffusion 24 -8 24 -8 0 cellNo=278
rlabel pdiffusion 31 -8 31 -8 0 cellNo=60
rlabel pdiffusion 38 -8 38 -8 0 cellNo=335
rlabel pdiffusion 45 -8 45 -8 0 cellNo=473
rlabel pdiffusion 52 -8 52 -8 0 cellNo=381
rlabel pdiffusion 59 -8 59 -8 0 cellNo=595
rlabel pdiffusion 66 -8 66 -8 0 cellNo=795
rlabel pdiffusion 136 -8 136 -8 0 cellNo=803
rlabel pdiffusion 143 -8 143 -8 0 cellNo=102
rlabel pdiffusion 150 -8 150 -8 0 feedthrough
rlabel pdiffusion 178 -8 178 -8 0 feedthrough
rlabel pdiffusion 185 -8 185 -8 0 cellNo=207
rlabel pdiffusion 192 -8 192 -8 0 cellNo=339
rlabel pdiffusion 199 -8 199 -8 0 feedthrough
rlabel pdiffusion 206 -8 206 -8 0 cellNo=619
rlabel pdiffusion 213 -8 213 -8 0 cellNo=14
rlabel pdiffusion 220 -8 220 -8 0 feedthrough
rlabel pdiffusion 227 -8 227 -8 0 cellNo=178
rlabel pdiffusion 234 -8 234 -8 0 cellNo=209
rlabel pdiffusion 241 -8 241 -8 0 feedthrough
rlabel pdiffusion 3 -27 3 -27 0 cellNo=35
rlabel pdiffusion 10 -27 10 -27 0 cellNo=475
rlabel pdiffusion 17 -27 17 -27 0 cellNo=47
rlabel pdiffusion 24 -27 24 -27 0 cellNo=49
rlabel pdiffusion 31 -27 31 -27 0 cellNo=267
rlabel pdiffusion 38 -27 38 -27 0 cellNo=322
rlabel pdiffusion 45 -27 45 -27 0 cellNo=293
rlabel pdiffusion 52 -27 52 -27 0 cellNo=441
rlabel pdiffusion 59 -27 59 -27 0 cellNo=671
rlabel pdiffusion 66 -27 66 -27 0 cellNo=764
rlabel pdiffusion 129 -27 129 -27 0 cellNo=17
rlabel pdiffusion 136 -27 136 -27 0 feedthrough
rlabel pdiffusion 143 -27 143 -27 0 feedthrough
rlabel pdiffusion 150 -27 150 -27 0 cellNo=575
rlabel pdiffusion 157 -27 157 -27 0 cellNo=480
rlabel pdiffusion 164 -27 164 -27 0 feedthrough
rlabel pdiffusion 171 -27 171 -27 0 cellNo=311
rlabel pdiffusion 178 -27 178 -27 0 feedthrough
rlabel pdiffusion 185 -27 185 -27 0 cellNo=80
rlabel pdiffusion 192 -27 192 -27 0 cellNo=606
rlabel pdiffusion 199 -27 199 -27 0 feedthrough
rlabel pdiffusion 206 -27 206 -27 0 feedthrough
rlabel pdiffusion 213 -27 213 -27 0 cellNo=413
rlabel pdiffusion 220 -27 220 -27 0 cellNo=642
rlabel pdiffusion 227 -27 227 -27 0 cellNo=783
rlabel pdiffusion 234 -27 234 -27 0 feedthrough
rlabel pdiffusion 241 -27 241 -27 0 feedthrough
rlabel pdiffusion 248 -27 248 -27 0 cellNo=711
rlabel pdiffusion 255 -27 255 -27 0 cellNo=26
rlabel pdiffusion 297 -27 297 -27 0 cellNo=53
rlabel pdiffusion 325 -27 325 -27 0 cellNo=784
rlabel pdiffusion 332 -27 332 -27 0 feedthrough
rlabel pdiffusion 3 -54 3 -54 0 cellNo=68
rlabel pdiffusion 10 -54 10 -54 0 cellNo=542
rlabel pdiffusion 17 -54 17 -54 0 cellNo=219
rlabel pdiffusion 24 -54 24 -54 0 cellNo=479
rlabel pdiffusion 31 -54 31 -54 0 cellNo=409
rlabel pdiffusion 38 -54 38 -54 0 cellNo=695
rlabel pdiffusion 45 -54 45 -54 0 cellNo=292
rlabel pdiffusion 52 -54 52 -54 0 cellNo=366
rlabel pdiffusion 59 -54 59 -54 0 cellNo=430
rlabel pdiffusion 66 -54 66 -54 0 cellNo=780
rlabel pdiffusion 73 -54 73 -54 0 cellNo=756
rlabel pdiffusion 136 -54 136 -54 0 feedthrough
rlabel pdiffusion 143 -54 143 -54 0 cellNo=66
rlabel pdiffusion 150 -54 150 -54 0 cellNo=252
rlabel pdiffusion 157 -54 157 -54 0 cellNo=222
rlabel pdiffusion 164 -54 164 -54 0 cellNo=894
rlabel pdiffusion 171 -54 171 -54 0 cellNo=86
rlabel pdiffusion 178 -54 178 -54 0 cellNo=208
rlabel pdiffusion 185 -54 185 -54 0 feedthrough
rlabel pdiffusion 192 -54 192 -54 0 feedthrough
rlabel pdiffusion 199 -54 199 -54 0 cellNo=215
rlabel pdiffusion 206 -54 206 -54 0 cellNo=376
rlabel pdiffusion 213 -54 213 -54 0 feedthrough
rlabel pdiffusion 220 -54 220 -54 0 cellNo=31
rlabel pdiffusion 227 -54 227 -54 0 cellNo=9
rlabel pdiffusion 234 -54 234 -54 0 feedthrough
rlabel pdiffusion 241 -54 241 -54 0 feedthrough
rlabel pdiffusion 248 -54 248 -54 0 feedthrough
rlabel pdiffusion 255 -54 255 -54 0 cellNo=538
rlabel pdiffusion 262 -54 262 -54 0 feedthrough
rlabel pdiffusion 269 -54 269 -54 0 cellNo=844
rlabel pdiffusion 276 -54 276 -54 0 cellNo=808
rlabel pdiffusion 283 -54 283 -54 0 feedthrough
rlabel pdiffusion 290 -54 290 -54 0 feedthrough
rlabel pdiffusion 297 -54 297 -54 0 cellNo=128
rlabel pdiffusion 304 -54 304 -54 0 feedthrough
rlabel pdiffusion 325 -54 325 -54 0 feedthrough
rlabel pdiffusion 332 -54 332 -54 0 feedthrough
rlabel pdiffusion 3 -77 3 -77 0 cellNo=73
rlabel pdiffusion 10 -77 10 -77 0 cellNo=372
rlabel pdiffusion 17 -77 17 -77 0 cellNo=91
rlabel pdiffusion 24 -77 24 -77 0 cellNo=838
rlabel pdiffusion 31 -77 31 -77 0 cellNo=109
rlabel pdiffusion 38 -77 38 -77 0 cellNo=262
rlabel pdiffusion 45 -77 45 -77 0 cellNo=365
rlabel pdiffusion 52 -77 52 -77 0 cellNo=424
rlabel pdiffusion 87 -77 87 -77 0 cellNo=116
rlabel pdiffusion 101 -77 101 -77 0 cellNo=82
rlabel pdiffusion 108 -77 108 -77 0 feedthrough
rlabel pdiffusion 115 -77 115 -77 0 cellNo=87
rlabel pdiffusion 122 -77 122 -77 0 feedthrough
rlabel pdiffusion 129 -77 129 -77 0 feedthrough
rlabel pdiffusion 136 -77 136 -77 0 cellNo=503
rlabel pdiffusion 143 -77 143 -77 0 cellNo=744
rlabel pdiffusion 150 -77 150 -77 0 feedthrough
rlabel pdiffusion 157 -77 157 -77 0 cellNo=285
rlabel pdiffusion 164 -77 164 -77 0 cellNo=225
rlabel pdiffusion 171 -77 171 -77 0 feedthrough
rlabel pdiffusion 178 -77 178 -77 0 feedthrough
rlabel pdiffusion 185 -77 185 -77 0 cellNo=297
rlabel pdiffusion 192 -77 192 -77 0 feedthrough
rlabel pdiffusion 199 -77 199 -77 0 cellNo=246
rlabel pdiffusion 206 -77 206 -77 0 feedthrough
rlabel pdiffusion 213 -77 213 -77 0 cellNo=5
rlabel pdiffusion 220 -77 220 -77 0 cellNo=440
rlabel pdiffusion 227 -77 227 -77 0 cellNo=343
rlabel pdiffusion 234 -77 234 -77 0 cellNo=351
rlabel pdiffusion 241 -77 241 -77 0 feedthrough
rlabel pdiffusion 248 -77 248 -77 0 cellNo=257
rlabel pdiffusion 255 -77 255 -77 0 feedthrough
rlabel pdiffusion 262 -77 262 -77 0 feedthrough
rlabel pdiffusion 269 -77 269 -77 0 cellNo=593
rlabel pdiffusion 276 -77 276 -77 0 feedthrough
rlabel pdiffusion 283 -77 283 -77 0 feedthrough
rlabel pdiffusion 290 -77 290 -77 0 cellNo=407
rlabel pdiffusion 297 -77 297 -77 0 feedthrough
rlabel pdiffusion 304 -77 304 -77 0 cellNo=305
rlabel pdiffusion 311 -77 311 -77 0 cellNo=747
rlabel pdiffusion 318 -77 318 -77 0 cellNo=327
rlabel pdiffusion 325 -77 325 -77 0 feedthrough
rlabel pdiffusion 332 -77 332 -77 0 feedthrough
rlabel pdiffusion 3 -102 3 -102 0 cellNo=99
rlabel pdiffusion 10 -102 10 -102 0 cellNo=871
rlabel pdiffusion 17 -102 17 -102 0 cellNo=281
rlabel pdiffusion 24 -102 24 -102 0 cellNo=801
rlabel pdiffusion 31 -102 31 -102 0 cellNo=228
rlabel pdiffusion 38 -102 38 -102 0 cellNo=354
rlabel pdiffusion 45 -102 45 -102 0 cellNo=857
rlabel pdiffusion 52 -102 52 -102 0 cellNo=561
rlabel pdiffusion 87 -102 87 -102 0 cellNo=94
rlabel pdiffusion 101 -102 101 -102 0 cellNo=348
rlabel pdiffusion 108 -102 108 -102 0 feedthrough
rlabel pdiffusion 115 -102 115 -102 0 feedthrough
rlabel pdiffusion 122 -102 122 -102 0 cellNo=146
rlabel pdiffusion 129 -102 129 -102 0 cellNo=180
rlabel pdiffusion 136 -102 136 -102 0 feedthrough
rlabel pdiffusion 143 -102 143 -102 0 cellNo=417
rlabel pdiffusion 150 -102 150 -102 0 feedthrough
rlabel pdiffusion 157 -102 157 -102 0 cellNo=179
rlabel pdiffusion 164 -102 164 -102 0 cellNo=571
rlabel pdiffusion 171 -102 171 -102 0 cellNo=644
rlabel pdiffusion 178 -102 178 -102 0 cellNo=419
rlabel pdiffusion 185 -102 185 -102 0 feedthrough
rlabel pdiffusion 192 -102 192 -102 0 cellNo=504
rlabel pdiffusion 199 -102 199 -102 0 feedthrough
rlabel pdiffusion 206 -102 206 -102 0 cellNo=617
rlabel pdiffusion 213 -102 213 -102 0 cellNo=646
rlabel pdiffusion 220 -102 220 -102 0 cellNo=570
rlabel pdiffusion 227 -102 227 -102 0 cellNo=481
rlabel pdiffusion 234 -102 234 -102 0 feedthrough
rlabel pdiffusion 241 -102 241 -102 0 cellNo=12
rlabel pdiffusion 248 -102 248 -102 0 feedthrough
rlabel pdiffusion 255 -102 255 -102 0 feedthrough
rlabel pdiffusion 262 -102 262 -102 0 feedthrough
rlabel pdiffusion 269 -102 269 -102 0 cellNo=133
rlabel pdiffusion 276 -102 276 -102 0 feedthrough
rlabel pdiffusion 283 -102 283 -102 0 cellNo=467
rlabel pdiffusion 290 -102 290 -102 0 cellNo=229
rlabel pdiffusion 297 -102 297 -102 0 feedthrough
rlabel pdiffusion 304 -102 304 -102 0 feedthrough
rlabel pdiffusion 311 -102 311 -102 0 feedthrough
rlabel pdiffusion 318 -102 318 -102 0 feedthrough
rlabel pdiffusion 325 -102 325 -102 0 cellNo=63
rlabel pdiffusion 381 -102 381 -102 0 cellNo=898
rlabel pdiffusion 3 -127 3 -127 0 cellNo=167
rlabel pdiffusion 10 -127 10 -127 0 cellNo=469
rlabel pdiffusion 17 -127 17 -127 0 cellNo=536
rlabel pdiffusion 24 -127 24 -127 0 cellNo=195
rlabel pdiffusion 31 -127 31 -127 0 cellNo=416
rlabel pdiffusion 38 -127 38 -127 0 cellNo=408
rlabel pdiffusion 45 -127 45 -127 0 cellNo=559
rlabel pdiffusion 80 -127 80 -127 0 cellNo=300
rlabel pdiffusion 87 -127 87 -127 0 cellNo=449
rlabel pdiffusion 101 -127 101 -127 0 cellNo=177
rlabel pdiffusion 108 -127 108 -127 0 feedthrough
rlabel pdiffusion 115 -127 115 -127 0 cellNo=224
rlabel pdiffusion 122 -127 122 -127 0 cellNo=718
rlabel pdiffusion 129 -127 129 -127 0 cellNo=43
rlabel pdiffusion 136 -127 136 -127 0 feedthrough
rlabel pdiffusion 143 -127 143 -127 0 cellNo=338
rlabel pdiffusion 150 -127 150 -127 0 cellNo=615
rlabel pdiffusion 157 -127 157 -127 0 feedthrough
rlabel pdiffusion 164 -127 164 -127 0 feedthrough
rlabel pdiffusion 171 -127 171 -127 0 cellNo=221
rlabel pdiffusion 178 -127 178 -127 0 cellNo=142
rlabel pdiffusion 185 -127 185 -127 0 feedthrough
rlabel pdiffusion 192 -127 192 -127 0 cellNo=410
rlabel pdiffusion 199 -127 199 -127 0 feedthrough
rlabel pdiffusion 206 -127 206 -127 0 feedthrough
rlabel pdiffusion 213 -127 213 -127 0 cellNo=93
rlabel pdiffusion 220 -127 220 -127 0 feedthrough
rlabel pdiffusion 227 -127 227 -127 0 cellNo=582
rlabel pdiffusion 234 -127 234 -127 0 cellNo=727
rlabel pdiffusion 241 -127 241 -127 0 feedthrough
rlabel pdiffusion 255 -127 255 -127 0 feedthrough
rlabel pdiffusion 262 -127 262 -127 0 feedthrough
rlabel pdiffusion 269 -127 269 -127 0 feedthrough
rlabel pdiffusion 297 -127 297 -127 0 cellNo=876
rlabel pdiffusion 304 -127 304 -127 0 feedthrough
rlabel pdiffusion 311 -127 311 -127 0 cellNo=332
rlabel pdiffusion 318 -127 318 -127 0 feedthrough
rlabel pdiffusion 381 -127 381 -127 0 feedthrough
rlabel pdiffusion 3 -152 3 -152 0 cellNo=156
rlabel pdiffusion 10 -152 10 -152 0 cellNo=245
rlabel pdiffusion 17 -152 17 -152 0 cellNo=517
rlabel pdiffusion 24 -152 24 -152 0 cellNo=820
rlabel pdiffusion 31 -152 31 -152 0 cellNo=401
rlabel pdiffusion 38 -152 38 -152 0 cellNo=556
rlabel pdiffusion 45 -152 45 -152 0 cellNo=730
rlabel pdiffusion 80 -152 80 -152 0 cellNo=317
rlabel pdiffusion 108 -152 108 -152 0 feedthrough
rlabel pdiffusion 115 -152 115 -152 0 feedthrough
rlabel pdiffusion 122 -152 122 -152 0 feedthrough
rlabel pdiffusion 129 -152 129 -152 0 cellNo=653
rlabel pdiffusion 136 -152 136 -152 0 cellNo=85
rlabel pdiffusion 143 -152 143 -152 0 cellNo=129
rlabel pdiffusion 150 -152 150 -152 0 cellNo=144
rlabel pdiffusion 157 -152 157 -152 0 cellNo=766
rlabel pdiffusion 164 -152 164 -152 0 feedthrough
rlabel pdiffusion 171 -152 171 -152 0 cellNo=388
rlabel pdiffusion 178 -152 178 -152 0 feedthrough
rlabel pdiffusion 185 -152 185 -152 0 cellNo=641
rlabel pdiffusion 192 -152 192 -152 0 feedthrough
rlabel pdiffusion 199 -152 199 -152 0 cellNo=635
rlabel pdiffusion 206 -152 206 -152 0 cellNo=147
rlabel pdiffusion 213 -152 213 -152 0 cellNo=119
rlabel pdiffusion 220 -152 220 -152 0 feedthrough
rlabel pdiffusion 227 -152 227 -152 0 feedthrough
rlabel pdiffusion 234 -152 234 -152 0 feedthrough
rlabel pdiffusion 241 -152 241 -152 0 cellNo=217
rlabel pdiffusion 255 -152 255 -152 0 cellNo=22
rlabel pdiffusion 262 -152 262 -152 0 feedthrough
rlabel pdiffusion 269 -152 269 -152 0 cellNo=123
rlabel pdiffusion 276 -152 276 -152 0 feedthrough
rlabel pdiffusion 311 -152 311 -152 0 cellNo=20
rlabel pdiffusion 318 -152 318 -152 0 cellNo=547
rlabel pdiffusion 325 -152 325 -152 0 feedthrough
rlabel pdiffusion 381 -152 381 -152 0 cellNo=452
rlabel pdiffusion 388 -152 388 -152 0 feedthrough
rlabel pdiffusion 3 -175 3 -175 0 cellNo=233
rlabel pdiffusion 10 -175 10 -175 0 cellNo=347
rlabel pdiffusion 17 -175 17 -175 0 cellNo=588
rlabel pdiffusion 24 -175 24 -175 0 cellNo=541
rlabel pdiffusion 31 -175 31 -175 0 cellNo=696
rlabel pdiffusion 80 -175 80 -175 0 cellNo=266
rlabel pdiffusion 115 -175 115 -175 0 cellNo=81
rlabel pdiffusion 122 -175 122 -175 0 cellNo=218
rlabel pdiffusion 129 -175 129 -175 0 cellNo=282
rlabel pdiffusion 136 -175 136 -175 0 feedthrough
rlabel pdiffusion 143 -175 143 -175 0 cellNo=304
rlabel pdiffusion 150 -175 150 -175 0 cellNo=751
rlabel pdiffusion 157 -175 157 -175 0 cellNo=150
rlabel pdiffusion 164 -175 164 -175 0 feedthrough
rlabel pdiffusion 171 -175 171 -175 0 feedthrough
rlabel pdiffusion 178 -175 178 -175 0 feedthrough
rlabel pdiffusion 185 -175 185 -175 0 cellNo=394
rlabel pdiffusion 192 -175 192 -175 0 cellNo=592
rlabel pdiffusion 199 -175 199 -175 0 feedthrough
rlabel pdiffusion 206 -175 206 -175 0 feedthrough
rlabel pdiffusion 213 -175 213 -175 0 cellNo=205
rlabel pdiffusion 220 -175 220 -175 0 feedthrough
rlabel pdiffusion 227 -175 227 -175 0 cellNo=537
rlabel pdiffusion 234 -175 234 -175 0 cellNo=140
rlabel pdiffusion 241 -175 241 -175 0 feedthrough
rlabel pdiffusion 248 -175 248 -175 0 feedthrough
rlabel pdiffusion 255 -175 255 -175 0 feedthrough
rlabel pdiffusion 262 -175 262 -175 0 feedthrough
rlabel pdiffusion 269 -175 269 -175 0 cellNo=640
rlabel pdiffusion 276 -175 276 -175 0 cellNo=519
rlabel pdiffusion 283 -175 283 -175 0 cellNo=896
rlabel pdiffusion 290 -175 290 -175 0 feedthrough
rlabel pdiffusion 297 -175 297 -175 0 feedthrough
rlabel pdiffusion 304 -175 304 -175 0 feedthrough
rlabel pdiffusion 311 -175 311 -175 0 cellNo=97
rlabel pdiffusion 318 -175 318 -175 0 feedthrough
rlabel pdiffusion 325 -175 325 -175 0 feedthrough
rlabel pdiffusion 332 -175 332 -175 0 feedthrough
rlabel pdiffusion 339 -175 339 -175 0 cellNo=143
rlabel pdiffusion 346 -175 346 -175 0 feedthrough
rlabel pdiffusion 353 -175 353 -175 0 cellNo=321
rlabel pdiffusion 360 -175 360 -175 0 cellNo=141
rlabel pdiffusion 367 -175 367 -175 0 feedthrough
rlabel pdiffusion 374 -175 374 -175 0 feedthrough
rlabel pdiffusion 381 -175 381 -175 0 cellNo=360
rlabel pdiffusion 388 -175 388 -175 0 feedthrough
rlabel pdiffusion 395 -175 395 -175 0 feedthrough
rlabel pdiffusion 409 -175 409 -175 0 cellNo=591
rlabel pdiffusion 416 -175 416 -175 0 feedthrough
rlabel pdiffusion 437 -175 437 -175 0 cellNo=235
rlabel pdiffusion 444 -175 444 -175 0 feedthrough
rlabel pdiffusion 3 -202 3 -202 0 cellNo=148
rlabel pdiffusion 10 -202 10 -202 0 cellNo=345
rlabel pdiffusion 17 -202 17 -202 0 cellNo=889
rlabel pdiffusion 24 -202 24 -202 0 cellNo=683
rlabel pdiffusion 73 -202 73 -202 0 cellNo=36
rlabel pdiffusion 80 -202 80 -202 0 feedthrough
rlabel pdiffusion 87 -202 87 -202 0 cellNo=654
rlabel pdiffusion 94 -202 94 -202 0 cellNo=601
rlabel pdiffusion 101 -202 101 -202 0 cellNo=201
rlabel pdiffusion 108 -202 108 -202 0 feedthrough
rlabel pdiffusion 115 -202 115 -202 0 cellNo=157
rlabel pdiffusion 122 -202 122 -202 0 feedthrough
rlabel pdiffusion 129 -202 129 -202 0 cellNo=170
rlabel pdiffusion 136 -202 136 -202 0 cellNo=135
rlabel pdiffusion 143 -202 143 -202 0 cellNo=426
rlabel pdiffusion 150 -202 150 -202 0 feedthrough
rlabel pdiffusion 157 -202 157 -202 0 feedthrough
rlabel pdiffusion 164 -202 164 -202 0 feedthrough
rlabel pdiffusion 171 -202 171 -202 0 feedthrough
rlabel pdiffusion 178 -202 178 -202 0 feedthrough
rlabel pdiffusion 185 -202 185 -202 0 feedthrough
rlabel pdiffusion 192 -202 192 -202 0 feedthrough
rlabel pdiffusion 199 -202 199 -202 0 cellNo=255
rlabel pdiffusion 206 -202 206 -202 0 cellNo=737
rlabel pdiffusion 213 -202 213 -202 0 cellNo=598
rlabel pdiffusion 220 -202 220 -202 0 cellNo=816
rlabel pdiffusion 227 -202 227 -202 0 cellNo=77
rlabel pdiffusion 234 -202 234 -202 0 feedthrough
rlabel pdiffusion 241 -202 241 -202 0 feedthrough
rlabel pdiffusion 248 -202 248 -202 0 cellNo=839
rlabel pdiffusion 255 -202 255 -202 0 feedthrough
rlabel pdiffusion 262 -202 262 -202 0 cellNo=16
rlabel pdiffusion 269 -202 269 -202 0 feedthrough
rlabel pdiffusion 276 -202 276 -202 0 feedthrough
rlabel pdiffusion 283 -202 283 -202 0 cellNo=579
rlabel pdiffusion 290 -202 290 -202 0 feedthrough
rlabel pdiffusion 297 -202 297 -202 0 feedthrough
rlabel pdiffusion 304 -202 304 -202 0 cellNo=628
rlabel pdiffusion 311 -202 311 -202 0 feedthrough
rlabel pdiffusion 318 -202 318 -202 0 feedthrough
rlabel pdiffusion 325 -202 325 -202 0 feedthrough
rlabel pdiffusion 332 -202 332 -202 0 feedthrough
rlabel pdiffusion 339 -202 339 -202 0 feedthrough
rlabel pdiffusion 346 -202 346 -202 0 feedthrough
rlabel pdiffusion 353 -202 353 -202 0 feedthrough
rlabel pdiffusion 360 -202 360 -202 0 feedthrough
rlabel pdiffusion 367 -202 367 -202 0 cellNo=183
rlabel pdiffusion 374 -202 374 -202 0 feedthrough
rlabel pdiffusion 381 -202 381 -202 0 cellNo=67
rlabel pdiffusion 395 -202 395 -202 0 feedthrough
rlabel pdiffusion 402 -202 402 -202 0 cellNo=632
rlabel pdiffusion 409 -202 409 -202 0 feedthrough
rlabel pdiffusion 416 -202 416 -202 0 feedthrough
rlabel pdiffusion 423 -202 423 -202 0 cellNo=692
rlabel pdiffusion 430 -202 430 -202 0 cellNo=508
rlabel pdiffusion 437 -202 437 -202 0 feedthrough
rlabel pdiffusion 444 -202 444 -202 0 cellNo=237
rlabel pdiffusion 3 -235 3 -235 0 cellNo=342
rlabel pdiffusion 10 -235 10 -235 0 cellNo=581
rlabel pdiffusion 17 -235 17 -235 0 cellNo=474
rlabel pdiffusion 24 -235 24 -235 0 cellNo=673
rlabel pdiffusion 31 -235 31 -235 0 cellNo=895
rlabel pdiffusion 66 -235 66 -235 0 cellNo=785
rlabel pdiffusion 73 -235 73 -235 0 cellNo=52
rlabel pdiffusion 80 -235 80 -235 0 feedthrough
rlabel pdiffusion 87 -235 87 -235 0 feedthrough
rlabel pdiffusion 94 -235 94 -235 0 feedthrough
rlabel pdiffusion 101 -235 101 -235 0 feedthrough
rlabel pdiffusion 108 -235 108 -235 0 feedthrough
rlabel pdiffusion 115 -235 115 -235 0 feedthrough
rlabel pdiffusion 122 -235 122 -235 0 feedthrough
rlabel pdiffusion 129 -235 129 -235 0 feedthrough
rlabel pdiffusion 136 -235 136 -235 0 cellNo=395
rlabel pdiffusion 143 -235 143 -235 0 feedthrough
rlabel pdiffusion 150 -235 150 -235 0 cellNo=573
rlabel pdiffusion 157 -235 157 -235 0 cellNo=344
rlabel pdiffusion 164 -235 164 -235 0 cellNo=238
rlabel pdiffusion 171 -235 171 -235 0 feedthrough
rlabel pdiffusion 178 -235 178 -235 0 cellNo=794
rlabel pdiffusion 185 -235 185 -235 0 cellNo=643
rlabel pdiffusion 192 -235 192 -235 0 feedthrough
rlabel pdiffusion 199 -235 199 -235 0 cellNo=137
rlabel pdiffusion 206 -235 206 -235 0 cellNo=486
rlabel pdiffusion 213 -235 213 -235 0 feedthrough
rlabel pdiffusion 220 -235 220 -235 0 cellNo=689
rlabel pdiffusion 227 -235 227 -235 0 cellNo=466
rlabel pdiffusion 234 -235 234 -235 0 cellNo=48
rlabel pdiffusion 241 -235 241 -235 0 cellNo=726
rlabel pdiffusion 248 -235 248 -235 0 cellNo=39
rlabel pdiffusion 255 -235 255 -235 0 cellNo=800
rlabel pdiffusion 262 -235 262 -235 0 cellNo=8
rlabel pdiffusion 269 -235 269 -235 0 feedthrough
rlabel pdiffusion 276 -235 276 -235 0 feedthrough
rlabel pdiffusion 283 -235 283 -235 0 feedthrough
rlabel pdiffusion 290 -235 290 -235 0 feedthrough
rlabel pdiffusion 297 -235 297 -235 0 feedthrough
rlabel pdiffusion 304 -235 304 -235 0 feedthrough
rlabel pdiffusion 311 -235 311 -235 0 feedthrough
rlabel pdiffusion 318 -235 318 -235 0 feedthrough
rlabel pdiffusion 325 -235 325 -235 0 cellNo=638
rlabel pdiffusion 332 -235 332 -235 0 feedthrough
rlabel pdiffusion 339 -235 339 -235 0 feedthrough
rlabel pdiffusion 346 -235 346 -235 0 feedthrough
rlabel pdiffusion 353 -235 353 -235 0 feedthrough
rlabel pdiffusion 360 -235 360 -235 0 feedthrough
rlabel pdiffusion 367 -235 367 -235 0 cellNo=274
rlabel pdiffusion 374 -235 374 -235 0 feedthrough
rlabel pdiffusion 381 -235 381 -235 0 cellNo=568
rlabel pdiffusion 388 -235 388 -235 0 feedthrough
rlabel pdiffusion 416 -235 416 -235 0 cellNo=380
rlabel pdiffusion 423 -235 423 -235 0 feedthrough
rlabel pdiffusion 437 -235 437 -235 0 cellNo=710
rlabel pdiffusion 3 -278 3 -278 0 cellNo=399
rlabel pdiffusion 10 -278 10 -278 0 cellNo=470
rlabel pdiffusion 17 -278 17 -278 0 cellNo=670
rlabel pdiffusion 24 -278 24 -278 0 cellNo=830
rlabel pdiffusion 31 -278 31 -278 0 cellNo=371
rlabel pdiffusion 38 -278 38 -278 0 cellNo=709
rlabel pdiffusion 52 -278 52 -278 0 cellNo=577
rlabel pdiffusion 73 -278 73 -278 0 cellNo=191
rlabel pdiffusion 80 -278 80 -278 0 feedthrough
rlabel pdiffusion 87 -278 87 -278 0 cellNo=819
rlabel pdiffusion 94 -278 94 -278 0 feedthrough
rlabel pdiffusion 101 -278 101 -278 0 cellNo=668
rlabel pdiffusion 108 -278 108 -278 0 feedthrough
rlabel pdiffusion 115 -278 115 -278 0 feedthrough
rlabel pdiffusion 122 -278 122 -278 0 cellNo=513
rlabel pdiffusion 129 -278 129 -278 0 cellNo=576
rlabel pdiffusion 136 -278 136 -278 0 cellNo=161
rlabel pdiffusion 143 -278 143 -278 0 cellNo=341
rlabel pdiffusion 150 -278 150 -278 0 cellNo=621
rlabel pdiffusion 157 -278 157 -278 0 feedthrough
rlabel pdiffusion 164 -278 164 -278 0 feedthrough
rlabel pdiffusion 171 -278 171 -278 0 feedthrough
rlabel pdiffusion 178 -278 178 -278 0 feedthrough
rlabel pdiffusion 185 -278 185 -278 0 cellNo=484
rlabel pdiffusion 192 -278 192 -278 0 cellNo=487
rlabel pdiffusion 199 -278 199 -278 0 feedthrough
rlabel pdiffusion 206 -278 206 -278 0 cellNo=136
rlabel pdiffusion 213 -278 213 -278 0 cellNo=882
rlabel pdiffusion 220 -278 220 -278 0 cellNo=525
rlabel pdiffusion 227 -278 227 -278 0 cellNo=500
rlabel pdiffusion 234 -278 234 -278 0 feedthrough
rlabel pdiffusion 241 -278 241 -278 0 feedthrough
rlabel pdiffusion 248 -278 248 -278 0 feedthrough
rlabel pdiffusion 255 -278 255 -278 0 cellNo=71
rlabel pdiffusion 262 -278 262 -278 0 feedthrough
rlabel pdiffusion 269 -278 269 -278 0 cellNo=185
rlabel pdiffusion 276 -278 276 -278 0 feedthrough
rlabel pdiffusion 283 -278 283 -278 0 feedthrough
rlabel pdiffusion 290 -278 290 -278 0 cellNo=810
rlabel pdiffusion 297 -278 297 -278 0 cellNo=437
rlabel pdiffusion 304 -278 304 -278 0 cellNo=539
rlabel pdiffusion 311 -278 311 -278 0 feedthrough
rlabel pdiffusion 318 -278 318 -278 0 feedthrough
rlabel pdiffusion 325 -278 325 -278 0 feedthrough
rlabel pdiffusion 332 -278 332 -278 0 feedthrough
rlabel pdiffusion 339 -278 339 -278 0 feedthrough
rlabel pdiffusion 346 -278 346 -278 0 feedthrough
rlabel pdiffusion 353 -278 353 -278 0 feedthrough
rlabel pdiffusion 360 -278 360 -278 0 feedthrough
rlabel pdiffusion 367 -278 367 -278 0 feedthrough
rlabel pdiffusion 374 -278 374 -278 0 feedthrough
rlabel pdiffusion 381 -278 381 -278 0 feedthrough
rlabel pdiffusion 388 -278 388 -278 0 feedthrough
rlabel pdiffusion 395 -278 395 -278 0 feedthrough
rlabel pdiffusion 402 -278 402 -278 0 feedthrough
rlabel pdiffusion 409 -278 409 -278 0 feedthrough
rlabel pdiffusion 416 -278 416 -278 0 cellNo=422
rlabel pdiffusion 423 -278 423 -278 0 feedthrough
rlabel pdiffusion 430 -278 430 -278 0 feedthrough
rlabel pdiffusion 437 -278 437 -278 0 cellNo=103
rlabel pdiffusion 444 -278 444 -278 0 feedthrough
rlabel pdiffusion 451 -278 451 -278 0 cellNo=412
rlabel pdiffusion 458 -278 458 -278 0 feedthrough
rlabel pdiffusion 528 -278 528 -278 0 cellNo=258
rlabel pdiffusion 535 -278 535 -278 0 feedthrough
rlabel pdiffusion 3 -319 3 -319 0 cellNo=438
rlabel pdiffusion 10 -319 10 -319 0 cellNo=662
rlabel pdiffusion 17 -319 17 -319 0 cellNo=827
rlabel pdiffusion 31 -319 31 -319 0 cellNo=378
rlabel pdiffusion 45 -319 45 -319 0 cellNo=72
rlabel pdiffusion 52 -319 52 -319 0 cellNo=392
rlabel pdiffusion 59 -319 59 -319 0 feedthrough
rlabel pdiffusion 66 -319 66 -319 0 cellNo=624
rlabel pdiffusion 73 -319 73 -319 0 cellNo=350
rlabel pdiffusion 80 -319 80 -319 0 cellNo=92
rlabel pdiffusion 87 -319 87 -319 0 feedthrough
rlabel pdiffusion 94 -319 94 -319 0 feedthrough
rlabel pdiffusion 101 -319 101 -319 0 feedthrough
rlabel pdiffusion 108 -319 108 -319 0 cellNo=182
rlabel pdiffusion 115 -319 115 -319 0 feedthrough
rlabel pdiffusion 122 -319 122 -319 0 feedthrough
rlabel pdiffusion 129 -319 129 -319 0 feedthrough
rlabel pdiffusion 136 -319 136 -319 0 feedthrough
rlabel pdiffusion 143 -319 143 -319 0 cellNo=313
rlabel pdiffusion 150 -319 150 -319 0 cellNo=138
rlabel pdiffusion 157 -319 157 -319 0 cellNo=42
rlabel pdiffusion 164 -319 164 -319 0 feedthrough
rlabel pdiffusion 171 -319 171 -319 0 cellNo=236
rlabel pdiffusion 178 -319 178 -319 0 feedthrough
rlabel pdiffusion 185 -319 185 -319 0 feedthrough
rlabel pdiffusion 192 -319 192 -319 0 cellNo=58
rlabel pdiffusion 199 -319 199 -319 0 feedthrough
rlabel pdiffusion 206 -319 206 -319 0 cellNo=664
rlabel pdiffusion 213 -319 213 -319 0 feedthrough
rlabel pdiffusion 220 -319 220 -319 0 feedthrough
rlabel pdiffusion 227 -319 227 -319 0 cellNo=203
rlabel pdiffusion 234 -319 234 -319 0 feedthrough
rlabel pdiffusion 241 -319 241 -319 0 cellNo=658
rlabel pdiffusion 248 -319 248 -319 0 cellNo=154
rlabel pdiffusion 255 -319 255 -319 0 cellNo=384
rlabel pdiffusion 262 -319 262 -319 0 cellNo=283
rlabel pdiffusion 269 -319 269 -319 0 feedthrough
rlabel pdiffusion 276 -319 276 -319 0 feedthrough
rlabel pdiffusion 283 -319 283 -319 0 cellNo=667
rlabel pdiffusion 290 -319 290 -319 0 feedthrough
rlabel pdiffusion 297 -319 297 -319 0 cellNo=574
rlabel pdiffusion 304 -319 304 -319 0 feedthrough
rlabel pdiffusion 311 -319 311 -319 0 feedthrough
rlabel pdiffusion 318 -319 318 -319 0 feedthrough
rlabel pdiffusion 325 -319 325 -319 0 cellNo=680
rlabel pdiffusion 332 -319 332 -319 0 feedthrough
rlabel pdiffusion 339 -319 339 -319 0 feedthrough
rlabel pdiffusion 346 -319 346 -319 0 feedthrough
rlabel pdiffusion 353 -319 353 -319 0 feedthrough
rlabel pdiffusion 360 -319 360 -319 0 feedthrough
rlabel pdiffusion 367 -319 367 -319 0 feedthrough
rlabel pdiffusion 374 -319 374 -319 0 cellNo=331
rlabel pdiffusion 381 -319 381 -319 0 feedthrough
rlabel pdiffusion 388 -319 388 -319 0 feedthrough
rlabel pdiffusion 395 -319 395 -319 0 feedthrough
rlabel pdiffusion 402 -319 402 -319 0 feedthrough
rlabel pdiffusion 409 -319 409 -319 0 feedthrough
rlabel pdiffusion 416 -319 416 -319 0 cellNo=312
rlabel pdiffusion 423 -319 423 -319 0 feedthrough
rlabel pdiffusion 430 -319 430 -319 0 cellNo=397
rlabel pdiffusion 437 -319 437 -319 0 feedthrough
rlabel pdiffusion 451 -319 451 -319 0 cellNo=271
rlabel pdiffusion 521 -319 521 -319 0 cellNo=623
rlabel pdiffusion 528 -319 528 -319 0 feedthrough
rlabel pdiffusion 3 -366 3 -366 0 cellNo=657
rlabel pdiffusion 10 -366 10 -366 0 cellNo=825
rlabel pdiffusion 17 -366 17 -366 0 cellNo=774
rlabel pdiffusion 24 -366 24 -366 0 cellNo=566
rlabel pdiffusion 31 -366 31 -366 0 cellNo=403
rlabel pdiffusion 38 -366 38 -366 0 feedthrough
rlabel pdiffusion 45 -366 45 -366 0 feedthrough
rlabel pdiffusion 52 -366 52 -366 0 feedthrough
rlabel pdiffusion 59 -366 59 -366 0 feedthrough
rlabel pdiffusion 66 -366 66 -366 0 feedthrough
rlabel pdiffusion 73 -366 73 -366 0 feedthrough
rlabel pdiffusion 80 -366 80 -366 0 cellNo=708
rlabel pdiffusion 87 -366 87 -366 0 cellNo=565
rlabel pdiffusion 94 -366 94 -366 0 cellNo=428
rlabel pdiffusion 101 -366 101 -366 0 feedthrough
rlabel pdiffusion 108 -366 108 -366 0 cellNo=899
rlabel pdiffusion 115 -366 115 -366 0 cellNo=383
rlabel pdiffusion 122 -366 122 -366 0 cellNo=352
rlabel pdiffusion 129 -366 129 -366 0 cellNo=421
rlabel pdiffusion 136 -366 136 -366 0 cellNo=461
rlabel pdiffusion 143 -366 143 -366 0 cellNo=181
rlabel pdiffusion 150 -366 150 -366 0 feedthrough
rlabel pdiffusion 157 -366 157 -366 0 feedthrough
rlabel pdiffusion 164 -366 164 -366 0 cellNo=189
rlabel pdiffusion 171 -366 171 -366 0 cellNo=319
rlabel pdiffusion 178 -366 178 -366 0 feedthrough
rlabel pdiffusion 185 -366 185 -366 0 feedthrough
rlabel pdiffusion 192 -366 192 -366 0 cellNo=76
rlabel pdiffusion 199 -366 199 -366 0 cellNo=631
rlabel pdiffusion 206 -366 206 -366 0 feedthrough
rlabel pdiffusion 213 -366 213 -366 0 cellNo=552
rlabel pdiffusion 220 -366 220 -366 0 feedthrough
rlabel pdiffusion 227 -366 227 -366 0 feedthrough
rlabel pdiffusion 234 -366 234 -366 0 feedthrough
rlabel pdiffusion 241 -366 241 -366 0 cellNo=445
rlabel pdiffusion 248 -366 248 -366 0 cellNo=540
rlabel pdiffusion 255 -366 255 -366 0 cellNo=324
rlabel pdiffusion 262 -366 262 -366 0 cellNo=716
rlabel pdiffusion 269 -366 269 -366 0 cellNo=655
rlabel pdiffusion 276 -366 276 -366 0 cellNo=158
rlabel pdiffusion 283 -366 283 -366 0 cellNo=231
rlabel pdiffusion 290 -366 290 -366 0 feedthrough
rlabel pdiffusion 297 -366 297 -366 0 feedthrough
rlabel pdiffusion 304 -366 304 -366 0 cellNo=762
rlabel pdiffusion 311 -366 311 -366 0 feedthrough
rlabel pdiffusion 318 -366 318 -366 0 cellNo=596
rlabel pdiffusion 325 -366 325 -366 0 cellNo=162
rlabel pdiffusion 332 -366 332 -366 0 feedthrough
rlabel pdiffusion 339 -366 339 -366 0 feedthrough
rlabel pdiffusion 346 -366 346 -366 0 feedthrough
rlabel pdiffusion 353 -366 353 -366 0 feedthrough
rlabel pdiffusion 360 -366 360 -366 0 feedthrough
rlabel pdiffusion 367 -366 367 -366 0 feedthrough
rlabel pdiffusion 374 -366 374 -366 0 feedthrough
rlabel pdiffusion 381 -366 381 -366 0 feedthrough
rlabel pdiffusion 388 -366 388 -366 0 cellNo=286
rlabel pdiffusion 395 -366 395 -366 0 feedthrough
rlabel pdiffusion 402 -366 402 -366 0 feedthrough
rlabel pdiffusion 409 -366 409 -366 0 feedthrough
rlabel pdiffusion 416 -366 416 -366 0 feedthrough
rlabel pdiffusion 423 -366 423 -366 0 feedthrough
rlabel pdiffusion 430 -366 430 -366 0 feedthrough
rlabel pdiffusion 437 -366 437 -366 0 feedthrough
rlabel pdiffusion 444 -366 444 -366 0 feedthrough
rlabel pdiffusion 451 -366 451 -366 0 feedthrough
rlabel pdiffusion 458 -366 458 -366 0 feedthrough
rlabel pdiffusion 465 -366 465 -366 0 cellNo=609
rlabel pdiffusion 472 -366 472 -366 0 feedthrough
rlabel pdiffusion 514 -366 514 -366 0 feedthrough
rlabel pdiffusion 3 -417 3 -417 0 cellNo=818
rlabel pdiffusion 17 -417 17 -417 0 cellNo=431
rlabel pdiffusion 24 -417 24 -417 0 feedthrough
rlabel pdiffusion 31 -417 31 -417 0 feedthrough
rlabel pdiffusion 38 -417 38 -417 0 cellNo=447
rlabel pdiffusion 45 -417 45 -417 0 cellNo=302
rlabel pdiffusion 52 -417 52 -417 0 cellNo=64
rlabel pdiffusion 59 -417 59 -417 0 cellNo=251
rlabel pdiffusion 66 -417 66 -417 0 cellNo=420
rlabel pdiffusion 73 -417 73 -417 0 feedthrough
rlabel pdiffusion 80 -417 80 -417 0 feedthrough
rlabel pdiffusion 87 -417 87 -417 0 feedthrough
rlabel pdiffusion 94 -417 94 -417 0 feedthrough
rlabel pdiffusion 101 -417 101 -417 0 cellNo=496
rlabel pdiffusion 108 -417 108 -417 0 cellNo=841
rlabel pdiffusion 115 -417 115 -417 0 feedthrough
rlabel pdiffusion 122 -417 122 -417 0 feedthrough
rlabel pdiffusion 129 -417 129 -417 0 feedthrough
rlabel pdiffusion 136 -417 136 -417 0 cellNo=346
rlabel pdiffusion 143 -417 143 -417 0 cellNo=543
rlabel pdiffusion 150 -417 150 -417 0 cellNo=24
rlabel pdiffusion 157 -417 157 -417 0 cellNo=220
rlabel pdiffusion 164 -417 164 -417 0 cellNo=448
rlabel pdiffusion 171 -417 171 -417 0 feedthrough
rlabel pdiffusion 178 -417 178 -417 0 feedthrough
rlabel pdiffusion 185 -417 185 -417 0 feedthrough
rlabel pdiffusion 192 -417 192 -417 0 cellNo=622
rlabel pdiffusion 199 -417 199 -417 0 feedthrough
rlabel pdiffusion 206 -417 206 -417 0 cellNo=328
rlabel pdiffusion 213 -417 213 -417 0 cellNo=767
rlabel pdiffusion 220 -417 220 -417 0 feedthrough
rlabel pdiffusion 227 -417 227 -417 0 cellNo=110
rlabel pdiffusion 234 -417 234 -417 0 feedthrough
rlabel pdiffusion 241 -417 241 -417 0 feedthrough
rlabel pdiffusion 248 -417 248 -417 0 feedthrough
rlabel pdiffusion 255 -417 255 -417 0 feedthrough
rlabel pdiffusion 262 -417 262 -417 0 cellNo=186
rlabel pdiffusion 269 -417 269 -417 0 cellNo=652
rlabel pdiffusion 276 -417 276 -417 0 feedthrough
rlabel pdiffusion 283 -417 283 -417 0 cellNo=11
rlabel pdiffusion 290 -417 290 -417 0 feedthrough
rlabel pdiffusion 297 -417 297 -417 0 feedthrough
rlabel pdiffusion 304 -417 304 -417 0 feedthrough
rlabel pdiffusion 311 -417 311 -417 0 cellNo=316
rlabel pdiffusion 318 -417 318 -417 0 cellNo=160
rlabel pdiffusion 325 -417 325 -417 0 cellNo=124
rlabel pdiffusion 332 -417 332 -417 0 feedthrough
rlabel pdiffusion 339 -417 339 -417 0 cellNo=719
rlabel pdiffusion 346 -417 346 -417 0 cellNo=131
rlabel pdiffusion 353 -417 353 -417 0 feedthrough
rlabel pdiffusion 360 -417 360 -417 0 feedthrough
rlabel pdiffusion 367 -417 367 -417 0 feedthrough
rlabel pdiffusion 374 -417 374 -417 0 feedthrough
rlabel pdiffusion 381 -417 381 -417 0 feedthrough
rlabel pdiffusion 388 -417 388 -417 0 feedthrough
rlabel pdiffusion 395 -417 395 -417 0 feedthrough
rlabel pdiffusion 402 -417 402 -417 0 feedthrough
rlabel pdiffusion 409 -417 409 -417 0 feedthrough
rlabel pdiffusion 416 -417 416 -417 0 cellNo=851
rlabel pdiffusion 423 -417 423 -417 0 feedthrough
rlabel pdiffusion 430 -417 430 -417 0 feedthrough
rlabel pdiffusion 437 -417 437 -417 0 feedthrough
rlabel pdiffusion 444 -417 444 -417 0 feedthrough
rlabel pdiffusion 451 -417 451 -417 0 feedthrough
rlabel pdiffusion 458 -417 458 -417 0 feedthrough
rlabel pdiffusion 465 -417 465 -417 0 feedthrough
rlabel pdiffusion 472 -417 472 -417 0 feedthrough
rlabel pdiffusion 479 -417 479 -417 0 cellNo=368
rlabel pdiffusion 486 -417 486 -417 0 cellNo=760
rlabel pdiffusion 493 -417 493 -417 0 feedthrough
rlabel pdiffusion 500 -417 500 -417 0 feedthrough
rlabel pdiffusion 507 -417 507 -417 0 cellNo=535
rlabel pdiffusion 514 -417 514 -417 0 feedthrough
rlabel pdiffusion 521 -417 521 -417 0 feedthrough
rlabel pdiffusion 528 -417 528 -417 0 feedthrough
rlabel pdiffusion 3 -468 3 -468 0 feedthrough
rlabel pdiffusion 10 -468 10 -468 0 feedthrough
rlabel pdiffusion 17 -468 17 -468 0 feedthrough
rlabel pdiffusion 24 -468 24 -468 0 cellNo=502
rlabel pdiffusion 31 -468 31 -468 0 cellNo=105
rlabel pdiffusion 38 -468 38 -468 0 feedthrough
rlabel pdiffusion 45 -468 45 -468 0 feedthrough
rlabel pdiffusion 52 -468 52 -468 0 cellNo=69
rlabel pdiffusion 59 -468 59 -468 0 feedthrough
rlabel pdiffusion 66 -468 66 -468 0 feedthrough
rlabel pdiffusion 73 -468 73 -468 0 feedthrough
rlabel pdiffusion 80 -468 80 -468 0 feedthrough
rlabel pdiffusion 87 -468 87 -468 0 feedthrough
rlabel pdiffusion 94 -468 94 -468 0 cellNo=788
rlabel pdiffusion 101 -468 101 -468 0 feedthrough
rlabel pdiffusion 108 -468 108 -468 0 feedthrough
rlabel pdiffusion 115 -468 115 -468 0 cellNo=518
rlabel pdiffusion 122 -468 122 -468 0 cellNo=603
rlabel pdiffusion 129 -468 129 -468 0 cellNo=456
rlabel pdiffusion 136 -468 136 -468 0 feedthrough
rlabel pdiffusion 143 -468 143 -468 0 feedthrough
rlabel pdiffusion 150 -468 150 -468 0 cellNo=44
rlabel pdiffusion 157 -468 157 -468 0 cellNo=334
rlabel pdiffusion 164 -468 164 -468 0 cellNo=489
rlabel pdiffusion 171 -468 171 -468 0 cellNo=572
rlabel pdiffusion 178 -468 178 -468 0 feedthrough
rlabel pdiffusion 185 -468 185 -468 0 feedthrough
rlabel pdiffusion 192 -468 192 -468 0 cellNo=682
rlabel pdiffusion 199 -468 199 -468 0 cellNo=65
rlabel pdiffusion 206 -468 206 -468 0 feedthrough
rlabel pdiffusion 213 -468 213 -468 0 feedthrough
rlabel pdiffusion 220 -468 220 -468 0 cellNo=355
rlabel pdiffusion 227 -468 227 -468 0 cellNo=531
rlabel pdiffusion 234 -468 234 -468 0 feedthrough
rlabel pdiffusion 241 -468 241 -468 0 cellNo=152
rlabel pdiffusion 248 -468 248 -468 0 feedthrough
rlabel pdiffusion 255 -468 255 -468 0 cellNo=118
rlabel pdiffusion 262 -468 262 -468 0 cellNo=738
rlabel pdiffusion 269 -468 269 -468 0 feedthrough
rlabel pdiffusion 276 -468 276 -468 0 cellNo=55
rlabel pdiffusion 283 -468 283 -468 0 cellNo=100
rlabel pdiffusion 290 -468 290 -468 0 feedthrough
rlabel pdiffusion 297 -468 297 -468 0 feedthrough
rlabel pdiffusion 304 -468 304 -468 0 feedthrough
rlabel pdiffusion 311 -468 311 -468 0 cellNo=522
rlabel pdiffusion 318 -468 318 -468 0 cellNo=78
rlabel pdiffusion 325 -468 325 -468 0 feedthrough
rlabel pdiffusion 332 -468 332 -468 0 feedthrough
rlabel pdiffusion 339 -468 339 -468 0 feedthrough
rlabel pdiffusion 346 -468 346 -468 0 cellNo=847
rlabel pdiffusion 353 -468 353 -468 0 cellNo=791
rlabel pdiffusion 360 -468 360 -468 0 cellNo=594
rlabel pdiffusion 367 -468 367 -468 0 cellNo=544
rlabel pdiffusion 374 -468 374 -468 0 cellNo=757
rlabel pdiffusion 381 -468 381 -468 0 feedthrough
rlabel pdiffusion 388 -468 388 -468 0 feedthrough
rlabel pdiffusion 395 -468 395 -468 0 feedthrough
rlabel pdiffusion 402 -468 402 -468 0 feedthrough
rlabel pdiffusion 409 -468 409 -468 0 feedthrough
rlabel pdiffusion 416 -468 416 -468 0 feedthrough
rlabel pdiffusion 423 -468 423 -468 0 feedthrough
rlabel pdiffusion 430 -468 430 -468 0 feedthrough
rlabel pdiffusion 437 -468 437 -468 0 feedthrough
rlabel pdiffusion 444 -468 444 -468 0 feedthrough
rlabel pdiffusion 451 -468 451 -468 0 feedthrough
rlabel pdiffusion 458 -468 458 -468 0 feedthrough
rlabel pdiffusion 465 -468 465 -468 0 feedthrough
rlabel pdiffusion 472 -468 472 -468 0 feedthrough
rlabel pdiffusion 479 -468 479 -468 0 feedthrough
rlabel pdiffusion 486 -468 486 -468 0 feedthrough
rlabel pdiffusion 493 -468 493 -468 0 feedthrough
rlabel pdiffusion 500 -468 500 -468 0 feedthrough
rlabel pdiffusion 507 -468 507 -468 0 feedthrough
rlabel pdiffusion 514 -468 514 -468 0 feedthrough
rlabel pdiffusion 521 -468 521 -468 0 feedthrough
rlabel pdiffusion 528 -468 528 -468 0 feedthrough
rlabel pdiffusion 535 -468 535 -468 0 feedthrough
rlabel pdiffusion 542 -468 542 -468 0 feedthrough
rlabel pdiffusion 549 -468 549 -468 0 feedthrough
rlabel pdiffusion 556 -468 556 -468 0 cellNo=862
rlabel pdiffusion 563 -468 563 -468 0 feedthrough
rlabel pdiffusion 570 -468 570 -468 0 cellNo=608
rlabel pdiffusion 577 -468 577 -468 0 feedthrough
rlabel pdiffusion 17 -525 17 -525 0 feedthrough
rlabel pdiffusion 24 -525 24 -525 0 feedthrough
rlabel pdiffusion 31 -525 31 -525 0 feedthrough
rlabel pdiffusion 38 -525 38 -525 0 feedthrough
rlabel pdiffusion 45 -525 45 -525 0 feedthrough
rlabel pdiffusion 52 -525 52 -525 0 feedthrough
rlabel pdiffusion 59 -525 59 -525 0 feedthrough
rlabel pdiffusion 66 -525 66 -525 0 cellNo=848
rlabel pdiffusion 73 -525 73 -525 0 cellNo=806
rlabel pdiffusion 80 -525 80 -525 0 cellNo=269
rlabel pdiffusion 87 -525 87 -525 0 cellNo=600
rlabel pdiffusion 94 -525 94 -525 0 feedthrough
rlabel pdiffusion 101 -525 101 -525 0 feedthrough
rlabel pdiffusion 108 -525 108 -525 0 feedthrough
rlabel pdiffusion 115 -525 115 -525 0 cellNo=824
rlabel pdiffusion 122 -525 122 -525 0 cellNo=555
rlabel pdiffusion 129 -525 129 -525 0 cellNo=2
rlabel pdiffusion 136 -525 136 -525 0 cellNo=298
rlabel pdiffusion 143 -525 143 -525 0 cellNo=460
rlabel pdiffusion 150 -525 150 -525 0 feedthrough
rlabel pdiffusion 157 -525 157 -525 0 cellNo=450
rlabel pdiffusion 164 -525 164 -525 0 feedthrough
rlabel pdiffusion 171 -525 171 -525 0 feedthrough
rlabel pdiffusion 178 -525 178 -525 0 feedthrough
rlabel pdiffusion 185 -525 185 -525 0 cellNo=755
rlabel pdiffusion 192 -525 192 -525 0 feedthrough
rlabel pdiffusion 199 -525 199 -525 0 cellNo=382
rlabel pdiffusion 206 -525 206 -525 0 feedthrough
rlabel pdiffusion 213 -525 213 -525 0 feedthrough
rlabel pdiffusion 220 -525 220 -525 0 cellNo=234
rlabel pdiffusion 227 -525 227 -525 0 cellNo=227
rlabel pdiffusion 234 -525 234 -525 0 feedthrough
rlabel pdiffusion 241 -525 241 -525 0 cellNo=309
rlabel pdiffusion 248 -525 248 -525 0 feedthrough
rlabel pdiffusion 255 -525 255 -525 0 feedthrough
rlabel pdiffusion 262 -525 262 -525 0 cellNo=411
rlabel pdiffusion 269 -525 269 -525 0 feedthrough
rlabel pdiffusion 276 -525 276 -525 0 cellNo=57
rlabel pdiffusion 283 -525 283 -525 0 cellNo=279
rlabel pdiffusion 290 -525 290 -525 0 cellNo=253
rlabel pdiffusion 297 -525 297 -525 0 cellNo=465
rlabel pdiffusion 304 -525 304 -525 0 feedthrough
rlabel pdiffusion 311 -525 311 -525 0 cellNo=506
rlabel pdiffusion 318 -525 318 -525 0 feedthrough
rlabel pdiffusion 325 -525 325 -525 0 cellNo=546
rlabel pdiffusion 332 -525 332 -525 0 feedthrough
rlabel pdiffusion 339 -525 339 -525 0 feedthrough
rlabel pdiffusion 346 -525 346 -525 0 cellNo=782
rlabel pdiffusion 353 -525 353 -525 0 cellNo=106
rlabel pdiffusion 360 -525 360 -525 0 feedthrough
rlabel pdiffusion 367 -525 367 -525 0 cellNo=497
rlabel pdiffusion 374 -525 374 -525 0 cellNo=557
rlabel pdiffusion 381 -525 381 -525 0 feedthrough
rlabel pdiffusion 388 -525 388 -525 0 cellNo=892
rlabel pdiffusion 395 -525 395 -525 0 feedthrough
rlabel pdiffusion 402 -525 402 -525 0 feedthrough
rlabel pdiffusion 409 -525 409 -525 0 feedthrough
rlabel pdiffusion 416 -525 416 -525 0 feedthrough
rlabel pdiffusion 423 -525 423 -525 0 cellNo=318
rlabel pdiffusion 430 -525 430 -525 0 feedthrough
rlabel pdiffusion 437 -525 437 -525 0 feedthrough
rlabel pdiffusion 444 -525 444 -525 0 feedthrough
rlabel pdiffusion 451 -525 451 -525 0 feedthrough
rlabel pdiffusion 458 -525 458 -525 0 feedthrough
rlabel pdiffusion 465 -525 465 -525 0 feedthrough
rlabel pdiffusion 472 -525 472 -525 0 feedthrough
rlabel pdiffusion 479 -525 479 -525 0 feedthrough
rlabel pdiffusion 486 -525 486 -525 0 feedthrough
rlabel pdiffusion 493 -525 493 -525 0 feedthrough
rlabel pdiffusion 500 -525 500 -525 0 feedthrough
rlabel pdiffusion 507 -525 507 -525 0 cellNo=314
rlabel pdiffusion 514 -525 514 -525 0 cellNo=620
rlabel pdiffusion 521 -525 521 -525 0 feedthrough
rlabel pdiffusion 542 -525 542 -525 0 feedthrough
rlabel pdiffusion 563 -525 563 -525 0 feedthrough
rlabel pdiffusion 10 -574 10 -574 0 feedthrough
rlabel pdiffusion 17 -574 17 -574 0 cellNo=736
rlabel pdiffusion 24 -574 24 -574 0 cellNo=247
rlabel pdiffusion 31 -574 31 -574 0 feedthrough
rlabel pdiffusion 38 -574 38 -574 0 cellNo=691
rlabel pdiffusion 45 -574 45 -574 0 cellNo=464
rlabel pdiffusion 52 -574 52 -574 0 feedthrough
rlabel pdiffusion 59 -574 59 -574 0 cellNo=423
rlabel pdiffusion 66 -574 66 -574 0 cellNo=387
rlabel pdiffusion 73 -574 73 -574 0 feedthrough
rlabel pdiffusion 80 -574 80 -574 0 feedthrough
rlabel pdiffusion 87 -574 87 -574 0 cellNo=153
rlabel pdiffusion 94 -574 94 -574 0 feedthrough
rlabel pdiffusion 101 -574 101 -574 0 cellNo=656
rlabel pdiffusion 108 -574 108 -574 0 cellNo=599
rlabel pdiffusion 115 -574 115 -574 0 cellNo=612
rlabel pdiffusion 122 -574 122 -574 0 feedthrough
rlabel pdiffusion 129 -574 129 -574 0 feedthrough
rlabel pdiffusion 136 -574 136 -574 0 feedthrough
rlabel pdiffusion 143 -574 143 -574 0 feedthrough
rlabel pdiffusion 150 -574 150 -574 0 feedthrough
rlabel pdiffusion 157 -574 157 -574 0 feedthrough
rlabel pdiffusion 164 -574 164 -574 0 feedthrough
rlabel pdiffusion 171 -574 171 -574 0 cellNo=163
rlabel pdiffusion 178 -574 178 -574 0 feedthrough
rlabel pdiffusion 185 -574 185 -574 0 cellNo=511
rlabel pdiffusion 192 -574 192 -574 0 feedthrough
rlabel pdiffusion 199 -574 199 -574 0 feedthrough
rlabel pdiffusion 206 -574 206 -574 0 cellNo=307
rlabel pdiffusion 213 -574 213 -574 0 cellNo=527
rlabel pdiffusion 220 -574 220 -574 0 cellNo=115
rlabel pdiffusion 227 -574 227 -574 0 cellNo=38
rlabel pdiffusion 234 -574 234 -574 0 cellNo=114
rlabel pdiffusion 241 -574 241 -574 0 cellNo=418
rlabel pdiffusion 248 -574 248 -574 0 feedthrough
rlabel pdiffusion 255 -574 255 -574 0 cellNo=405
rlabel pdiffusion 262 -574 262 -574 0 feedthrough
rlabel pdiffusion 269 -574 269 -574 0 cellNo=173
rlabel pdiffusion 276 -574 276 -574 0 feedthrough
rlabel pdiffusion 283 -574 283 -574 0 cellNo=139
rlabel pdiffusion 290 -574 290 -574 0 feedthrough
rlabel pdiffusion 297 -574 297 -574 0 feedthrough
rlabel pdiffusion 304 -574 304 -574 0 cellNo=89
rlabel pdiffusion 311 -574 311 -574 0 cellNo=859
rlabel pdiffusion 318 -574 318 -574 0 feedthrough
rlabel pdiffusion 325 -574 325 -574 0 feedthrough
rlabel pdiffusion 332 -574 332 -574 0 feedthrough
rlabel pdiffusion 339 -574 339 -574 0 cellNo=514
rlabel pdiffusion 346 -574 346 -574 0 feedthrough
rlabel pdiffusion 353 -574 353 -574 0 feedthrough
rlabel pdiffusion 360 -574 360 -574 0 cellNo=754
rlabel pdiffusion 367 -574 367 -574 0 cellNo=393
rlabel pdiffusion 374 -574 374 -574 0 feedthrough
rlabel pdiffusion 381 -574 381 -574 0 feedthrough
rlabel pdiffusion 388 -574 388 -574 0 feedthrough
rlabel pdiffusion 395 -574 395 -574 0 feedthrough
rlabel pdiffusion 402 -574 402 -574 0 feedthrough
rlabel pdiffusion 409 -574 409 -574 0 feedthrough
rlabel pdiffusion 416 -574 416 -574 0 feedthrough
rlabel pdiffusion 423 -574 423 -574 0 feedthrough
rlabel pdiffusion 430 -574 430 -574 0 cellNo=590
rlabel pdiffusion 437 -574 437 -574 0 feedthrough
rlabel pdiffusion 444 -574 444 -574 0 feedthrough
rlabel pdiffusion 451 -574 451 -574 0 feedthrough
rlabel pdiffusion 458 -574 458 -574 0 feedthrough
rlabel pdiffusion 465 -574 465 -574 0 feedthrough
rlabel pdiffusion 472 -574 472 -574 0 feedthrough
rlabel pdiffusion 479 -574 479 -574 0 feedthrough
rlabel pdiffusion 486 -574 486 -574 0 feedthrough
rlabel pdiffusion 493 -574 493 -574 0 feedthrough
rlabel pdiffusion 500 -574 500 -574 0 cellNo=439
rlabel pdiffusion 507 -574 507 -574 0 feedthrough
rlabel pdiffusion 514 -574 514 -574 0 cellNo=773
rlabel pdiffusion 521 -574 521 -574 0 feedthrough
rlabel pdiffusion 528 -574 528 -574 0 cellNo=204
rlabel pdiffusion 535 -574 535 -574 0 feedthrough
rlabel pdiffusion 542 -574 542 -574 0 feedthrough
rlabel pdiffusion 549 -574 549 -574 0 cellNo=250
rlabel pdiffusion 556 -574 556 -574 0 feedthrough
rlabel pdiffusion 563 -574 563 -574 0 feedthrough
rlabel pdiffusion 10 -617 10 -617 0 feedthrough
rlabel pdiffusion 17 -617 17 -617 0 feedthrough
rlabel pdiffusion 24 -617 24 -617 0 feedthrough
rlabel pdiffusion 31 -617 31 -617 0 feedthrough
rlabel pdiffusion 38 -617 38 -617 0 feedthrough
rlabel pdiffusion 45 -617 45 -617 0 cellNo=375
rlabel pdiffusion 52 -617 52 -617 0 cellNo=214
rlabel pdiffusion 59 -617 59 -617 0 feedthrough
rlabel pdiffusion 66 -617 66 -617 0 cellNo=550
rlabel pdiffusion 73 -617 73 -617 0 feedthrough
rlabel pdiffusion 80 -617 80 -617 0 cellNo=442
rlabel pdiffusion 87 -617 87 -617 0 cellNo=374
rlabel pdiffusion 94 -617 94 -617 0 feedthrough
rlabel pdiffusion 101 -617 101 -617 0 cellNo=822
rlabel pdiffusion 108 -617 108 -617 0 feedthrough
rlabel pdiffusion 115 -617 115 -617 0 cellNo=230
rlabel pdiffusion 122 -617 122 -617 0 feedthrough
rlabel pdiffusion 129 -617 129 -617 0 cellNo=303
rlabel pdiffusion 136 -617 136 -617 0 cellNo=564
rlabel pdiffusion 143 -617 143 -617 0 cellNo=184
rlabel pdiffusion 150 -617 150 -617 0 feedthrough
rlabel pdiffusion 157 -617 157 -617 0 feedthrough
rlabel pdiffusion 164 -617 164 -617 0 feedthrough
rlabel pdiffusion 171 -617 171 -617 0 feedthrough
rlabel pdiffusion 178 -617 178 -617 0 cellNo=515
rlabel pdiffusion 185 -617 185 -617 0 cellNo=117
rlabel pdiffusion 192 -617 192 -617 0 feedthrough
rlabel pdiffusion 199 -617 199 -617 0 feedthrough
rlabel pdiffusion 206 -617 206 -617 0 feedthrough
rlabel pdiffusion 213 -617 213 -617 0 cellNo=805
rlabel pdiffusion 220 -617 220 -617 0 cellNo=95
rlabel pdiffusion 227 -617 227 -617 0 cellNo=323
rlabel pdiffusion 234 -617 234 -617 0 feedthrough
rlabel pdiffusion 241 -617 241 -617 0 feedthrough
rlabel pdiffusion 248 -617 248 -617 0 feedthrough
rlabel pdiffusion 255 -617 255 -617 0 feedthrough
rlabel pdiffusion 262 -617 262 -617 0 feedthrough
rlabel pdiffusion 269 -617 269 -617 0 feedthrough
rlabel pdiffusion 276 -617 276 -617 0 feedthrough
rlabel pdiffusion 283 -617 283 -617 0 feedthrough
rlabel pdiffusion 290 -617 290 -617 0 cellNo=98
rlabel pdiffusion 297 -617 297 -617 0 cellNo=223
rlabel pdiffusion 304 -617 304 -617 0 feedthrough
rlabel pdiffusion 311 -617 311 -617 0 cellNo=444
rlabel pdiffusion 318 -617 318 -617 0 feedthrough
rlabel pdiffusion 325 -617 325 -617 0 cellNo=777
rlabel pdiffusion 332 -617 332 -617 0 feedthrough
rlabel pdiffusion 339 -617 339 -617 0 cellNo=618
rlabel pdiffusion 346 -617 346 -617 0 feedthrough
rlabel pdiffusion 353 -617 353 -617 0 cellNo=83
rlabel pdiffusion 360 -617 360 -617 0 feedthrough
rlabel pdiffusion 367 -617 367 -617 0 feedthrough
rlabel pdiffusion 374 -617 374 -617 0 feedthrough
rlabel pdiffusion 381 -617 381 -617 0 feedthrough
rlabel pdiffusion 388 -617 388 -617 0 feedthrough
rlabel pdiffusion 395 -617 395 -617 0 cellNo=491
rlabel pdiffusion 402 -617 402 -617 0 feedthrough
rlabel pdiffusion 409 -617 409 -617 0 feedthrough
rlabel pdiffusion 416 -617 416 -617 0 cellNo=358
rlabel pdiffusion 423 -617 423 -617 0 feedthrough
rlabel pdiffusion 430 -617 430 -617 0 feedthrough
rlabel pdiffusion 437 -617 437 -617 0 feedthrough
rlabel pdiffusion 444 -617 444 -617 0 feedthrough
rlabel pdiffusion 451 -617 451 -617 0 feedthrough
rlabel pdiffusion 458 -617 458 -617 0 feedthrough
rlabel pdiffusion 465 -617 465 -617 0 feedthrough
rlabel pdiffusion 472 -617 472 -617 0 feedthrough
rlabel pdiffusion 479 -617 479 -617 0 cellNo=748
rlabel pdiffusion 486 -617 486 -617 0 feedthrough
rlabel pdiffusion 493 -617 493 -617 0 feedthrough
rlabel pdiffusion 500 -617 500 -617 0 feedthrough
rlabel pdiffusion 507 -617 507 -617 0 cellNo=459
rlabel pdiffusion 514 -617 514 -617 0 cellNo=665
rlabel pdiffusion 521 -617 521 -617 0 cellNo=74
rlabel pdiffusion 528 -617 528 -617 0 feedthrough
rlabel pdiffusion 535 -617 535 -617 0 feedthrough
rlabel pdiffusion 542 -617 542 -617 0 feedthrough
rlabel pdiffusion 549 -617 549 -617 0 feedthrough
rlabel pdiffusion 556 -617 556 -617 0 feedthrough
rlabel pdiffusion 563 -617 563 -617 0 cellNo=415
rlabel pdiffusion 38 -664 38 -664 0 cellNo=505
rlabel pdiffusion 45 -664 45 -664 0 feedthrough
rlabel pdiffusion 52 -664 52 -664 0 feedthrough
rlabel pdiffusion 59 -664 59 -664 0 cellNo=404
rlabel pdiffusion 66 -664 66 -664 0 feedthrough
rlabel pdiffusion 73 -664 73 -664 0 cellNo=356
rlabel pdiffusion 80 -664 80 -664 0 feedthrough
rlabel pdiffusion 87 -664 87 -664 0 feedthrough
rlabel pdiffusion 94 -664 94 -664 0 cellNo=21
rlabel pdiffusion 101 -664 101 -664 0 cellNo=856
rlabel pdiffusion 108 -664 108 -664 0 feedthrough
rlabel pdiffusion 115 -664 115 -664 0 cellNo=530
rlabel pdiffusion 122 -664 122 -664 0 feedthrough
rlabel pdiffusion 129 -664 129 -664 0 cellNo=634
rlabel pdiffusion 136 -664 136 -664 0 feedthrough
rlabel pdiffusion 143 -664 143 -664 0 cellNo=244
rlabel pdiffusion 150 -664 150 -664 0 feedthrough
rlabel pdiffusion 157 -664 157 -664 0 feedthrough
rlabel pdiffusion 164 -664 164 -664 0 feedthrough
rlabel pdiffusion 171 -664 171 -664 0 cellNo=175
rlabel pdiffusion 178 -664 178 -664 0 feedthrough
rlabel pdiffusion 185 -664 185 -664 0 feedthrough
rlabel pdiffusion 192 -664 192 -664 0 feedthrough
rlabel pdiffusion 199 -664 199 -664 0 cellNo=202
rlabel pdiffusion 206 -664 206 -664 0 cellNo=320
rlabel pdiffusion 213 -664 213 -664 0 feedthrough
rlabel pdiffusion 220 -664 220 -664 0 feedthrough
rlabel pdiffusion 227 -664 227 -664 0 feedthrough
rlabel pdiffusion 234 -664 234 -664 0 feedthrough
rlabel pdiffusion 241 -664 241 -664 0 cellNo=684
rlabel pdiffusion 248 -664 248 -664 0 cellNo=704
rlabel pdiffusion 255 -664 255 -664 0 feedthrough
rlabel pdiffusion 262 -664 262 -664 0 feedthrough
rlabel pdiffusion 269 -664 269 -664 0 cellNo=30
rlabel pdiffusion 276 -664 276 -664 0 feedthrough
rlabel pdiffusion 283 -664 283 -664 0 feedthrough
rlabel pdiffusion 290 -664 290 -664 0 feedthrough
rlabel pdiffusion 297 -664 297 -664 0 feedthrough
rlabel pdiffusion 304 -664 304 -664 0 feedthrough
rlabel pdiffusion 311 -664 311 -664 0 feedthrough
rlabel pdiffusion 318 -664 318 -664 0 cellNo=56
rlabel pdiffusion 325 -664 325 -664 0 feedthrough
rlabel pdiffusion 332 -664 332 -664 0 cellNo=389
rlabel pdiffusion 339 -664 339 -664 0 cellNo=526
rlabel pdiffusion 346 -664 346 -664 0 cellNo=206
rlabel pdiffusion 353 -664 353 -664 0 cellNo=690
rlabel pdiffusion 360 -664 360 -664 0 feedthrough
rlabel pdiffusion 367 -664 367 -664 0 feedthrough
rlabel pdiffusion 374 -664 374 -664 0 cellNo=54
rlabel pdiffusion 381 -664 381 -664 0 feedthrough
rlabel pdiffusion 388 -664 388 -664 0 feedthrough
rlabel pdiffusion 395 -664 395 -664 0 cellNo=686
rlabel pdiffusion 402 -664 402 -664 0 cellNo=427
rlabel pdiffusion 409 -664 409 -664 0 feedthrough
rlabel pdiffusion 416 -664 416 -664 0 feedthrough
rlabel pdiffusion 423 -664 423 -664 0 feedthrough
rlabel pdiffusion 430 -664 430 -664 0 feedthrough
rlabel pdiffusion 437 -664 437 -664 0 feedthrough
rlabel pdiffusion 444 -664 444 -664 0 feedthrough
rlabel pdiffusion 451 -664 451 -664 0 feedthrough
rlabel pdiffusion 458 -664 458 -664 0 feedthrough
rlabel pdiffusion 465 -664 465 -664 0 feedthrough
rlabel pdiffusion 472 -664 472 -664 0 cellNo=745
rlabel pdiffusion 479 -664 479 -664 0 feedthrough
rlabel pdiffusion 486 -664 486 -664 0 cellNo=273
rlabel pdiffusion 493 -664 493 -664 0 feedthrough
rlabel pdiffusion 500 -664 500 -664 0 feedthrough
rlabel pdiffusion 507 -664 507 -664 0 feedthrough
rlabel pdiffusion 514 -664 514 -664 0 cellNo=735
rlabel pdiffusion 521 -664 521 -664 0 feedthrough
rlabel pdiffusion 528 -664 528 -664 0 cellNo=287
rlabel pdiffusion 535 -664 535 -664 0 feedthrough
rlabel pdiffusion 542 -664 542 -664 0 cellNo=436
rlabel pdiffusion 549 -664 549 -664 0 feedthrough
rlabel pdiffusion 556 -664 556 -664 0 feedthrough
rlabel pdiffusion 563 -664 563 -664 0 cellNo=551
rlabel pdiffusion 584 -664 584 -664 0 feedthrough
rlabel pdiffusion 17 -713 17 -713 0 feedthrough
rlabel pdiffusion 24 -713 24 -713 0 feedthrough
rlabel pdiffusion 31 -713 31 -713 0 cellNo=213
rlabel pdiffusion 38 -713 38 -713 0 feedthrough
rlabel pdiffusion 45 -713 45 -713 0 feedthrough
rlabel pdiffusion 52 -713 52 -713 0 feedthrough
rlabel pdiffusion 59 -713 59 -713 0 cellNo=276
rlabel pdiffusion 66 -713 66 -713 0 cellNo=866
rlabel pdiffusion 73 -713 73 -713 0 cellNo=814
rlabel pdiffusion 80 -713 80 -713 0 feedthrough
rlabel pdiffusion 87 -713 87 -713 0 feedthrough
rlabel pdiffusion 94 -713 94 -713 0 feedthrough
rlabel pdiffusion 101 -713 101 -713 0 cellNo=879
rlabel pdiffusion 108 -713 108 -713 0 cellNo=336
rlabel pdiffusion 115 -713 115 -713 0 feedthrough
rlabel pdiffusion 122 -713 122 -713 0 feedthrough
rlabel pdiffusion 129 -713 129 -713 0 feedthrough
rlabel pdiffusion 136 -713 136 -713 0 cellNo=364
rlabel pdiffusion 143 -713 143 -713 0 feedthrough
rlabel pdiffusion 150 -713 150 -713 0 cellNo=149
rlabel pdiffusion 157 -713 157 -713 0 feedthrough
rlabel pdiffusion 164 -713 164 -713 0 cellNo=498
rlabel pdiffusion 171 -713 171 -713 0 feedthrough
rlabel pdiffusion 178 -713 178 -713 0 feedthrough
rlabel pdiffusion 185 -713 185 -713 0 cellNo=367
rlabel pdiffusion 192 -713 192 -713 0 cellNo=849
rlabel pdiffusion 199 -713 199 -713 0 cellNo=361
rlabel pdiffusion 206 -713 206 -713 0 feedthrough
rlabel pdiffusion 213 -713 213 -713 0 feedthrough
rlabel pdiffusion 220 -713 220 -713 0 cellNo=471
rlabel pdiffusion 227 -713 227 -713 0 feedthrough
rlabel pdiffusion 234 -713 234 -713 0 feedthrough
rlabel pdiffusion 241 -713 241 -713 0 feedthrough
rlabel pdiffusion 248 -713 248 -713 0 feedthrough
rlabel pdiffusion 255 -713 255 -713 0 feedthrough
rlabel pdiffusion 262 -713 262 -713 0 feedthrough
rlabel pdiffusion 269 -713 269 -713 0 feedthrough
rlabel pdiffusion 276 -713 276 -713 0 feedthrough
rlabel pdiffusion 283 -713 283 -713 0 cellNo=51
rlabel pdiffusion 290 -713 290 -713 0 feedthrough
rlabel pdiffusion 297 -713 297 -713 0 cellNo=776
rlabel pdiffusion 304 -713 304 -713 0 feedthrough
rlabel pdiffusion 311 -713 311 -713 0 cellNo=88
rlabel pdiffusion 318 -713 318 -713 0 feedthrough
rlabel pdiffusion 325 -713 325 -713 0 feedthrough
rlabel pdiffusion 332 -713 332 -713 0 cellNo=113
rlabel pdiffusion 339 -713 339 -713 0 cellNo=567
rlabel pdiffusion 346 -713 346 -713 0 cellNo=337
rlabel pdiffusion 353 -713 353 -713 0 feedthrough
rlabel pdiffusion 360 -713 360 -713 0 feedthrough
rlabel pdiffusion 367 -713 367 -713 0 feedthrough
rlabel pdiffusion 374 -713 374 -713 0 feedthrough
rlabel pdiffusion 381 -713 381 -713 0 cellNo=893
rlabel pdiffusion 388 -713 388 -713 0 cellNo=254
rlabel pdiffusion 395 -713 395 -713 0 cellNo=633
rlabel pdiffusion 402 -713 402 -713 0 feedthrough
rlabel pdiffusion 409 -713 409 -713 0 feedthrough
rlabel pdiffusion 416 -713 416 -713 0 feedthrough
rlabel pdiffusion 423 -713 423 -713 0 cellNo=843
rlabel pdiffusion 430 -713 430 -713 0 feedthrough
rlabel pdiffusion 437 -713 437 -713 0 feedthrough
rlabel pdiffusion 444 -713 444 -713 0 feedthrough
rlabel pdiffusion 451 -713 451 -713 0 feedthrough
rlabel pdiffusion 458 -713 458 -713 0 feedthrough
rlabel pdiffusion 465 -713 465 -713 0 feedthrough
rlabel pdiffusion 472 -713 472 -713 0 feedthrough
rlabel pdiffusion 479 -713 479 -713 0 feedthrough
rlabel pdiffusion 486 -713 486 -713 0 feedthrough
rlabel pdiffusion 493 -713 493 -713 0 cellNo=753
rlabel pdiffusion 500 -713 500 -713 0 feedthrough
rlabel pdiffusion 507 -713 507 -713 0 feedthrough
rlabel pdiffusion 514 -713 514 -713 0 feedthrough
rlabel pdiffusion 521 -713 521 -713 0 feedthrough
rlabel pdiffusion 528 -713 528 -713 0 feedthrough
rlabel pdiffusion 535 -713 535 -713 0 feedthrough
rlabel pdiffusion 542 -713 542 -713 0 feedthrough
rlabel pdiffusion 549 -713 549 -713 0 feedthrough
rlabel pdiffusion 556 -713 556 -713 0 feedthrough
rlabel pdiffusion 563 -713 563 -713 0 feedthrough
rlabel pdiffusion 570 -713 570 -713 0 cellNo=270
rlabel pdiffusion 577 -713 577 -713 0 feedthrough
rlabel pdiffusion 584 -713 584 -713 0 feedthrough
rlabel pdiffusion 591 -713 591 -713 0 cellNo=326
rlabel pdiffusion 598 -713 598 -713 0 cellNo=865
rlabel pdiffusion 605 -713 605 -713 0 feedthrough
rlabel pdiffusion 612 -713 612 -713 0 cellNo=402
rlabel pdiffusion 619 -713 619 -713 0 feedthrough
rlabel pdiffusion 626 -713 626 -713 0 cellNo=700
rlabel pdiffusion 633 -713 633 -713 0 feedthrough
rlabel pdiffusion 640 -713 640 -713 0 feedthrough
rlabel pdiffusion 647 -713 647 -713 0 feedthrough
rlabel pdiffusion 31 -764 31 -764 0 cellNo=400
rlabel pdiffusion 38 -764 38 -764 0 cellNo=817
rlabel pdiffusion 45 -764 45 -764 0 feedthrough
rlabel pdiffusion 52 -764 52 -764 0 feedthrough
rlabel pdiffusion 59 -764 59 -764 0 feedthrough
rlabel pdiffusion 66 -764 66 -764 0 feedthrough
rlabel pdiffusion 73 -764 73 -764 0 feedthrough
rlabel pdiffusion 80 -764 80 -764 0 feedthrough
rlabel pdiffusion 87 -764 87 -764 0 feedthrough
rlabel pdiffusion 94 -764 94 -764 0 feedthrough
rlabel pdiffusion 101 -764 101 -764 0 cellNo=485
rlabel pdiffusion 108 -764 108 -764 0 feedthrough
rlabel pdiffusion 115 -764 115 -764 0 cellNo=739
rlabel pdiffusion 122 -764 122 -764 0 feedthrough
rlabel pdiffusion 129 -764 129 -764 0 feedthrough
rlabel pdiffusion 136 -764 136 -764 0 cellNo=586
rlabel pdiffusion 143 -764 143 -764 0 cellNo=650
rlabel pdiffusion 150 -764 150 -764 0 cellNo=584
rlabel pdiffusion 157 -764 157 -764 0 feedthrough
rlabel pdiffusion 164 -764 164 -764 0 feedthrough
rlabel pdiffusion 171 -764 171 -764 0 feedthrough
rlabel pdiffusion 178 -764 178 -764 0 feedthrough
rlabel pdiffusion 185 -764 185 -764 0 feedthrough
rlabel pdiffusion 192 -764 192 -764 0 cellNo=701
rlabel pdiffusion 199 -764 199 -764 0 feedthrough
rlabel pdiffusion 206 -764 206 -764 0 cellNo=759
rlabel pdiffusion 213 -764 213 -764 0 cellNo=687
rlabel pdiffusion 220 -764 220 -764 0 cellNo=166
rlabel pdiffusion 227 -764 227 -764 0 cellNo=499
rlabel pdiffusion 234 -764 234 -764 0 feedthrough
rlabel pdiffusion 241 -764 241 -764 0 feedthrough
rlabel pdiffusion 248 -764 248 -764 0 cellNo=734
rlabel pdiffusion 255 -764 255 -764 0 cellNo=291
rlabel pdiffusion 262 -764 262 -764 0 feedthrough
rlabel pdiffusion 269 -764 269 -764 0 feedthrough
rlabel pdiffusion 276 -764 276 -764 0 cellNo=705
rlabel pdiffusion 283 -764 283 -764 0 cellNo=41
rlabel pdiffusion 290 -764 290 -764 0 cellNo=867
rlabel pdiffusion 297 -764 297 -764 0 feedthrough
rlabel pdiffusion 304 -764 304 -764 0 cellNo=126
rlabel pdiffusion 311 -764 311 -764 0 feedthrough
rlabel pdiffusion 318 -764 318 -764 0 feedthrough
rlabel pdiffusion 325 -764 325 -764 0 feedthrough
rlabel pdiffusion 332 -764 332 -764 0 cellNo=679
rlabel pdiffusion 339 -764 339 -764 0 cellNo=10
rlabel pdiffusion 346 -764 346 -764 0 cellNo=249
rlabel pdiffusion 353 -764 353 -764 0 feedthrough
rlabel pdiffusion 360 -764 360 -764 0 cellNo=111
rlabel pdiffusion 367 -764 367 -764 0 feedthrough
rlabel pdiffusion 374 -764 374 -764 0 cellNo=200
rlabel pdiffusion 381 -764 381 -764 0 feedthrough
rlabel pdiffusion 388 -764 388 -764 0 feedthrough
rlabel pdiffusion 395 -764 395 -764 0 cellNo=560
rlabel pdiffusion 402 -764 402 -764 0 feedthrough
rlabel pdiffusion 409 -764 409 -764 0 feedthrough
rlabel pdiffusion 416 -764 416 -764 0 feedthrough
rlabel pdiffusion 423 -764 423 -764 0 feedthrough
rlabel pdiffusion 430 -764 430 -764 0 feedthrough
rlabel pdiffusion 437 -764 437 -764 0 feedthrough
rlabel pdiffusion 444 -764 444 -764 0 cellNo=33
rlabel pdiffusion 451 -764 451 -764 0 feedthrough
rlabel pdiffusion 458 -764 458 -764 0 feedthrough
rlabel pdiffusion 465 -764 465 -764 0 feedthrough
rlabel pdiffusion 472 -764 472 -764 0 cellNo=23
rlabel pdiffusion 479 -764 479 -764 0 feedthrough
rlabel pdiffusion 486 -764 486 -764 0 cellNo=164
rlabel pdiffusion 493 -764 493 -764 0 feedthrough
rlabel pdiffusion 500 -764 500 -764 0 feedthrough
rlabel pdiffusion 507 -764 507 -764 0 feedthrough
rlabel pdiffusion 514 -764 514 -764 0 feedthrough
rlabel pdiffusion 521 -764 521 -764 0 feedthrough
rlabel pdiffusion 528 -764 528 -764 0 cellNo=272
rlabel pdiffusion 535 -764 535 -764 0 feedthrough
rlabel pdiffusion 542 -764 542 -764 0 feedthrough
rlabel pdiffusion 556 -764 556 -764 0 feedthrough
rlabel pdiffusion 612 -764 612 -764 0 cellNo=648
rlabel pdiffusion 24 -821 24 -821 0 cellNo=578
rlabel pdiffusion 31 -821 31 -821 0 cellNo=786
rlabel pdiffusion 38 -821 38 -821 0 feedthrough
rlabel pdiffusion 45 -821 45 -821 0 feedthrough
rlabel pdiffusion 52 -821 52 -821 0 feedthrough
rlabel pdiffusion 59 -821 59 -821 0 cellNo=295
rlabel pdiffusion 66 -821 66 -821 0 feedthrough
rlabel pdiffusion 73 -821 73 -821 0 cellNo=833
rlabel pdiffusion 80 -821 80 -821 0 feedthrough
rlabel pdiffusion 87 -821 87 -821 0 feedthrough
rlabel pdiffusion 94 -821 94 -821 0 feedthrough
rlabel pdiffusion 101 -821 101 -821 0 cellNo=804
rlabel pdiffusion 108 -821 108 -821 0 cellNo=799
rlabel pdiffusion 115 -821 115 -821 0 cellNo=275
rlabel pdiffusion 122 -821 122 -821 0 cellNo=694
rlabel pdiffusion 129 -821 129 -821 0 feedthrough
rlabel pdiffusion 136 -821 136 -821 0 feedthrough
rlabel pdiffusion 143 -821 143 -821 0 cellNo=134
rlabel pdiffusion 150 -821 150 -821 0 cellNo=666
rlabel pdiffusion 157 -821 157 -821 0 cellNo=492
rlabel pdiffusion 164 -821 164 -821 0 cellNo=828
rlabel pdiffusion 171 -821 171 -821 0 feedthrough
rlabel pdiffusion 178 -821 178 -821 0 feedthrough
rlabel pdiffusion 185 -821 185 -821 0 cellNo=1
rlabel pdiffusion 192 -821 192 -821 0 feedthrough
rlabel pdiffusion 199 -821 199 -821 0 cellNo=807
rlabel pdiffusion 206 -821 206 -821 0 feedthrough
rlabel pdiffusion 213 -821 213 -821 0 cellNo=268
rlabel pdiffusion 220 -821 220 -821 0 feedthrough
rlabel pdiffusion 227 -821 227 -821 0 feedthrough
rlabel pdiffusion 234 -821 234 -821 0 cellNo=741
rlabel pdiffusion 241 -821 241 -821 0 feedthrough
rlabel pdiffusion 248 -821 248 -821 0 cellNo=651
rlabel pdiffusion 255 -821 255 -821 0 cellNo=563
rlabel pdiffusion 262 -821 262 -821 0 cellNo=232
rlabel pdiffusion 269 -821 269 -821 0 feedthrough
rlabel pdiffusion 276 -821 276 -821 0 feedthrough
rlabel pdiffusion 283 -821 283 -821 0 feedthrough
rlabel pdiffusion 290 -821 290 -821 0 feedthrough
rlabel pdiffusion 297 -821 297 -821 0 cellNo=463
rlabel pdiffusion 304 -821 304 -821 0 feedthrough
rlabel pdiffusion 311 -821 311 -821 0 cellNo=778
rlabel pdiffusion 318 -821 318 -821 0 cellNo=385
rlabel pdiffusion 325 -821 325 -821 0 feedthrough
rlabel pdiffusion 332 -821 332 -821 0 cellNo=476
rlabel pdiffusion 339 -821 339 -821 0 feedthrough
rlabel pdiffusion 346 -821 346 -821 0 cellNo=835
rlabel pdiffusion 353 -821 353 -821 0 cellNo=425
rlabel pdiffusion 360 -821 360 -821 0 feedthrough
rlabel pdiffusion 367 -821 367 -821 0 feedthrough
rlabel pdiffusion 374 -821 374 -821 0 cellNo=721
rlabel pdiffusion 381 -821 381 -821 0 feedthrough
rlabel pdiffusion 388 -821 388 -821 0 feedthrough
rlabel pdiffusion 395 -821 395 -821 0 feedthrough
rlabel pdiffusion 402 -821 402 -821 0 cellNo=688
rlabel pdiffusion 409 -821 409 -821 0 feedthrough
rlabel pdiffusion 416 -821 416 -821 0 feedthrough
rlabel pdiffusion 423 -821 423 -821 0 feedthrough
rlabel pdiffusion 430 -821 430 -821 0 feedthrough
rlabel pdiffusion 437 -821 437 -821 0 feedthrough
rlabel pdiffusion 444 -821 444 -821 0 feedthrough
rlabel pdiffusion 451 -821 451 -821 0 feedthrough
rlabel pdiffusion 458 -821 458 -821 0 cellNo=888
rlabel pdiffusion 465 -821 465 -821 0 feedthrough
rlabel pdiffusion 472 -821 472 -821 0 feedthrough
rlabel pdiffusion 479 -821 479 -821 0 feedthrough
rlabel pdiffusion 486 -821 486 -821 0 feedthrough
rlabel pdiffusion 493 -821 493 -821 0 feedthrough
rlabel pdiffusion 500 -821 500 -821 0 feedthrough
rlabel pdiffusion 507 -821 507 -821 0 feedthrough
rlabel pdiffusion 514 -821 514 -821 0 feedthrough
rlabel pdiffusion 521 -821 521 -821 0 feedthrough
rlabel pdiffusion 528 -821 528 -821 0 feedthrough
rlabel pdiffusion 535 -821 535 -821 0 feedthrough
rlabel pdiffusion 542 -821 542 -821 0 feedthrough
rlabel pdiffusion 549 -821 549 -821 0 feedthrough
rlabel pdiffusion 556 -821 556 -821 0 cellNo=698
rlabel pdiffusion 24 -884 24 -884 0 cellNo=812
rlabel pdiffusion 31 -884 31 -884 0 cellNo=429
rlabel pdiffusion 38 -884 38 -884 0 cellNo=733
rlabel pdiffusion 45 -884 45 -884 0 cellNo=122
rlabel pdiffusion 52 -884 52 -884 0 feedthrough
rlabel pdiffusion 59 -884 59 -884 0 feedthrough
rlabel pdiffusion 66 -884 66 -884 0 feedthrough
rlabel pdiffusion 73 -884 73 -884 0 cellNo=32
rlabel pdiffusion 80 -884 80 -884 0 feedthrough
rlabel pdiffusion 87 -884 87 -884 0 feedthrough
rlabel pdiffusion 94 -884 94 -884 0 feedthrough
rlabel pdiffusion 101 -884 101 -884 0 feedthrough
rlabel pdiffusion 108 -884 108 -884 0 feedthrough
rlabel pdiffusion 115 -884 115 -884 0 cellNo=717
rlabel pdiffusion 122 -884 122 -884 0 cellNo=187
rlabel pdiffusion 129 -884 129 -884 0 cellNo=301
rlabel pdiffusion 136 -884 136 -884 0 cellNo=580
rlabel pdiffusion 143 -884 143 -884 0 feedthrough
rlabel pdiffusion 150 -884 150 -884 0 feedthrough
rlabel pdiffusion 157 -884 157 -884 0 cellNo=256
rlabel pdiffusion 164 -884 164 -884 0 cellNo=809
rlabel pdiffusion 171 -884 171 -884 0 cellNo=787
rlabel pdiffusion 178 -884 178 -884 0 cellNo=263
rlabel pdiffusion 185 -884 185 -884 0 feedthrough
rlabel pdiffusion 192 -884 192 -884 0 cellNo=414
rlabel pdiffusion 199 -884 199 -884 0 cellNo=190
rlabel pdiffusion 206 -884 206 -884 0 cellNo=884
rlabel pdiffusion 213 -884 213 -884 0 feedthrough
rlabel pdiffusion 220 -884 220 -884 0 feedthrough
rlabel pdiffusion 227 -884 227 -884 0 feedthrough
rlabel pdiffusion 234 -884 234 -884 0 feedthrough
rlabel pdiffusion 241 -884 241 -884 0 feedthrough
rlabel pdiffusion 248 -884 248 -884 0 feedthrough
rlabel pdiffusion 255 -884 255 -884 0 feedthrough
rlabel pdiffusion 262 -884 262 -884 0 feedthrough
rlabel pdiffusion 269 -884 269 -884 0 feedthrough
rlabel pdiffusion 276 -884 276 -884 0 feedthrough
rlabel pdiffusion 283 -884 283 -884 0 cellNo=823
rlabel pdiffusion 290 -884 290 -884 0 feedthrough
rlabel pdiffusion 297 -884 297 -884 0 cellNo=602
rlabel pdiffusion 304 -884 304 -884 0 cellNo=765
rlabel pdiffusion 311 -884 311 -884 0 cellNo=746
rlabel pdiffusion 318 -884 318 -884 0 feedthrough
rlabel pdiffusion 325 -884 325 -884 0 feedthrough
rlabel pdiffusion 332 -884 332 -884 0 cellNo=890
rlabel pdiffusion 339 -884 339 -884 0 feedthrough
rlabel pdiffusion 346 -884 346 -884 0 cellNo=672
rlabel pdiffusion 353 -884 353 -884 0 cellNo=70
rlabel pdiffusion 360 -884 360 -884 0 feedthrough
rlabel pdiffusion 367 -884 367 -884 0 feedthrough
rlabel pdiffusion 374 -884 374 -884 0 cellNo=626
rlabel pdiffusion 381 -884 381 -884 0 cellNo=558
rlabel pdiffusion 388 -884 388 -884 0 feedthrough
rlabel pdiffusion 395 -884 395 -884 0 feedthrough
rlabel pdiffusion 402 -884 402 -884 0 feedthrough
rlabel pdiffusion 409 -884 409 -884 0 feedthrough
rlabel pdiffusion 416 -884 416 -884 0 feedthrough
rlabel pdiffusion 423 -884 423 -884 0 feedthrough
rlabel pdiffusion 430 -884 430 -884 0 feedthrough
rlabel pdiffusion 437 -884 437 -884 0 feedthrough
rlabel pdiffusion 444 -884 444 -884 0 feedthrough
rlabel pdiffusion 451 -884 451 -884 0 feedthrough
rlabel pdiffusion 458 -884 458 -884 0 feedthrough
rlabel pdiffusion 465 -884 465 -884 0 cellNo=743
rlabel pdiffusion 472 -884 472 -884 0 cellNo=261
rlabel pdiffusion 479 -884 479 -884 0 feedthrough
rlabel pdiffusion 486 -884 486 -884 0 feedthrough
rlabel pdiffusion 493 -884 493 -884 0 feedthrough
rlabel pdiffusion 500 -884 500 -884 0 feedthrough
rlabel pdiffusion 507 -884 507 -884 0 feedthrough
rlabel pdiffusion 514 -884 514 -884 0 feedthrough
rlabel pdiffusion 521 -884 521 -884 0 cellNo=288
rlabel pdiffusion 528 -884 528 -884 0 feedthrough
rlabel pdiffusion 535 -884 535 -884 0 feedthrough
rlabel pdiffusion 10 -939 10 -939 0 feedthrough
rlabel pdiffusion 17 -939 17 -939 0 feedthrough
rlabel pdiffusion 24 -939 24 -939 0 feedthrough
rlabel pdiffusion 31 -939 31 -939 0 cellNo=524
rlabel pdiffusion 38 -939 38 -939 0 feedthrough
rlabel pdiffusion 45 -939 45 -939 0 cellNo=771
rlabel pdiffusion 52 -939 52 -939 0 feedthrough
rlabel pdiffusion 59 -939 59 -939 0 feedthrough
rlabel pdiffusion 66 -939 66 -939 0 feedthrough
rlabel pdiffusion 73 -939 73 -939 0 cellNo=216
rlabel pdiffusion 80 -939 80 -939 0 cellNo=359
rlabel pdiffusion 87 -939 87 -939 0 cellNo=647
rlabel pdiffusion 94 -939 94 -939 0 feedthrough
rlabel pdiffusion 101 -939 101 -939 0 cellNo=752
rlabel pdiffusion 108 -939 108 -939 0 feedthrough
rlabel pdiffusion 115 -939 115 -939 0 feedthrough
rlabel pdiffusion 122 -939 122 -939 0 feedthrough
rlabel pdiffusion 129 -939 129 -939 0 feedthrough
rlabel pdiffusion 136 -939 136 -939 0 cellNo=3
rlabel pdiffusion 143 -939 143 -939 0 feedthrough
rlabel pdiffusion 150 -939 150 -939 0 cellNo=872
rlabel pdiffusion 157 -939 157 -939 0 cellNo=589
rlabel pdiffusion 164 -939 164 -939 0 cellNo=386
rlabel pdiffusion 171 -939 171 -939 0 feedthrough
rlabel pdiffusion 178 -939 178 -939 0 feedthrough
rlabel pdiffusion 185 -939 185 -939 0 feedthrough
rlabel pdiffusion 192 -939 192 -939 0 cellNo=379
rlabel pdiffusion 199 -939 199 -939 0 cellNo=289
rlabel pdiffusion 206 -939 206 -939 0 cellNo=529
rlabel pdiffusion 213 -939 213 -939 0 cellNo=340
rlabel pdiffusion 220 -939 220 -939 0 cellNo=370
rlabel pdiffusion 227 -939 227 -939 0 cellNo=210
rlabel pdiffusion 234 -939 234 -939 0 feedthrough
rlabel pdiffusion 241 -939 241 -939 0 feedthrough
rlabel pdiffusion 248 -939 248 -939 0 feedthrough
rlabel pdiffusion 255 -939 255 -939 0 feedthrough
rlabel pdiffusion 262 -939 262 -939 0 cellNo=636
rlabel pdiffusion 269 -939 269 -939 0 feedthrough
rlabel pdiffusion 276 -939 276 -939 0 feedthrough
rlabel pdiffusion 283 -939 283 -939 0 feedthrough
rlabel pdiffusion 290 -939 290 -939 0 cellNo=197
rlabel pdiffusion 297 -939 297 -939 0 feedthrough
rlabel pdiffusion 304 -939 304 -939 0 cellNo=728
rlabel pdiffusion 311 -939 311 -939 0 feedthrough
rlabel pdiffusion 318 -939 318 -939 0 feedthrough
rlabel pdiffusion 325 -939 325 -939 0 cellNo=846
rlabel pdiffusion 332 -939 332 -939 0 cellNo=165
rlabel pdiffusion 339 -939 339 -939 0 feedthrough
rlabel pdiffusion 346 -939 346 -939 0 feedthrough
rlabel pdiffusion 353 -939 353 -939 0 cellNo=769
rlabel pdiffusion 360 -939 360 -939 0 feedthrough
rlabel pdiffusion 367 -939 367 -939 0 feedthrough
rlabel pdiffusion 374 -939 374 -939 0 feedthrough
rlabel pdiffusion 381 -939 381 -939 0 cellNo=130
rlabel pdiffusion 388 -939 388 -939 0 feedthrough
rlabel pdiffusion 395 -939 395 -939 0 cellNo=454
rlabel pdiffusion 402 -939 402 -939 0 feedthrough
rlabel pdiffusion 409 -939 409 -939 0 cellNo=455
rlabel pdiffusion 416 -939 416 -939 0 feedthrough
rlabel pdiffusion 423 -939 423 -939 0 feedthrough
rlabel pdiffusion 430 -939 430 -939 0 feedthrough
rlabel pdiffusion 437 -939 437 -939 0 feedthrough
rlabel pdiffusion 444 -939 444 -939 0 cellNo=501
rlabel pdiffusion 451 -939 451 -939 0 feedthrough
rlabel pdiffusion 458 -939 458 -939 0 feedthrough
rlabel pdiffusion 465 -939 465 -939 0 cellNo=616
rlabel pdiffusion 472 -939 472 -939 0 feedthrough
rlabel pdiffusion 479 -939 479 -939 0 feedthrough
rlabel pdiffusion 486 -939 486 -939 0 feedthrough
rlabel pdiffusion 493 -939 493 -939 0 feedthrough
rlabel pdiffusion 500 -939 500 -939 0 feedthrough
rlabel pdiffusion 507 -939 507 -939 0 feedthrough
rlabel pdiffusion 514 -939 514 -939 0 feedthrough
rlabel pdiffusion 521 -939 521 -939 0 feedthrough
rlabel pdiffusion 3 -988 3 -988 0 feedthrough
rlabel pdiffusion 10 -988 10 -988 0 feedthrough
rlabel pdiffusion 17 -988 17 -988 0 cellNo=712
rlabel pdiffusion 24 -988 24 -988 0 cellNo=90
rlabel pdiffusion 31 -988 31 -988 0 cellNo=127
rlabel pdiffusion 38 -988 38 -988 0 cellNo=259
rlabel pdiffusion 45 -988 45 -988 0 feedthrough
rlabel pdiffusion 52 -988 52 -988 0 feedthrough
rlabel pdiffusion 59 -988 59 -988 0 cellNo=151
rlabel pdiffusion 66 -988 66 -988 0 feedthrough
rlabel pdiffusion 73 -988 73 -988 0 cellNo=858
rlabel pdiffusion 80 -988 80 -988 0 cellNo=863
rlabel pdiffusion 87 -988 87 -988 0 feedthrough
rlabel pdiffusion 94 -988 94 -988 0 cellNo=194
rlabel pdiffusion 101 -988 101 -988 0 cellNo=699
rlabel pdiffusion 108 -988 108 -988 0 feedthrough
rlabel pdiffusion 115 -988 115 -988 0 feedthrough
rlabel pdiffusion 122 -988 122 -988 0 feedthrough
rlabel pdiffusion 129 -988 129 -988 0 cellNo=649
rlabel pdiffusion 136 -988 136 -988 0 cellNo=585
rlabel pdiffusion 143 -988 143 -988 0 feedthrough
rlabel pdiffusion 150 -988 150 -988 0 feedthrough
rlabel pdiffusion 157 -988 157 -988 0 cellNo=676
rlabel pdiffusion 164 -988 164 -988 0 cellNo=125
rlabel pdiffusion 171 -988 171 -988 0 feedthrough
rlabel pdiffusion 178 -988 178 -988 0 cellNo=854
rlabel pdiffusion 185 -988 185 -988 0 cellNo=50
rlabel pdiffusion 192 -988 192 -988 0 cellNo=520
rlabel pdiffusion 199 -988 199 -988 0 cellNo=614
rlabel pdiffusion 206 -988 206 -988 0 feedthrough
rlabel pdiffusion 213 -988 213 -988 0 feedthrough
rlabel pdiffusion 220 -988 220 -988 0 cellNo=610
rlabel pdiffusion 227 -988 227 -988 0 cellNo=813
rlabel pdiffusion 234 -988 234 -988 0 cellNo=265
rlabel pdiffusion 241 -988 241 -988 0 cellNo=169
rlabel pdiffusion 248 -988 248 -988 0 feedthrough
rlabel pdiffusion 255 -988 255 -988 0 cellNo=790
rlabel pdiffusion 262 -988 262 -988 0 cellNo=604
rlabel pdiffusion 269 -988 269 -988 0 feedthrough
rlabel pdiffusion 276 -988 276 -988 0 feedthrough
rlabel pdiffusion 283 -988 283 -988 0 feedthrough
rlabel pdiffusion 290 -988 290 -988 0 cellNo=299
rlabel pdiffusion 297 -988 297 -988 0 cellNo=435
rlabel pdiffusion 304 -988 304 -988 0 feedthrough
rlabel pdiffusion 311 -988 311 -988 0 feedthrough
rlabel pdiffusion 318 -988 318 -988 0 feedthrough
rlabel pdiffusion 325 -988 325 -988 0 feedthrough
rlabel pdiffusion 332 -988 332 -988 0 cellNo=62
rlabel pdiffusion 339 -988 339 -988 0 cellNo=27
rlabel pdiffusion 346 -988 346 -988 0 feedthrough
rlabel pdiffusion 353 -988 353 -988 0 cellNo=112
rlabel pdiffusion 360 -988 360 -988 0 feedthrough
rlabel pdiffusion 367 -988 367 -988 0 feedthrough
rlabel pdiffusion 374 -988 374 -988 0 feedthrough
rlabel pdiffusion 381 -988 381 -988 0 feedthrough
rlabel pdiffusion 388 -988 388 -988 0 feedthrough
rlabel pdiffusion 395 -988 395 -988 0 feedthrough
rlabel pdiffusion 402 -988 402 -988 0 feedthrough
rlabel pdiffusion 409 -988 409 -988 0 feedthrough
rlabel pdiffusion 416 -988 416 -988 0 feedthrough
rlabel pdiffusion 423 -988 423 -988 0 feedthrough
rlabel pdiffusion 430 -988 430 -988 0 feedthrough
rlabel pdiffusion 437 -988 437 -988 0 feedthrough
rlabel pdiffusion 444 -988 444 -988 0 feedthrough
rlabel pdiffusion 451 -988 451 -988 0 feedthrough
rlabel pdiffusion 458 -988 458 -988 0 feedthrough
rlabel pdiffusion 465 -988 465 -988 0 cellNo=779
rlabel pdiffusion 472 -988 472 -988 0 cellNo=583
rlabel pdiffusion 479 -988 479 -988 0 feedthrough
rlabel pdiffusion 493 -988 493 -988 0 feedthrough
rlabel pdiffusion 507 -988 507 -988 0 feedthrough
rlabel pdiffusion 17 -1035 17 -1035 0 cellNo=597
rlabel pdiffusion 24 -1035 24 -1035 0 feedthrough
rlabel pdiffusion 31 -1035 31 -1035 0 cellNo=850
rlabel pdiffusion 38 -1035 38 -1035 0 feedthrough
rlabel pdiffusion 45 -1035 45 -1035 0 cellNo=861
rlabel pdiffusion 59 -1035 59 -1035 0 feedthrough
rlabel pdiffusion 80 -1035 80 -1035 0 cellNo=675
rlabel pdiffusion 87 -1035 87 -1035 0 feedthrough
rlabel pdiffusion 94 -1035 94 -1035 0 cellNo=605
rlabel pdiffusion 101 -1035 101 -1035 0 cellNo=390
rlabel pdiffusion 108 -1035 108 -1035 0 feedthrough
rlabel pdiffusion 115 -1035 115 -1035 0 feedthrough
rlabel pdiffusion 122 -1035 122 -1035 0 feedthrough
rlabel pdiffusion 129 -1035 129 -1035 0 feedthrough
rlabel pdiffusion 136 -1035 136 -1035 0 cellNo=533
rlabel pdiffusion 143 -1035 143 -1035 0 feedthrough
rlabel pdiffusion 150 -1035 150 -1035 0 cellNo=507
rlabel pdiffusion 157 -1035 157 -1035 0 cellNo=396
rlabel pdiffusion 164 -1035 164 -1035 0 cellNo=483
rlabel pdiffusion 171 -1035 171 -1035 0 feedthrough
rlabel pdiffusion 178 -1035 178 -1035 0 feedthrough
rlabel pdiffusion 185 -1035 185 -1035 0 cellNo=468
rlabel pdiffusion 192 -1035 192 -1035 0 feedthrough
rlabel pdiffusion 199 -1035 199 -1035 0 feedthrough
rlabel pdiffusion 206 -1035 206 -1035 0 feedthrough
rlabel pdiffusion 213 -1035 213 -1035 0 cellNo=132
rlabel pdiffusion 220 -1035 220 -1035 0 cellNo=729
rlabel pdiffusion 227 -1035 227 -1035 0 cellNo=855
rlabel pdiffusion 234 -1035 234 -1035 0 feedthrough
rlabel pdiffusion 241 -1035 241 -1035 0 feedthrough
rlabel pdiffusion 248 -1035 248 -1035 0 feedthrough
rlabel pdiffusion 255 -1035 255 -1035 0 feedthrough
rlabel pdiffusion 262 -1035 262 -1035 0 feedthrough
rlabel pdiffusion 269 -1035 269 -1035 0 feedthrough
rlabel pdiffusion 276 -1035 276 -1035 0 cellNo=6
rlabel pdiffusion 283 -1035 283 -1035 0 cellNo=681
rlabel pdiffusion 290 -1035 290 -1035 0 feedthrough
rlabel pdiffusion 297 -1035 297 -1035 0 cellNo=545
rlabel pdiffusion 304 -1035 304 -1035 0 cellNo=308
rlabel pdiffusion 311 -1035 311 -1035 0 feedthrough
rlabel pdiffusion 318 -1035 318 -1035 0 feedthrough
rlabel pdiffusion 325 -1035 325 -1035 0 cellNo=873
rlabel pdiffusion 332 -1035 332 -1035 0 cellNo=458
rlabel pdiffusion 339 -1035 339 -1035 0 cellNo=363
rlabel pdiffusion 346 -1035 346 -1035 0 feedthrough
rlabel pdiffusion 353 -1035 353 -1035 0 feedthrough
rlabel pdiffusion 360 -1035 360 -1035 0 feedthrough
rlabel pdiffusion 367 -1035 367 -1035 0 feedthrough
rlabel pdiffusion 374 -1035 374 -1035 0 feedthrough
rlabel pdiffusion 381 -1035 381 -1035 0 feedthrough
rlabel pdiffusion 388 -1035 388 -1035 0 feedthrough
rlabel pdiffusion 395 -1035 395 -1035 0 feedthrough
rlabel pdiffusion 402 -1035 402 -1035 0 feedthrough
rlabel pdiffusion 409 -1035 409 -1035 0 feedthrough
rlabel pdiffusion 416 -1035 416 -1035 0 cellNo=325
rlabel pdiffusion 423 -1035 423 -1035 0 cellNo=306
rlabel pdiffusion 430 -1035 430 -1035 0 feedthrough
rlabel pdiffusion 437 -1035 437 -1035 0 cellNo=742
rlabel pdiffusion 444 -1035 444 -1035 0 cellNo=715
rlabel pdiffusion 451 -1035 451 -1035 0 feedthrough
rlabel pdiffusion 458 -1035 458 -1035 0 cellNo=713
rlabel pdiffusion 465 -1035 465 -1035 0 cellNo=19
rlabel pdiffusion 472 -1035 472 -1035 0 feedthrough
rlabel pdiffusion 479 -1035 479 -1035 0 feedthrough
rlabel pdiffusion 486 -1035 486 -1035 0 cellNo=4
rlabel pdiffusion 31 -1080 31 -1080 0 feedthrough
rlabel pdiffusion 38 -1080 38 -1080 0 feedthrough
rlabel pdiffusion 45 -1080 45 -1080 0 cellNo=212
rlabel pdiffusion 52 -1080 52 -1080 0 feedthrough
rlabel pdiffusion 59 -1080 59 -1080 0 cellNo=172
rlabel pdiffusion 66 -1080 66 -1080 0 cellNo=840
rlabel pdiffusion 73 -1080 73 -1080 0 feedthrough
rlabel pdiffusion 80 -1080 80 -1080 0 feedthrough
rlabel pdiffusion 87 -1080 87 -1080 0 feedthrough
rlabel pdiffusion 94 -1080 94 -1080 0 cellNo=523
rlabel pdiffusion 101 -1080 101 -1080 0 feedthrough
rlabel pdiffusion 108 -1080 108 -1080 0 cellNo=353
rlabel pdiffusion 115 -1080 115 -1080 0 cellNo=587
rlabel pdiffusion 122 -1080 122 -1080 0 feedthrough
rlabel pdiffusion 129 -1080 129 -1080 0 feedthrough
rlabel pdiffusion 136 -1080 136 -1080 0 feedthrough
rlabel pdiffusion 143 -1080 143 -1080 0 cellNo=406
rlabel pdiffusion 150 -1080 150 -1080 0 cellNo=611
rlabel pdiffusion 157 -1080 157 -1080 0 cellNo=188
rlabel pdiffusion 164 -1080 164 -1080 0 cellNo=749
rlabel pdiffusion 171 -1080 171 -1080 0 cellNo=482
rlabel pdiffusion 178 -1080 178 -1080 0 feedthrough
rlabel pdiffusion 185 -1080 185 -1080 0 feedthrough
rlabel pdiffusion 192 -1080 192 -1080 0 cellNo=193
rlabel pdiffusion 199 -1080 199 -1080 0 cellNo=18
rlabel pdiffusion 206 -1080 206 -1080 0 feedthrough
rlabel pdiffusion 213 -1080 213 -1080 0 cellNo=874
rlabel pdiffusion 220 -1080 220 -1080 0 cellNo=168
rlabel pdiffusion 227 -1080 227 -1080 0 cellNo=7
rlabel pdiffusion 234 -1080 234 -1080 0 cellNo=329
rlabel pdiffusion 241 -1080 241 -1080 0 feedthrough
rlabel pdiffusion 248 -1080 248 -1080 0 feedthrough
rlabel pdiffusion 255 -1080 255 -1080 0 feedthrough
rlabel pdiffusion 262 -1080 262 -1080 0 feedthrough
rlabel pdiffusion 269 -1080 269 -1080 0 cellNo=155
rlabel pdiffusion 276 -1080 276 -1080 0 cellNo=75
rlabel pdiffusion 283 -1080 283 -1080 0 cellNo=176
rlabel pdiffusion 290 -1080 290 -1080 0 cellNo=528
rlabel pdiffusion 297 -1080 297 -1080 0 feedthrough
rlabel pdiffusion 304 -1080 304 -1080 0 cellNo=107
rlabel pdiffusion 311 -1080 311 -1080 0 feedthrough
rlabel pdiffusion 318 -1080 318 -1080 0 feedthrough
rlabel pdiffusion 325 -1080 325 -1080 0 feedthrough
rlabel pdiffusion 332 -1080 332 -1080 0 feedthrough
rlabel pdiffusion 339 -1080 339 -1080 0 cellNo=815
rlabel pdiffusion 346 -1080 346 -1080 0 cellNo=192
rlabel pdiffusion 353 -1080 353 -1080 0 feedthrough
rlabel pdiffusion 360 -1080 360 -1080 0 feedthrough
rlabel pdiffusion 367 -1080 367 -1080 0 feedthrough
rlabel pdiffusion 374 -1080 374 -1080 0 feedthrough
rlabel pdiffusion 381 -1080 381 -1080 0 feedthrough
rlabel pdiffusion 388 -1080 388 -1080 0 feedthrough
rlabel pdiffusion 395 -1080 395 -1080 0 feedthrough
rlabel pdiffusion 402 -1080 402 -1080 0 feedthrough
rlabel pdiffusion 409 -1080 409 -1080 0 feedthrough
rlabel pdiffusion 416 -1080 416 -1080 0 feedthrough
rlabel pdiffusion 423 -1080 423 -1080 0 feedthrough
rlabel pdiffusion 430 -1080 430 -1080 0 feedthrough
rlabel pdiffusion 437 -1080 437 -1080 0 feedthrough
rlabel pdiffusion 444 -1080 444 -1080 0 feedthrough
rlabel pdiffusion 451 -1080 451 -1080 0 feedthrough
rlabel pdiffusion 458 -1080 458 -1080 0 feedthrough
rlabel pdiffusion 465 -1080 465 -1080 0 feedthrough
rlabel pdiffusion 472 -1080 472 -1080 0 cellNo=451
rlabel pdiffusion 479 -1080 479 -1080 0 cellNo=663
rlabel pdiffusion 486 -1080 486 -1080 0 feedthrough
rlabel pdiffusion 493 -1080 493 -1080 0 cellNo=639
rlabel pdiffusion 500 -1080 500 -1080 0 feedthrough
rlabel pdiffusion 45 -1113 45 -1113 0 cellNo=294
rlabel pdiffusion 66 -1113 66 -1113 0 feedthrough
rlabel pdiffusion 73 -1113 73 -1113 0 feedthrough
rlabel pdiffusion 80 -1113 80 -1113 0 cellNo=897
rlabel pdiffusion 87 -1113 87 -1113 0 cellNo=860
rlabel pdiffusion 94 -1113 94 -1113 0 cellNo=46
rlabel pdiffusion 101 -1113 101 -1113 0 feedthrough
rlabel pdiffusion 108 -1113 108 -1113 0 cellNo=373
rlabel pdiffusion 115 -1113 115 -1113 0 feedthrough
rlabel pdiffusion 122 -1113 122 -1113 0 cellNo=722
rlabel pdiffusion 129 -1113 129 -1113 0 feedthrough
rlabel pdiffusion 136 -1113 136 -1113 0 feedthrough
rlabel pdiffusion 143 -1113 143 -1113 0 cellNo=493
rlabel pdiffusion 150 -1113 150 -1113 0 feedthrough
rlabel pdiffusion 157 -1113 157 -1113 0 feedthrough
rlabel pdiffusion 164 -1113 164 -1113 0 cellNo=731
rlabel pdiffusion 171 -1113 171 -1113 0 feedthrough
rlabel pdiffusion 178 -1113 178 -1113 0 feedthrough
rlabel pdiffusion 185 -1113 185 -1113 0 feedthrough
rlabel pdiffusion 192 -1113 192 -1113 0 cellNo=674
rlabel pdiffusion 199 -1113 199 -1113 0 cellNo=562
rlabel pdiffusion 206 -1113 206 -1113 0 cellNo=472
rlabel pdiffusion 213 -1113 213 -1113 0 cellNo=171
rlabel pdiffusion 220 -1113 220 -1113 0 cellNo=37
rlabel pdiffusion 227 -1113 227 -1113 0 cellNo=877
rlabel pdiffusion 234 -1113 234 -1113 0 cellNo=310
rlabel pdiffusion 241 -1113 241 -1113 0 feedthrough
rlabel pdiffusion 248 -1113 248 -1113 0 cellNo=239
rlabel pdiffusion 255 -1113 255 -1113 0 feedthrough
rlabel pdiffusion 262 -1113 262 -1113 0 feedthrough
rlabel pdiffusion 269 -1113 269 -1113 0 cellNo=645
rlabel pdiffusion 276 -1113 276 -1113 0 feedthrough
rlabel pdiffusion 283 -1113 283 -1113 0 cellNo=377
rlabel pdiffusion 290 -1113 290 -1113 0 feedthrough
rlabel pdiffusion 297 -1113 297 -1113 0 feedthrough
rlabel pdiffusion 304 -1113 304 -1113 0 feedthrough
rlabel pdiffusion 311 -1113 311 -1113 0 cellNo=706
rlabel pdiffusion 318 -1113 318 -1113 0 feedthrough
rlabel pdiffusion 325 -1113 325 -1113 0 feedthrough
rlabel pdiffusion 332 -1113 332 -1113 0 cellNo=864
rlabel pdiffusion 339 -1113 339 -1113 0 feedthrough
rlabel pdiffusion 346 -1113 346 -1113 0 feedthrough
rlabel pdiffusion 353 -1113 353 -1113 0 cellNo=685
rlabel pdiffusion 360 -1113 360 -1113 0 feedthrough
rlabel pdiffusion 367 -1113 367 -1113 0 cellNo=280
rlabel pdiffusion 374 -1113 374 -1113 0 feedthrough
rlabel pdiffusion 381 -1113 381 -1113 0 feedthrough
rlabel pdiffusion 388 -1113 388 -1113 0 feedthrough
rlabel pdiffusion 395 -1113 395 -1113 0 cellNo=446
rlabel pdiffusion 402 -1113 402 -1113 0 feedthrough
rlabel pdiffusion 409 -1113 409 -1113 0 cellNo=725
rlabel pdiffusion 416 -1113 416 -1113 0 feedthrough
rlabel pdiffusion 423 -1113 423 -1113 0 feedthrough
rlabel pdiffusion 430 -1113 430 -1113 0 cellNo=723
rlabel pdiffusion 437 -1113 437 -1113 0 feedthrough
rlabel pdiffusion 444 -1113 444 -1113 0 feedthrough
rlabel pdiffusion 451 -1113 451 -1113 0 cellNo=707
rlabel pdiffusion 458 -1113 458 -1113 0 feedthrough
rlabel pdiffusion 45 -1146 45 -1146 0 cellNo=243
rlabel pdiffusion 52 -1146 52 -1146 0 feedthrough
rlabel pdiffusion 59 -1146 59 -1146 0 cellNo=79
rlabel pdiffusion 66 -1146 66 -1146 0 feedthrough
rlabel pdiffusion 73 -1146 73 -1146 0 cellNo=829
rlabel pdiffusion 80 -1146 80 -1146 0 cellNo=443
rlabel pdiffusion 87 -1146 87 -1146 0 cellNo=330
rlabel pdiffusion 94 -1146 94 -1146 0 cellNo=490
rlabel pdiffusion 101 -1146 101 -1146 0 feedthrough
rlabel pdiffusion 108 -1146 108 -1146 0 cellNo=763
rlabel pdiffusion 115 -1146 115 -1146 0 feedthrough
rlabel pdiffusion 122 -1146 122 -1146 0 feedthrough
rlabel pdiffusion 129 -1146 129 -1146 0 cellNo=510
rlabel pdiffusion 136 -1146 136 -1146 0 cellNo=703
rlabel pdiffusion 143 -1146 143 -1146 0 feedthrough
rlabel pdiffusion 150 -1146 150 -1146 0 feedthrough
rlabel pdiffusion 157 -1146 157 -1146 0 feedthrough
rlabel pdiffusion 164 -1146 164 -1146 0 feedthrough
rlabel pdiffusion 171 -1146 171 -1146 0 feedthrough
rlabel pdiffusion 178 -1146 178 -1146 0 feedthrough
rlabel pdiffusion 185 -1146 185 -1146 0 cellNo=637
rlabel pdiffusion 192 -1146 192 -1146 0 cellNo=29
rlabel pdiffusion 199 -1146 199 -1146 0 feedthrough
rlabel pdiffusion 206 -1146 206 -1146 0 cellNo=96
rlabel pdiffusion 213 -1146 213 -1146 0 cellNo=104
rlabel pdiffusion 220 -1146 220 -1146 0 cellNo=869
rlabel pdiffusion 227 -1146 227 -1146 0 cellNo=462
rlabel pdiffusion 234 -1146 234 -1146 0 feedthrough
rlabel pdiffusion 241 -1146 241 -1146 0 cellNo=240
rlabel pdiffusion 248 -1146 248 -1146 0 cellNo=678
rlabel pdiffusion 255 -1146 255 -1146 0 cellNo=242
rlabel pdiffusion 262 -1146 262 -1146 0 feedthrough
rlabel pdiffusion 269 -1146 269 -1146 0 cellNo=883
rlabel pdiffusion 276 -1146 276 -1146 0 feedthrough
rlabel pdiffusion 283 -1146 283 -1146 0 feedthrough
rlabel pdiffusion 290 -1146 290 -1146 0 feedthrough
rlabel pdiffusion 297 -1146 297 -1146 0 feedthrough
rlabel pdiffusion 304 -1146 304 -1146 0 cellNo=677
rlabel pdiffusion 311 -1146 311 -1146 0 cellNo=199
rlabel pdiffusion 318 -1146 318 -1146 0 feedthrough
rlabel pdiffusion 325 -1146 325 -1146 0 feedthrough
rlabel pdiffusion 332 -1146 332 -1146 0 feedthrough
rlabel pdiffusion 339 -1146 339 -1146 0 feedthrough
rlabel pdiffusion 346 -1146 346 -1146 0 feedthrough
rlabel pdiffusion 353 -1146 353 -1146 0 feedthrough
rlabel pdiffusion 360 -1146 360 -1146 0 feedthrough
rlabel pdiffusion 367 -1146 367 -1146 0 feedthrough
rlabel pdiffusion 374 -1146 374 -1146 0 feedthrough
rlabel pdiffusion 381 -1146 381 -1146 0 cellNo=891
rlabel pdiffusion 388 -1146 388 -1146 0 cellNo=521
rlabel pdiffusion 395 -1146 395 -1146 0 feedthrough
rlabel pdiffusion 402 -1146 402 -1146 0 cellNo=532
rlabel pdiffusion 409 -1146 409 -1146 0 feedthrough
rlabel pdiffusion 416 -1146 416 -1146 0 feedthrough
rlabel pdiffusion 423 -1146 423 -1146 0 feedthrough
rlabel pdiffusion 444 -1146 444 -1146 0 cellNo=569
rlabel pdiffusion 451 -1146 451 -1146 0 feedthrough
rlabel pdiffusion 45 -1183 45 -1183 0 cellNo=702
rlabel pdiffusion 52 -1183 52 -1183 0 feedthrough
rlabel pdiffusion 59 -1183 59 -1183 0 cellNo=34
rlabel pdiffusion 66 -1183 66 -1183 0 cellNo=750
rlabel pdiffusion 73 -1183 73 -1183 0 cellNo=811
rlabel pdiffusion 80 -1183 80 -1183 0 cellNo=772
rlabel pdiffusion 87 -1183 87 -1183 0 cellNo=660
rlabel pdiffusion 94 -1183 94 -1183 0 cellNo=478
rlabel pdiffusion 101 -1183 101 -1183 0 feedthrough
rlabel pdiffusion 108 -1183 108 -1183 0 feedthrough
rlabel pdiffusion 115 -1183 115 -1183 0 cellNo=886
rlabel pdiffusion 122 -1183 122 -1183 0 feedthrough
rlabel pdiffusion 129 -1183 129 -1183 0 feedthrough
rlabel pdiffusion 136 -1183 136 -1183 0 feedthrough
rlabel pdiffusion 143 -1183 143 -1183 0 cellNo=781
rlabel pdiffusion 150 -1183 150 -1183 0 cellNo=826
rlabel pdiffusion 157 -1183 157 -1183 0 feedthrough
rlabel pdiffusion 164 -1183 164 -1183 0 cellNo=290
rlabel pdiffusion 171 -1183 171 -1183 0 cellNo=45
rlabel pdiffusion 178 -1183 178 -1183 0 cellNo=277
rlabel pdiffusion 185 -1183 185 -1183 0 feedthrough
rlabel pdiffusion 192 -1183 192 -1183 0 cellNo=101
rlabel pdiffusion 199 -1183 199 -1183 0 cellNo=613
rlabel pdiffusion 206 -1183 206 -1183 0 feedthrough
rlabel pdiffusion 213 -1183 213 -1183 0 feedthrough
rlabel pdiffusion 220 -1183 220 -1183 0 cellNo=770
rlabel pdiffusion 227 -1183 227 -1183 0 cellNo=714
rlabel pdiffusion 234 -1183 234 -1183 0 cellNo=789
rlabel pdiffusion 241 -1183 241 -1183 0 cellNo=853
rlabel pdiffusion 248 -1183 248 -1183 0 cellNo=433
rlabel pdiffusion 255 -1183 255 -1183 0 cellNo=669
rlabel pdiffusion 262 -1183 262 -1183 0 feedthrough
rlabel pdiffusion 269 -1183 269 -1183 0 feedthrough
rlabel pdiffusion 276 -1183 276 -1183 0 feedthrough
rlabel pdiffusion 283 -1183 283 -1183 0 feedthrough
rlabel pdiffusion 290 -1183 290 -1183 0 cellNo=768
rlabel pdiffusion 297 -1183 297 -1183 0 cellNo=887
rlabel pdiffusion 304 -1183 304 -1183 0 cellNo=495
rlabel pdiffusion 311 -1183 311 -1183 0 feedthrough
rlabel pdiffusion 318 -1183 318 -1183 0 feedthrough
rlabel pdiffusion 325 -1183 325 -1183 0 feedthrough
rlabel pdiffusion 332 -1183 332 -1183 0 feedthrough
rlabel pdiffusion 339 -1183 339 -1183 0 feedthrough
rlabel pdiffusion 346 -1183 346 -1183 0 cellNo=453
rlabel pdiffusion 353 -1183 353 -1183 0 feedthrough
rlabel pdiffusion 360 -1183 360 -1183 0 feedthrough
rlabel pdiffusion 367 -1183 367 -1183 0 feedthrough
rlabel pdiffusion 374 -1183 374 -1183 0 feedthrough
rlabel pdiffusion 381 -1183 381 -1183 0 feedthrough
rlabel pdiffusion 388 -1183 388 -1183 0 feedthrough
rlabel pdiffusion 395 -1183 395 -1183 0 feedthrough
rlabel pdiffusion 402 -1183 402 -1183 0 feedthrough
rlabel pdiffusion 416 -1183 416 -1183 0 cellNo=630
rlabel pdiffusion 423 -1183 423 -1183 0 feedthrough
rlabel pdiffusion 430 -1183 430 -1183 0 feedthrough
rlabel pdiffusion 45 -1210 45 -1210 0 cellNo=821
rlabel pdiffusion 66 -1210 66 -1210 0 cellNo=13
rlabel pdiffusion 73 -1210 73 -1210 0 feedthrough
rlabel pdiffusion 80 -1210 80 -1210 0 cellNo=84
rlabel pdiffusion 87 -1210 87 -1210 0 cellNo=625
rlabel pdiffusion 94 -1210 94 -1210 0 cellNo=880
rlabel pdiffusion 101 -1210 101 -1210 0 feedthrough
rlabel pdiffusion 108 -1210 108 -1210 0 feedthrough
rlabel pdiffusion 115 -1210 115 -1210 0 cellNo=488
rlabel pdiffusion 122 -1210 122 -1210 0 feedthrough
rlabel pdiffusion 129 -1210 129 -1210 0 feedthrough
rlabel pdiffusion 136 -1210 136 -1210 0 cellNo=836
rlabel pdiffusion 143 -1210 143 -1210 0 cellNo=120
rlabel pdiffusion 150 -1210 150 -1210 0 cellNo=549
rlabel pdiffusion 157 -1210 157 -1210 0 cellNo=264
rlabel pdiffusion 164 -1210 164 -1210 0 cellNo=25
rlabel pdiffusion 171 -1210 171 -1210 0 feedthrough
rlabel pdiffusion 178 -1210 178 -1210 0 feedthrough
rlabel pdiffusion 185 -1210 185 -1210 0 cellNo=145
rlabel pdiffusion 192 -1210 192 -1210 0 cellNo=494
rlabel pdiffusion 199 -1210 199 -1210 0 feedthrough
rlabel pdiffusion 206 -1210 206 -1210 0 feedthrough
rlabel pdiffusion 213 -1210 213 -1210 0 feedthrough
rlabel pdiffusion 220 -1210 220 -1210 0 cellNo=661
rlabel pdiffusion 227 -1210 227 -1210 0 cellNo=627
rlabel pdiffusion 234 -1210 234 -1210 0 feedthrough
rlabel pdiffusion 241 -1210 241 -1210 0 cellNo=852
rlabel pdiffusion 248 -1210 248 -1210 0 feedthrough
rlabel pdiffusion 255 -1210 255 -1210 0 feedthrough
rlabel pdiffusion 283 -1210 283 -1210 0 feedthrough
rlabel pdiffusion 290 -1210 290 -1210 0 cellNo=434
rlabel pdiffusion 297 -1210 297 -1210 0 feedthrough
rlabel pdiffusion 304 -1210 304 -1210 0 cellNo=15
rlabel pdiffusion 311 -1210 311 -1210 0 cellNo=457
rlabel pdiffusion 318 -1210 318 -1210 0 feedthrough
rlabel pdiffusion 325 -1210 325 -1210 0 feedthrough
rlabel pdiffusion 332 -1210 332 -1210 0 feedthrough
rlabel pdiffusion 339 -1210 339 -1210 0 cellNo=315
rlabel pdiffusion 346 -1210 346 -1210 0 feedthrough
rlabel pdiffusion 353 -1210 353 -1210 0 cellNo=837
rlabel pdiffusion 360 -1210 360 -1210 0 feedthrough
rlabel pdiffusion 367 -1210 367 -1210 0 feedthrough
rlabel pdiffusion 374 -1210 374 -1210 0 cellNo=211
rlabel pdiffusion 381 -1210 381 -1210 0 feedthrough
rlabel pdiffusion 409 -1210 409 -1210 0 feedthrough
rlabel pdiffusion 423 -1210 423 -1210 0 cellNo=834
rlabel pdiffusion 430 -1210 430 -1210 0 feedthrough
rlabel pdiffusion 24 -1233 24 -1233 0 cellNo=697
rlabel pdiffusion 31 -1233 31 -1233 0 cellNo=797
rlabel pdiffusion 38 -1233 38 -1233 0 feedthrough
rlabel pdiffusion 45 -1233 45 -1233 0 cellNo=398
rlabel pdiffusion 52 -1233 52 -1233 0 feedthrough
rlabel pdiffusion 59 -1233 59 -1233 0 feedthrough
rlabel pdiffusion 66 -1233 66 -1233 0 cellNo=477
rlabel pdiffusion 73 -1233 73 -1233 0 cellNo=761
rlabel pdiffusion 80 -1233 80 -1233 0 feedthrough
rlabel pdiffusion 94 -1233 94 -1233 0 feedthrough
rlabel pdiffusion 101 -1233 101 -1233 0 feedthrough
rlabel pdiffusion 108 -1233 108 -1233 0 cellNo=878
rlabel pdiffusion 115 -1233 115 -1233 0 cellNo=629
rlabel pdiffusion 122 -1233 122 -1233 0 cellNo=881
rlabel pdiffusion 129 -1233 129 -1233 0 cellNo=732
rlabel pdiffusion 136 -1233 136 -1233 0 cellNo=59
rlabel pdiffusion 143 -1233 143 -1233 0 feedthrough
rlabel pdiffusion 150 -1233 150 -1233 0 feedthrough
rlabel pdiffusion 157 -1233 157 -1233 0 cellNo=775
rlabel pdiffusion 164 -1233 164 -1233 0 feedthrough
rlabel pdiffusion 171 -1233 171 -1233 0 cellNo=248
rlabel pdiffusion 178 -1233 178 -1233 0 cellNo=362
rlabel pdiffusion 185 -1233 185 -1233 0 feedthrough
rlabel pdiffusion 192 -1233 192 -1233 0 feedthrough
rlabel pdiffusion 199 -1233 199 -1233 0 cellNo=241
rlabel pdiffusion 206 -1233 206 -1233 0 cellNo=196
rlabel pdiffusion 213 -1233 213 -1233 0 cellNo=740
rlabel pdiffusion 220 -1233 220 -1233 0 cellNo=260
rlabel pdiffusion 227 -1233 227 -1233 0 cellNo=724
rlabel pdiffusion 234 -1233 234 -1233 0 feedthrough
rlabel pdiffusion 241 -1233 241 -1233 0 feedthrough
rlabel pdiffusion 248 -1233 248 -1233 0 cellNo=693
rlabel pdiffusion 255 -1233 255 -1233 0 feedthrough
rlabel pdiffusion 262 -1233 262 -1233 0 cellNo=607
rlabel pdiffusion 269 -1233 269 -1233 0 feedthrough
rlabel pdiffusion 276 -1233 276 -1233 0 feedthrough
rlabel pdiffusion 283 -1233 283 -1233 0 feedthrough
rlabel pdiffusion 290 -1233 290 -1233 0 cellNo=516
rlabel pdiffusion 297 -1233 297 -1233 0 cellNo=802
rlabel pdiffusion 304 -1233 304 -1233 0 feedthrough
rlabel pdiffusion 311 -1233 311 -1233 0 feedthrough
rlabel pdiffusion 318 -1233 318 -1233 0 cellNo=333
rlabel pdiffusion 325 -1233 325 -1233 0 cellNo=108
rlabel pdiffusion 339 -1233 339 -1233 0 feedthrough
rlabel pdiffusion 346 -1233 346 -1233 0 cellNo=758
rlabel pdiffusion 353 -1233 353 -1233 0 feedthrough
rlabel pdiffusion 360 -1233 360 -1233 0 feedthrough
rlabel pdiffusion 367 -1233 367 -1233 0 cellNo=798
rlabel pdiffusion 374 -1233 374 -1233 0 feedthrough
rlabel pdiffusion 402 -1233 402 -1233 0 feedthrough
rlabel pdiffusion 409 -1233 409 -1233 0 cellNo=720
rlabel pdiffusion 416 -1233 416 -1233 0 cellNo=349
rlabel pdiffusion 423 -1233 423 -1233 0 feedthrough
rlabel pdiffusion 430 -1233 430 -1233 0 cellNo=432
rlabel pdiffusion 24 -1258 24 -1258 0 cellNo=61
rlabel pdiffusion 31 -1258 31 -1258 0 feedthrough
rlabel pdiffusion 38 -1258 38 -1258 0 cellNo=512
rlabel pdiffusion 45 -1258 45 -1258 0 cellNo=868
rlabel pdiffusion 59 -1258 59 -1258 0 feedthrough
rlabel pdiffusion 66 -1258 66 -1258 0 cellNo=900
rlabel pdiffusion 73 -1258 73 -1258 0 cellNo=357
rlabel pdiffusion 80 -1258 80 -1258 0 feedthrough
rlabel pdiffusion 101 -1258 101 -1258 0 cellNo=534
rlabel pdiffusion 108 -1258 108 -1258 0 cellNo=870
rlabel pdiffusion 115 -1258 115 -1258 0 feedthrough
rlabel pdiffusion 122 -1258 122 -1258 0 feedthrough
rlabel pdiffusion 129 -1258 129 -1258 0 feedthrough
rlabel pdiffusion 136 -1258 136 -1258 0 cellNo=509
rlabel pdiffusion 143 -1258 143 -1258 0 cellNo=159
rlabel pdiffusion 150 -1258 150 -1258 0 cellNo=793
rlabel pdiffusion 157 -1258 157 -1258 0 cellNo=174
rlabel pdiffusion 164 -1258 164 -1258 0 cellNo=796
rlabel pdiffusion 171 -1258 171 -1258 0 feedthrough
rlabel pdiffusion 178 -1258 178 -1258 0 feedthrough
rlabel pdiffusion 185 -1258 185 -1258 0 cellNo=553
rlabel pdiffusion 192 -1258 192 -1258 0 cellNo=554
rlabel pdiffusion 199 -1258 199 -1258 0 cellNo=296
rlabel pdiffusion 206 -1258 206 -1258 0 cellNo=391
rlabel pdiffusion 213 -1258 213 -1258 0 feedthrough
rlabel pdiffusion 220 -1258 220 -1258 0 cellNo=226
rlabel pdiffusion 227 -1258 227 -1258 0 cellNo=875
rlabel pdiffusion 234 -1258 234 -1258 0 feedthrough
rlabel pdiffusion 241 -1258 241 -1258 0 cellNo=792
rlabel pdiffusion 248 -1258 248 -1258 0 cellNo=659
rlabel pdiffusion 255 -1258 255 -1258 0 cellNo=845
rlabel pdiffusion 262 -1258 262 -1258 0 feedthrough
rlabel pdiffusion 269 -1258 269 -1258 0 feedthrough
rlabel pdiffusion 276 -1258 276 -1258 0 cellNo=842
rlabel pdiffusion 283 -1258 283 -1258 0 cellNo=198
rlabel pdiffusion 290 -1258 290 -1258 0 feedthrough
rlabel pdiffusion 297 -1258 297 -1258 0 cellNo=369
rlabel pdiffusion 304 -1258 304 -1258 0 feedthrough
rlabel pdiffusion 318 -1258 318 -1258 0 cellNo=831
rlabel pdiffusion 325 -1258 325 -1258 0 feedthrough
rlabel pdiffusion 332 -1258 332 -1258 0 cellNo=284
rlabel pdiffusion 339 -1258 339 -1258 0 feedthrough
rlabel pdiffusion 346 -1258 346 -1258 0 cellNo=832
rlabel pdiffusion 353 -1258 353 -1258 0 cellNo=548
rlabel pdiffusion 360 -1258 360 -1258 0 feedthrough
rlabel pdiffusion 367 -1258 367 -1258 0 cellNo=885
rlabel polysilicon 138 -4 138 -4 0 2
rlabel polysilicon 142 -10 142 -10 0 3
rlabel polysilicon 145 -10 145 -10 0 4
rlabel polysilicon 149 -4 149 -4 0 1
rlabel polysilicon 149 -10 149 -10 0 3
rlabel polysilicon 177 -4 177 -4 0 1
rlabel polysilicon 177 -10 177 -10 0 3
rlabel polysilicon 187 -4 187 -4 0 2
rlabel polysilicon 184 -10 184 -10 0 3
rlabel polysilicon 187 -10 187 -10 0 4
rlabel polysilicon 191 -4 191 -4 0 1
rlabel polysilicon 198 -4 198 -4 0 1
rlabel polysilicon 198 -10 198 -10 0 3
rlabel polysilicon 205 -4 205 -4 0 1
rlabel polysilicon 208 -10 208 -10 0 4
rlabel polysilicon 212 -4 212 -4 0 1
rlabel polysilicon 215 -4 215 -4 0 2
rlabel polysilicon 219 -4 219 -4 0 1
rlabel polysilicon 219 -10 219 -10 0 3
rlabel polysilicon 226 -4 226 -4 0 1
rlabel polysilicon 229 -10 229 -10 0 4
rlabel polysilicon 236 -10 236 -10 0 4
rlabel polysilicon 240 -4 240 -4 0 1
rlabel polysilicon 240 -10 240 -10 0 3
rlabel polysilicon 128 -29 128 -29 0 3
rlabel polysilicon 135 -23 135 -23 0 1
rlabel polysilicon 135 -29 135 -29 0 3
rlabel polysilicon 142 -23 142 -23 0 1
rlabel polysilicon 142 -29 142 -29 0 3
rlabel polysilicon 152 -29 152 -29 0 4
rlabel polysilicon 156 -23 156 -23 0 1
rlabel polysilicon 159 -29 159 -29 0 4
rlabel polysilicon 163 -23 163 -23 0 1
rlabel polysilicon 163 -29 163 -29 0 3
rlabel polysilicon 170 -23 170 -23 0 1
rlabel polysilicon 177 -23 177 -23 0 1
rlabel polysilicon 177 -29 177 -29 0 3
rlabel polysilicon 184 -23 184 -23 0 1
rlabel polysilicon 191 -23 191 -23 0 1
rlabel polysilicon 198 -23 198 -23 0 1
rlabel polysilicon 198 -29 198 -29 0 3
rlabel polysilicon 205 -23 205 -23 0 1
rlabel polysilicon 205 -29 205 -29 0 3
rlabel polysilicon 215 -23 215 -23 0 2
rlabel polysilicon 219 -23 219 -23 0 1
rlabel polysilicon 226 -23 226 -23 0 1
rlabel polysilicon 229 -23 229 -23 0 2
rlabel polysilicon 226 -29 226 -29 0 3
rlabel polysilicon 229 -29 229 -29 0 4
rlabel polysilicon 233 -23 233 -23 0 1
rlabel polysilicon 233 -29 233 -29 0 3
rlabel polysilicon 240 -23 240 -23 0 1
rlabel polysilicon 240 -29 240 -29 0 3
rlabel polysilicon 247 -23 247 -23 0 1
rlabel polysilicon 254 -23 254 -23 0 1
rlabel polysilicon 296 -29 296 -29 0 3
rlabel polysilicon 324 -23 324 -23 0 1
rlabel polysilicon 327 -29 327 -29 0 4
rlabel polysilicon 331 -23 331 -23 0 1
rlabel polysilicon 331 -29 331 -29 0 3
rlabel polysilicon 135 -50 135 -50 0 1
rlabel polysilicon 135 -56 135 -56 0 3
rlabel polysilicon 145 -50 145 -50 0 2
rlabel polysilicon 142 -56 142 -56 0 3
rlabel polysilicon 152 -50 152 -50 0 2
rlabel polysilicon 159 -50 159 -50 0 2
rlabel polysilicon 163 -50 163 -50 0 1
rlabel polysilicon 173 -50 173 -50 0 2
rlabel polysilicon 170 -56 170 -56 0 3
rlabel polysilicon 177 -50 177 -50 0 1
rlabel polysilicon 184 -50 184 -50 0 1
rlabel polysilicon 184 -56 184 -56 0 3
rlabel polysilicon 191 -50 191 -50 0 1
rlabel polysilicon 191 -56 191 -56 0 3
rlabel polysilicon 198 -50 198 -50 0 1
rlabel polysilicon 201 -50 201 -50 0 2
rlabel polysilicon 205 -50 205 -50 0 1
rlabel polysilicon 208 -50 208 -50 0 2
rlabel polysilicon 212 -50 212 -50 0 1
rlabel polysilicon 212 -56 212 -56 0 3
rlabel polysilicon 219 -50 219 -50 0 1
rlabel polysilicon 222 -50 222 -50 0 2
rlabel polysilicon 219 -56 219 -56 0 3
rlabel polysilicon 226 -50 226 -50 0 1
rlabel polysilicon 229 -50 229 -50 0 2
rlabel polysilicon 229 -56 229 -56 0 4
rlabel polysilicon 233 -50 233 -50 0 1
rlabel polysilicon 233 -56 233 -56 0 3
rlabel polysilicon 240 -50 240 -50 0 1
rlabel polysilicon 240 -56 240 -56 0 3
rlabel polysilicon 247 -50 247 -50 0 1
rlabel polysilicon 247 -56 247 -56 0 3
rlabel polysilicon 254 -56 254 -56 0 3
rlabel polysilicon 261 -50 261 -50 0 1
rlabel polysilicon 261 -56 261 -56 0 3
rlabel polysilicon 268 -50 268 -50 0 1
rlabel polysilicon 268 -56 268 -56 0 3
rlabel polysilicon 278 -56 278 -56 0 4
rlabel polysilicon 282 -50 282 -50 0 1
rlabel polysilicon 282 -56 282 -56 0 3
rlabel polysilicon 289 -50 289 -50 0 1
rlabel polysilicon 289 -56 289 -56 0 3
rlabel polysilicon 296 -56 296 -56 0 3
rlabel polysilicon 299 -56 299 -56 0 4
rlabel polysilicon 303 -50 303 -50 0 1
rlabel polysilicon 303 -56 303 -56 0 3
rlabel polysilicon 324 -50 324 -50 0 1
rlabel polysilicon 324 -56 324 -56 0 3
rlabel polysilicon 331 -50 331 -50 0 1
rlabel polysilicon 331 -56 331 -56 0 3
rlabel polysilicon 89 -79 89 -79 0 4
rlabel polysilicon 103 -73 103 -73 0 2
rlabel polysilicon 107 -73 107 -73 0 1
rlabel polysilicon 107 -79 107 -79 0 3
rlabel polysilicon 117 -79 117 -79 0 4
rlabel polysilicon 121 -73 121 -73 0 1
rlabel polysilicon 121 -79 121 -79 0 3
rlabel polysilicon 128 -73 128 -73 0 1
rlabel polysilicon 128 -79 128 -79 0 3
rlabel polysilicon 138 -79 138 -79 0 4
rlabel polysilicon 142 -73 142 -73 0 1
rlabel polysilicon 142 -79 142 -79 0 3
rlabel polysilicon 145 -79 145 -79 0 4
rlabel polysilicon 149 -73 149 -73 0 1
rlabel polysilicon 149 -79 149 -79 0 3
rlabel polysilicon 159 -73 159 -73 0 2
rlabel polysilicon 163 -73 163 -73 0 1
rlabel polysilicon 166 -73 166 -73 0 2
rlabel polysilicon 170 -73 170 -73 0 1
rlabel polysilicon 170 -79 170 -79 0 3
rlabel polysilicon 177 -73 177 -73 0 1
rlabel polysilicon 177 -79 177 -79 0 3
rlabel polysilicon 184 -73 184 -73 0 1
rlabel polysilicon 191 -73 191 -73 0 1
rlabel polysilicon 191 -79 191 -79 0 3
rlabel polysilicon 201 -73 201 -73 0 2
rlabel polysilicon 198 -79 198 -79 0 3
rlabel polysilicon 205 -73 205 -73 0 1
rlabel polysilicon 205 -79 205 -79 0 3
rlabel polysilicon 215 -79 215 -79 0 4
rlabel polysilicon 219 -73 219 -73 0 1
rlabel polysilicon 222 -79 222 -79 0 4
rlabel polysilicon 226 -73 226 -73 0 1
rlabel polysilicon 229 -79 229 -79 0 4
rlabel polysilicon 236 -79 236 -79 0 4
rlabel polysilicon 240 -73 240 -73 0 1
rlabel polysilicon 240 -79 240 -79 0 3
rlabel polysilicon 247 -79 247 -79 0 3
rlabel polysilicon 254 -73 254 -73 0 1
rlabel polysilicon 254 -79 254 -79 0 3
rlabel polysilicon 261 -73 261 -73 0 1
rlabel polysilicon 261 -79 261 -79 0 3
rlabel polysilicon 271 -79 271 -79 0 4
rlabel polysilicon 275 -73 275 -73 0 1
rlabel polysilicon 275 -79 275 -79 0 3
rlabel polysilicon 282 -73 282 -73 0 1
rlabel polysilicon 282 -79 282 -79 0 3
rlabel polysilicon 292 -73 292 -73 0 2
rlabel polysilicon 292 -79 292 -79 0 4
rlabel polysilicon 296 -73 296 -73 0 1
rlabel polysilicon 296 -79 296 -79 0 3
rlabel polysilicon 306 -73 306 -73 0 2
rlabel polysilicon 313 -73 313 -73 0 2
rlabel polysilicon 317 -79 317 -79 0 3
rlabel polysilicon 320 -79 320 -79 0 4
rlabel polysilicon 324 -73 324 -73 0 1
rlabel polysilicon 324 -79 324 -79 0 3
rlabel polysilicon 331 -73 331 -73 0 1
rlabel polysilicon 331 -79 331 -79 0 3
rlabel polysilicon 89 -98 89 -98 0 2
rlabel polysilicon 100 -98 100 -98 0 1
rlabel polysilicon 103 -104 103 -104 0 4
rlabel polysilicon 107 -98 107 -98 0 1
rlabel polysilicon 107 -104 107 -104 0 3
rlabel polysilicon 114 -98 114 -98 0 1
rlabel polysilicon 114 -104 114 -104 0 3
rlabel polysilicon 121 -98 121 -98 0 1
rlabel polysilicon 124 -104 124 -104 0 4
rlabel polysilicon 128 -98 128 -98 0 1
rlabel polysilicon 131 -98 131 -98 0 2
rlabel polysilicon 128 -104 128 -104 0 3
rlabel polysilicon 135 -98 135 -98 0 1
rlabel polysilicon 135 -104 135 -104 0 3
rlabel polysilicon 145 -98 145 -98 0 2
rlabel polysilicon 149 -98 149 -98 0 1
rlabel polysilicon 149 -104 149 -104 0 3
rlabel polysilicon 159 -98 159 -98 0 2
rlabel polysilicon 163 -98 163 -98 0 1
rlabel polysilicon 166 -98 166 -98 0 2
rlabel polysilicon 163 -104 163 -104 0 3
rlabel polysilicon 170 -104 170 -104 0 3
rlabel polysilicon 177 -104 177 -104 0 3
rlabel polysilicon 180 -104 180 -104 0 4
rlabel polysilicon 184 -98 184 -98 0 1
rlabel polysilicon 184 -104 184 -104 0 3
rlabel polysilicon 194 -98 194 -98 0 2
rlabel polysilicon 198 -98 198 -98 0 1
rlabel polysilicon 198 -104 198 -104 0 3
rlabel polysilicon 205 -104 205 -104 0 3
rlabel polysilicon 208 -104 208 -104 0 4
rlabel polysilicon 212 -98 212 -98 0 1
rlabel polysilicon 212 -104 212 -104 0 3
rlabel polysilicon 215 -104 215 -104 0 4
rlabel polysilicon 219 -98 219 -98 0 1
rlabel polysilicon 222 -98 222 -98 0 2
rlabel polysilicon 219 -104 219 -104 0 3
rlabel polysilicon 226 -98 226 -98 0 1
rlabel polysilicon 229 -98 229 -98 0 2
rlabel polysilicon 229 -104 229 -104 0 4
rlabel polysilicon 233 -98 233 -98 0 1
rlabel polysilicon 233 -104 233 -104 0 3
rlabel polysilicon 240 -104 240 -104 0 3
rlabel polysilicon 243 -104 243 -104 0 4
rlabel polysilicon 247 -98 247 -98 0 1
rlabel polysilicon 247 -104 247 -104 0 3
rlabel polysilicon 254 -98 254 -98 0 1
rlabel polysilicon 254 -104 254 -104 0 3
rlabel polysilicon 261 -98 261 -98 0 1
rlabel polysilicon 261 -104 261 -104 0 3
rlabel polysilicon 268 -104 268 -104 0 3
rlabel polysilicon 271 -104 271 -104 0 4
rlabel polysilicon 275 -98 275 -98 0 1
rlabel polysilicon 275 -104 275 -104 0 3
rlabel polysilicon 282 -104 282 -104 0 3
rlabel polysilicon 289 -104 289 -104 0 3
rlabel polysilicon 296 -98 296 -98 0 1
rlabel polysilicon 296 -104 296 -104 0 3
rlabel polysilicon 303 -98 303 -98 0 1
rlabel polysilicon 303 -104 303 -104 0 3
rlabel polysilicon 310 -98 310 -98 0 1
rlabel polysilicon 310 -104 310 -104 0 3
rlabel polysilicon 317 -98 317 -98 0 1
rlabel polysilicon 317 -104 317 -104 0 3
rlabel polysilicon 324 -98 324 -98 0 1
rlabel polysilicon 324 -104 324 -104 0 3
rlabel polysilicon 383 -104 383 -104 0 4
rlabel polysilicon 79 -129 79 -129 0 3
rlabel polysilicon 86 -123 86 -123 0 1
rlabel polysilicon 86 -129 86 -129 0 3
rlabel polysilicon 103 -123 103 -123 0 2
rlabel polysilicon 107 -123 107 -123 0 1
rlabel polysilicon 107 -129 107 -129 0 3
rlabel polysilicon 114 -123 114 -123 0 1
rlabel polysilicon 117 -129 117 -129 0 4
rlabel polysilicon 124 -123 124 -123 0 2
rlabel polysilicon 121 -129 121 -129 0 3
rlabel polysilicon 128 -129 128 -129 0 3
rlabel polysilicon 131 -129 131 -129 0 4
rlabel polysilicon 135 -123 135 -123 0 1
rlabel polysilicon 135 -129 135 -129 0 3
rlabel polysilicon 145 -123 145 -123 0 2
rlabel polysilicon 152 -129 152 -129 0 4
rlabel polysilicon 156 -123 156 -123 0 1
rlabel polysilicon 156 -129 156 -129 0 3
rlabel polysilicon 163 -123 163 -123 0 1
rlabel polysilicon 163 -129 163 -129 0 3
rlabel polysilicon 173 -129 173 -129 0 4
rlabel polysilicon 180 -123 180 -123 0 2
rlabel polysilicon 177 -129 177 -129 0 3
rlabel polysilicon 184 -123 184 -123 0 1
rlabel polysilicon 184 -129 184 -129 0 3
rlabel polysilicon 191 -123 191 -123 0 1
rlabel polysilicon 194 -129 194 -129 0 4
rlabel polysilicon 198 -123 198 -123 0 1
rlabel polysilicon 198 -129 198 -129 0 3
rlabel polysilicon 205 -123 205 -123 0 1
rlabel polysilicon 205 -129 205 -129 0 3
rlabel polysilicon 212 -123 212 -123 0 1
rlabel polysilicon 215 -123 215 -123 0 2
rlabel polysilicon 215 -129 215 -129 0 4
rlabel polysilicon 219 -123 219 -123 0 1
rlabel polysilicon 219 -129 219 -129 0 3
rlabel polysilicon 226 -123 226 -123 0 1
rlabel polysilicon 229 -129 229 -129 0 4
rlabel polysilicon 236 -123 236 -123 0 2
rlabel polysilicon 240 -123 240 -123 0 1
rlabel polysilicon 240 -129 240 -129 0 3
rlabel polysilicon 254 -123 254 -123 0 1
rlabel polysilicon 254 -129 254 -129 0 3
rlabel polysilicon 261 -123 261 -123 0 1
rlabel polysilicon 261 -129 261 -129 0 3
rlabel polysilicon 268 -123 268 -123 0 1
rlabel polysilicon 268 -129 268 -129 0 3
rlabel polysilicon 299 -123 299 -123 0 2
rlabel polysilicon 296 -129 296 -129 0 3
rlabel polysilicon 299 -129 299 -129 0 4
rlabel polysilicon 303 -123 303 -123 0 1
rlabel polysilicon 303 -129 303 -129 0 3
rlabel polysilicon 310 -123 310 -123 0 1
rlabel polysilicon 317 -123 317 -123 0 1
rlabel polysilicon 317 -129 317 -129 0 3
rlabel polysilicon 380 -123 380 -123 0 1
rlabel polysilicon 380 -129 380 -129 0 3
rlabel polysilicon 79 -148 79 -148 0 1
rlabel polysilicon 82 -148 82 -148 0 2
rlabel polysilicon 82 -154 82 -154 0 4
rlabel polysilicon 107 -148 107 -148 0 1
rlabel polysilicon 107 -154 107 -154 0 3
rlabel polysilicon 114 -148 114 -148 0 1
rlabel polysilicon 114 -154 114 -154 0 3
rlabel polysilicon 121 -148 121 -148 0 1
rlabel polysilicon 121 -154 121 -154 0 3
rlabel polysilicon 128 -148 128 -148 0 1
rlabel polysilicon 131 -148 131 -148 0 2
rlabel polysilicon 138 -148 138 -148 0 2
rlabel polysilicon 135 -154 135 -154 0 3
rlabel polysilicon 138 -154 138 -154 0 4
rlabel polysilicon 142 -148 142 -148 0 1
rlabel polysilicon 145 -148 145 -148 0 2
rlabel polysilicon 152 -148 152 -148 0 2
rlabel polysilicon 152 -154 152 -154 0 4
rlabel polysilicon 156 -148 156 -148 0 1
rlabel polysilicon 159 -148 159 -148 0 2
rlabel polysilicon 163 -148 163 -148 0 1
rlabel polysilicon 163 -154 163 -154 0 3
rlabel polysilicon 170 -148 170 -148 0 1
rlabel polysilicon 173 -148 173 -148 0 2
rlabel polysilicon 173 -154 173 -154 0 4
rlabel polysilicon 177 -148 177 -148 0 1
rlabel polysilicon 177 -154 177 -154 0 3
rlabel polysilicon 184 -154 184 -154 0 3
rlabel polysilicon 187 -154 187 -154 0 4
rlabel polysilicon 191 -148 191 -148 0 1
rlabel polysilicon 191 -154 191 -154 0 3
rlabel polysilicon 198 -148 198 -148 0 1
rlabel polysilicon 201 -154 201 -154 0 4
rlabel polysilicon 205 -148 205 -148 0 1
rlabel polysilicon 208 -148 208 -148 0 2
rlabel polysilicon 205 -154 205 -154 0 3
rlabel polysilicon 215 -148 215 -148 0 2
rlabel polysilicon 212 -154 212 -154 0 3
rlabel polysilicon 215 -154 215 -154 0 4
rlabel polysilicon 219 -148 219 -148 0 1
rlabel polysilicon 219 -154 219 -154 0 3
rlabel polysilicon 226 -148 226 -148 0 1
rlabel polysilicon 226 -154 226 -154 0 3
rlabel polysilicon 233 -148 233 -148 0 1
rlabel polysilicon 233 -154 233 -154 0 3
rlabel polysilicon 243 -154 243 -154 0 4
rlabel polysilicon 254 -148 254 -148 0 1
rlabel polysilicon 257 -148 257 -148 0 2
rlabel polysilicon 254 -154 254 -154 0 3
rlabel polysilicon 261 -148 261 -148 0 1
rlabel polysilicon 261 -154 261 -154 0 3
rlabel polysilicon 268 -148 268 -148 0 1
rlabel polysilicon 271 -148 271 -148 0 2
rlabel polysilicon 268 -154 268 -154 0 3
rlabel polysilicon 271 -154 271 -154 0 4
rlabel polysilicon 275 -148 275 -148 0 1
rlabel polysilicon 275 -154 275 -154 0 3
rlabel polysilicon 310 -148 310 -148 0 1
rlabel polysilicon 313 -154 313 -154 0 4
rlabel polysilicon 317 -148 317 -148 0 1
rlabel polysilicon 317 -154 317 -154 0 3
rlabel polysilicon 320 -154 320 -154 0 4
rlabel polysilicon 324 -148 324 -148 0 1
rlabel polysilicon 324 -154 324 -154 0 3
rlabel polysilicon 383 -154 383 -154 0 4
rlabel polysilicon 387 -148 387 -148 0 1
rlabel polysilicon 387 -154 387 -154 0 3
rlabel polysilicon 82 -171 82 -171 0 2
rlabel polysilicon 117 -171 117 -171 0 2
rlabel polysilicon 124 -171 124 -171 0 2
rlabel polysilicon 121 -177 121 -177 0 3
rlabel polysilicon 131 -177 131 -177 0 4
rlabel polysilicon 135 -171 135 -171 0 1
rlabel polysilicon 135 -177 135 -177 0 3
rlabel polysilicon 145 -171 145 -171 0 2
rlabel polysilicon 152 -171 152 -171 0 2
rlabel polysilicon 156 -171 156 -171 0 1
rlabel polysilicon 159 -177 159 -177 0 4
rlabel polysilicon 163 -171 163 -171 0 1
rlabel polysilicon 163 -177 163 -177 0 3
rlabel polysilicon 170 -171 170 -171 0 1
rlabel polysilicon 170 -177 170 -177 0 3
rlabel polysilicon 177 -171 177 -171 0 1
rlabel polysilicon 177 -177 177 -177 0 3
rlabel polysilicon 184 -177 184 -177 0 3
rlabel polysilicon 191 -171 191 -171 0 1
rlabel polysilicon 198 -171 198 -171 0 1
rlabel polysilicon 198 -177 198 -177 0 3
rlabel polysilicon 205 -171 205 -171 0 1
rlabel polysilicon 205 -177 205 -177 0 3
rlabel polysilicon 212 -171 212 -171 0 1
rlabel polysilicon 215 -171 215 -171 0 2
rlabel polysilicon 219 -171 219 -171 0 1
rlabel polysilicon 219 -177 219 -177 0 3
rlabel polysilicon 226 -171 226 -171 0 1
rlabel polysilicon 229 -171 229 -171 0 2
rlabel polysilicon 229 -177 229 -177 0 4
rlabel polysilicon 233 -171 233 -171 0 1
rlabel polysilicon 233 -177 233 -177 0 3
rlabel polysilicon 240 -171 240 -171 0 1
rlabel polysilicon 240 -177 240 -177 0 3
rlabel polysilicon 247 -171 247 -171 0 1
rlabel polysilicon 247 -177 247 -177 0 3
rlabel polysilicon 254 -171 254 -171 0 1
rlabel polysilicon 254 -177 254 -177 0 3
rlabel polysilicon 261 -171 261 -171 0 1
rlabel polysilicon 261 -177 261 -177 0 3
rlabel polysilicon 271 -177 271 -177 0 4
rlabel polysilicon 278 -171 278 -171 0 2
rlabel polysilicon 275 -177 275 -177 0 3
rlabel polysilicon 282 -171 282 -171 0 1
rlabel polysilicon 285 -177 285 -177 0 4
rlabel polysilicon 289 -171 289 -171 0 1
rlabel polysilicon 289 -177 289 -177 0 3
rlabel polysilicon 296 -171 296 -171 0 1
rlabel polysilicon 296 -177 296 -177 0 3
rlabel polysilicon 303 -171 303 -171 0 1
rlabel polysilicon 303 -177 303 -177 0 3
rlabel polysilicon 313 -177 313 -177 0 4
rlabel polysilicon 317 -171 317 -171 0 1
rlabel polysilicon 317 -177 317 -177 0 3
rlabel polysilicon 324 -171 324 -171 0 1
rlabel polysilicon 324 -177 324 -177 0 3
rlabel polysilicon 331 -171 331 -171 0 1
rlabel polysilicon 331 -177 331 -177 0 3
rlabel polysilicon 341 -171 341 -171 0 2
rlabel polysilicon 345 -171 345 -171 0 1
rlabel polysilicon 345 -177 345 -177 0 3
rlabel polysilicon 352 -171 352 -171 0 1
rlabel polysilicon 355 -177 355 -177 0 4
rlabel polysilicon 359 -171 359 -171 0 1
rlabel polysilicon 362 -171 362 -171 0 2
rlabel polysilicon 366 -171 366 -171 0 1
rlabel polysilicon 366 -177 366 -177 0 3
rlabel polysilicon 373 -171 373 -171 0 1
rlabel polysilicon 373 -177 373 -177 0 3
rlabel polysilicon 380 -171 380 -171 0 1
rlabel polysilicon 383 -171 383 -171 0 2
rlabel polysilicon 387 -171 387 -171 0 1
rlabel polysilicon 387 -177 387 -177 0 3
rlabel polysilicon 394 -171 394 -171 0 1
rlabel polysilicon 394 -177 394 -177 0 3
rlabel polysilicon 408 -171 408 -171 0 1
rlabel polysilicon 408 -177 408 -177 0 3
rlabel polysilicon 415 -171 415 -171 0 1
rlabel polysilicon 415 -177 415 -177 0 3
rlabel polysilicon 436 -171 436 -171 0 1
rlabel polysilicon 443 -171 443 -171 0 1
rlabel polysilicon 443 -177 443 -177 0 3
rlabel polysilicon 75 -198 75 -198 0 2
rlabel polysilicon 79 -198 79 -198 0 1
rlabel polysilicon 79 -204 79 -204 0 3
rlabel polysilicon 86 -198 86 -198 0 1
rlabel polysilicon 89 -198 89 -198 0 2
rlabel polysilicon 86 -204 86 -204 0 3
rlabel polysilicon 93 -198 93 -198 0 1
rlabel polysilicon 96 -204 96 -204 0 4
rlabel polysilicon 103 -204 103 -204 0 4
rlabel polysilicon 107 -198 107 -198 0 1
rlabel polysilicon 107 -204 107 -204 0 3
rlabel polysilicon 114 -204 114 -204 0 3
rlabel polysilicon 121 -198 121 -198 0 1
rlabel polysilicon 121 -204 121 -204 0 3
rlabel polysilicon 128 -198 128 -198 0 1
rlabel polysilicon 131 -198 131 -198 0 2
rlabel polysilicon 131 -204 131 -204 0 4
rlabel polysilicon 135 -198 135 -198 0 1
rlabel polysilicon 142 -198 142 -198 0 1
rlabel polysilicon 145 -204 145 -204 0 4
rlabel polysilicon 149 -198 149 -198 0 1
rlabel polysilicon 149 -204 149 -204 0 3
rlabel polysilicon 156 -198 156 -198 0 1
rlabel polysilicon 156 -204 156 -204 0 3
rlabel polysilicon 163 -198 163 -198 0 1
rlabel polysilicon 163 -204 163 -204 0 3
rlabel polysilicon 170 -198 170 -198 0 1
rlabel polysilicon 170 -204 170 -204 0 3
rlabel polysilicon 177 -198 177 -198 0 1
rlabel polysilicon 177 -204 177 -204 0 3
rlabel polysilicon 184 -198 184 -198 0 1
rlabel polysilicon 184 -204 184 -204 0 3
rlabel polysilicon 191 -198 191 -198 0 1
rlabel polysilicon 191 -204 191 -204 0 3
rlabel polysilicon 201 -198 201 -198 0 2
rlabel polysilicon 205 -198 205 -198 0 1
rlabel polysilicon 205 -204 205 -204 0 3
rlabel polysilicon 212 -198 212 -198 0 1
rlabel polysilicon 215 -198 215 -198 0 2
rlabel polysilicon 212 -204 212 -204 0 3
rlabel polysilicon 219 -198 219 -198 0 1
rlabel polysilicon 219 -204 219 -204 0 3
rlabel polysilicon 229 -198 229 -198 0 2
rlabel polysilicon 229 -204 229 -204 0 4
rlabel polysilicon 233 -198 233 -198 0 1
rlabel polysilicon 233 -204 233 -204 0 3
rlabel polysilicon 240 -198 240 -198 0 1
rlabel polysilicon 240 -204 240 -204 0 3
rlabel polysilicon 250 -198 250 -198 0 2
rlabel polysilicon 247 -204 247 -204 0 3
rlabel polysilicon 254 -198 254 -198 0 1
rlabel polysilicon 254 -204 254 -204 0 3
rlabel polysilicon 261 -198 261 -198 0 1
rlabel polysilicon 264 -204 264 -204 0 4
rlabel polysilicon 268 -198 268 -198 0 1
rlabel polysilicon 268 -204 268 -204 0 3
rlabel polysilicon 275 -198 275 -198 0 1
rlabel polysilicon 275 -204 275 -204 0 3
rlabel polysilicon 282 -198 282 -198 0 1
rlabel polysilicon 285 -198 285 -198 0 2
rlabel polysilicon 289 -198 289 -198 0 1
rlabel polysilicon 289 -204 289 -204 0 3
rlabel polysilicon 296 -198 296 -198 0 1
rlabel polysilicon 296 -204 296 -204 0 3
rlabel polysilicon 303 -198 303 -198 0 1
rlabel polysilicon 306 -204 306 -204 0 4
rlabel polysilicon 310 -198 310 -198 0 1
rlabel polysilicon 310 -204 310 -204 0 3
rlabel polysilicon 317 -198 317 -198 0 1
rlabel polysilicon 317 -204 317 -204 0 3
rlabel polysilicon 324 -198 324 -198 0 1
rlabel polysilicon 324 -204 324 -204 0 3
rlabel polysilicon 331 -198 331 -198 0 1
rlabel polysilicon 331 -204 331 -204 0 3
rlabel polysilicon 338 -198 338 -198 0 1
rlabel polysilicon 338 -204 338 -204 0 3
rlabel polysilicon 345 -198 345 -198 0 1
rlabel polysilicon 345 -204 345 -204 0 3
rlabel polysilicon 352 -198 352 -198 0 1
rlabel polysilicon 352 -204 352 -204 0 3
rlabel polysilicon 359 -198 359 -198 0 1
rlabel polysilicon 359 -204 359 -204 0 3
rlabel polysilicon 369 -198 369 -198 0 2
rlabel polysilicon 369 -204 369 -204 0 4
rlabel polysilicon 373 -198 373 -198 0 1
rlabel polysilicon 373 -204 373 -204 0 3
rlabel polysilicon 380 -198 380 -198 0 1
rlabel polysilicon 383 -198 383 -198 0 2
rlabel polysilicon 380 -204 380 -204 0 3
rlabel polysilicon 383 -204 383 -204 0 4
rlabel polysilicon 394 -198 394 -198 0 1
rlabel polysilicon 394 -204 394 -204 0 3
rlabel polysilicon 401 -198 401 -198 0 1
rlabel polysilicon 401 -204 401 -204 0 3
rlabel polysilicon 404 -204 404 -204 0 4
rlabel polysilicon 408 -198 408 -198 0 1
rlabel polysilicon 408 -204 408 -204 0 3
rlabel polysilicon 415 -198 415 -198 0 1
rlabel polysilicon 415 -204 415 -204 0 3
rlabel polysilicon 422 -198 422 -198 0 1
rlabel polysilicon 432 -198 432 -198 0 2
rlabel polysilicon 436 -198 436 -198 0 1
rlabel polysilicon 436 -204 436 -204 0 3
rlabel polysilicon 443 -198 443 -198 0 1
rlabel polysilicon 68 -237 68 -237 0 4
rlabel polysilicon 72 -231 72 -231 0 1
rlabel polysilicon 79 -231 79 -231 0 1
rlabel polysilicon 79 -237 79 -237 0 3
rlabel polysilicon 86 -231 86 -231 0 1
rlabel polysilicon 86 -237 86 -237 0 3
rlabel polysilicon 93 -231 93 -231 0 1
rlabel polysilicon 93 -237 93 -237 0 3
rlabel polysilicon 100 -231 100 -231 0 1
rlabel polysilicon 100 -237 100 -237 0 3
rlabel polysilicon 107 -231 107 -231 0 1
rlabel polysilicon 107 -237 107 -237 0 3
rlabel polysilicon 114 -231 114 -231 0 1
rlabel polysilicon 114 -237 114 -237 0 3
rlabel polysilicon 121 -231 121 -231 0 1
rlabel polysilicon 121 -237 121 -237 0 3
rlabel polysilicon 128 -231 128 -231 0 1
rlabel polysilicon 128 -237 128 -237 0 3
rlabel polysilicon 135 -237 135 -237 0 3
rlabel polysilicon 138 -237 138 -237 0 4
rlabel polysilicon 142 -231 142 -231 0 1
rlabel polysilicon 142 -237 142 -237 0 3
rlabel polysilicon 149 -231 149 -231 0 1
rlabel polysilicon 149 -237 149 -237 0 3
rlabel polysilicon 152 -237 152 -237 0 4
rlabel polysilicon 159 -231 159 -231 0 2
rlabel polysilicon 156 -237 156 -237 0 3
rlabel polysilicon 159 -237 159 -237 0 4
rlabel polysilicon 166 -237 166 -237 0 4
rlabel polysilicon 170 -231 170 -231 0 1
rlabel polysilicon 170 -237 170 -237 0 3
rlabel polysilicon 177 -231 177 -231 0 1
rlabel polysilicon 180 -231 180 -231 0 2
rlabel polysilicon 180 -237 180 -237 0 4
rlabel polysilicon 187 -231 187 -231 0 2
rlabel polysilicon 187 -237 187 -237 0 4
rlabel polysilicon 191 -231 191 -231 0 1
rlabel polysilicon 191 -237 191 -237 0 3
rlabel polysilicon 198 -231 198 -231 0 1
rlabel polysilicon 201 -231 201 -231 0 2
rlabel polysilicon 205 -231 205 -231 0 1
rlabel polysilicon 205 -237 205 -237 0 3
rlabel polysilicon 212 -231 212 -231 0 1
rlabel polysilicon 212 -237 212 -237 0 3
rlabel polysilicon 219 -231 219 -231 0 1
rlabel polysilicon 222 -231 222 -231 0 2
rlabel polysilicon 219 -237 219 -237 0 3
rlabel polysilicon 226 -231 226 -231 0 1
rlabel polysilicon 229 -231 229 -231 0 2
rlabel polysilicon 226 -237 226 -237 0 3
rlabel polysilicon 233 -231 233 -231 0 1
rlabel polysilicon 236 -231 236 -231 0 2
rlabel polysilicon 240 -231 240 -231 0 1
rlabel polysilicon 240 -237 240 -237 0 3
rlabel polysilicon 243 -237 243 -237 0 4
rlabel polysilicon 247 -231 247 -231 0 1
rlabel polysilicon 250 -237 250 -237 0 4
rlabel polysilicon 257 -231 257 -231 0 2
rlabel polysilicon 254 -237 254 -237 0 3
rlabel polysilicon 261 -231 261 -231 0 1
rlabel polysilicon 261 -237 261 -237 0 3
rlabel polysilicon 264 -237 264 -237 0 4
rlabel polysilicon 268 -231 268 -231 0 1
rlabel polysilicon 268 -237 268 -237 0 3
rlabel polysilicon 275 -231 275 -231 0 1
rlabel polysilicon 275 -237 275 -237 0 3
rlabel polysilicon 282 -231 282 -231 0 1
rlabel polysilicon 282 -237 282 -237 0 3
rlabel polysilicon 289 -231 289 -231 0 1
rlabel polysilicon 289 -237 289 -237 0 3
rlabel polysilicon 296 -231 296 -231 0 1
rlabel polysilicon 296 -237 296 -237 0 3
rlabel polysilicon 303 -231 303 -231 0 1
rlabel polysilicon 303 -237 303 -237 0 3
rlabel polysilicon 310 -231 310 -231 0 1
rlabel polysilicon 310 -237 310 -237 0 3
rlabel polysilicon 317 -231 317 -231 0 1
rlabel polysilicon 317 -237 317 -237 0 3
rlabel polysilicon 324 -231 324 -231 0 1
rlabel polysilicon 331 -231 331 -231 0 1
rlabel polysilicon 331 -237 331 -237 0 3
rlabel polysilicon 338 -231 338 -231 0 1
rlabel polysilicon 338 -237 338 -237 0 3
rlabel polysilicon 345 -231 345 -231 0 1
rlabel polysilicon 345 -237 345 -237 0 3
rlabel polysilicon 352 -231 352 -231 0 1
rlabel polysilicon 352 -237 352 -237 0 3
rlabel polysilicon 359 -231 359 -231 0 1
rlabel polysilicon 359 -237 359 -237 0 3
rlabel polysilicon 366 -237 366 -237 0 3
rlabel polysilicon 369 -237 369 -237 0 4
rlabel polysilicon 373 -231 373 -231 0 1
rlabel polysilicon 373 -237 373 -237 0 3
rlabel polysilicon 380 -231 380 -231 0 1
rlabel polysilicon 387 -231 387 -231 0 1
rlabel polysilicon 387 -237 387 -237 0 3
rlabel polysilicon 418 -237 418 -237 0 4
rlabel polysilicon 422 -231 422 -231 0 1
rlabel polysilicon 422 -237 422 -237 0 3
rlabel polysilicon 439 -231 439 -231 0 2
rlabel polysilicon 30 -280 30 -280 0 3
rlabel polysilicon 33 -280 33 -280 0 4
rlabel polysilicon 37 -280 37 -280 0 3
rlabel polysilicon 54 -280 54 -280 0 4
rlabel polysilicon 72 -274 72 -274 0 1
rlabel polysilicon 79 -274 79 -274 0 1
rlabel polysilicon 79 -280 79 -280 0 3
rlabel polysilicon 86 -274 86 -274 0 1
rlabel polysilicon 93 -274 93 -274 0 1
rlabel polysilicon 93 -280 93 -280 0 3
rlabel polysilicon 103 -280 103 -280 0 4
rlabel polysilicon 107 -274 107 -274 0 1
rlabel polysilicon 107 -280 107 -280 0 3
rlabel polysilicon 114 -274 114 -274 0 1
rlabel polysilicon 114 -280 114 -280 0 3
rlabel polysilicon 121 -274 121 -274 0 1
rlabel polysilicon 121 -280 121 -280 0 3
rlabel polysilicon 131 -274 131 -274 0 2
rlabel polysilicon 131 -280 131 -280 0 4
rlabel polysilicon 135 -274 135 -274 0 1
rlabel polysilicon 145 -274 145 -274 0 2
rlabel polysilicon 149 -274 149 -274 0 1
rlabel polysilicon 152 -274 152 -274 0 2
rlabel polysilicon 149 -280 149 -280 0 3
rlabel polysilicon 152 -280 152 -280 0 4
rlabel polysilicon 156 -274 156 -274 0 1
rlabel polysilicon 156 -280 156 -280 0 3
rlabel polysilicon 163 -274 163 -274 0 1
rlabel polysilicon 163 -280 163 -280 0 3
rlabel polysilicon 170 -274 170 -274 0 1
rlabel polysilicon 170 -280 170 -280 0 3
rlabel polysilicon 177 -274 177 -274 0 1
rlabel polysilicon 177 -280 177 -280 0 3
rlabel polysilicon 184 -274 184 -274 0 1
rlabel polysilicon 187 -274 187 -274 0 2
rlabel polysilicon 184 -280 184 -280 0 3
rlabel polysilicon 187 -280 187 -280 0 4
rlabel polysilicon 194 -274 194 -274 0 2
rlabel polysilicon 194 -280 194 -280 0 4
rlabel polysilicon 198 -274 198 -274 0 1
rlabel polysilicon 198 -280 198 -280 0 3
rlabel polysilicon 205 -274 205 -274 0 1
rlabel polysilicon 208 -274 208 -274 0 2
rlabel polysilicon 212 -274 212 -274 0 1
rlabel polysilicon 215 -274 215 -274 0 2
rlabel polysilicon 219 -280 219 -280 0 3
rlabel polysilicon 222 -280 222 -280 0 4
rlabel polysilicon 226 -274 226 -274 0 1
rlabel polysilicon 229 -274 229 -274 0 2
rlabel polysilicon 226 -280 226 -280 0 3
rlabel polysilicon 233 -274 233 -274 0 1
rlabel polysilicon 233 -280 233 -280 0 3
rlabel polysilicon 240 -274 240 -274 0 1
rlabel polysilicon 240 -280 240 -280 0 3
rlabel polysilicon 247 -274 247 -274 0 1
rlabel polysilicon 247 -280 247 -280 0 3
rlabel polysilicon 254 -274 254 -274 0 1
rlabel polysilicon 257 -274 257 -274 0 2
rlabel polysilicon 254 -280 254 -280 0 3
rlabel polysilicon 261 -274 261 -274 0 1
rlabel polysilicon 261 -280 261 -280 0 3
rlabel polysilicon 268 -274 268 -274 0 1
rlabel polysilicon 271 -274 271 -274 0 2
rlabel polysilicon 268 -280 268 -280 0 3
rlabel polysilicon 275 -274 275 -274 0 1
rlabel polysilicon 275 -280 275 -280 0 3
rlabel polysilicon 282 -274 282 -274 0 1
rlabel polysilicon 282 -280 282 -280 0 3
rlabel polysilicon 292 -274 292 -274 0 2
rlabel polysilicon 292 -280 292 -280 0 4
rlabel polysilicon 296 -274 296 -274 0 1
rlabel polysilicon 299 -274 299 -274 0 2
rlabel polysilicon 296 -280 296 -280 0 3
rlabel polysilicon 303 -274 303 -274 0 1
rlabel polysilicon 306 -280 306 -280 0 4
rlabel polysilicon 310 -274 310 -274 0 1
rlabel polysilicon 310 -280 310 -280 0 3
rlabel polysilicon 317 -274 317 -274 0 1
rlabel polysilicon 317 -280 317 -280 0 3
rlabel polysilicon 324 -274 324 -274 0 1
rlabel polysilicon 324 -280 324 -280 0 3
rlabel polysilicon 331 -274 331 -274 0 1
rlabel polysilicon 331 -280 331 -280 0 3
rlabel polysilicon 338 -274 338 -274 0 1
rlabel polysilicon 338 -280 338 -280 0 3
rlabel polysilicon 345 -274 345 -274 0 1
rlabel polysilicon 345 -280 345 -280 0 3
rlabel polysilicon 352 -274 352 -274 0 1
rlabel polysilicon 352 -280 352 -280 0 3
rlabel polysilicon 359 -274 359 -274 0 1
rlabel polysilicon 359 -280 359 -280 0 3
rlabel polysilicon 366 -274 366 -274 0 1
rlabel polysilicon 366 -280 366 -280 0 3
rlabel polysilicon 373 -274 373 -274 0 1
rlabel polysilicon 373 -280 373 -280 0 3
rlabel polysilicon 380 -274 380 -274 0 1
rlabel polysilicon 380 -280 380 -280 0 3
rlabel polysilicon 387 -274 387 -274 0 1
rlabel polysilicon 387 -280 387 -280 0 3
rlabel polysilicon 394 -274 394 -274 0 1
rlabel polysilicon 394 -280 394 -280 0 3
rlabel polysilicon 401 -274 401 -274 0 1
rlabel polysilicon 401 -280 401 -280 0 3
rlabel polysilicon 408 -274 408 -274 0 1
rlabel polysilicon 408 -280 408 -280 0 3
rlabel polysilicon 415 -274 415 -274 0 1
rlabel polysilicon 418 -274 418 -274 0 2
rlabel polysilicon 415 -280 415 -280 0 3
rlabel polysilicon 422 -274 422 -274 0 1
rlabel polysilicon 422 -280 422 -280 0 3
rlabel polysilicon 429 -274 429 -274 0 1
rlabel polysilicon 429 -280 429 -280 0 3
rlabel polysilicon 439 -274 439 -274 0 2
rlabel polysilicon 443 -274 443 -274 0 1
rlabel polysilicon 443 -280 443 -280 0 3
rlabel polysilicon 450 -274 450 -274 0 1
rlabel polysilicon 453 -274 453 -274 0 2
rlabel polysilicon 450 -280 450 -280 0 3
rlabel polysilicon 457 -274 457 -274 0 1
rlabel polysilicon 457 -280 457 -280 0 3
rlabel polysilicon 530 -274 530 -274 0 2
rlabel polysilicon 534 -274 534 -274 0 1
rlabel polysilicon 534 -280 534 -280 0 3
rlabel polysilicon 30 -315 30 -315 0 1
rlabel polysilicon 47 -315 47 -315 0 2
rlabel polysilicon 51 -315 51 -315 0 1
rlabel polysilicon 58 -315 58 -315 0 1
rlabel polysilicon 58 -321 58 -321 0 3
rlabel polysilicon 68 -315 68 -315 0 2
rlabel polysilicon 75 -315 75 -315 0 2
rlabel polysilicon 82 -315 82 -315 0 2
rlabel polysilicon 82 -321 82 -321 0 4
rlabel polysilicon 86 -315 86 -315 0 1
rlabel polysilicon 86 -321 86 -321 0 3
rlabel polysilicon 93 -315 93 -315 0 1
rlabel polysilicon 93 -321 93 -321 0 3
rlabel polysilicon 100 -315 100 -315 0 1
rlabel polysilicon 100 -321 100 -321 0 3
rlabel polysilicon 107 -321 107 -321 0 3
rlabel polysilicon 110 -321 110 -321 0 4
rlabel polysilicon 114 -315 114 -315 0 1
rlabel polysilicon 114 -321 114 -321 0 3
rlabel polysilicon 121 -315 121 -315 0 1
rlabel polysilicon 121 -321 121 -321 0 3
rlabel polysilicon 128 -315 128 -315 0 1
rlabel polysilicon 128 -321 128 -321 0 3
rlabel polysilicon 135 -315 135 -315 0 1
rlabel polysilicon 135 -321 135 -321 0 3
rlabel polysilicon 142 -315 142 -315 0 1
rlabel polysilicon 145 -315 145 -315 0 2
rlabel polysilicon 142 -321 142 -321 0 3
rlabel polysilicon 149 -315 149 -315 0 1
rlabel polysilicon 149 -321 149 -321 0 3
rlabel polysilicon 152 -321 152 -321 0 4
rlabel polysilicon 159 -321 159 -321 0 4
rlabel polysilicon 163 -315 163 -315 0 1
rlabel polysilicon 163 -321 163 -321 0 3
rlabel polysilicon 170 -315 170 -315 0 1
rlabel polysilicon 170 -321 170 -321 0 3
rlabel polysilicon 177 -315 177 -315 0 1
rlabel polysilicon 177 -321 177 -321 0 3
rlabel polysilicon 184 -315 184 -315 0 1
rlabel polysilicon 184 -321 184 -321 0 3
rlabel polysilicon 191 -315 191 -315 0 1
rlabel polysilicon 194 -321 194 -321 0 4
rlabel polysilicon 198 -315 198 -315 0 1
rlabel polysilicon 198 -321 198 -321 0 3
rlabel polysilicon 205 -315 205 -315 0 1
rlabel polysilicon 208 -315 208 -315 0 2
rlabel polysilicon 212 -315 212 -315 0 1
rlabel polysilicon 212 -321 212 -321 0 3
rlabel polysilicon 219 -315 219 -315 0 1
rlabel polysilicon 219 -321 219 -321 0 3
rlabel polysilicon 226 -315 226 -315 0 1
rlabel polysilicon 229 -315 229 -315 0 2
rlabel polysilicon 229 -321 229 -321 0 4
rlabel polysilicon 233 -315 233 -315 0 1
rlabel polysilicon 233 -321 233 -321 0 3
rlabel polysilicon 243 -315 243 -315 0 2
rlabel polysilicon 240 -321 240 -321 0 3
rlabel polysilicon 243 -321 243 -321 0 4
rlabel polysilicon 247 -315 247 -315 0 1
rlabel polysilicon 247 -321 247 -321 0 3
rlabel polysilicon 250 -321 250 -321 0 4
rlabel polysilicon 254 -321 254 -321 0 3
rlabel polysilicon 261 -315 261 -315 0 1
rlabel polysilicon 264 -321 264 -321 0 4
rlabel polysilicon 268 -315 268 -315 0 1
rlabel polysilicon 268 -321 268 -321 0 3
rlabel polysilicon 275 -315 275 -315 0 1
rlabel polysilicon 275 -321 275 -321 0 3
rlabel polysilicon 282 -315 282 -315 0 1
rlabel polysilicon 282 -321 282 -321 0 3
rlabel polysilicon 285 -321 285 -321 0 4
rlabel polysilicon 289 -315 289 -315 0 1
rlabel polysilicon 289 -321 289 -321 0 3
rlabel polysilicon 296 -315 296 -315 0 1
rlabel polysilicon 299 -315 299 -315 0 2
rlabel polysilicon 299 -321 299 -321 0 4
rlabel polysilicon 303 -315 303 -315 0 1
rlabel polysilicon 303 -321 303 -321 0 3
rlabel polysilicon 310 -315 310 -315 0 1
rlabel polysilicon 310 -321 310 -321 0 3
rlabel polysilicon 317 -315 317 -315 0 1
rlabel polysilicon 317 -321 317 -321 0 3
rlabel polysilicon 324 -321 324 -321 0 3
rlabel polysilicon 331 -315 331 -315 0 1
rlabel polysilicon 331 -321 331 -321 0 3
rlabel polysilicon 338 -315 338 -315 0 1
rlabel polysilicon 338 -321 338 -321 0 3
rlabel polysilicon 345 -315 345 -315 0 1
rlabel polysilicon 345 -321 345 -321 0 3
rlabel polysilicon 352 -315 352 -315 0 1
rlabel polysilicon 352 -321 352 -321 0 3
rlabel polysilicon 359 -315 359 -315 0 1
rlabel polysilicon 359 -321 359 -321 0 3
rlabel polysilicon 366 -315 366 -315 0 1
rlabel polysilicon 366 -321 366 -321 0 3
rlabel polysilicon 376 -315 376 -315 0 2
rlabel polysilicon 373 -321 373 -321 0 3
rlabel polysilicon 380 -315 380 -315 0 1
rlabel polysilicon 380 -321 380 -321 0 3
rlabel polysilicon 387 -315 387 -315 0 1
rlabel polysilicon 387 -321 387 -321 0 3
rlabel polysilicon 394 -315 394 -315 0 1
rlabel polysilicon 394 -321 394 -321 0 3
rlabel polysilicon 401 -315 401 -315 0 1
rlabel polysilicon 401 -321 401 -321 0 3
rlabel polysilicon 408 -315 408 -315 0 1
rlabel polysilicon 408 -321 408 -321 0 3
rlabel polysilicon 418 -315 418 -315 0 2
rlabel polysilicon 422 -315 422 -315 0 1
rlabel polysilicon 422 -321 422 -321 0 3
rlabel polysilicon 429 -321 429 -321 0 3
rlabel polysilicon 436 -315 436 -315 0 1
rlabel polysilicon 436 -321 436 -321 0 3
rlabel polysilicon 453 -315 453 -315 0 2
rlabel polysilicon 520 -321 520 -321 0 3
rlabel polysilicon 523 -321 523 -321 0 4
rlabel polysilicon 527 -315 527 -315 0 1
rlabel polysilicon 527 -321 527 -321 0 3
rlabel polysilicon 19 -362 19 -362 0 2
rlabel polysilicon 16 -368 16 -368 0 3
rlabel polysilicon 23 -362 23 -362 0 1
rlabel polysilicon 30 -368 30 -368 0 3
rlabel polysilicon 37 -362 37 -362 0 1
rlabel polysilicon 37 -368 37 -368 0 3
rlabel polysilicon 44 -362 44 -362 0 1
rlabel polysilicon 44 -368 44 -368 0 3
rlabel polysilicon 51 -362 51 -362 0 1
rlabel polysilicon 51 -368 51 -368 0 3
rlabel polysilicon 58 -362 58 -362 0 1
rlabel polysilicon 58 -368 58 -368 0 3
rlabel polysilicon 65 -362 65 -362 0 1
rlabel polysilicon 65 -368 65 -368 0 3
rlabel polysilicon 72 -362 72 -362 0 1
rlabel polysilicon 72 -368 72 -368 0 3
rlabel polysilicon 82 -362 82 -362 0 2
rlabel polysilicon 82 -368 82 -368 0 4
rlabel polysilicon 86 -362 86 -362 0 1
rlabel polysilicon 89 -368 89 -368 0 4
rlabel polysilicon 96 -362 96 -362 0 2
rlabel polysilicon 93 -368 93 -368 0 3
rlabel polysilicon 100 -362 100 -362 0 1
rlabel polysilicon 100 -368 100 -368 0 3
rlabel polysilicon 107 -362 107 -362 0 1
rlabel polysilicon 110 -362 110 -362 0 2
rlabel polysilicon 107 -368 107 -368 0 3
rlabel polysilicon 110 -368 110 -368 0 4
rlabel polysilicon 114 -362 114 -362 0 1
rlabel polysilicon 117 -362 117 -362 0 2
rlabel polysilicon 114 -368 114 -368 0 3
rlabel polysilicon 117 -368 117 -368 0 4
rlabel polysilicon 124 -362 124 -362 0 2
rlabel polysilicon 124 -368 124 -368 0 4
rlabel polysilicon 131 -362 131 -362 0 2
rlabel polysilicon 131 -368 131 -368 0 4
rlabel polysilicon 135 -362 135 -362 0 1
rlabel polysilicon 138 -362 138 -362 0 2
rlabel polysilicon 135 -368 135 -368 0 3
rlabel polysilicon 145 -362 145 -362 0 2
rlabel polysilicon 142 -368 142 -368 0 3
rlabel polysilicon 149 -362 149 -362 0 1
rlabel polysilicon 149 -368 149 -368 0 3
rlabel polysilicon 156 -362 156 -362 0 1
rlabel polysilicon 156 -368 156 -368 0 3
rlabel polysilicon 166 -362 166 -362 0 2
rlabel polysilicon 166 -368 166 -368 0 4
rlabel polysilicon 170 -362 170 -362 0 1
rlabel polysilicon 173 -368 173 -368 0 4
rlabel polysilicon 177 -362 177 -362 0 1
rlabel polysilicon 177 -368 177 -368 0 3
rlabel polysilicon 184 -362 184 -362 0 1
rlabel polysilicon 184 -368 184 -368 0 3
rlabel polysilicon 194 -362 194 -362 0 2
rlabel polysilicon 191 -368 191 -368 0 3
rlabel polysilicon 198 -362 198 -362 0 1
rlabel polysilicon 201 -362 201 -362 0 2
rlabel polysilicon 205 -362 205 -362 0 1
rlabel polysilicon 205 -368 205 -368 0 3
rlabel polysilicon 212 -362 212 -362 0 1
rlabel polysilicon 215 -362 215 -362 0 2
rlabel polysilicon 212 -368 212 -368 0 3
rlabel polysilicon 219 -362 219 -362 0 1
rlabel polysilicon 219 -368 219 -368 0 3
rlabel polysilicon 226 -362 226 -362 0 1
rlabel polysilicon 226 -368 226 -368 0 3
rlabel polysilicon 233 -362 233 -362 0 1
rlabel polysilicon 233 -368 233 -368 0 3
rlabel polysilicon 240 -362 240 -362 0 1
rlabel polysilicon 243 -362 243 -362 0 2
rlabel polysilicon 240 -368 240 -368 0 3
rlabel polysilicon 243 -368 243 -368 0 4
rlabel polysilicon 250 -362 250 -362 0 2
rlabel polysilicon 247 -368 247 -368 0 3
rlabel polysilicon 250 -368 250 -368 0 4
rlabel polysilicon 254 -368 254 -368 0 3
rlabel polysilicon 261 -362 261 -362 0 1
rlabel polysilicon 264 -362 264 -362 0 2
rlabel polysilicon 261 -368 261 -368 0 3
rlabel polysilicon 271 -362 271 -362 0 2
rlabel polysilicon 268 -368 268 -368 0 3
rlabel polysilicon 271 -368 271 -368 0 4
rlabel polysilicon 275 -368 275 -368 0 3
rlabel polysilicon 278 -368 278 -368 0 4
rlabel polysilicon 285 -362 285 -362 0 2
rlabel polysilicon 282 -368 282 -368 0 3
rlabel polysilicon 289 -362 289 -362 0 1
rlabel polysilicon 289 -368 289 -368 0 3
rlabel polysilicon 296 -362 296 -362 0 1
rlabel polysilicon 296 -368 296 -368 0 3
rlabel polysilicon 306 -362 306 -362 0 2
rlabel polysilicon 310 -362 310 -362 0 1
rlabel polysilicon 310 -368 310 -368 0 3
rlabel polysilicon 317 -368 317 -368 0 3
rlabel polysilicon 320 -368 320 -368 0 4
rlabel polysilicon 324 -362 324 -362 0 1
rlabel polysilicon 327 -362 327 -362 0 2
rlabel polysilicon 324 -368 324 -368 0 3
rlabel polysilicon 331 -362 331 -362 0 1
rlabel polysilicon 331 -368 331 -368 0 3
rlabel polysilicon 338 -362 338 -362 0 1
rlabel polysilicon 338 -368 338 -368 0 3
rlabel polysilicon 345 -362 345 -362 0 1
rlabel polysilicon 345 -368 345 -368 0 3
rlabel polysilicon 352 -362 352 -362 0 1
rlabel polysilicon 352 -368 352 -368 0 3
rlabel polysilicon 359 -362 359 -362 0 1
rlabel polysilicon 359 -368 359 -368 0 3
rlabel polysilicon 366 -362 366 -362 0 1
rlabel polysilicon 366 -368 366 -368 0 3
rlabel polysilicon 373 -362 373 -362 0 1
rlabel polysilicon 373 -368 373 -368 0 3
rlabel polysilicon 380 -362 380 -362 0 1
rlabel polysilicon 380 -368 380 -368 0 3
rlabel polysilicon 390 -362 390 -362 0 2
rlabel polysilicon 387 -368 387 -368 0 3
rlabel polysilicon 390 -368 390 -368 0 4
rlabel polysilicon 394 -362 394 -362 0 1
rlabel polysilicon 394 -368 394 -368 0 3
rlabel polysilicon 401 -362 401 -362 0 1
rlabel polysilicon 401 -368 401 -368 0 3
rlabel polysilicon 408 -362 408 -362 0 1
rlabel polysilicon 408 -368 408 -368 0 3
rlabel polysilicon 415 -362 415 -362 0 1
rlabel polysilicon 415 -368 415 -368 0 3
rlabel polysilicon 422 -362 422 -362 0 1
rlabel polysilicon 422 -368 422 -368 0 3
rlabel polysilicon 429 -362 429 -362 0 1
rlabel polysilicon 429 -368 429 -368 0 3
rlabel polysilicon 436 -362 436 -362 0 1
rlabel polysilicon 436 -368 436 -368 0 3
rlabel polysilicon 443 -362 443 -362 0 1
rlabel polysilicon 443 -368 443 -368 0 3
rlabel polysilicon 450 -362 450 -362 0 1
rlabel polysilicon 450 -368 450 -368 0 3
rlabel polysilicon 457 -362 457 -362 0 1
rlabel polysilicon 457 -368 457 -368 0 3
rlabel polysilicon 467 -362 467 -362 0 2
rlabel polysilicon 471 -362 471 -362 0 1
rlabel polysilicon 471 -368 471 -368 0 3
rlabel polysilicon 513 -362 513 -362 0 1
rlabel polysilicon 513 -368 513 -368 0 3
rlabel polysilicon 16 -413 16 -413 0 1
rlabel polysilicon 23 -413 23 -413 0 1
rlabel polysilicon 23 -419 23 -419 0 3
rlabel polysilicon 30 -413 30 -413 0 1
rlabel polysilicon 30 -419 30 -419 0 3
rlabel polysilicon 37 -413 37 -413 0 1
rlabel polysilicon 44 -413 44 -413 0 1
rlabel polysilicon 51 -419 51 -419 0 3
rlabel polysilicon 58 -413 58 -413 0 1
rlabel polysilicon 65 -413 65 -413 0 1
rlabel polysilicon 72 -413 72 -413 0 1
rlabel polysilicon 72 -419 72 -419 0 3
rlabel polysilicon 79 -413 79 -413 0 1
rlabel polysilicon 79 -419 79 -419 0 3
rlabel polysilicon 86 -413 86 -413 0 1
rlabel polysilicon 86 -419 86 -419 0 3
rlabel polysilicon 93 -413 93 -413 0 1
rlabel polysilicon 93 -419 93 -419 0 3
rlabel polysilicon 100 -413 100 -413 0 1
rlabel polysilicon 103 -413 103 -413 0 2
rlabel polysilicon 107 -413 107 -413 0 1
rlabel polysilicon 110 -413 110 -413 0 2
rlabel polysilicon 110 -419 110 -419 0 4
rlabel polysilicon 114 -413 114 -413 0 1
rlabel polysilicon 114 -419 114 -419 0 3
rlabel polysilicon 121 -413 121 -413 0 1
rlabel polysilicon 121 -419 121 -419 0 3
rlabel polysilicon 128 -413 128 -413 0 1
rlabel polysilicon 128 -419 128 -419 0 3
rlabel polysilicon 138 -413 138 -413 0 2
rlabel polysilicon 142 -419 142 -419 0 3
rlabel polysilicon 145 -419 145 -419 0 4
rlabel polysilicon 152 -413 152 -413 0 2
rlabel polysilicon 156 -413 156 -413 0 1
rlabel polysilicon 159 -413 159 -413 0 2
rlabel polysilicon 166 -413 166 -413 0 2
rlabel polysilicon 170 -413 170 -413 0 1
rlabel polysilicon 170 -419 170 -419 0 3
rlabel polysilicon 177 -413 177 -413 0 1
rlabel polysilicon 177 -419 177 -419 0 3
rlabel polysilicon 184 -413 184 -413 0 1
rlabel polysilicon 191 -413 191 -413 0 1
rlabel polysilicon 194 -413 194 -413 0 2
rlabel polysilicon 198 -413 198 -413 0 1
rlabel polysilicon 198 -419 198 -419 0 3
rlabel polysilicon 208 -413 208 -413 0 2
rlabel polysilicon 212 -413 212 -413 0 1
rlabel polysilicon 215 -413 215 -413 0 2
rlabel polysilicon 215 -419 215 -419 0 4
rlabel polysilicon 219 -413 219 -413 0 1
rlabel polysilicon 219 -419 219 -419 0 3
rlabel polysilicon 226 -413 226 -413 0 1
rlabel polysilicon 229 -413 229 -413 0 2
rlabel polysilicon 226 -419 226 -419 0 3
rlabel polysilicon 229 -419 229 -419 0 4
rlabel polysilicon 233 -413 233 -413 0 1
rlabel polysilicon 233 -419 233 -419 0 3
rlabel polysilicon 240 -413 240 -413 0 1
rlabel polysilicon 240 -419 240 -419 0 3
rlabel polysilicon 247 -413 247 -413 0 1
rlabel polysilicon 247 -419 247 -419 0 3
rlabel polysilicon 254 -413 254 -413 0 1
rlabel polysilicon 254 -419 254 -419 0 3
rlabel polysilicon 261 -413 261 -413 0 1
rlabel polysilicon 261 -419 261 -419 0 3
rlabel polysilicon 264 -419 264 -419 0 4
rlabel polysilicon 268 -413 268 -413 0 1
rlabel polysilicon 275 -413 275 -413 0 1
rlabel polysilicon 275 -419 275 -419 0 3
rlabel polysilicon 282 -413 282 -413 0 1
rlabel polysilicon 285 -419 285 -419 0 4
rlabel polysilicon 289 -413 289 -413 0 1
rlabel polysilicon 289 -419 289 -419 0 3
rlabel polysilicon 296 -413 296 -413 0 1
rlabel polysilicon 296 -419 296 -419 0 3
rlabel polysilicon 303 -413 303 -413 0 1
rlabel polysilicon 303 -419 303 -419 0 3
rlabel polysilicon 310 -413 310 -413 0 1
rlabel polysilicon 313 -413 313 -413 0 2
rlabel polysilicon 317 -413 317 -413 0 1
rlabel polysilicon 320 -419 320 -419 0 4
rlabel polysilicon 324 -413 324 -413 0 1
rlabel polysilicon 327 -413 327 -413 0 2
rlabel polysilicon 324 -419 324 -419 0 3
rlabel polysilicon 327 -419 327 -419 0 4
rlabel polysilicon 331 -413 331 -413 0 1
rlabel polysilicon 331 -419 331 -419 0 3
rlabel polysilicon 341 -419 341 -419 0 4
rlabel polysilicon 348 -413 348 -413 0 2
rlabel polysilicon 352 -413 352 -413 0 1
rlabel polysilicon 352 -419 352 -419 0 3
rlabel polysilicon 359 -413 359 -413 0 1
rlabel polysilicon 359 -419 359 -419 0 3
rlabel polysilicon 366 -413 366 -413 0 1
rlabel polysilicon 366 -419 366 -419 0 3
rlabel polysilicon 373 -413 373 -413 0 1
rlabel polysilicon 373 -419 373 -419 0 3
rlabel polysilicon 380 -413 380 -413 0 1
rlabel polysilicon 380 -419 380 -419 0 3
rlabel polysilicon 387 -413 387 -413 0 1
rlabel polysilicon 387 -419 387 -419 0 3
rlabel polysilicon 394 -413 394 -413 0 1
rlabel polysilicon 394 -419 394 -419 0 3
rlabel polysilicon 397 -419 397 -419 0 4
rlabel polysilicon 401 -413 401 -413 0 1
rlabel polysilicon 401 -419 401 -419 0 3
rlabel polysilicon 408 -413 408 -413 0 1
rlabel polysilicon 408 -419 408 -419 0 3
rlabel polysilicon 415 -413 415 -413 0 1
rlabel polysilicon 418 -413 418 -413 0 2
rlabel polysilicon 415 -419 415 -419 0 3
rlabel polysilicon 422 -413 422 -413 0 1
rlabel polysilicon 422 -419 422 -419 0 3
rlabel polysilicon 429 -413 429 -413 0 1
rlabel polysilicon 429 -419 429 -419 0 3
rlabel polysilicon 436 -413 436 -413 0 1
rlabel polysilicon 436 -419 436 -419 0 3
rlabel polysilicon 443 -413 443 -413 0 1
rlabel polysilicon 443 -419 443 -419 0 3
rlabel polysilicon 450 -413 450 -413 0 1
rlabel polysilicon 450 -419 450 -419 0 3
rlabel polysilicon 457 -413 457 -413 0 1
rlabel polysilicon 457 -419 457 -419 0 3
rlabel polysilicon 464 -413 464 -413 0 1
rlabel polysilicon 464 -419 464 -419 0 3
rlabel polysilicon 471 -413 471 -413 0 1
rlabel polysilicon 471 -419 471 -419 0 3
rlabel polysilicon 481 -413 481 -413 0 2
rlabel polysilicon 485 -419 485 -419 0 3
rlabel polysilicon 492 -413 492 -413 0 1
rlabel polysilicon 492 -419 492 -419 0 3
rlabel polysilicon 499 -413 499 -413 0 1
rlabel polysilicon 499 -419 499 -419 0 3
rlabel polysilicon 506 -413 506 -413 0 1
rlabel polysilicon 506 -419 506 -419 0 3
rlabel polysilicon 513 -413 513 -413 0 1
rlabel polysilicon 513 -419 513 -419 0 3
rlabel polysilicon 520 -413 520 -413 0 1
rlabel polysilicon 520 -419 520 -419 0 3
rlabel polysilicon 527 -413 527 -413 0 1
rlabel polysilicon 527 -419 527 -419 0 3
rlabel polysilicon 2 -464 2 -464 0 1
rlabel polysilicon 2 -470 2 -470 0 3
rlabel polysilicon 9 -464 9 -464 0 1
rlabel polysilicon 9 -470 9 -470 0 3
rlabel polysilicon 16 -464 16 -464 0 1
rlabel polysilicon 16 -470 16 -470 0 3
rlabel polysilicon 23 -470 23 -470 0 3
rlabel polysilicon 30 -464 30 -464 0 1
rlabel polysilicon 37 -464 37 -464 0 1
rlabel polysilicon 37 -470 37 -470 0 3
rlabel polysilicon 44 -464 44 -464 0 1
rlabel polysilicon 44 -470 44 -470 0 3
rlabel polysilicon 54 -464 54 -464 0 2
rlabel polysilicon 54 -470 54 -470 0 4
rlabel polysilicon 58 -464 58 -464 0 1
rlabel polysilicon 58 -470 58 -470 0 3
rlabel polysilicon 65 -464 65 -464 0 1
rlabel polysilicon 65 -470 65 -470 0 3
rlabel polysilicon 72 -464 72 -464 0 1
rlabel polysilicon 72 -470 72 -470 0 3
rlabel polysilicon 79 -464 79 -464 0 1
rlabel polysilicon 79 -470 79 -470 0 3
rlabel polysilicon 86 -464 86 -464 0 1
rlabel polysilicon 86 -470 86 -470 0 3
rlabel polysilicon 96 -464 96 -464 0 2
rlabel polysilicon 93 -470 93 -470 0 3
rlabel polysilicon 96 -470 96 -470 0 4
rlabel polysilicon 100 -464 100 -464 0 1
rlabel polysilicon 100 -470 100 -470 0 3
rlabel polysilicon 107 -464 107 -464 0 1
rlabel polysilicon 107 -470 107 -470 0 3
rlabel polysilicon 114 -470 114 -470 0 3
rlabel polysilicon 121 -464 121 -464 0 1
rlabel polysilicon 121 -470 121 -470 0 3
rlabel polysilicon 124 -470 124 -470 0 4
rlabel polysilicon 128 -470 128 -470 0 3
rlabel polysilicon 131 -470 131 -470 0 4
rlabel polysilicon 135 -464 135 -464 0 1
rlabel polysilicon 135 -470 135 -470 0 3
rlabel polysilicon 142 -464 142 -464 0 1
rlabel polysilicon 142 -470 142 -470 0 3
rlabel polysilicon 149 -470 149 -470 0 3
rlabel polysilicon 152 -470 152 -470 0 4
rlabel polysilicon 159 -464 159 -464 0 2
rlabel polysilicon 156 -470 156 -470 0 3
rlabel polysilicon 166 -464 166 -464 0 2
rlabel polysilicon 163 -470 163 -470 0 3
rlabel polysilicon 170 -464 170 -464 0 1
rlabel polysilicon 173 -464 173 -464 0 2
rlabel polysilicon 170 -470 170 -470 0 3
rlabel polysilicon 177 -464 177 -464 0 1
rlabel polysilicon 177 -470 177 -470 0 3
rlabel polysilicon 184 -470 184 -470 0 3
rlabel polysilicon 191 -464 191 -464 0 1
rlabel polysilicon 191 -470 191 -470 0 3
rlabel polysilicon 198 -464 198 -464 0 1
rlabel polysilicon 201 -464 201 -464 0 2
rlabel polysilicon 201 -470 201 -470 0 4
rlabel polysilicon 205 -464 205 -464 0 1
rlabel polysilicon 205 -470 205 -470 0 3
rlabel polysilicon 212 -464 212 -464 0 1
rlabel polysilicon 212 -470 212 -470 0 3
rlabel polysilicon 219 -464 219 -464 0 1
rlabel polysilicon 222 -464 222 -464 0 2
rlabel polysilicon 219 -470 219 -470 0 3
rlabel polysilicon 229 -464 229 -464 0 2
rlabel polysilicon 229 -470 229 -470 0 4
rlabel polysilicon 233 -464 233 -464 0 1
rlabel polysilicon 233 -470 233 -470 0 3
rlabel polysilicon 240 -464 240 -464 0 1
rlabel polysilicon 243 -464 243 -464 0 2
rlabel polysilicon 240 -470 240 -470 0 3
rlabel polysilicon 247 -464 247 -464 0 1
rlabel polysilicon 247 -470 247 -470 0 3
rlabel polysilicon 254 -464 254 -464 0 1
rlabel polysilicon 261 -470 261 -470 0 3
rlabel polysilicon 264 -470 264 -470 0 4
rlabel polysilicon 268 -464 268 -464 0 1
rlabel polysilicon 268 -470 268 -470 0 3
rlabel polysilicon 275 -464 275 -464 0 1
rlabel polysilicon 278 -464 278 -464 0 2
rlabel polysilicon 278 -470 278 -470 0 4
rlabel polysilicon 282 -464 282 -464 0 1
rlabel polysilicon 285 -464 285 -464 0 2
rlabel polysilicon 282 -470 282 -470 0 3
rlabel polysilicon 285 -470 285 -470 0 4
rlabel polysilicon 289 -464 289 -464 0 1
rlabel polysilicon 289 -470 289 -470 0 3
rlabel polysilicon 296 -464 296 -464 0 1
rlabel polysilicon 296 -470 296 -470 0 3
rlabel polysilicon 303 -464 303 -464 0 1
rlabel polysilicon 303 -470 303 -470 0 3
rlabel polysilicon 313 -464 313 -464 0 2
rlabel polysilicon 310 -470 310 -470 0 3
rlabel polysilicon 313 -470 313 -470 0 4
rlabel polysilicon 317 -470 317 -470 0 3
rlabel polysilicon 320 -470 320 -470 0 4
rlabel polysilicon 324 -464 324 -464 0 1
rlabel polysilicon 324 -470 324 -470 0 3
rlabel polysilicon 331 -464 331 -464 0 1
rlabel polysilicon 331 -470 331 -470 0 3
rlabel polysilicon 338 -464 338 -464 0 1
rlabel polysilicon 338 -470 338 -470 0 3
rlabel polysilicon 345 -464 345 -464 0 1
rlabel polysilicon 348 -464 348 -464 0 2
rlabel polysilicon 352 -464 352 -464 0 1
rlabel polysilicon 359 -464 359 -464 0 1
rlabel polysilicon 359 -470 359 -470 0 3
rlabel polysilicon 366 -470 366 -470 0 3
rlabel polysilicon 373 -470 373 -470 0 3
rlabel polysilicon 380 -464 380 -464 0 1
rlabel polysilicon 380 -470 380 -470 0 3
rlabel polysilicon 387 -464 387 -464 0 1
rlabel polysilicon 387 -470 387 -470 0 3
rlabel polysilicon 394 -464 394 -464 0 1
rlabel polysilicon 397 -464 397 -464 0 2
rlabel polysilicon 394 -470 394 -470 0 3
rlabel polysilicon 401 -464 401 -464 0 1
rlabel polysilicon 401 -470 401 -470 0 3
rlabel polysilicon 408 -464 408 -464 0 1
rlabel polysilicon 408 -470 408 -470 0 3
rlabel polysilicon 415 -464 415 -464 0 1
rlabel polysilicon 415 -470 415 -470 0 3
rlabel polysilicon 422 -464 422 -464 0 1
rlabel polysilicon 422 -470 422 -470 0 3
rlabel polysilicon 429 -464 429 -464 0 1
rlabel polysilicon 429 -470 429 -470 0 3
rlabel polysilicon 436 -464 436 -464 0 1
rlabel polysilicon 436 -470 436 -470 0 3
rlabel polysilicon 443 -464 443 -464 0 1
rlabel polysilicon 443 -470 443 -470 0 3
rlabel polysilicon 450 -464 450 -464 0 1
rlabel polysilicon 450 -470 450 -470 0 3
rlabel polysilicon 457 -464 457 -464 0 1
rlabel polysilicon 457 -470 457 -470 0 3
rlabel polysilicon 464 -464 464 -464 0 1
rlabel polysilicon 464 -470 464 -470 0 3
rlabel polysilicon 471 -464 471 -464 0 1
rlabel polysilicon 471 -470 471 -470 0 3
rlabel polysilicon 478 -464 478 -464 0 1
rlabel polysilicon 478 -470 478 -470 0 3
rlabel polysilicon 485 -464 485 -464 0 1
rlabel polysilicon 485 -470 485 -470 0 3
rlabel polysilicon 492 -464 492 -464 0 1
rlabel polysilicon 492 -470 492 -470 0 3
rlabel polysilicon 499 -464 499 -464 0 1
rlabel polysilicon 499 -470 499 -470 0 3
rlabel polysilicon 506 -464 506 -464 0 1
rlabel polysilicon 506 -470 506 -470 0 3
rlabel polysilicon 513 -464 513 -464 0 1
rlabel polysilicon 513 -470 513 -470 0 3
rlabel polysilicon 520 -464 520 -464 0 1
rlabel polysilicon 520 -470 520 -470 0 3
rlabel polysilicon 527 -464 527 -464 0 1
rlabel polysilicon 527 -470 527 -470 0 3
rlabel polysilicon 534 -464 534 -464 0 1
rlabel polysilicon 534 -470 534 -470 0 3
rlabel polysilicon 541 -464 541 -464 0 1
rlabel polysilicon 541 -470 541 -470 0 3
rlabel polysilicon 548 -464 548 -464 0 1
rlabel polysilicon 548 -470 548 -470 0 3
rlabel polysilicon 555 -470 555 -470 0 3
rlabel polysilicon 558 -470 558 -470 0 4
rlabel polysilicon 562 -464 562 -464 0 1
rlabel polysilicon 562 -470 562 -470 0 3
rlabel polysilicon 572 -470 572 -470 0 4
rlabel polysilicon 576 -464 576 -464 0 1
rlabel polysilicon 576 -470 576 -470 0 3
rlabel polysilicon 16 -521 16 -521 0 1
rlabel polysilicon 16 -527 16 -527 0 3
rlabel polysilicon 23 -521 23 -521 0 1
rlabel polysilicon 23 -527 23 -527 0 3
rlabel polysilicon 30 -521 30 -521 0 1
rlabel polysilicon 30 -527 30 -527 0 3
rlabel polysilicon 37 -521 37 -521 0 1
rlabel polysilicon 37 -527 37 -527 0 3
rlabel polysilicon 44 -521 44 -521 0 1
rlabel polysilicon 44 -527 44 -527 0 3
rlabel polysilicon 51 -521 51 -521 0 1
rlabel polysilicon 51 -527 51 -527 0 3
rlabel polysilicon 58 -521 58 -521 0 1
rlabel polysilicon 58 -527 58 -527 0 3
rlabel polysilicon 65 -521 65 -521 0 1
rlabel polysilicon 68 -527 68 -527 0 4
rlabel polysilicon 75 -521 75 -521 0 2
rlabel polysilicon 75 -527 75 -527 0 4
rlabel polysilicon 79 -521 79 -521 0 1
rlabel polysilicon 82 -521 82 -521 0 2
rlabel polysilicon 86 -521 86 -521 0 1
rlabel polysilicon 89 -521 89 -521 0 2
rlabel polysilicon 89 -527 89 -527 0 4
rlabel polysilicon 93 -521 93 -521 0 1
rlabel polysilicon 93 -527 93 -527 0 3
rlabel polysilicon 100 -521 100 -521 0 1
rlabel polysilicon 100 -527 100 -527 0 3
rlabel polysilicon 107 -521 107 -521 0 1
rlabel polysilicon 107 -527 107 -527 0 3
rlabel polysilicon 117 -521 117 -521 0 2
rlabel polysilicon 114 -527 114 -527 0 3
rlabel polysilicon 124 -521 124 -521 0 2
rlabel polysilicon 121 -527 121 -527 0 3
rlabel polysilicon 124 -527 124 -527 0 4
rlabel polysilicon 128 -527 128 -527 0 3
rlabel polysilicon 131 -527 131 -527 0 4
rlabel polysilicon 138 -527 138 -527 0 4
rlabel polysilicon 145 -527 145 -527 0 4
rlabel polysilicon 149 -521 149 -521 0 1
rlabel polysilicon 149 -527 149 -527 0 3
rlabel polysilicon 159 -521 159 -521 0 2
rlabel polysilicon 156 -527 156 -527 0 3
rlabel polysilicon 159 -527 159 -527 0 4
rlabel polysilicon 163 -521 163 -521 0 1
rlabel polysilicon 163 -527 163 -527 0 3
rlabel polysilicon 170 -521 170 -521 0 1
rlabel polysilicon 170 -527 170 -527 0 3
rlabel polysilicon 177 -521 177 -521 0 1
rlabel polysilicon 177 -527 177 -527 0 3
rlabel polysilicon 184 -521 184 -521 0 1
rlabel polysilicon 187 -527 187 -527 0 4
rlabel polysilicon 191 -521 191 -521 0 1
rlabel polysilicon 191 -527 191 -527 0 3
rlabel polysilicon 201 -521 201 -521 0 2
rlabel polysilicon 201 -527 201 -527 0 4
rlabel polysilicon 205 -521 205 -521 0 1
rlabel polysilicon 205 -527 205 -527 0 3
rlabel polysilicon 212 -521 212 -521 0 1
rlabel polysilicon 212 -527 212 -527 0 3
rlabel polysilicon 219 -521 219 -521 0 1
rlabel polysilicon 222 -521 222 -521 0 2
rlabel polysilicon 219 -527 219 -527 0 3
rlabel polysilicon 226 -521 226 -521 0 1
rlabel polysilicon 229 -521 229 -521 0 2
rlabel polysilicon 226 -527 226 -527 0 3
rlabel polysilicon 233 -521 233 -521 0 1
rlabel polysilicon 233 -527 233 -527 0 3
rlabel polysilicon 240 -521 240 -521 0 1
rlabel polysilicon 243 -521 243 -521 0 2
rlabel polysilicon 240 -527 240 -527 0 3
rlabel polysilicon 247 -521 247 -521 0 1
rlabel polysilicon 247 -527 247 -527 0 3
rlabel polysilicon 254 -521 254 -521 0 1
rlabel polysilicon 254 -527 254 -527 0 3
rlabel polysilicon 261 -521 261 -521 0 1
rlabel polysilicon 264 -521 264 -521 0 2
rlabel polysilicon 261 -527 261 -527 0 3
rlabel polysilicon 264 -527 264 -527 0 4
rlabel polysilicon 268 -521 268 -521 0 1
rlabel polysilicon 268 -527 268 -527 0 3
rlabel polysilicon 275 -521 275 -521 0 1
rlabel polysilicon 278 -527 278 -527 0 4
rlabel polysilicon 282 -521 282 -521 0 1
rlabel polysilicon 285 -521 285 -521 0 2
rlabel polysilicon 285 -527 285 -527 0 4
rlabel polysilicon 289 -521 289 -521 0 1
rlabel polysilicon 292 -521 292 -521 0 2
rlabel polysilicon 292 -527 292 -527 0 4
rlabel polysilicon 296 -521 296 -521 0 1
rlabel polysilicon 299 -521 299 -521 0 2
rlabel polysilicon 299 -527 299 -527 0 4
rlabel polysilicon 303 -521 303 -521 0 1
rlabel polysilicon 303 -527 303 -527 0 3
rlabel polysilicon 310 -521 310 -521 0 1
rlabel polysilicon 310 -527 310 -527 0 3
rlabel polysilicon 313 -527 313 -527 0 4
rlabel polysilicon 317 -521 317 -521 0 1
rlabel polysilicon 317 -527 317 -527 0 3
rlabel polysilicon 324 -527 324 -527 0 3
rlabel polysilicon 331 -521 331 -521 0 1
rlabel polysilicon 331 -527 331 -527 0 3
rlabel polysilicon 338 -521 338 -521 0 1
rlabel polysilicon 338 -527 338 -527 0 3
rlabel polysilicon 345 -521 345 -521 0 1
rlabel polysilicon 348 -527 348 -527 0 4
rlabel polysilicon 355 -521 355 -521 0 2
rlabel polysilicon 352 -527 352 -527 0 3
rlabel polysilicon 359 -521 359 -521 0 1
rlabel polysilicon 359 -527 359 -527 0 3
rlabel polysilicon 366 -521 366 -521 0 1
rlabel polysilicon 369 -521 369 -521 0 2
rlabel polysilicon 373 -527 373 -527 0 3
rlabel polysilicon 376 -527 376 -527 0 4
rlabel polysilicon 380 -521 380 -521 0 1
rlabel polysilicon 380 -527 380 -527 0 3
rlabel polysilicon 390 -521 390 -521 0 2
rlabel polysilicon 394 -521 394 -521 0 1
rlabel polysilicon 394 -527 394 -527 0 3
rlabel polysilicon 401 -521 401 -521 0 1
rlabel polysilicon 401 -527 401 -527 0 3
rlabel polysilicon 408 -521 408 -521 0 1
rlabel polysilicon 408 -527 408 -527 0 3
rlabel polysilicon 415 -521 415 -521 0 1
rlabel polysilicon 415 -527 415 -527 0 3
rlabel polysilicon 425 -521 425 -521 0 2
rlabel polysilicon 429 -521 429 -521 0 1
rlabel polysilicon 429 -527 429 -527 0 3
rlabel polysilicon 436 -521 436 -521 0 1
rlabel polysilicon 436 -527 436 -527 0 3
rlabel polysilicon 443 -521 443 -521 0 1
rlabel polysilicon 443 -527 443 -527 0 3
rlabel polysilicon 450 -521 450 -521 0 1
rlabel polysilicon 450 -527 450 -527 0 3
rlabel polysilicon 457 -521 457 -521 0 1
rlabel polysilicon 457 -527 457 -527 0 3
rlabel polysilicon 464 -521 464 -521 0 1
rlabel polysilicon 464 -527 464 -527 0 3
rlabel polysilicon 471 -521 471 -521 0 1
rlabel polysilicon 471 -527 471 -527 0 3
rlabel polysilicon 478 -521 478 -521 0 1
rlabel polysilicon 478 -527 478 -527 0 3
rlabel polysilicon 485 -521 485 -521 0 1
rlabel polysilicon 485 -527 485 -527 0 3
rlabel polysilicon 492 -521 492 -521 0 1
rlabel polysilicon 492 -527 492 -527 0 3
rlabel polysilicon 499 -521 499 -521 0 1
rlabel polysilicon 499 -527 499 -527 0 3
rlabel polysilicon 509 -521 509 -521 0 2
rlabel polysilicon 506 -527 506 -527 0 3
rlabel polysilicon 509 -527 509 -527 0 4
rlabel polysilicon 513 -521 513 -521 0 1
rlabel polysilicon 513 -527 513 -527 0 3
rlabel polysilicon 520 -521 520 -521 0 1
rlabel polysilicon 520 -527 520 -527 0 3
rlabel polysilicon 541 -521 541 -521 0 1
rlabel polysilicon 541 -527 541 -527 0 3
rlabel polysilicon 562 -521 562 -521 0 1
rlabel polysilicon 562 -527 562 -527 0 3
rlabel polysilicon 9 -570 9 -570 0 1
rlabel polysilicon 9 -576 9 -576 0 3
rlabel polysilicon 16 -570 16 -570 0 1
rlabel polysilicon 23 -576 23 -576 0 3
rlabel polysilicon 30 -570 30 -570 0 1
rlabel polysilicon 30 -576 30 -576 0 3
rlabel polysilicon 40 -570 40 -570 0 2
rlabel polysilicon 44 -576 44 -576 0 3
rlabel polysilicon 51 -570 51 -570 0 1
rlabel polysilicon 51 -576 51 -576 0 3
rlabel polysilicon 58 -570 58 -570 0 1
rlabel polysilicon 58 -576 58 -576 0 3
rlabel polysilicon 68 -570 68 -570 0 2
rlabel polysilicon 65 -576 65 -576 0 3
rlabel polysilicon 72 -570 72 -570 0 1
rlabel polysilicon 72 -576 72 -576 0 3
rlabel polysilicon 79 -570 79 -570 0 1
rlabel polysilicon 79 -576 79 -576 0 3
rlabel polysilicon 86 -576 86 -576 0 3
rlabel polysilicon 89 -576 89 -576 0 4
rlabel polysilicon 93 -570 93 -570 0 1
rlabel polysilicon 93 -576 93 -576 0 3
rlabel polysilicon 103 -570 103 -570 0 2
rlabel polysilicon 100 -576 100 -576 0 3
rlabel polysilicon 107 -570 107 -570 0 1
rlabel polysilicon 110 -576 110 -576 0 4
rlabel polysilicon 117 -570 117 -570 0 2
rlabel polysilicon 114 -576 114 -576 0 3
rlabel polysilicon 117 -576 117 -576 0 4
rlabel polysilicon 121 -570 121 -570 0 1
rlabel polysilicon 121 -576 121 -576 0 3
rlabel polysilicon 128 -570 128 -570 0 1
rlabel polysilicon 128 -576 128 -576 0 3
rlabel polysilicon 135 -570 135 -570 0 1
rlabel polysilicon 135 -576 135 -576 0 3
rlabel polysilicon 142 -570 142 -570 0 1
rlabel polysilicon 142 -576 142 -576 0 3
rlabel polysilicon 149 -570 149 -570 0 1
rlabel polysilicon 149 -576 149 -576 0 3
rlabel polysilicon 156 -570 156 -570 0 1
rlabel polysilicon 156 -576 156 -576 0 3
rlabel polysilicon 163 -570 163 -570 0 1
rlabel polysilicon 163 -576 163 -576 0 3
rlabel polysilicon 170 -570 170 -570 0 1
rlabel polysilicon 173 -576 173 -576 0 4
rlabel polysilicon 177 -570 177 -570 0 1
rlabel polysilicon 177 -576 177 -576 0 3
rlabel polysilicon 184 -570 184 -570 0 1
rlabel polysilicon 187 -576 187 -576 0 4
rlabel polysilicon 191 -570 191 -570 0 1
rlabel polysilicon 191 -576 191 -576 0 3
rlabel polysilicon 198 -570 198 -570 0 1
rlabel polysilicon 198 -576 198 -576 0 3
rlabel polysilicon 205 -570 205 -570 0 1
rlabel polysilicon 208 -570 208 -570 0 2
rlabel polysilicon 205 -576 205 -576 0 3
rlabel polysilicon 208 -576 208 -576 0 4
rlabel polysilicon 215 -570 215 -570 0 2
rlabel polysilicon 219 -570 219 -570 0 1
rlabel polysilicon 222 -570 222 -570 0 2
rlabel polysilicon 219 -576 219 -576 0 3
rlabel polysilicon 229 -570 229 -570 0 2
rlabel polysilicon 229 -576 229 -576 0 4
rlabel polysilicon 236 -570 236 -570 0 2
rlabel polysilicon 233 -576 233 -576 0 3
rlabel polysilicon 236 -576 236 -576 0 4
rlabel polysilicon 240 -570 240 -570 0 1
rlabel polysilicon 247 -570 247 -570 0 1
rlabel polysilicon 247 -576 247 -576 0 3
rlabel polysilicon 254 -570 254 -570 0 1
rlabel polysilicon 257 -570 257 -570 0 2
rlabel polysilicon 261 -570 261 -570 0 1
rlabel polysilicon 261 -576 261 -576 0 3
rlabel polysilicon 268 -570 268 -570 0 1
rlabel polysilicon 271 -570 271 -570 0 2
rlabel polysilicon 268 -576 268 -576 0 3
rlabel polysilicon 271 -576 271 -576 0 4
rlabel polysilicon 275 -570 275 -570 0 1
rlabel polysilicon 275 -576 275 -576 0 3
rlabel polysilicon 282 -570 282 -570 0 1
rlabel polysilicon 285 -576 285 -576 0 4
rlabel polysilicon 289 -570 289 -570 0 1
rlabel polysilicon 289 -576 289 -576 0 3
rlabel polysilicon 296 -570 296 -570 0 1
rlabel polysilicon 296 -576 296 -576 0 3
rlabel polysilicon 306 -570 306 -570 0 2
rlabel polysilicon 306 -576 306 -576 0 4
rlabel polysilicon 313 -570 313 -570 0 2
rlabel polysilicon 313 -576 313 -576 0 4
rlabel polysilicon 317 -570 317 -570 0 1
rlabel polysilicon 317 -576 317 -576 0 3
rlabel polysilicon 324 -570 324 -570 0 1
rlabel polysilicon 324 -576 324 -576 0 3
rlabel polysilicon 331 -570 331 -570 0 1
rlabel polysilicon 331 -576 331 -576 0 3
rlabel polysilicon 338 -570 338 -570 0 1
rlabel polysilicon 341 -570 341 -570 0 2
rlabel polysilicon 338 -576 338 -576 0 3
rlabel polysilicon 345 -570 345 -570 0 1
rlabel polysilicon 345 -576 345 -576 0 3
rlabel polysilicon 352 -570 352 -570 0 1
rlabel polysilicon 352 -576 352 -576 0 3
rlabel polysilicon 359 -570 359 -570 0 1
rlabel polysilicon 362 -570 362 -570 0 2
rlabel polysilicon 359 -576 359 -576 0 3
rlabel polysilicon 362 -576 362 -576 0 4
rlabel polysilicon 366 -570 366 -570 0 1
rlabel polysilicon 369 -570 369 -570 0 2
rlabel polysilicon 373 -570 373 -570 0 1
rlabel polysilicon 373 -576 373 -576 0 3
rlabel polysilicon 380 -570 380 -570 0 1
rlabel polysilicon 380 -576 380 -576 0 3
rlabel polysilicon 387 -570 387 -570 0 1
rlabel polysilicon 387 -576 387 -576 0 3
rlabel polysilicon 394 -570 394 -570 0 1
rlabel polysilicon 394 -576 394 -576 0 3
rlabel polysilicon 401 -570 401 -570 0 1
rlabel polysilicon 401 -576 401 -576 0 3
rlabel polysilicon 408 -570 408 -570 0 1
rlabel polysilicon 408 -576 408 -576 0 3
rlabel polysilicon 415 -570 415 -570 0 1
rlabel polysilicon 415 -576 415 -576 0 3
rlabel polysilicon 422 -570 422 -570 0 1
rlabel polysilicon 422 -576 422 -576 0 3
rlabel polysilicon 429 -570 429 -570 0 1
rlabel polysilicon 432 -576 432 -576 0 4
rlabel polysilicon 436 -570 436 -570 0 1
rlabel polysilicon 436 -576 436 -576 0 3
rlabel polysilicon 443 -570 443 -570 0 1
rlabel polysilicon 443 -576 443 -576 0 3
rlabel polysilicon 450 -570 450 -570 0 1
rlabel polysilicon 450 -576 450 -576 0 3
rlabel polysilicon 457 -570 457 -570 0 1
rlabel polysilicon 457 -576 457 -576 0 3
rlabel polysilicon 464 -570 464 -570 0 1
rlabel polysilicon 464 -576 464 -576 0 3
rlabel polysilicon 471 -570 471 -570 0 1
rlabel polysilicon 471 -576 471 -576 0 3
rlabel polysilicon 478 -570 478 -570 0 1
rlabel polysilicon 478 -576 478 -576 0 3
rlabel polysilicon 485 -570 485 -570 0 1
rlabel polysilicon 485 -576 485 -576 0 3
rlabel polysilicon 492 -570 492 -570 0 1
rlabel polysilicon 492 -576 492 -576 0 3
rlabel polysilicon 499 -576 499 -576 0 3
rlabel polysilicon 506 -570 506 -570 0 1
rlabel polysilicon 506 -576 506 -576 0 3
rlabel polysilicon 513 -576 513 -576 0 3
rlabel polysilicon 520 -570 520 -570 0 1
rlabel polysilicon 520 -576 520 -576 0 3
rlabel polysilicon 527 -570 527 -570 0 1
rlabel polysilicon 530 -570 530 -570 0 2
rlabel polysilicon 527 -576 527 -576 0 3
rlabel polysilicon 530 -576 530 -576 0 4
rlabel polysilicon 534 -570 534 -570 0 1
rlabel polysilicon 534 -576 534 -576 0 3
rlabel polysilicon 541 -570 541 -570 0 1
rlabel polysilicon 541 -576 541 -576 0 3
rlabel polysilicon 548 -576 548 -576 0 3
rlabel polysilicon 555 -570 555 -570 0 1
rlabel polysilicon 555 -576 555 -576 0 3
rlabel polysilicon 562 -570 562 -570 0 1
rlabel polysilicon 562 -576 562 -576 0 3
rlabel polysilicon 9 -613 9 -613 0 1
rlabel polysilicon 9 -619 9 -619 0 3
rlabel polysilicon 16 -613 16 -613 0 1
rlabel polysilicon 16 -619 16 -619 0 3
rlabel polysilicon 23 -613 23 -613 0 1
rlabel polysilicon 23 -619 23 -619 0 3
rlabel polysilicon 30 -613 30 -613 0 1
rlabel polysilicon 30 -619 30 -619 0 3
rlabel polysilicon 37 -613 37 -613 0 1
rlabel polysilicon 37 -619 37 -619 0 3
rlabel polysilicon 44 -619 44 -619 0 3
rlabel polysilicon 47 -619 47 -619 0 4
rlabel polysilicon 51 -613 51 -613 0 1
rlabel polysilicon 54 -613 54 -613 0 2
rlabel polysilicon 58 -613 58 -613 0 1
rlabel polysilicon 58 -619 58 -619 0 3
rlabel polysilicon 65 -613 65 -613 0 1
rlabel polysilicon 68 -619 68 -619 0 4
rlabel polysilicon 72 -613 72 -613 0 1
rlabel polysilicon 72 -619 72 -619 0 3
rlabel polysilicon 79 -613 79 -613 0 1
rlabel polysilicon 82 -613 82 -613 0 2
rlabel polysilicon 86 -619 86 -619 0 3
rlabel polysilicon 89 -619 89 -619 0 4
rlabel polysilicon 93 -613 93 -613 0 1
rlabel polysilicon 93 -619 93 -619 0 3
rlabel polysilicon 103 -613 103 -613 0 2
rlabel polysilicon 103 -619 103 -619 0 4
rlabel polysilicon 107 -613 107 -613 0 1
rlabel polysilicon 107 -619 107 -619 0 3
rlabel polysilicon 114 -619 114 -619 0 3
rlabel polysilicon 121 -613 121 -613 0 1
rlabel polysilicon 121 -619 121 -619 0 3
rlabel polysilicon 131 -613 131 -613 0 2
rlabel polysilicon 131 -619 131 -619 0 4
rlabel polysilicon 135 -613 135 -613 0 1
rlabel polysilicon 138 -613 138 -613 0 2
rlabel polysilicon 142 -613 142 -613 0 1
rlabel polysilicon 145 -613 145 -613 0 2
rlabel polysilicon 142 -619 142 -619 0 3
rlabel polysilicon 149 -613 149 -613 0 1
rlabel polysilicon 149 -619 149 -619 0 3
rlabel polysilicon 156 -613 156 -613 0 1
rlabel polysilicon 156 -619 156 -619 0 3
rlabel polysilicon 163 -613 163 -613 0 1
rlabel polysilicon 163 -619 163 -619 0 3
rlabel polysilicon 170 -613 170 -613 0 1
rlabel polysilicon 170 -619 170 -619 0 3
rlabel polysilicon 177 -619 177 -619 0 3
rlabel polysilicon 180 -619 180 -619 0 4
rlabel polysilicon 187 -619 187 -619 0 4
rlabel polysilicon 191 -613 191 -613 0 1
rlabel polysilicon 191 -619 191 -619 0 3
rlabel polysilicon 198 -613 198 -613 0 1
rlabel polysilicon 198 -619 198 -619 0 3
rlabel polysilicon 205 -613 205 -613 0 1
rlabel polysilicon 205 -619 205 -619 0 3
rlabel polysilicon 212 -613 212 -613 0 1
rlabel polysilicon 212 -619 212 -619 0 3
rlabel polysilicon 219 -613 219 -613 0 1
rlabel polysilicon 222 -613 222 -613 0 2
rlabel polysilicon 219 -619 219 -619 0 3
rlabel polysilicon 222 -619 222 -619 0 4
rlabel polysilicon 226 -613 226 -613 0 1
rlabel polysilicon 229 -613 229 -613 0 2
rlabel polysilicon 226 -619 226 -619 0 3
rlabel polysilicon 233 -613 233 -613 0 1
rlabel polysilicon 233 -619 233 -619 0 3
rlabel polysilicon 240 -613 240 -613 0 1
rlabel polysilicon 240 -619 240 -619 0 3
rlabel polysilicon 247 -613 247 -613 0 1
rlabel polysilicon 247 -619 247 -619 0 3
rlabel polysilicon 254 -613 254 -613 0 1
rlabel polysilicon 254 -619 254 -619 0 3
rlabel polysilicon 261 -613 261 -613 0 1
rlabel polysilicon 261 -619 261 -619 0 3
rlabel polysilicon 268 -613 268 -613 0 1
rlabel polysilicon 268 -619 268 -619 0 3
rlabel polysilicon 275 -613 275 -613 0 1
rlabel polysilicon 275 -619 275 -619 0 3
rlabel polysilicon 282 -613 282 -613 0 1
rlabel polysilicon 282 -619 282 -619 0 3
rlabel polysilicon 289 -613 289 -613 0 1
rlabel polysilicon 289 -619 289 -619 0 3
rlabel polysilicon 292 -619 292 -619 0 4
rlabel polysilicon 299 -613 299 -613 0 2
rlabel polysilicon 296 -619 296 -619 0 3
rlabel polysilicon 299 -619 299 -619 0 4
rlabel polysilicon 303 -613 303 -613 0 1
rlabel polysilicon 303 -619 303 -619 0 3
rlabel polysilicon 310 -613 310 -613 0 1
rlabel polysilicon 310 -619 310 -619 0 3
rlabel polysilicon 317 -613 317 -613 0 1
rlabel polysilicon 317 -619 317 -619 0 3
rlabel polysilicon 327 -613 327 -613 0 2
rlabel polysilicon 324 -619 324 -619 0 3
rlabel polysilicon 327 -619 327 -619 0 4
rlabel polysilicon 331 -613 331 -613 0 1
rlabel polysilicon 331 -619 331 -619 0 3
rlabel polysilicon 338 -613 338 -613 0 1
rlabel polysilicon 341 -613 341 -613 0 2
rlabel polysilicon 341 -619 341 -619 0 4
rlabel polysilicon 345 -613 345 -613 0 1
rlabel polysilicon 345 -619 345 -619 0 3
rlabel polysilicon 352 -613 352 -613 0 1
rlabel polysilicon 352 -619 352 -619 0 3
rlabel polysilicon 355 -619 355 -619 0 4
rlabel polysilicon 359 -613 359 -613 0 1
rlabel polysilicon 359 -619 359 -619 0 3
rlabel polysilicon 366 -613 366 -613 0 1
rlabel polysilicon 366 -619 366 -619 0 3
rlabel polysilicon 373 -613 373 -613 0 1
rlabel polysilicon 373 -619 373 -619 0 3
rlabel polysilicon 380 -613 380 -613 0 1
rlabel polysilicon 380 -619 380 -619 0 3
rlabel polysilicon 387 -613 387 -613 0 1
rlabel polysilicon 387 -619 387 -619 0 3
rlabel polysilicon 394 -613 394 -613 0 1
rlabel polysilicon 394 -619 394 -619 0 3
rlabel polysilicon 397 -619 397 -619 0 4
rlabel polysilicon 401 -613 401 -613 0 1
rlabel polysilicon 401 -619 401 -619 0 3
rlabel polysilicon 408 -613 408 -613 0 1
rlabel polysilicon 408 -619 408 -619 0 3
rlabel polysilicon 418 -619 418 -619 0 4
rlabel polysilicon 422 -613 422 -613 0 1
rlabel polysilicon 422 -619 422 -619 0 3
rlabel polysilicon 429 -613 429 -613 0 1
rlabel polysilicon 429 -619 429 -619 0 3
rlabel polysilicon 436 -613 436 -613 0 1
rlabel polysilicon 436 -619 436 -619 0 3
rlabel polysilicon 443 -613 443 -613 0 1
rlabel polysilicon 443 -619 443 -619 0 3
rlabel polysilicon 450 -613 450 -613 0 1
rlabel polysilicon 450 -619 450 -619 0 3
rlabel polysilicon 457 -613 457 -613 0 1
rlabel polysilicon 457 -619 457 -619 0 3
rlabel polysilicon 464 -613 464 -613 0 1
rlabel polysilicon 464 -619 464 -619 0 3
rlabel polysilicon 471 -613 471 -613 0 1
rlabel polysilicon 471 -619 471 -619 0 3
rlabel polysilicon 481 -613 481 -613 0 2
rlabel polysilicon 481 -619 481 -619 0 4
rlabel polysilicon 485 -613 485 -613 0 1
rlabel polysilicon 485 -619 485 -619 0 3
rlabel polysilicon 492 -613 492 -613 0 1
rlabel polysilicon 492 -619 492 -619 0 3
rlabel polysilicon 499 -613 499 -613 0 1
rlabel polysilicon 499 -619 499 -619 0 3
rlabel polysilicon 509 -613 509 -613 0 2
rlabel polysilicon 513 -613 513 -613 0 1
rlabel polysilicon 516 -613 516 -613 0 2
rlabel polysilicon 516 -619 516 -619 0 4
rlabel polysilicon 520 -613 520 -613 0 1
rlabel polysilicon 523 -613 523 -613 0 2
rlabel polysilicon 527 -613 527 -613 0 1
rlabel polysilicon 527 -619 527 -619 0 3
rlabel polysilicon 534 -613 534 -613 0 1
rlabel polysilicon 534 -619 534 -619 0 3
rlabel polysilicon 541 -613 541 -613 0 1
rlabel polysilicon 541 -619 541 -619 0 3
rlabel polysilicon 548 -613 548 -613 0 1
rlabel polysilicon 548 -619 548 -619 0 3
rlabel polysilicon 555 -613 555 -613 0 1
rlabel polysilicon 555 -619 555 -619 0 3
rlabel polysilicon 562 -613 562 -613 0 1
rlabel polysilicon 40 -660 40 -660 0 2
rlabel polysilicon 44 -660 44 -660 0 1
rlabel polysilicon 44 -666 44 -666 0 3
rlabel polysilicon 51 -660 51 -660 0 1
rlabel polysilicon 51 -666 51 -666 0 3
rlabel polysilicon 61 -660 61 -660 0 2
rlabel polysilicon 58 -666 58 -666 0 3
rlabel polysilicon 65 -660 65 -660 0 1
rlabel polysilicon 65 -666 65 -666 0 3
rlabel polysilicon 72 -660 72 -660 0 1
rlabel polysilicon 75 -660 75 -660 0 2
rlabel polysilicon 79 -660 79 -660 0 1
rlabel polysilicon 79 -666 79 -666 0 3
rlabel polysilicon 86 -660 86 -660 0 1
rlabel polysilicon 86 -666 86 -666 0 3
rlabel polysilicon 96 -660 96 -660 0 2
rlabel polysilicon 100 -660 100 -660 0 1
rlabel polysilicon 100 -666 100 -666 0 3
rlabel polysilicon 103 -666 103 -666 0 4
rlabel polysilicon 107 -660 107 -660 0 1
rlabel polysilicon 107 -666 107 -666 0 3
rlabel polysilicon 114 -660 114 -660 0 1
rlabel polysilicon 117 -660 117 -660 0 2
rlabel polysilicon 114 -666 114 -666 0 3
rlabel polysilicon 121 -660 121 -660 0 1
rlabel polysilicon 121 -666 121 -666 0 3
rlabel polysilicon 128 -660 128 -660 0 1
rlabel polysilicon 131 -660 131 -660 0 2
rlabel polysilicon 135 -660 135 -660 0 1
rlabel polysilicon 135 -666 135 -666 0 3
rlabel polysilicon 142 -666 142 -666 0 3
rlabel polysilicon 149 -660 149 -660 0 1
rlabel polysilicon 149 -666 149 -666 0 3
rlabel polysilicon 156 -660 156 -660 0 1
rlabel polysilicon 156 -666 156 -666 0 3
rlabel polysilicon 163 -660 163 -660 0 1
rlabel polysilicon 163 -666 163 -666 0 3
rlabel polysilicon 170 -660 170 -660 0 1
rlabel polysilicon 170 -666 170 -666 0 3
rlabel polysilicon 177 -660 177 -660 0 1
rlabel polysilicon 177 -666 177 -666 0 3
rlabel polysilicon 184 -660 184 -660 0 1
rlabel polysilicon 184 -666 184 -666 0 3
rlabel polysilicon 191 -660 191 -660 0 1
rlabel polysilicon 191 -666 191 -666 0 3
rlabel polysilicon 201 -666 201 -666 0 4
rlabel polysilicon 208 -660 208 -660 0 2
rlabel polysilicon 205 -666 205 -666 0 3
rlabel polysilicon 212 -660 212 -660 0 1
rlabel polysilicon 212 -666 212 -666 0 3
rlabel polysilicon 219 -660 219 -660 0 1
rlabel polysilicon 219 -666 219 -666 0 3
rlabel polysilicon 226 -660 226 -660 0 1
rlabel polysilicon 226 -666 226 -666 0 3
rlabel polysilicon 233 -660 233 -660 0 1
rlabel polysilicon 233 -666 233 -666 0 3
rlabel polysilicon 243 -666 243 -666 0 4
rlabel polysilicon 247 -660 247 -660 0 1
rlabel polysilicon 250 -660 250 -660 0 2
rlabel polysilicon 247 -666 247 -666 0 3
rlabel polysilicon 250 -666 250 -666 0 4
rlabel polysilicon 254 -660 254 -660 0 1
rlabel polysilicon 254 -666 254 -666 0 3
rlabel polysilicon 261 -660 261 -660 0 1
rlabel polysilicon 261 -666 261 -666 0 3
rlabel polysilicon 268 -666 268 -666 0 3
rlabel polysilicon 271 -666 271 -666 0 4
rlabel polysilicon 275 -660 275 -660 0 1
rlabel polysilicon 275 -666 275 -666 0 3
rlabel polysilicon 282 -660 282 -660 0 1
rlabel polysilicon 282 -666 282 -666 0 3
rlabel polysilicon 289 -660 289 -660 0 1
rlabel polysilicon 289 -666 289 -666 0 3
rlabel polysilicon 296 -660 296 -660 0 1
rlabel polysilicon 296 -666 296 -666 0 3
rlabel polysilicon 303 -660 303 -660 0 1
rlabel polysilicon 303 -666 303 -666 0 3
rlabel polysilicon 310 -660 310 -660 0 1
rlabel polysilicon 310 -666 310 -666 0 3
rlabel polysilicon 320 -660 320 -660 0 2
rlabel polysilicon 320 -666 320 -666 0 4
rlabel polysilicon 324 -660 324 -660 0 1
rlabel polysilicon 324 -666 324 -666 0 3
rlabel polysilicon 331 -660 331 -660 0 1
rlabel polysilicon 334 -660 334 -660 0 2
rlabel polysilicon 338 -660 338 -660 0 1
rlabel polysilicon 341 -660 341 -660 0 2
rlabel polysilicon 338 -666 338 -666 0 3
rlabel polysilicon 345 -660 345 -660 0 1
rlabel polysilicon 348 -660 348 -660 0 2
rlabel polysilicon 345 -666 345 -666 0 3
rlabel polysilicon 348 -666 348 -666 0 4
rlabel polysilicon 352 -660 352 -660 0 1
rlabel polysilicon 359 -660 359 -660 0 1
rlabel polysilicon 359 -666 359 -666 0 3
rlabel polysilicon 366 -660 366 -660 0 1
rlabel polysilicon 366 -666 366 -666 0 3
rlabel polysilicon 373 -666 373 -666 0 3
rlabel polysilicon 376 -666 376 -666 0 4
rlabel polysilicon 380 -660 380 -660 0 1
rlabel polysilicon 380 -666 380 -666 0 3
rlabel polysilicon 387 -660 387 -660 0 1
rlabel polysilicon 387 -666 387 -666 0 3
rlabel polysilicon 397 -660 397 -660 0 2
rlabel polysilicon 394 -666 394 -666 0 3
rlabel polysilicon 397 -666 397 -666 0 4
rlabel polysilicon 401 -660 401 -660 0 1
rlabel polysilicon 401 -666 401 -666 0 3
rlabel polysilicon 404 -666 404 -666 0 4
rlabel polysilicon 408 -660 408 -660 0 1
rlabel polysilicon 408 -666 408 -666 0 3
rlabel polysilicon 415 -660 415 -660 0 1
rlabel polysilicon 415 -666 415 -666 0 3
rlabel polysilicon 422 -660 422 -660 0 1
rlabel polysilicon 422 -666 422 -666 0 3
rlabel polysilicon 429 -660 429 -660 0 1
rlabel polysilicon 429 -666 429 -666 0 3
rlabel polysilicon 436 -660 436 -660 0 1
rlabel polysilicon 436 -666 436 -666 0 3
rlabel polysilicon 443 -660 443 -660 0 1
rlabel polysilicon 443 -666 443 -666 0 3
rlabel polysilicon 450 -660 450 -660 0 1
rlabel polysilicon 450 -666 450 -666 0 3
rlabel polysilicon 457 -660 457 -660 0 1
rlabel polysilicon 457 -666 457 -666 0 3
rlabel polysilicon 464 -660 464 -660 0 1
rlabel polysilicon 464 -666 464 -666 0 3
rlabel polysilicon 471 -660 471 -660 0 1
rlabel polysilicon 474 -660 474 -660 0 2
rlabel polysilicon 471 -666 471 -666 0 3
rlabel polysilicon 474 -666 474 -666 0 4
rlabel polysilicon 478 -660 478 -660 0 1
rlabel polysilicon 478 -666 478 -666 0 3
rlabel polysilicon 488 -660 488 -660 0 2
rlabel polysilicon 488 -666 488 -666 0 4
rlabel polysilicon 492 -660 492 -660 0 1
rlabel polysilicon 492 -666 492 -666 0 3
rlabel polysilicon 499 -660 499 -660 0 1
rlabel polysilicon 499 -666 499 -666 0 3
rlabel polysilicon 506 -660 506 -660 0 1
rlabel polysilicon 506 -666 506 -666 0 3
rlabel polysilicon 513 -660 513 -660 0 1
rlabel polysilicon 516 -660 516 -660 0 2
rlabel polysilicon 516 -666 516 -666 0 4
rlabel polysilicon 520 -660 520 -660 0 1
rlabel polysilicon 520 -666 520 -666 0 3
rlabel polysilicon 530 -660 530 -660 0 2
rlabel polysilicon 530 -666 530 -666 0 4
rlabel polysilicon 534 -660 534 -660 0 1
rlabel polysilicon 534 -666 534 -666 0 3
rlabel polysilicon 544 -660 544 -660 0 2
rlabel polysilicon 544 -666 544 -666 0 4
rlabel polysilicon 548 -660 548 -660 0 1
rlabel polysilicon 548 -666 548 -666 0 3
rlabel polysilicon 555 -660 555 -660 0 1
rlabel polysilicon 555 -666 555 -666 0 3
rlabel polysilicon 562 -660 562 -660 0 1
rlabel polysilicon 583 -660 583 -660 0 1
rlabel polysilicon 583 -666 583 -666 0 3
rlabel polysilicon 16 -709 16 -709 0 1
rlabel polysilicon 16 -715 16 -715 0 3
rlabel polysilicon 23 -709 23 -709 0 1
rlabel polysilicon 23 -715 23 -715 0 3
rlabel polysilicon 30 -709 30 -709 0 1
rlabel polysilicon 37 -709 37 -709 0 1
rlabel polysilicon 37 -715 37 -715 0 3
rlabel polysilicon 44 -709 44 -709 0 1
rlabel polysilicon 44 -715 44 -715 0 3
rlabel polysilicon 51 -709 51 -709 0 1
rlabel polysilicon 51 -715 51 -715 0 3
rlabel polysilicon 58 -715 58 -715 0 3
rlabel polysilicon 65 -709 65 -709 0 1
rlabel polysilicon 65 -715 65 -715 0 3
rlabel polysilicon 72 -709 72 -709 0 1
rlabel polysilicon 72 -715 72 -715 0 3
rlabel polysilicon 75 -715 75 -715 0 4
rlabel polysilicon 79 -709 79 -709 0 1
rlabel polysilicon 79 -715 79 -715 0 3
rlabel polysilicon 86 -709 86 -709 0 1
rlabel polysilicon 86 -715 86 -715 0 3
rlabel polysilicon 93 -709 93 -709 0 1
rlabel polysilicon 93 -715 93 -715 0 3
rlabel polysilicon 103 -709 103 -709 0 2
rlabel polysilicon 103 -715 103 -715 0 4
rlabel polysilicon 110 -709 110 -709 0 2
rlabel polysilicon 107 -715 107 -715 0 3
rlabel polysilicon 114 -709 114 -709 0 1
rlabel polysilicon 114 -715 114 -715 0 3
rlabel polysilicon 121 -709 121 -709 0 1
rlabel polysilicon 121 -715 121 -715 0 3
rlabel polysilicon 128 -709 128 -709 0 1
rlabel polysilicon 128 -715 128 -715 0 3
rlabel polysilicon 135 -709 135 -709 0 1
rlabel polysilicon 142 -709 142 -709 0 1
rlabel polysilicon 142 -715 142 -715 0 3
rlabel polysilicon 149 -709 149 -709 0 1
rlabel polysilicon 149 -715 149 -715 0 3
rlabel polysilicon 152 -715 152 -715 0 4
rlabel polysilicon 156 -709 156 -709 0 1
rlabel polysilicon 156 -715 156 -715 0 3
rlabel polysilicon 163 -709 163 -709 0 1
rlabel polysilicon 166 -709 166 -709 0 2
rlabel polysilicon 163 -715 163 -715 0 3
rlabel polysilicon 170 -709 170 -709 0 1
rlabel polysilicon 170 -715 170 -715 0 3
rlabel polysilicon 177 -709 177 -709 0 1
rlabel polysilicon 177 -715 177 -715 0 3
rlabel polysilicon 184 -709 184 -709 0 1
rlabel polysilicon 184 -715 184 -715 0 3
rlabel polysilicon 187 -715 187 -715 0 4
rlabel polysilicon 194 -709 194 -709 0 2
rlabel polysilicon 191 -715 191 -715 0 3
rlabel polysilicon 194 -715 194 -715 0 4
rlabel polysilicon 198 -709 198 -709 0 1
rlabel polysilicon 201 -709 201 -709 0 2
rlabel polysilicon 198 -715 198 -715 0 3
rlabel polysilicon 201 -715 201 -715 0 4
rlabel polysilicon 205 -709 205 -709 0 1
rlabel polysilicon 205 -715 205 -715 0 3
rlabel polysilicon 212 -709 212 -709 0 1
rlabel polysilicon 212 -715 212 -715 0 3
rlabel polysilicon 219 -709 219 -709 0 1
rlabel polysilicon 219 -715 219 -715 0 3
rlabel polysilicon 222 -715 222 -715 0 4
rlabel polysilicon 226 -709 226 -709 0 1
rlabel polysilicon 226 -715 226 -715 0 3
rlabel polysilicon 233 -709 233 -709 0 1
rlabel polysilicon 233 -715 233 -715 0 3
rlabel polysilicon 240 -709 240 -709 0 1
rlabel polysilicon 240 -715 240 -715 0 3
rlabel polysilicon 247 -709 247 -709 0 1
rlabel polysilicon 247 -715 247 -715 0 3
rlabel polysilicon 254 -709 254 -709 0 1
rlabel polysilicon 254 -715 254 -715 0 3
rlabel polysilicon 261 -709 261 -709 0 1
rlabel polysilicon 261 -715 261 -715 0 3
rlabel polysilicon 268 -709 268 -709 0 1
rlabel polysilicon 268 -715 268 -715 0 3
rlabel polysilicon 275 -709 275 -709 0 1
rlabel polysilicon 275 -715 275 -715 0 3
rlabel polysilicon 282 -715 282 -715 0 3
rlabel polysilicon 289 -709 289 -709 0 1
rlabel polysilicon 289 -715 289 -715 0 3
rlabel polysilicon 296 -709 296 -709 0 1
rlabel polysilicon 299 -709 299 -709 0 2
rlabel polysilicon 296 -715 296 -715 0 3
rlabel polysilicon 303 -709 303 -709 0 1
rlabel polysilicon 303 -715 303 -715 0 3
rlabel polysilicon 310 -709 310 -709 0 1
rlabel polysilicon 310 -715 310 -715 0 3
rlabel polysilicon 317 -709 317 -709 0 1
rlabel polysilicon 317 -715 317 -715 0 3
rlabel polysilicon 324 -709 324 -709 0 1
rlabel polysilicon 324 -715 324 -715 0 3
rlabel polysilicon 331 -709 331 -709 0 1
rlabel polysilicon 334 -709 334 -709 0 2
rlabel polysilicon 331 -715 331 -715 0 3
rlabel polysilicon 334 -715 334 -715 0 4
rlabel polysilicon 338 -709 338 -709 0 1
rlabel polysilicon 338 -715 338 -715 0 3
rlabel polysilicon 345 -709 345 -709 0 1
rlabel polysilicon 345 -715 345 -715 0 3
rlabel polysilicon 348 -715 348 -715 0 4
rlabel polysilicon 352 -709 352 -709 0 1
rlabel polysilicon 352 -715 352 -715 0 3
rlabel polysilicon 359 -709 359 -709 0 1
rlabel polysilicon 359 -715 359 -715 0 3
rlabel polysilicon 366 -709 366 -709 0 1
rlabel polysilicon 366 -715 366 -715 0 3
rlabel polysilicon 373 -709 373 -709 0 1
rlabel polysilicon 373 -715 373 -715 0 3
rlabel polysilicon 380 -709 380 -709 0 1
rlabel polysilicon 380 -715 380 -715 0 3
rlabel polysilicon 383 -715 383 -715 0 4
rlabel polysilicon 387 -709 387 -709 0 1
rlabel polysilicon 387 -715 387 -715 0 3
rlabel polysilicon 394 -715 394 -715 0 3
rlabel polysilicon 397 -715 397 -715 0 4
rlabel polysilicon 401 -709 401 -709 0 1
rlabel polysilicon 401 -715 401 -715 0 3
rlabel polysilicon 408 -709 408 -709 0 1
rlabel polysilicon 408 -715 408 -715 0 3
rlabel polysilicon 415 -709 415 -709 0 1
rlabel polysilicon 415 -715 415 -715 0 3
rlabel polysilicon 422 -709 422 -709 0 1
rlabel polysilicon 425 -715 425 -715 0 4
rlabel polysilicon 429 -709 429 -709 0 1
rlabel polysilicon 429 -715 429 -715 0 3
rlabel polysilicon 436 -709 436 -709 0 1
rlabel polysilicon 436 -715 436 -715 0 3
rlabel polysilicon 443 -709 443 -709 0 1
rlabel polysilicon 443 -715 443 -715 0 3
rlabel polysilicon 450 -709 450 -709 0 1
rlabel polysilicon 450 -715 450 -715 0 3
rlabel polysilicon 457 -709 457 -709 0 1
rlabel polysilicon 457 -715 457 -715 0 3
rlabel polysilicon 464 -709 464 -709 0 1
rlabel polysilicon 464 -715 464 -715 0 3
rlabel polysilicon 471 -709 471 -709 0 1
rlabel polysilicon 471 -715 471 -715 0 3
rlabel polysilicon 478 -709 478 -709 0 1
rlabel polysilicon 478 -715 478 -715 0 3
rlabel polysilicon 485 -709 485 -709 0 1
rlabel polysilicon 485 -715 485 -715 0 3
rlabel polysilicon 495 -715 495 -715 0 4
rlabel polysilicon 499 -709 499 -709 0 1
rlabel polysilicon 499 -715 499 -715 0 3
rlabel polysilicon 506 -709 506 -709 0 1
rlabel polysilicon 506 -715 506 -715 0 3
rlabel polysilicon 513 -709 513 -709 0 1
rlabel polysilicon 513 -715 513 -715 0 3
rlabel polysilicon 520 -709 520 -709 0 1
rlabel polysilicon 520 -715 520 -715 0 3
rlabel polysilicon 527 -709 527 -709 0 1
rlabel polysilicon 527 -715 527 -715 0 3
rlabel polysilicon 534 -709 534 -709 0 1
rlabel polysilicon 534 -715 534 -715 0 3
rlabel polysilicon 541 -709 541 -709 0 1
rlabel polysilicon 541 -715 541 -715 0 3
rlabel polysilicon 548 -709 548 -709 0 1
rlabel polysilicon 548 -715 548 -715 0 3
rlabel polysilicon 555 -709 555 -709 0 1
rlabel polysilicon 555 -715 555 -715 0 3
rlabel polysilicon 562 -709 562 -709 0 1
rlabel polysilicon 562 -715 562 -715 0 3
rlabel polysilicon 572 -709 572 -709 0 2
rlabel polysilicon 569 -715 569 -715 0 3
rlabel polysilicon 572 -715 572 -715 0 4
rlabel polysilicon 576 -709 576 -709 0 1
rlabel polysilicon 576 -715 576 -715 0 3
rlabel polysilicon 583 -709 583 -709 0 1
rlabel polysilicon 583 -715 583 -715 0 3
rlabel polysilicon 593 -709 593 -709 0 2
rlabel polysilicon 593 -715 593 -715 0 4
rlabel polysilicon 597 -715 597 -715 0 3
rlabel polysilicon 600 -715 600 -715 0 4
rlabel polysilicon 604 -709 604 -709 0 1
rlabel polysilicon 604 -715 604 -715 0 3
rlabel polysilicon 611 -709 611 -709 0 1
rlabel polysilicon 614 -715 614 -715 0 4
rlabel polysilicon 618 -709 618 -709 0 1
rlabel polysilicon 618 -715 618 -715 0 3
rlabel polysilicon 628 -709 628 -709 0 2
rlabel polysilicon 632 -709 632 -709 0 1
rlabel polysilicon 632 -715 632 -715 0 3
rlabel polysilicon 639 -709 639 -709 0 1
rlabel polysilicon 639 -715 639 -715 0 3
rlabel polysilicon 646 -709 646 -709 0 1
rlabel polysilicon 646 -715 646 -715 0 3
rlabel polysilicon 33 -760 33 -760 0 2
rlabel polysilicon 33 -766 33 -766 0 4
rlabel polysilicon 40 -766 40 -766 0 4
rlabel polysilicon 44 -760 44 -760 0 1
rlabel polysilicon 44 -766 44 -766 0 3
rlabel polysilicon 51 -760 51 -760 0 1
rlabel polysilicon 51 -766 51 -766 0 3
rlabel polysilicon 58 -760 58 -760 0 1
rlabel polysilicon 58 -766 58 -766 0 3
rlabel polysilicon 65 -760 65 -760 0 1
rlabel polysilicon 65 -766 65 -766 0 3
rlabel polysilicon 72 -760 72 -760 0 1
rlabel polysilicon 72 -766 72 -766 0 3
rlabel polysilicon 79 -760 79 -760 0 1
rlabel polysilicon 79 -766 79 -766 0 3
rlabel polysilicon 86 -760 86 -760 0 1
rlabel polysilicon 86 -766 86 -766 0 3
rlabel polysilicon 93 -760 93 -760 0 1
rlabel polysilicon 93 -766 93 -766 0 3
rlabel polysilicon 103 -760 103 -760 0 2
rlabel polysilicon 107 -760 107 -760 0 1
rlabel polysilicon 107 -766 107 -766 0 3
rlabel polysilicon 114 -760 114 -760 0 1
rlabel polysilicon 117 -766 117 -766 0 4
rlabel polysilicon 121 -760 121 -760 0 1
rlabel polysilicon 121 -766 121 -766 0 3
rlabel polysilicon 128 -760 128 -760 0 1
rlabel polysilicon 128 -766 128 -766 0 3
rlabel polysilicon 135 -760 135 -760 0 1
rlabel polysilicon 135 -766 135 -766 0 3
rlabel polysilicon 142 -760 142 -760 0 1
rlabel polysilicon 145 -766 145 -766 0 4
rlabel polysilicon 149 -760 149 -760 0 1
rlabel polysilicon 152 -760 152 -760 0 2
rlabel polysilicon 149 -766 149 -766 0 3
rlabel polysilicon 152 -766 152 -766 0 4
rlabel polysilicon 156 -760 156 -760 0 1
rlabel polysilicon 156 -766 156 -766 0 3
rlabel polysilicon 163 -760 163 -760 0 1
rlabel polysilicon 163 -766 163 -766 0 3
rlabel polysilicon 170 -760 170 -760 0 1
rlabel polysilicon 170 -766 170 -766 0 3
rlabel polysilicon 177 -760 177 -760 0 1
rlabel polysilicon 177 -766 177 -766 0 3
rlabel polysilicon 184 -760 184 -760 0 1
rlabel polysilicon 184 -766 184 -766 0 3
rlabel polysilicon 194 -760 194 -760 0 2
rlabel polysilicon 191 -766 191 -766 0 3
rlabel polysilicon 194 -766 194 -766 0 4
rlabel polysilicon 198 -760 198 -760 0 1
rlabel polysilicon 198 -766 198 -766 0 3
rlabel polysilicon 205 -760 205 -760 0 1
rlabel polysilicon 205 -766 205 -766 0 3
rlabel polysilicon 215 -760 215 -760 0 2
rlabel polysilicon 212 -766 212 -766 0 3
rlabel polysilicon 215 -766 215 -766 0 4
rlabel polysilicon 222 -760 222 -760 0 2
rlabel polysilicon 219 -766 219 -766 0 3
rlabel polysilicon 222 -766 222 -766 0 4
rlabel polysilicon 229 -760 229 -760 0 2
rlabel polysilicon 226 -766 226 -766 0 3
rlabel polysilicon 229 -766 229 -766 0 4
rlabel polysilicon 233 -760 233 -760 0 1
rlabel polysilicon 233 -766 233 -766 0 3
rlabel polysilicon 240 -760 240 -760 0 1
rlabel polysilicon 240 -766 240 -766 0 3
rlabel polysilicon 250 -760 250 -760 0 2
rlabel polysilicon 247 -766 247 -766 0 3
rlabel polysilicon 254 -760 254 -760 0 1
rlabel polysilicon 257 -760 257 -760 0 2
rlabel polysilicon 257 -766 257 -766 0 4
rlabel polysilicon 261 -760 261 -760 0 1
rlabel polysilicon 261 -766 261 -766 0 3
rlabel polysilicon 268 -760 268 -760 0 1
rlabel polysilicon 268 -766 268 -766 0 3
rlabel polysilicon 278 -760 278 -760 0 2
rlabel polysilicon 275 -766 275 -766 0 3
rlabel polysilicon 285 -760 285 -760 0 2
rlabel polysilicon 285 -766 285 -766 0 4
rlabel polysilicon 292 -760 292 -760 0 2
rlabel polysilicon 292 -766 292 -766 0 4
rlabel polysilicon 296 -760 296 -760 0 1
rlabel polysilicon 296 -766 296 -766 0 3
rlabel polysilicon 303 -760 303 -760 0 1
rlabel polysilicon 303 -766 303 -766 0 3
rlabel polysilicon 306 -766 306 -766 0 4
rlabel polysilicon 310 -760 310 -760 0 1
rlabel polysilicon 310 -766 310 -766 0 3
rlabel polysilicon 317 -760 317 -760 0 1
rlabel polysilicon 317 -766 317 -766 0 3
rlabel polysilicon 324 -760 324 -760 0 1
rlabel polysilicon 324 -766 324 -766 0 3
rlabel polysilicon 331 -760 331 -760 0 1
rlabel polysilicon 334 -760 334 -760 0 2
rlabel polysilicon 331 -766 331 -766 0 3
rlabel polysilicon 338 -760 338 -760 0 1
rlabel polysilicon 338 -766 338 -766 0 3
rlabel polysilicon 341 -766 341 -766 0 4
rlabel polysilicon 348 -760 348 -760 0 2
rlabel polysilicon 352 -760 352 -760 0 1
rlabel polysilicon 352 -766 352 -766 0 3
rlabel polysilicon 359 -760 359 -760 0 1
rlabel polysilicon 362 -760 362 -760 0 2
rlabel polysilicon 359 -766 359 -766 0 3
rlabel polysilicon 366 -760 366 -760 0 1
rlabel polysilicon 366 -766 366 -766 0 3
rlabel polysilicon 373 -766 373 -766 0 3
rlabel polysilicon 376 -766 376 -766 0 4
rlabel polysilicon 380 -760 380 -760 0 1
rlabel polysilicon 380 -766 380 -766 0 3
rlabel polysilicon 387 -760 387 -760 0 1
rlabel polysilicon 387 -766 387 -766 0 3
rlabel polysilicon 394 -760 394 -760 0 1
rlabel polysilicon 397 -766 397 -766 0 4
rlabel polysilicon 401 -760 401 -760 0 1
rlabel polysilicon 401 -766 401 -766 0 3
rlabel polysilicon 408 -760 408 -760 0 1
rlabel polysilicon 408 -766 408 -766 0 3
rlabel polysilicon 415 -760 415 -760 0 1
rlabel polysilicon 415 -766 415 -766 0 3
rlabel polysilicon 422 -760 422 -760 0 1
rlabel polysilicon 422 -766 422 -766 0 3
rlabel polysilicon 429 -760 429 -760 0 1
rlabel polysilicon 429 -766 429 -766 0 3
rlabel polysilicon 436 -760 436 -760 0 1
rlabel polysilicon 436 -766 436 -766 0 3
rlabel polysilicon 443 -766 443 -766 0 3
rlabel polysilicon 446 -766 446 -766 0 4
rlabel polysilicon 450 -760 450 -760 0 1
rlabel polysilicon 450 -766 450 -766 0 3
rlabel polysilicon 457 -760 457 -760 0 1
rlabel polysilicon 457 -766 457 -766 0 3
rlabel polysilicon 464 -760 464 -760 0 1
rlabel polysilicon 464 -766 464 -766 0 3
rlabel polysilicon 471 -760 471 -760 0 1
rlabel polysilicon 474 -760 474 -760 0 2
rlabel polysilicon 471 -766 471 -766 0 3
rlabel polysilicon 478 -760 478 -760 0 1
rlabel polysilicon 478 -766 478 -766 0 3
rlabel polysilicon 485 -760 485 -760 0 1
rlabel polysilicon 488 -760 488 -760 0 2
rlabel polysilicon 492 -760 492 -760 0 1
rlabel polysilicon 492 -766 492 -766 0 3
rlabel polysilicon 499 -760 499 -760 0 1
rlabel polysilicon 499 -766 499 -766 0 3
rlabel polysilicon 506 -760 506 -760 0 1
rlabel polysilicon 506 -766 506 -766 0 3
rlabel polysilicon 513 -760 513 -760 0 1
rlabel polysilicon 513 -766 513 -766 0 3
rlabel polysilicon 520 -760 520 -760 0 1
rlabel polysilicon 520 -766 520 -766 0 3
rlabel polysilicon 527 -760 527 -760 0 1
rlabel polysilicon 530 -760 530 -760 0 2
rlabel polysilicon 530 -766 530 -766 0 4
rlabel polysilicon 534 -760 534 -760 0 1
rlabel polysilicon 534 -766 534 -766 0 3
rlabel polysilicon 541 -760 541 -760 0 1
rlabel polysilicon 541 -766 541 -766 0 3
rlabel polysilicon 555 -760 555 -760 0 1
rlabel polysilicon 555 -766 555 -766 0 3
rlabel polysilicon 611 -760 611 -760 0 1
rlabel polysilicon 26 -817 26 -817 0 2
rlabel polysilicon 30 -817 30 -817 0 1
rlabel polysilicon 37 -817 37 -817 0 1
rlabel polysilicon 37 -823 37 -823 0 3
rlabel polysilicon 44 -817 44 -817 0 1
rlabel polysilicon 44 -823 44 -823 0 3
rlabel polysilicon 51 -817 51 -817 0 1
rlabel polysilicon 51 -823 51 -823 0 3
rlabel polysilicon 58 -817 58 -817 0 1
rlabel polysilicon 65 -817 65 -817 0 1
rlabel polysilicon 65 -823 65 -823 0 3
rlabel polysilicon 72 -817 72 -817 0 1
rlabel polysilicon 79 -817 79 -817 0 1
rlabel polysilicon 79 -823 79 -823 0 3
rlabel polysilicon 86 -817 86 -817 0 1
rlabel polysilicon 86 -823 86 -823 0 3
rlabel polysilicon 93 -817 93 -817 0 1
rlabel polysilicon 93 -823 93 -823 0 3
rlabel polysilicon 103 -817 103 -817 0 2
rlabel polysilicon 107 -817 107 -817 0 1
rlabel polysilicon 110 -823 110 -823 0 4
rlabel polysilicon 114 -817 114 -817 0 1
rlabel polysilicon 121 -817 121 -817 0 1
rlabel polysilicon 124 -823 124 -823 0 4
rlabel polysilicon 128 -817 128 -817 0 1
rlabel polysilicon 128 -823 128 -823 0 3
rlabel polysilicon 135 -817 135 -817 0 1
rlabel polysilicon 135 -823 135 -823 0 3
rlabel polysilicon 142 -817 142 -817 0 1
rlabel polysilicon 145 -817 145 -817 0 2
rlabel polysilicon 145 -823 145 -823 0 4
rlabel polysilicon 152 -817 152 -817 0 2
rlabel polysilicon 149 -823 149 -823 0 3
rlabel polysilicon 152 -823 152 -823 0 4
rlabel polysilicon 156 -817 156 -817 0 1
rlabel polysilicon 159 -823 159 -823 0 4
rlabel polysilicon 163 -817 163 -817 0 1
rlabel polysilicon 166 -817 166 -817 0 2
rlabel polysilicon 163 -823 163 -823 0 3
rlabel polysilicon 170 -817 170 -817 0 1
rlabel polysilicon 170 -823 170 -823 0 3
rlabel polysilicon 177 -817 177 -817 0 1
rlabel polysilicon 177 -823 177 -823 0 3
rlabel polysilicon 187 -817 187 -817 0 2
rlabel polysilicon 187 -823 187 -823 0 4
rlabel polysilicon 191 -817 191 -817 0 1
rlabel polysilicon 191 -823 191 -823 0 3
rlabel polysilicon 198 -823 198 -823 0 3
rlabel polysilicon 201 -823 201 -823 0 4
rlabel polysilicon 205 -817 205 -817 0 1
rlabel polysilicon 205 -823 205 -823 0 3
rlabel polysilicon 212 -817 212 -817 0 1
rlabel polysilicon 215 -817 215 -817 0 2
rlabel polysilicon 219 -817 219 -817 0 1
rlabel polysilicon 219 -823 219 -823 0 3
rlabel polysilicon 226 -817 226 -817 0 1
rlabel polysilicon 226 -823 226 -823 0 3
rlabel polysilicon 236 -817 236 -817 0 2
rlabel polysilicon 233 -823 233 -823 0 3
rlabel polysilicon 236 -823 236 -823 0 4
rlabel polysilicon 240 -817 240 -817 0 1
rlabel polysilicon 240 -823 240 -823 0 3
rlabel polysilicon 247 -817 247 -817 0 1
rlabel polysilicon 247 -823 247 -823 0 3
rlabel polysilicon 254 -817 254 -817 0 1
rlabel polysilicon 257 -817 257 -817 0 2
rlabel polysilicon 257 -823 257 -823 0 4
rlabel polysilicon 261 -817 261 -817 0 1
rlabel polysilicon 261 -823 261 -823 0 3
rlabel polysilicon 268 -817 268 -817 0 1
rlabel polysilicon 268 -823 268 -823 0 3
rlabel polysilicon 275 -817 275 -817 0 1
rlabel polysilicon 275 -823 275 -823 0 3
rlabel polysilicon 282 -817 282 -817 0 1
rlabel polysilicon 282 -823 282 -823 0 3
rlabel polysilicon 289 -817 289 -817 0 1
rlabel polysilicon 289 -823 289 -823 0 3
rlabel polysilicon 296 -817 296 -817 0 1
rlabel polysilicon 296 -823 296 -823 0 3
rlabel polysilicon 303 -817 303 -817 0 1
rlabel polysilicon 303 -823 303 -823 0 3
rlabel polysilicon 313 -817 313 -817 0 2
rlabel polysilicon 310 -823 310 -823 0 3
rlabel polysilicon 313 -823 313 -823 0 4
rlabel polysilicon 317 -817 317 -817 0 1
rlabel polysilicon 317 -823 317 -823 0 3
rlabel polysilicon 320 -823 320 -823 0 4
rlabel polysilicon 324 -817 324 -817 0 1
rlabel polysilicon 324 -823 324 -823 0 3
rlabel polysilicon 331 -817 331 -817 0 1
rlabel polysilicon 334 -817 334 -817 0 2
rlabel polysilicon 338 -817 338 -817 0 1
rlabel polysilicon 338 -823 338 -823 0 3
rlabel polysilicon 348 -823 348 -823 0 4
rlabel polysilicon 352 -817 352 -817 0 1
rlabel polysilicon 355 -823 355 -823 0 4
rlabel polysilicon 359 -817 359 -817 0 1
rlabel polysilicon 359 -823 359 -823 0 3
rlabel polysilicon 366 -817 366 -817 0 1
rlabel polysilicon 366 -823 366 -823 0 3
rlabel polysilicon 376 -817 376 -817 0 2
rlabel polysilicon 373 -823 373 -823 0 3
rlabel polysilicon 376 -823 376 -823 0 4
rlabel polysilicon 380 -817 380 -817 0 1
rlabel polysilicon 380 -823 380 -823 0 3
rlabel polysilicon 387 -817 387 -817 0 1
rlabel polysilicon 387 -823 387 -823 0 3
rlabel polysilicon 394 -817 394 -817 0 1
rlabel polysilicon 394 -823 394 -823 0 3
rlabel polysilicon 404 -817 404 -817 0 2
rlabel polysilicon 401 -823 401 -823 0 3
rlabel polysilicon 404 -823 404 -823 0 4
rlabel polysilicon 408 -817 408 -817 0 1
rlabel polysilicon 408 -823 408 -823 0 3
rlabel polysilicon 415 -817 415 -817 0 1
rlabel polysilicon 415 -823 415 -823 0 3
rlabel polysilicon 422 -817 422 -817 0 1
rlabel polysilicon 422 -823 422 -823 0 3
rlabel polysilicon 429 -817 429 -817 0 1
rlabel polysilicon 429 -823 429 -823 0 3
rlabel polysilicon 436 -817 436 -817 0 1
rlabel polysilicon 436 -823 436 -823 0 3
rlabel polysilicon 443 -817 443 -817 0 1
rlabel polysilicon 443 -823 443 -823 0 3
rlabel polysilicon 450 -817 450 -817 0 1
rlabel polysilicon 450 -823 450 -823 0 3
rlabel polysilicon 460 -817 460 -817 0 2
rlabel polysilicon 464 -817 464 -817 0 1
rlabel polysilicon 464 -823 464 -823 0 3
rlabel polysilicon 471 -817 471 -817 0 1
rlabel polysilicon 471 -823 471 -823 0 3
rlabel polysilicon 478 -817 478 -817 0 1
rlabel polysilicon 478 -823 478 -823 0 3
rlabel polysilicon 485 -817 485 -817 0 1
rlabel polysilicon 485 -823 485 -823 0 3
rlabel polysilicon 492 -817 492 -817 0 1
rlabel polysilicon 492 -823 492 -823 0 3
rlabel polysilicon 499 -817 499 -817 0 1
rlabel polysilicon 499 -823 499 -823 0 3
rlabel polysilicon 506 -817 506 -817 0 1
rlabel polysilicon 506 -823 506 -823 0 3
rlabel polysilicon 513 -817 513 -817 0 1
rlabel polysilicon 513 -823 513 -823 0 3
rlabel polysilicon 520 -817 520 -817 0 1
rlabel polysilicon 520 -823 520 -823 0 3
rlabel polysilicon 527 -817 527 -817 0 1
rlabel polysilicon 527 -823 527 -823 0 3
rlabel polysilicon 534 -817 534 -817 0 1
rlabel polysilicon 534 -823 534 -823 0 3
rlabel polysilicon 541 -817 541 -817 0 1
rlabel polysilicon 541 -823 541 -823 0 3
rlabel polysilicon 548 -817 548 -817 0 1
rlabel polysilicon 548 -823 548 -823 0 3
rlabel polysilicon 555 -817 555 -817 0 1
rlabel polysilicon 558 -817 558 -817 0 2
rlabel polysilicon 558 -823 558 -823 0 4
rlabel polysilicon 26 -880 26 -880 0 2
rlabel polysilicon 30 -880 30 -880 0 1
rlabel polysilicon 37 -880 37 -880 0 1
rlabel polysilicon 40 -880 40 -880 0 2
rlabel polysilicon 44 -880 44 -880 0 1
rlabel polysilicon 44 -886 44 -886 0 3
rlabel polysilicon 51 -880 51 -880 0 1
rlabel polysilicon 51 -886 51 -886 0 3
rlabel polysilicon 58 -880 58 -880 0 1
rlabel polysilicon 58 -886 58 -886 0 3
rlabel polysilicon 65 -880 65 -880 0 1
rlabel polysilicon 65 -886 65 -886 0 3
rlabel polysilicon 72 -880 72 -880 0 1
rlabel polysilicon 75 -880 75 -880 0 2
rlabel polysilicon 79 -880 79 -880 0 1
rlabel polysilicon 79 -886 79 -886 0 3
rlabel polysilicon 86 -880 86 -880 0 1
rlabel polysilicon 86 -886 86 -886 0 3
rlabel polysilicon 93 -880 93 -880 0 1
rlabel polysilicon 93 -886 93 -886 0 3
rlabel polysilicon 100 -880 100 -880 0 1
rlabel polysilicon 100 -886 100 -886 0 3
rlabel polysilicon 107 -880 107 -880 0 1
rlabel polysilicon 107 -886 107 -886 0 3
rlabel polysilicon 114 -880 114 -880 0 1
rlabel polysilicon 117 -880 117 -880 0 2
rlabel polysilicon 121 -880 121 -880 0 1
rlabel polysilicon 124 -886 124 -886 0 4
rlabel polysilicon 128 -880 128 -880 0 1
rlabel polysilicon 128 -886 128 -886 0 3
rlabel polysilicon 138 -886 138 -886 0 4
rlabel polysilicon 142 -880 142 -880 0 1
rlabel polysilicon 142 -886 142 -886 0 3
rlabel polysilicon 149 -880 149 -880 0 1
rlabel polysilicon 149 -886 149 -886 0 3
rlabel polysilicon 156 -880 156 -880 0 1
rlabel polysilicon 156 -886 156 -886 0 3
rlabel polysilicon 159 -886 159 -886 0 4
rlabel polysilicon 163 -880 163 -880 0 1
rlabel polysilicon 163 -886 163 -886 0 3
rlabel polysilicon 166 -886 166 -886 0 4
rlabel polysilicon 173 -880 173 -880 0 2
rlabel polysilicon 170 -886 170 -886 0 3
rlabel polysilicon 180 -880 180 -880 0 2
rlabel polysilicon 180 -886 180 -886 0 4
rlabel polysilicon 184 -880 184 -880 0 1
rlabel polysilicon 184 -886 184 -886 0 3
rlabel polysilicon 194 -880 194 -880 0 2
rlabel polysilicon 191 -886 191 -886 0 3
rlabel polysilicon 194 -886 194 -886 0 4
rlabel polysilicon 201 -880 201 -880 0 2
rlabel polysilicon 201 -886 201 -886 0 4
rlabel polysilicon 205 -886 205 -886 0 3
rlabel polysilicon 208 -886 208 -886 0 4
rlabel polysilicon 212 -880 212 -880 0 1
rlabel polysilicon 212 -886 212 -886 0 3
rlabel polysilicon 219 -880 219 -880 0 1
rlabel polysilicon 219 -886 219 -886 0 3
rlabel polysilicon 226 -880 226 -880 0 1
rlabel polysilicon 226 -886 226 -886 0 3
rlabel polysilicon 233 -880 233 -880 0 1
rlabel polysilicon 233 -886 233 -886 0 3
rlabel polysilicon 240 -880 240 -880 0 1
rlabel polysilicon 240 -886 240 -886 0 3
rlabel polysilicon 247 -880 247 -880 0 1
rlabel polysilicon 247 -886 247 -886 0 3
rlabel polysilicon 254 -880 254 -880 0 1
rlabel polysilicon 254 -886 254 -886 0 3
rlabel polysilicon 261 -880 261 -880 0 1
rlabel polysilicon 261 -886 261 -886 0 3
rlabel polysilicon 268 -880 268 -880 0 1
rlabel polysilicon 268 -886 268 -886 0 3
rlabel polysilicon 275 -880 275 -880 0 1
rlabel polysilicon 275 -886 275 -886 0 3
rlabel polysilicon 285 -880 285 -880 0 2
rlabel polysilicon 282 -886 282 -886 0 3
rlabel polysilicon 285 -886 285 -886 0 4
rlabel polysilicon 289 -880 289 -880 0 1
rlabel polysilicon 289 -886 289 -886 0 3
rlabel polysilicon 296 -880 296 -880 0 1
rlabel polysilicon 296 -886 296 -886 0 3
rlabel polysilicon 306 -880 306 -880 0 2
rlabel polysilicon 306 -886 306 -886 0 4
rlabel polysilicon 310 -880 310 -880 0 1
rlabel polysilicon 313 -880 313 -880 0 2
rlabel polysilicon 310 -886 310 -886 0 3
rlabel polysilicon 313 -886 313 -886 0 4
rlabel polysilicon 317 -880 317 -880 0 1
rlabel polysilicon 317 -886 317 -886 0 3
rlabel polysilicon 324 -880 324 -880 0 1
rlabel polysilicon 324 -886 324 -886 0 3
rlabel polysilicon 331 -880 331 -880 0 1
rlabel polysilicon 334 -880 334 -880 0 2
rlabel polysilicon 334 -886 334 -886 0 4
rlabel polysilicon 338 -880 338 -880 0 1
rlabel polysilicon 338 -886 338 -886 0 3
rlabel polysilicon 348 -880 348 -880 0 2
rlabel polysilicon 345 -886 345 -886 0 3
rlabel polysilicon 348 -886 348 -886 0 4
rlabel polysilicon 352 -880 352 -880 0 1
rlabel polysilicon 355 -880 355 -880 0 2
rlabel polysilicon 352 -886 352 -886 0 3
rlabel polysilicon 355 -886 355 -886 0 4
rlabel polysilicon 359 -880 359 -880 0 1
rlabel polysilicon 359 -886 359 -886 0 3
rlabel polysilicon 366 -880 366 -880 0 1
rlabel polysilicon 366 -886 366 -886 0 3
rlabel polysilicon 373 -880 373 -880 0 1
rlabel polysilicon 373 -886 373 -886 0 3
rlabel polysilicon 380 -886 380 -886 0 3
rlabel polysilicon 383 -886 383 -886 0 4
rlabel polysilicon 387 -880 387 -880 0 1
rlabel polysilicon 387 -886 387 -886 0 3
rlabel polysilicon 394 -880 394 -880 0 1
rlabel polysilicon 394 -886 394 -886 0 3
rlabel polysilicon 401 -880 401 -880 0 1
rlabel polysilicon 401 -886 401 -886 0 3
rlabel polysilicon 408 -880 408 -880 0 1
rlabel polysilicon 408 -886 408 -886 0 3
rlabel polysilicon 415 -880 415 -880 0 1
rlabel polysilicon 415 -886 415 -886 0 3
rlabel polysilicon 422 -880 422 -880 0 1
rlabel polysilicon 422 -886 422 -886 0 3
rlabel polysilicon 429 -880 429 -880 0 1
rlabel polysilicon 429 -886 429 -886 0 3
rlabel polysilicon 436 -880 436 -880 0 1
rlabel polysilicon 436 -886 436 -886 0 3
rlabel polysilicon 443 -880 443 -880 0 1
rlabel polysilicon 443 -886 443 -886 0 3
rlabel polysilicon 450 -880 450 -880 0 1
rlabel polysilicon 450 -886 450 -886 0 3
rlabel polysilicon 457 -880 457 -880 0 1
rlabel polysilicon 457 -886 457 -886 0 3
rlabel polysilicon 464 -880 464 -880 0 1
rlabel polysilicon 467 -880 467 -880 0 2
rlabel polysilicon 474 -880 474 -880 0 2
rlabel polysilicon 474 -886 474 -886 0 4
rlabel polysilicon 478 -880 478 -880 0 1
rlabel polysilicon 478 -886 478 -886 0 3
rlabel polysilicon 485 -880 485 -880 0 1
rlabel polysilicon 485 -886 485 -886 0 3
rlabel polysilicon 492 -880 492 -880 0 1
rlabel polysilicon 492 -886 492 -886 0 3
rlabel polysilicon 499 -880 499 -880 0 1
rlabel polysilicon 499 -886 499 -886 0 3
rlabel polysilicon 506 -880 506 -880 0 1
rlabel polysilicon 506 -886 506 -886 0 3
rlabel polysilicon 513 -880 513 -880 0 1
rlabel polysilicon 513 -886 513 -886 0 3
rlabel polysilicon 520 -886 520 -886 0 3
rlabel polysilicon 523 -886 523 -886 0 4
rlabel polysilicon 527 -880 527 -880 0 1
rlabel polysilicon 527 -886 527 -886 0 3
rlabel polysilicon 534 -880 534 -880 0 1
rlabel polysilicon 534 -886 534 -886 0 3
rlabel polysilicon 9 -935 9 -935 0 1
rlabel polysilicon 9 -941 9 -941 0 3
rlabel polysilicon 16 -935 16 -935 0 1
rlabel polysilicon 16 -941 16 -941 0 3
rlabel polysilicon 23 -935 23 -935 0 1
rlabel polysilicon 23 -941 23 -941 0 3
rlabel polysilicon 30 -941 30 -941 0 3
rlabel polysilicon 37 -935 37 -935 0 1
rlabel polysilicon 37 -941 37 -941 0 3
rlabel polysilicon 44 -935 44 -935 0 1
rlabel polysilicon 51 -935 51 -935 0 1
rlabel polysilicon 51 -941 51 -941 0 3
rlabel polysilicon 58 -935 58 -935 0 1
rlabel polysilicon 58 -941 58 -941 0 3
rlabel polysilicon 65 -935 65 -935 0 1
rlabel polysilicon 65 -941 65 -941 0 3
rlabel polysilicon 72 -935 72 -935 0 1
rlabel polysilicon 82 -941 82 -941 0 4
rlabel polysilicon 86 -941 86 -941 0 3
rlabel polysilicon 93 -935 93 -935 0 1
rlabel polysilicon 93 -941 93 -941 0 3
rlabel polysilicon 100 -941 100 -941 0 3
rlabel polysilicon 103 -941 103 -941 0 4
rlabel polysilicon 107 -935 107 -935 0 1
rlabel polysilicon 107 -941 107 -941 0 3
rlabel polysilicon 114 -935 114 -935 0 1
rlabel polysilicon 114 -941 114 -941 0 3
rlabel polysilicon 121 -935 121 -935 0 1
rlabel polysilicon 121 -941 121 -941 0 3
rlabel polysilicon 128 -935 128 -935 0 1
rlabel polysilicon 128 -941 128 -941 0 3
rlabel polysilicon 135 -935 135 -935 0 1
rlabel polysilicon 142 -935 142 -935 0 1
rlabel polysilicon 142 -941 142 -941 0 3
rlabel polysilicon 149 -935 149 -935 0 1
rlabel polysilicon 152 -935 152 -935 0 2
rlabel polysilicon 159 -935 159 -935 0 2
rlabel polysilicon 156 -941 156 -941 0 3
rlabel polysilicon 159 -941 159 -941 0 4
rlabel polysilicon 166 -935 166 -935 0 2
rlabel polysilicon 163 -941 163 -941 0 3
rlabel polysilicon 166 -941 166 -941 0 4
rlabel polysilicon 170 -935 170 -935 0 1
rlabel polysilicon 170 -941 170 -941 0 3
rlabel polysilicon 177 -935 177 -935 0 1
rlabel polysilicon 177 -941 177 -941 0 3
rlabel polysilicon 184 -935 184 -935 0 1
rlabel polysilicon 184 -941 184 -941 0 3
rlabel polysilicon 194 -935 194 -935 0 2
rlabel polysilicon 191 -941 191 -941 0 3
rlabel polysilicon 201 -935 201 -935 0 2
rlabel polysilicon 198 -941 198 -941 0 3
rlabel polysilicon 201 -941 201 -941 0 4
rlabel polysilicon 205 -935 205 -935 0 1
rlabel polysilicon 208 -935 208 -935 0 2
rlabel polysilicon 205 -941 205 -941 0 3
rlabel polysilicon 212 -935 212 -935 0 1
rlabel polysilicon 212 -941 212 -941 0 3
rlabel polysilicon 219 -935 219 -935 0 1
rlabel polysilicon 222 -935 222 -935 0 2
rlabel polysilicon 219 -941 219 -941 0 3
rlabel polysilicon 226 -935 226 -935 0 1
rlabel polysilicon 229 -935 229 -935 0 2
rlabel polysilicon 226 -941 226 -941 0 3
rlabel polysilicon 229 -941 229 -941 0 4
rlabel polysilicon 233 -935 233 -935 0 1
rlabel polysilicon 233 -941 233 -941 0 3
rlabel polysilicon 240 -935 240 -935 0 1
rlabel polysilicon 240 -941 240 -941 0 3
rlabel polysilicon 247 -935 247 -935 0 1
rlabel polysilicon 247 -941 247 -941 0 3
rlabel polysilicon 254 -935 254 -935 0 1
rlabel polysilicon 254 -941 254 -941 0 3
rlabel polysilicon 264 -935 264 -935 0 2
rlabel polysilicon 264 -941 264 -941 0 4
rlabel polysilicon 268 -935 268 -935 0 1
rlabel polysilicon 268 -941 268 -941 0 3
rlabel polysilicon 275 -935 275 -935 0 1
rlabel polysilicon 275 -941 275 -941 0 3
rlabel polysilicon 282 -935 282 -935 0 1
rlabel polysilicon 282 -941 282 -941 0 3
rlabel polysilicon 292 -935 292 -935 0 2
rlabel polysilicon 289 -941 289 -941 0 3
rlabel polysilicon 296 -935 296 -935 0 1
rlabel polysilicon 296 -941 296 -941 0 3
rlabel polysilicon 306 -935 306 -935 0 2
rlabel polysilicon 306 -941 306 -941 0 4
rlabel polysilicon 310 -935 310 -935 0 1
rlabel polysilicon 310 -941 310 -941 0 3
rlabel polysilicon 317 -935 317 -935 0 1
rlabel polysilicon 317 -941 317 -941 0 3
rlabel polysilicon 324 -935 324 -935 0 1
rlabel polysilicon 324 -941 324 -941 0 3
rlabel polysilicon 327 -941 327 -941 0 4
rlabel polysilicon 331 -935 331 -935 0 1
rlabel polysilicon 334 -935 334 -935 0 2
rlabel polysilicon 334 -941 334 -941 0 4
rlabel polysilicon 338 -935 338 -935 0 1
rlabel polysilicon 338 -941 338 -941 0 3
rlabel polysilicon 345 -935 345 -935 0 1
rlabel polysilicon 345 -941 345 -941 0 3
rlabel polysilicon 352 -941 352 -941 0 3
rlabel polysilicon 359 -935 359 -935 0 1
rlabel polysilicon 359 -941 359 -941 0 3
rlabel polysilicon 366 -935 366 -935 0 1
rlabel polysilicon 366 -941 366 -941 0 3
rlabel polysilicon 373 -935 373 -935 0 1
rlabel polysilicon 373 -941 373 -941 0 3
rlabel polysilicon 380 -935 380 -935 0 1
rlabel polysilicon 387 -935 387 -935 0 1
rlabel polysilicon 387 -941 387 -941 0 3
rlabel polysilicon 397 -935 397 -935 0 2
rlabel polysilicon 394 -941 394 -941 0 3
rlabel polysilicon 401 -935 401 -935 0 1
rlabel polysilicon 401 -941 401 -941 0 3
rlabel polysilicon 408 -935 408 -935 0 1
rlabel polysilicon 415 -935 415 -935 0 1
rlabel polysilicon 415 -941 415 -941 0 3
rlabel polysilicon 422 -935 422 -935 0 1
rlabel polysilicon 422 -941 422 -941 0 3
rlabel polysilicon 429 -935 429 -935 0 1
rlabel polysilicon 429 -941 429 -941 0 3
rlabel polysilicon 436 -935 436 -935 0 1
rlabel polysilicon 436 -941 436 -941 0 3
rlabel polysilicon 443 -941 443 -941 0 3
rlabel polysilicon 450 -935 450 -935 0 1
rlabel polysilicon 450 -941 450 -941 0 3
rlabel polysilicon 457 -935 457 -935 0 1
rlabel polysilicon 457 -941 457 -941 0 3
rlabel polysilicon 464 -941 464 -941 0 3
rlabel polysilicon 471 -935 471 -935 0 1
rlabel polysilicon 471 -941 471 -941 0 3
rlabel polysilicon 478 -935 478 -935 0 1
rlabel polysilicon 478 -941 478 -941 0 3
rlabel polysilicon 485 -935 485 -935 0 1
rlabel polysilicon 485 -941 485 -941 0 3
rlabel polysilicon 492 -935 492 -935 0 1
rlabel polysilicon 492 -941 492 -941 0 3
rlabel polysilicon 499 -935 499 -935 0 1
rlabel polysilicon 499 -941 499 -941 0 3
rlabel polysilicon 506 -935 506 -935 0 1
rlabel polysilicon 506 -941 506 -941 0 3
rlabel polysilicon 513 -935 513 -935 0 1
rlabel polysilicon 513 -941 513 -941 0 3
rlabel polysilicon 520 -935 520 -935 0 1
rlabel polysilicon 520 -941 520 -941 0 3
rlabel polysilicon 2 -984 2 -984 0 1
rlabel polysilicon 2 -990 2 -990 0 3
rlabel polysilicon 9 -984 9 -984 0 1
rlabel polysilicon 9 -990 9 -990 0 3
rlabel polysilicon 16 -984 16 -984 0 1
rlabel polysilicon 16 -990 16 -990 0 3
rlabel polysilicon 23 -984 23 -984 0 1
rlabel polysilicon 30 -984 30 -984 0 1
rlabel polysilicon 33 -990 33 -990 0 4
rlabel polysilicon 37 -990 37 -990 0 3
rlabel polysilicon 40 -990 40 -990 0 4
rlabel polysilicon 44 -984 44 -984 0 1
rlabel polysilicon 44 -990 44 -990 0 3
rlabel polysilicon 51 -984 51 -984 0 1
rlabel polysilicon 51 -990 51 -990 0 3
rlabel polysilicon 58 -990 58 -990 0 3
rlabel polysilicon 61 -990 61 -990 0 4
rlabel polysilicon 65 -984 65 -984 0 1
rlabel polysilicon 65 -990 65 -990 0 3
rlabel polysilicon 75 -984 75 -984 0 2
rlabel polysilicon 79 -990 79 -990 0 3
rlabel polysilicon 82 -990 82 -990 0 4
rlabel polysilicon 86 -984 86 -984 0 1
rlabel polysilicon 86 -990 86 -990 0 3
rlabel polysilicon 96 -984 96 -984 0 2
rlabel polysilicon 93 -990 93 -990 0 3
rlabel polysilicon 96 -990 96 -990 0 4
rlabel polysilicon 103 -984 103 -984 0 2
rlabel polysilicon 103 -990 103 -990 0 4
rlabel polysilicon 107 -984 107 -984 0 1
rlabel polysilicon 107 -990 107 -990 0 3
rlabel polysilicon 114 -984 114 -984 0 1
rlabel polysilicon 114 -990 114 -990 0 3
rlabel polysilicon 121 -984 121 -984 0 1
rlabel polysilicon 121 -990 121 -990 0 3
rlabel polysilicon 128 -990 128 -990 0 3
rlabel polysilicon 131 -990 131 -990 0 4
rlabel polysilicon 135 -984 135 -984 0 1
rlabel polysilicon 138 -984 138 -984 0 2
rlabel polysilicon 142 -984 142 -984 0 1
rlabel polysilicon 142 -990 142 -990 0 3
rlabel polysilicon 149 -984 149 -984 0 1
rlabel polysilicon 149 -990 149 -990 0 3
rlabel polysilicon 159 -984 159 -984 0 2
rlabel polysilicon 159 -990 159 -990 0 4
rlabel polysilicon 163 -984 163 -984 0 1
rlabel polysilicon 166 -984 166 -984 0 2
rlabel polysilicon 163 -990 163 -990 0 3
rlabel polysilicon 170 -984 170 -984 0 1
rlabel polysilicon 170 -990 170 -990 0 3
rlabel polysilicon 177 -984 177 -984 0 1
rlabel polysilicon 177 -990 177 -990 0 3
rlabel polysilicon 184 -984 184 -984 0 1
rlabel polysilicon 187 -984 187 -984 0 2
rlabel polysilicon 184 -990 184 -990 0 3
rlabel polysilicon 187 -990 187 -990 0 4
rlabel polysilicon 191 -984 191 -984 0 1
rlabel polysilicon 194 -984 194 -984 0 2
rlabel polysilicon 191 -990 191 -990 0 3
rlabel polysilicon 194 -990 194 -990 0 4
rlabel polysilicon 198 -984 198 -984 0 1
rlabel polysilicon 201 -984 201 -984 0 2
rlabel polysilicon 198 -990 198 -990 0 3
rlabel polysilicon 205 -984 205 -984 0 1
rlabel polysilicon 205 -990 205 -990 0 3
rlabel polysilicon 212 -984 212 -984 0 1
rlabel polysilicon 212 -990 212 -990 0 3
rlabel polysilicon 219 -984 219 -984 0 1
rlabel polysilicon 222 -984 222 -984 0 2
rlabel polysilicon 219 -990 219 -990 0 3
rlabel polysilicon 222 -990 222 -990 0 4
rlabel polysilicon 226 -990 226 -990 0 3
rlabel polysilicon 229 -990 229 -990 0 4
rlabel polysilicon 233 -984 233 -984 0 1
rlabel polysilicon 243 -990 243 -990 0 4
rlabel polysilicon 247 -984 247 -984 0 1
rlabel polysilicon 247 -990 247 -990 0 3
rlabel polysilicon 257 -984 257 -984 0 2
rlabel polysilicon 254 -990 254 -990 0 3
rlabel polysilicon 261 -984 261 -984 0 1
rlabel polysilicon 264 -984 264 -984 0 2
rlabel polysilicon 261 -990 261 -990 0 3
rlabel polysilicon 268 -984 268 -984 0 1
rlabel polysilicon 268 -990 268 -990 0 3
rlabel polysilicon 275 -984 275 -984 0 1
rlabel polysilicon 275 -990 275 -990 0 3
rlabel polysilicon 282 -984 282 -984 0 1
rlabel polysilicon 282 -990 282 -990 0 3
rlabel polysilicon 292 -984 292 -984 0 2
rlabel polysilicon 289 -990 289 -990 0 3
rlabel polysilicon 292 -990 292 -990 0 4
rlabel polysilicon 296 -984 296 -984 0 1
rlabel polysilicon 299 -984 299 -984 0 2
rlabel polysilicon 303 -984 303 -984 0 1
rlabel polysilicon 303 -990 303 -990 0 3
rlabel polysilicon 310 -984 310 -984 0 1
rlabel polysilicon 310 -990 310 -990 0 3
rlabel polysilicon 317 -984 317 -984 0 1
rlabel polysilicon 317 -990 317 -990 0 3
rlabel polysilicon 324 -984 324 -984 0 1
rlabel polysilicon 324 -990 324 -990 0 3
rlabel polysilicon 331 -984 331 -984 0 1
rlabel polysilicon 334 -984 334 -984 0 2
rlabel polysilicon 338 -984 338 -984 0 1
rlabel polysilicon 338 -990 338 -990 0 3
rlabel polysilicon 341 -990 341 -990 0 4
rlabel polysilicon 345 -984 345 -984 0 1
rlabel polysilicon 345 -990 345 -990 0 3
rlabel polysilicon 355 -984 355 -984 0 2
rlabel polysilicon 352 -990 352 -990 0 3
rlabel polysilicon 359 -984 359 -984 0 1
rlabel polysilicon 359 -990 359 -990 0 3
rlabel polysilicon 366 -984 366 -984 0 1
rlabel polysilicon 366 -990 366 -990 0 3
rlabel polysilicon 373 -984 373 -984 0 1
rlabel polysilicon 373 -990 373 -990 0 3
rlabel polysilicon 380 -984 380 -984 0 1
rlabel polysilicon 380 -990 380 -990 0 3
rlabel polysilicon 387 -984 387 -984 0 1
rlabel polysilicon 387 -990 387 -990 0 3
rlabel polysilicon 394 -984 394 -984 0 1
rlabel polysilicon 394 -990 394 -990 0 3
rlabel polysilicon 401 -984 401 -984 0 1
rlabel polysilicon 401 -990 401 -990 0 3
rlabel polysilicon 408 -984 408 -984 0 1
rlabel polysilicon 408 -990 408 -990 0 3
rlabel polysilicon 415 -984 415 -984 0 1
rlabel polysilicon 415 -990 415 -990 0 3
rlabel polysilicon 422 -984 422 -984 0 1
rlabel polysilicon 422 -990 422 -990 0 3
rlabel polysilicon 429 -984 429 -984 0 1
rlabel polysilicon 429 -990 429 -990 0 3
rlabel polysilicon 436 -984 436 -984 0 1
rlabel polysilicon 436 -990 436 -990 0 3
rlabel polysilicon 443 -984 443 -984 0 1
rlabel polysilicon 443 -990 443 -990 0 3
rlabel polysilicon 450 -984 450 -984 0 1
rlabel polysilicon 450 -990 450 -990 0 3
rlabel polysilicon 457 -984 457 -984 0 1
rlabel polysilicon 457 -990 457 -990 0 3
rlabel polysilicon 467 -984 467 -984 0 2
rlabel polysilicon 464 -990 464 -990 0 3
rlabel polysilicon 471 -984 471 -984 0 1
rlabel polysilicon 474 -990 474 -990 0 4
rlabel polysilicon 478 -984 478 -984 0 1
rlabel polysilicon 478 -990 478 -990 0 3
rlabel polysilicon 492 -984 492 -984 0 1
rlabel polysilicon 492 -990 492 -990 0 3
rlabel polysilicon 506 -984 506 -984 0 1
rlabel polysilicon 506 -990 506 -990 0 3
rlabel polysilicon 16 -1031 16 -1031 0 1
rlabel polysilicon 23 -1031 23 -1031 0 1
rlabel polysilicon 23 -1037 23 -1037 0 3
rlabel polysilicon 33 -1037 33 -1037 0 4
rlabel polysilicon 37 -1031 37 -1031 0 1
rlabel polysilicon 37 -1037 37 -1037 0 3
rlabel polysilicon 47 -1031 47 -1031 0 2
rlabel polysilicon 58 -1031 58 -1031 0 1
rlabel polysilicon 58 -1037 58 -1037 0 3
rlabel polysilicon 82 -1031 82 -1031 0 2
rlabel polysilicon 79 -1037 79 -1037 0 3
rlabel polysilicon 86 -1031 86 -1031 0 1
rlabel polysilicon 86 -1037 86 -1037 0 3
rlabel polysilicon 93 -1031 93 -1031 0 1
rlabel polysilicon 96 -1037 96 -1037 0 4
rlabel polysilicon 100 -1037 100 -1037 0 3
rlabel polysilicon 107 -1031 107 -1031 0 1
rlabel polysilicon 107 -1037 107 -1037 0 3
rlabel polysilicon 114 -1031 114 -1031 0 1
rlabel polysilicon 114 -1037 114 -1037 0 3
rlabel polysilicon 121 -1031 121 -1031 0 1
rlabel polysilicon 121 -1037 121 -1037 0 3
rlabel polysilicon 128 -1031 128 -1031 0 1
rlabel polysilicon 128 -1037 128 -1037 0 3
rlabel polysilicon 135 -1037 135 -1037 0 3
rlabel polysilicon 138 -1037 138 -1037 0 4
rlabel polysilicon 142 -1031 142 -1031 0 1
rlabel polysilicon 142 -1037 142 -1037 0 3
rlabel polysilicon 149 -1031 149 -1031 0 1
rlabel polysilicon 149 -1037 149 -1037 0 3
rlabel polysilicon 156 -1031 156 -1031 0 1
rlabel polysilicon 156 -1037 156 -1037 0 3
rlabel polysilicon 166 -1031 166 -1031 0 2
rlabel polysilicon 170 -1031 170 -1031 0 1
rlabel polysilicon 170 -1037 170 -1037 0 3
rlabel polysilicon 177 -1031 177 -1031 0 1
rlabel polysilicon 177 -1037 177 -1037 0 3
rlabel polysilicon 184 -1037 184 -1037 0 3
rlabel polysilicon 191 -1031 191 -1031 0 1
rlabel polysilicon 191 -1037 191 -1037 0 3
rlabel polysilicon 198 -1031 198 -1031 0 1
rlabel polysilicon 198 -1037 198 -1037 0 3
rlabel polysilicon 205 -1031 205 -1031 0 1
rlabel polysilicon 205 -1037 205 -1037 0 3
rlabel polysilicon 212 -1031 212 -1031 0 1
rlabel polysilicon 215 -1031 215 -1031 0 2
rlabel polysilicon 222 -1031 222 -1031 0 2
rlabel polysilicon 219 -1037 219 -1037 0 3
rlabel polysilicon 229 -1031 229 -1031 0 2
rlabel polysilicon 226 -1037 226 -1037 0 3
rlabel polysilicon 229 -1037 229 -1037 0 4
rlabel polysilicon 233 -1031 233 -1031 0 1
rlabel polysilicon 233 -1037 233 -1037 0 3
rlabel polysilicon 240 -1031 240 -1031 0 1
rlabel polysilicon 240 -1037 240 -1037 0 3
rlabel polysilicon 247 -1031 247 -1031 0 1
rlabel polysilicon 247 -1037 247 -1037 0 3
rlabel polysilicon 254 -1031 254 -1031 0 1
rlabel polysilicon 254 -1037 254 -1037 0 3
rlabel polysilicon 261 -1031 261 -1031 0 1
rlabel polysilicon 261 -1037 261 -1037 0 3
rlabel polysilicon 268 -1031 268 -1031 0 1
rlabel polysilicon 268 -1037 268 -1037 0 3
rlabel polysilicon 278 -1031 278 -1031 0 2
rlabel polysilicon 278 -1037 278 -1037 0 4
rlabel polysilicon 285 -1031 285 -1031 0 2
rlabel polysilicon 285 -1037 285 -1037 0 4
rlabel polysilicon 289 -1031 289 -1031 0 1
rlabel polysilicon 289 -1037 289 -1037 0 3
rlabel polysilicon 299 -1037 299 -1037 0 4
rlabel polysilicon 303 -1037 303 -1037 0 3
rlabel polysilicon 310 -1031 310 -1031 0 1
rlabel polysilicon 310 -1037 310 -1037 0 3
rlabel polysilicon 317 -1031 317 -1031 0 1
rlabel polysilicon 317 -1037 317 -1037 0 3
rlabel polysilicon 327 -1031 327 -1031 0 2
rlabel polysilicon 324 -1037 324 -1037 0 3
rlabel polysilicon 327 -1037 327 -1037 0 4
rlabel polysilicon 334 -1031 334 -1031 0 2
rlabel polysilicon 338 -1031 338 -1031 0 1
rlabel polysilicon 338 -1037 338 -1037 0 3
rlabel polysilicon 345 -1031 345 -1031 0 1
rlabel polysilicon 345 -1037 345 -1037 0 3
rlabel polysilicon 352 -1031 352 -1031 0 1
rlabel polysilicon 352 -1037 352 -1037 0 3
rlabel polysilicon 359 -1031 359 -1031 0 1
rlabel polysilicon 359 -1037 359 -1037 0 3
rlabel polysilicon 366 -1031 366 -1031 0 1
rlabel polysilicon 366 -1037 366 -1037 0 3
rlabel polysilicon 373 -1031 373 -1031 0 1
rlabel polysilicon 373 -1037 373 -1037 0 3
rlabel polysilicon 380 -1031 380 -1031 0 1
rlabel polysilicon 380 -1037 380 -1037 0 3
rlabel polysilicon 387 -1031 387 -1031 0 1
rlabel polysilicon 387 -1037 387 -1037 0 3
rlabel polysilicon 394 -1031 394 -1031 0 1
rlabel polysilicon 394 -1037 394 -1037 0 3
rlabel polysilicon 401 -1031 401 -1031 0 1
rlabel polysilicon 401 -1037 401 -1037 0 3
rlabel polysilicon 408 -1031 408 -1031 0 1
rlabel polysilicon 408 -1037 408 -1037 0 3
rlabel polysilicon 415 -1031 415 -1031 0 1
rlabel polysilicon 418 -1031 418 -1031 0 2
rlabel polysilicon 418 -1037 418 -1037 0 4
rlabel polysilicon 422 -1037 422 -1037 0 3
rlabel polysilicon 429 -1031 429 -1031 0 1
rlabel polysilicon 429 -1037 429 -1037 0 3
rlabel polysilicon 439 -1031 439 -1031 0 2
rlabel polysilicon 436 -1037 436 -1037 0 3
rlabel polysilicon 446 -1031 446 -1031 0 2
rlabel polysilicon 443 -1037 443 -1037 0 3
rlabel polysilicon 450 -1031 450 -1031 0 1
rlabel polysilicon 450 -1037 450 -1037 0 3
rlabel polysilicon 460 -1031 460 -1031 0 2
rlabel polysilicon 457 -1037 457 -1037 0 3
rlabel polysilicon 460 -1037 460 -1037 0 4
rlabel polysilicon 467 -1031 467 -1031 0 2
rlabel polysilicon 467 -1037 467 -1037 0 4
rlabel polysilicon 471 -1031 471 -1031 0 1
rlabel polysilicon 471 -1037 471 -1037 0 3
rlabel polysilicon 478 -1031 478 -1031 0 1
rlabel polysilicon 478 -1037 478 -1037 0 3
rlabel polysilicon 488 -1031 488 -1031 0 2
rlabel polysilicon 485 -1037 485 -1037 0 3
rlabel polysilicon 488 -1037 488 -1037 0 4
rlabel polysilicon 30 -1076 30 -1076 0 1
rlabel polysilicon 30 -1082 30 -1082 0 3
rlabel polysilicon 37 -1076 37 -1076 0 1
rlabel polysilicon 37 -1082 37 -1082 0 3
rlabel polysilicon 44 -1082 44 -1082 0 3
rlabel polysilicon 47 -1082 47 -1082 0 4
rlabel polysilicon 51 -1076 51 -1076 0 1
rlabel polysilicon 51 -1082 51 -1082 0 3
rlabel polysilicon 58 -1082 58 -1082 0 3
rlabel polysilicon 61 -1082 61 -1082 0 4
rlabel polysilicon 68 -1076 68 -1076 0 2
rlabel polysilicon 65 -1082 65 -1082 0 3
rlabel polysilicon 72 -1076 72 -1076 0 1
rlabel polysilicon 72 -1082 72 -1082 0 3
rlabel polysilicon 79 -1076 79 -1076 0 1
rlabel polysilicon 79 -1082 79 -1082 0 3
rlabel polysilicon 86 -1076 86 -1076 0 1
rlabel polysilicon 86 -1082 86 -1082 0 3
rlabel polysilicon 96 -1076 96 -1076 0 2
rlabel polysilicon 96 -1082 96 -1082 0 4
rlabel polysilicon 100 -1076 100 -1076 0 1
rlabel polysilicon 100 -1082 100 -1082 0 3
rlabel polysilicon 110 -1076 110 -1076 0 2
rlabel polysilicon 110 -1082 110 -1082 0 4
rlabel polysilicon 114 -1076 114 -1076 0 1
rlabel polysilicon 117 -1076 117 -1076 0 2
rlabel polysilicon 121 -1076 121 -1076 0 1
rlabel polysilicon 121 -1082 121 -1082 0 3
rlabel polysilicon 128 -1076 128 -1076 0 1
rlabel polysilicon 128 -1082 128 -1082 0 3
rlabel polysilicon 135 -1076 135 -1076 0 1
rlabel polysilicon 135 -1082 135 -1082 0 3
rlabel polysilicon 142 -1076 142 -1076 0 1
rlabel polysilicon 145 -1082 145 -1082 0 4
rlabel polysilicon 149 -1076 149 -1076 0 1
rlabel polysilicon 149 -1082 149 -1082 0 3
rlabel polysilicon 156 -1076 156 -1076 0 1
rlabel polysilicon 159 -1076 159 -1076 0 2
rlabel polysilicon 156 -1082 156 -1082 0 3
rlabel polysilicon 159 -1082 159 -1082 0 4
rlabel polysilicon 163 -1076 163 -1076 0 1
rlabel polysilicon 163 -1082 163 -1082 0 3
rlabel polysilicon 173 -1076 173 -1076 0 2
rlabel polysilicon 170 -1082 170 -1082 0 3
rlabel polysilicon 173 -1082 173 -1082 0 4
rlabel polysilicon 177 -1076 177 -1076 0 1
rlabel polysilicon 177 -1082 177 -1082 0 3
rlabel polysilicon 184 -1076 184 -1076 0 1
rlabel polysilicon 184 -1082 184 -1082 0 3
rlabel polysilicon 191 -1076 191 -1076 0 1
rlabel polysilicon 191 -1082 191 -1082 0 3
rlabel polysilicon 194 -1082 194 -1082 0 4
rlabel polysilicon 198 -1076 198 -1076 0 1
rlabel polysilicon 201 -1082 201 -1082 0 4
rlabel polysilicon 205 -1076 205 -1076 0 1
rlabel polysilicon 205 -1082 205 -1082 0 3
rlabel polysilicon 215 -1076 215 -1076 0 2
rlabel polysilicon 212 -1082 212 -1082 0 3
rlabel polysilicon 215 -1082 215 -1082 0 4
rlabel polysilicon 222 -1076 222 -1076 0 2
rlabel polysilicon 222 -1082 222 -1082 0 4
rlabel polysilicon 226 -1082 226 -1082 0 3
rlabel polysilicon 229 -1082 229 -1082 0 4
rlabel polysilicon 233 -1076 233 -1076 0 1
rlabel polysilicon 236 -1082 236 -1082 0 4
rlabel polysilicon 240 -1076 240 -1076 0 1
rlabel polysilicon 240 -1082 240 -1082 0 3
rlabel polysilicon 247 -1076 247 -1076 0 1
rlabel polysilicon 247 -1082 247 -1082 0 3
rlabel polysilicon 254 -1076 254 -1076 0 1
rlabel polysilicon 254 -1082 254 -1082 0 3
rlabel polysilicon 261 -1076 261 -1076 0 1
rlabel polysilicon 261 -1082 261 -1082 0 3
rlabel polysilicon 268 -1076 268 -1076 0 1
rlabel polysilicon 271 -1082 271 -1082 0 4
rlabel polysilicon 275 -1076 275 -1076 0 1
rlabel polysilicon 278 -1076 278 -1076 0 2
rlabel polysilicon 278 -1082 278 -1082 0 4
rlabel polysilicon 282 -1076 282 -1076 0 1
rlabel polysilicon 289 -1076 289 -1076 0 1
rlabel polysilicon 296 -1076 296 -1076 0 1
rlabel polysilicon 296 -1082 296 -1082 0 3
rlabel polysilicon 303 -1076 303 -1076 0 1
rlabel polysilicon 306 -1076 306 -1076 0 2
rlabel polysilicon 303 -1082 303 -1082 0 3
rlabel polysilicon 310 -1076 310 -1076 0 1
rlabel polysilicon 310 -1082 310 -1082 0 3
rlabel polysilicon 317 -1076 317 -1076 0 1
rlabel polysilicon 317 -1082 317 -1082 0 3
rlabel polysilicon 324 -1076 324 -1076 0 1
rlabel polysilicon 324 -1082 324 -1082 0 3
rlabel polysilicon 331 -1076 331 -1076 0 1
rlabel polysilicon 331 -1082 331 -1082 0 3
rlabel polysilicon 338 -1076 338 -1076 0 1
rlabel polysilicon 341 -1076 341 -1076 0 2
rlabel polysilicon 338 -1082 338 -1082 0 3
rlabel polysilicon 341 -1082 341 -1082 0 4
rlabel polysilicon 345 -1076 345 -1076 0 1
rlabel polysilicon 348 -1076 348 -1076 0 2
rlabel polysilicon 348 -1082 348 -1082 0 4
rlabel polysilicon 352 -1076 352 -1076 0 1
rlabel polysilicon 352 -1082 352 -1082 0 3
rlabel polysilicon 359 -1076 359 -1076 0 1
rlabel polysilicon 359 -1082 359 -1082 0 3
rlabel polysilicon 366 -1076 366 -1076 0 1
rlabel polysilicon 366 -1082 366 -1082 0 3
rlabel polysilicon 373 -1076 373 -1076 0 1
rlabel polysilicon 373 -1082 373 -1082 0 3
rlabel polysilicon 380 -1076 380 -1076 0 1
rlabel polysilicon 380 -1082 380 -1082 0 3
rlabel polysilicon 387 -1076 387 -1076 0 1
rlabel polysilicon 387 -1082 387 -1082 0 3
rlabel polysilicon 394 -1076 394 -1076 0 1
rlabel polysilicon 394 -1082 394 -1082 0 3
rlabel polysilicon 401 -1076 401 -1076 0 1
rlabel polysilicon 401 -1082 401 -1082 0 3
rlabel polysilicon 408 -1076 408 -1076 0 1
rlabel polysilicon 408 -1082 408 -1082 0 3
rlabel polysilicon 415 -1076 415 -1076 0 1
rlabel polysilicon 415 -1082 415 -1082 0 3
rlabel polysilicon 422 -1076 422 -1076 0 1
rlabel polysilicon 422 -1082 422 -1082 0 3
rlabel polysilicon 429 -1076 429 -1076 0 1
rlabel polysilicon 429 -1082 429 -1082 0 3
rlabel polysilicon 436 -1076 436 -1076 0 1
rlabel polysilicon 436 -1082 436 -1082 0 3
rlabel polysilicon 443 -1076 443 -1076 0 1
rlabel polysilicon 443 -1082 443 -1082 0 3
rlabel polysilicon 450 -1076 450 -1076 0 1
rlabel polysilicon 450 -1082 450 -1082 0 3
rlabel polysilicon 457 -1076 457 -1076 0 1
rlabel polysilicon 457 -1082 457 -1082 0 3
rlabel polysilicon 464 -1076 464 -1076 0 1
rlabel polysilicon 464 -1082 464 -1082 0 3
rlabel polysilicon 471 -1082 471 -1082 0 3
rlabel polysilicon 478 -1082 478 -1082 0 3
rlabel polysilicon 481 -1082 481 -1082 0 4
rlabel polysilicon 485 -1076 485 -1076 0 1
rlabel polysilicon 485 -1082 485 -1082 0 3
rlabel polysilicon 495 -1076 495 -1076 0 2
rlabel polysilicon 495 -1082 495 -1082 0 4
rlabel polysilicon 499 -1076 499 -1076 0 1
rlabel polysilicon 499 -1082 499 -1082 0 3
rlabel polysilicon 47 -1115 47 -1115 0 4
rlabel polysilicon 65 -1109 65 -1109 0 1
rlabel polysilicon 65 -1115 65 -1115 0 3
rlabel polysilicon 72 -1109 72 -1109 0 1
rlabel polysilicon 72 -1115 72 -1115 0 3
rlabel polysilicon 79 -1109 79 -1109 0 1
rlabel polysilicon 82 -1109 82 -1109 0 2
rlabel polysilicon 86 -1109 86 -1109 0 1
rlabel polysilicon 89 -1109 89 -1109 0 2
rlabel polysilicon 93 -1115 93 -1115 0 3
rlabel polysilicon 100 -1109 100 -1109 0 1
rlabel polysilicon 100 -1115 100 -1115 0 3
rlabel polysilicon 107 -1109 107 -1109 0 1
rlabel polysilicon 114 -1109 114 -1109 0 1
rlabel polysilicon 114 -1115 114 -1115 0 3
rlabel polysilicon 121 -1109 121 -1109 0 1
rlabel polysilicon 124 -1109 124 -1109 0 2
rlabel polysilicon 124 -1115 124 -1115 0 4
rlabel polysilicon 128 -1109 128 -1109 0 1
rlabel polysilicon 128 -1115 128 -1115 0 3
rlabel polysilicon 135 -1109 135 -1109 0 1
rlabel polysilicon 135 -1115 135 -1115 0 3
rlabel polysilicon 142 -1115 142 -1115 0 3
rlabel polysilicon 149 -1109 149 -1109 0 1
rlabel polysilicon 149 -1115 149 -1115 0 3
rlabel polysilicon 156 -1109 156 -1109 0 1
rlabel polysilicon 156 -1115 156 -1115 0 3
rlabel polysilicon 163 -1109 163 -1109 0 1
rlabel polysilicon 170 -1109 170 -1109 0 1
rlabel polysilicon 170 -1115 170 -1115 0 3
rlabel polysilicon 177 -1109 177 -1109 0 1
rlabel polysilicon 177 -1115 177 -1115 0 3
rlabel polysilicon 184 -1109 184 -1109 0 1
rlabel polysilicon 184 -1115 184 -1115 0 3
rlabel polysilicon 191 -1115 191 -1115 0 3
rlabel polysilicon 194 -1115 194 -1115 0 4
rlabel polysilicon 201 -1115 201 -1115 0 4
rlabel polysilicon 208 -1109 208 -1109 0 2
rlabel polysilicon 208 -1115 208 -1115 0 4
rlabel polysilicon 212 -1109 212 -1109 0 1
rlabel polysilicon 215 -1109 215 -1109 0 2
rlabel polysilicon 212 -1115 212 -1115 0 3
rlabel polysilicon 222 -1109 222 -1109 0 2
rlabel polysilicon 226 -1109 226 -1109 0 1
rlabel polysilicon 226 -1115 226 -1115 0 3
rlabel polysilicon 229 -1115 229 -1115 0 4
rlabel polysilicon 233 -1109 233 -1109 0 1
rlabel polysilicon 236 -1109 236 -1109 0 2
rlabel polysilicon 233 -1115 233 -1115 0 3
rlabel polysilicon 240 -1109 240 -1109 0 1
rlabel polysilicon 240 -1115 240 -1115 0 3
rlabel polysilicon 247 -1109 247 -1109 0 1
rlabel polysilicon 250 -1115 250 -1115 0 4
rlabel polysilicon 254 -1109 254 -1109 0 1
rlabel polysilicon 254 -1115 254 -1115 0 3
rlabel polysilicon 261 -1109 261 -1109 0 1
rlabel polysilicon 261 -1115 261 -1115 0 3
rlabel polysilicon 268 -1109 268 -1109 0 1
rlabel polysilicon 271 -1109 271 -1109 0 2
rlabel polysilicon 268 -1115 268 -1115 0 3
rlabel polysilicon 271 -1115 271 -1115 0 4
rlabel polysilicon 275 -1109 275 -1109 0 1
rlabel polysilicon 275 -1115 275 -1115 0 3
rlabel polysilicon 285 -1115 285 -1115 0 4
rlabel polysilicon 289 -1109 289 -1109 0 1
rlabel polysilicon 289 -1115 289 -1115 0 3
rlabel polysilicon 296 -1109 296 -1109 0 1
rlabel polysilicon 296 -1115 296 -1115 0 3
rlabel polysilicon 303 -1109 303 -1109 0 1
rlabel polysilicon 303 -1115 303 -1115 0 3
rlabel polysilicon 310 -1109 310 -1109 0 1
rlabel polysilicon 310 -1115 310 -1115 0 3
rlabel polysilicon 313 -1115 313 -1115 0 4
rlabel polysilicon 317 -1109 317 -1109 0 1
rlabel polysilicon 317 -1115 317 -1115 0 3
rlabel polysilicon 324 -1109 324 -1109 0 1
rlabel polysilicon 324 -1115 324 -1115 0 3
rlabel polysilicon 331 -1109 331 -1109 0 1
rlabel polysilicon 331 -1115 331 -1115 0 3
rlabel polysilicon 334 -1115 334 -1115 0 4
rlabel polysilicon 338 -1109 338 -1109 0 1
rlabel polysilicon 338 -1115 338 -1115 0 3
rlabel polysilicon 345 -1109 345 -1109 0 1
rlabel polysilicon 345 -1115 345 -1115 0 3
rlabel polysilicon 352 -1115 352 -1115 0 3
rlabel polysilicon 359 -1109 359 -1109 0 1
rlabel polysilicon 359 -1115 359 -1115 0 3
rlabel polysilicon 366 -1109 366 -1109 0 1
rlabel polysilicon 369 -1109 369 -1109 0 2
rlabel polysilicon 369 -1115 369 -1115 0 4
rlabel polysilicon 373 -1109 373 -1109 0 1
rlabel polysilicon 373 -1115 373 -1115 0 3
rlabel polysilicon 380 -1109 380 -1109 0 1
rlabel polysilicon 380 -1115 380 -1115 0 3
rlabel polysilicon 387 -1109 387 -1109 0 1
rlabel polysilicon 387 -1115 387 -1115 0 3
rlabel polysilicon 394 -1109 394 -1109 0 1
rlabel polysilicon 397 -1115 397 -1115 0 4
rlabel polysilicon 401 -1109 401 -1109 0 1
rlabel polysilicon 401 -1115 401 -1115 0 3
rlabel polysilicon 408 -1115 408 -1115 0 3
rlabel polysilicon 415 -1109 415 -1109 0 1
rlabel polysilicon 415 -1115 415 -1115 0 3
rlabel polysilicon 422 -1109 422 -1109 0 1
rlabel polysilicon 422 -1115 422 -1115 0 3
rlabel polysilicon 432 -1109 432 -1109 0 2
rlabel polysilicon 432 -1115 432 -1115 0 4
rlabel polysilicon 436 -1109 436 -1109 0 1
rlabel polysilicon 436 -1115 436 -1115 0 3
rlabel polysilicon 443 -1109 443 -1109 0 1
rlabel polysilicon 443 -1115 443 -1115 0 3
rlabel polysilicon 450 -1115 450 -1115 0 3
rlabel polysilicon 457 -1109 457 -1109 0 1
rlabel polysilicon 457 -1115 457 -1115 0 3
rlabel polysilicon 47 -1148 47 -1148 0 4
rlabel polysilicon 51 -1142 51 -1142 0 1
rlabel polysilicon 51 -1148 51 -1148 0 3
rlabel polysilicon 58 -1148 58 -1148 0 3
rlabel polysilicon 65 -1142 65 -1142 0 1
rlabel polysilicon 65 -1148 65 -1148 0 3
rlabel polysilicon 72 -1142 72 -1142 0 1
rlabel polysilicon 75 -1142 75 -1142 0 2
rlabel polysilicon 82 -1142 82 -1142 0 2
rlabel polysilicon 82 -1148 82 -1148 0 4
rlabel polysilicon 86 -1148 86 -1148 0 3
rlabel polysilicon 89 -1148 89 -1148 0 4
rlabel polysilicon 93 -1142 93 -1142 0 1
rlabel polysilicon 100 -1142 100 -1142 0 1
rlabel polysilicon 100 -1148 100 -1148 0 3
rlabel polysilicon 110 -1142 110 -1142 0 2
rlabel polysilicon 107 -1148 107 -1148 0 3
rlabel polysilicon 114 -1142 114 -1142 0 1
rlabel polysilicon 114 -1148 114 -1148 0 3
rlabel polysilicon 121 -1142 121 -1142 0 1
rlabel polysilicon 121 -1148 121 -1148 0 3
rlabel polysilicon 128 -1148 128 -1148 0 3
rlabel polysilicon 135 -1148 135 -1148 0 3
rlabel polysilicon 142 -1142 142 -1142 0 1
rlabel polysilicon 142 -1148 142 -1148 0 3
rlabel polysilicon 149 -1142 149 -1142 0 1
rlabel polysilicon 149 -1148 149 -1148 0 3
rlabel polysilicon 156 -1142 156 -1142 0 1
rlabel polysilicon 156 -1148 156 -1148 0 3
rlabel polysilicon 163 -1142 163 -1142 0 1
rlabel polysilicon 163 -1148 163 -1148 0 3
rlabel polysilicon 170 -1142 170 -1142 0 1
rlabel polysilicon 170 -1148 170 -1148 0 3
rlabel polysilicon 177 -1142 177 -1142 0 1
rlabel polysilicon 177 -1148 177 -1148 0 3
rlabel polysilicon 184 -1148 184 -1148 0 3
rlabel polysilicon 187 -1148 187 -1148 0 4
rlabel polysilicon 191 -1142 191 -1142 0 1
rlabel polysilicon 194 -1142 194 -1142 0 2
rlabel polysilicon 198 -1142 198 -1142 0 1
rlabel polysilicon 198 -1148 198 -1148 0 3
rlabel polysilicon 205 -1142 205 -1142 0 1
rlabel polysilicon 208 -1148 208 -1148 0 4
rlabel polysilicon 212 -1148 212 -1148 0 3
rlabel polysilicon 215 -1148 215 -1148 0 4
rlabel polysilicon 222 -1142 222 -1142 0 2
rlabel polysilicon 222 -1148 222 -1148 0 4
rlabel polysilicon 226 -1142 226 -1142 0 1
rlabel polysilicon 229 -1142 229 -1142 0 2
rlabel polysilicon 226 -1148 226 -1148 0 3
rlabel polysilicon 229 -1148 229 -1148 0 4
rlabel polysilicon 233 -1142 233 -1142 0 1
rlabel polysilicon 233 -1148 233 -1148 0 3
rlabel polysilicon 240 -1142 240 -1142 0 1
rlabel polysilicon 243 -1142 243 -1142 0 2
rlabel polysilicon 240 -1148 240 -1148 0 3
rlabel polysilicon 243 -1148 243 -1148 0 4
rlabel polysilicon 247 -1142 247 -1142 0 1
rlabel polysilicon 247 -1148 247 -1148 0 3
rlabel polysilicon 254 -1142 254 -1142 0 1
rlabel polysilicon 257 -1142 257 -1142 0 2
rlabel polysilicon 257 -1148 257 -1148 0 4
rlabel polysilicon 261 -1142 261 -1142 0 1
rlabel polysilicon 261 -1148 261 -1148 0 3
rlabel polysilicon 268 -1142 268 -1142 0 1
rlabel polysilicon 268 -1148 268 -1148 0 3
rlabel polysilicon 271 -1148 271 -1148 0 4
rlabel polysilicon 275 -1142 275 -1142 0 1
rlabel polysilicon 275 -1148 275 -1148 0 3
rlabel polysilicon 282 -1142 282 -1142 0 1
rlabel polysilicon 282 -1148 282 -1148 0 3
rlabel polysilicon 289 -1142 289 -1142 0 1
rlabel polysilicon 289 -1148 289 -1148 0 3
rlabel polysilicon 296 -1142 296 -1142 0 1
rlabel polysilicon 296 -1148 296 -1148 0 3
rlabel polysilicon 303 -1142 303 -1142 0 1
rlabel polysilicon 306 -1142 306 -1142 0 2
rlabel polysilicon 306 -1148 306 -1148 0 4
rlabel polysilicon 310 -1142 310 -1142 0 1
rlabel polysilicon 310 -1148 310 -1148 0 3
rlabel polysilicon 313 -1148 313 -1148 0 4
rlabel polysilicon 317 -1142 317 -1142 0 1
rlabel polysilicon 317 -1148 317 -1148 0 3
rlabel polysilicon 324 -1142 324 -1142 0 1
rlabel polysilicon 324 -1148 324 -1148 0 3
rlabel polysilicon 331 -1142 331 -1142 0 1
rlabel polysilicon 331 -1148 331 -1148 0 3
rlabel polysilicon 338 -1142 338 -1142 0 1
rlabel polysilicon 338 -1148 338 -1148 0 3
rlabel polysilicon 345 -1142 345 -1142 0 1
rlabel polysilicon 345 -1148 345 -1148 0 3
rlabel polysilicon 352 -1142 352 -1142 0 1
rlabel polysilicon 352 -1148 352 -1148 0 3
rlabel polysilicon 359 -1142 359 -1142 0 1
rlabel polysilicon 359 -1148 359 -1148 0 3
rlabel polysilicon 366 -1142 366 -1142 0 1
rlabel polysilicon 366 -1148 366 -1148 0 3
rlabel polysilicon 373 -1142 373 -1142 0 1
rlabel polysilicon 373 -1148 373 -1148 0 3
rlabel polysilicon 383 -1142 383 -1142 0 2
rlabel polysilicon 387 -1142 387 -1142 0 1
rlabel polysilicon 394 -1142 394 -1142 0 1
rlabel polysilicon 394 -1148 394 -1148 0 3
rlabel polysilicon 401 -1142 401 -1142 0 1
rlabel polysilicon 404 -1142 404 -1142 0 2
rlabel polysilicon 401 -1148 401 -1148 0 3
rlabel polysilicon 404 -1148 404 -1148 0 4
rlabel polysilicon 408 -1142 408 -1142 0 1
rlabel polysilicon 408 -1148 408 -1148 0 3
rlabel polysilicon 415 -1142 415 -1142 0 1
rlabel polysilicon 415 -1148 415 -1148 0 3
rlabel polysilicon 422 -1142 422 -1142 0 1
rlabel polysilicon 422 -1148 422 -1148 0 3
rlabel polysilicon 446 -1148 446 -1148 0 4
rlabel polysilicon 450 -1142 450 -1142 0 1
rlabel polysilicon 450 -1148 450 -1148 0 3
rlabel polysilicon 47 -1185 47 -1185 0 4
rlabel polysilicon 51 -1179 51 -1179 0 1
rlabel polysilicon 51 -1185 51 -1185 0 3
rlabel polysilicon 61 -1179 61 -1179 0 2
rlabel polysilicon 65 -1179 65 -1179 0 1
rlabel polysilicon 75 -1185 75 -1185 0 4
rlabel polysilicon 79 -1185 79 -1185 0 3
rlabel polysilicon 89 -1185 89 -1185 0 4
rlabel polysilicon 93 -1185 93 -1185 0 3
rlabel polysilicon 100 -1179 100 -1179 0 1
rlabel polysilicon 100 -1185 100 -1185 0 3
rlabel polysilicon 107 -1179 107 -1179 0 1
rlabel polysilicon 107 -1185 107 -1185 0 3
rlabel polysilicon 117 -1179 117 -1179 0 2
rlabel polysilicon 121 -1179 121 -1179 0 1
rlabel polysilicon 121 -1185 121 -1185 0 3
rlabel polysilicon 128 -1179 128 -1179 0 1
rlabel polysilicon 128 -1185 128 -1185 0 3
rlabel polysilicon 135 -1179 135 -1179 0 1
rlabel polysilicon 135 -1185 135 -1185 0 3
rlabel polysilicon 145 -1179 145 -1179 0 2
rlabel polysilicon 142 -1185 142 -1185 0 3
rlabel polysilicon 149 -1185 149 -1185 0 3
rlabel polysilicon 152 -1185 152 -1185 0 4
rlabel polysilicon 156 -1179 156 -1179 0 1
rlabel polysilicon 156 -1185 156 -1185 0 3
rlabel polysilicon 166 -1185 166 -1185 0 4
rlabel polysilicon 173 -1185 173 -1185 0 4
rlabel polysilicon 177 -1185 177 -1185 0 3
rlabel polysilicon 184 -1179 184 -1179 0 1
rlabel polysilicon 184 -1185 184 -1185 0 3
rlabel polysilicon 191 -1179 191 -1179 0 1
rlabel polysilicon 194 -1179 194 -1179 0 2
rlabel polysilicon 191 -1185 191 -1185 0 3
rlabel polysilicon 201 -1185 201 -1185 0 4
rlabel polysilicon 205 -1179 205 -1179 0 1
rlabel polysilicon 205 -1185 205 -1185 0 3
rlabel polysilicon 212 -1179 212 -1179 0 1
rlabel polysilicon 212 -1185 212 -1185 0 3
rlabel polysilicon 222 -1185 222 -1185 0 4
rlabel polysilicon 226 -1179 226 -1179 0 1
rlabel polysilicon 226 -1185 226 -1185 0 3
rlabel polysilicon 229 -1185 229 -1185 0 4
rlabel polysilicon 233 -1179 233 -1179 0 1
rlabel polysilicon 236 -1179 236 -1179 0 2
rlabel polysilicon 236 -1185 236 -1185 0 4
rlabel polysilicon 243 -1179 243 -1179 0 2
rlabel polysilicon 240 -1185 240 -1185 0 3
rlabel polysilicon 247 -1179 247 -1179 0 1
rlabel polysilicon 254 -1179 254 -1179 0 1
rlabel polysilicon 261 -1179 261 -1179 0 1
rlabel polysilicon 261 -1185 261 -1185 0 3
rlabel polysilicon 268 -1179 268 -1179 0 1
rlabel polysilicon 268 -1185 268 -1185 0 3
rlabel polysilicon 275 -1179 275 -1179 0 1
rlabel polysilicon 275 -1185 275 -1185 0 3
rlabel polysilicon 282 -1179 282 -1179 0 1
rlabel polysilicon 282 -1185 282 -1185 0 3
rlabel polysilicon 289 -1185 289 -1185 0 3
rlabel polysilicon 292 -1185 292 -1185 0 4
rlabel polysilicon 296 -1179 296 -1179 0 1
rlabel polysilicon 299 -1179 299 -1179 0 2
rlabel polysilicon 303 -1179 303 -1179 0 1
rlabel polysilicon 303 -1185 303 -1185 0 3
rlabel polysilicon 310 -1179 310 -1179 0 1
rlabel polysilicon 310 -1185 310 -1185 0 3
rlabel polysilicon 317 -1179 317 -1179 0 1
rlabel polysilicon 317 -1185 317 -1185 0 3
rlabel polysilicon 324 -1179 324 -1179 0 1
rlabel polysilicon 324 -1185 324 -1185 0 3
rlabel polysilicon 331 -1179 331 -1179 0 1
rlabel polysilicon 331 -1185 331 -1185 0 3
rlabel polysilicon 338 -1179 338 -1179 0 1
rlabel polysilicon 338 -1185 338 -1185 0 3
rlabel polysilicon 345 -1185 345 -1185 0 3
rlabel polysilicon 348 -1185 348 -1185 0 4
rlabel polysilicon 352 -1179 352 -1179 0 1
rlabel polysilicon 352 -1185 352 -1185 0 3
rlabel polysilicon 359 -1179 359 -1179 0 1
rlabel polysilicon 359 -1185 359 -1185 0 3
rlabel polysilicon 366 -1179 366 -1179 0 1
rlabel polysilicon 366 -1185 366 -1185 0 3
rlabel polysilicon 373 -1179 373 -1179 0 1
rlabel polysilicon 373 -1185 373 -1185 0 3
rlabel polysilicon 380 -1179 380 -1179 0 1
rlabel polysilicon 380 -1185 380 -1185 0 3
rlabel polysilicon 387 -1179 387 -1179 0 1
rlabel polysilicon 387 -1185 387 -1185 0 3
rlabel polysilicon 394 -1179 394 -1179 0 1
rlabel polysilicon 394 -1185 394 -1185 0 3
rlabel polysilicon 401 -1179 401 -1179 0 1
rlabel polysilicon 401 -1185 401 -1185 0 3
rlabel polysilicon 415 -1179 415 -1179 0 1
rlabel polysilicon 418 -1179 418 -1179 0 2
rlabel polysilicon 415 -1185 415 -1185 0 3
rlabel polysilicon 422 -1179 422 -1179 0 1
rlabel polysilicon 422 -1185 422 -1185 0 3
rlabel polysilicon 429 -1179 429 -1179 0 1
rlabel polysilicon 429 -1185 429 -1185 0 3
rlabel polysilicon 47 -1206 47 -1206 0 2
rlabel polysilicon 65 -1206 65 -1206 0 1
rlabel polysilicon 68 -1206 68 -1206 0 2
rlabel polysilicon 72 -1206 72 -1206 0 1
rlabel polysilicon 72 -1212 72 -1212 0 3
rlabel polysilicon 79 -1206 79 -1206 0 1
rlabel polysilicon 82 -1206 82 -1206 0 2
rlabel polysilicon 79 -1212 79 -1212 0 3
rlabel polysilicon 89 -1212 89 -1212 0 4
rlabel polysilicon 96 -1206 96 -1206 0 2
rlabel polysilicon 100 -1206 100 -1206 0 1
rlabel polysilicon 100 -1212 100 -1212 0 3
rlabel polysilicon 107 -1206 107 -1206 0 1
rlabel polysilicon 107 -1212 107 -1212 0 3
rlabel polysilicon 114 -1206 114 -1206 0 1
rlabel polysilicon 114 -1212 114 -1212 0 3
rlabel polysilicon 121 -1206 121 -1206 0 1
rlabel polysilicon 121 -1212 121 -1212 0 3
rlabel polysilicon 128 -1206 128 -1206 0 1
rlabel polysilicon 128 -1212 128 -1212 0 3
rlabel polysilicon 135 -1206 135 -1206 0 1
rlabel polysilicon 138 -1206 138 -1206 0 2
rlabel polysilicon 135 -1212 135 -1212 0 3
rlabel polysilicon 138 -1212 138 -1212 0 4
rlabel polysilicon 145 -1206 145 -1206 0 2
rlabel polysilicon 142 -1212 142 -1212 0 3
rlabel polysilicon 149 -1206 149 -1206 0 1
rlabel polysilicon 152 -1212 152 -1212 0 4
rlabel polysilicon 156 -1206 156 -1206 0 1
rlabel polysilicon 159 -1206 159 -1206 0 2
rlabel polysilicon 156 -1212 156 -1212 0 3
rlabel polysilicon 159 -1212 159 -1212 0 4
rlabel polysilicon 166 -1206 166 -1206 0 2
rlabel polysilicon 163 -1212 163 -1212 0 3
rlabel polysilicon 170 -1206 170 -1206 0 1
rlabel polysilicon 170 -1212 170 -1212 0 3
rlabel polysilicon 177 -1206 177 -1206 0 1
rlabel polysilicon 177 -1212 177 -1212 0 3
rlabel polysilicon 184 -1206 184 -1206 0 1
rlabel polysilicon 187 -1212 187 -1212 0 4
rlabel polysilicon 194 -1212 194 -1212 0 4
rlabel polysilicon 198 -1206 198 -1206 0 1
rlabel polysilicon 198 -1212 198 -1212 0 3
rlabel polysilicon 205 -1206 205 -1206 0 1
rlabel polysilicon 205 -1212 205 -1212 0 3
rlabel polysilicon 212 -1206 212 -1206 0 1
rlabel polysilicon 212 -1212 212 -1212 0 3
rlabel polysilicon 219 -1206 219 -1206 0 1
rlabel polysilicon 222 -1206 222 -1206 0 2
rlabel polysilicon 222 -1212 222 -1212 0 4
rlabel polysilicon 226 -1206 226 -1206 0 1
rlabel polysilicon 229 -1206 229 -1206 0 2
rlabel polysilicon 229 -1212 229 -1212 0 4
rlabel polysilicon 233 -1206 233 -1206 0 1
rlabel polysilicon 233 -1212 233 -1212 0 3
rlabel polysilicon 240 -1206 240 -1206 0 1
rlabel polysilicon 243 -1212 243 -1212 0 4
rlabel polysilicon 247 -1206 247 -1206 0 1
rlabel polysilicon 247 -1212 247 -1212 0 3
rlabel polysilicon 254 -1206 254 -1206 0 1
rlabel polysilicon 254 -1212 254 -1212 0 3
rlabel polysilicon 282 -1206 282 -1206 0 1
rlabel polysilicon 282 -1212 282 -1212 0 3
rlabel polysilicon 289 -1206 289 -1206 0 1
rlabel polysilicon 292 -1206 292 -1206 0 2
rlabel polysilicon 292 -1212 292 -1212 0 4
rlabel polysilicon 296 -1206 296 -1206 0 1
rlabel polysilicon 296 -1212 296 -1212 0 3
rlabel polysilicon 303 -1206 303 -1206 0 1
rlabel polysilicon 303 -1212 303 -1212 0 3
rlabel polysilicon 306 -1212 306 -1212 0 4
rlabel polysilicon 310 -1212 310 -1212 0 3
rlabel polysilicon 313 -1212 313 -1212 0 4
rlabel polysilicon 317 -1206 317 -1206 0 1
rlabel polysilicon 317 -1212 317 -1212 0 3
rlabel polysilicon 324 -1206 324 -1206 0 1
rlabel polysilicon 324 -1212 324 -1212 0 3
rlabel polysilicon 331 -1206 331 -1206 0 1
rlabel polysilicon 331 -1212 331 -1212 0 3
rlabel polysilicon 341 -1206 341 -1206 0 2
rlabel polysilicon 341 -1212 341 -1212 0 4
rlabel polysilicon 345 -1206 345 -1206 0 1
rlabel polysilicon 345 -1212 345 -1212 0 3
rlabel polysilicon 352 -1212 352 -1212 0 3
rlabel polysilicon 359 -1206 359 -1206 0 1
rlabel polysilicon 359 -1212 359 -1212 0 3
rlabel polysilicon 366 -1206 366 -1206 0 1
rlabel polysilicon 366 -1212 366 -1212 0 3
rlabel polysilicon 373 -1212 373 -1212 0 3
rlabel polysilicon 380 -1206 380 -1206 0 1
rlabel polysilicon 380 -1212 380 -1212 0 3
rlabel polysilicon 408 -1206 408 -1206 0 1
rlabel polysilicon 408 -1212 408 -1212 0 3
rlabel polysilicon 422 -1206 422 -1206 0 1
rlabel polysilicon 425 -1212 425 -1212 0 4
rlabel polysilicon 429 -1206 429 -1206 0 1
rlabel polysilicon 429 -1212 429 -1212 0 3
rlabel polysilicon 23 -1235 23 -1235 0 3
rlabel polysilicon 33 -1229 33 -1229 0 2
rlabel polysilicon 37 -1229 37 -1229 0 1
rlabel polysilicon 37 -1235 37 -1235 0 3
rlabel polysilicon 44 -1229 44 -1229 0 1
rlabel polysilicon 51 -1229 51 -1229 0 1
rlabel polysilicon 51 -1235 51 -1235 0 3
rlabel polysilicon 58 -1229 58 -1229 0 1
rlabel polysilicon 58 -1235 58 -1235 0 3
rlabel polysilicon 65 -1229 65 -1229 0 1
rlabel polysilicon 65 -1235 65 -1235 0 3
rlabel polysilicon 72 -1229 72 -1229 0 1
rlabel polysilicon 79 -1229 79 -1229 0 1
rlabel polysilicon 79 -1235 79 -1235 0 3
rlabel polysilicon 93 -1229 93 -1229 0 1
rlabel polysilicon 93 -1235 93 -1235 0 3
rlabel polysilicon 100 -1229 100 -1229 0 1
rlabel polysilicon 100 -1235 100 -1235 0 3
rlabel polysilicon 110 -1235 110 -1235 0 4
rlabel polysilicon 114 -1235 114 -1235 0 3
rlabel polysilicon 117 -1235 117 -1235 0 4
rlabel polysilicon 121 -1229 121 -1229 0 1
rlabel polysilicon 124 -1229 124 -1229 0 2
rlabel polysilicon 128 -1229 128 -1229 0 1
rlabel polysilicon 128 -1235 128 -1235 0 3
rlabel polysilicon 138 -1235 138 -1235 0 4
rlabel polysilicon 142 -1229 142 -1229 0 1
rlabel polysilicon 142 -1235 142 -1235 0 3
rlabel polysilicon 149 -1229 149 -1229 0 1
rlabel polysilicon 149 -1235 149 -1235 0 3
rlabel polysilicon 159 -1235 159 -1235 0 4
rlabel polysilicon 163 -1229 163 -1229 0 1
rlabel polysilicon 163 -1235 163 -1235 0 3
rlabel polysilicon 173 -1229 173 -1229 0 2
rlabel polysilicon 170 -1235 170 -1235 0 3
rlabel polysilicon 180 -1229 180 -1229 0 2
rlabel polysilicon 184 -1229 184 -1229 0 1
rlabel polysilicon 184 -1235 184 -1235 0 3
rlabel polysilicon 191 -1229 191 -1229 0 1
rlabel polysilicon 191 -1235 191 -1235 0 3
rlabel polysilicon 201 -1229 201 -1229 0 2
rlabel polysilicon 205 -1235 205 -1235 0 3
rlabel polysilicon 208 -1235 208 -1235 0 4
rlabel polysilicon 212 -1229 212 -1229 0 1
rlabel polysilicon 215 -1229 215 -1229 0 2
rlabel polysilicon 215 -1235 215 -1235 0 4
rlabel polysilicon 219 -1229 219 -1229 0 1
rlabel polysilicon 222 -1229 222 -1229 0 2
rlabel polysilicon 222 -1235 222 -1235 0 4
rlabel polysilicon 229 -1229 229 -1229 0 2
rlabel polysilicon 233 -1229 233 -1229 0 1
rlabel polysilicon 233 -1235 233 -1235 0 3
rlabel polysilicon 240 -1229 240 -1229 0 1
rlabel polysilicon 240 -1235 240 -1235 0 3
rlabel polysilicon 250 -1235 250 -1235 0 4
rlabel polysilicon 254 -1229 254 -1229 0 1
rlabel polysilicon 254 -1235 254 -1235 0 3
rlabel polysilicon 261 -1235 261 -1235 0 3
rlabel polysilicon 268 -1229 268 -1229 0 1
rlabel polysilicon 268 -1235 268 -1235 0 3
rlabel polysilicon 275 -1229 275 -1229 0 1
rlabel polysilicon 275 -1235 275 -1235 0 3
rlabel polysilicon 282 -1229 282 -1229 0 1
rlabel polysilicon 282 -1235 282 -1235 0 3
rlabel polysilicon 292 -1229 292 -1229 0 2
rlabel polysilicon 299 -1235 299 -1235 0 4
rlabel polysilicon 303 -1229 303 -1229 0 1
rlabel polysilicon 303 -1235 303 -1235 0 3
rlabel polysilicon 310 -1229 310 -1229 0 1
rlabel polysilicon 310 -1235 310 -1235 0 3
rlabel polysilicon 317 -1229 317 -1229 0 1
rlabel polysilicon 320 -1229 320 -1229 0 2
rlabel polysilicon 327 -1235 327 -1235 0 4
rlabel polysilicon 338 -1229 338 -1229 0 1
rlabel polysilicon 338 -1235 338 -1235 0 3
rlabel polysilicon 345 -1229 345 -1229 0 1
rlabel polysilicon 352 -1229 352 -1229 0 1
rlabel polysilicon 352 -1235 352 -1235 0 3
rlabel polysilicon 359 -1229 359 -1229 0 1
rlabel polysilicon 359 -1235 359 -1235 0 3
rlabel polysilicon 366 -1229 366 -1229 0 1
rlabel polysilicon 373 -1229 373 -1229 0 1
rlabel polysilicon 373 -1235 373 -1235 0 3
rlabel polysilicon 401 -1229 401 -1229 0 1
rlabel polysilicon 401 -1235 401 -1235 0 3
rlabel polysilicon 408 -1235 408 -1235 0 3
rlabel polysilicon 415 -1235 415 -1235 0 3
rlabel polysilicon 422 -1229 422 -1229 0 1
rlabel polysilicon 422 -1235 422 -1235 0 3
rlabel polysilicon 432 -1229 432 -1229 0 2
rlabel polysilicon 23 -1254 23 -1254 0 1
rlabel polysilicon 30 -1254 30 -1254 0 1
rlabel polysilicon 30 -1260 30 -1260 0 3
rlabel polysilicon 37 -1260 37 -1260 0 3
rlabel polysilicon 44 -1254 44 -1254 0 1
rlabel polysilicon 58 -1254 58 -1254 0 1
rlabel polysilicon 58 -1260 58 -1260 0 3
rlabel polysilicon 68 -1260 68 -1260 0 4
rlabel polysilicon 75 -1254 75 -1254 0 2
rlabel polysilicon 72 -1260 72 -1260 0 3
rlabel polysilicon 79 -1254 79 -1254 0 1
rlabel polysilicon 79 -1260 79 -1260 0 3
rlabel polysilicon 103 -1254 103 -1254 0 2
rlabel polysilicon 107 -1260 107 -1260 0 3
rlabel polysilicon 114 -1254 114 -1254 0 1
rlabel polysilicon 114 -1260 114 -1260 0 3
rlabel polysilicon 121 -1254 121 -1254 0 1
rlabel polysilicon 121 -1260 121 -1260 0 3
rlabel polysilicon 128 -1254 128 -1254 0 1
rlabel polysilicon 128 -1260 128 -1260 0 3
rlabel polysilicon 138 -1260 138 -1260 0 4
rlabel polysilicon 145 -1254 145 -1254 0 2
rlabel polysilicon 142 -1260 142 -1260 0 3
rlabel polysilicon 152 -1254 152 -1254 0 2
rlabel polysilicon 152 -1260 152 -1260 0 4
rlabel polysilicon 159 -1254 159 -1254 0 2
rlabel polysilicon 163 -1260 163 -1260 0 3
rlabel polysilicon 170 -1254 170 -1254 0 1
rlabel polysilicon 170 -1260 170 -1260 0 3
rlabel polysilicon 177 -1254 177 -1254 0 1
rlabel polysilicon 177 -1260 177 -1260 0 3
rlabel polysilicon 187 -1260 187 -1260 0 4
rlabel polysilicon 194 -1254 194 -1254 0 2
rlabel polysilicon 198 -1260 198 -1260 0 3
rlabel polysilicon 208 -1254 208 -1254 0 2
rlabel polysilicon 205 -1260 205 -1260 0 3
rlabel polysilicon 208 -1260 208 -1260 0 4
rlabel polysilicon 212 -1254 212 -1254 0 1
rlabel polysilicon 212 -1260 212 -1260 0 3
rlabel polysilicon 219 -1254 219 -1254 0 1
rlabel polysilicon 222 -1254 222 -1254 0 2
rlabel polysilicon 226 -1254 226 -1254 0 1
rlabel polysilicon 226 -1260 226 -1260 0 3
rlabel polysilicon 233 -1254 233 -1254 0 1
rlabel polysilicon 233 -1260 233 -1260 0 3
rlabel polysilicon 240 -1254 240 -1254 0 1
rlabel polysilicon 250 -1260 250 -1260 0 4
rlabel polysilicon 257 -1254 257 -1254 0 2
rlabel polysilicon 261 -1254 261 -1254 0 1
rlabel polysilicon 261 -1260 261 -1260 0 3
rlabel polysilicon 268 -1254 268 -1254 0 1
rlabel polysilicon 268 -1260 268 -1260 0 3
rlabel polysilicon 278 -1254 278 -1254 0 2
rlabel polysilicon 285 -1260 285 -1260 0 4
rlabel polysilicon 289 -1254 289 -1254 0 1
rlabel polysilicon 289 -1260 289 -1260 0 3
rlabel polysilicon 296 -1260 296 -1260 0 3
rlabel polysilicon 303 -1254 303 -1254 0 1
rlabel polysilicon 303 -1260 303 -1260 0 3
rlabel polysilicon 317 -1260 317 -1260 0 3
rlabel polysilicon 324 -1254 324 -1254 0 1
rlabel polysilicon 324 -1260 324 -1260 0 3
rlabel polysilicon 334 -1254 334 -1254 0 2
rlabel polysilicon 338 -1254 338 -1254 0 1
rlabel polysilicon 338 -1260 338 -1260 0 3
rlabel polysilicon 348 -1260 348 -1260 0 4
rlabel polysilicon 355 -1260 355 -1260 0 4
rlabel polysilicon 359 -1254 359 -1254 0 1
rlabel polysilicon 359 -1260 359 -1260 0 3
rlabel polysilicon 369 -1254 369 -1254 0 2
rlabel metal2 138 1 138 1 0 net=1615
rlabel metal2 177 1 177 1 0 net=1189
rlabel metal2 198 1 198 1 0 net=1019
rlabel metal2 226 1 226 1 0 net=1495
rlabel metal2 187 -1 187 -1 0 net=265
rlabel metal2 212 -1 212 -1 0 net=1667
rlabel metal2 135 -12 135 -12 0 net=2955
rlabel metal2 187 -12 187 -12 0 net=727
rlabel metal2 240 -12 240 -12 0 net=1496
rlabel metal2 324 -12 324 -12 0 net=2469
rlabel metal2 142 -14 142 -14 0 net=1747
rlabel metal2 142 -14 142 -14 0 net=1747
rlabel metal2 145 -14 145 -14 0 net=1616
rlabel metal2 163 -14 163 -14 0 net=1525
rlabel metal2 177 -14 177 -14 0 net=1190
rlabel metal2 191 -14 191 -14 0 net=2057
rlabel metal2 156 -16 156 -16 0 net=1791
rlabel metal2 198 -16 198 -16 0 net=1021
rlabel metal2 208 -16 208 -16 0 net=1668
rlabel metal2 226 -16 226 -16 0 net=251
rlabel metal2 198 -18 198 -18 0 net=1421
rlabel metal2 219 -18 219 -18 0 net=2259
rlabel metal2 229 -20 229 -20 0 net=217
rlabel metal2 128 -31 128 -31 0 net=244
rlabel metal2 198 -31 198 -31 0 net=1422
rlabel metal2 222 -31 222 -31 0 net=873
rlabel metal2 268 -31 268 -31 0 net=2987
rlabel metal2 296 -31 296 -31 0 net=2981
rlabel metal2 324 -31 324 -31 0 net=2471
rlabel metal2 135 -33 135 -33 0 net=2956
rlabel metal2 198 -33 198 -33 0 net=1969
rlabel metal2 327 -33 327 -33 0 net=2043
rlabel metal2 135 -35 135 -35 0 net=1925
rlabel metal2 201 -35 201 -35 0 net=2058
rlabel metal2 142 -37 142 -37 0 net=1748
rlabel metal2 173 -37 173 -37 0 net=1127
rlabel metal2 159 -39 159 -39 0 net=1792
rlabel metal2 205 -39 205 -39 0 net=1022
rlabel metal2 163 -41 163 -41 0 net=1526
rlabel metal2 205 -41 205 -41 0 net=2260
rlabel metal2 163 -43 163 -43 0 net=1363
rlabel metal2 208 -43 208 -43 0 net=1307
rlabel metal2 226 -43 226 -43 0 net=2617
rlabel metal2 229 -45 229 -45 0 net=941
rlabel metal2 191 -47 191 -47 0 net=1501
rlabel metal2 103 -58 103 -58 0 net=2171
rlabel metal2 121 -58 121 -58 0 net=1927
rlabel metal2 142 -58 142 -58 0 net=60
rlabel metal2 205 -58 205 -58 0 net=1309
rlabel metal2 226 -58 226 -58 0 net=1970
rlabel metal2 261 -58 261 -58 0 net=874
rlabel metal2 324 -58 324 -58 0 net=2473
rlabel metal2 324 -58 324 -58 0 net=2473
rlabel metal2 331 -58 331 -58 0 net=2045
rlabel metal2 331 -58 331 -58 0 net=2045
rlabel metal2 128 -60 128 -60 0 net=2451
rlabel metal2 191 -60 191 -60 0 net=1503
rlabel metal2 268 -60 268 -60 0 net=2618
rlabel metal2 289 -60 289 -60 0 net=2988
rlabel metal2 142 -62 142 -62 0 net=1087
rlabel metal2 184 -62 184 -62 0 net=1365
rlabel metal2 229 -62 229 -62 0 net=1128
rlabel metal2 240 -62 240 -62 0 net=942
rlabel metal2 275 -62 275 -62 0 net=2583
rlabel metal2 282 -62 282 -62 0 net=1997
rlabel metal2 177 -64 177 -64 0 net=1033
rlabel metal2 201 -64 201 -64 0 net=2187
rlabel metal2 296 -64 296 -64 0 net=2982
rlabel metal2 219 -66 219 -66 0 net=1955
rlabel metal2 292 -66 292 -66 0 net=2651
rlabel metal2 170 -68 170 -68 0 net=228
rlabel metal2 166 -70 166 -70 0 net=2279
rlabel metal2 89 -81 89 -81 0 net=527
rlabel metal2 89 -81 89 -81 0 net=527
rlabel metal2 100 -81 100 -81 0 net=2172
rlabel metal2 114 -81 114 -81 0 net=2557
rlabel metal2 138 -81 138 -81 0 net=1088
rlabel metal2 159 -81 159 -81 0 net=24
rlabel metal2 166 -81 166 -81 0 net=1034
rlabel metal2 184 -81 184 -81 0 net=1151
rlabel metal2 205 -81 205 -81 0 net=1310
rlabel metal2 229 -81 229 -81 0 net=1956
rlabel metal2 275 -81 275 -81 0 net=2585
rlabel metal2 317 -81 317 -81 0 net=2474
rlabel metal2 107 -83 107 -83 0 net=2453
rlabel metal2 149 -83 149 -83 0 net=2281
rlabel metal2 191 -83 191 -83 0 net=1366
rlabel metal2 222 -83 222 -83 0 net=716
rlabel metal2 233 -83 233 -83 0 net=859
rlabel metal2 282 -83 282 -83 0 net=1998
rlabel metal2 296 -83 296 -83 0 net=2653
rlabel metal2 317 -83 317 -83 0 net=2707
rlabel metal2 324 -83 324 -83 0 net=2046
rlabel metal2 121 -85 121 -85 0 net=1928
rlabel metal2 198 -85 198 -85 0 net=899
rlabel metal2 219 -85 219 -85 0 net=2121
rlabel metal2 117 -87 117 -87 0 net=118
rlabel metal2 128 -87 128 -87 0 net=1031
rlabel metal2 142 -87 142 -87 0 net=798
rlabel metal2 222 -87 222 -87 0 net=2293
rlabel metal2 226 -89 226 -89 0 net=2219
rlabel metal2 236 -91 236 -91 0 net=1504
rlabel metal2 240 -93 240 -93 0 net=2189
rlabel metal2 261 -95 261 -95 0 net=1371
rlabel metal2 86 -106 86 -106 0 net=559
rlabel metal2 107 -106 107 -106 0 net=2454
rlabel metal2 135 -106 135 -106 0 net=1032
rlabel metal2 149 -106 149 -106 0 net=2282
rlabel metal2 198 -106 198 -106 0 net=900
rlabel metal2 229 -106 229 -106 0 net=2190
rlabel metal2 282 -106 282 -106 0 net=2294
rlabel metal2 380 -106 380 -106 0 net=2991
rlabel metal2 114 -108 114 -108 0 net=2558
rlabel metal2 135 -108 135 -108 0 net=1589
rlabel metal2 198 -108 198 -108 0 net=2587
rlabel metal2 215 -108 215 -108 0 net=860
rlabel metal2 240 -108 240 -108 0 net=2299
rlabel metal2 240 -108 240 -108 0 net=2299
rlabel metal2 243 -108 243 -108 0 net=2586
rlabel metal2 103 -110 103 -110 0 net=450
rlabel metal2 156 -110 156 -110 0 net=1153
rlabel metal2 205 -110 205 -110 0 net=257
rlabel metal2 247 -110 247 -110 0 net=2122
rlabel metal2 289 -110 289 -110 0 net=2654
rlabel metal2 107 -112 107 -112 0 net=2897
rlabel metal2 163 -112 163 -112 0 net=801
rlabel metal2 177 -112 177 -112 0 net=666
rlabel metal2 268 -112 268 -112 0 net=2708
rlabel metal2 180 -114 180 -114 0 net=1325
rlabel metal2 208 -114 208 -114 0 net=1001
rlabel metal2 261 -114 261 -114 0 net=1373
rlabel metal2 303 -114 303 -114 0 net=2755
rlabel metal2 184 -116 184 -116 0 net=1285
rlabel metal2 212 -116 212 -116 0 net=752
rlabel metal2 310 -116 310 -116 0 net=2673
rlabel metal2 254 -118 254 -118 0 net=2221
rlabel metal2 226 -120 226 -120 0 net=2191
rlabel metal2 79 -131 79 -131 0 net=471
rlabel metal2 107 -131 107 -131 0 net=2898
rlabel metal2 156 -131 156 -131 0 net=1154
rlabel metal2 198 -131 198 -131 0 net=2588
rlabel metal2 198 -131 198 -131 0 net=2588
rlabel metal2 219 -131 219 -131 0 net=1003
rlabel metal2 257 -131 257 -131 0 net=2222
rlabel metal2 268 -131 268 -131 0 net=1374
rlabel metal2 296 -131 296 -131 0 net=2756
rlabel metal2 310 -131 310 -131 0 net=2674
rlabel metal2 380 -131 380 -131 0 net=2993
rlabel metal2 79 -133 79 -133 0 net=593
rlabel metal2 107 -133 107 -133 0 net=2921
rlabel metal2 131 -133 131 -133 0 net=319
rlabel metal2 159 -133 159 -133 0 net=491
rlabel metal2 226 -133 226 -133 0 net=2973
rlabel metal2 275 -133 275 -133 0 net=2035
rlabel metal2 114 -135 114 -135 0 net=2223
rlabel metal2 128 -135 128 -135 0 net=525
rlabel metal2 135 -135 135 -135 0 net=1590
rlabel metal2 163 -135 163 -135 0 net=802
rlabel metal2 184 -135 184 -135 0 net=1286
rlabel metal2 254 -135 254 -135 0 net=2193
rlabel metal2 299 -135 299 -135 0 net=2253
rlabel metal2 128 -137 128 -137 0 net=313
rlabel metal2 170 -137 170 -137 0 net=147
rlabel metal2 145 -139 145 -139 0 net=1867
rlabel metal2 173 -139 173 -139 0 net=2309
rlabel metal2 191 -139 191 -139 0 net=2229
rlabel metal2 121 -141 121 -141 0 net=2821
rlabel metal2 205 -141 205 -141 0 net=1327
rlabel metal2 152 -143 152 -143 0 net=800
rlabel metal2 205 -145 205 -145 0 net=2300
rlabel metal2 82 -156 82 -156 0 net=197
rlabel metal2 82 -156 82 -156 0 net=197
rlabel metal2 107 -156 107 -156 0 net=2922
rlabel metal2 156 -156 156 -156 0 net=1868
rlabel metal2 173 -156 173 -156 0 net=2310
rlabel metal2 187 -156 187 -156 0 net=2230
rlabel metal2 198 -156 198 -156 0 net=2975
rlabel metal2 233 -156 233 -156 0 net=1005
rlabel metal2 254 -156 254 -156 0 net=1971
rlabel metal2 317 -156 317 -156 0 net=680
rlabel metal2 359 -156 359 -156 0 net=2877
rlabel metal2 387 -156 387 -156 0 net=2995
rlabel metal2 408 -156 408 -156 0 net=2277
rlabel metal2 436 -156 436 -156 0 net=2503
rlabel metal2 114 -158 114 -158 0 net=2224
rlabel metal2 121 -158 121 -158 0 net=2822
rlabel metal2 152 -158 152 -158 0 net=473
rlabel metal2 212 -158 212 -158 0 net=1145
rlabel metal2 261 -158 261 -158 0 net=2194
rlabel metal2 296 -158 296 -158 0 net=1797
rlabel metal2 317 -158 317 -158 0 net=2255
rlabel metal2 331 -158 331 -158 0 net=2263
rlabel metal2 362 -158 362 -158 0 net=608
rlabel metal2 383 -158 383 -158 0 net=2581
rlabel metal2 124 -160 124 -160 0 net=436
rlabel metal2 163 -160 163 -160 0 net=1597
rlabel metal2 205 -160 205 -160 0 net=362
rlabel metal2 215 -160 215 -160 0 net=1328
rlabel metal2 226 -160 226 -160 0 net=2613
rlabel metal2 135 -162 135 -162 0 net=1113
rlabel metal2 170 -162 170 -162 0 net=1417
rlabel metal2 205 -162 205 -162 0 net=869
rlabel metal2 219 -162 219 -162 0 net=971
rlabel metal2 233 -162 233 -162 0 net=1685
rlabel metal2 320 -162 320 -162 0 net=2403
rlabel metal2 177 -164 177 -164 0 net=2019
rlabel metal2 261 -164 261 -164 0 net=2037
rlabel metal2 278 -164 278 -164 0 net=2521
rlabel metal2 240 -166 240 -166 0 net=1479
rlabel metal2 268 -168 268 -168 0 net=360
rlabel metal2 75 -179 75 -179 0 net=2007
rlabel metal2 86 -179 86 -179 0 net=438
rlabel metal2 131 -179 131 -179 0 net=234
rlabel metal2 131 -179 131 -179 0 net=234
rlabel metal2 135 -179 135 -179 0 net=1114
rlabel metal2 149 -179 149 -179 0 net=2977
rlabel metal2 229 -179 229 -179 0 net=1006
rlabel metal2 250 -179 250 -179 0 net=2979
rlabel metal2 369 -179 369 -179 0 net=2582
rlabel metal2 408 -179 408 -179 0 net=2823
rlabel metal2 408 -179 408 -179 0 net=2823
rlabel metal2 415 -179 415 -179 0 net=2278
rlabel metal2 432 -179 432 -179 0 net=2504
rlabel metal2 89 -181 89 -181 0 net=255
rlabel metal2 107 -181 107 -181 0 net=875
rlabel metal2 156 -181 156 -181 0 net=1893
rlabel metal2 163 -181 163 -181 0 net=1599
rlabel metal2 271 -181 271 -181 0 net=2522
rlabel metal2 338 -181 338 -181 0 net=2879
rlabel metal2 383 -181 383 -181 0 net=2996
rlabel metal2 401 -181 401 -181 0 net=1139
rlabel metal2 436 -181 436 -181 0 net=2363
rlabel metal2 121 -183 121 -183 0 net=1339
rlabel metal2 170 -183 170 -183 0 net=1418
rlabel metal2 233 -183 233 -183 0 net=2038
rlabel metal2 289 -183 289 -183 0 net=1687
rlabel metal2 289 -183 289 -183 0 net=1687
rlabel metal2 296 -183 296 -183 0 net=1798
rlabel metal2 317 -183 317 -183 0 net=2256
rlabel metal2 380 -183 380 -183 0 net=1995
rlabel metal2 170 -185 170 -185 0 net=973
rlabel metal2 229 -185 229 -185 0 net=1549
rlabel metal2 254 -185 254 -185 0 net=1146
rlabel metal2 303 -185 303 -185 0 net=1973
rlabel metal2 317 -185 317 -185 0 net=2265
rlabel metal2 345 -185 345 -185 0 net=2405
rlabel metal2 177 -187 177 -187 0 net=2020
rlabel metal2 219 -187 219 -187 0 net=1649
rlabel metal2 285 -187 285 -187 0 net=2211
rlabel metal2 177 -189 177 -189 0 net=1181
rlabel metal2 191 -189 191 -189 0 net=871
rlabel metal2 254 -189 254 -189 0 net=1115
rlabel metal2 285 -189 285 -189 0 net=2889
rlabel metal2 163 -191 163 -191 0 net=923
rlabel metal2 261 -191 261 -191 0 net=2129
rlabel metal2 331 -191 331 -191 0 net=2615
rlabel metal2 184 -193 184 -193 0 net=1481
rlabel metal2 296 -193 296 -193 0 net=1807
rlabel metal2 201 -195 201 -195 0 net=1099
rlabel metal2 72 -206 72 -206 0 net=37
rlabel metal2 100 -206 100 -206 0 net=1341
rlabel metal2 128 -206 128 -206 0 net=1173
rlabel metal2 261 -206 261 -206 0 net=2616
rlabel metal2 345 -206 345 -206 0 net=2213
rlabel metal2 394 -206 394 -206 0 net=1996
rlabel metal2 404 -206 404 -206 0 net=2824
rlabel metal2 415 -206 415 -206 0 net=1141
rlabel metal2 436 -206 436 -206 0 net=2364
rlabel metal2 79 -208 79 -208 0 net=2008
rlabel metal2 103 -208 103 -208 0 net=876
rlabel metal2 114 -208 114 -208 0 net=1155
rlabel metal2 114 -208 114 -208 0 net=1155
rlabel metal2 121 -208 121 -208 0 net=957
rlabel metal2 268 -208 268 -208 0 net=1601
rlabel metal2 306 -208 306 -208 0 net=2266
rlabel metal2 373 -208 373 -208 0 net=2406
rlabel metal2 79 -210 79 -210 0 net=1935
rlabel metal2 149 -210 149 -210 0 net=2978
rlabel metal2 236 -210 236 -210 0 net=2543
rlabel metal2 373 -210 373 -210 0 net=2691
rlabel metal2 86 -212 86 -212 0 net=1465
rlabel metal2 191 -212 191 -212 0 net=872
rlabel metal2 222 -212 222 -212 0 net=1100
rlabel metal2 257 -212 257 -212 0 net=1163
rlabel metal2 275 -212 275 -212 0 net=1651
rlabel metal2 359 -212 359 -212 0 net=2980
rlabel metal2 93 -214 93 -214 0 net=2175
rlabel metal2 156 -214 156 -214 0 net=1894
rlabel metal2 198 -214 198 -214 0 net=202
rlabel metal2 289 -214 289 -214 0 net=1689
rlabel metal2 289 -214 289 -214 0 net=1689
rlabel metal2 310 -214 310 -214 0 net=1975
rlabel metal2 107 -216 107 -216 0 net=955
rlabel metal2 229 -216 229 -216 0 net=2880
rlabel metal2 142 -218 142 -218 0 net=925
rlabel metal2 170 -218 170 -218 0 net=974
rlabel metal2 296 -218 296 -218 0 net=1809
rlabel metal2 324 -218 324 -218 0 net=2131
rlabel metal2 159 -220 159 -220 0 net=837
rlabel metal2 201 -220 201 -220 0 net=1263
rlabel metal2 324 -220 324 -220 0 net=2890
rlabel metal2 170 -222 170 -222 0 net=1183
rlabel metal2 205 -222 205 -222 0 net=1116
rlabel metal2 352 -222 352 -222 0 net=2009
rlabel metal2 131 -224 131 -224 0 net=677
rlabel metal2 184 -224 184 -224 0 net=1482
rlabel metal2 212 -224 212 -224 0 net=1769
rlabel metal2 212 -226 212 -226 0 net=1551
rlabel metal2 240 -226 240 -226 0 net=2059
rlabel metal2 233 -228 233 -228 0 net=1419
rlabel metal2 68 -239 68 -239 0 net=679
rlabel metal2 170 -239 170 -239 0 net=1184
rlabel metal2 229 -239 229 -239 0 net=1652
rlabel metal2 359 -239 359 -239 0 net=2061
rlabel metal2 450 -239 450 -239 0 net=2319
rlabel metal2 530 -239 530 -239 0 net=1631
rlabel metal2 86 -241 86 -241 0 net=1466
rlabel metal2 170 -241 170 -241 0 net=2239
rlabel metal2 240 -241 240 -241 0 net=1264
rlabel metal2 292 -241 292 -241 0 net=2047
rlabel metal2 366 -241 366 -241 0 net=86
rlabel metal2 79 -243 79 -243 0 net=1936
rlabel metal2 243 -243 243 -243 0 net=1602
rlabel metal2 331 -243 331 -243 0 net=1977
rlabel metal2 369 -243 369 -243 0 net=2214
rlabel metal2 394 -243 394 -243 0 net=2179
rlabel metal2 72 -245 72 -245 0 net=1565
rlabel metal2 93 -245 93 -245 0 net=2176
rlabel metal2 194 -245 194 -245 0 net=995
rlabel metal2 250 -245 250 -245 0 net=2544
rlabel metal2 418 -245 418 -245 0 net=1142
rlabel metal2 93 -247 93 -247 0 net=1553
rlabel metal2 254 -247 254 -247 0 net=178
rlabel metal2 271 -247 271 -247 0 net=2132
rlabel metal2 345 -247 345 -247 0 net=2011
rlabel metal2 373 -247 373 -247 0 net=2693
rlabel metal2 100 -249 100 -249 0 net=1342
rlabel metal2 138 -249 138 -249 0 net=373
rlabel metal2 208 -249 208 -249 0 net=2247
rlabel metal2 408 -249 408 -249 0 net=2575
rlabel metal2 107 -251 107 -251 0 net=956
rlabel metal2 177 -251 177 -251 0 net=839
rlabel metal2 212 -251 212 -251 0 net=1393
rlabel metal2 254 -251 254 -251 0 net=2347
rlabel metal2 107 -253 107 -253 0 net=1157
rlabel metal2 121 -253 121 -253 0 net=958
rlabel metal2 257 -253 257 -253 0 net=1701
rlabel metal2 338 -253 338 -253 0 net=2619
rlabel metal2 114 -255 114 -255 0 net=2905
rlabel metal2 180 -255 180 -255 0 net=2505
rlabel metal2 261 -255 261 -255 0 net=1783
rlabel metal2 121 -257 121 -257 0 net=401
rlabel metal2 198 -257 198 -257 0 net=1347
rlabel metal2 261 -257 261 -257 0 net=1165
rlabel metal2 275 -257 275 -257 0 net=1013
rlabel metal2 303 -257 303 -257 0 net=2925
rlabel metal2 128 -259 128 -259 0 net=1175
rlabel metal2 268 -259 268 -259 0 net=1897
rlabel metal2 131 -261 131 -261 0 net=590
rlabel metal2 296 -261 296 -261 0 net=1771
rlabel metal2 135 -263 135 -263 0 net=821
rlabel metal2 296 -263 296 -263 0 net=2655
rlabel metal2 142 -265 142 -265 0 net=926
rlabel metal2 310 -265 310 -265 0 net=1811
rlabel metal2 86 -267 86 -267 0 net=572
rlabel metal2 219 -267 219 -267 0 net=989
rlabel metal2 149 -269 149 -269 0 net=1420
rlabel metal2 282 -271 282 -271 0 net=1691
rlabel metal2 30 -282 30 -282 0 net=589
rlabel metal2 47 -282 47 -282 0 net=154
rlabel metal2 177 -282 177 -282 0 net=841
rlabel metal2 222 -282 222 -282 0 net=1166
rlabel metal2 268 -282 268 -282 0 net=2656
rlabel metal2 415 -282 415 -282 0 net=1457
rlabel metal2 453 -282 453 -282 0 net=2320
rlabel metal2 527 -282 527 -282 0 net=1633
rlabel metal2 30 -284 30 -284 0 net=304
rlabel metal2 51 -284 51 -284 0 net=406
rlabel metal2 58 -284 58 -284 0 net=1853
rlabel metal2 135 -284 135 -284 0 net=1177
rlabel metal2 184 -284 184 -284 0 net=691
rlabel metal2 243 -284 243 -284 0 net=632
rlabel metal2 68 -286 68 -286 0 net=1221
rlabel metal2 194 -286 194 -286 0 net=2180
rlabel metal2 401 -286 401 -286 0 net=2695
rlabel metal2 75 -288 75 -288 0 net=1566
rlabel metal2 82 -288 82 -288 0 net=582
rlabel metal2 205 -288 205 -288 0 net=1289
rlabel metal2 247 -288 247 -288 0 net=1395
rlabel metal2 292 -288 292 -288 0 net=1978
rlabel metal2 387 -288 387 -288 0 net=2927
rlabel metal2 86 -290 86 -290 0 net=2295
rlabel metal2 107 -290 107 -290 0 net=1158
rlabel metal2 149 -290 149 -290 0 net=2240
rlabel metal2 208 -290 208 -290 0 net=996
rlabel metal2 254 -290 254 -290 0 net=1812
rlabel metal2 380 -290 380 -290 0 net=2349
rlabel metal2 394 -290 394 -290 0 net=2577
rlabel metal2 93 -292 93 -292 0 net=1554
rlabel metal2 268 -292 268 -292 0 net=1015
rlabel metal2 282 -292 282 -292 0 net=1693
rlabel metal2 306 -292 306 -292 0 net=990
rlabel metal2 338 -292 338 -292 0 net=2621
rlabel metal2 408 -292 408 -292 0 net=2657
rlabel metal2 93 -294 93 -294 0 net=2907
rlabel metal2 121 -294 121 -294 0 net=987
rlabel metal2 156 -294 156 -294 0 net=823
rlabel metal2 226 -294 226 -294 0 net=2721
rlabel metal2 296 -294 296 -294 0 net=1772
rlabel metal2 100 -296 100 -296 0 net=1843
rlabel metal2 163 -296 163 -296 0 net=1785
rlabel metal2 352 -296 352 -296 0 net=1983
rlabel metal2 114 -298 114 -298 0 net=1349
rlabel metal2 226 -298 226 -298 0 net=117
rlabel metal2 299 -298 299 -298 0 net=2062
rlabel metal2 128 -300 128 -300 0 net=2127
rlabel metal2 310 -300 310 -300 0 net=1703
rlabel metal2 142 -302 142 -302 0 net=182
rlabel metal2 317 -302 317 -302 0 net=2013
rlabel metal2 170 -304 170 -304 0 net=2531
rlabel metal2 198 -306 198 -306 0 net=2507
rlabel metal2 331 -306 331 -306 0 net=1899
rlabel metal2 187 -308 187 -308 0 net=1451
rlabel metal2 331 -308 331 -308 0 net=2049
rlabel metal2 229 -310 229 -310 0 net=2323
rlabel metal2 359 -312 359 -312 0 net=2249
rlabel metal2 19 -323 19 -323 0 net=69
rlabel metal2 37 -323 37 -323 0 net=2909
rlabel metal2 96 -323 96 -323 0 net=396
rlabel metal2 194 -323 194 -323 0 net=2722
rlabel metal2 282 -323 282 -323 0 net=2622
rlabel metal2 373 -323 373 -323 0 net=1875
rlabel metal2 513 -323 513 -323 0 net=2675
rlabel metal2 523 -323 523 -323 0 net=1634
rlabel metal2 51 -325 51 -325 0 net=1895
rlabel metal2 219 -325 219 -325 0 net=1291
rlabel metal2 324 -325 324 -325 0 net=335
rlabel metal2 324 -325 324 -325 0 net=335
rlabel metal2 327 -325 327 -325 0 net=2050
rlabel metal2 408 -325 408 -325 0 net=2659
rlabel metal2 422 -325 422 -325 0 net=2929
rlabel metal2 58 -327 58 -327 0 net=1854
rlabel metal2 110 -327 110 -327 0 net=88
rlabel metal2 145 -327 145 -327 0 net=943
rlabel metal2 159 -327 159 -327 0 net=824
rlabel metal2 198 -327 198 -327 0 net=2508
rlabel metal2 247 -327 247 -327 0 net=2014
rlabel metal2 331 -327 331 -327 0 net=2325
rlabel metal2 390 -327 390 -327 0 net=2625
rlabel metal2 436 -327 436 -327 0 net=1458
rlabel metal2 58 -329 58 -329 0 net=2297
rlabel metal2 100 -329 100 -329 0 net=1844
rlabel metal2 177 -329 177 -329 0 net=1223
rlabel metal2 198 -329 198 -329 0 net=2367
rlabel metal2 387 -329 387 -329 0 net=2351
rlabel metal2 65 -331 65 -331 0 net=1179
rlabel metal2 149 -331 149 -331 0 net=1023
rlabel metal2 184 -331 184 -331 0 net=963
rlabel metal2 254 -331 254 -331 0 net=2063
rlabel metal2 401 -331 401 -331 0 net=2697
rlabel metal2 82 -333 82 -333 0 net=150
rlabel metal2 212 -333 212 -333 0 net=843
rlabel metal2 243 -333 243 -333 0 net=2532
rlabel metal2 72 -335 72 -335 0 net=1723
rlabel metal2 86 -335 86 -335 0 net=988
rlabel metal2 124 -335 124 -335 0 net=565
rlabel metal2 250 -335 250 -335 0 net=1694
rlabel metal2 100 -337 100 -337 0 net=2641
rlabel metal2 110 -337 110 -337 0 net=318
rlabel metal2 163 -337 163 -337 0 net=1786
rlabel metal2 261 -337 261 -337 0 net=1704
rlabel metal2 114 -339 114 -339 0 net=1351
rlabel metal2 264 -339 264 -339 0 net=2715
rlabel metal2 44 -341 44 -341 0 net=2033
rlabel metal2 117 -341 117 -341 0 net=1411
rlabel metal2 264 -341 264 -341 0 net=2427
rlabel metal2 128 -343 128 -343 0 net=2128
rlabel metal2 268 -343 268 -343 0 net=1016
rlabel metal2 285 -343 285 -343 0 net=1396
rlabel metal2 299 -343 299 -343 0 net=2923
rlabel metal2 131 -345 131 -345 0 net=649
rlabel metal2 194 -345 194 -345 0 net=2537
rlabel metal2 233 -347 233 -347 0 net=1452
rlabel metal2 289 -347 289 -347 0 net=1295
rlabel metal2 310 -347 310 -347 0 net=2251
rlabel metal2 170 -349 170 -349 0 net=1143
rlabel metal2 352 -349 352 -349 0 net=1985
rlabel metal2 345 -351 345 -351 0 net=1901
rlabel metal2 345 -353 345 -353 0 net=1979
rlabel metal2 394 -355 394 -355 0 net=2579
rlabel metal2 240 -357 240 -357 0 net=1505
rlabel metal2 240 -359 240 -359 0 net=2727
rlabel metal2 16 -370 16 -370 0 net=120
rlabel metal2 16 -370 16 -370 0 net=120
rlabel metal2 23 -370 23 -370 0 net=2643
rlabel metal2 121 -370 121 -370 0 net=1215
rlabel metal2 198 -370 198 -370 0 net=1251
rlabel metal2 275 -370 275 -370 0 net=2352
rlabel metal2 443 -370 443 -370 0 net=2429
rlabel metal2 30 -372 30 -372 0 net=98
rlabel metal2 135 -372 135 -372 0 net=699
rlabel metal2 219 -372 219 -372 0 net=845
rlabel metal2 219 -372 219 -372 0 net=845
rlabel metal2 226 -372 226 -372 0 net=1353
rlabel metal2 317 -372 317 -372 0 net=2064
rlabel metal2 387 -372 387 -372 0 net=2930
rlabel metal2 481 -372 481 -372 0 net=2963
rlabel metal2 513 -372 513 -372 0 net=2677
rlabel metal2 513 -372 513 -372 0 net=2677
rlabel metal2 30 -374 30 -374 0 net=2051
rlabel metal2 226 -374 226 -374 0 net=2252
rlabel metal2 331 -374 331 -374 0 net=2327
rlabel metal2 37 -376 37 -376 0 net=2910
rlabel metal2 128 -376 128 -376 0 net=1655
rlabel metal2 233 -376 233 -376 0 net=1144
rlabel metal2 282 -376 282 -376 0 net=2885
rlabel metal2 44 -378 44 -378 0 net=2034
rlabel metal2 138 -378 138 -378 0 net=1343
rlabel metal2 233 -378 233 -378 0 net=901
rlabel metal2 338 -378 338 -378 0 net=2539
rlabel metal2 390 -378 390 -378 0 net=2660
rlabel metal2 418 -378 418 -378 0 net=2743
rlabel metal2 44 -380 44 -380 0 net=712
rlabel metal2 149 -380 149 -380 0 net=1024
rlabel metal2 240 -380 240 -380 0 net=1292
rlabel metal2 310 -380 310 -380 0 net=2924
rlabel metal2 415 -380 415 -380 0 net=2481
rlabel metal2 450 -380 450 -380 0 net=2729
rlabel metal2 51 -382 51 -382 0 net=1896
rlabel metal2 243 -382 243 -382 0 net=1980
rlabel metal2 348 -382 348 -382 0 net=1813
rlabel metal2 394 -382 394 -382 0 net=1506
rlabel metal2 58 -384 58 -384 0 net=2298
rlabel metal2 254 -384 254 -384 0 net=545
rlabel metal2 296 -384 296 -384 0 net=1937
rlabel metal2 352 -384 352 -384 0 net=1903
rlabel metal2 408 -384 408 -384 0 net=2627
rlabel metal2 58 -386 58 -386 0 net=371
rlabel metal2 254 -386 254 -386 0 net=1297
rlabel metal2 352 -386 352 -386 0 net=1877
rlabel metal2 65 -388 65 -388 0 net=1180
rlabel metal2 250 -388 250 -388 0 net=2965
rlabel metal2 65 -390 65 -390 0 net=430
rlabel metal2 86 -390 86 -390 0 net=865
rlabel metal2 261 -390 261 -390 0 net=2368
rlabel metal2 408 -390 408 -390 0 net=2699
rlabel metal2 72 -392 72 -392 0 net=1724
rlabel metal2 110 -392 110 -392 0 net=105
rlabel metal2 261 -392 261 -392 0 net=2181
rlabel metal2 72 -394 72 -394 0 net=2245
rlabel metal2 268 -394 268 -394 0 net=2580
rlabel metal2 79 -396 79 -396 0 net=2161
rlabel metal2 131 -396 131 -396 0 net=1329
rlabel metal2 324 -396 324 -396 0 net=2383
rlabel metal2 37 -398 37 -398 0 net=672
rlabel metal2 114 -398 114 -398 0 net=1381
rlabel metal2 359 -398 359 -398 0 net=1987
rlabel metal2 89 -400 89 -400 0 net=1
rlabel metal2 156 -400 156 -400 0 net=944
rlabel metal2 212 -400 212 -400 0 net=1705
rlabel metal2 373 -400 373 -400 0 net=2717
rlabel metal2 93 -402 93 -402 0 net=965
rlabel metal2 229 -402 229 -402 0 net=2305
rlabel metal2 156 -404 156 -404 0 net=2807
rlabel metal2 177 -406 177 -406 0 net=1225
rlabel metal2 275 -406 275 -406 0 net=2401
rlabel metal2 177 -408 177 -408 0 net=2267
rlabel metal2 240 -408 240 -408 0 net=1781
rlabel metal2 317 -408 317 -408 0 net=1999
rlabel metal2 184 -410 184 -410 0 net=1413
rlabel metal2 16 -421 16 -421 0 net=2163
rlabel metal2 86 -421 86 -421 0 net=867
rlabel metal2 93 -421 93 -421 0 net=966
rlabel metal2 233 -421 233 -421 0 net=903
rlabel metal2 233 -421 233 -421 0 net=903
rlabel metal2 247 -421 247 -421 0 net=1226
rlabel metal2 268 -421 268 -421 0 net=831
rlabel metal2 289 -421 289 -421 0 net=1331
rlabel metal2 324 -421 324 -421 0 net=2964
rlabel metal2 513 -421 513 -421 0 net=2679
rlabel metal2 513 -421 513 -421 0 net=2679
rlabel metal2 520 -421 520 -421 0 net=2745
rlabel metal2 30 -423 30 -423 0 net=2052
rlabel metal2 159 -423 159 -423 0 net=2328
rlabel metal2 464 -423 464 -423 0 net=2887
rlabel metal2 30 -425 30 -425 0 net=487
rlabel metal2 114 -425 114 -425 0 net=1383
rlabel metal2 219 -425 219 -425 0 net=847
rlabel metal2 254 -425 254 -425 0 net=1299
rlabel metal2 327 -425 327 -425 0 net=2700
rlabel metal2 415 -425 415 -425 0 net=1293
rlabel metal2 44 -427 44 -427 0 net=1591
rlabel metal2 240 -427 240 -427 0 net=1782
rlabel metal2 261 -427 261 -427 0 net=2730
rlabel metal2 527 -427 527 -427 0 net=2431
rlabel metal2 2 -429 2 -429 0 net=2761
rlabel metal2 278 -429 278 -429 0 net=1938
rlabel metal2 331 -429 331 -429 0 net=1707
rlabel metal2 331 -429 331 -429 0 net=1707
rlabel metal2 338 -429 338 -429 0 net=1805
rlabel metal2 51 -431 51 -431 0 net=793
rlabel metal2 58 -431 58 -431 0 net=1217
rlabel metal2 128 -431 128 -431 0 net=1656
rlabel metal2 219 -431 219 -431 0 net=2681
rlabel metal2 37 -433 37 -433 0 net=1639
rlabel metal2 135 -433 135 -433 0 net=927
rlabel metal2 173 -433 173 -433 0 net=2339
rlabel metal2 471 -433 471 -433 0 net=2967
rlabel metal2 65 -435 65 -435 0 net=1253
rlabel metal2 226 -435 226 -435 0 net=2737
rlabel metal2 72 -437 72 -437 0 net=2246
rlabel metal2 341 -437 341 -437 0 net=1904
rlabel metal2 429 -437 429 -437 0 net=2719
rlabel metal2 72 -439 72 -439 0 net=1345
rlabel metal2 191 -439 191 -439 0 net=2402
rlabel metal2 285 -439 285 -439 0 net=2341
rlabel metal2 9 -441 9 -441 0 net=2217
rlabel metal2 177 -441 177 -441 0 net=2268
rlabel metal2 289 -441 289 -441 0 net=1355
rlabel metal2 348 -441 348 -441 0 net=2725
rlabel metal2 79 -443 79 -443 0 net=945
rlabel metal2 352 -443 352 -443 0 net=1879
rlabel metal2 436 -443 436 -443 0 net=2809
rlabel metal2 86 -445 86 -445 0 net=1415
rlabel metal2 198 -445 198 -445 0 net=286
rlabel metal2 296 -445 296 -445 0 net=1743
rlabel metal2 359 -445 359 -445 0 net=2307
rlabel metal2 96 -447 96 -447 0 net=1541
rlabel metal2 107 -447 107 -447 0 net=1101
rlabel metal2 177 -447 177 -447 0 net=1147
rlabel metal2 366 -447 366 -447 0 net=1815
rlabel metal2 436 -447 436 -447 0 net=2483
rlabel metal2 450 -447 450 -447 0 net=2629
rlabel metal2 450 -447 450 -447 0 net=2629
rlabel metal2 142 -449 142 -449 0 net=803
rlabel metal2 380 -449 380 -449 0 net=1989
rlabel metal2 443 -449 443 -449 0 net=2093
rlabel metal2 23 -451 23 -451 0 net=2645
rlabel metal2 205 -453 205 -453 0 net=879
rlabel metal2 373 -453 373 -453 0 net=2001
rlabel metal2 387 -453 387 -453 0 net=2541
rlabel metal2 229 -455 229 -455 0 net=1885
rlabel metal2 275 -457 275 -457 0 net=1749
rlabel metal2 394 -457 394 -457 0 net=2183
rlabel metal2 394 -459 394 -459 0 net=2385
rlabel metal2 397 -461 397 -461 0 net=1
rlabel metal2 9 -472 9 -472 0 net=2218
rlabel metal2 131 -472 131 -472 0 net=332
rlabel metal2 219 -472 219 -472 0 net=848
rlabel metal2 275 -472 275 -472 0 net=2342
rlabel metal2 513 -472 513 -472 0 net=2680
rlabel metal2 513 -472 513 -472 0 net=2680
rlabel metal2 555 -472 555 -472 0 net=2432
rlabel metal2 16 -474 16 -474 0 net=2164
rlabel metal2 152 -474 152 -474 0 net=1148
rlabel metal2 184 -474 184 -474 0 net=868
rlabel metal2 355 -474 355 -474 0 net=2810
rlabel metal2 558 -474 558 -474 0 net=2547
rlabel metal2 16 -476 16 -476 0 net=1483
rlabel metal2 100 -476 100 -476 0 net=1543
rlabel metal2 100 -476 100 -476 0 net=1543
rlabel metal2 107 -476 107 -476 0 net=1102
rlabel metal2 282 -476 282 -476 0 net=2853
rlabel metal2 23 -478 23 -478 0 net=614
rlabel metal2 159 -478 159 -478 0 net=2184
rlabel metal2 425 -478 425 -478 0 net=2726
rlabel metal2 30 -480 30 -480 0 net=1671
rlabel metal2 58 -480 58 -480 0 net=1218
rlabel metal2 107 -480 107 -480 0 net=905
rlabel metal2 240 -480 240 -480 0 net=1806
rlabel metal2 359 -480 359 -480 0 net=2888
rlabel metal2 37 -482 37 -482 0 net=1640
rlabel metal2 285 -482 285 -482 0 net=1880
rlabel metal2 464 -482 464 -482 0 net=2340
rlabel metal2 2 -484 2 -484 0 net=2762
rlabel metal2 299 -484 299 -484 0 net=2021
rlabel metal2 373 -484 373 -484 0 net=2308
rlabel metal2 541 -484 541 -484 0 net=2747
rlabel metal2 37 -486 37 -486 0 net=1359
rlabel metal2 142 -486 142 -486 0 net=805
rlabel metal2 163 -486 163 -486 0 net=2646
rlabel metal2 44 -488 44 -488 0 net=1592
rlabel metal2 135 -488 135 -488 0 net=929
rlabel metal2 170 -488 170 -488 0 net=2173
rlabel metal2 184 -488 184 -488 0 net=832
rlabel metal2 303 -488 303 -488 0 net=1332
rlabel metal2 331 -488 331 -488 0 net=1709
rlabel metal2 394 -488 394 -488 0 net=2387
rlabel metal2 51 -490 51 -490 0 net=1187
rlabel metal2 380 -490 380 -490 0 net=2003
rlabel metal2 408 -490 408 -490 0 net=1887
rlabel metal2 436 -490 436 -490 0 net=2485
rlabel metal2 72 -492 72 -492 0 net=1346
rlabel metal2 233 -492 233 -492 0 net=1583
rlabel metal2 380 -492 380 -492 0 net=1817
rlabel metal2 457 -492 457 -492 0 net=2683
rlabel metal2 44 -494 44 -494 0 net=1193
rlabel metal2 289 -494 289 -494 0 net=1357
rlabel metal2 310 -494 310 -494 0 net=2738
rlabel metal2 75 -496 75 -496 0 net=1257
rlabel metal2 124 -496 124 -496 0 net=637
rlabel metal2 222 -496 222 -496 0 net=1294
rlabel metal2 86 -498 86 -498 0 net=1416
rlabel metal2 289 -498 289 -498 0 net=1744
rlabel metal2 310 -498 310 -498 0 net=1300
rlabel metal2 331 -498 331 -498 0 net=2631
rlabel metal2 82 -500 82 -500 0 net=548
rlabel metal2 89 -500 89 -500 0 net=103
rlabel metal2 156 -500 156 -500 0 net=2073
rlabel metal2 429 -500 429 -500 0 net=1991
rlabel metal2 170 -502 170 -502 0 net=863
rlabel metal2 264 -502 264 -502 0 net=1389
rlabel metal2 296 -502 296 -502 0 net=2542
rlabel metal2 191 -504 191 -504 0 net=1081
rlabel metal2 320 -504 320 -504 0 net=2379
rlabel metal2 429 -504 429 -504 0 net=2095
rlabel metal2 478 -504 478 -504 0 net=2969
rlabel metal2 65 -506 65 -506 0 net=1254
rlabel metal2 282 -506 282 -506 0 net=2499
rlabel metal2 58 -508 58 -508 0 net=1471
rlabel metal2 201 -508 201 -508 0 net=1535
rlabel metal2 292 -508 292 -508 0 net=2827
rlabel metal2 201 -510 201 -510 0 net=799
rlabel metal2 212 -512 212 -512 0 net=1385
rlabel metal2 366 -512 366 -512 0 net=2811
rlabel metal2 205 -514 205 -514 0 net=881
rlabel metal2 226 -514 226 -514 0 net=2243
rlabel metal2 366 -514 366 -514 0 net=2720
rlabel metal2 79 -516 79 -516 0 net=947
rlabel metal2 387 -516 387 -516 0 net=1751
rlabel metal2 23 -518 23 -518 0 net=2491
rlabel metal2 390 -518 390 -518 0 net=2867
rlabel metal2 9 -529 9 -529 0 net=1485
rlabel metal2 23 -529 23 -529 0 net=2492
rlabel metal2 131 -529 131 -529 0 net=864
rlabel metal2 177 -529 177 -529 0 net=2174
rlabel metal2 198 -529 198 -529 0 net=883
rlabel metal2 215 -529 215 -529 0 net=574
rlabel metal2 226 -529 226 -529 0 net=2868
rlabel metal2 509 -529 509 -529 0 net=1467
rlabel metal2 562 -529 562 -529 0 net=2549
rlabel metal2 562 -529 562 -529 0 net=2549
rlabel metal2 16 -531 16 -531 0 net=705
rlabel metal2 268 -531 268 -531 0 net=1390
rlabel metal2 275 -531 275 -531 0 net=1201
rlabel metal2 373 -531 373 -531 0 net=299
rlabel metal2 541 -531 541 -531 0 net=2749
rlabel metal2 541 -531 541 -531 0 net=2749
rlabel metal2 30 -533 30 -533 0 net=1672
rlabel metal2 79 -533 79 -533 0 net=1545
rlabel metal2 107 -533 107 -533 0 net=907
rlabel metal2 205 -533 205 -533 0 net=948
rlabel metal2 296 -533 296 -533 0 net=1387
rlabel metal2 331 -533 331 -533 0 net=2632
rlabel metal2 373 -533 373 -533 0 net=1753
rlabel metal2 30 -535 30 -535 0 net=2461
rlabel metal2 93 -535 93 -535 0 net=1259
rlabel metal2 93 -535 93 -535 0 net=1259
rlabel metal2 103 -535 103 -535 0 net=167
rlabel metal2 219 -535 219 -535 0 net=181
rlabel metal2 37 -537 37 -537 0 net=1360
rlabel metal2 247 -537 247 -537 0 net=1537
rlabel metal2 247 -537 247 -537 0 net=1537
rlabel metal2 254 -537 254 -537 0 net=2244
rlabel metal2 306 -537 306 -537 0 net=1888
rlabel metal2 478 -537 478 -537 0 net=2501
rlabel metal2 40 -539 40 -539 0 net=472
rlabel metal2 107 -539 107 -539 0 net=930
rlabel metal2 254 -539 254 -539 0 net=1911
rlabel metal2 464 -539 464 -539 0 net=2487
rlabel metal2 485 -539 485 -539 0 net=2388
rlabel metal2 44 -541 44 -541 0 net=1194
rlabel metal2 156 -541 156 -541 0 net=511
rlabel metal2 289 -541 289 -541 0 net=1317
rlabel metal2 380 -541 380 -541 0 net=1819
rlabel metal2 380 -541 380 -541 0 net=1819
rlabel metal2 492 -541 492 -541 0 net=2971
rlabel metal2 51 -543 51 -543 0 net=1188
rlabel metal2 208 -543 208 -543 0 net=2957
rlabel metal2 51 -545 51 -545 0 net=2015
rlabel metal2 114 -545 114 -545 0 net=420
rlabel metal2 268 -545 268 -545 0 net=1358
rlabel metal2 313 -545 313 -545 0 net=2079
rlabel metal2 492 -545 492 -545 0 net=2415
rlabel metal2 58 -547 58 -547 0 net=1472
rlabel metal2 124 -547 124 -547 0 net=555
rlabel metal2 149 -547 149 -547 0 net=807
rlabel metal2 163 -547 163 -547 0 net=1409
rlabel metal2 282 -547 282 -547 0 net=2854
rlabel metal2 58 -549 58 -549 0 net=1923
rlabel metal2 117 -549 117 -549 0 net=131
rlabel metal2 313 -549 313 -549 0 net=2828
rlabel metal2 121 -551 121 -551 0 net=1397
rlabel metal2 317 -551 317 -551 0 net=1429
rlabel metal2 331 -551 331 -551 0 net=2091
rlabel metal2 345 -551 345 -551 0 net=1993
rlabel metal2 128 -553 128 -553 0 net=1507
rlabel metal2 229 -553 229 -553 0 net=1679
rlabel metal2 348 -553 348 -553 0 net=2812
rlabel metal2 443 -553 443 -553 0 net=2685
rlabel metal2 135 -555 135 -555 0 net=1585
rlabel metal2 240 -555 240 -555 0 net=2953
rlabel metal2 149 -557 149 -557 0 net=1083
rlabel metal2 240 -557 240 -557 0 net=1055
rlabel metal2 352 -557 352 -557 0 net=1869
rlabel metal2 159 -559 159 -559 0 net=967
rlabel metal2 338 -559 338 -559 0 net=1711
rlabel metal2 359 -559 359 -559 0 net=2023
rlabel metal2 415 -559 415 -559 0 net=2075
rlabel metal2 142 -561 142 -561 0 net=1831
rlabel metal2 362 -561 362 -561 0 net=2563
rlabel metal2 236 -563 236 -563 0 net=160
rlabel metal2 394 -563 394 -563 0 net=2005
rlabel metal2 429 -563 429 -563 0 net=2097
rlabel metal2 394 -565 394 -565 0 net=2381
rlabel metal2 429 -565 429 -565 0 net=2177
rlabel metal2 264 -567 264 -567 0 net=1957
rlabel metal2 9 -578 9 -578 0 net=1486
rlabel metal2 93 -578 93 -578 0 net=1261
rlabel metal2 93 -578 93 -578 0 net=1261
rlabel metal2 121 -578 121 -578 0 net=1399
rlabel metal2 289 -578 289 -578 0 net=1319
rlabel metal2 338 -578 338 -578 0 net=2382
rlabel metal2 408 -578 408 -578 0 net=2025
rlabel metal2 408 -578 408 -578 0 net=2025
rlabel metal2 429 -578 429 -578 0 net=2077
rlabel metal2 464 -578 464 -578 0 net=2564
rlabel metal2 530 -578 530 -578 0 net=2750
rlabel metal2 555 -578 555 -578 0 net=1469
rlabel metal2 555 -578 555 -578 0 net=1469
rlabel metal2 562 -578 562 -578 0 net=2550
rlabel metal2 562 -578 562 -578 0 net=2550
rlabel metal2 9 -580 9 -580 0 net=2989
rlabel metal2 121 -580 121 -580 0 net=1423
rlabel metal2 135 -580 135 -580 0 net=1586
rlabel metal2 222 -580 222 -580 0 net=2092
rlabel metal2 338 -580 338 -580 0 net=1994
rlabel metal2 359 -580 359 -580 0 net=2006
rlabel metal2 432 -580 432 -580 0 net=2972
rlabel metal2 534 -580 534 -580 0 net=2502
rlabel metal2 23 -582 23 -582 0 net=683
rlabel metal2 72 -582 72 -582 0 net=1924
rlabel metal2 86 -582 86 -582 0 net=703
rlabel metal2 233 -582 233 -582 0 net=1538
rlabel metal2 254 -582 254 -582 0 net=1203
rlabel metal2 324 -582 324 -582 0 net=1681
rlabel metal2 341 -582 341 -582 0 net=1659
rlabel metal2 352 -582 352 -582 0 net=1713
rlabel metal2 366 -582 366 -582 0 net=1821
rlabel metal2 436 -582 436 -582 0 net=2954
rlabel metal2 520 -582 520 -582 0 net=2155
rlabel metal2 23 -584 23 -584 0 net=2709
rlabel metal2 135 -584 135 -584 0 net=496
rlabel metal2 380 -584 380 -584 0 net=1913
rlabel metal2 436 -584 436 -584 0 net=1929
rlabel metal2 523 -584 523 -584 0 net=1883
rlabel metal2 30 -586 30 -586 0 net=2462
rlabel metal2 138 -586 138 -586 0 net=1410
rlabel metal2 170 -586 170 -586 0 net=1011
rlabel metal2 191 -586 191 -586 0 net=968
rlabel metal2 236 -586 236 -586 0 net=678
rlabel metal2 30 -588 30 -588 0 net=2017
rlabel metal2 54 -588 54 -588 0 net=83
rlabel metal2 72 -588 72 -588 0 net=1509
rlabel metal2 145 -588 145 -588 0 net=808
rlabel metal2 191 -588 191 -588 0 net=1103
rlabel metal2 352 -588 352 -588 0 net=1459
rlabel metal2 16 -590 16 -590 0 net=2713
rlabel metal2 58 -590 58 -590 0 net=2551
rlabel metal2 79 -590 79 -590 0 net=1546
rlabel metal2 142 -590 142 -590 0 net=1833
rlabel metal2 198 -590 198 -590 0 net=884
rlabel metal2 240 -590 240 -590 0 net=2789
rlabel metal2 443 -590 443 -590 0 net=2687
rlabel metal2 471 -590 471 -590 0 net=1871
rlabel metal2 37 -592 37 -592 0 net=1881
rlabel metal2 79 -592 79 -592 0 net=1051
rlabel metal2 149 -592 149 -592 0 net=1084
rlabel metal2 198 -592 198 -592 0 net=1333
rlabel metal2 275 -592 275 -592 0 net=1431
rlabel metal2 387 -592 387 -592 0 net=2081
rlabel metal2 443 -592 443 -592 0 net=2099
rlabel metal2 481 -592 481 -592 0 net=2958
rlabel metal2 103 -594 103 -594 0 net=1907
rlabel metal2 205 -594 205 -594 0 net=1388
rlabel metal2 373 -594 373 -594 0 net=1755
rlabel metal2 485 -594 485 -594 0 net=2178
rlabel metal2 142 -596 142 -596 0 net=1823
rlabel metal2 401 -596 401 -596 0 net=1959
rlabel metal2 485 -596 485 -596 0 net=2417
rlabel metal2 499 -596 499 -596 0 net=2509
rlabel metal2 149 -598 149 -598 0 net=1235
rlabel metal2 450 -598 450 -598 0 net=2489
rlabel metal2 205 -600 205 -600 0 net=983
rlabel metal2 208 -602 208 -602 0 net=1379
rlabel metal2 247 -602 247 -602 0 net=1057
rlabel metal2 268 -602 268 -602 0 net=2849
rlabel metal2 177 -604 177 -604 0 net=909
rlabel metal2 289 -604 289 -604 0 net=2301
rlabel metal2 219 -606 219 -606 0 net=440
rlabel metal2 306 -606 306 -606 0 net=2101
rlabel metal2 229 -608 229 -608 0 net=2115
rlabel metal2 261 -610 261 -610 0 net=1301
rlabel metal2 9 -621 9 -621 0 net=2990
rlabel metal2 72 -621 72 -621 0 net=1510
rlabel metal2 142 -621 142 -621 0 net=492
rlabel metal2 233 -621 233 -621 0 net=1380
rlabel metal2 296 -621 296 -621 0 net=1914
rlabel metal2 394 -621 394 -621 0 net=1930
rlabel metal2 443 -621 443 -621 0 net=2100
rlabel metal2 499 -621 499 -621 0 net=2511
rlabel metal2 513 -621 513 -621 0 net=2411
rlabel metal2 16 -623 16 -623 0 net=2714
rlabel metal2 65 -623 65 -623 0 net=2571
rlabel metal2 121 -623 121 -623 0 net=1425
rlabel metal2 121 -623 121 -623 0 net=1425
rlabel metal2 163 -623 163 -623 0 net=1908
rlabel metal2 184 -623 184 -623 0 net=1335
rlabel metal2 219 -623 219 -623 0 net=1058
rlabel metal2 261 -623 261 -623 0 net=1302
rlabel metal2 422 -623 422 -623 0 net=2303
rlabel metal2 450 -623 450 -623 0 net=2490
rlabel metal2 516 -623 516 -623 0 net=1884
rlabel metal2 544 -623 544 -623 0 net=1470
rlabel metal2 23 -625 23 -625 0 net=2710
rlabel metal2 93 -625 93 -625 0 net=1262
rlabel metal2 103 -625 103 -625 0 net=474
rlabel metal2 310 -625 310 -625 0 net=1714
rlabel metal2 401 -625 401 -625 0 net=2103
rlabel metal2 520 -625 520 -625 0 net=2157
rlabel metal2 555 -625 555 -625 0 net=2435
rlabel metal2 30 -627 30 -627 0 net=2018
rlabel metal2 51 -627 51 -627 0 net=2553
rlabel metal2 72 -627 72 -627 0 net=1137
rlabel metal2 96 -627 96 -627 0 net=754
rlabel metal2 222 -627 222 -627 0 net=1245
rlabel metal2 275 -627 275 -627 0 net=1433
rlabel metal2 317 -627 317 -627 0 net=2117
rlabel metal2 527 -627 527 -627 0 net=1873
rlabel metal2 37 -629 37 -629 0 net=1882
rlabel metal2 107 -629 107 -629 0 net=1053
rlabel metal2 149 -629 149 -629 0 net=1237
rlabel metal2 226 -629 226 -629 0 net=1321
rlabel metal2 327 -629 327 -629 0 net=2078
rlabel metal2 44 -631 44 -631 0 net=2565
rlabel metal2 334 -631 334 -631 0 net=2082
rlabel metal2 397 -631 397 -631 0 net=2159
rlabel metal2 86 -633 86 -633 0 net=877
rlabel metal2 114 -633 114 -633 0 net=817
rlabel metal2 233 -633 233 -633 0 net=2545
rlabel metal2 275 -633 275 -633 0 net=1107
rlabel metal2 352 -633 352 -633 0 net=1756
rlabel metal2 75 -635 75 -635 0 net=1511
rlabel metal2 114 -635 114 -635 0 net=258
rlabel metal2 282 -635 282 -635 0 net=1401
rlabel metal2 282 -635 282 -635 0 net=1401
rlabel metal2 296 -635 296 -635 0 net=1825
rlabel metal2 380 -635 380 -635 0 net=1981
rlabel metal2 408 -635 408 -635 0 net=2027
rlabel metal2 422 -635 422 -635 0 net=1961
rlabel metal2 131 -637 131 -637 0 net=1837
rlabel metal2 366 -637 366 -637 0 net=1822
rlabel metal2 149 -639 149 -639 0 net=1835
rlabel metal2 163 -639 163 -639 0 net=1219
rlabel metal2 240 -639 240 -639 0 net=2790
rlabel metal2 324 -639 324 -639 0 net=2203
rlabel metal2 128 -641 128 -641 0 net=1287
rlabel metal2 170 -641 170 -641 0 net=1012
rlabel metal2 191 -641 191 -641 0 net=1105
rlabel metal2 324 -641 324 -641 0 net=1557
rlabel metal2 40 -643 40 -643 0 net=748
rlabel metal2 180 -643 180 -643 0 net=1039
rlabel metal2 205 -643 205 -643 0 net=985
rlabel metal2 254 -643 254 -643 0 net=1205
rlabel metal2 331 -643 331 -643 0 net=1683
rlabel metal2 401 -643 401 -643 0 net=2053
rlabel metal2 254 -645 254 -645 0 net=1461
rlabel metal2 331 -647 331 -647 0 net=1801
rlabel metal2 481 -647 481 -647 0 net=2647
rlabel metal2 338 -649 338 -649 0 net=2329
rlabel metal2 341 -651 341 -651 0 net=2455
rlabel metal2 268 -653 268 -653 0 net=910
rlabel metal2 345 -653 345 -653 0 net=1660
rlabel metal2 355 -653 355 -653 0 net=2850
rlabel metal2 345 -655 345 -655 0 net=2688
rlabel metal2 485 -655 485 -655 0 net=2419
rlabel metal2 464 -657 464 -657 0 net=2783
rlabel metal2 16 -668 16 -668 0 net=2573
rlabel metal2 107 -668 107 -668 0 net=878
rlabel metal2 114 -668 114 -668 0 net=1054
rlabel metal2 142 -668 142 -668 0 net=1677
rlabel metal2 142 -668 142 -668 0 net=1677
rlabel metal2 156 -668 156 -668 0 net=1288
rlabel metal2 296 -668 296 -668 0 net=1827
rlabel metal2 320 -668 320 -668 0 net=2160
rlabel metal2 471 -668 471 -668 0 net=2859
rlabel metal2 628 -668 628 -668 0 net=2423
rlabel metal2 23 -670 23 -670 0 net=2603
rlabel metal2 156 -670 156 -670 0 net=1239
rlabel metal2 205 -670 205 -670 0 net=986
rlabel metal2 240 -670 240 -670 0 net=1207
rlabel metal2 303 -670 303 -670 0 net=1106
rlabel metal2 471 -670 471 -670 0 net=2331
rlabel metal2 485 -670 485 -670 0 net=1653
rlabel metal2 499 -670 499 -670 0 net=2457
rlabel metal2 516 -670 516 -670 0 net=2158
rlabel metal2 527 -670 527 -670 0 net=2589
rlabel metal2 30 -672 30 -672 0 net=2333
rlabel metal2 44 -672 44 -672 0 net=2566
rlabel metal2 163 -672 163 -672 0 net=1220
rlabel metal2 170 -672 170 -672 0 net=2546
rlabel metal2 247 -672 247 -672 0 net=1097
rlabel metal2 345 -672 345 -672 0 net=2843
rlabel metal2 583 -672 583 -672 0 net=2413
rlabel metal2 44 -674 44 -674 0 net=2555
rlabel metal2 58 -674 58 -674 0 net=1138
rlabel metal2 93 -674 93 -674 0 net=1073
rlabel metal2 114 -674 114 -674 0 net=1121
rlabel metal2 170 -674 170 -674 0 net=1323
rlabel metal2 247 -674 247 -674 0 net=937
rlabel metal2 348 -674 348 -674 0 net=1684
rlabel metal2 376 -674 376 -674 0 net=2028
rlabel metal2 478 -674 478 -674 0 net=2421
rlabel metal2 499 -674 499 -674 0 net=2437
rlabel metal2 593 -674 593 -674 0 net=2185
rlabel metal2 51 -676 51 -676 0 net=1065
rlabel metal2 352 -676 352 -676 0 net=1367
rlabel metal2 380 -676 380 -676 0 net=1982
rlabel metal2 415 -676 415 -676 0 net=2205
rlabel metal2 506 -676 506 -676 0 net=2513
rlabel metal2 530 -676 530 -676 0 net=1874
rlabel metal2 548 -676 548 -676 0 net=2649
rlabel metal2 65 -678 65 -678 0 net=1512
rlabel metal2 191 -678 191 -678 0 net=1041
rlabel metal2 250 -678 250 -678 0 net=2784
rlabel metal2 72 -680 72 -680 0 net=939
rlabel metal2 86 -680 86 -680 0 net=1427
rlabel metal2 201 -680 201 -680 0 net=2315
rlabel metal2 212 -680 212 -680 0 net=1109
rlabel metal2 296 -680 296 -680 0 net=2637
rlabel metal2 121 -682 121 -682 0 net=1603
rlabel metal2 219 -682 219 -682 0 net=819
rlabel metal2 324 -682 324 -682 0 net=1559
rlabel metal2 380 -682 380 -682 0 net=1061
rlabel metal2 177 -684 177 -684 0 net=861
rlabel metal2 219 -684 219 -684 0 net=289
rlabel metal2 254 -684 254 -684 0 net=1463
rlabel metal2 331 -684 331 -684 0 net=2935
rlabel metal2 184 -686 184 -686 0 net=1337
rlabel metal2 261 -686 261 -686 0 net=1247
rlabel metal2 338 -686 338 -686 0 net=2493
rlabel metal2 135 -688 135 -688 0 net=969
rlabel metal2 268 -688 268 -688 0 net=2515
rlabel metal2 149 -690 149 -690 0 net=1836
rlabel metal2 194 -690 194 -690 0 net=1035
rlabel metal2 310 -690 310 -690 0 net=1434
rlabel metal2 359 -690 359 -690 0 net=1839
rlabel metal2 443 -690 443 -690 0 net=2105
rlabel metal2 128 -692 128 -692 0 net=2527
rlabel metal2 233 -692 233 -692 0 net=1227
rlabel metal2 366 -692 366 -692 0 net=2055
rlabel metal2 443 -692 443 -692 0 net=2369
rlabel metal2 282 -694 282 -694 0 net=1403
rlabel metal2 387 -694 387 -694 0 net=1803
rlabel metal2 387 -696 387 -696 0 net=2304
rlabel metal2 450 -696 450 -696 0 net=2119
rlabel metal2 345 -698 345 -698 0 net=1915
rlabel metal2 450 -698 450 -698 0 net=2447
rlabel metal2 394 -700 394 -700 0 net=2791
rlabel metal2 397 -702 397 -702 0 net=1962
rlabel metal2 408 -704 408 -704 0 net=1313
rlabel metal2 422 -706 422 -706 0 net=2947
rlabel metal2 16 -717 16 -717 0 net=2574
rlabel metal2 86 -717 86 -717 0 net=1428
rlabel metal2 142 -717 142 -717 0 net=1678
rlabel metal2 152 -717 152 -717 0 net=337
rlabel metal2 194 -717 194 -717 0 net=2316
rlabel metal2 219 -717 219 -717 0 net=1338
rlabel metal2 261 -717 261 -717 0 net=970
rlabel metal2 348 -717 348 -717 0 net=2206
rlabel metal2 422 -717 422 -717 0 net=2133
rlabel metal2 495 -717 495 -717 0 net=2936
rlabel metal2 541 -717 541 -717 0 net=2948
rlabel metal2 23 -719 23 -719 0 net=2604
rlabel metal2 79 -719 79 -719 0 net=940
rlabel metal2 156 -719 156 -719 0 net=1241
rlabel metal2 268 -719 268 -719 0 net=1036
rlabel metal2 334 -719 334 -719 0 net=2332
rlabel metal2 474 -719 474 -719 0 net=1669
rlabel metal2 562 -719 562 -719 0 net=2650
rlabel metal2 611 -719 611 -719 0 net=2186
rlabel metal2 33 -721 33 -721 0 net=2334
rlabel metal2 44 -721 44 -721 0 net=2556
rlabel metal2 79 -721 79 -721 0 net=1123
rlabel metal2 156 -721 156 -721 0 net=931
rlabel metal2 296 -721 296 -721 0 net=1464
rlabel metal2 338 -721 338 -721 0 net=2120
rlabel metal2 485 -721 485 -721 0 net=1654
rlabel metal2 485 -721 485 -721 0 net=1654
rlabel metal2 499 -721 499 -721 0 net=2438
rlabel metal2 593 -721 593 -721 0 net=2414
rlabel metal2 44 -723 44 -723 0 net=1605
rlabel metal2 163 -723 163 -723 0 net=862
rlabel metal2 194 -723 194 -723 0 net=1098
rlabel metal2 310 -723 310 -723 0 net=2494
rlabel metal2 527 -723 527 -723 0 net=2590
rlabel metal2 569 -723 569 -723 0 net=1062
rlabel metal2 51 -725 51 -725 0 net=1066
rlabel metal2 268 -725 268 -725 0 net=1249
rlabel metal2 310 -725 310 -725 0 net=1405
rlabel metal2 366 -725 366 -725 0 net=2056
rlabel metal2 597 -725 597 -725 0 net=2424
rlabel metal2 51 -727 51 -727 0 net=2529
rlabel metal2 163 -727 163 -727 0 net=1085
rlabel metal2 233 -727 233 -727 0 net=1229
rlabel metal2 233 -727 233 -727 0 net=1229
rlabel metal2 240 -727 240 -727 0 net=1208
rlabel metal2 317 -727 317 -727 0 net=1829
rlabel metal2 352 -727 352 -727 0 net=1369
rlabel metal2 65 -729 65 -729 0 net=1191
rlabel metal2 86 -729 86 -729 0 net=1075
rlabel metal2 103 -729 103 -729 0 net=2106
rlabel metal2 464 -729 464 -729 0 net=2639
rlabel metal2 58 -731 58 -731 0 net=1391
rlabel metal2 114 -731 114 -731 0 net=895
rlabel metal2 170 -731 170 -731 0 net=1324
rlabel metal2 205 -731 205 -731 0 net=2871
rlabel metal2 317 -731 317 -731 0 net=2389
rlabel metal2 352 -731 352 -731 0 net=1657
rlabel metal2 366 -731 366 -731 0 net=2459
rlabel metal2 555 -731 555 -731 0 net=2861
rlabel metal2 72 -733 72 -733 0 net=1059
rlabel metal2 121 -733 121 -733 0 net=1641
rlabel metal2 226 -733 226 -733 0 net=1043
rlabel metal2 247 -733 247 -733 0 net=938
rlabel metal2 397 -733 397 -733 0 net=2514
rlabel metal2 93 -735 93 -735 0 net=1513
rlabel metal2 170 -735 170 -735 0 net=1111
rlabel metal2 250 -735 250 -735 0 net=573
rlabel metal2 408 -735 408 -735 0 net=1315
rlabel metal2 107 -737 107 -737 0 net=2911
rlabel metal2 222 -737 222 -737 0 net=2231
rlabel metal2 408 -737 408 -737 0 net=2371
rlabel metal2 450 -737 450 -737 0 net=2449
rlabel metal2 506 -737 506 -737 0 net=2845
rlabel metal2 177 -739 177 -739 0 net=1611
rlabel metal2 222 -739 222 -739 0 net=653
rlabel metal2 373 -739 373 -739 0 net=1561
rlabel metal2 184 -741 184 -741 0 net=833
rlabel metal2 254 -741 254 -741 0 net=187
rlabel metal2 380 -741 380 -741 0 net=2422
rlabel metal2 142 -743 142 -743 0 net=1625
rlabel metal2 275 -743 275 -743 0 net=820
rlabel metal2 282 -743 282 -743 0 net=1840
rlabel metal2 415 -743 415 -743 0 net=2731
rlabel metal2 478 -743 478 -743 0 net=2517
rlabel metal2 292 -745 292 -745 0 net=2767
rlabel metal2 425 -745 425 -745 0 net=1804
rlabel metal2 334 -747 334 -747 0 net=2949
rlabel metal2 338 -749 338 -749 0 net=2931
rlabel metal2 380 -751 380 -751 0 net=1917
rlabel metal2 429 -753 429 -753 0 net=2793
rlabel metal2 394 -755 394 -755 0 net=2407
rlabel metal2 394 -757 394 -757 0 net=2399
rlabel metal2 26 -768 26 -768 0 net=369
rlabel metal2 40 -768 40 -768 0 net=291
rlabel metal2 152 -768 152 -768 0 net=759
rlabel metal2 387 -768 387 -768 0 net=2233
rlabel metal2 397 -768 397 -768 0 net=2450
rlabel metal2 471 -768 471 -768 0 net=1316
rlabel metal2 534 -768 534 -768 0 net=1670
rlabel metal2 30 -770 30 -770 0 net=1863
rlabel metal2 44 -770 44 -770 0 net=1606
rlabel metal2 128 -770 128 -770 0 net=896
rlabel metal2 170 -770 170 -770 0 net=1112
rlabel metal2 212 -770 212 -770 0 net=1250
rlabel metal2 275 -770 275 -770 0 net=2400
rlabel metal2 446 -770 446 -770 0 net=2518
rlabel metal2 492 -770 492 -770 0 net=1563
rlabel metal2 44 -772 44 -772 0 net=1515
rlabel metal2 128 -772 128 -772 0 net=1661
rlabel metal2 212 -772 212 -772 0 net=1406
rlabel metal2 324 -772 324 -772 0 net=1830
rlabel metal2 352 -772 352 -772 0 net=1658
rlabel metal2 513 -772 513 -772 0 net=2951
rlabel metal2 51 -774 51 -774 0 net=2530
rlabel metal2 156 -774 156 -774 0 net=932
rlabel metal2 219 -774 219 -774 0 net=1242
rlabel metal2 285 -774 285 -774 0 net=2390
rlabel metal2 334 -774 334 -774 0 net=2519
rlabel metal2 499 -774 499 -774 0 net=2795
rlabel metal2 520 -774 520 -774 0 net=2863
rlabel metal2 51 -776 51 -776 0 net=1643
rlabel metal2 135 -776 135 -776 0 net=1007
rlabel metal2 135 -776 135 -776 0 net=1007
rlabel metal2 156 -776 156 -776 0 net=1273
rlabel metal2 222 -776 222 -776 0 net=1735
rlabel metal2 292 -776 292 -776 0 net=52
rlabel metal2 401 -776 401 -776 0 net=2769
rlabel metal2 58 -778 58 -778 0 net=1392
rlabel metal2 163 -778 163 -778 0 net=1086
rlabel metal2 338 -778 338 -778 0 net=2917
rlabel metal2 492 -778 492 -778 0 net=2771
rlabel metal2 58 -780 58 -780 0 net=1192
rlabel metal2 72 -780 72 -780 0 net=1060
rlabel metal2 163 -780 163 -780 0 net=1277
rlabel metal2 303 -780 303 -780 0 net=1119
rlabel metal2 429 -780 429 -780 0 net=2409
rlabel metal2 65 -782 65 -782 0 net=2855
rlabel metal2 359 -782 359 -782 0 net=2640
rlabel metal2 72 -784 72 -784 0 net=194
rlabel metal2 170 -784 170 -784 0 net=933
rlabel metal2 261 -784 261 -784 0 net=2134
rlabel metal2 443 -784 443 -784 0 net=2669
rlabel metal2 86 -786 86 -786 0 net=1076
rlabel metal2 121 -786 121 -786 0 net=2353
rlabel metal2 464 -786 464 -786 0 net=2847
rlabel metal2 86 -788 86 -788 0 net=1049
rlabel metal2 226 -788 226 -788 0 net=1067
rlabel metal2 303 -788 303 -788 0 net=1211
rlabel metal2 359 -788 359 -788 0 net=1919
rlabel metal2 404 -788 404 -788 0 net=2343
rlabel metal2 93 -790 93 -790 0 net=1185
rlabel metal2 306 -790 306 -790 0 net=2701
rlabel metal2 177 -792 177 -792 0 net=1613
rlabel metal2 103 -794 103 -794 0 net=1265
rlabel metal2 184 -794 184 -794 0 net=1627
rlabel metal2 229 -794 229 -794 0 net=2460
rlabel metal2 205 -796 205 -796 0 net=1093
rlabel metal2 233 -796 233 -796 0 net=1231
rlabel metal2 313 -796 313 -796 0 net=2197
rlabel metal2 215 -798 215 -798 0 net=885
rlabel metal2 236 -798 236 -798 0 net=702
rlabel metal2 366 -798 366 -798 0 net=2373
rlabel metal2 240 -800 240 -800 0 net=1045
rlabel metal2 240 -800 240 -800 0 net=1045
rlabel metal2 247 -800 247 -800 0 net=2872
rlabel metal2 317 -800 317 -800 0 net=2623
rlabel metal2 247 -802 247 -802 0 net=2289
rlabel metal2 254 -804 254 -804 0 net=1370
rlabel metal2 296 -806 296 -806 0 net=1727
rlabel metal2 450 -806 450 -806 0 net=2933
rlabel metal2 376 -808 376 -808 0 net=2143
rlabel metal2 415 -808 415 -808 0 net=2733
rlabel metal2 107 -810 107 -810 0 net=2913
rlabel metal2 79 -812 79 -812 0 net=1124
rlabel metal2 79 -814 79 -814 0 net=835
rlabel metal2 26 -825 26 -825 0 net=93
rlabel metal2 44 -825 44 -825 0 net=1516
rlabel metal2 240 -825 240 -825 0 net=1046
rlabel metal2 254 -825 254 -825 0 net=949
rlabel metal2 306 -825 306 -825 0 net=2520
rlabel metal2 30 -827 30 -827 0 net=1864
rlabel metal2 44 -827 44 -827 0 net=285
rlabel metal2 75 -827 75 -827 0 net=563
rlabel metal2 114 -827 114 -827 0 net=2031
rlabel metal2 145 -827 145 -827 0 net=640
rlabel metal2 320 -827 320 -827 0 net=1120
rlabel metal2 401 -827 401 -827 0 net=2848
rlabel metal2 467 -827 467 -827 0 net=2934
rlabel metal2 51 -829 51 -829 0 net=1644
rlabel metal2 173 -829 173 -829 0 net=121
rlabel metal2 201 -829 201 -829 0 net=110
rlabel metal2 450 -829 450 -829 0 net=2735
rlabel metal2 37 -831 37 -831 0 net=825
rlabel metal2 58 -831 58 -831 0 net=2445
rlabel metal2 187 -831 187 -831 0 net=586
rlabel metal2 313 -831 313 -831 0 net=2952
rlabel metal2 79 -833 79 -833 0 net=836
rlabel metal2 212 -833 212 -833 0 net=887
rlabel metal2 240 -833 240 -833 0 net=1069
rlabel metal2 296 -833 296 -833 0 net=2595
rlabel metal2 457 -833 457 -833 0 net=2813
rlabel metal2 79 -835 79 -835 0 net=935
rlabel metal2 177 -835 177 -835 0 net=1267
rlabel metal2 261 -835 261 -835 0 net=1614
rlabel metal2 331 -835 331 -835 0 net=2374
rlabel metal2 373 -835 373 -835 0 net=2796
rlabel metal2 86 -837 86 -837 0 net=1050
rlabel metal2 205 -837 205 -837 0 net=1095
rlabel metal2 310 -837 310 -837 0 net=1963
rlabel metal2 324 -837 324 -837 0 net=1921
rlabel metal2 366 -837 366 -837 0 net=2345
rlabel metal2 86 -839 86 -839 0 net=1009
rlabel metal2 149 -839 149 -839 0 net=57
rlabel metal2 100 -841 100 -841 0 net=1629
rlabel metal2 257 -841 257 -841 0 net=1305
rlabel metal2 107 -843 107 -843 0 net=1275
rlabel metal2 226 -843 226 -843 0 net=1279
rlabel metal2 313 -843 313 -843 0 net=2624
rlabel metal2 117 -845 117 -845 0 net=2311
rlabel metal2 121 -847 121 -847 0 net=1212
rlabel metal2 348 -847 348 -847 0 net=2770
rlabel metal2 124 -849 124 -849 0 net=1662
rlabel metal2 149 -849 149 -849 0 net=1487
rlabel metal2 338 -849 338 -849 0 net=2919
rlabel metal2 93 -851 93 -851 0 net=1186
rlabel metal2 156 -851 156 -851 0 net=1847
rlabel metal2 289 -851 289 -851 0 net=1737
rlabel metal2 355 -851 355 -851 0 net=2410
rlabel metal2 65 -853 65 -853 0 net=2857
rlabel metal2 163 -853 163 -853 0 net=1169
rlabel metal2 247 -853 247 -853 0 net=1435
rlabel metal2 359 -853 359 -853 0 net=2145
rlabel metal2 520 -853 520 -853 0 net=2865
rlabel metal2 65 -855 65 -855 0 net=2215
rlabel metal2 268 -855 268 -855 0 net=1233
rlabel metal2 373 -855 373 -855 0 net=2198
rlabel metal2 268 -857 268 -857 0 net=1729
rlabel metal2 387 -857 387 -857 0 net=1931
rlabel metal2 492 -857 492 -857 0 net=2773
rlabel metal2 376 -859 376 -859 0 net=1564
rlabel metal2 348 -861 348 -861 0 net=1577
rlabel metal2 401 -863 401 -863 0 net=2355
rlabel metal2 408 -865 408 -865 0 net=2291
rlabel metal2 436 -865 436 -865 0 net=2703
rlabel metal2 352 -867 352 -867 0 net=2763
rlabel metal2 415 -869 415 -869 0 net=2915
rlabel metal2 394 -871 394 -871 0 net=2235
rlabel metal2 422 -871 422 -871 0 net=2671
rlabel metal2 152 -873 152 -873 0 net=2335
rlabel metal2 233 -875 233 -875 0 net=1949
rlabel metal2 233 -877 233 -877 0 net=1841
rlabel metal2 9 -888 9 -888 0 net=2711
rlabel metal2 142 -888 142 -888 0 net=2032
rlabel metal2 159 -888 159 -888 0 net=2916
rlabel metal2 520 -888 520 -888 0 net=2866
rlabel metal2 16 -890 16 -890 0 net=1063
rlabel metal2 240 -890 240 -890 0 net=1070
rlabel metal2 268 -890 268 -890 0 net=1730
rlabel metal2 348 -890 348 -890 0 net=2736
rlabel metal2 520 -890 520 -890 0 net=2609
rlabel metal2 23 -892 23 -892 0 net=2601
rlabel metal2 58 -892 58 -892 0 net=2446
rlabel metal2 355 -892 355 -892 0 net=2704
rlabel metal2 457 -892 457 -892 0 net=2815
rlabel metal2 44 -894 44 -894 0 net=826
rlabel metal2 58 -894 58 -894 0 net=1731
rlabel metal2 79 -894 79 -894 0 net=936
rlabel metal2 177 -894 177 -894 0 net=889
rlabel metal2 240 -894 240 -894 0 net=1243
rlabel metal2 359 -894 359 -894 0 net=2147
rlabel metal2 373 -894 373 -894 0 net=2069
rlabel metal2 373 -894 373 -894 0 net=2069
rlabel metal2 380 -894 380 -894 0 net=1306
rlabel metal2 37 -896 37 -896 0 net=2425
rlabel metal2 233 -896 233 -896 0 net=1842
rlabel metal2 383 -896 383 -896 0 net=2739
rlabel metal2 51 -898 51 -898 0 net=1195
rlabel metal2 313 -898 313 -898 0 net=2292
rlabel metal2 422 -898 422 -898 0 net=2672
rlabel metal2 478 -898 478 -898 0 net=2765
rlabel metal2 65 -900 65 -900 0 net=2216
rlabel metal2 142 -900 142 -900 0 net=951
rlabel metal2 282 -900 282 -900 0 net=1922
rlabel metal2 331 -900 331 -900 0 net=2920
rlabel metal2 65 -902 65 -902 0 net=2201
rlabel metal2 194 -902 194 -902 0 net=1096
rlabel metal2 282 -902 282 -902 0 net=1939
rlabel metal2 352 -902 352 -902 0 net=2851
rlabel metal2 86 -904 86 -904 0 net=1010
rlabel metal2 296 -904 296 -904 0 net=1779
rlabel metal2 436 -904 436 -904 0 net=2337
rlabel metal2 478 -904 478 -904 0 net=2775
rlabel metal2 93 -906 93 -906 0 net=2858
rlabel metal2 201 -906 201 -906 0 net=490
rlabel metal2 317 -906 317 -906 0 net=1965
rlabel metal2 359 -906 359 -906 0 net=2357
rlabel metal2 506 -906 506 -906 0 net=1579
rlabel metal2 93 -908 93 -908 0 net=1715
rlabel metal2 149 -908 149 -908 0 net=1489
rlabel metal2 317 -908 317 -908 0 net=1739
rlabel metal2 394 -908 394 -908 0 net=1950
rlabel metal2 100 -910 100 -910 0 net=1630
rlabel metal2 205 -910 205 -910 0 net=1234
rlabel metal2 397 -910 397 -910 0 net=2689
rlabel metal2 107 -912 107 -912 0 net=1276
rlabel metal2 401 -912 401 -912 0 net=2237
rlabel metal2 107 -914 107 -914 0 net=1437
rlabel metal2 275 -914 275 -914 0 net=1849
rlabel metal2 415 -914 415 -914 0 net=2313
rlabel metal2 114 -916 114 -916 0 net=1619
rlabel metal2 152 -916 152 -916 0 net=1645
rlabel metal2 201 -916 201 -916 0 net=1635
rlabel metal2 306 -916 306 -916 0 net=2346
rlabel metal2 429 -916 429 -916 0 net=2597
rlabel metal2 121 -918 121 -918 0 net=1171
rlabel metal2 208 -918 208 -918 0 net=1311
rlabel metal2 387 -918 387 -918 0 net=1933
rlabel metal2 124 -920 124 -920 0 net=615
rlabel metal2 184 -920 184 -920 0 net=1531
rlabel metal2 226 -920 226 -920 0 net=1281
rlabel metal2 128 -922 128 -922 0 net=849
rlabel metal2 219 -922 219 -922 0 net=1269
rlabel metal2 159 -924 159 -924 0 net=59
rlabel metal2 166 -926 166 -926 0 net=1763
rlabel metal2 205 -928 205 -928 0 net=2273
rlabel metal2 219 -930 219 -930 0 net=2495
rlabel metal2 226 -932 226 -932 0 net=2467
rlabel metal2 2 -943 2 -943 0 net=2441
rlabel metal2 201 -943 201 -943 0 net=1780
rlabel metal2 443 -943 443 -943 0 net=2852
rlabel metal2 16 -945 16 -945 0 net=1064
rlabel metal2 107 -945 107 -945 0 net=1439
rlabel metal2 114 -945 114 -945 0 net=1620
rlabel metal2 142 -945 142 -945 0 net=952
rlabel metal2 212 -945 212 -945 0 net=1244
rlabel metal2 257 -945 257 -945 0 net=1312
rlabel metal2 299 -945 299 -945 0 net=2314
rlabel metal2 429 -945 429 -945 0 net=2599
rlabel metal2 464 -945 464 -945 0 net=2766
rlabel metal2 9 -947 9 -947 0 net=2712
rlabel metal2 222 -947 222 -947 0 net=531
rlabel metal2 268 -947 268 -947 0 net=1491
rlabel metal2 310 -947 310 -947 0 net=2275
rlabel metal2 467 -947 467 -947 0 net=2816
rlabel metal2 23 -949 23 -949 0 net=2602
rlabel metal2 37 -949 37 -949 0 net=2426
rlabel metal2 254 -949 254 -949 0 net=1765
rlabel metal2 317 -949 317 -949 0 net=1741
rlabel metal2 317 -949 317 -949 0 net=1741
rlabel metal2 324 -949 324 -949 0 net=2238
rlabel metal2 492 -949 492 -949 0 net=2741
rlabel metal2 9 -951 9 -951 0 net=2287
rlabel metal2 44 -951 44 -951 0 net=1533
rlabel metal2 187 -951 187 -951 0 net=911
rlabel metal2 268 -951 268 -951 0 net=1271
rlabel metal2 296 -951 296 -951 0 net=1761
rlabel metal2 327 -951 327 -951 0 net=2559
rlabel metal2 16 -953 16 -953 0 net=311
rlabel metal2 51 -953 51 -953 0 net=1196
rlabel metal2 198 -953 198 -953 0 net=2365
rlabel metal2 51 -955 51 -955 0 net=1733
rlabel metal2 65 -955 65 -955 0 net=2202
rlabel metal2 247 -955 247 -955 0 net=1637
rlabel metal2 338 -955 338 -955 0 net=1851
rlabel metal2 394 -955 394 -955 0 net=2776
rlabel metal2 65 -957 65 -957 0 net=809
rlabel metal2 306 -957 306 -957 0 net=2803
rlabel metal2 478 -957 478 -957 0 net=1581
rlabel metal2 75 -959 75 -959 0 net=7
rlabel metal2 107 -959 107 -959 0 net=1647
rlabel metal2 177 -959 177 -959 0 net=891
rlabel metal2 331 -959 331 -959 0 net=479
rlabel metal2 345 -959 345 -959 0 net=1967
rlabel metal2 506 -959 506 -959 0 net=2611
rlabel metal2 86 -961 86 -961 0 net=661
rlabel metal2 163 -961 163 -961 0 net=1940
rlabel metal2 289 -961 289 -961 0 net=2873
rlabel metal2 352 -961 352 -961 0 net=1934
rlabel metal2 86 -963 86 -963 0 net=1453
rlabel metal2 373 -963 373 -963 0 net=2071
rlabel metal2 93 -965 93 -965 0 net=1716
rlabel metal2 177 -965 177 -965 0 net=488
rlabel metal2 373 -965 373 -965 0 net=2149
rlabel metal2 96 -967 96 -967 0 net=2690
rlabel metal2 114 -969 114 -969 0 net=999
rlabel metal2 194 -969 194 -969 0 net=1695
rlabel metal2 264 -969 264 -969 0 net=2338
rlabel metal2 457 -969 457 -969 0 net=2468
rlabel metal2 121 -971 121 -971 0 net=1172
rlabel metal2 226 -971 226 -971 0 net=2817
rlabel metal2 128 -973 128 -973 0 net=850
rlabel metal2 233 -973 233 -973 0 net=1283
rlabel metal2 359 -973 359 -973 0 net=2359
rlabel metal2 82 -975 82 -975 0 net=452
rlabel metal2 355 -975 355 -975 0 net=1757
rlabel metal2 366 -975 366 -975 0 net=2497
rlabel metal2 135 -977 135 -977 0 net=1077
rlabel metal2 149 -977 149 -977 0 net=1149
rlabel metal2 334 -977 334 -977 0 net=2751
rlabel metal2 159 -979 159 -979 0 net=348
rlabel metal2 334 -979 334 -979 0 net=2723
rlabel metal2 121 -981 121 -981 0 net=2463
rlabel metal2 9 -992 9 -992 0 net=2288
rlabel metal2 44 -992 44 -992 0 net=1534
rlabel metal2 229 -992 229 -992 0 net=1017
rlabel metal2 247 -992 247 -992 0 net=1697
rlabel metal2 247 -992 247 -992 0 net=1697
rlabel metal2 278 -992 278 -992 0 net=1852
rlabel metal2 418 -992 418 -992 0 net=2498
rlabel metal2 439 -992 439 -992 0 net=1582
rlabel metal2 488 -992 488 -992 0 net=2612
rlabel metal2 16 -994 16 -994 0 net=180
rlabel metal2 16 -994 16 -994 0 net=180
rlabel metal2 23 -994 23 -994 0 net=1361
rlabel metal2 37 -994 37 -994 0 net=2881
rlabel metal2 51 -994 51 -994 0 net=1734
rlabel metal2 65 -994 65 -994 0 net=810
rlabel metal2 107 -994 107 -994 0 net=1648
rlabel metal2 187 -994 187 -994 0 net=1638
rlabel metal2 289 -994 289 -994 0 net=1742
rlabel metal2 341 -994 341 -994 0 net=2600
rlabel metal2 446 -994 446 -994 0 net=1521
rlabel metal2 40 -996 40 -996 0 net=275
rlabel metal2 107 -996 107 -996 0 net=2869
rlabel metal2 205 -996 205 -996 0 net=893
rlabel metal2 205 -996 205 -996 0 net=893
rlabel metal2 215 -996 215 -996 0 net=18
rlabel metal2 233 -996 233 -996 0 net=2875
rlabel metal2 352 -996 352 -996 0 net=2724
rlabel metal2 467 -996 467 -996 0 net=1447
rlabel metal2 474 -996 474 -996 0 net=2742
rlabel metal2 58 -998 58 -998 0 net=991
rlabel metal2 79 -998 79 -998 0 net=1000
rlabel metal2 121 -998 121 -998 0 net=2465
rlabel metal2 121 -998 121 -998 0 net=2465
rlabel metal2 131 -998 131 -998 0 net=1762
rlabel metal2 327 -998 327 -998 0 net=2085
rlabel metal2 359 -998 359 -998 0 net=1759
rlabel metal2 359 -998 359 -998 0 net=1759
rlabel metal2 380 -998 380 -998 0 net=2361
rlabel metal2 415 -998 415 -998 0 net=2561
rlabel metal2 82 -1000 82 -1000 0 net=2818
rlabel metal2 2 -1002 2 -1002 0 net=2442
rlabel metal2 86 -1002 86 -1002 0 net=1454
rlabel metal2 285 -1002 285 -1002 0 net=1441
rlabel metal2 303 -1002 303 -1002 0 net=1493
rlabel metal2 334 -1002 334 -1002 0 net=1745
rlabel metal2 366 -1002 366 -1002 0 net=2753
rlabel metal2 422 -1002 422 -1002 0 net=2072
rlabel metal2 86 -1004 86 -1004 0 net=1125
rlabel metal2 142 -1004 142 -1004 0 net=1079
rlabel metal2 142 -1004 142 -1004 0 net=1079
rlabel metal2 149 -1004 149 -1004 0 net=1150
rlabel metal2 163 -1004 163 -1004 0 net=704
rlabel metal2 170 -1004 170 -1004 0 net=1440
rlabel metal2 310 -1004 310 -1004 0 net=1767
rlabel metal2 96 -1006 96 -1006 0 net=1375
rlabel metal2 149 -1006 149 -1006 0 net=2366
rlabel metal2 156 -1008 156 -1008 0 net=1477
rlabel metal2 191 -1008 191 -1008 0 net=1284
rlabel metal2 415 -1008 415 -1008 0 net=2391
rlabel metal2 191 -1010 191 -1010 0 net=913
rlabel metal2 222 -1010 222 -1010 0 net=2107
rlabel metal2 212 -1012 212 -1012 0 net=1272
rlabel metal2 128 -1014 128 -1014 0 net=1889
rlabel metal2 128 -1016 128 -1016 0 net=2433
rlabel metal2 222 -1016 222 -1016 0 net=2276
rlabel metal2 177 -1018 177 -1018 0 net=1407
rlabel metal2 394 -1018 394 -1018 0 net=2805
rlabel metal2 198 -1020 198 -1020 0 net=1593
rlabel metal2 373 -1020 373 -1020 0 net=2151
rlabel metal2 254 -1022 254 -1022 0 net=2825
rlabel metal2 373 -1022 373 -1022 0 net=1951
rlabel metal2 254 -1024 254 -1024 0 net=1555
rlabel metal2 338 -1026 338 -1026 0 net=1968
rlabel metal2 292 -1028 292 -1028 0 net=2663
rlabel metal2 23 -1039 23 -1039 0 net=1362
rlabel metal2 51 -1039 51 -1039 0 net=993
rlabel metal2 72 -1039 72 -1039 0 net=2283
rlabel metal2 86 -1039 86 -1039 0 net=1126
rlabel metal2 117 -1039 117 -1039 0 net=2466
rlabel metal2 128 -1039 128 -1039 0 net=2434
rlabel metal2 159 -1039 159 -1039 0 net=1773
rlabel metal2 299 -1039 299 -1039 0 net=1760
rlabel metal2 408 -1039 408 -1039 0 net=2806
rlabel metal2 443 -1039 443 -1039 0 net=2562
rlabel metal2 460 -1039 460 -1039 0 net=609
rlabel metal2 488 -1039 488 -1039 0 net=953
rlabel metal2 30 -1041 30 -1041 0 net=2883
rlabel metal2 68 -1041 68 -1041 0 net=2199
rlabel metal2 100 -1041 100 -1041 0 net=1377
rlabel metal2 121 -1041 121 -1041 0 net=1197
rlabel metal2 149 -1041 149 -1041 0 net=1478
rlabel metal2 177 -1041 177 -1041 0 net=1408
rlabel metal2 205 -1041 205 -1041 0 net=894
rlabel metal2 233 -1041 233 -1041 0 net=2876
rlabel metal2 285 -1041 285 -1041 0 net=1494
rlabel metal2 324 -1041 324 -1041 0 net=2754
rlabel metal2 401 -1041 401 -1041 0 net=2665
rlabel metal2 429 -1041 429 -1041 0 net=2393
rlabel metal2 464 -1041 464 -1041 0 net=1449
rlabel metal2 37 -1043 37 -1043 0 net=981
rlabel metal2 110 -1043 110 -1043 0 net=514
rlabel metal2 163 -1043 163 -1043 0 net=1556
rlabel metal2 261 -1043 261 -1043 0 net=2826
rlabel metal2 331 -1043 331 -1043 0 net=2067
rlabel metal2 345 -1043 345 -1043 0 net=2087
rlabel metal2 394 -1043 394 -1043 0 net=2153
rlabel metal2 408 -1043 408 -1043 0 net=2135
rlabel metal2 86 -1045 86 -1045 0 net=1859
rlabel metal2 128 -1045 128 -1045 0 net=811
rlabel metal2 135 -1047 135 -1047 0 net=1080
rlabel metal2 177 -1047 177 -1047 0 net=1047
rlabel metal2 222 -1047 222 -1047 0 net=99
rlabel metal2 303 -1047 303 -1047 0 net=1768
rlabel metal2 418 -1047 418 -1047 0 net=750
rlabel metal2 478 -1047 478 -1047 0 net=1523
rlabel metal2 107 -1049 107 -1049 0 net=2870
rlabel metal2 184 -1049 184 -1049 0 net=915
rlabel metal2 198 -1049 198 -1049 0 net=1595
rlabel metal2 215 -1049 215 -1049 0 net=2591
rlabel metal2 96 -1051 96 -1051 0 net=437
rlabel metal2 198 -1051 198 -1051 0 net=2165
rlabel metal2 135 -1053 135 -1053 0 net=975
rlabel metal2 233 -1053 233 -1053 0 net=1473
rlabel metal2 268 -1053 268 -1053 0 net=1891
rlabel metal2 338 -1053 338 -1053 0 net=2321
rlabel metal2 240 -1055 240 -1055 0 net=1018
rlabel metal2 303 -1055 303 -1055 0 net=2535
rlabel metal2 240 -1057 240 -1057 0 net=853
rlabel metal2 341 -1057 341 -1057 0 net=2891
rlabel metal2 247 -1059 247 -1059 0 net=1699
rlabel metal2 268 -1059 268 -1059 0 net=2039
rlabel metal2 149 -1061 149 -1061 0 net=1167
rlabel metal2 278 -1061 278 -1061 0 net=1499
rlabel metal2 348 -1061 348 -1061 0 net=2362
rlabel metal2 310 -1063 310 -1063 0 net=2109
rlabel metal2 289 -1065 289 -1065 0 net=1443
rlabel metal2 373 -1065 373 -1065 0 net=1953
rlabel metal2 229 -1067 229 -1067 0 net=2785
rlabel metal2 289 -1069 289 -1069 0 net=1746
rlabel metal2 352 -1071 352 -1071 0 net=1607
rlabel metal2 345 -1073 345 -1073 0 net=2829
rlabel metal2 30 -1084 30 -1084 0 net=2884
rlabel metal2 47 -1084 47 -1084 0 net=526
rlabel metal2 79 -1084 79 -1084 0 net=2200
rlabel metal2 79 -1084 79 -1084 0 net=2200
rlabel metal2 86 -1084 86 -1084 0 net=1860
rlabel metal2 96 -1084 96 -1084 0 net=1048
rlabel metal2 184 -1084 184 -1084 0 net=917
rlabel metal2 184 -1084 184 -1084 0 net=917
rlabel metal2 191 -1084 191 -1084 0 net=468
rlabel metal2 212 -1084 212 -1084 0 net=1892
rlabel metal2 338 -1084 338 -1084 0 net=2154
rlabel metal2 432 -1084 432 -1084 0 net=1450
rlabel metal2 471 -1084 471 -1084 0 net=68
rlabel metal2 481 -1084 481 -1084 0 net=1524
rlabel metal2 495 -1084 495 -1084 0 net=954
rlabel metal2 37 -1086 37 -1086 0 net=982
rlabel metal2 212 -1086 212 -1086 0 net=411
rlabel metal2 345 -1086 345 -1086 0 net=2593
rlabel metal2 401 -1086 401 -1086 0 net=2893
rlabel metal2 51 -1088 51 -1088 0 net=994
rlabel metal2 100 -1088 100 -1088 0 net=1378
rlabel metal2 170 -1088 170 -1088 0 net=1168
rlabel metal2 271 -1088 271 -1088 0 net=1444
rlabel metal2 338 -1088 338 -1088 0 net=2787
rlabel metal2 436 -1088 436 -1088 0 net=2831
rlabel metal2 436 -1088 436 -1088 0 net=2831
rlabel metal2 450 -1088 450 -1088 0 net=2395
rlabel metal2 58 -1090 58 -1090 0 net=53
rlabel metal2 114 -1090 114 -1090 0 net=977
rlabel metal2 149 -1090 149 -1090 0 net=854
rlabel metal2 271 -1090 271 -1090 0 net=2068
rlabel metal2 348 -1090 348 -1090 0 net=1954
rlabel metal2 65 -1092 65 -1092 0 net=2285
rlabel metal2 100 -1092 100 -1092 0 net=1199
rlabel metal2 124 -1092 124 -1092 0 net=1793
rlabel metal2 149 -1092 149 -1092 0 net=2113
rlabel metal2 229 -1092 229 -1092 0 net=1500
rlabel metal2 352 -1092 352 -1092 0 net=1609
rlabel metal2 72 -1094 72 -1094 0 net=1209
rlabel metal2 128 -1094 128 -1094 0 net=813
rlabel metal2 128 -1094 128 -1094 0 net=813
rlabel metal2 163 -1094 163 -1094 0 net=1567
rlabel metal2 173 -1094 173 -1094 0 net=571
rlabel metal2 240 -1094 240 -1094 0 net=829
rlabel metal2 268 -1094 268 -1094 0 net=2225
rlabel metal2 366 -1094 366 -1094 0 net=2041
rlabel metal2 380 -1094 380 -1094 0 net=2167
rlabel metal2 82 -1096 82 -1096 0 net=611
rlabel metal2 156 -1096 156 -1096 0 net=709
rlabel metal2 177 -1096 177 -1096 0 net=1455
rlabel metal2 226 -1096 226 -1096 0 net=126
rlabel metal2 366 -1096 366 -1096 0 net=2536
rlabel metal2 156 -1098 156 -1098 0 net=1799
rlabel metal2 289 -1098 289 -1098 0 net=2089
rlabel metal2 369 -1098 369 -1098 0 net=2322
rlabel metal2 194 -1100 194 -1100 0 net=599
rlabel metal2 236 -1100 236 -1100 0 net=1700
rlabel metal2 275 -1100 275 -1100 0 net=1775
rlabel metal2 303 -1100 303 -1100 0 net=1029
rlabel metal2 303 -1100 303 -1100 0 net=1029
rlabel metal2 310 -1100 310 -1100 0 net=2757
rlabel metal2 359 -1100 359 -1100 0 net=2111
rlabel metal2 422 -1100 422 -1100 0 net=2667
rlabel metal2 107 -1102 107 -1102 0 net=106
rlabel metal2 233 -1102 233 -1102 0 net=1717
rlabel metal2 261 -1102 261 -1102 0 net=1475
rlabel metal2 373 -1102 373 -1102 0 net=2137
rlabel metal2 145 -1104 145 -1104 0 net=1159
rlabel metal2 205 -1106 205 -1106 0 net=1596
rlabel metal2 394 -1106 394 -1106 0 net=2983
rlabel metal2 47 -1117 47 -1117 0 net=827
rlabel metal2 72 -1117 72 -1117 0 net=1210
rlabel metal2 93 -1117 93 -1117 0 net=613
rlabel metal2 93 -1117 93 -1117 0 net=613
rlabel metal2 100 -1117 100 -1117 0 net=1200
rlabel metal2 149 -1117 149 -1117 0 net=2114
rlabel metal2 212 -1117 212 -1117 0 net=454
rlabel metal2 229 -1117 229 -1117 0 net=84
rlabel metal2 334 -1117 334 -1117 0 net=1610
rlabel metal2 394 -1117 394 -1117 0 net=2895
rlabel metal2 408 -1117 408 -1117 0 net=2668
rlabel metal2 65 -1119 65 -1119 0 net=2286
rlabel metal2 100 -1119 100 -1119 0 net=1517
rlabel metal2 285 -1119 285 -1119 0 net=1476
rlabel metal2 306 -1119 306 -1119 0 net=747
rlabel metal2 338 -1119 338 -1119 0 net=2788
rlabel metal2 408 -1119 408 -1119 0 net=2985
rlabel metal2 422 -1119 422 -1119 0 net=2042
rlabel metal2 65 -1121 65 -1121 0 net=2195
rlabel metal2 110 -1121 110 -1121 0 net=2479
rlabel metal2 149 -1121 149 -1121 0 net=2269
rlabel metal2 233 -1121 233 -1121 0 net=394
rlabel metal2 261 -1121 261 -1121 0 net=1161
rlabel metal2 261 -1121 261 -1121 0 net=1161
rlabel metal2 275 -1121 275 -1121 0 net=1777
rlabel metal2 317 -1121 317 -1121 0 net=2227
rlabel metal2 352 -1121 352 -1121 0 net=2112
rlabel metal2 366 -1121 366 -1121 0 net=2375
rlabel metal2 415 -1121 415 -1121 0 net=1497
rlabel metal2 450 -1121 450 -1121 0 net=2397
rlabel metal2 114 -1123 114 -1123 0 net=978
rlabel metal2 170 -1123 170 -1123 0 net=1569
rlabel metal2 289 -1123 289 -1123 0 net=2090
rlabel metal2 317 -1123 317 -1123 0 net=2169
rlabel metal2 387 -1123 387 -1123 0 net=266
rlabel metal2 422 -1123 422 -1123 0 net=2833
rlabel metal2 114 -1125 114 -1125 0 net=815
rlabel metal2 135 -1125 135 -1125 0 net=1795
rlabel metal2 170 -1125 170 -1125 0 net=1527
rlabel metal2 240 -1125 240 -1125 0 net=830
rlabel metal2 310 -1125 310 -1125 0 net=2594
rlabel metal2 177 -1127 177 -1127 0 net=1456
rlabel metal2 205 -1127 205 -1127 0 net=1303
rlabel metal2 243 -1127 243 -1127 0 net=2797
rlabel metal2 184 -1129 184 -1129 0 net=918
rlabel metal2 198 -1129 198 -1129 0 net=855
rlabel metal2 247 -1129 247 -1129 0 net=1030
rlabel metal2 331 -1129 331 -1129 0 net=2139
rlabel metal2 163 -1131 163 -1131 0 net=919
rlabel metal2 226 -1131 226 -1131 0 net=583
rlabel metal2 254 -1133 254 -1133 0 net=1719
rlabel metal2 303 -1133 303 -1133 0 net=2937
rlabel metal2 156 -1135 156 -1135 0 net=1800
rlabel metal2 268 -1135 268 -1135 0 net=1665
rlabel metal2 324 -1135 324 -1135 0 net=2759
rlabel metal2 156 -1137 156 -1137 0 net=1673
rlabel metal2 250 -1137 250 -1137 0 net=2123
rlabel metal2 345 -1137 345 -1137 0 net=2439
rlabel metal2 177 -1139 177 -1139 0 net=1539
rlabel metal2 47 -1150 47 -1150 0 net=828
rlabel metal2 58 -1150 58 -1150 0 net=320
rlabel metal2 89 -1150 89 -1150 0 net=384
rlabel metal2 114 -1150 114 -1150 0 net=816
rlabel metal2 191 -1150 191 -1150 0 net=1129
rlabel metal2 212 -1150 212 -1150 0 net=1778
rlabel metal2 299 -1150 299 -1150 0 net=2841
rlabel metal2 394 -1150 394 -1150 0 net=2896
rlabel metal2 408 -1150 408 -1150 0 net=2986
rlabel metal2 422 -1150 422 -1150 0 net=2835
rlabel metal2 422 -1150 422 -1150 0 net=2835
rlabel metal2 446 -1150 446 -1150 0 net=2398
rlabel metal2 51 -1152 51 -1152 0 net=2443
rlabel metal2 65 -1152 65 -1152 0 net=2196
rlabel metal2 107 -1152 107 -1152 0 net=2029
rlabel metal2 135 -1152 135 -1152 0 net=2270
rlabel metal2 170 -1152 170 -1152 0 net=1529
rlabel metal2 194 -1152 194 -1152 0 net=1570
rlabel metal2 303 -1152 303 -1152 0 net=2760
rlabel metal2 65 -1154 65 -1154 0 net=220
rlabel metal2 212 -1154 212 -1154 0 net=1133
rlabel metal2 240 -1154 240 -1154 0 net=2228
rlabel metal2 100 -1156 100 -1156 0 net=1519
rlabel metal2 142 -1156 142 -1156 0 net=1796
rlabel metal2 177 -1156 177 -1156 0 net=1540
rlabel metal2 222 -1156 222 -1156 0 net=1304
rlabel metal2 243 -1156 243 -1156 0 net=1162
rlabel metal2 271 -1156 271 -1156 0 net=2170
rlabel metal2 324 -1156 324 -1156 0 net=2125
rlabel metal2 338 -1156 338 -1156 0 net=2377
rlabel metal2 100 -1158 100 -1158 0 net=1865
rlabel metal2 226 -1158 226 -1158 0 net=2440
rlabel metal2 359 -1158 359 -1158 0 net=2939
rlabel metal2 117 -1160 117 -1160 0 net=2480
rlabel metal2 128 -1160 128 -1160 0 net=1037
rlabel metal2 247 -1160 247 -1160 0 net=2605
rlabel metal2 121 -1162 121 -1162 0 net=1675
rlabel metal2 226 -1162 226 -1162 0 net=1845
rlabel metal2 306 -1162 306 -1162 0 net=2567
rlabel metal2 156 -1164 156 -1164 0 net=921
rlabel metal2 229 -1164 229 -1164 0 net=710
rlabel metal2 275 -1164 275 -1164 0 net=1721
rlabel metal2 275 -1164 275 -1164 0 net=1721
rlabel metal2 310 -1164 310 -1164 0 net=2777
rlabel metal2 198 -1166 198 -1166 0 net=857
rlabel metal2 296 -1166 296 -1166 0 net=2065
rlabel metal2 313 -1166 313 -1166 0 net=1498
rlabel metal2 233 -1168 233 -1168 0 net=1666
rlabel metal2 317 -1168 317 -1168 0 net=1725
rlabel metal2 415 -1168 415 -1168 0 net=2705
rlabel metal2 254 -1170 254 -1170 0 net=2207
rlabel metal2 324 -1170 324 -1170 0 net=2141
rlabel metal2 352 -1170 352 -1170 0 net=2799
rlabel metal2 247 -1172 247 -1172 0 net=2475
rlabel metal2 257 -1174 257 -1174 0 net=1941
rlabel metal2 47 -1187 47 -1187 0 net=412
rlabel metal2 47 -1187 47 -1187 0 net=412
rlabel metal2 51 -1187 51 -1187 0 net=2444
rlabel metal2 72 -1187 72 -1187 0 net=1255
rlabel metal2 89 -1187 89 -1187 0 net=721
rlabel metal2 100 -1187 100 -1187 0 net=1866
rlabel metal2 156 -1187 156 -1187 0 net=922
rlabel metal2 229 -1187 229 -1187 0 net=1722
rlabel metal2 289 -1187 289 -1187 0 net=2142
rlabel metal2 338 -1187 338 -1187 0 net=2378
rlabel metal2 380 -1187 380 -1187 0 net=2779
rlabel metal2 380 -1187 380 -1187 0 net=2779
rlabel metal2 408 -1187 408 -1187 0 net=2959
rlabel metal2 422 -1187 422 -1187 0 net=2837
rlabel metal2 65 -1189 65 -1189 0 net=134
rlabel metal2 93 -1189 93 -1189 0 net=1587
rlabel metal2 107 -1189 107 -1189 0 net=2030
rlabel metal2 166 -1189 166 -1189 0 net=1071
rlabel metal2 205 -1189 205 -1189 0 net=1131
rlabel metal2 205 -1189 205 -1189 0 net=1131
rlabel metal2 212 -1189 212 -1189 0 net=1135
rlabel metal2 212 -1189 212 -1189 0 net=1135
rlabel metal2 219 -1189 219 -1189 0 net=2066
rlabel metal2 324 -1189 324 -1189 0 net=2477
rlabel metal2 422 -1189 422 -1189 0 net=2706
rlabel metal2 79 -1191 79 -1191 0 net=174
rlabel metal2 170 -1191 170 -1191 0 net=2083
rlabel metal2 184 -1191 184 -1191 0 net=1530
rlabel metal2 229 -1191 229 -1191 0 net=1089
rlabel metal2 268 -1191 268 -1191 0 net=858
rlabel metal2 303 -1191 303 -1191 0 net=2126
rlabel metal2 345 -1191 345 -1191 0 net=2842
rlabel metal2 79 -1193 79 -1193 0 net=347
rlabel metal2 121 -1193 121 -1193 0 net=1676
rlabel metal2 159 -1193 159 -1193 0 net=1621
rlabel metal2 240 -1193 240 -1193 0 net=1726
rlabel metal2 331 -1193 331 -1193 0 net=1547
rlabel metal2 345 -1193 345 -1193 0 net=2801
rlabel metal2 107 -1195 107 -1195 0 net=2607
rlabel metal2 149 -1195 149 -1195 0 net=494
rlabel metal2 233 -1195 233 -1195 0 net=2317
rlabel metal2 247 -1195 247 -1195 0 net=2209
rlabel metal2 282 -1195 282 -1195 0 net=1846
rlabel metal2 317 -1195 317 -1195 0 net=2569
rlabel metal2 128 -1197 128 -1197 0 net=1038
rlabel metal2 236 -1197 236 -1197 0 net=2633
rlabel metal2 289 -1197 289 -1197 0 net=2606
rlabel metal2 128 -1199 128 -1199 0 net=979
rlabel metal2 184 -1199 184 -1199 0 net=353
rlabel metal2 292 -1199 292 -1199 0 net=2899
rlabel metal2 359 -1199 359 -1199 0 net=2941
rlabel metal2 135 -1201 135 -1201 0 net=1520
rlabel metal2 366 -1201 366 -1201 0 net=1943
rlabel metal2 121 -1203 121 -1203 0 net=1213
rlabel metal2 138 -1203 138 -1203 0 net=184
rlabel metal2 33 -1214 33 -1214 0 net=2523
rlabel metal2 44 -1214 44 -1214 0 net=2261
rlabel metal2 58 -1214 58 -1214 0 net=959
rlabel metal2 72 -1214 72 -1214 0 net=1256
rlabel metal2 89 -1214 89 -1214 0 net=1588
rlabel metal2 107 -1214 107 -1214 0 net=2608
rlabel metal2 180 -1214 180 -1214 0 net=1132
rlabel metal2 229 -1214 229 -1214 0 net=2210
rlabel metal2 254 -1214 254 -1214 0 net=1091
rlabel metal2 303 -1214 303 -1214 0 net=26
rlabel metal2 359 -1214 359 -1214 0 net=2943
rlabel metal2 359 -1214 359 -1214 0 net=2943
rlabel metal2 373 -1214 373 -1214 0 net=2780
rlabel metal2 401 -1214 401 -1214 0 net=2961
rlabel metal2 422 -1214 422 -1214 0 net=2839
rlabel metal2 72 -1216 72 -1216 0 net=1787
rlabel metal2 93 -1216 93 -1216 0 net=2271
rlabel metal2 152 -1216 152 -1216 0 net=681
rlabel metal2 163 -1216 163 -1216 0 net=1136
rlabel metal2 229 -1216 229 -1216 0 net=1117
rlabel metal2 243 -1216 243 -1216 0 net=342
rlabel metal2 296 -1216 296 -1216 0 net=2901
rlabel metal2 306 -1216 306 -1216 0 net=2478
rlabel metal2 331 -1216 331 -1216 0 net=1548
rlabel metal2 425 -1216 425 -1216 0 net=89
rlabel metal2 114 -1218 114 -1218 0 net=1214
rlabel metal2 128 -1218 128 -1218 0 net=980
rlabel metal2 163 -1218 163 -1218 0 net=1623
rlabel metal2 184 -1218 184 -1218 0 net=1573
rlabel metal2 212 -1218 212 -1218 0 net=1663
rlabel metal2 275 -1218 275 -1218 0 net=1855
rlabel metal2 310 -1218 310 -1218 0 net=2802
rlabel metal2 352 -1218 352 -1218 0 net=1945
rlabel metal2 100 -1220 100 -1220 0 net=851
rlabel metal2 135 -1220 135 -1220 0 net=235
rlabel metal2 170 -1220 170 -1220 0 net=2084
rlabel metal2 191 -1220 191 -1220 0 net=1025
rlabel metal2 282 -1220 282 -1220 0 net=2635
rlabel metal2 317 -1220 317 -1220 0 net=2570
rlabel metal2 338 -1220 338 -1220 0 net=2257
rlabel metal2 366 -1220 366 -1220 0 net=2819
rlabel metal2 121 -1222 121 -1222 0 net=1909
rlabel metal2 194 -1222 194 -1222 0 net=1072
rlabel metal2 215 -1222 215 -1222 0 net=80
rlabel metal2 124 -1224 124 -1224 0 net=2533
rlabel metal2 222 -1224 222 -1224 0 net=2318
rlabel metal2 282 -1224 282 -1224 0 net=1861
rlabel metal2 219 -1226 219 -1226 0 net=1571
rlabel metal2 23 -1237 23 -1237 0 net=198
rlabel metal2 23 -1237 23 -1237 0 net=198
rlabel metal2 30 -1237 30 -1237 0 net=2525
rlabel metal2 44 -1237 44 -1237 0 net=2262
rlabel metal2 58 -1237 58 -1237 0 net=961
rlabel metal2 58 -1237 58 -1237 0 net=961
rlabel metal2 65 -1237 65 -1237 0 net=364
rlabel metal2 79 -1237 79 -1237 0 net=1789
rlabel metal2 79 -1237 79 -1237 0 net=1789
rlabel metal2 93 -1237 93 -1237 0 net=2272
rlabel metal2 128 -1237 128 -1237 0 net=1910
rlabel metal2 152 -1237 152 -1237 0 net=247
rlabel metal2 222 -1237 222 -1237 0 net=1092
rlabel metal2 275 -1237 275 -1237 0 net=1857
rlabel metal2 299 -1237 299 -1237 0 net=2636
rlabel metal2 324 -1237 324 -1237 0 net=2661
rlabel metal2 334 -1237 334 -1237 0 net=2258
rlabel metal2 359 -1237 359 -1237 0 net=2945
rlabel metal2 359 -1237 359 -1237 0 net=2945
rlabel metal2 369 -1237 369 -1237 0 net=2820
rlabel metal2 401 -1237 401 -1237 0 net=2962
rlabel metal2 415 -1237 415 -1237 0 net=2840
rlabel metal2 100 -1239 100 -1239 0 net=852
rlabel metal2 128 -1239 128 -1239 0 net=997
rlabel metal2 142 -1239 142 -1239 0 net=2534
rlabel metal2 159 -1239 159 -1239 0 net=201
rlabel metal2 159 -1239 159 -1239 0 net=201
rlabel metal2 163 -1239 163 -1239 0 net=1624
rlabel metal2 226 -1239 226 -1239 0 net=267
rlabel metal2 303 -1239 303 -1239 0 net=2903
rlabel metal2 303 -1239 303 -1239 0 net=2903
rlabel metal2 338 -1239 338 -1239 0 net=1947
rlabel metal2 103 -1241 103 -1241 0 net=1445
rlabel metal2 177 -1241 177 -1241 0 net=1027
rlabel metal2 194 -1241 194 -1241 0 net=1118
rlabel metal2 250 -1241 250 -1241 0 net=2781
rlabel metal2 110 -1243 110 -1243 0 net=897
rlabel metal2 205 -1243 205 -1243 0 net=1862
rlabel metal2 208 -1245 208 -1245 0 net=1664
rlabel metal2 261 -1245 261 -1245 0 net=1905
rlabel metal2 261 -1245 261 -1245 0 net=1905
rlabel metal2 212 -1247 212 -1247 0 net=2241
rlabel metal2 233 -1247 233 -1247 0 net=1572
rlabel metal2 170 -1249 170 -1249 0 net=1617
rlabel metal2 170 -1251 170 -1251 0 net=1575
rlabel metal2 219 -1251 219 -1251 0 net=314
rlabel metal2 30 -1262 30 -1262 0 net=2526
rlabel metal2 58 -1262 58 -1262 0 net=962
rlabel metal2 72 -1262 72 -1262 0 net=1790
rlabel metal2 107 -1262 107 -1262 0 net=898
rlabel metal2 121 -1262 121 -1262 0 net=1446
rlabel metal2 170 -1262 170 -1262 0 net=1576
rlabel metal2 208 -1262 208 -1262 0 net=2242
rlabel metal2 226 -1262 226 -1262 0 net=2782
rlabel metal2 285 -1262 285 -1262 0 net=1858
rlabel metal2 296 -1262 296 -1262 0 net=2904
rlabel metal2 317 -1262 317 -1262 0 net=2662
rlabel metal2 338 -1262 338 -1262 0 net=1948
rlabel metal2 355 -1262 355 -1262 0 net=2946
rlabel metal2 128 -1264 128 -1264 0 net=998
rlabel metal2 142 -1264 142 -1264 0 net=66
rlabel metal2 177 -1264 177 -1264 0 net=1028
rlabel metal2 198 -1264 198 -1264 0 net=1618
rlabel metal2 250 -1264 250 -1264 0 net=1906
<< end >>
