magic
tech scmos
timestamp 1555071848 
<< pdiffusion >>
rect 1 -14 7 -8
rect 8 -14 14 -8
rect 15 -14 21 -8
rect 22 -14 28 -8
rect 29 -14 35 -8
rect 36 -14 42 -8
rect 43 -14 49 -8
rect 50 -14 56 -8
rect 57 -14 63 -8
rect 64 -14 70 -8
rect 71 -14 77 -8
rect 78 -14 84 -8
rect 85 -14 91 -8
rect 92 -14 98 -8
rect 99 -14 105 -8
rect 106 -14 112 -8
rect 113 -14 119 -8
rect 120 -14 126 -8
rect 127 -14 133 -8
rect 134 -14 140 -8
rect 141 -14 147 -8
rect 148 -14 154 -8
rect 155 -14 161 -8
rect 162 -14 168 -8
rect 169 -14 175 -8
rect 225 -14 228 -8
rect 253 -14 256 -8
rect 274 -14 277 -8
rect 316 -14 319 -8
rect 330 -14 336 -8
rect 365 -14 368 -8
rect 372 -14 378 -8
rect 379 -14 385 -8
rect 393 -14 399 -8
rect 400 -14 406 -8
rect 414 -14 417 -8
rect 428 -14 434 -8
rect 435 -14 438 -8
rect 442 -14 448 -8
rect 449 -14 452 -8
rect 456 -14 462 -8
rect 470 -14 473 -8
rect 491 -14 494 -8
rect 505 -14 508 -8
rect 512 -14 518 -8
rect 526 -14 529 -8
rect 533 -14 539 -8
rect 540 -14 546 -8
rect 561 -14 567 -8
rect 568 -14 571 -8
rect 589 -14 592 -8
rect 617 -14 623 -8
rect 638 -14 644 -8
rect 666 -14 672 -8
rect 673 -14 676 -8
rect 701 -14 707 -8
rect 764 -14 767 -8
rect 799 -14 805 -8
rect 827 -14 830 -8
rect 841 -14 844 -8
rect 1 -43 7 -37
rect 8 -43 14 -37
rect 15 -43 21 -37
rect 22 -43 28 -37
rect 29 -43 35 -37
rect 36 -43 42 -37
rect 43 -43 49 -37
rect 50 -43 56 -37
rect 57 -43 63 -37
rect 64 -43 70 -37
rect 71 -43 77 -37
rect 78 -43 84 -37
rect 85 -43 91 -37
rect 92 -43 98 -37
rect 99 -43 105 -37
rect 106 -43 112 -37
rect 113 -43 119 -37
rect 120 -43 126 -37
rect 127 -43 133 -37
rect 134 -43 137 -37
rect 141 -43 147 -37
rect 148 -43 154 -37
rect 176 -43 182 -37
rect 190 -43 193 -37
rect 204 -43 207 -37
rect 211 -43 214 -37
rect 218 -43 224 -37
rect 225 -43 228 -37
rect 232 -43 238 -37
rect 253 -43 256 -37
rect 295 -43 301 -37
rect 302 -43 305 -37
rect 309 -43 315 -37
rect 316 -43 319 -37
rect 323 -43 329 -37
rect 330 -43 333 -37
rect 337 -43 340 -37
rect 344 -43 347 -37
rect 351 -43 354 -37
rect 358 -43 361 -37
rect 365 -43 371 -37
rect 372 -43 375 -37
rect 379 -43 382 -37
rect 386 -43 389 -37
rect 393 -43 399 -37
rect 400 -43 406 -37
rect 407 -43 410 -37
rect 414 -43 417 -37
rect 421 -43 424 -37
rect 442 -43 448 -37
rect 449 -43 455 -37
rect 456 -43 459 -37
rect 463 -43 469 -37
rect 470 -43 473 -37
rect 477 -43 480 -37
rect 484 -43 490 -37
rect 491 -43 494 -37
rect 512 -43 515 -37
rect 519 -43 522 -37
rect 526 -43 529 -37
rect 533 -43 536 -37
rect 540 -43 543 -37
rect 547 -43 550 -37
rect 554 -43 557 -37
rect 568 -43 571 -37
rect 575 -43 578 -37
rect 582 -43 585 -37
rect 589 -43 595 -37
rect 617 -43 623 -37
rect 631 -43 637 -37
rect 638 -43 641 -37
rect 645 -43 648 -37
rect 652 -43 655 -37
rect 659 -43 662 -37
rect 666 -43 669 -37
rect 680 -43 686 -37
rect 694 -43 697 -37
rect 701 -43 704 -37
rect 708 -43 711 -37
rect 757 -43 763 -37
rect 764 -43 767 -37
rect 771 -43 777 -37
rect 778 -43 784 -37
rect 785 -43 788 -37
rect 792 -43 795 -37
rect 799 -43 802 -37
rect 820 -43 826 -37
rect 855 -43 858 -37
rect 876 -43 879 -37
rect 918 -43 921 -37
rect 1 -92 7 -86
rect 8 -92 14 -86
rect 15 -92 21 -86
rect 22 -92 28 -86
rect 29 -92 35 -86
rect 36 -92 42 -86
rect 43 -92 49 -86
rect 50 -92 56 -86
rect 57 -92 63 -86
rect 64 -92 70 -86
rect 71 -92 77 -86
rect 78 -92 81 -86
rect 85 -92 91 -86
rect 92 -92 98 -86
rect 99 -92 102 -86
rect 106 -92 112 -86
rect 113 -92 119 -86
rect 120 -92 126 -86
rect 127 -92 130 -86
rect 134 -92 140 -86
rect 141 -92 147 -86
rect 148 -92 151 -86
rect 155 -92 158 -86
rect 162 -92 165 -86
rect 169 -92 172 -86
rect 176 -92 182 -86
rect 183 -92 186 -86
rect 190 -92 193 -86
rect 197 -92 200 -86
rect 204 -92 207 -86
rect 211 -92 217 -86
rect 218 -92 221 -86
rect 225 -92 231 -86
rect 232 -92 238 -86
rect 239 -92 245 -86
rect 246 -92 252 -86
rect 253 -92 256 -86
rect 260 -92 263 -86
rect 267 -92 270 -86
rect 274 -92 280 -86
rect 281 -92 287 -86
rect 288 -92 291 -86
rect 295 -92 301 -86
rect 302 -92 305 -86
rect 309 -92 312 -86
rect 316 -92 319 -86
rect 323 -92 326 -86
rect 330 -92 336 -86
rect 337 -92 340 -86
rect 344 -92 347 -86
rect 351 -92 354 -86
rect 358 -92 361 -86
rect 365 -92 371 -86
rect 372 -92 375 -86
rect 379 -92 382 -86
rect 386 -92 392 -86
rect 393 -92 399 -86
rect 400 -92 403 -86
rect 407 -92 410 -86
rect 414 -92 417 -86
rect 421 -92 424 -86
rect 428 -92 431 -86
rect 435 -92 438 -86
rect 442 -92 448 -86
rect 449 -92 455 -86
rect 456 -92 459 -86
rect 463 -92 466 -86
rect 470 -92 476 -86
rect 477 -92 480 -86
rect 484 -92 487 -86
rect 491 -92 494 -86
rect 498 -92 501 -86
rect 505 -92 508 -86
rect 512 -92 515 -86
rect 519 -92 522 -86
rect 526 -92 529 -86
rect 533 -92 536 -86
rect 540 -92 543 -86
rect 547 -92 550 -86
rect 554 -92 557 -86
rect 561 -92 564 -86
rect 568 -92 574 -86
rect 575 -92 578 -86
rect 582 -92 585 -86
rect 589 -92 595 -86
rect 596 -92 599 -86
rect 603 -92 606 -86
rect 610 -92 613 -86
rect 617 -92 620 -86
rect 624 -92 630 -86
rect 631 -92 634 -86
rect 638 -92 644 -86
rect 645 -92 648 -86
rect 652 -92 655 -86
rect 659 -92 662 -86
rect 666 -92 669 -86
rect 673 -92 676 -86
rect 680 -92 683 -86
rect 687 -92 690 -86
rect 694 -92 697 -86
rect 701 -92 704 -86
rect 708 -92 711 -86
rect 715 -92 718 -86
rect 722 -92 725 -86
rect 729 -92 735 -86
rect 736 -92 742 -86
rect 743 -92 746 -86
rect 750 -92 753 -86
rect 757 -92 763 -86
rect 764 -92 767 -86
rect 771 -92 774 -86
rect 778 -92 784 -86
rect 785 -92 788 -86
rect 792 -92 795 -86
rect 799 -92 802 -86
rect 806 -92 809 -86
rect 813 -92 816 -86
rect 820 -92 823 -86
rect 855 -92 858 -86
rect 862 -92 865 -86
rect 869 -92 872 -86
rect 890 -92 893 -86
rect 904 -92 907 -86
rect 967 -92 970 -86
rect 1 -163 7 -157
rect 8 -163 14 -157
rect 15 -163 21 -157
rect 22 -163 28 -157
rect 29 -163 35 -157
rect 36 -163 42 -157
rect 43 -163 49 -157
rect 50 -163 56 -157
rect 57 -163 63 -157
rect 64 -163 70 -157
rect 71 -163 77 -157
rect 78 -163 84 -157
rect 85 -163 91 -157
rect 92 -163 98 -157
rect 99 -163 105 -157
rect 106 -163 112 -157
rect 113 -163 116 -157
rect 120 -163 126 -157
rect 127 -163 133 -157
rect 148 -163 151 -157
rect 155 -163 161 -157
rect 162 -163 165 -157
rect 169 -163 172 -157
rect 176 -163 179 -157
rect 183 -163 186 -157
rect 190 -163 193 -157
rect 197 -163 200 -157
rect 204 -163 207 -157
rect 211 -163 214 -157
rect 218 -163 221 -157
rect 225 -163 228 -157
rect 232 -163 235 -157
rect 239 -163 242 -157
rect 246 -163 252 -157
rect 253 -163 259 -157
rect 260 -163 263 -157
rect 267 -163 273 -157
rect 274 -163 280 -157
rect 281 -163 287 -157
rect 288 -163 294 -157
rect 295 -163 301 -157
rect 302 -163 305 -157
rect 309 -163 312 -157
rect 316 -163 319 -157
rect 323 -163 326 -157
rect 330 -163 333 -157
rect 337 -163 340 -157
rect 344 -163 347 -157
rect 351 -163 354 -157
rect 358 -163 361 -157
rect 365 -163 368 -157
rect 372 -163 375 -157
rect 379 -163 382 -157
rect 386 -163 392 -157
rect 393 -163 396 -157
rect 400 -163 403 -157
rect 407 -163 410 -157
rect 414 -163 420 -157
rect 421 -163 424 -157
rect 428 -163 434 -157
rect 435 -163 438 -157
rect 442 -163 445 -157
rect 449 -163 452 -157
rect 456 -163 459 -157
rect 463 -163 469 -157
rect 470 -163 476 -157
rect 477 -163 480 -157
rect 484 -163 490 -157
rect 491 -163 494 -157
rect 498 -163 501 -157
rect 505 -163 511 -157
rect 512 -163 515 -157
rect 519 -163 522 -157
rect 526 -163 529 -157
rect 533 -163 536 -157
rect 540 -163 543 -157
rect 547 -163 550 -157
rect 554 -163 560 -157
rect 561 -163 564 -157
rect 568 -163 571 -157
rect 575 -163 578 -157
rect 582 -163 585 -157
rect 589 -163 592 -157
rect 596 -163 599 -157
rect 603 -163 606 -157
rect 610 -163 613 -157
rect 617 -163 623 -157
rect 624 -163 627 -157
rect 631 -163 634 -157
rect 638 -163 641 -157
rect 645 -163 648 -157
rect 652 -163 655 -157
rect 659 -163 662 -157
rect 666 -163 669 -157
rect 673 -163 676 -157
rect 680 -163 686 -157
rect 687 -163 690 -157
rect 694 -163 700 -157
rect 701 -163 707 -157
rect 708 -163 711 -157
rect 715 -163 718 -157
rect 722 -163 725 -157
rect 729 -163 732 -157
rect 736 -163 739 -157
rect 743 -163 746 -157
rect 750 -163 756 -157
rect 757 -163 760 -157
rect 764 -163 767 -157
rect 771 -163 774 -157
rect 778 -163 781 -157
rect 785 -163 788 -157
rect 792 -163 795 -157
rect 799 -163 802 -157
rect 806 -163 809 -157
rect 813 -163 816 -157
rect 820 -163 823 -157
rect 827 -163 830 -157
rect 834 -163 837 -157
rect 841 -163 844 -157
rect 848 -163 851 -157
rect 855 -163 858 -157
rect 862 -163 865 -157
rect 869 -163 872 -157
rect 876 -163 879 -157
rect 883 -163 886 -157
rect 890 -163 893 -157
rect 897 -163 900 -157
rect 904 -163 907 -157
rect 911 -163 914 -157
rect 918 -163 921 -157
rect 925 -163 928 -157
rect 932 -163 935 -157
rect 939 -163 945 -157
rect 946 -163 952 -157
rect 953 -163 956 -157
rect 960 -163 963 -157
rect 967 -163 970 -157
rect 974 -163 977 -157
rect 981 -163 984 -157
rect 988 -163 991 -157
rect 995 -163 1001 -157
rect 1002 -163 1005 -157
rect 1 -258 7 -252
rect 8 -258 14 -252
rect 15 -258 21 -252
rect 22 -258 28 -252
rect 29 -258 35 -252
rect 36 -258 42 -252
rect 43 -258 49 -252
rect 50 -258 56 -252
rect 57 -258 63 -252
rect 64 -258 70 -252
rect 71 -258 74 -252
rect 78 -258 84 -252
rect 85 -258 91 -252
rect 92 -258 98 -252
rect 99 -258 102 -252
rect 106 -258 112 -252
rect 113 -258 116 -252
rect 120 -258 126 -252
rect 127 -258 130 -252
rect 134 -258 137 -252
rect 141 -258 147 -252
rect 148 -258 154 -252
rect 155 -258 161 -252
rect 162 -258 168 -252
rect 169 -258 175 -252
rect 176 -258 179 -252
rect 183 -258 186 -252
rect 190 -258 193 -252
rect 197 -258 200 -252
rect 204 -258 210 -252
rect 211 -258 214 -252
rect 218 -258 224 -252
rect 225 -258 228 -252
rect 232 -258 235 -252
rect 239 -258 245 -252
rect 246 -258 249 -252
rect 253 -258 256 -252
rect 260 -258 263 -252
rect 267 -258 270 -252
rect 274 -258 277 -252
rect 281 -258 287 -252
rect 288 -258 291 -252
rect 295 -258 298 -252
rect 302 -258 305 -252
rect 309 -258 312 -252
rect 316 -258 322 -252
rect 323 -258 326 -252
rect 330 -258 333 -252
rect 337 -258 343 -252
rect 344 -258 347 -252
rect 351 -258 354 -252
rect 358 -258 361 -252
rect 365 -258 368 -252
rect 372 -258 375 -252
rect 379 -258 382 -252
rect 386 -258 389 -252
rect 393 -258 396 -252
rect 400 -258 406 -252
rect 407 -258 410 -252
rect 414 -258 417 -252
rect 421 -258 424 -252
rect 428 -258 434 -252
rect 435 -258 438 -252
rect 442 -258 448 -252
rect 449 -258 455 -252
rect 456 -258 459 -252
rect 463 -258 466 -252
rect 470 -258 473 -252
rect 477 -258 483 -252
rect 484 -258 490 -252
rect 491 -258 497 -252
rect 498 -258 501 -252
rect 505 -258 508 -252
rect 512 -258 518 -252
rect 519 -258 522 -252
rect 526 -258 529 -252
rect 533 -258 539 -252
rect 540 -258 546 -252
rect 547 -258 550 -252
rect 554 -258 557 -252
rect 561 -258 564 -252
rect 568 -258 571 -252
rect 575 -258 578 -252
rect 582 -258 588 -252
rect 589 -258 592 -252
rect 596 -258 599 -252
rect 603 -258 606 -252
rect 610 -258 616 -252
rect 617 -258 620 -252
rect 624 -258 627 -252
rect 631 -258 634 -252
rect 638 -258 641 -252
rect 645 -258 648 -252
rect 652 -258 655 -252
rect 659 -258 662 -252
rect 666 -258 669 -252
rect 673 -258 676 -252
rect 680 -258 686 -252
rect 687 -258 690 -252
rect 694 -258 697 -252
rect 701 -258 704 -252
rect 708 -258 711 -252
rect 715 -258 718 -252
rect 722 -258 725 -252
rect 729 -258 732 -252
rect 736 -258 739 -252
rect 743 -258 746 -252
rect 750 -258 753 -252
rect 757 -258 760 -252
rect 764 -258 770 -252
rect 771 -258 774 -252
rect 778 -258 781 -252
rect 785 -258 788 -252
rect 792 -258 795 -252
rect 799 -258 802 -252
rect 806 -258 809 -252
rect 813 -258 816 -252
rect 820 -258 823 -252
rect 827 -258 833 -252
rect 834 -258 837 -252
rect 841 -258 847 -252
rect 848 -258 851 -252
rect 855 -258 858 -252
rect 862 -258 865 -252
rect 869 -258 872 -252
rect 876 -258 879 -252
rect 883 -258 886 -252
rect 890 -258 893 -252
rect 897 -258 900 -252
rect 904 -258 907 -252
rect 911 -258 914 -252
rect 918 -258 921 -252
rect 925 -258 928 -252
rect 932 -258 935 -252
rect 939 -258 942 -252
rect 946 -258 949 -252
rect 953 -258 956 -252
rect 960 -258 963 -252
rect 967 -258 970 -252
rect 974 -258 977 -252
rect 981 -258 984 -252
rect 988 -258 991 -252
rect 995 -258 998 -252
rect 1002 -258 1005 -252
rect 1009 -258 1012 -252
rect 1016 -258 1019 -252
rect 1023 -258 1026 -252
rect 1030 -258 1033 -252
rect 1037 -258 1040 -252
rect 1044 -258 1047 -252
rect 1051 -258 1054 -252
rect 1058 -258 1061 -252
rect 1065 -258 1068 -252
rect 1072 -258 1075 -252
rect 1079 -258 1082 -252
rect 1086 -258 1089 -252
rect 1093 -258 1096 -252
rect 1100 -258 1103 -252
rect 1107 -258 1110 -252
rect 1114 -258 1117 -252
rect 1121 -258 1124 -252
rect 1128 -258 1131 -252
rect 1 -361 7 -355
rect 8 -361 14 -355
rect 15 -361 21 -355
rect 22 -361 28 -355
rect 29 -361 35 -355
rect 36 -361 42 -355
rect 43 -361 49 -355
rect 50 -361 53 -355
rect 57 -361 63 -355
rect 64 -361 70 -355
rect 71 -361 77 -355
rect 78 -361 84 -355
rect 85 -361 88 -355
rect 92 -361 95 -355
rect 99 -361 102 -355
rect 106 -361 109 -355
rect 113 -361 116 -355
rect 120 -361 126 -355
rect 127 -361 130 -355
rect 134 -361 137 -355
rect 141 -361 144 -355
rect 148 -361 151 -355
rect 155 -361 161 -355
rect 162 -361 165 -355
rect 169 -361 175 -355
rect 176 -361 179 -355
rect 183 -361 186 -355
rect 190 -361 193 -355
rect 197 -361 200 -355
rect 204 -361 207 -355
rect 211 -361 214 -355
rect 218 -361 221 -355
rect 225 -361 228 -355
rect 232 -361 238 -355
rect 239 -361 242 -355
rect 246 -361 252 -355
rect 253 -361 256 -355
rect 260 -361 266 -355
rect 267 -361 270 -355
rect 274 -361 277 -355
rect 281 -361 287 -355
rect 288 -361 291 -355
rect 295 -361 298 -355
rect 302 -361 305 -355
rect 309 -361 312 -355
rect 316 -361 319 -355
rect 323 -361 326 -355
rect 330 -361 336 -355
rect 337 -361 340 -355
rect 344 -361 347 -355
rect 351 -361 354 -355
rect 358 -361 364 -355
rect 365 -361 371 -355
rect 372 -361 375 -355
rect 379 -361 382 -355
rect 386 -361 389 -355
rect 393 -361 396 -355
rect 400 -361 403 -355
rect 407 -361 410 -355
rect 414 -361 417 -355
rect 421 -361 424 -355
rect 428 -361 431 -355
rect 435 -361 438 -355
rect 442 -361 445 -355
rect 449 -361 452 -355
rect 456 -361 459 -355
rect 463 -361 469 -355
rect 470 -361 476 -355
rect 477 -361 483 -355
rect 484 -361 490 -355
rect 491 -361 497 -355
rect 498 -361 501 -355
rect 505 -361 508 -355
rect 512 -361 518 -355
rect 519 -361 522 -355
rect 526 -361 532 -355
rect 533 -361 536 -355
rect 540 -361 543 -355
rect 547 -361 550 -355
rect 554 -361 557 -355
rect 561 -361 567 -355
rect 568 -361 574 -355
rect 575 -361 581 -355
rect 582 -361 588 -355
rect 589 -361 595 -355
rect 596 -361 599 -355
rect 603 -361 609 -355
rect 610 -361 613 -355
rect 617 -361 620 -355
rect 624 -361 627 -355
rect 631 -361 637 -355
rect 638 -361 641 -355
rect 645 -361 648 -355
rect 652 -361 655 -355
rect 659 -361 665 -355
rect 666 -361 669 -355
rect 673 -361 676 -355
rect 680 -361 686 -355
rect 687 -361 690 -355
rect 694 -361 697 -355
rect 701 -361 704 -355
rect 708 -361 711 -355
rect 715 -361 721 -355
rect 722 -361 728 -355
rect 729 -361 732 -355
rect 736 -361 739 -355
rect 743 -361 746 -355
rect 750 -361 753 -355
rect 757 -361 760 -355
rect 764 -361 767 -355
rect 771 -361 777 -355
rect 778 -361 781 -355
rect 785 -361 791 -355
rect 792 -361 795 -355
rect 799 -361 802 -355
rect 806 -361 809 -355
rect 813 -361 816 -355
rect 820 -361 823 -355
rect 827 -361 830 -355
rect 834 -361 837 -355
rect 841 -361 844 -355
rect 848 -361 851 -355
rect 855 -361 858 -355
rect 862 -361 865 -355
rect 869 -361 872 -355
rect 876 -361 879 -355
rect 883 -361 886 -355
rect 890 -361 893 -355
rect 897 -361 900 -355
rect 904 -361 907 -355
rect 911 -361 914 -355
rect 918 -361 921 -355
rect 925 -361 928 -355
rect 932 -361 935 -355
rect 939 -361 942 -355
rect 946 -361 949 -355
rect 953 -361 956 -355
rect 960 -361 963 -355
rect 967 -361 970 -355
rect 974 -361 977 -355
rect 981 -361 984 -355
rect 988 -361 991 -355
rect 995 -361 998 -355
rect 1002 -361 1005 -355
rect 1009 -361 1012 -355
rect 1016 -361 1019 -355
rect 1023 -361 1026 -355
rect 1030 -361 1033 -355
rect 1037 -361 1040 -355
rect 1044 -361 1047 -355
rect 1051 -361 1054 -355
rect 1058 -361 1061 -355
rect 1065 -361 1068 -355
rect 1072 -361 1075 -355
rect 1079 -361 1082 -355
rect 1086 -361 1089 -355
rect 1093 -361 1096 -355
rect 1100 -361 1103 -355
rect 1107 -361 1110 -355
rect 1114 -361 1117 -355
rect 1121 -361 1124 -355
rect 1128 -361 1131 -355
rect 1135 -361 1138 -355
rect 1142 -361 1145 -355
rect 1149 -361 1152 -355
rect 1156 -361 1159 -355
rect 1163 -361 1166 -355
rect 1170 -361 1173 -355
rect 1177 -361 1180 -355
rect 1184 -361 1187 -355
rect 1191 -361 1194 -355
rect 1198 -361 1201 -355
rect 1205 -361 1208 -355
rect 1212 -361 1215 -355
rect 1219 -361 1222 -355
rect 1226 -361 1229 -355
rect 1233 -361 1236 -355
rect 1240 -361 1243 -355
rect 1247 -361 1250 -355
rect 1254 -361 1257 -355
rect 1261 -361 1264 -355
rect 1268 -361 1271 -355
rect 1275 -361 1278 -355
rect 1282 -361 1285 -355
rect 1289 -361 1292 -355
rect 1296 -361 1302 -355
rect 1 -486 7 -480
rect 8 -486 14 -480
rect 15 -486 21 -480
rect 22 -486 28 -480
rect 29 -486 35 -480
rect 36 -486 42 -480
rect 43 -486 49 -480
rect 50 -486 56 -480
rect 57 -486 63 -480
rect 64 -486 67 -480
rect 71 -486 74 -480
rect 78 -486 81 -480
rect 85 -486 88 -480
rect 92 -486 98 -480
rect 99 -486 102 -480
rect 106 -486 109 -480
rect 113 -486 119 -480
rect 120 -486 126 -480
rect 127 -486 133 -480
rect 134 -486 137 -480
rect 141 -486 144 -480
rect 148 -486 154 -480
rect 155 -486 158 -480
rect 162 -486 165 -480
rect 169 -486 172 -480
rect 176 -486 179 -480
rect 183 -486 186 -480
rect 190 -486 193 -480
rect 197 -486 200 -480
rect 204 -486 207 -480
rect 211 -486 217 -480
rect 218 -486 221 -480
rect 225 -486 228 -480
rect 232 -486 235 -480
rect 239 -486 242 -480
rect 246 -486 249 -480
rect 253 -486 256 -480
rect 260 -486 263 -480
rect 267 -486 273 -480
rect 274 -486 280 -480
rect 281 -486 287 -480
rect 288 -486 294 -480
rect 295 -486 298 -480
rect 302 -486 305 -480
rect 309 -486 312 -480
rect 316 -486 319 -480
rect 323 -486 326 -480
rect 330 -486 333 -480
rect 337 -486 340 -480
rect 344 -486 347 -480
rect 351 -486 357 -480
rect 358 -486 361 -480
rect 365 -486 368 -480
rect 372 -486 375 -480
rect 379 -486 382 -480
rect 386 -486 389 -480
rect 393 -486 396 -480
rect 400 -486 403 -480
rect 407 -486 410 -480
rect 414 -486 417 -480
rect 421 -486 424 -480
rect 428 -486 431 -480
rect 435 -486 438 -480
rect 442 -486 445 -480
rect 449 -486 452 -480
rect 456 -486 462 -480
rect 463 -486 466 -480
rect 470 -486 473 -480
rect 477 -486 480 -480
rect 484 -486 487 -480
rect 491 -486 494 -480
rect 498 -486 504 -480
rect 505 -486 508 -480
rect 512 -486 518 -480
rect 519 -486 522 -480
rect 526 -486 529 -480
rect 533 -486 539 -480
rect 540 -486 543 -480
rect 547 -486 550 -480
rect 554 -486 560 -480
rect 561 -486 564 -480
rect 568 -486 571 -480
rect 575 -486 581 -480
rect 582 -486 585 -480
rect 589 -486 592 -480
rect 596 -486 602 -480
rect 603 -486 606 -480
rect 610 -486 616 -480
rect 617 -486 620 -480
rect 624 -486 627 -480
rect 631 -486 637 -480
rect 638 -486 644 -480
rect 645 -486 648 -480
rect 652 -486 655 -480
rect 659 -486 662 -480
rect 666 -486 669 -480
rect 673 -486 679 -480
rect 680 -486 686 -480
rect 687 -486 693 -480
rect 694 -486 700 -480
rect 701 -486 704 -480
rect 708 -486 711 -480
rect 715 -486 721 -480
rect 722 -486 725 -480
rect 729 -486 732 -480
rect 736 -486 739 -480
rect 743 -486 746 -480
rect 750 -486 756 -480
rect 757 -486 763 -480
rect 764 -486 767 -480
rect 771 -486 777 -480
rect 778 -486 781 -480
rect 785 -486 791 -480
rect 792 -486 795 -480
rect 799 -486 802 -480
rect 806 -486 809 -480
rect 813 -486 816 -480
rect 820 -486 823 -480
rect 827 -486 833 -480
rect 834 -486 837 -480
rect 841 -486 844 -480
rect 848 -486 851 -480
rect 855 -486 858 -480
rect 862 -486 865 -480
rect 869 -486 872 -480
rect 876 -486 879 -480
rect 883 -486 889 -480
rect 890 -486 893 -480
rect 897 -486 900 -480
rect 904 -486 907 -480
rect 911 -486 914 -480
rect 918 -486 921 -480
rect 925 -486 928 -480
rect 932 -486 935 -480
rect 939 -486 942 -480
rect 946 -486 949 -480
rect 953 -486 956 -480
rect 960 -486 963 -480
rect 967 -486 970 -480
rect 974 -486 977 -480
rect 981 -486 984 -480
rect 988 -486 991 -480
rect 995 -486 998 -480
rect 1002 -486 1005 -480
rect 1009 -486 1012 -480
rect 1016 -486 1019 -480
rect 1023 -486 1026 -480
rect 1030 -486 1033 -480
rect 1037 -486 1040 -480
rect 1044 -486 1047 -480
rect 1051 -486 1054 -480
rect 1058 -486 1061 -480
rect 1065 -486 1068 -480
rect 1072 -486 1075 -480
rect 1079 -486 1082 -480
rect 1086 -486 1089 -480
rect 1093 -486 1096 -480
rect 1100 -486 1103 -480
rect 1107 -486 1110 -480
rect 1114 -486 1117 -480
rect 1121 -486 1124 -480
rect 1128 -486 1131 -480
rect 1135 -486 1138 -480
rect 1142 -486 1145 -480
rect 1149 -486 1152 -480
rect 1156 -486 1159 -480
rect 1163 -486 1166 -480
rect 1170 -486 1173 -480
rect 1177 -486 1180 -480
rect 1184 -486 1187 -480
rect 1191 -486 1194 -480
rect 1198 -486 1201 -480
rect 1205 -486 1208 -480
rect 1212 -486 1215 -480
rect 1219 -486 1222 -480
rect 1226 -486 1229 -480
rect 1233 -486 1236 -480
rect 1240 -486 1243 -480
rect 1247 -486 1250 -480
rect 1254 -486 1257 -480
rect 1261 -486 1264 -480
rect 1268 -486 1271 -480
rect 1275 -486 1278 -480
rect 1282 -486 1285 -480
rect 1289 -486 1292 -480
rect 1296 -486 1299 -480
rect 1303 -486 1306 -480
rect 1310 -486 1313 -480
rect 1317 -486 1320 -480
rect 1324 -486 1327 -480
rect 1331 -486 1334 -480
rect 1338 -486 1341 -480
rect 1345 -486 1348 -480
rect 1352 -486 1355 -480
rect 1359 -486 1362 -480
rect 1366 -486 1369 -480
rect 1373 -486 1379 -480
rect 1 -619 7 -613
rect 8 -619 14 -613
rect 15 -619 21 -613
rect 22 -619 28 -613
rect 29 -619 35 -613
rect 36 -619 42 -613
rect 43 -619 49 -613
rect 50 -619 53 -613
rect 57 -619 60 -613
rect 64 -619 70 -613
rect 71 -619 74 -613
rect 78 -619 84 -613
rect 85 -619 88 -613
rect 92 -619 98 -613
rect 99 -619 102 -613
rect 106 -619 109 -613
rect 113 -619 119 -613
rect 120 -619 123 -613
rect 127 -619 130 -613
rect 134 -619 140 -613
rect 141 -619 144 -613
rect 148 -619 154 -613
rect 155 -619 161 -613
rect 162 -619 165 -613
rect 169 -619 175 -613
rect 176 -619 179 -613
rect 183 -619 186 -613
rect 190 -619 193 -613
rect 197 -619 203 -613
rect 204 -619 207 -613
rect 211 -619 214 -613
rect 218 -619 224 -613
rect 225 -619 228 -613
rect 232 -619 238 -613
rect 239 -619 245 -613
rect 246 -619 252 -613
rect 253 -619 259 -613
rect 260 -619 263 -613
rect 267 -619 270 -613
rect 274 -619 277 -613
rect 281 -619 284 -613
rect 288 -619 291 -613
rect 295 -619 298 -613
rect 302 -619 305 -613
rect 309 -619 312 -613
rect 316 -619 319 -613
rect 323 -619 326 -613
rect 330 -619 333 -613
rect 337 -619 340 -613
rect 344 -619 347 -613
rect 351 -619 354 -613
rect 358 -619 361 -613
rect 365 -619 371 -613
rect 372 -619 375 -613
rect 379 -619 382 -613
rect 386 -619 389 -613
rect 393 -619 399 -613
rect 400 -619 403 -613
rect 407 -619 410 -613
rect 414 -619 417 -613
rect 421 -619 424 -613
rect 428 -619 431 -613
rect 435 -619 438 -613
rect 442 -619 445 -613
rect 449 -619 452 -613
rect 456 -619 459 -613
rect 463 -619 466 -613
rect 470 -619 473 -613
rect 477 -619 480 -613
rect 484 -619 487 -613
rect 491 -619 494 -613
rect 498 -619 504 -613
rect 505 -619 508 -613
rect 512 -619 518 -613
rect 519 -619 522 -613
rect 526 -619 532 -613
rect 533 -619 536 -613
rect 540 -619 546 -613
rect 547 -619 550 -613
rect 554 -619 557 -613
rect 561 -619 564 -613
rect 568 -619 571 -613
rect 575 -619 578 -613
rect 582 -619 588 -613
rect 589 -619 592 -613
rect 596 -619 599 -613
rect 603 -619 606 -613
rect 610 -619 613 -613
rect 617 -619 620 -613
rect 624 -619 627 -613
rect 631 -619 634 -613
rect 638 -619 641 -613
rect 645 -619 648 -613
rect 652 -619 655 -613
rect 659 -619 662 -613
rect 666 -619 672 -613
rect 673 -619 676 -613
rect 680 -619 686 -613
rect 687 -619 690 -613
rect 694 -619 700 -613
rect 701 -619 707 -613
rect 708 -619 711 -613
rect 715 -619 721 -613
rect 722 -619 725 -613
rect 729 -619 735 -613
rect 736 -619 739 -613
rect 743 -619 746 -613
rect 750 -619 753 -613
rect 757 -619 760 -613
rect 764 -619 770 -613
rect 771 -619 777 -613
rect 778 -619 784 -613
rect 785 -619 788 -613
rect 792 -619 798 -613
rect 799 -619 802 -613
rect 806 -619 812 -613
rect 813 -619 816 -613
rect 820 -619 823 -613
rect 827 -619 830 -613
rect 834 -619 837 -613
rect 841 -619 844 -613
rect 848 -619 851 -613
rect 855 -619 858 -613
rect 862 -619 865 -613
rect 869 -619 872 -613
rect 876 -619 879 -613
rect 883 -619 886 -613
rect 890 -619 893 -613
rect 897 -619 903 -613
rect 904 -619 907 -613
rect 911 -619 914 -613
rect 918 -619 921 -613
rect 925 -619 928 -613
rect 932 -619 935 -613
rect 939 -619 942 -613
rect 946 -619 949 -613
rect 953 -619 956 -613
rect 960 -619 963 -613
rect 967 -619 970 -613
rect 974 -619 980 -613
rect 981 -619 984 -613
rect 988 -619 991 -613
rect 995 -619 998 -613
rect 1002 -619 1005 -613
rect 1009 -619 1012 -613
rect 1016 -619 1019 -613
rect 1023 -619 1026 -613
rect 1030 -619 1033 -613
rect 1037 -619 1040 -613
rect 1044 -619 1047 -613
rect 1051 -619 1054 -613
rect 1058 -619 1061 -613
rect 1065 -619 1068 -613
rect 1072 -619 1075 -613
rect 1079 -619 1082 -613
rect 1086 -619 1089 -613
rect 1093 -619 1096 -613
rect 1100 -619 1103 -613
rect 1107 -619 1110 -613
rect 1114 -619 1117 -613
rect 1121 -619 1124 -613
rect 1128 -619 1131 -613
rect 1135 -619 1138 -613
rect 1142 -619 1145 -613
rect 1149 -619 1152 -613
rect 1156 -619 1159 -613
rect 1163 -619 1166 -613
rect 1170 -619 1173 -613
rect 1177 -619 1180 -613
rect 1184 -619 1187 -613
rect 1191 -619 1194 -613
rect 1198 -619 1201 -613
rect 1205 -619 1208 -613
rect 1212 -619 1215 -613
rect 1219 -619 1222 -613
rect 1226 -619 1229 -613
rect 1233 -619 1236 -613
rect 1240 -619 1243 -613
rect 1247 -619 1250 -613
rect 1254 -619 1257 -613
rect 1261 -619 1264 -613
rect 1268 -619 1271 -613
rect 1275 -619 1278 -613
rect 1282 -619 1285 -613
rect 1289 -619 1292 -613
rect 1296 -619 1299 -613
rect 1303 -619 1306 -613
rect 1310 -619 1313 -613
rect 1317 -619 1320 -613
rect 1324 -619 1327 -613
rect 1331 -619 1334 -613
rect 1338 -619 1341 -613
rect 1345 -619 1348 -613
rect 1352 -619 1358 -613
rect 1359 -619 1362 -613
rect 1366 -619 1369 -613
rect 1373 -619 1376 -613
rect 1380 -619 1383 -613
rect 1387 -619 1390 -613
rect 1471 -619 1474 -613
rect 1 -742 7 -736
rect 8 -742 14 -736
rect 15 -742 21 -736
rect 22 -742 28 -736
rect 29 -742 35 -736
rect 36 -742 42 -736
rect 43 -742 46 -736
rect 50 -742 53 -736
rect 57 -742 60 -736
rect 64 -742 67 -736
rect 71 -742 74 -736
rect 78 -742 84 -736
rect 85 -742 88 -736
rect 92 -742 98 -736
rect 99 -742 102 -736
rect 106 -742 109 -736
rect 113 -742 116 -736
rect 120 -742 126 -736
rect 127 -742 130 -736
rect 134 -742 137 -736
rect 141 -742 147 -736
rect 148 -742 151 -736
rect 155 -742 158 -736
rect 162 -742 165 -736
rect 169 -742 172 -736
rect 176 -742 179 -736
rect 183 -742 189 -736
rect 190 -742 193 -736
rect 197 -742 200 -736
rect 204 -742 207 -736
rect 211 -742 214 -736
rect 218 -742 221 -736
rect 225 -742 228 -736
rect 232 -742 235 -736
rect 239 -742 242 -736
rect 246 -742 252 -736
rect 253 -742 256 -736
rect 260 -742 263 -736
rect 267 -742 270 -736
rect 274 -742 280 -736
rect 281 -742 284 -736
rect 288 -742 294 -736
rect 295 -742 298 -736
rect 302 -742 305 -736
rect 309 -742 312 -736
rect 316 -742 319 -736
rect 323 -742 326 -736
rect 330 -742 333 -736
rect 337 -742 340 -736
rect 344 -742 347 -736
rect 351 -742 354 -736
rect 358 -742 361 -736
rect 365 -742 368 -736
rect 372 -742 375 -736
rect 379 -742 382 -736
rect 386 -742 389 -736
rect 393 -742 396 -736
rect 400 -742 403 -736
rect 407 -742 410 -736
rect 414 -742 417 -736
rect 421 -742 424 -736
rect 428 -742 434 -736
rect 435 -742 441 -736
rect 442 -742 445 -736
rect 449 -742 452 -736
rect 456 -742 459 -736
rect 463 -742 466 -736
rect 470 -742 473 -736
rect 477 -742 480 -736
rect 484 -742 490 -736
rect 491 -742 494 -736
rect 498 -742 504 -736
rect 505 -742 508 -736
rect 512 -742 515 -736
rect 519 -742 522 -736
rect 526 -742 529 -736
rect 533 -742 539 -736
rect 540 -742 543 -736
rect 547 -742 550 -736
rect 554 -742 560 -736
rect 561 -742 567 -736
rect 568 -742 571 -736
rect 575 -742 581 -736
rect 582 -742 585 -736
rect 589 -742 595 -736
rect 596 -742 599 -736
rect 603 -742 609 -736
rect 610 -742 613 -736
rect 617 -742 620 -736
rect 624 -742 627 -736
rect 631 -742 637 -736
rect 638 -742 641 -736
rect 645 -742 651 -736
rect 652 -742 658 -736
rect 659 -742 662 -736
rect 666 -742 669 -736
rect 673 -742 676 -736
rect 680 -742 683 -736
rect 687 -742 690 -736
rect 694 -742 697 -736
rect 701 -742 704 -736
rect 708 -742 714 -736
rect 715 -742 718 -736
rect 722 -742 728 -736
rect 729 -742 735 -736
rect 736 -742 739 -736
rect 743 -742 746 -736
rect 750 -742 753 -736
rect 757 -742 760 -736
rect 764 -742 767 -736
rect 771 -742 774 -736
rect 778 -742 781 -736
rect 785 -742 788 -736
rect 792 -742 798 -736
rect 799 -742 802 -736
rect 806 -742 809 -736
rect 813 -742 816 -736
rect 820 -742 823 -736
rect 827 -742 833 -736
rect 834 -742 837 -736
rect 841 -742 844 -736
rect 848 -742 851 -736
rect 855 -742 861 -736
rect 862 -742 865 -736
rect 869 -742 875 -736
rect 876 -742 879 -736
rect 883 -742 889 -736
rect 890 -742 893 -736
rect 897 -742 900 -736
rect 904 -742 910 -736
rect 911 -742 917 -736
rect 918 -742 924 -736
rect 925 -742 928 -736
rect 932 -742 935 -736
rect 939 -742 942 -736
rect 946 -742 949 -736
rect 953 -742 956 -736
rect 960 -742 963 -736
rect 967 -742 970 -736
rect 974 -742 977 -736
rect 981 -742 984 -736
rect 988 -742 994 -736
rect 995 -742 998 -736
rect 1002 -742 1008 -736
rect 1009 -742 1012 -736
rect 1016 -742 1019 -736
rect 1023 -742 1026 -736
rect 1030 -742 1033 -736
rect 1037 -742 1040 -736
rect 1044 -742 1047 -736
rect 1051 -742 1054 -736
rect 1058 -742 1064 -736
rect 1065 -742 1068 -736
rect 1072 -742 1075 -736
rect 1079 -742 1082 -736
rect 1086 -742 1089 -736
rect 1093 -742 1096 -736
rect 1100 -742 1103 -736
rect 1107 -742 1110 -736
rect 1114 -742 1117 -736
rect 1121 -742 1124 -736
rect 1128 -742 1131 -736
rect 1135 -742 1138 -736
rect 1142 -742 1145 -736
rect 1149 -742 1152 -736
rect 1156 -742 1159 -736
rect 1163 -742 1166 -736
rect 1170 -742 1173 -736
rect 1177 -742 1180 -736
rect 1184 -742 1187 -736
rect 1191 -742 1194 -736
rect 1198 -742 1201 -736
rect 1205 -742 1208 -736
rect 1212 -742 1215 -736
rect 1219 -742 1222 -736
rect 1226 -742 1229 -736
rect 1233 -742 1236 -736
rect 1240 -742 1243 -736
rect 1247 -742 1250 -736
rect 1254 -742 1257 -736
rect 1261 -742 1264 -736
rect 1268 -742 1271 -736
rect 1275 -742 1278 -736
rect 1282 -742 1285 -736
rect 1289 -742 1292 -736
rect 1296 -742 1299 -736
rect 1303 -742 1306 -736
rect 1310 -742 1313 -736
rect 1317 -742 1320 -736
rect 1324 -742 1327 -736
rect 1331 -742 1334 -736
rect 1338 -742 1341 -736
rect 1345 -742 1348 -736
rect 1352 -742 1355 -736
rect 1359 -742 1362 -736
rect 1366 -742 1369 -736
rect 1373 -742 1376 -736
rect 1380 -742 1383 -736
rect 1387 -742 1390 -736
rect 1394 -742 1397 -736
rect 1401 -742 1404 -736
rect 1408 -742 1411 -736
rect 1415 -742 1418 -736
rect 1422 -742 1428 -736
rect 1429 -742 1432 -736
rect 1499 -742 1502 -736
rect 1520 -742 1523 -736
rect 1569 -742 1572 -736
rect 1632 -742 1635 -736
rect 1 -881 7 -875
rect 8 -881 14 -875
rect 15 -881 21 -875
rect 22 -881 25 -875
rect 29 -881 35 -875
rect 36 -881 39 -875
rect 43 -881 46 -875
rect 50 -881 56 -875
rect 57 -881 60 -875
rect 64 -881 67 -875
rect 71 -881 74 -875
rect 78 -881 81 -875
rect 85 -881 91 -875
rect 92 -881 95 -875
rect 99 -881 105 -875
rect 106 -881 112 -875
rect 113 -881 116 -875
rect 120 -881 123 -875
rect 127 -881 130 -875
rect 134 -881 140 -875
rect 141 -881 144 -875
rect 148 -881 151 -875
rect 155 -881 158 -875
rect 162 -881 168 -875
rect 169 -881 172 -875
rect 176 -881 179 -875
rect 183 -881 186 -875
rect 190 -881 193 -875
rect 197 -881 200 -875
rect 204 -881 210 -875
rect 211 -881 214 -875
rect 218 -881 221 -875
rect 225 -881 231 -875
rect 232 -881 238 -875
rect 239 -881 242 -875
rect 246 -881 252 -875
rect 253 -881 256 -875
rect 260 -881 263 -875
rect 267 -881 270 -875
rect 274 -881 277 -875
rect 281 -881 284 -875
rect 288 -881 291 -875
rect 295 -881 301 -875
rect 302 -881 305 -875
rect 309 -881 312 -875
rect 316 -881 322 -875
rect 323 -881 326 -875
rect 330 -881 333 -875
rect 337 -881 340 -875
rect 344 -881 347 -875
rect 351 -881 354 -875
rect 358 -881 361 -875
rect 365 -881 368 -875
rect 372 -881 375 -875
rect 379 -881 382 -875
rect 386 -881 389 -875
rect 393 -881 396 -875
rect 400 -881 403 -875
rect 407 -881 410 -875
rect 414 -881 417 -875
rect 421 -881 424 -875
rect 428 -881 431 -875
rect 435 -881 438 -875
rect 442 -881 445 -875
rect 449 -881 452 -875
rect 456 -881 459 -875
rect 463 -881 469 -875
rect 470 -881 473 -875
rect 477 -881 483 -875
rect 484 -881 487 -875
rect 491 -881 494 -875
rect 498 -881 501 -875
rect 505 -881 508 -875
rect 512 -881 515 -875
rect 519 -881 522 -875
rect 526 -881 529 -875
rect 533 -881 536 -875
rect 540 -881 543 -875
rect 547 -881 550 -875
rect 554 -881 557 -875
rect 561 -881 567 -875
rect 568 -881 571 -875
rect 575 -881 581 -875
rect 582 -881 588 -875
rect 589 -881 592 -875
rect 596 -881 599 -875
rect 603 -881 606 -875
rect 610 -881 616 -875
rect 617 -881 620 -875
rect 624 -881 630 -875
rect 631 -881 634 -875
rect 638 -881 644 -875
rect 645 -881 648 -875
rect 652 -881 658 -875
rect 659 -881 665 -875
rect 666 -881 669 -875
rect 673 -881 676 -875
rect 680 -881 683 -875
rect 687 -881 693 -875
rect 694 -881 697 -875
rect 701 -881 707 -875
rect 708 -881 711 -875
rect 715 -881 718 -875
rect 722 -881 725 -875
rect 729 -881 732 -875
rect 736 -881 742 -875
rect 743 -881 746 -875
rect 750 -881 753 -875
rect 757 -881 763 -875
rect 764 -881 767 -875
rect 771 -881 774 -875
rect 778 -881 784 -875
rect 785 -881 791 -875
rect 792 -881 798 -875
rect 799 -881 802 -875
rect 806 -881 809 -875
rect 813 -881 816 -875
rect 820 -881 823 -875
rect 827 -881 833 -875
rect 834 -881 837 -875
rect 841 -881 844 -875
rect 848 -881 851 -875
rect 855 -881 858 -875
rect 862 -881 865 -875
rect 869 -881 872 -875
rect 876 -881 882 -875
rect 883 -881 886 -875
rect 890 -881 893 -875
rect 897 -881 900 -875
rect 904 -881 910 -875
rect 911 -881 914 -875
rect 918 -881 921 -875
rect 925 -881 931 -875
rect 932 -881 935 -875
rect 939 -881 942 -875
rect 946 -881 949 -875
rect 953 -881 956 -875
rect 960 -881 966 -875
rect 967 -881 970 -875
rect 974 -881 977 -875
rect 981 -881 984 -875
rect 988 -881 991 -875
rect 995 -881 998 -875
rect 1002 -881 1005 -875
rect 1009 -881 1012 -875
rect 1016 -881 1019 -875
rect 1023 -881 1026 -875
rect 1030 -881 1033 -875
rect 1037 -881 1040 -875
rect 1044 -881 1047 -875
rect 1051 -881 1054 -875
rect 1058 -881 1064 -875
rect 1065 -881 1068 -875
rect 1072 -881 1075 -875
rect 1079 -881 1082 -875
rect 1086 -881 1089 -875
rect 1093 -881 1096 -875
rect 1100 -881 1103 -875
rect 1107 -881 1110 -875
rect 1114 -881 1117 -875
rect 1121 -881 1124 -875
rect 1128 -881 1131 -875
rect 1135 -881 1138 -875
rect 1142 -881 1145 -875
rect 1149 -881 1152 -875
rect 1156 -881 1159 -875
rect 1163 -881 1166 -875
rect 1170 -881 1173 -875
rect 1177 -881 1180 -875
rect 1184 -881 1187 -875
rect 1191 -881 1194 -875
rect 1198 -881 1201 -875
rect 1205 -881 1208 -875
rect 1212 -881 1215 -875
rect 1219 -881 1222 -875
rect 1226 -881 1229 -875
rect 1233 -881 1236 -875
rect 1240 -881 1243 -875
rect 1247 -881 1250 -875
rect 1254 -881 1257 -875
rect 1261 -881 1264 -875
rect 1268 -881 1271 -875
rect 1275 -881 1278 -875
rect 1282 -881 1285 -875
rect 1289 -881 1292 -875
rect 1296 -881 1299 -875
rect 1303 -881 1306 -875
rect 1310 -881 1313 -875
rect 1317 -881 1320 -875
rect 1324 -881 1327 -875
rect 1331 -881 1334 -875
rect 1338 -881 1341 -875
rect 1345 -881 1348 -875
rect 1352 -881 1355 -875
rect 1359 -881 1362 -875
rect 1366 -881 1369 -875
rect 1373 -881 1376 -875
rect 1380 -881 1383 -875
rect 1387 -881 1390 -875
rect 1394 -881 1397 -875
rect 1401 -881 1404 -875
rect 1408 -881 1411 -875
rect 1415 -881 1418 -875
rect 1422 -881 1425 -875
rect 1429 -881 1432 -875
rect 1436 -881 1439 -875
rect 1443 -881 1446 -875
rect 1450 -881 1453 -875
rect 1457 -881 1460 -875
rect 1464 -881 1467 -875
rect 1471 -881 1474 -875
rect 1478 -881 1481 -875
rect 1485 -881 1488 -875
rect 1492 -881 1495 -875
rect 1499 -881 1502 -875
rect 1506 -881 1509 -875
rect 1513 -881 1516 -875
rect 1520 -881 1523 -875
rect 1527 -881 1530 -875
rect 1534 -881 1537 -875
rect 1541 -881 1544 -875
rect 1548 -881 1551 -875
rect 1555 -881 1558 -875
rect 1562 -881 1565 -875
rect 1569 -881 1572 -875
rect 1576 -881 1579 -875
rect 1583 -881 1586 -875
rect 1590 -881 1593 -875
rect 1597 -881 1603 -875
rect 1604 -881 1610 -875
rect 1611 -881 1614 -875
rect 1618 -881 1621 -875
rect 1625 -881 1628 -875
rect 1632 -881 1635 -875
rect 1695 -881 1698 -875
rect 1 -1042 7 -1036
rect 8 -1042 14 -1036
rect 15 -1042 21 -1036
rect 22 -1042 28 -1036
rect 29 -1042 32 -1036
rect 36 -1042 39 -1036
rect 43 -1042 49 -1036
rect 50 -1042 56 -1036
rect 57 -1042 60 -1036
rect 64 -1042 67 -1036
rect 71 -1042 74 -1036
rect 78 -1042 81 -1036
rect 85 -1042 91 -1036
rect 92 -1042 95 -1036
rect 99 -1042 102 -1036
rect 106 -1042 112 -1036
rect 113 -1042 116 -1036
rect 120 -1042 126 -1036
rect 127 -1042 130 -1036
rect 134 -1042 137 -1036
rect 141 -1042 144 -1036
rect 148 -1042 151 -1036
rect 155 -1042 158 -1036
rect 162 -1042 165 -1036
rect 169 -1042 172 -1036
rect 176 -1042 179 -1036
rect 183 -1042 186 -1036
rect 190 -1042 193 -1036
rect 197 -1042 203 -1036
rect 204 -1042 207 -1036
rect 211 -1042 214 -1036
rect 218 -1042 224 -1036
rect 225 -1042 228 -1036
rect 232 -1042 235 -1036
rect 239 -1042 242 -1036
rect 246 -1042 249 -1036
rect 253 -1042 256 -1036
rect 260 -1042 263 -1036
rect 267 -1042 270 -1036
rect 274 -1042 277 -1036
rect 281 -1042 284 -1036
rect 288 -1042 294 -1036
rect 295 -1042 298 -1036
rect 302 -1042 305 -1036
rect 309 -1042 315 -1036
rect 316 -1042 319 -1036
rect 323 -1042 326 -1036
rect 330 -1042 333 -1036
rect 337 -1042 340 -1036
rect 344 -1042 347 -1036
rect 351 -1042 354 -1036
rect 358 -1042 361 -1036
rect 365 -1042 368 -1036
rect 372 -1042 375 -1036
rect 379 -1042 382 -1036
rect 386 -1042 389 -1036
rect 393 -1042 396 -1036
rect 400 -1042 403 -1036
rect 407 -1042 410 -1036
rect 414 -1042 417 -1036
rect 421 -1042 424 -1036
rect 428 -1042 431 -1036
rect 435 -1042 438 -1036
rect 442 -1042 445 -1036
rect 449 -1042 452 -1036
rect 456 -1042 459 -1036
rect 463 -1042 469 -1036
rect 470 -1042 476 -1036
rect 477 -1042 480 -1036
rect 484 -1042 487 -1036
rect 491 -1042 494 -1036
rect 498 -1042 501 -1036
rect 505 -1042 508 -1036
rect 512 -1042 515 -1036
rect 519 -1042 522 -1036
rect 526 -1042 529 -1036
rect 533 -1042 539 -1036
rect 540 -1042 543 -1036
rect 547 -1042 553 -1036
rect 554 -1042 557 -1036
rect 561 -1042 564 -1036
rect 568 -1042 571 -1036
rect 575 -1042 578 -1036
rect 582 -1042 585 -1036
rect 589 -1042 595 -1036
rect 596 -1042 602 -1036
rect 603 -1042 609 -1036
rect 610 -1042 613 -1036
rect 617 -1042 623 -1036
rect 624 -1042 630 -1036
rect 631 -1042 637 -1036
rect 638 -1042 641 -1036
rect 645 -1042 648 -1036
rect 652 -1042 655 -1036
rect 659 -1042 662 -1036
rect 666 -1042 669 -1036
rect 673 -1042 676 -1036
rect 680 -1042 686 -1036
rect 687 -1042 690 -1036
rect 694 -1042 697 -1036
rect 701 -1042 704 -1036
rect 708 -1042 711 -1036
rect 715 -1042 718 -1036
rect 722 -1042 728 -1036
rect 729 -1042 735 -1036
rect 736 -1042 739 -1036
rect 743 -1042 746 -1036
rect 750 -1042 753 -1036
rect 757 -1042 763 -1036
rect 764 -1042 770 -1036
rect 771 -1042 774 -1036
rect 778 -1042 781 -1036
rect 785 -1042 788 -1036
rect 792 -1042 798 -1036
rect 799 -1042 802 -1036
rect 806 -1042 812 -1036
rect 813 -1042 816 -1036
rect 820 -1042 823 -1036
rect 827 -1042 833 -1036
rect 834 -1042 837 -1036
rect 841 -1042 847 -1036
rect 848 -1042 851 -1036
rect 855 -1042 861 -1036
rect 862 -1042 865 -1036
rect 869 -1042 875 -1036
rect 876 -1042 882 -1036
rect 883 -1042 886 -1036
rect 890 -1042 893 -1036
rect 897 -1042 903 -1036
rect 904 -1042 907 -1036
rect 911 -1042 914 -1036
rect 918 -1042 921 -1036
rect 925 -1042 928 -1036
rect 932 -1042 935 -1036
rect 939 -1042 942 -1036
rect 946 -1042 949 -1036
rect 953 -1042 959 -1036
rect 960 -1042 963 -1036
rect 967 -1042 970 -1036
rect 974 -1042 980 -1036
rect 981 -1042 984 -1036
rect 988 -1042 994 -1036
rect 995 -1042 998 -1036
rect 1002 -1042 1005 -1036
rect 1009 -1042 1012 -1036
rect 1016 -1042 1019 -1036
rect 1023 -1042 1026 -1036
rect 1030 -1042 1033 -1036
rect 1037 -1042 1040 -1036
rect 1044 -1042 1047 -1036
rect 1051 -1042 1054 -1036
rect 1058 -1042 1064 -1036
rect 1065 -1042 1071 -1036
rect 1072 -1042 1075 -1036
rect 1079 -1042 1082 -1036
rect 1086 -1042 1089 -1036
rect 1093 -1042 1096 -1036
rect 1100 -1042 1103 -1036
rect 1107 -1042 1110 -1036
rect 1114 -1042 1117 -1036
rect 1121 -1042 1124 -1036
rect 1128 -1042 1131 -1036
rect 1135 -1042 1138 -1036
rect 1142 -1042 1145 -1036
rect 1149 -1042 1152 -1036
rect 1156 -1042 1159 -1036
rect 1163 -1042 1166 -1036
rect 1170 -1042 1173 -1036
rect 1177 -1042 1180 -1036
rect 1184 -1042 1187 -1036
rect 1191 -1042 1194 -1036
rect 1198 -1042 1201 -1036
rect 1205 -1042 1208 -1036
rect 1212 -1042 1215 -1036
rect 1219 -1042 1222 -1036
rect 1226 -1042 1229 -1036
rect 1233 -1042 1236 -1036
rect 1240 -1042 1243 -1036
rect 1247 -1042 1250 -1036
rect 1254 -1042 1257 -1036
rect 1261 -1042 1264 -1036
rect 1268 -1042 1271 -1036
rect 1275 -1042 1278 -1036
rect 1282 -1042 1285 -1036
rect 1289 -1042 1292 -1036
rect 1296 -1042 1299 -1036
rect 1303 -1042 1306 -1036
rect 1310 -1042 1313 -1036
rect 1317 -1042 1320 -1036
rect 1324 -1042 1327 -1036
rect 1331 -1042 1334 -1036
rect 1338 -1042 1341 -1036
rect 1345 -1042 1348 -1036
rect 1352 -1042 1355 -1036
rect 1359 -1042 1362 -1036
rect 1366 -1042 1369 -1036
rect 1373 -1042 1376 -1036
rect 1380 -1042 1383 -1036
rect 1387 -1042 1390 -1036
rect 1394 -1042 1397 -1036
rect 1401 -1042 1404 -1036
rect 1408 -1042 1411 -1036
rect 1415 -1042 1418 -1036
rect 1422 -1042 1425 -1036
rect 1429 -1042 1432 -1036
rect 1436 -1042 1439 -1036
rect 1443 -1042 1446 -1036
rect 1450 -1042 1453 -1036
rect 1457 -1042 1460 -1036
rect 1464 -1042 1467 -1036
rect 1471 -1042 1474 -1036
rect 1478 -1042 1481 -1036
rect 1485 -1042 1488 -1036
rect 1492 -1042 1495 -1036
rect 1499 -1042 1502 -1036
rect 1506 -1042 1509 -1036
rect 1513 -1042 1516 -1036
rect 1520 -1042 1523 -1036
rect 1527 -1042 1530 -1036
rect 1534 -1042 1537 -1036
rect 1541 -1042 1544 -1036
rect 1548 -1042 1551 -1036
rect 1555 -1042 1558 -1036
rect 1562 -1042 1565 -1036
rect 1569 -1042 1572 -1036
rect 1576 -1042 1579 -1036
rect 1583 -1042 1586 -1036
rect 1590 -1042 1593 -1036
rect 1597 -1042 1600 -1036
rect 1604 -1042 1607 -1036
rect 1611 -1042 1614 -1036
rect 1618 -1042 1621 -1036
rect 1625 -1042 1628 -1036
rect 1632 -1042 1635 -1036
rect 1639 -1042 1642 -1036
rect 1646 -1042 1649 -1036
rect 1653 -1042 1656 -1036
rect 1660 -1042 1663 -1036
rect 1667 -1042 1670 -1036
rect 1674 -1042 1677 -1036
rect 1681 -1042 1684 -1036
rect 1688 -1042 1691 -1036
rect 1695 -1042 1698 -1036
rect 1702 -1042 1705 -1036
rect 1709 -1042 1712 -1036
rect 1716 -1042 1719 -1036
rect 1723 -1042 1726 -1036
rect 1 -1193 7 -1187
rect 8 -1193 14 -1187
rect 15 -1193 21 -1187
rect 22 -1193 28 -1187
rect 29 -1193 32 -1187
rect 36 -1193 39 -1187
rect 43 -1193 46 -1187
rect 50 -1193 53 -1187
rect 57 -1193 60 -1187
rect 64 -1193 67 -1187
rect 71 -1193 77 -1187
rect 78 -1193 84 -1187
rect 85 -1193 91 -1187
rect 92 -1193 95 -1187
rect 99 -1193 105 -1187
rect 106 -1193 109 -1187
rect 113 -1193 116 -1187
rect 120 -1193 126 -1187
rect 127 -1193 130 -1187
rect 134 -1193 137 -1187
rect 141 -1193 144 -1187
rect 148 -1193 154 -1187
rect 155 -1193 158 -1187
rect 162 -1193 168 -1187
rect 169 -1193 172 -1187
rect 176 -1193 179 -1187
rect 183 -1193 189 -1187
rect 190 -1193 193 -1187
rect 197 -1193 203 -1187
rect 204 -1193 210 -1187
rect 211 -1193 214 -1187
rect 218 -1193 221 -1187
rect 225 -1193 228 -1187
rect 232 -1193 238 -1187
rect 239 -1193 242 -1187
rect 246 -1193 249 -1187
rect 253 -1193 259 -1187
rect 260 -1193 263 -1187
rect 267 -1193 270 -1187
rect 274 -1193 280 -1187
rect 281 -1193 284 -1187
rect 288 -1193 291 -1187
rect 295 -1193 298 -1187
rect 302 -1193 305 -1187
rect 309 -1193 312 -1187
rect 316 -1193 319 -1187
rect 323 -1193 326 -1187
rect 330 -1193 333 -1187
rect 337 -1193 340 -1187
rect 344 -1193 347 -1187
rect 351 -1193 354 -1187
rect 358 -1193 361 -1187
rect 365 -1193 368 -1187
rect 372 -1193 375 -1187
rect 379 -1193 382 -1187
rect 386 -1193 389 -1187
rect 393 -1193 396 -1187
rect 400 -1193 403 -1187
rect 407 -1193 410 -1187
rect 414 -1193 417 -1187
rect 421 -1193 424 -1187
rect 428 -1193 431 -1187
rect 435 -1193 438 -1187
rect 442 -1193 445 -1187
rect 449 -1193 452 -1187
rect 456 -1193 459 -1187
rect 463 -1193 469 -1187
rect 470 -1193 473 -1187
rect 477 -1193 480 -1187
rect 484 -1193 490 -1187
rect 491 -1193 494 -1187
rect 498 -1193 501 -1187
rect 505 -1193 511 -1187
rect 512 -1193 518 -1187
rect 519 -1193 522 -1187
rect 526 -1193 529 -1187
rect 533 -1193 536 -1187
rect 540 -1193 546 -1187
rect 547 -1193 550 -1187
rect 554 -1193 557 -1187
rect 561 -1193 564 -1187
rect 568 -1193 571 -1187
rect 575 -1193 581 -1187
rect 582 -1193 585 -1187
rect 589 -1193 592 -1187
rect 596 -1193 602 -1187
rect 603 -1193 606 -1187
rect 610 -1193 616 -1187
rect 617 -1193 623 -1187
rect 624 -1193 627 -1187
rect 631 -1193 634 -1187
rect 638 -1193 641 -1187
rect 645 -1193 648 -1187
rect 652 -1193 655 -1187
rect 659 -1193 665 -1187
rect 666 -1193 669 -1187
rect 673 -1193 676 -1187
rect 680 -1193 683 -1187
rect 687 -1193 690 -1187
rect 694 -1193 697 -1187
rect 701 -1193 704 -1187
rect 708 -1193 711 -1187
rect 715 -1193 721 -1187
rect 722 -1193 728 -1187
rect 729 -1193 732 -1187
rect 736 -1193 739 -1187
rect 743 -1193 749 -1187
rect 750 -1193 756 -1187
rect 757 -1193 760 -1187
rect 764 -1193 767 -1187
rect 771 -1193 774 -1187
rect 778 -1193 781 -1187
rect 785 -1193 788 -1187
rect 792 -1193 795 -1187
rect 799 -1193 802 -1187
rect 806 -1193 809 -1187
rect 813 -1193 816 -1187
rect 820 -1193 823 -1187
rect 827 -1193 833 -1187
rect 834 -1193 837 -1187
rect 841 -1193 844 -1187
rect 848 -1193 851 -1187
rect 855 -1193 858 -1187
rect 862 -1193 865 -1187
rect 869 -1193 875 -1187
rect 876 -1193 879 -1187
rect 883 -1193 886 -1187
rect 890 -1193 896 -1187
rect 897 -1193 903 -1187
rect 904 -1193 907 -1187
rect 911 -1193 914 -1187
rect 918 -1193 921 -1187
rect 925 -1193 928 -1187
rect 932 -1193 935 -1187
rect 939 -1193 942 -1187
rect 946 -1193 949 -1187
rect 953 -1193 959 -1187
rect 960 -1193 963 -1187
rect 967 -1193 973 -1187
rect 974 -1193 977 -1187
rect 981 -1193 984 -1187
rect 988 -1193 994 -1187
rect 995 -1193 998 -1187
rect 1002 -1193 1005 -1187
rect 1009 -1193 1012 -1187
rect 1016 -1193 1019 -1187
rect 1023 -1193 1026 -1187
rect 1030 -1193 1033 -1187
rect 1037 -1193 1040 -1187
rect 1044 -1193 1050 -1187
rect 1051 -1193 1054 -1187
rect 1058 -1193 1061 -1187
rect 1065 -1193 1068 -1187
rect 1072 -1193 1075 -1187
rect 1079 -1193 1082 -1187
rect 1086 -1193 1089 -1187
rect 1093 -1193 1096 -1187
rect 1100 -1193 1103 -1187
rect 1107 -1193 1110 -1187
rect 1114 -1193 1117 -1187
rect 1121 -1193 1124 -1187
rect 1128 -1193 1131 -1187
rect 1135 -1193 1138 -1187
rect 1142 -1193 1145 -1187
rect 1149 -1193 1152 -1187
rect 1156 -1193 1159 -1187
rect 1163 -1193 1166 -1187
rect 1170 -1193 1173 -1187
rect 1177 -1193 1180 -1187
rect 1184 -1193 1187 -1187
rect 1191 -1193 1194 -1187
rect 1198 -1193 1201 -1187
rect 1205 -1193 1208 -1187
rect 1212 -1193 1215 -1187
rect 1219 -1193 1222 -1187
rect 1226 -1193 1229 -1187
rect 1233 -1193 1236 -1187
rect 1240 -1193 1243 -1187
rect 1247 -1193 1250 -1187
rect 1254 -1193 1257 -1187
rect 1261 -1193 1264 -1187
rect 1268 -1193 1271 -1187
rect 1275 -1193 1278 -1187
rect 1282 -1193 1285 -1187
rect 1289 -1193 1292 -1187
rect 1296 -1193 1299 -1187
rect 1303 -1193 1306 -1187
rect 1310 -1193 1313 -1187
rect 1317 -1193 1320 -1187
rect 1324 -1193 1327 -1187
rect 1331 -1193 1334 -1187
rect 1338 -1193 1341 -1187
rect 1345 -1193 1348 -1187
rect 1352 -1193 1355 -1187
rect 1359 -1193 1362 -1187
rect 1366 -1193 1369 -1187
rect 1373 -1193 1376 -1187
rect 1380 -1193 1383 -1187
rect 1387 -1193 1390 -1187
rect 1394 -1193 1397 -1187
rect 1401 -1193 1404 -1187
rect 1408 -1193 1411 -1187
rect 1415 -1193 1418 -1187
rect 1422 -1193 1425 -1187
rect 1429 -1193 1432 -1187
rect 1436 -1193 1439 -1187
rect 1443 -1193 1446 -1187
rect 1450 -1193 1453 -1187
rect 1457 -1193 1460 -1187
rect 1464 -1193 1467 -1187
rect 1471 -1193 1474 -1187
rect 1478 -1193 1481 -1187
rect 1485 -1193 1488 -1187
rect 1492 -1193 1495 -1187
rect 1499 -1193 1502 -1187
rect 1506 -1193 1509 -1187
rect 1513 -1193 1516 -1187
rect 1520 -1193 1523 -1187
rect 1527 -1193 1530 -1187
rect 1534 -1193 1537 -1187
rect 1541 -1193 1544 -1187
rect 1548 -1193 1551 -1187
rect 1555 -1193 1558 -1187
rect 1562 -1193 1565 -1187
rect 1569 -1193 1572 -1187
rect 1576 -1193 1579 -1187
rect 1583 -1193 1586 -1187
rect 1590 -1193 1593 -1187
rect 1597 -1193 1600 -1187
rect 1604 -1193 1607 -1187
rect 1611 -1193 1614 -1187
rect 1618 -1193 1621 -1187
rect 1625 -1193 1628 -1187
rect 1632 -1193 1635 -1187
rect 1639 -1193 1642 -1187
rect 1646 -1193 1652 -1187
rect 1653 -1193 1656 -1187
rect 1660 -1193 1666 -1187
rect 1674 -1193 1677 -1187
rect 1723 -1193 1726 -1187
rect 1730 -1193 1733 -1187
rect 1 -1324 7 -1318
rect 8 -1324 14 -1318
rect 15 -1324 21 -1318
rect 22 -1324 25 -1318
rect 29 -1324 32 -1318
rect 36 -1324 39 -1318
rect 43 -1324 46 -1318
rect 50 -1324 53 -1318
rect 57 -1324 60 -1318
rect 64 -1324 67 -1318
rect 71 -1324 77 -1318
rect 78 -1324 84 -1318
rect 85 -1324 88 -1318
rect 92 -1324 98 -1318
rect 99 -1324 102 -1318
rect 106 -1324 109 -1318
rect 113 -1324 116 -1318
rect 120 -1324 126 -1318
rect 127 -1324 130 -1318
rect 134 -1324 137 -1318
rect 141 -1324 147 -1318
rect 148 -1324 151 -1318
rect 155 -1324 158 -1318
rect 162 -1324 168 -1318
rect 169 -1324 172 -1318
rect 176 -1324 179 -1318
rect 183 -1324 186 -1318
rect 190 -1324 193 -1318
rect 197 -1324 200 -1318
rect 204 -1324 207 -1318
rect 211 -1324 214 -1318
rect 218 -1324 221 -1318
rect 225 -1324 228 -1318
rect 232 -1324 238 -1318
rect 239 -1324 242 -1318
rect 246 -1324 252 -1318
rect 253 -1324 256 -1318
rect 260 -1324 263 -1318
rect 267 -1324 270 -1318
rect 274 -1324 280 -1318
rect 281 -1324 284 -1318
rect 288 -1324 291 -1318
rect 295 -1324 298 -1318
rect 302 -1324 305 -1318
rect 309 -1324 312 -1318
rect 316 -1324 319 -1318
rect 323 -1324 326 -1318
rect 330 -1324 333 -1318
rect 337 -1324 340 -1318
rect 344 -1324 347 -1318
rect 351 -1324 354 -1318
rect 358 -1324 361 -1318
rect 365 -1324 368 -1318
rect 372 -1324 375 -1318
rect 379 -1324 382 -1318
rect 386 -1324 389 -1318
rect 393 -1324 396 -1318
rect 400 -1324 403 -1318
rect 407 -1324 410 -1318
rect 414 -1324 417 -1318
rect 421 -1324 427 -1318
rect 428 -1324 431 -1318
rect 435 -1324 438 -1318
rect 442 -1324 445 -1318
rect 449 -1324 452 -1318
rect 456 -1324 462 -1318
rect 463 -1324 466 -1318
rect 470 -1324 473 -1318
rect 477 -1324 483 -1318
rect 484 -1324 487 -1318
rect 491 -1324 494 -1318
rect 498 -1324 501 -1318
rect 505 -1324 511 -1318
rect 512 -1324 518 -1318
rect 519 -1324 522 -1318
rect 526 -1324 532 -1318
rect 533 -1324 536 -1318
rect 540 -1324 543 -1318
rect 547 -1324 550 -1318
rect 554 -1324 557 -1318
rect 561 -1324 564 -1318
rect 568 -1324 571 -1318
rect 575 -1324 581 -1318
rect 582 -1324 585 -1318
rect 589 -1324 595 -1318
rect 596 -1324 599 -1318
rect 603 -1324 606 -1318
rect 610 -1324 616 -1318
rect 617 -1324 620 -1318
rect 624 -1324 630 -1318
rect 631 -1324 634 -1318
rect 638 -1324 641 -1318
rect 645 -1324 648 -1318
rect 652 -1324 655 -1318
rect 659 -1324 665 -1318
rect 666 -1324 669 -1318
rect 673 -1324 676 -1318
rect 680 -1324 683 -1318
rect 687 -1324 693 -1318
rect 694 -1324 697 -1318
rect 701 -1324 704 -1318
rect 708 -1324 711 -1318
rect 715 -1324 718 -1318
rect 722 -1324 725 -1318
rect 729 -1324 732 -1318
rect 736 -1324 739 -1318
rect 743 -1324 746 -1318
rect 750 -1324 753 -1318
rect 757 -1324 760 -1318
rect 764 -1324 770 -1318
rect 771 -1324 774 -1318
rect 778 -1324 781 -1318
rect 785 -1324 791 -1318
rect 792 -1324 798 -1318
rect 799 -1324 802 -1318
rect 806 -1324 812 -1318
rect 813 -1324 819 -1318
rect 820 -1324 826 -1318
rect 827 -1324 833 -1318
rect 834 -1324 837 -1318
rect 841 -1324 844 -1318
rect 848 -1324 851 -1318
rect 855 -1324 858 -1318
rect 862 -1324 865 -1318
rect 869 -1324 872 -1318
rect 876 -1324 879 -1318
rect 883 -1324 886 -1318
rect 890 -1324 893 -1318
rect 897 -1324 900 -1318
rect 904 -1324 907 -1318
rect 911 -1324 914 -1318
rect 918 -1324 921 -1318
rect 925 -1324 928 -1318
rect 932 -1324 938 -1318
rect 939 -1324 942 -1318
rect 946 -1324 952 -1318
rect 953 -1324 956 -1318
rect 960 -1324 963 -1318
rect 967 -1324 970 -1318
rect 974 -1324 980 -1318
rect 981 -1324 987 -1318
rect 988 -1324 991 -1318
rect 995 -1324 998 -1318
rect 1002 -1324 1005 -1318
rect 1009 -1324 1015 -1318
rect 1016 -1324 1019 -1318
rect 1023 -1324 1026 -1318
rect 1030 -1324 1033 -1318
rect 1037 -1324 1040 -1318
rect 1044 -1324 1047 -1318
rect 1051 -1324 1057 -1318
rect 1058 -1324 1061 -1318
rect 1065 -1324 1068 -1318
rect 1072 -1324 1075 -1318
rect 1079 -1324 1082 -1318
rect 1086 -1324 1089 -1318
rect 1093 -1324 1096 -1318
rect 1100 -1324 1103 -1318
rect 1107 -1324 1110 -1318
rect 1114 -1324 1117 -1318
rect 1121 -1324 1124 -1318
rect 1128 -1324 1131 -1318
rect 1135 -1324 1138 -1318
rect 1142 -1324 1145 -1318
rect 1149 -1324 1152 -1318
rect 1156 -1324 1159 -1318
rect 1163 -1324 1166 -1318
rect 1170 -1324 1173 -1318
rect 1177 -1324 1180 -1318
rect 1184 -1324 1187 -1318
rect 1191 -1324 1194 -1318
rect 1198 -1324 1201 -1318
rect 1205 -1324 1208 -1318
rect 1212 -1324 1215 -1318
rect 1219 -1324 1222 -1318
rect 1226 -1324 1229 -1318
rect 1233 -1324 1236 -1318
rect 1240 -1324 1243 -1318
rect 1247 -1324 1250 -1318
rect 1254 -1324 1257 -1318
rect 1261 -1324 1264 -1318
rect 1268 -1324 1271 -1318
rect 1275 -1324 1278 -1318
rect 1282 -1324 1285 -1318
rect 1289 -1324 1292 -1318
rect 1296 -1324 1299 -1318
rect 1303 -1324 1306 -1318
rect 1310 -1324 1313 -1318
rect 1317 -1324 1320 -1318
rect 1324 -1324 1327 -1318
rect 1331 -1324 1334 -1318
rect 1338 -1324 1341 -1318
rect 1345 -1324 1348 -1318
rect 1352 -1324 1358 -1318
rect 1359 -1324 1362 -1318
rect 1366 -1324 1369 -1318
rect 1373 -1324 1376 -1318
rect 1380 -1324 1383 -1318
rect 1387 -1324 1390 -1318
rect 1394 -1324 1397 -1318
rect 1401 -1324 1404 -1318
rect 1408 -1324 1411 -1318
rect 1415 -1324 1418 -1318
rect 1422 -1324 1425 -1318
rect 1429 -1324 1432 -1318
rect 1436 -1324 1439 -1318
rect 1443 -1324 1446 -1318
rect 1450 -1324 1453 -1318
rect 1457 -1324 1460 -1318
rect 1464 -1324 1467 -1318
rect 1471 -1324 1474 -1318
rect 1478 -1324 1481 -1318
rect 1485 -1324 1488 -1318
rect 1492 -1324 1495 -1318
rect 1499 -1324 1502 -1318
rect 1506 -1324 1509 -1318
rect 1513 -1324 1516 -1318
rect 1520 -1324 1523 -1318
rect 1527 -1324 1530 -1318
rect 1534 -1324 1537 -1318
rect 1541 -1324 1544 -1318
rect 1548 -1324 1551 -1318
rect 1555 -1324 1558 -1318
rect 1562 -1324 1565 -1318
rect 1569 -1324 1572 -1318
rect 1576 -1324 1579 -1318
rect 1583 -1324 1586 -1318
rect 1590 -1324 1593 -1318
rect 1597 -1324 1600 -1318
rect 1604 -1324 1607 -1318
rect 1611 -1324 1614 -1318
rect 1618 -1324 1621 -1318
rect 1625 -1324 1628 -1318
rect 1632 -1324 1635 -1318
rect 1639 -1324 1642 -1318
rect 1646 -1324 1649 -1318
rect 1653 -1324 1656 -1318
rect 1660 -1324 1663 -1318
rect 1667 -1324 1670 -1318
rect 1674 -1324 1677 -1318
rect 1681 -1324 1684 -1318
rect 1688 -1324 1691 -1318
rect 1695 -1324 1698 -1318
rect 1702 -1324 1708 -1318
rect 1709 -1324 1715 -1318
rect 1716 -1324 1719 -1318
rect 1723 -1324 1726 -1318
rect 1730 -1324 1736 -1318
rect 1737 -1324 1740 -1318
rect 1 -1479 7 -1473
rect 8 -1479 14 -1473
rect 15 -1479 18 -1473
rect 22 -1479 28 -1473
rect 29 -1479 32 -1473
rect 36 -1479 39 -1473
rect 43 -1479 46 -1473
rect 50 -1479 53 -1473
rect 57 -1479 63 -1473
rect 64 -1479 67 -1473
rect 71 -1479 77 -1473
rect 78 -1479 84 -1473
rect 85 -1479 88 -1473
rect 92 -1479 98 -1473
rect 99 -1479 102 -1473
rect 106 -1479 112 -1473
rect 113 -1479 119 -1473
rect 120 -1479 123 -1473
rect 127 -1479 130 -1473
rect 134 -1479 137 -1473
rect 141 -1479 144 -1473
rect 148 -1479 151 -1473
rect 155 -1479 161 -1473
rect 162 -1479 165 -1473
rect 169 -1479 172 -1473
rect 176 -1479 179 -1473
rect 183 -1479 186 -1473
rect 190 -1479 193 -1473
rect 197 -1479 200 -1473
rect 204 -1479 207 -1473
rect 211 -1479 214 -1473
rect 218 -1479 224 -1473
rect 225 -1479 231 -1473
rect 232 -1479 235 -1473
rect 239 -1479 242 -1473
rect 246 -1479 249 -1473
rect 253 -1479 256 -1473
rect 260 -1479 266 -1473
rect 267 -1479 270 -1473
rect 274 -1479 277 -1473
rect 281 -1479 284 -1473
rect 288 -1479 291 -1473
rect 295 -1479 301 -1473
rect 302 -1479 305 -1473
rect 309 -1479 312 -1473
rect 316 -1479 319 -1473
rect 323 -1479 326 -1473
rect 330 -1479 333 -1473
rect 337 -1479 340 -1473
rect 344 -1479 347 -1473
rect 351 -1479 354 -1473
rect 358 -1479 361 -1473
rect 365 -1479 368 -1473
rect 372 -1479 375 -1473
rect 379 -1479 382 -1473
rect 386 -1479 392 -1473
rect 393 -1479 396 -1473
rect 400 -1479 403 -1473
rect 407 -1479 413 -1473
rect 414 -1479 420 -1473
rect 421 -1479 424 -1473
rect 428 -1479 431 -1473
rect 435 -1479 438 -1473
rect 442 -1479 445 -1473
rect 449 -1479 452 -1473
rect 456 -1479 459 -1473
rect 463 -1479 466 -1473
rect 470 -1479 473 -1473
rect 477 -1479 480 -1473
rect 484 -1479 487 -1473
rect 491 -1479 494 -1473
rect 498 -1479 504 -1473
rect 505 -1479 508 -1473
rect 512 -1479 515 -1473
rect 519 -1479 522 -1473
rect 526 -1479 529 -1473
rect 533 -1479 536 -1473
rect 540 -1479 543 -1473
rect 547 -1479 550 -1473
rect 554 -1479 560 -1473
rect 561 -1479 564 -1473
rect 568 -1479 571 -1473
rect 575 -1479 578 -1473
rect 582 -1479 585 -1473
rect 589 -1479 595 -1473
rect 596 -1479 602 -1473
rect 603 -1479 606 -1473
rect 610 -1479 616 -1473
rect 617 -1479 620 -1473
rect 624 -1479 627 -1473
rect 631 -1479 637 -1473
rect 638 -1479 644 -1473
rect 645 -1479 648 -1473
rect 652 -1479 655 -1473
rect 659 -1479 662 -1473
rect 666 -1479 669 -1473
rect 673 -1479 679 -1473
rect 680 -1479 683 -1473
rect 687 -1479 690 -1473
rect 694 -1479 697 -1473
rect 701 -1479 704 -1473
rect 708 -1479 711 -1473
rect 715 -1479 721 -1473
rect 722 -1479 728 -1473
rect 729 -1479 735 -1473
rect 736 -1479 739 -1473
rect 743 -1479 746 -1473
rect 750 -1479 753 -1473
rect 757 -1479 760 -1473
rect 764 -1479 770 -1473
rect 771 -1479 774 -1473
rect 778 -1479 781 -1473
rect 785 -1479 788 -1473
rect 792 -1479 795 -1473
rect 799 -1479 802 -1473
rect 806 -1479 809 -1473
rect 813 -1479 816 -1473
rect 820 -1479 823 -1473
rect 827 -1479 830 -1473
rect 834 -1479 837 -1473
rect 841 -1479 844 -1473
rect 848 -1479 851 -1473
rect 855 -1479 858 -1473
rect 862 -1479 868 -1473
rect 869 -1479 875 -1473
rect 876 -1479 879 -1473
rect 883 -1479 886 -1473
rect 890 -1479 896 -1473
rect 897 -1479 903 -1473
rect 904 -1479 907 -1473
rect 911 -1479 914 -1473
rect 918 -1479 921 -1473
rect 925 -1479 928 -1473
rect 932 -1479 938 -1473
rect 939 -1479 942 -1473
rect 946 -1479 949 -1473
rect 953 -1479 956 -1473
rect 960 -1479 963 -1473
rect 967 -1479 970 -1473
rect 974 -1479 977 -1473
rect 981 -1479 984 -1473
rect 988 -1479 991 -1473
rect 995 -1479 998 -1473
rect 1002 -1479 1005 -1473
rect 1009 -1479 1012 -1473
rect 1016 -1479 1019 -1473
rect 1023 -1479 1029 -1473
rect 1030 -1479 1033 -1473
rect 1037 -1479 1040 -1473
rect 1044 -1479 1047 -1473
rect 1051 -1479 1054 -1473
rect 1058 -1479 1061 -1473
rect 1065 -1479 1071 -1473
rect 1072 -1479 1075 -1473
rect 1079 -1479 1082 -1473
rect 1086 -1479 1089 -1473
rect 1093 -1479 1096 -1473
rect 1100 -1479 1103 -1473
rect 1107 -1479 1110 -1473
rect 1114 -1479 1117 -1473
rect 1121 -1479 1127 -1473
rect 1128 -1479 1131 -1473
rect 1135 -1479 1141 -1473
rect 1142 -1479 1148 -1473
rect 1149 -1479 1152 -1473
rect 1156 -1479 1159 -1473
rect 1163 -1479 1166 -1473
rect 1170 -1479 1173 -1473
rect 1177 -1479 1180 -1473
rect 1184 -1479 1187 -1473
rect 1191 -1479 1194 -1473
rect 1198 -1479 1201 -1473
rect 1205 -1479 1208 -1473
rect 1212 -1479 1215 -1473
rect 1219 -1479 1222 -1473
rect 1226 -1479 1229 -1473
rect 1233 -1479 1236 -1473
rect 1240 -1479 1243 -1473
rect 1247 -1479 1250 -1473
rect 1254 -1479 1257 -1473
rect 1261 -1479 1264 -1473
rect 1268 -1479 1271 -1473
rect 1275 -1479 1278 -1473
rect 1282 -1479 1285 -1473
rect 1289 -1479 1292 -1473
rect 1296 -1479 1299 -1473
rect 1303 -1479 1306 -1473
rect 1310 -1479 1313 -1473
rect 1317 -1479 1320 -1473
rect 1324 -1479 1327 -1473
rect 1331 -1479 1334 -1473
rect 1338 -1479 1341 -1473
rect 1345 -1479 1348 -1473
rect 1352 -1479 1355 -1473
rect 1359 -1479 1362 -1473
rect 1366 -1479 1369 -1473
rect 1373 -1479 1376 -1473
rect 1380 -1479 1383 -1473
rect 1387 -1479 1390 -1473
rect 1394 -1479 1397 -1473
rect 1401 -1479 1404 -1473
rect 1408 -1479 1411 -1473
rect 1415 -1479 1418 -1473
rect 1422 -1479 1425 -1473
rect 1429 -1479 1432 -1473
rect 1436 -1479 1439 -1473
rect 1443 -1479 1446 -1473
rect 1450 -1479 1453 -1473
rect 1457 -1479 1460 -1473
rect 1464 -1479 1467 -1473
rect 1471 -1479 1474 -1473
rect 1478 -1479 1481 -1473
rect 1485 -1479 1488 -1473
rect 1492 -1479 1495 -1473
rect 1499 -1479 1502 -1473
rect 1506 -1479 1509 -1473
rect 1513 -1479 1516 -1473
rect 1520 -1479 1523 -1473
rect 1527 -1479 1530 -1473
rect 1534 -1479 1537 -1473
rect 1541 -1479 1544 -1473
rect 1548 -1479 1551 -1473
rect 1555 -1479 1558 -1473
rect 1562 -1479 1565 -1473
rect 1569 -1479 1572 -1473
rect 1576 -1479 1579 -1473
rect 1583 -1479 1586 -1473
rect 1590 -1479 1593 -1473
rect 1597 -1479 1600 -1473
rect 1604 -1479 1607 -1473
rect 1611 -1479 1614 -1473
rect 1618 -1479 1621 -1473
rect 1625 -1479 1628 -1473
rect 1632 -1479 1635 -1473
rect 1639 -1479 1642 -1473
rect 1646 -1479 1649 -1473
rect 1653 -1479 1656 -1473
rect 1660 -1479 1663 -1473
rect 1667 -1479 1670 -1473
rect 1674 -1479 1677 -1473
rect 1681 -1479 1684 -1473
rect 1688 -1479 1691 -1473
rect 1695 -1479 1701 -1473
rect 1702 -1479 1705 -1473
rect 1709 -1479 1712 -1473
rect 1716 -1479 1722 -1473
rect 1723 -1479 1726 -1473
rect 1744 -1479 1747 -1473
rect 1 -1616 7 -1610
rect 8 -1616 14 -1610
rect 15 -1616 21 -1610
rect 22 -1616 25 -1610
rect 29 -1616 32 -1610
rect 36 -1616 42 -1610
rect 43 -1616 46 -1610
rect 50 -1616 53 -1610
rect 57 -1616 63 -1610
rect 64 -1616 70 -1610
rect 71 -1616 74 -1610
rect 78 -1616 81 -1610
rect 85 -1616 88 -1610
rect 92 -1616 98 -1610
rect 99 -1616 102 -1610
rect 106 -1616 109 -1610
rect 113 -1616 116 -1610
rect 120 -1616 123 -1610
rect 127 -1616 130 -1610
rect 134 -1616 137 -1610
rect 141 -1616 144 -1610
rect 148 -1616 151 -1610
rect 155 -1616 158 -1610
rect 162 -1616 165 -1610
rect 169 -1616 172 -1610
rect 176 -1616 179 -1610
rect 183 -1616 186 -1610
rect 190 -1616 196 -1610
rect 197 -1616 200 -1610
rect 204 -1616 210 -1610
rect 211 -1616 214 -1610
rect 218 -1616 221 -1610
rect 225 -1616 228 -1610
rect 232 -1616 235 -1610
rect 239 -1616 242 -1610
rect 246 -1616 249 -1610
rect 253 -1616 259 -1610
rect 260 -1616 263 -1610
rect 267 -1616 273 -1610
rect 274 -1616 277 -1610
rect 281 -1616 284 -1610
rect 288 -1616 294 -1610
rect 295 -1616 298 -1610
rect 302 -1616 305 -1610
rect 309 -1616 312 -1610
rect 316 -1616 322 -1610
rect 323 -1616 326 -1610
rect 330 -1616 333 -1610
rect 337 -1616 340 -1610
rect 344 -1616 347 -1610
rect 351 -1616 354 -1610
rect 358 -1616 361 -1610
rect 365 -1616 371 -1610
rect 372 -1616 375 -1610
rect 379 -1616 385 -1610
rect 386 -1616 389 -1610
rect 393 -1616 396 -1610
rect 400 -1616 403 -1610
rect 407 -1616 410 -1610
rect 414 -1616 417 -1610
rect 421 -1616 424 -1610
rect 428 -1616 431 -1610
rect 435 -1616 438 -1610
rect 442 -1616 445 -1610
rect 449 -1616 452 -1610
rect 456 -1616 459 -1610
rect 463 -1616 466 -1610
rect 470 -1616 476 -1610
rect 477 -1616 480 -1610
rect 484 -1616 487 -1610
rect 491 -1616 497 -1610
rect 498 -1616 501 -1610
rect 505 -1616 508 -1610
rect 512 -1616 515 -1610
rect 519 -1616 522 -1610
rect 526 -1616 532 -1610
rect 533 -1616 536 -1610
rect 540 -1616 546 -1610
rect 547 -1616 550 -1610
rect 554 -1616 557 -1610
rect 561 -1616 567 -1610
rect 568 -1616 571 -1610
rect 575 -1616 578 -1610
rect 582 -1616 585 -1610
rect 589 -1616 592 -1610
rect 596 -1616 599 -1610
rect 603 -1616 609 -1610
rect 610 -1616 616 -1610
rect 617 -1616 623 -1610
rect 624 -1616 627 -1610
rect 631 -1616 634 -1610
rect 638 -1616 641 -1610
rect 645 -1616 648 -1610
rect 652 -1616 655 -1610
rect 659 -1616 662 -1610
rect 666 -1616 672 -1610
rect 673 -1616 676 -1610
rect 680 -1616 683 -1610
rect 687 -1616 690 -1610
rect 694 -1616 697 -1610
rect 701 -1616 704 -1610
rect 708 -1616 714 -1610
rect 715 -1616 721 -1610
rect 722 -1616 728 -1610
rect 729 -1616 732 -1610
rect 736 -1616 742 -1610
rect 743 -1616 749 -1610
rect 750 -1616 753 -1610
rect 757 -1616 763 -1610
rect 764 -1616 767 -1610
rect 771 -1616 774 -1610
rect 778 -1616 781 -1610
rect 785 -1616 788 -1610
rect 792 -1616 798 -1610
rect 799 -1616 802 -1610
rect 806 -1616 812 -1610
rect 813 -1616 816 -1610
rect 820 -1616 823 -1610
rect 827 -1616 830 -1610
rect 834 -1616 837 -1610
rect 841 -1616 844 -1610
rect 848 -1616 851 -1610
rect 855 -1616 858 -1610
rect 862 -1616 865 -1610
rect 869 -1616 872 -1610
rect 876 -1616 879 -1610
rect 883 -1616 886 -1610
rect 890 -1616 893 -1610
rect 897 -1616 900 -1610
rect 904 -1616 907 -1610
rect 911 -1616 914 -1610
rect 918 -1616 921 -1610
rect 925 -1616 931 -1610
rect 932 -1616 935 -1610
rect 939 -1616 942 -1610
rect 946 -1616 949 -1610
rect 953 -1616 956 -1610
rect 960 -1616 963 -1610
rect 967 -1616 970 -1610
rect 974 -1616 977 -1610
rect 981 -1616 984 -1610
rect 988 -1616 991 -1610
rect 995 -1616 998 -1610
rect 1002 -1616 1005 -1610
rect 1009 -1616 1012 -1610
rect 1016 -1616 1022 -1610
rect 1023 -1616 1026 -1610
rect 1030 -1616 1033 -1610
rect 1037 -1616 1040 -1610
rect 1044 -1616 1050 -1610
rect 1051 -1616 1054 -1610
rect 1058 -1616 1064 -1610
rect 1065 -1616 1068 -1610
rect 1072 -1616 1075 -1610
rect 1079 -1616 1082 -1610
rect 1086 -1616 1089 -1610
rect 1093 -1616 1096 -1610
rect 1100 -1616 1106 -1610
rect 1107 -1616 1110 -1610
rect 1114 -1616 1120 -1610
rect 1121 -1616 1124 -1610
rect 1128 -1616 1131 -1610
rect 1135 -1616 1138 -1610
rect 1142 -1616 1145 -1610
rect 1149 -1616 1155 -1610
rect 1156 -1616 1159 -1610
rect 1163 -1616 1166 -1610
rect 1170 -1616 1173 -1610
rect 1177 -1616 1180 -1610
rect 1184 -1616 1187 -1610
rect 1191 -1616 1194 -1610
rect 1198 -1616 1201 -1610
rect 1205 -1616 1208 -1610
rect 1212 -1616 1215 -1610
rect 1219 -1616 1222 -1610
rect 1226 -1616 1229 -1610
rect 1233 -1616 1236 -1610
rect 1240 -1616 1243 -1610
rect 1247 -1616 1250 -1610
rect 1254 -1616 1260 -1610
rect 1261 -1616 1264 -1610
rect 1268 -1616 1271 -1610
rect 1275 -1616 1278 -1610
rect 1282 -1616 1285 -1610
rect 1289 -1616 1292 -1610
rect 1296 -1616 1299 -1610
rect 1303 -1616 1306 -1610
rect 1310 -1616 1313 -1610
rect 1317 -1616 1320 -1610
rect 1324 -1616 1327 -1610
rect 1331 -1616 1334 -1610
rect 1338 -1616 1341 -1610
rect 1345 -1616 1348 -1610
rect 1352 -1616 1355 -1610
rect 1359 -1616 1362 -1610
rect 1366 -1616 1369 -1610
rect 1373 -1616 1376 -1610
rect 1380 -1616 1383 -1610
rect 1387 -1616 1390 -1610
rect 1394 -1616 1397 -1610
rect 1401 -1616 1404 -1610
rect 1408 -1616 1411 -1610
rect 1415 -1616 1418 -1610
rect 1422 -1616 1425 -1610
rect 1429 -1616 1432 -1610
rect 1436 -1616 1439 -1610
rect 1443 -1616 1446 -1610
rect 1450 -1616 1453 -1610
rect 1457 -1616 1460 -1610
rect 1464 -1616 1467 -1610
rect 1471 -1616 1474 -1610
rect 1478 -1616 1481 -1610
rect 1485 -1616 1488 -1610
rect 1492 -1616 1495 -1610
rect 1499 -1616 1502 -1610
rect 1506 -1616 1509 -1610
rect 1513 -1616 1516 -1610
rect 1520 -1616 1523 -1610
rect 1527 -1616 1530 -1610
rect 1534 -1616 1537 -1610
rect 1541 -1616 1544 -1610
rect 1548 -1616 1551 -1610
rect 1555 -1616 1558 -1610
rect 1562 -1616 1565 -1610
rect 1569 -1616 1572 -1610
rect 1576 -1616 1579 -1610
rect 1583 -1616 1586 -1610
rect 1590 -1616 1593 -1610
rect 1597 -1616 1600 -1610
rect 1604 -1616 1607 -1610
rect 1611 -1616 1614 -1610
rect 1618 -1616 1621 -1610
rect 1625 -1616 1628 -1610
rect 1632 -1616 1635 -1610
rect 1639 -1616 1642 -1610
rect 1646 -1616 1649 -1610
rect 1653 -1616 1656 -1610
rect 1660 -1616 1663 -1610
rect 1667 -1616 1670 -1610
rect 1674 -1616 1677 -1610
rect 1681 -1616 1684 -1610
rect 1688 -1616 1691 -1610
rect 1695 -1616 1698 -1610
rect 1702 -1616 1708 -1610
rect 1709 -1616 1715 -1610
rect 1716 -1616 1719 -1610
rect 1751 -1616 1754 -1610
rect 1 -1743 7 -1737
rect 8 -1743 14 -1737
rect 15 -1743 21 -1737
rect 22 -1743 28 -1737
rect 29 -1743 35 -1737
rect 36 -1743 39 -1737
rect 43 -1743 46 -1737
rect 50 -1743 53 -1737
rect 57 -1743 63 -1737
rect 64 -1743 67 -1737
rect 71 -1743 74 -1737
rect 78 -1743 81 -1737
rect 85 -1743 88 -1737
rect 92 -1743 95 -1737
rect 99 -1743 102 -1737
rect 106 -1743 109 -1737
rect 113 -1743 116 -1737
rect 120 -1743 123 -1737
rect 127 -1743 130 -1737
rect 134 -1743 137 -1737
rect 141 -1743 144 -1737
rect 148 -1743 151 -1737
rect 155 -1743 161 -1737
rect 162 -1743 165 -1737
rect 169 -1743 175 -1737
rect 176 -1743 182 -1737
rect 183 -1743 186 -1737
rect 190 -1743 196 -1737
rect 197 -1743 200 -1737
rect 204 -1743 207 -1737
rect 211 -1743 214 -1737
rect 218 -1743 221 -1737
rect 225 -1743 228 -1737
rect 232 -1743 235 -1737
rect 239 -1743 242 -1737
rect 246 -1743 249 -1737
rect 253 -1743 259 -1737
rect 260 -1743 266 -1737
rect 267 -1743 270 -1737
rect 274 -1743 280 -1737
rect 281 -1743 284 -1737
rect 288 -1743 291 -1737
rect 295 -1743 298 -1737
rect 302 -1743 305 -1737
rect 309 -1743 312 -1737
rect 316 -1743 319 -1737
rect 323 -1743 326 -1737
rect 330 -1743 333 -1737
rect 337 -1743 340 -1737
rect 344 -1743 350 -1737
rect 351 -1743 354 -1737
rect 358 -1743 361 -1737
rect 365 -1743 368 -1737
rect 372 -1743 375 -1737
rect 379 -1743 382 -1737
rect 386 -1743 389 -1737
rect 393 -1743 396 -1737
rect 400 -1743 403 -1737
rect 407 -1743 413 -1737
rect 414 -1743 417 -1737
rect 421 -1743 424 -1737
rect 428 -1743 434 -1737
rect 435 -1743 438 -1737
rect 442 -1743 445 -1737
rect 449 -1743 452 -1737
rect 456 -1743 459 -1737
rect 463 -1743 466 -1737
rect 470 -1743 473 -1737
rect 477 -1743 483 -1737
rect 484 -1743 487 -1737
rect 491 -1743 494 -1737
rect 498 -1743 501 -1737
rect 505 -1743 508 -1737
rect 512 -1743 515 -1737
rect 519 -1743 522 -1737
rect 526 -1743 532 -1737
rect 533 -1743 536 -1737
rect 540 -1743 546 -1737
rect 547 -1743 550 -1737
rect 554 -1743 557 -1737
rect 561 -1743 564 -1737
rect 568 -1743 571 -1737
rect 575 -1743 578 -1737
rect 582 -1743 585 -1737
rect 589 -1743 592 -1737
rect 596 -1743 599 -1737
rect 603 -1743 606 -1737
rect 610 -1743 613 -1737
rect 617 -1743 620 -1737
rect 624 -1743 627 -1737
rect 631 -1743 634 -1737
rect 638 -1743 641 -1737
rect 645 -1743 648 -1737
rect 652 -1743 655 -1737
rect 659 -1743 662 -1737
rect 666 -1743 669 -1737
rect 673 -1743 679 -1737
rect 680 -1743 683 -1737
rect 687 -1743 693 -1737
rect 694 -1743 697 -1737
rect 701 -1743 707 -1737
rect 708 -1743 711 -1737
rect 715 -1743 718 -1737
rect 722 -1743 728 -1737
rect 729 -1743 735 -1737
rect 736 -1743 742 -1737
rect 743 -1743 746 -1737
rect 750 -1743 753 -1737
rect 757 -1743 760 -1737
rect 764 -1743 767 -1737
rect 771 -1743 774 -1737
rect 778 -1743 784 -1737
rect 785 -1743 791 -1737
rect 792 -1743 795 -1737
rect 799 -1743 805 -1737
rect 806 -1743 812 -1737
rect 813 -1743 816 -1737
rect 820 -1743 823 -1737
rect 827 -1743 833 -1737
rect 834 -1743 837 -1737
rect 841 -1743 844 -1737
rect 848 -1743 851 -1737
rect 855 -1743 858 -1737
rect 862 -1743 865 -1737
rect 869 -1743 875 -1737
rect 876 -1743 879 -1737
rect 883 -1743 889 -1737
rect 890 -1743 896 -1737
rect 897 -1743 900 -1737
rect 904 -1743 907 -1737
rect 911 -1743 917 -1737
rect 918 -1743 924 -1737
rect 925 -1743 931 -1737
rect 932 -1743 935 -1737
rect 939 -1743 942 -1737
rect 946 -1743 949 -1737
rect 953 -1743 956 -1737
rect 960 -1743 963 -1737
rect 967 -1743 970 -1737
rect 974 -1743 980 -1737
rect 981 -1743 984 -1737
rect 988 -1743 994 -1737
rect 995 -1743 998 -1737
rect 1002 -1743 1005 -1737
rect 1009 -1743 1012 -1737
rect 1016 -1743 1019 -1737
rect 1023 -1743 1026 -1737
rect 1030 -1743 1033 -1737
rect 1037 -1743 1040 -1737
rect 1044 -1743 1047 -1737
rect 1051 -1743 1054 -1737
rect 1058 -1743 1061 -1737
rect 1065 -1743 1071 -1737
rect 1072 -1743 1075 -1737
rect 1079 -1743 1082 -1737
rect 1086 -1743 1089 -1737
rect 1093 -1743 1096 -1737
rect 1100 -1743 1103 -1737
rect 1107 -1743 1110 -1737
rect 1114 -1743 1120 -1737
rect 1121 -1743 1124 -1737
rect 1128 -1743 1131 -1737
rect 1135 -1743 1138 -1737
rect 1142 -1743 1145 -1737
rect 1149 -1743 1152 -1737
rect 1156 -1743 1159 -1737
rect 1163 -1743 1166 -1737
rect 1170 -1743 1173 -1737
rect 1177 -1743 1180 -1737
rect 1184 -1743 1187 -1737
rect 1191 -1743 1194 -1737
rect 1198 -1743 1201 -1737
rect 1205 -1743 1208 -1737
rect 1212 -1743 1215 -1737
rect 1219 -1743 1222 -1737
rect 1226 -1743 1229 -1737
rect 1233 -1743 1236 -1737
rect 1240 -1743 1243 -1737
rect 1247 -1743 1253 -1737
rect 1254 -1743 1257 -1737
rect 1261 -1743 1264 -1737
rect 1268 -1743 1271 -1737
rect 1275 -1743 1278 -1737
rect 1282 -1743 1285 -1737
rect 1289 -1743 1292 -1737
rect 1296 -1743 1299 -1737
rect 1303 -1743 1306 -1737
rect 1310 -1743 1313 -1737
rect 1317 -1743 1320 -1737
rect 1324 -1743 1327 -1737
rect 1331 -1743 1334 -1737
rect 1338 -1743 1341 -1737
rect 1345 -1743 1348 -1737
rect 1352 -1743 1355 -1737
rect 1359 -1743 1362 -1737
rect 1366 -1743 1369 -1737
rect 1373 -1743 1376 -1737
rect 1380 -1743 1383 -1737
rect 1387 -1743 1390 -1737
rect 1394 -1743 1397 -1737
rect 1401 -1743 1404 -1737
rect 1408 -1743 1411 -1737
rect 1415 -1743 1418 -1737
rect 1422 -1743 1425 -1737
rect 1429 -1743 1432 -1737
rect 1436 -1743 1439 -1737
rect 1443 -1743 1446 -1737
rect 1450 -1743 1453 -1737
rect 1457 -1743 1460 -1737
rect 1464 -1743 1467 -1737
rect 1471 -1743 1474 -1737
rect 1478 -1743 1481 -1737
rect 1485 -1743 1488 -1737
rect 1492 -1743 1495 -1737
rect 1499 -1743 1502 -1737
rect 1506 -1743 1509 -1737
rect 1513 -1743 1516 -1737
rect 1520 -1743 1523 -1737
rect 1527 -1743 1530 -1737
rect 1534 -1743 1537 -1737
rect 1541 -1743 1544 -1737
rect 1548 -1743 1551 -1737
rect 1555 -1743 1558 -1737
rect 1562 -1743 1565 -1737
rect 1569 -1743 1572 -1737
rect 1576 -1743 1579 -1737
rect 1583 -1743 1586 -1737
rect 1590 -1743 1593 -1737
rect 1597 -1743 1600 -1737
rect 1604 -1743 1607 -1737
rect 1611 -1743 1614 -1737
rect 1618 -1743 1621 -1737
rect 1625 -1743 1628 -1737
rect 1632 -1743 1635 -1737
rect 1639 -1743 1642 -1737
rect 1646 -1743 1649 -1737
rect 1653 -1743 1656 -1737
rect 1660 -1743 1663 -1737
rect 1667 -1743 1670 -1737
rect 1674 -1743 1677 -1737
rect 1681 -1743 1684 -1737
rect 1688 -1743 1691 -1737
rect 1695 -1743 1698 -1737
rect 1702 -1743 1705 -1737
rect 1709 -1743 1712 -1737
rect 1716 -1743 1719 -1737
rect 1723 -1743 1726 -1737
rect 1730 -1743 1733 -1737
rect 1737 -1743 1740 -1737
rect 1744 -1743 1750 -1737
rect 1751 -1743 1754 -1737
rect 1758 -1743 1761 -1737
rect 1765 -1743 1768 -1737
rect 1772 -1743 1775 -1737
rect 1779 -1743 1782 -1737
rect 1 -1890 7 -1884
rect 8 -1890 14 -1884
rect 15 -1890 21 -1884
rect 22 -1890 28 -1884
rect 29 -1890 32 -1884
rect 36 -1890 39 -1884
rect 43 -1890 46 -1884
rect 50 -1890 53 -1884
rect 57 -1890 60 -1884
rect 64 -1890 67 -1884
rect 71 -1890 74 -1884
rect 78 -1890 81 -1884
rect 85 -1890 88 -1884
rect 92 -1890 95 -1884
rect 99 -1890 102 -1884
rect 106 -1890 112 -1884
rect 113 -1890 116 -1884
rect 120 -1890 123 -1884
rect 127 -1890 130 -1884
rect 134 -1890 137 -1884
rect 141 -1890 144 -1884
rect 148 -1890 151 -1884
rect 155 -1890 161 -1884
rect 162 -1890 165 -1884
rect 169 -1890 172 -1884
rect 176 -1890 182 -1884
rect 183 -1890 186 -1884
rect 190 -1890 196 -1884
rect 197 -1890 200 -1884
rect 204 -1890 210 -1884
rect 211 -1890 214 -1884
rect 218 -1890 221 -1884
rect 225 -1890 228 -1884
rect 232 -1890 235 -1884
rect 239 -1890 242 -1884
rect 246 -1890 252 -1884
rect 253 -1890 256 -1884
rect 260 -1890 266 -1884
rect 267 -1890 270 -1884
rect 274 -1890 277 -1884
rect 281 -1890 284 -1884
rect 288 -1890 291 -1884
rect 295 -1890 298 -1884
rect 302 -1890 305 -1884
rect 309 -1890 312 -1884
rect 316 -1890 319 -1884
rect 323 -1890 326 -1884
rect 330 -1890 333 -1884
rect 337 -1890 343 -1884
rect 344 -1890 347 -1884
rect 351 -1890 354 -1884
rect 358 -1890 361 -1884
rect 365 -1890 368 -1884
rect 372 -1890 375 -1884
rect 379 -1890 382 -1884
rect 386 -1890 389 -1884
rect 393 -1890 396 -1884
rect 400 -1890 403 -1884
rect 407 -1890 410 -1884
rect 414 -1890 417 -1884
rect 421 -1890 424 -1884
rect 428 -1890 431 -1884
rect 435 -1890 438 -1884
rect 442 -1890 448 -1884
rect 449 -1890 452 -1884
rect 456 -1890 459 -1884
rect 463 -1890 469 -1884
rect 470 -1890 476 -1884
rect 477 -1890 480 -1884
rect 484 -1890 487 -1884
rect 491 -1890 494 -1884
rect 498 -1890 504 -1884
rect 505 -1890 508 -1884
rect 512 -1890 515 -1884
rect 519 -1890 522 -1884
rect 526 -1890 532 -1884
rect 533 -1890 536 -1884
rect 540 -1890 543 -1884
rect 547 -1890 550 -1884
rect 554 -1890 557 -1884
rect 561 -1890 564 -1884
rect 568 -1890 574 -1884
rect 575 -1890 578 -1884
rect 582 -1890 585 -1884
rect 589 -1890 592 -1884
rect 596 -1890 599 -1884
rect 603 -1890 606 -1884
rect 610 -1890 613 -1884
rect 617 -1890 620 -1884
rect 624 -1890 627 -1884
rect 631 -1890 634 -1884
rect 638 -1890 641 -1884
rect 645 -1890 651 -1884
rect 652 -1890 658 -1884
rect 659 -1890 662 -1884
rect 666 -1890 669 -1884
rect 673 -1890 676 -1884
rect 680 -1890 683 -1884
rect 687 -1890 690 -1884
rect 694 -1890 697 -1884
rect 701 -1890 704 -1884
rect 708 -1890 711 -1884
rect 715 -1890 718 -1884
rect 722 -1890 725 -1884
rect 729 -1890 732 -1884
rect 736 -1890 739 -1884
rect 743 -1890 746 -1884
rect 750 -1890 753 -1884
rect 757 -1890 760 -1884
rect 764 -1890 767 -1884
rect 771 -1890 774 -1884
rect 778 -1890 781 -1884
rect 785 -1890 788 -1884
rect 792 -1890 795 -1884
rect 799 -1890 805 -1884
rect 806 -1890 812 -1884
rect 813 -1890 816 -1884
rect 820 -1890 826 -1884
rect 827 -1890 833 -1884
rect 834 -1890 840 -1884
rect 841 -1890 844 -1884
rect 848 -1890 851 -1884
rect 855 -1890 858 -1884
rect 862 -1890 868 -1884
rect 869 -1890 872 -1884
rect 876 -1890 879 -1884
rect 883 -1890 886 -1884
rect 890 -1890 893 -1884
rect 897 -1890 900 -1884
rect 904 -1890 910 -1884
rect 911 -1890 914 -1884
rect 918 -1890 921 -1884
rect 925 -1890 931 -1884
rect 932 -1890 938 -1884
rect 939 -1890 942 -1884
rect 946 -1890 949 -1884
rect 953 -1890 959 -1884
rect 960 -1890 963 -1884
rect 967 -1890 970 -1884
rect 974 -1890 977 -1884
rect 981 -1890 987 -1884
rect 988 -1890 991 -1884
rect 995 -1890 998 -1884
rect 1002 -1890 1005 -1884
rect 1009 -1890 1012 -1884
rect 1016 -1890 1022 -1884
rect 1023 -1890 1029 -1884
rect 1030 -1890 1033 -1884
rect 1037 -1890 1043 -1884
rect 1044 -1890 1050 -1884
rect 1051 -1890 1054 -1884
rect 1058 -1890 1061 -1884
rect 1065 -1890 1068 -1884
rect 1072 -1890 1075 -1884
rect 1079 -1890 1082 -1884
rect 1086 -1890 1089 -1884
rect 1093 -1890 1096 -1884
rect 1100 -1890 1103 -1884
rect 1107 -1890 1113 -1884
rect 1114 -1890 1117 -1884
rect 1121 -1890 1124 -1884
rect 1128 -1890 1131 -1884
rect 1135 -1890 1138 -1884
rect 1142 -1890 1145 -1884
rect 1149 -1890 1155 -1884
rect 1156 -1890 1162 -1884
rect 1163 -1890 1166 -1884
rect 1170 -1890 1173 -1884
rect 1177 -1890 1180 -1884
rect 1184 -1890 1187 -1884
rect 1191 -1890 1194 -1884
rect 1198 -1890 1201 -1884
rect 1205 -1890 1208 -1884
rect 1212 -1890 1215 -1884
rect 1219 -1890 1222 -1884
rect 1226 -1890 1229 -1884
rect 1233 -1890 1236 -1884
rect 1240 -1890 1243 -1884
rect 1247 -1890 1250 -1884
rect 1254 -1890 1257 -1884
rect 1261 -1890 1264 -1884
rect 1268 -1890 1271 -1884
rect 1275 -1890 1281 -1884
rect 1282 -1890 1285 -1884
rect 1289 -1890 1292 -1884
rect 1296 -1890 1299 -1884
rect 1303 -1890 1306 -1884
rect 1310 -1890 1316 -1884
rect 1317 -1890 1320 -1884
rect 1324 -1890 1327 -1884
rect 1331 -1890 1334 -1884
rect 1338 -1890 1341 -1884
rect 1345 -1890 1348 -1884
rect 1352 -1890 1355 -1884
rect 1359 -1890 1362 -1884
rect 1366 -1890 1369 -1884
rect 1373 -1890 1376 -1884
rect 1380 -1890 1383 -1884
rect 1387 -1890 1390 -1884
rect 1394 -1890 1397 -1884
rect 1401 -1890 1404 -1884
rect 1408 -1890 1411 -1884
rect 1415 -1890 1418 -1884
rect 1422 -1890 1425 -1884
rect 1429 -1890 1432 -1884
rect 1436 -1890 1439 -1884
rect 1443 -1890 1446 -1884
rect 1450 -1890 1453 -1884
rect 1457 -1890 1460 -1884
rect 1464 -1890 1467 -1884
rect 1471 -1890 1474 -1884
rect 1478 -1890 1481 -1884
rect 1485 -1890 1488 -1884
rect 1492 -1890 1495 -1884
rect 1499 -1890 1502 -1884
rect 1506 -1890 1509 -1884
rect 1513 -1890 1516 -1884
rect 1520 -1890 1523 -1884
rect 1527 -1890 1530 -1884
rect 1534 -1890 1537 -1884
rect 1541 -1890 1544 -1884
rect 1548 -1890 1551 -1884
rect 1555 -1890 1558 -1884
rect 1562 -1890 1565 -1884
rect 1569 -1890 1572 -1884
rect 1576 -1890 1579 -1884
rect 1583 -1890 1586 -1884
rect 1590 -1890 1593 -1884
rect 1597 -1890 1600 -1884
rect 1604 -1890 1607 -1884
rect 1611 -1890 1614 -1884
rect 1618 -1890 1621 -1884
rect 1625 -1890 1628 -1884
rect 1632 -1890 1635 -1884
rect 1639 -1890 1642 -1884
rect 1646 -1890 1649 -1884
rect 1653 -1890 1656 -1884
rect 1660 -1890 1663 -1884
rect 1667 -1890 1670 -1884
rect 1674 -1890 1677 -1884
rect 1681 -1890 1684 -1884
rect 1688 -1890 1691 -1884
rect 1695 -1890 1698 -1884
rect 1702 -1890 1705 -1884
rect 1709 -1890 1712 -1884
rect 1716 -1890 1719 -1884
rect 1723 -1890 1726 -1884
rect 1730 -1890 1733 -1884
rect 1737 -1890 1740 -1884
rect 1744 -1890 1747 -1884
rect 1751 -1890 1754 -1884
rect 1758 -1890 1761 -1884
rect 1765 -1890 1768 -1884
rect 1772 -1890 1778 -1884
rect 1779 -1890 1782 -1884
rect 1786 -1890 1789 -1884
rect 1793 -1890 1796 -1884
rect 1800 -1890 1806 -1884
rect 1807 -1890 1810 -1884
rect 1814 -1890 1817 -1884
rect 1 -2023 7 -2017
rect 8 -2023 14 -2017
rect 15 -2023 21 -2017
rect 22 -2023 28 -2017
rect 29 -2023 32 -2017
rect 36 -2023 42 -2017
rect 43 -2023 46 -2017
rect 50 -2023 53 -2017
rect 57 -2023 60 -2017
rect 64 -2023 70 -2017
rect 71 -2023 74 -2017
rect 78 -2023 81 -2017
rect 85 -2023 91 -2017
rect 92 -2023 95 -2017
rect 99 -2023 105 -2017
rect 106 -2023 112 -2017
rect 113 -2023 116 -2017
rect 120 -2023 126 -2017
rect 127 -2023 133 -2017
rect 134 -2023 137 -2017
rect 141 -2023 147 -2017
rect 148 -2023 154 -2017
rect 155 -2023 158 -2017
rect 162 -2023 165 -2017
rect 169 -2023 172 -2017
rect 176 -2023 182 -2017
rect 183 -2023 186 -2017
rect 190 -2023 193 -2017
rect 197 -2023 200 -2017
rect 204 -2023 207 -2017
rect 211 -2023 217 -2017
rect 218 -2023 224 -2017
rect 225 -2023 228 -2017
rect 232 -2023 235 -2017
rect 239 -2023 242 -2017
rect 246 -2023 249 -2017
rect 253 -2023 256 -2017
rect 260 -2023 263 -2017
rect 267 -2023 270 -2017
rect 274 -2023 277 -2017
rect 281 -2023 284 -2017
rect 288 -2023 291 -2017
rect 295 -2023 298 -2017
rect 302 -2023 305 -2017
rect 309 -2023 312 -2017
rect 316 -2023 319 -2017
rect 323 -2023 326 -2017
rect 330 -2023 336 -2017
rect 337 -2023 340 -2017
rect 344 -2023 347 -2017
rect 351 -2023 354 -2017
rect 358 -2023 361 -2017
rect 365 -2023 368 -2017
rect 372 -2023 375 -2017
rect 379 -2023 382 -2017
rect 386 -2023 392 -2017
rect 393 -2023 396 -2017
rect 400 -2023 403 -2017
rect 407 -2023 410 -2017
rect 414 -2023 417 -2017
rect 421 -2023 424 -2017
rect 428 -2023 431 -2017
rect 435 -2023 438 -2017
rect 442 -2023 445 -2017
rect 449 -2023 452 -2017
rect 456 -2023 462 -2017
rect 463 -2023 466 -2017
rect 470 -2023 473 -2017
rect 477 -2023 480 -2017
rect 484 -2023 487 -2017
rect 491 -2023 494 -2017
rect 498 -2023 501 -2017
rect 505 -2023 511 -2017
rect 512 -2023 515 -2017
rect 519 -2023 522 -2017
rect 526 -2023 529 -2017
rect 533 -2023 536 -2017
rect 540 -2023 543 -2017
rect 547 -2023 553 -2017
rect 554 -2023 557 -2017
rect 561 -2023 564 -2017
rect 568 -2023 574 -2017
rect 575 -2023 578 -2017
rect 582 -2023 585 -2017
rect 589 -2023 595 -2017
rect 596 -2023 599 -2017
rect 603 -2023 606 -2017
rect 610 -2023 613 -2017
rect 617 -2023 620 -2017
rect 624 -2023 630 -2017
rect 631 -2023 634 -2017
rect 638 -2023 641 -2017
rect 645 -2023 648 -2017
rect 652 -2023 655 -2017
rect 659 -2023 662 -2017
rect 666 -2023 669 -2017
rect 673 -2023 676 -2017
rect 680 -2023 683 -2017
rect 687 -2023 690 -2017
rect 694 -2023 697 -2017
rect 701 -2023 704 -2017
rect 708 -2023 711 -2017
rect 715 -2023 721 -2017
rect 722 -2023 725 -2017
rect 729 -2023 732 -2017
rect 736 -2023 739 -2017
rect 743 -2023 746 -2017
rect 750 -2023 753 -2017
rect 757 -2023 763 -2017
rect 764 -2023 767 -2017
rect 771 -2023 774 -2017
rect 778 -2023 781 -2017
rect 785 -2023 788 -2017
rect 792 -2023 798 -2017
rect 799 -2023 802 -2017
rect 806 -2023 809 -2017
rect 813 -2023 816 -2017
rect 820 -2023 823 -2017
rect 827 -2023 830 -2017
rect 834 -2023 837 -2017
rect 841 -2023 844 -2017
rect 848 -2023 851 -2017
rect 855 -2023 858 -2017
rect 862 -2023 865 -2017
rect 869 -2023 872 -2017
rect 876 -2023 879 -2017
rect 883 -2023 889 -2017
rect 890 -2023 896 -2017
rect 897 -2023 903 -2017
rect 904 -2023 907 -2017
rect 911 -2023 914 -2017
rect 918 -2023 924 -2017
rect 925 -2023 928 -2017
rect 932 -2023 935 -2017
rect 939 -2023 942 -2017
rect 946 -2023 949 -2017
rect 953 -2023 959 -2017
rect 960 -2023 966 -2017
rect 967 -2023 970 -2017
rect 974 -2023 977 -2017
rect 981 -2023 984 -2017
rect 988 -2023 994 -2017
rect 995 -2023 1001 -2017
rect 1002 -2023 1005 -2017
rect 1009 -2023 1012 -2017
rect 1016 -2023 1019 -2017
rect 1023 -2023 1026 -2017
rect 1030 -2023 1033 -2017
rect 1037 -2023 1043 -2017
rect 1044 -2023 1047 -2017
rect 1051 -2023 1054 -2017
rect 1058 -2023 1061 -2017
rect 1065 -2023 1068 -2017
rect 1072 -2023 1075 -2017
rect 1079 -2023 1082 -2017
rect 1086 -2023 1089 -2017
rect 1093 -2023 1096 -2017
rect 1100 -2023 1103 -2017
rect 1107 -2023 1113 -2017
rect 1114 -2023 1117 -2017
rect 1121 -2023 1124 -2017
rect 1128 -2023 1131 -2017
rect 1135 -2023 1141 -2017
rect 1142 -2023 1145 -2017
rect 1149 -2023 1152 -2017
rect 1156 -2023 1159 -2017
rect 1163 -2023 1166 -2017
rect 1170 -2023 1173 -2017
rect 1177 -2023 1180 -2017
rect 1184 -2023 1187 -2017
rect 1191 -2023 1197 -2017
rect 1198 -2023 1201 -2017
rect 1205 -2023 1208 -2017
rect 1212 -2023 1218 -2017
rect 1219 -2023 1222 -2017
rect 1226 -2023 1229 -2017
rect 1233 -2023 1236 -2017
rect 1240 -2023 1243 -2017
rect 1247 -2023 1250 -2017
rect 1254 -2023 1257 -2017
rect 1261 -2023 1264 -2017
rect 1268 -2023 1271 -2017
rect 1275 -2023 1278 -2017
rect 1282 -2023 1285 -2017
rect 1289 -2023 1295 -2017
rect 1296 -2023 1299 -2017
rect 1303 -2023 1306 -2017
rect 1310 -2023 1313 -2017
rect 1317 -2023 1320 -2017
rect 1324 -2023 1327 -2017
rect 1331 -2023 1334 -2017
rect 1338 -2023 1341 -2017
rect 1345 -2023 1348 -2017
rect 1352 -2023 1355 -2017
rect 1359 -2023 1362 -2017
rect 1366 -2023 1369 -2017
rect 1373 -2023 1376 -2017
rect 1380 -2023 1383 -2017
rect 1387 -2023 1390 -2017
rect 1394 -2023 1397 -2017
rect 1401 -2023 1404 -2017
rect 1408 -2023 1411 -2017
rect 1415 -2023 1418 -2017
rect 1422 -2023 1425 -2017
rect 1429 -2023 1432 -2017
rect 1436 -2023 1439 -2017
rect 1443 -2023 1446 -2017
rect 1450 -2023 1453 -2017
rect 1457 -2023 1460 -2017
rect 1464 -2023 1467 -2017
rect 1471 -2023 1474 -2017
rect 1478 -2023 1481 -2017
rect 1485 -2023 1488 -2017
rect 1492 -2023 1495 -2017
rect 1499 -2023 1502 -2017
rect 1506 -2023 1509 -2017
rect 1513 -2023 1516 -2017
rect 1520 -2023 1523 -2017
rect 1527 -2023 1530 -2017
rect 1534 -2023 1537 -2017
rect 1541 -2023 1544 -2017
rect 1548 -2023 1551 -2017
rect 1555 -2023 1558 -2017
rect 1562 -2023 1565 -2017
rect 1569 -2023 1572 -2017
rect 1576 -2023 1579 -2017
rect 1583 -2023 1586 -2017
rect 1590 -2023 1593 -2017
rect 1597 -2023 1600 -2017
rect 1604 -2023 1607 -2017
rect 1611 -2023 1614 -2017
rect 1618 -2023 1621 -2017
rect 1625 -2023 1628 -2017
rect 1632 -2023 1635 -2017
rect 1639 -2023 1642 -2017
rect 1646 -2023 1649 -2017
rect 1653 -2023 1656 -2017
rect 1660 -2023 1663 -2017
rect 1667 -2023 1670 -2017
rect 1674 -2023 1677 -2017
rect 1681 -2023 1684 -2017
rect 1688 -2023 1691 -2017
rect 1695 -2023 1698 -2017
rect 1702 -2023 1705 -2017
rect 1709 -2023 1712 -2017
rect 1716 -2023 1719 -2017
rect 1723 -2023 1726 -2017
rect 1730 -2023 1733 -2017
rect 1737 -2023 1740 -2017
rect 1744 -2023 1750 -2017
rect 1751 -2023 1754 -2017
rect 1758 -2023 1761 -2017
rect 1765 -2023 1768 -2017
rect 1772 -2023 1775 -2017
rect 1779 -2023 1782 -2017
rect 1786 -2023 1789 -2017
rect 1793 -2023 1796 -2017
rect 1800 -2023 1803 -2017
rect 1807 -2023 1810 -2017
rect 1 -2178 7 -2172
rect 8 -2178 14 -2172
rect 15 -2178 21 -2172
rect 22 -2178 28 -2172
rect 29 -2178 32 -2172
rect 36 -2178 39 -2172
rect 43 -2178 46 -2172
rect 50 -2178 53 -2172
rect 57 -2178 63 -2172
rect 64 -2178 67 -2172
rect 71 -2178 74 -2172
rect 78 -2178 81 -2172
rect 85 -2178 88 -2172
rect 92 -2178 98 -2172
rect 99 -2178 105 -2172
rect 106 -2178 112 -2172
rect 113 -2178 116 -2172
rect 120 -2178 126 -2172
rect 127 -2178 133 -2172
rect 134 -2178 137 -2172
rect 141 -2178 144 -2172
rect 148 -2178 151 -2172
rect 155 -2178 158 -2172
rect 162 -2178 165 -2172
rect 169 -2178 172 -2172
rect 176 -2178 179 -2172
rect 183 -2178 186 -2172
rect 190 -2178 193 -2172
rect 197 -2178 203 -2172
rect 204 -2178 207 -2172
rect 211 -2178 214 -2172
rect 218 -2178 221 -2172
rect 225 -2178 231 -2172
rect 232 -2178 235 -2172
rect 239 -2178 242 -2172
rect 246 -2178 252 -2172
rect 253 -2178 259 -2172
rect 260 -2178 263 -2172
rect 267 -2178 270 -2172
rect 274 -2178 280 -2172
rect 281 -2178 284 -2172
rect 288 -2178 294 -2172
rect 295 -2178 298 -2172
rect 302 -2178 305 -2172
rect 309 -2178 312 -2172
rect 316 -2178 319 -2172
rect 323 -2178 326 -2172
rect 330 -2178 333 -2172
rect 337 -2178 340 -2172
rect 344 -2178 347 -2172
rect 351 -2178 354 -2172
rect 358 -2178 361 -2172
rect 365 -2178 368 -2172
rect 372 -2178 378 -2172
rect 379 -2178 382 -2172
rect 386 -2178 389 -2172
rect 393 -2178 396 -2172
rect 400 -2178 403 -2172
rect 407 -2178 410 -2172
rect 414 -2178 420 -2172
rect 421 -2178 424 -2172
rect 428 -2178 431 -2172
rect 435 -2178 438 -2172
rect 442 -2178 445 -2172
rect 449 -2178 452 -2172
rect 456 -2178 459 -2172
rect 463 -2178 466 -2172
rect 470 -2178 473 -2172
rect 477 -2178 480 -2172
rect 484 -2178 487 -2172
rect 491 -2178 494 -2172
rect 498 -2178 501 -2172
rect 505 -2178 508 -2172
rect 512 -2178 518 -2172
rect 519 -2178 522 -2172
rect 526 -2178 529 -2172
rect 533 -2178 536 -2172
rect 540 -2178 543 -2172
rect 547 -2178 550 -2172
rect 554 -2178 560 -2172
rect 561 -2178 564 -2172
rect 568 -2178 571 -2172
rect 575 -2178 578 -2172
rect 582 -2178 588 -2172
rect 589 -2178 592 -2172
rect 596 -2178 599 -2172
rect 603 -2178 606 -2172
rect 610 -2178 616 -2172
rect 617 -2178 620 -2172
rect 624 -2178 630 -2172
rect 631 -2178 634 -2172
rect 638 -2178 641 -2172
rect 645 -2178 648 -2172
rect 652 -2178 655 -2172
rect 659 -2178 662 -2172
rect 666 -2178 669 -2172
rect 673 -2178 676 -2172
rect 680 -2178 683 -2172
rect 687 -2178 690 -2172
rect 694 -2178 697 -2172
rect 701 -2178 707 -2172
rect 708 -2178 714 -2172
rect 715 -2178 718 -2172
rect 722 -2178 725 -2172
rect 729 -2178 732 -2172
rect 736 -2178 739 -2172
rect 743 -2178 746 -2172
rect 750 -2178 753 -2172
rect 757 -2178 760 -2172
rect 764 -2178 767 -2172
rect 771 -2178 774 -2172
rect 778 -2178 781 -2172
rect 785 -2178 788 -2172
rect 792 -2178 795 -2172
rect 799 -2178 805 -2172
rect 806 -2178 809 -2172
rect 813 -2178 819 -2172
rect 820 -2178 826 -2172
rect 827 -2178 833 -2172
rect 834 -2178 837 -2172
rect 841 -2178 844 -2172
rect 848 -2178 851 -2172
rect 855 -2178 858 -2172
rect 862 -2178 865 -2172
rect 869 -2178 875 -2172
rect 876 -2178 879 -2172
rect 883 -2178 886 -2172
rect 890 -2178 893 -2172
rect 897 -2178 900 -2172
rect 904 -2178 907 -2172
rect 911 -2178 914 -2172
rect 918 -2178 921 -2172
rect 925 -2178 931 -2172
rect 932 -2178 935 -2172
rect 939 -2178 942 -2172
rect 946 -2178 949 -2172
rect 953 -2178 956 -2172
rect 960 -2178 963 -2172
rect 967 -2178 970 -2172
rect 974 -2178 980 -2172
rect 981 -2178 984 -2172
rect 988 -2178 991 -2172
rect 995 -2178 1001 -2172
rect 1002 -2178 1005 -2172
rect 1009 -2178 1012 -2172
rect 1016 -2178 1019 -2172
rect 1023 -2178 1029 -2172
rect 1030 -2178 1033 -2172
rect 1037 -2178 1040 -2172
rect 1044 -2178 1047 -2172
rect 1051 -2178 1054 -2172
rect 1058 -2178 1064 -2172
rect 1065 -2178 1068 -2172
rect 1072 -2178 1075 -2172
rect 1079 -2178 1082 -2172
rect 1086 -2178 1089 -2172
rect 1093 -2178 1096 -2172
rect 1100 -2178 1103 -2172
rect 1107 -2178 1110 -2172
rect 1114 -2178 1117 -2172
rect 1121 -2178 1127 -2172
rect 1128 -2178 1134 -2172
rect 1135 -2178 1138 -2172
rect 1142 -2178 1145 -2172
rect 1149 -2178 1152 -2172
rect 1156 -2178 1159 -2172
rect 1163 -2178 1166 -2172
rect 1170 -2178 1173 -2172
rect 1177 -2178 1180 -2172
rect 1184 -2178 1187 -2172
rect 1191 -2178 1197 -2172
rect 1198 -2178 1201 -2172
rect 1205 -2178 1208 -2172
rect 1212 -2178 1215 -2172
rect 1219 -2178 1222 -2172
rect 1226 -2178 1229 -2172
rect 1233 -2178 1236 -2172
rect 1240 -2178 1243 -2172
rect 1247 -2178 1250 -2172
rect 1254 -2178 1257 -2172
rect 1261 -2178 1264 -2172
rect 1268 -2178 1271 -2172
rect 1275 -2178 1278 -2172
rect 1282 -2178 1285 -2172
rect 1289 -2178 1292 -2172
rect 1296 -2178 1299 -2172
rect 1303 -2178 1306 -2172
rect 1310 -2178 1316 -2172
rect 1317 -2178 1320 -2172
rect 1324 -2178 1327 -2172
rect 1331 -2178 1334 -2172
rect 1338 -2178 1341 -2172
rect 1345 -2178 1348 -2172
rect 1352 -2178 1355 -2172
rect 1359 -2178 1362 -2172
rect 1366 -2178 1369 -2172
rect 1373 -2178 1376 -2172
rect 1380 -2178 1383 -2172
rect 1387 -2178 1390 -2172
rect 1394 -2178 1397 -2172
rect 1401 -2178 1404 -2172
rect 1408 -2178 1411 -2172
rect 1415 -2178 1418 -2172
rect 1422 -2178 1425 -2172
rect 1429 -2178 1432 -2172
rect 1436 -2178 1439 -2172
rect 1443 -2178 1446 -2172
rect 1450 -2178 1453 -2172
rect 1457 -2178 1460 -2172
rect 1464 -2178 1467 -2172
rect 1471 -2178 1474 -2172
rect 1478 -2178 1481 -2172
rect 1485 -2178 1488 -2172
rect 1492 -2178 1495 -2172
rect 1499 -2178 1502 -2172
rect 1506 -2178 1509 -2172
rect 1513 -2178 1516 -2172
rect 1520 -2178 1523 -2172
rect 1527 -2178 1530 -2172
rect 1534 -2178 1537 -2172
rect 1541 -2178 1544 -2172
rect 1548 -2178 1551 -2172
rect 1555 -2178 1558 -2172
rect 1562 -2178 1565 -2172
rect 1569 -2178 1572 -2172
rect 1576 -2178 1579 -2172
rect 1583 -2178 1586 -2172
rect 1590 -2178 1593 -2172
rect 1597 -2178 1600 -2172
rect 1604 -2178 1607 -2172
rect 1611 -2178 1614 -2172
rect 1618 -2178 1621 -2172
rect 1625 -2178 1628 -2172
rect 1632 -2178 1635 -2172
rect 1639 -2178 1642 -2172
rect 1646 -2178 1649 -2172
rect 1653 -2178 1656 -2172
rect 1660 -2178 1663 -2172
rect 1667 -2178 1670 -2172
rect 1674 -2178 1677 -2172
rect 1681 -2178 1684 -2172
rect 1688 -2178 1691 -2172
rect 1695 -2178 1698 -2172
rect 1702 -2178 1705 -2172
rect 1709 -2178 1715 -2172
rect 1716 -2178 1722 -2172
rect 1723 -2178 1726 -2172
rect 1730 -2178 1733 -2172
rect 1737 -2178 1740 -2172
rect 1 -2307 7 -2301
rect 8 -2307 14 -2301
rect 15 -2307 21 -2301
rect 22 -2307 28 -2301
rect 29 -2307 32 -2301
rect 36 -2307 42 -2301
rect 43 -2307 46 -2301
rect 50 -2307 56 -2301
rect 57 -2307 60 -2301
rect 64 -2307 67 -2301
rect 71 -2307 74 -2301
rect 78 -2307 84 -2301
rect 85 -2307 88 -2301
rect 92 -2307 95 -2301
rect 99 -2307 102 -2301
rect 106 -2307 109 -2301
rect 113 -2307 116 -2301
rect 120 -2307 123 -2301
rect 127 -2307 130 -2301
rect 134 -2307 140 -2301
rect 141 -2307 147 -2301
rect 148 -2307 154 -2301
rect 155 -2307 158 -2301
rect 162 -2307 165 -2301
rect 169 -2307 172 -2301
rect 176 -2307 179 -2301
rect 183 -2307 186 -2301
rect 190 -2307 193 -2301
rect 197 -2307 200 -2301
rect 204 -2307 210 -2301
rect 211 -2307 217 -2301
rect 218 -2307 221 -2301
rect 225 -2307 228 -2301
rect 232 -2307 235 -2301
rect 239 -2307 242 -2301
rect 246 -2307 249 -2301
rect 253 -2307 256 -2301
rect 260 -2307 263 -2301
rect 267 -2307 270 -2301
rect 274 -2307 277 -2301
rect 281 -2307 287 -2301
rect 288 -2307 291 -2301
rect 295 -2307 298 -2301
rect 302 -2307 305 -2301
rect 309 -2307 312 -2301
rect 316 -2307 319 -2301
rect 323 -2307 326 -2301
rect 330 -2307 333 -2301
rect 337 -2307 340 -2301
rect 344 -2307 347 -2301
rect 351 -2307 354 -2301
rect 358 -2307 361 -2301
rect 365 -2307 368 -2301
rect 372 -2307 375 -2301
rect 379 -2307 382 -2301
rect 386 -2307 389 -2301
rect 393 -2307 396 -2301
rect 400 -2307 403 -2301
rect 407 -2307 410 -2301
rect 414 -2307 417 -2301
rect 421 -2307 424 -2301
rect 428 -2307 431 -2301
rect 435 -2307 438 -2301
rect 442 -2307 445 -2301
rect 449 -2307 455 -2301
rect 456 -2307 459 -2301
rect 463 -2307 466 -2301
rect 470 -2307 473 -2301
rect 477 -2307 480 -2301
rect 484 -2307 487 -2301
rect 491 -2307 497 -2301
rect 498 -2307 501 -2301
rect 505 -2307 511 -2301
rect 512 -2307 515 -2301
rect 519 -2307 522 -2301
rect 526 -2307 529 -2301
rect 533 -2307 536 -2301
rect 540 -2307 543 -2301
rect 547 -2307 550 -2301
rect 554 -2307 557 -2301
rect 561 -2307 564 -2301
rect 568 -2307 571 -2301
rect 575 -2307 581 -2301
rect 582 -2307 585 -2301
rect 589 -2307 592 -2301
rect 596 -2307 602 -2301
rect 603 -2307 606 -2301
rect 610 -2307 613 -2301
rect 617 -2307 620 -2301
rect 624 -2307 630 -2301
rect 631 -2307 634 -2301
rect 638 -2307 644 -2301
rect 645 -2307 648 -2301
rect 652 -2307 655 -2301
rect 659 -2307 662 -2301
rect 666 -2307 672 -2301
rect 673 -2307 679 -2301
rect 680 -2307 683 -2301
rect 687 -2307 693 -2301
rect 694 -2307 700 -2301
rect 701 -2307 707 -2301
rect 708 -2307 711 -2301
rect 715 -2307 718 -2301
rect 722 -2307 725 -2301
rect 729 -2307 732 -2301
rect 736 -2307 739 -2301
rect 743 -2307 746 -2301
rect 750 -2307 753 -2301
rect 757 -2307 763 -2301
rect 764 -2307 767 -2301
rect 771 -2307 774 -2301
rect 778 -2307 784 -2301
rect 785 -2307 788 -2301
rect 792 -2307 795 -2301
rect 799 -2307 802 -2301
rect 806 -2307 809 -2301
rect 813 -2307 816 -2301
rect 820 -2307 823 -2301
rect 827 -2307 830 -2301
rect 834 -2307 840 -2301
rect 841 -2307 844 -2301
rect 848 -2307 851 -2301
rect 855 -2307 858 -2301
rect 862 -2307 868 -2301
rect 869 -2307 875 -2301
rect 876 -2307 879 -2301
rect 883 -2307 886 -2301
rect 890 -2307 893 -2301
rect 897 -2307 900 -2301
rect 904 -2307 907 -2301
rect 911 -2307 917 -2301
rect 918 -2307 921 -2301
rect 925 -2307 928 -2301
rect 932 -2307 935 -2301
rect 939 -2307 945 -2301
rect 946 -2307 949 -2301
rect 953 -2307 956 -2301
rect 960 -2307 963 -2301
rect 967 -2307 970 -2301
rect 974 -2307 977 -2301
rect 981 -2307 984 -2301
rect 988 -2307 991 -2301
rect 995 -2307 998 -2301
rect 1002 -2307 1005 -2301
rect 1009 -2307 1012 -2301
rect 1016 -2307 1022 -2301
rect 1023 -2307 1029 -2301
rect 1030 -2307 1033 -2301
rect 1037 -2307 1043 -2301
rect 1044 -2307 1047 -2301
rect 1051 -2307 1054 -2301
rect 1058 -2307 1061 -2301
rect 1065 -2307 1068 -2301
rect 1072 -2307 1075 -2301
rect 1079 -2307 1082 -2301
rect 1086 -2307 1089 -2301
rect 1093 -2307 1096 -2301
rect 1100 -2307 1103 -2301
rect 1107 -2307 1110 -2301
rect 1114 -2307 1117 -2301
rect 1121 -2307 1124 -2301
rect 1128 -2307 1131 -2301
rect 1135 -2307 1138 -2301
rect 1142 -2307 1145 -2301
rect 1149 -2307 1152 -2301
rect 1156 -2307 1159 -2301
rect 1163 -2307 1166 -2301
rect 1170 -2307 1176 -2301
rect 1177 -2307 1180 -2301
rect 1184 -2307 1187 -2301
rect 1191 -2307 1194 -2301
rect 1198 -2307 1204 -2301
rect 1205 -2307 1208 -2301
rect 1212 -2307 1215 -2301
rect 1219 -2307 1222 -2301
rect 1226 -2307 1229 -2301
rect 1233 -2307 1236 -2301
rect 1240 -2307 1246 -2301
rect 1247 -2307 1250 -2301
rect 1254 -2307 1257 -2301
rect 1261 -2307 1264 -2301
rect 1268 -2307 1271 -2301
rect 1275 -2307 1278 -2301
rect 1282 -2307 1285 -2301
rect 1289 -2307 1292 -2301
rect 1296 -2307 1299 -2301
rect 1303 -2307 1306 -2301
rect 1310 -2307 1313 -2301
rect 1317 -2307 1320 -2301
rect 1324 -2307 1327 -2301
rect 1331 -2307 1334 -2301
rect 1338 -2307 1341 -2301
rect 1345 -2307 1348 -2301
rect 1352 -2307 1355 -2301
rect 1359 -2307 1362 -2301
rect 1366 -2307 1369 -2301
rect 1373 -2307 1376 -2301
rect 1380 -2307 1383 -2301
rect 1387 -2307 1390 -2301
rect 1394 -2307 1397 -2301
rect 1401 -2307 1404 -2301
rect 1408 -2307 1411 -2301
rect 1415 -2307 1418 -2301
rect 1422 -2307 1425 -2301
rect 1429 -2307 1432 -2301
rect 1436 -2307 1439 -2301
rect 1443 -2307 1446 -2301
rect 1450 -2307 1453 -2301
rect 1457 -2307 1460 -2301
rect 1464 -2307 1467 -2301
rect 1471 -2307 1474 -2301
rect 1478 -2307 1481 -2301
rect 1485 -2307 1488 -2301
rect 1492 -2307 1495 -2301
rect 1499 -2307 1502 -2301
rect 1506 -2307 1509 -2301
rect 1513 -2307 1516 -2301
rect 1520 -2307 1523 -2301
rect 1527 -2307 1530 -2301
rect 1534 -2307 1537 -2301
rect 1541 -2307 1544 -2301
rect 1548 -2307 1551 -2301
rect 1555 -2307 1558 -2301
rect 1562 -2307 1565 -2301
rect 1569 -2307 1572 -2301
rect 1576 -2307 1579 -2301
rect 1583 -2307 1586 -2301
rect 1590 -2307 1593 -2301
rect 1597 -2307 1600 -2301
rect 1604 -2307 1607 -2301
rect 1611 -2307 1614 -2301
rect 1618 -2307 1621 -2301
rect 1625 -2307 1628 -2301
rect 1632 -2307 1635 -2301
rect 1639 -2307 1642 -2301
rect 1646 -2307 1652 -2301
rect 1653 -2307 1659 -2301
rect 1660 -2307 1663 -2301
rect 1667 -2307 1673 -2301
rect 1674 -2307 1677 -2301
rect 1681 -2307 1684 -2301
rect 1688 -2307 1691 -2301
rect 1695 -2307 1698 -2301
rect 1 -2428 7 -2422
rect 8 -2428 14 -2422
rect 15 -2428 21 -2422
rect 22 -2428 28 -2422
rect 29 -2428 35 -2422
rect 36 -2428 42 -2422
rect 43 -2428 46 -2422
rect 50 -2428 53 -2422
rect 57 -2428 60 -2422
rect 64 -2428 67 -2422
rect 71 -2428 74 -2422
rect 78 -2428 81 -2422
rect 85 -2428 88 -2422
rect 92 -2428 95 -2422
rect 99 -2428 102 -2422
rect 106 -2428 112 -2422
rect 113 -2428 119 -2422
rect 120 -2428 123 -2422
rect 127 -2428 130 -2422
rect 134 -2428 137 -2422
rect 141 -2428 144 -2422
rect 148 -2428 151 -2422
rect 155 -2428 158 -2422
rect 162 -2428 165 -2422
rect 169 -2428 172 -2422
rect 176 -2428 179 -2422
rect 183 -2428 186 -2422
rect 190 -2428 193 -2422
rect 197 -2428 200 -2422
rect 204 -2428 207 -2422
rect 211 -2428 214 -2422
rect 218 -2428 221 -2422
rect 225 -2428 231 -2422
rect 232 -2428 235 -2422
rect 239 -2428 242 -2422
rect 246 -2428 249 -2422
rect 253 -2428 256 -2422
rect 260 -2428 263 -2422
rect 267 -2428 270 -2422
rect 274 -2428 277 -2422
rect 281 -2428 287 -2422
rect 288 -2428 291 -2422
rect 295 -2428 298 -2422
rect 302 -2428 305 -2422
rect 309 -2428 312 -2422
rect 316 -2428 319 -2422
rect 323 -2428 326 -2422
rect 330 -2428 333 -2422
rect 337 -2428 340 -2422
rect 344 -2428 347 -2422
rect 351 -2428 354 -2422
rect 358 -2428 361 -2422
rect 365 -2428 368 -2422
rect 372 -2428 375 -2422
rect 379 -2428 382 -2422
rect 386 -2428 389 -2422
rect 393 -2428 396 -2422
rect 400 -2428 406 -2422
rect 407 -2428 410 -2422
rect 414 -2428 417 -2422
rect 421 -2428 424 -2422
rect 428 -2428 431 -2422
rect 435 -2428 438 -2422
rect 442 -2428 445 -2422
rect 449 -2428 452 -2422
rect 456 -2428 459 -2422
rect 463 -2428 466 -2422
rect 470 -2428 473 -2422
rect 477 -2428 480 -2422
rect 484 -2428 487 -2422
rect 491 -2428 494 -2422
rect 498 -2428 501 -2422
rect 505 -2428 508 -2422
rect 512 -2428 515 -2422
rect 519 -2428 525 -2422
rect 526 -2428 529 -2422
rect 533 -2428 536 -2422
rect 540 -2428 543 -2422
rect 547 -2428 550 -2422
rect 554 -2428 557 -2422
rect 561 -2428 567 -2422
rect 568 -2428 571 -2422
rect 575 -2428 578 -2422
rect 582 -2428 588 -2422
rect 589 -2428 592 -2422
rect 596 -2428 599 -2422
rect 603 -2428 606 -2422
rect 610 -2428 616 -2422
rect 617 -2428 623 -2422
rect 624 -2428 627 -2422
rect 631 -2428 637 -2422
rect 638 -2428 641 -2422
rect 645 -2428 651 -2422
rect 652 -2428 655 -2422
rect 659 -2428 662 -2422
rect 666 -2428 669 -2422
rect 673 -2428 676 -2422
rect 680 -2428 686 -2422
rect 687 -2428 690 -2422
rect 694 -2428 697 -2422
rect 701 -2428 704 -2422
rect 708 -2428 711 -2422
rect 715 -2428 718 -2422
rect 722 -2428 725 -2422
rect 729 -2428 735 -2422
rect 736 -2428 742 -2422
rect 743 -2428 749 -2422
rect 750 -2428 753 -2422
rect 757 -2428 760 -2422
rect 764 -2428 767 -2422
rect 771 -2428 777 -2422
rect 778 -2428 781 -2422
rect 785 -2428 788 -2422
rect 792 -2428 795 -2422
rect 799 -2428 802 -2422
rect 806 -2428 809 -2422
rect 813 -2428 816 -2422
rect 820 -2428 823 -2422
rect 827 -2428 830 -2422
rect 834 -2428 840 -2422
rect 841 -2428 844 -2422
rect 848 -2428 854 -2422
rect 855 -2428 861 -2422
rect 862 -2428 865 -2422
rect 869 -2428 872 -2422
rect 876 -2428 879 -2422
rect 883 -2428 886 -2422
rect 890 -2428 893 -2422
rect 897 -2428 900 -2422
rect 904 -2428 907 -2422
rect 911 -2428 914 -2422
rect 918 -2428 924 -2422
rect 925 -2428 931 -2422
rect 932 -2428 935 -2422
rect 939 -2428 942 -2422
rect 946 -2428 949 -2422
rect 953 -2428 956 -2422
rect 960 -2428 963 -2422
rect 967 -2428 973 -2422
rect 974 -2428 977 -2422
rect 981 -2428 984 -2422
rect 988 -2428 991 -2422
rect 995 -2428 998 -2422
rect 1002 -2428 1005 -2422
rect 1009 -2428 1012 -2422
rect 1016 -2428 1019 -2422
rect 1023 -2428 1026 -2422
rect 1030 -2428 1033 -2422
rect 1037 -2428 1040 -2422
rect 1044 -2428 1047 -2422
rect 1051 -2428 1054 -2422
rect 1058 -2428 1061 -2422
rect 1065 -2428 1068 -2422
rect 1072 -2428 1075 -2422
rect 1079 -2428 1082 -2422
rect 1086 -2428 1089 -2422
rect 1093 -2428 1096 -2422
rect 1100 -2428 1106 -2422
rect 1107 -2428 1110 -2422
rect 1114 -2428 1117 -2422
rect 1121 -2428 1127 -2422
rect 1128 -2428 1131 -2422
rect 1135 -2428 1138 -2422
rect 1142 -2428 1145 -2422
rect 1149 -2428 1152 -2422
rect 1156 -2428 1159 -2422
rect 1163 -2428 1166 -2422
rect 1170 -2428 1173 -2422
rect 1177 -2428 1180 -2422
rect 1184 -2428 1190 -2422
rect 1191 -2428 1194 -2422
rect 1198 -2428 1204 -2422
rect 1205 -2428 1208 -2422
rect 1212 -2428 1215 -2422
rect 1219 -2428 1222 -2422
rect 1226 -2428 1229 -2422
rect 1233 -2428 1239 -2422
rect 1240 -2428 1243 -2422
rect 1247 -2428 1253 -2422
rect 1254 -2428 1257 -2422
rect 1261 -2428 1264 -2422
rect 1268 -2428 1271 -2422
rect 1275 -2428 1278 -2422
rect 1282 -2428 1285 -2422
rect 1289 -2428 1295 -2422
rect 1296 -2428 1299 -2422
rect 1303 -2428 1306 -2422
rect 1310 -2428 1313 -2422
rect 1317 -2428 1320 -2422
rect 1324 -2428 1327 -2422
rect 1331 -2428 1334 -2422
rect 1338 -2428 1341 -2422
rect 1345 -2428 1348 -2422
rect 1352 -2428 1355 -2422
rect 1359 -2428 1365 -2422
rect 1366 -2428 1369 -2422
rect 1373 -2428 1376 -2422
rect 1380 -2428 1386 -2422
rect 1387 -2428 1390 -2422
rect 1394 -2428 1397 -2422
rect 1401 -2428 1404 -2422
rect 1408 -2428 1411 -2422
rect 1415 -2428 1418 -2422
rect 1422 -2428 1425 -2422
rect 1429 -2428 1432 -2422
rect 1436 -2428 1439 -2422
rect 1443 -2428 1446 -2422
rect 1450 -2428 1453 -2422
rect 1457 -2428 1460 -2422
rect 1464 -2428 1467 -2422
rect 1471 -2428 1474 -2422
rect 1478 -2428 1481 -2422
rect 1485 -2428 1488 -2422
rect 1492 -2428 1495 -2422
rect 1499 -2428 1502 -2422
rect 1506 -2428 1509 -2422
rect 1513 -2428 1516 -2422
rect 1520 -2428 1523 -2422
rect 1527 -2428 1530 -2422
rect 1534 -2428 1537 -2422
rect 1541 -2428 1544 -2422
rect 1548 -2428 1551 -2422
rect 1555 -2428 1558 -2422
rect 1562 -2428 1565 -2422
rect 1569 -2428 1572 -2422
rect 1576 -2428 1579 -2422
rect 1583 -2428 1586 -2422
rect 1590 -2428 1593 -2422
rect 1597 -2428 1600 -2422
rect 1604 -2428 1607 -2422
rect 1611 -2428 1614 -2422
rect 1618 -2428 1624 -2422
rect 1625 -2428 1628 -2422
rect 1632 -2428 1635 -2422
rect 1639 -2428 1645 -2422
rect 1646 -2428 1652 -2422
rect 1653 -2428 1656 -2422
rect 1660 -2428 1663 -2422
rect 1 -2547 7 -2541
rect 8 -2547 14 -2541
rect 15 -2547 21 -2541
rect 22 -2547 28 -2541
rect 29 -2547 35 -2541
rect 36 -2547 42 -2541
rect 43 -2547 49 -2541
rect 50 -2547 53 -2541
rect 57 -2547 60 -2541
rect 64 -2547 67 -2541
rect 71 -2547 74 -2541
rect 78 -2547 81 -2541
rect 85 -2547 91 -2541
rect 92 -2547 95 -2541
rect 99 -2547 102 -2541
rect 106 -2547 109 -2541
rect 113 -2547 116 -2541
rect 120 -2547 123 -2541
rect 127 -2547 130 -2541
rect 134 -2547 137 -2541
rect 141 -2547 144 -2541
rect 148 -2547 151 -2541
rect 155 -2547 158 -2541
rect 162 -2547 165 -2541
rect 169 -2547 175 -2541
rect 176 -2547 179 -2541
rect 183 -2547 186 -2541
rect 190 -2547 193 -2541
rect 197 -2547 200 -2541
rect 204 -2547 207 -2541
rect 211 -2547 217 -2541
rect 218 -2547 221 -2541
rect 225 -2547 228 -2541
rect 232 -2547 235 -2541
rect 239 -2547 242 -2541
rect 246 -2547 249 -2541
rect 253 -2547 259 -2541
rect 260 -2547 263 -2541
rect 267 -2547 270 -2541
rect 274 -2547 280 -2541
rect 281 -2547 287 -2541
rect 288 -2547 294 -2541
rect 295 -2547 301 -2541
rect 302 -2547 305 -2541
rect 309 -2547 312 -2541
rect 316 -2547 319 -2541
rect 323 -2547 326 -2541
rect 330 -2547 333 -2541
rect 337 -2547 340 -2541
rect 344 -2547 347 -2541
rect 351 -2547 354 -2541
rect 358 -2547 361 -2541
rect 365 -2547 368 -2541
rect 372 -2547 375 -2541
rect 379 -2547 382 -2541
rect 386 -2547 392 -2541
rect 393 -2547 396 -2541
rect 400 -2547 403 -2541
rect 407 -2547 410 -2541
rect 414 -2547 420 -2541
rect 421 -2547 424 -2541
rect 428 -2547 431 -2541
rect 435 -2547 438 -2541
rect 442 -2547 445 -2541
rect 449 -2547 452 -2541
rect 456 -2547 459 -2541
rect 463 -2547 466 -2541
rect 470 -2547 473 -2541
rect 477 -2547 483 -2541
rect 484 -2547 487 -2541
rect 491 -2547 494 -2541
rect 498 -2547 501 -2541
rect 505 -2547 508 -2541
rect 512 -2547 515 -2541
rect 519 -2547 522 -2541
rect 526 -2547 532 -2541
rect 533 -2547 536 -2541
rect 540 -2547 546 -2541
rect 547 -2547 550 -2541
rect 554 -2547 557 -2541
rect 561 -2547 567 -2541
rect 568 -2547 574 -2541
rect 575 -2547 578 -2541
rect 582 -2547 585 -2541
rect 589 -2547 592 -2541
rect 596 -2547 602 -2541
rect 603 -2547 606 -2541
rect 610 -2547 613 -2541
rect 617 -2547 620 -2541
rect 624 -2547 627 -2541
rect 631 -2547 634 -2541
rect 638 -2547 641 -2541
rect 645 -2547 648 -2541
rect 652 -2547 655 -2541
rect 659 -2547 662 -2541
rect 666 -2547 672 -2541
rect 673 -2547 676 -2541
rect 680 -2547 683 -2541
rect 687 -2547 690 -2541
rect 694 -2547 697 -2541
rect 701 -2547 704 -2541
rect 708 -2547 711 -2541
rect 715 -2547 718 -2541
rect 722 -2547 725 -2541
rect 729 -2547 735 -2541
rect 736 -2547 742 -2541
rect 743 -2547 749 -2541
rect 750 -2547 756 -2541
rect 757 -2547 760 -2541
rect 764 -2547 767 -2541
rect 771 -2547 774 -2541
rect 778 -2547 781 -2541
rect 785 -2547 791 -2541
rect 792 -2547 795 -2541
rect 799 -2547 805 -2541
rect 806 -2547 812 -2541
rect 813 -2547 816 -2541
rect 820 -2547 823 -2541
rect 827 -2547 833 -2541
rect 834 -2547 837 -2541
rect 841 -2547 844 -2541
rect 848 -2547 851 -2541
rect 855 -2547 858 -2541
rect 862 -2547 865 -2541
rect 869 -2547 872 -2541
rect 876 -2547 879 -2541
rect 883 -2547 886 -2541
rect 890 -2547 893 -2541
rect 897 -2547 903 -2541
rect 904 -2547 907 -2541
rect 911 -2547 914 -2541
rect 918 -2547 921 -2541
rect 925 -2547 928 -2541
rect 932 -2547 935 -2541
rect 939 -2547 942 -2541
rect 946 -2547 949 -2541
rect 953 -2547 956 -2541
rect 960 -2547 963 -2541
rect 967 -2547 970 -2541
rect 974 -2547 977 -2541
rect 981 -2547 984 -2541
rect 988 -2547 991 -2541
rect 995 -2547 1001 -2541
rect 1002 -2547 1005 -2541
rect 1009 -2547 1015 -2541
rect 1016 -2547 1019 -2541
rect 1023 -2547 1029 -2541
rect 1030 -2547 1033 -2541
rect 1037 -2547 1040 -2541
rect 1044 -2547 1047 -2541
rect 1051 -2547 1054 -2541
rect 1058 -2547 1061 -2541
rect 1065 -2547 1068 -2541
rect 1072 -2547 1075 -2541
rect 1079 -2547 1082 -2541
rect 1086 -2547 1089 -2541
rect 1093 -2547 1096 -2541
rect 1100 -2547 1103 -2541
rect 1107 -2547 1110 -2541
rect 1114 -2547 1117 -2541
rect 1121 -2547 1124 -2541
rect 1128 -2547 1131 -2541
rect 1135 -2547 1138 -2541
rect 1142 -2547 1148 -2541
rect 1149 -2547 1152 -2541
rect 1156 -2547 1159 -2541
rect 1163 -2547 1166 -2541
rect 1170 -2547 1173 -2541
rect 1177 -2547 1180 -2541
rect 1184 -2547 1187 -2541
rect 1191 -2547 1194 -2541
rect 1198 -2547 1201 -2541
rect 1205 -2547 1208 -2541
rect 1212 -2547 1215 -2541
rect 1219 -2547 1222 -2541
rect 1226 -2547 1229 -2541
rect 1233 -2547 1236 -2541
rect 1240 -2547 1243 -2541
rect 1247 -2547 1253 -2541
rect 1254 -2547 1257 -2541
rect 1261 -2547 1264 -2541
rect 1268 -2547 1271 -2541
rect 1275 -2547 1278 -2541
rect 1282 -2547 1285 -2541
rect 1289 -2547 1292 -2541
rect 1296 -2547 1299 -2541
rect 1303 -2547 1306 -2541
rect 1310 -2547 1313 -2541
rect 1317 -2547 1320 -2541
rect 1324 -2547 1327 -2541
rect 1331 -2547 1334 -2541
rect 1338 -2547 1341 -2541
rect 1345 -2547 1348 -2541
rect 1352 -2547 1355 -2541
rect 1359 -2547 1362 -2541
rect 1366 -2547 1369 -2541
rect 1373 -2547 1376 -2541
rect 1380 -2547 1383 -2541
rect 1387 -2547 1390 -2541
rect 1394 -2547 1397 -2541
rect 1401 -2547 1407 -2541
rect 1408 -2547 1411 -2541
rect 1415 -2547 1418 -2541
rect 1422 -2547 1425 -2541
rect 1429 -2547 1432 -2541
rect 1436 -2547 1439 -2541
rect 1443 -2547 1446 -2541
rect 1450 -2547 1453 -2541
rect 1457 -2547 1460 -2541
rect 1464 -2547 1467 -2541
rect 1471 -2547 1474 -2541
rect 1478 -2547 1481 -2541
rect 1485 -2547 1488 -2541
rect 1492 -2547 1495 -2541
rect 1499 -2547 1502 -2541
rect 1506 -2547 1509 -2541
rect 1513 -2547 1516 -2541
rect 1520 -2547 1523 -2541
rect 1527 -2547 1530 -2541
rect 1534 -2547 1537 -2541
rect 1541 -2547 1544 -2541
rect 1548 -2547 1551 -2541
rect 1555 -2547 1558 -2541
rect 1562 -2547 1565 -2541
rect 1569 -2547 1572 -2541
rect 1576 -2547 1579 -2541
rect 1583 -2547 1589 -2541
rect 1590 -2547 1593 -2541
rect 1597 -2547 1600 -2541
rect 1604 -2547 1607 -2541
rect 1611 -2547 1617 -2541
rect 1639 -2547 1642 -2541
rect 1 -2676 7 -2670
rect 8 -2676 14 -2670
rect 15 -2676 21 -2670
rect 22 -2676 28 -2670
rect 29 -2676 35 -2670
rect 36 -2676 42 -2670
rect 43 -2676 46 -2670
rect 50 -2676 53 -2670
rect 57 -2676 60 -2670
rect 64 -2676 67 -2670
rect 71 -2676 74 -2670
rect 78 -2676 81 -2670
rect 85 -2676 88 -2670
rect 92 -2676 95 -2670
rect 99 -2676 102 -2670
rect 106 -2676 109 -2670
rect 113 -2676 116 -2670
rect 120 -2676 123 -2670
rect 127 -2676 133 -2670
rect 134 -2676 137 -2670
rect 141 -2676 144 -2670
rect 148 -2676 154 -2670
rect 155 -2676 161 -2670
rect 162 -2676 165 -2670
rect 169 -2676 172 -2670
rect 176 -2676 182 -2670
rect 183 -2676 186 -2670
rect 190 -2676 193 -2670
rect 197 -2676 203 -2670
rect 204 -2676 210 -2670
rect 211 -2676 214 -2670
rect 218 -2676 221 -2670
rect 225 -2676 228 -2670
rect 232 -2676 238 -2670
rect 239 -2676 242 -2670
rect 246 -2676 252 -2670
rect 253 -2676 256 -2670
rect 260 -2676 266 -2670
rect 267 -2676 270 -2670
rect 274 -2676 277 -2670
rect 281 -2676 284 -2670
rect 288 -2676 291 -2670
rect 295 -2676 298 -2670
rect 302 -2676 305 -2670
rect 309 -2676 312 -2670
rect 316 -2676 319 -2670
rect 323 -2676 326 -2670
rect 330 -2676 333 -2670
rect 337 -2676 340 -2670
rect 344 -2676 347 -2670
rect 351 -2676 354 -2670
rect 358 -2676 361 -2670
rect 365 -2676 368 -2670
rect 372 -2676 378 -2670
rect 379 -2676 382 -2670
rect 386 -2676 389 -2670
rect 393 -2676 399 -2670
rect 400 -2676 403 -2670
rect 407 -2676 410 -2670
rect 414 -2676 417 -2670
rect 421 -2676 427 -2670
rect 428 -2676 431 -2670
rect 435 -2676 438 -2670
rect 442 -2676 445 -2670
rect 449 -2676 452 -2670
rect 456 -2676 459 -2670
rect 463 -2676 466 -2670
rect 470 -2676 473 -2670
rect 477 -2676 480 -2670
rect 484 -2676 487 -2670
rect 491 -2676 494 -2670
rect 498 -2676 504 -2670
rect 505 -2676 508 -2670
rect 512 -2676 515 -2670
rect 519 -2676 522 -2670
rect 526 -2676 529 -2670
rect 533 -2676 536 -2670
rect 540 -2676 543 -2670
rect 547 -2676 550 -2670
rect 554 -2676 557 -2670
rect 561 -2676 564 -2670
rect 568 -2676 571 -2670
rect 575 -2676 578 -2670
rect 582 -2676 585 -2670
rect 589 -2676 592 -2670
rect 596 -2676 599 -2670
rect 603 -2676 606 -2670
rect 610 -2676 616 -2670
rect 617 -2676 620 -2670
rect 624 -2676 627 -2670
rect 631 -2676 634 -2670
rect 638 -2676 641 -2670
rect 645 -2676 651 -2670
rect 652 -2676 658 -2670
rect 659 -2676 662 -2670
rect 666 -2676 669 -2670
rect 673 -2676 676 -2670
rect 680 -2676 683 -2670
rect 687 -2676 690 -2670
rect 694 -2676 697 -2670
rect 701 -2676 704 -2670
rect 708 -2676 711 -2670
rect 715 -2676 721 -2670
rect 722 -2676 725 -2670
rect 729 -2676 735 -2670
rect 736 -2676 739 -2670
rect 743 -2676 746 -2670
rect 750 -2676 753 -2670
rect 757 -2676 760 -2670
rect 764 -2676 767 -2670
rect 771 -2676 774 -2670
rect 778 -2676 781 -2670
rect 785 -2676 788 -2670
rect 792 -2676 795 -2670
rect 799 -2676 805 -2670
rect 806 -2676 809 -2670
rect 813 -2676 816 -2670
rect 820 -2676 823 -2670
rect 827 -2676 830 -2670
rect 834 -2676 837 -2670
rect 841 -2676 844 -2670
rect 848 -2676 851 -2670
rect 855 -2676 861 -2670
rect 862 -2676 865 -2670
rect 869 -2676 872 -2670
rect 876 -2676 882 -2670
rect 883 -2676 889 -2670
rect 890 -2676 893 -2670
rect 897 -2676 903 -2670
rect 904 -2676 910 -2670
rect 911 -2676 914 -2670
rect 918 -2676 921 -2670
rect 925 -2676 928 -2670
rect 932 -2676 935 -2670
rect 939 -2676 942 -2670
rect 946 -2676 952 -2670
rect 953 -2676 959 -2670
rect 960 -2676 963 -2670
rect 967 -2676 973 -2670
rect 974 -2676 980 -2670
rect 981 -2676 984 -2670
rect 988 -2676 991 -2670
rect 995 -2676 998 -2670
rect 1002 -2676 1005 -2670
rect 1009 -2676 1012 -2670
rect 1016 -2676 1019 -2670
rect 1023 -2676 1029 -2670
rect 1030 -2676 1033 -2670
rect 1037 -2676 1040 -2670
rect 1044 -2676 1047 -2670
rect 1051 -2676 1054 -2670
rect 1058 -2676 1061 -2670
rect 1065 -2676 1068 -2670
rect 1072 -2676 1075 -2670
rect 1079 -2676 1082 -2670
rect 1086 -2676 1092 -2670
rect 1093 -2676 1096 -2670
rect 1100 -2676 1103 -2670
rect 1107 -2676 1110 -2670
rect 1114 -2676 1117 -2670
rect 1121 -2676 1124 -2670
rect 1128 -2676 1131 -2670
rect 1135 -2676 1138 -2670
rect 1142 -2676 1145 -2670
rect 1149 -2676 1155 -2670
rect 1156 -2676 1159 -2670
rect 1163 -2676 1166 -2670
rect 1170 -2676 1173 -2670
rect 1177 -2676 1180 -2670
rect 1184 -2676 1190 -2670
rect 1191 -2676 1194 -2670
rect 1198 -2676 1201 -2670
rect 1205 -2676 1208 -2670
rect 1212 -2676 1215 -2670
rect 1219 -2676 1222 -2670
rect 1226 -2676 1229 -2670
rect 1233 -2676 1236 -2670
rect 1240 -2676 1243 -2670
rect 1247 -2676 1250 -2670
rect 1254 -2676 1257 -2670
rect 1261 -2676 1264 -2670
rect 1268 -2676 1271 -2670
rect 1275 -2676 1278 -2670
rect 1282 -2676 1285 -2670
rect 1289 -2676 1292 -2670
rect 1296 -2676 1299 -2670
rect 1303 -2676 1306 -2670
rect 1310 -2676 1313 -2670
rect 1317 -2676 1320 -2670
rect 1324 -2676 1327 -2670
rect 1331 -2676 1334 -2670
rect 1338 -2676 1341 -2670
rect 1345 -2676 1348 -2670
rect 1352 -2676 1355 -2670
rect 1359 -2676 1362 -2670
rect 1366 -2676 1369 -2670
rect 1373 -2676 1376 -2670
rect 1380 -2676 1383 -2670
rect 1387 -2676 1390 -2670
rect 1394 -2676 1397 -2670
rect 1401 -2676 1404 -2670
rect 1408 -2676 1411 -2670
rect 1415 -2676 1418 -2670
rect 1422 -2676 1425 -2670
rect 1429 -2676 1432 -2670
rect 1436 -2676 1439 -2670
rect 1443 -2676 1446 -2670
rect 1450 -2676 1453 -2670
rect 1457 -2676 1460 -2670
rect 1464 -2676 1467 -2670
rect 1471 -2676 1474 -2670
rect 1478 -2676 1481 -2670
rect 1485 -2676 1488 -2670
rect 1492 -2676 1495 -2670
rect 1499 -2676 1502 -2670
rect 1506 -2676 1509 -2670
rect 1513 -2676 1516 -2670
rect 1520 -2676 1523 -2670
rect 1527 -2676 1530 -2670
rect 1534 -2676 1537 -2670
rect 1541 -2676 1544 -2670
rect 1548 -2676 1551 -2670
rect 1555 -2676 1558 -2670
rect 1562 -2676 1565 -2670
rect 1569 -2676 1572 -2670
rect 1576 -2676 1579 -2670
rect 1583 -2676 1586 -2670
rect 1590 -2676 1593 -2670
rect 1597 -2676 1600 -2670
rect 1604 -2676 1607 -2670
rect 1611 -2676 1614 -2670
rect 1618 -2676 1621 -2670
rect 1625 -2676 1631 -2670
rect 1632 -2676 1638 -2670
rect 1 -2789 7 -2783
rect 8 -2789 14 -2783
rect 15 -2789 21 -2783
rect 22 -2789 28 -2783
rect 29 -2789 35 -2783
rect 36 -2789 42 -2783
rect 43 -2789 46 -2783
rect 50 -2789 56 -2783
rect 57 -2789 60 -2783
rect 64 -2789 67 -2783
rect 71 -2789 74 -2783
rect 78 -2789 81 -2783
rect 85 -2789 88 -2783
rect 92 -2789 95 -2783
rect 99 -2789 102 -2783
rect 106 -2789 112 -2783
rect 113 -2789 116 -2783
rect 120 -2789 126 -2783
rect 127 -2789 133 -2783
rect 134 -2789 140 -2783
rect 141 -2789 144 -2783
rect 148 -2789 151 -2783
rect 155 -2789 161 -2783
rect 162 -2789 165 -2783
rect 169 -2789 172 -2783
rect 176 -2789 179 -2783
rect 183 -2789 186 -2783
rect 190 -2789 193 -2783
rect 197 -2789 200 -2783
rect 204 -2789 207 -2783
rect 211 -2789 217 -2783
rect 218 -2789 221 -2783
rect 225 -2789 228 -2783
rect 232 -2789 238 -2783
rect 239 -2789 242 -2783
rect 246 -2789 249 -2783
rect 253 -2789 256 -2783
rect 260 -2789 266 -2783
rect 267 -2789 270 -2783
rect 274 -2789 277 -2783
rect 281 -2789 287 -2783
rect 288 -2789 294 -2783
rect 295 -2789 298 -2783
rect 302 -2789 305 -2783
rect 309 -2789 312 -2783
rect 316 -2789 319 -2783
rect 323 -2789 326 -2783
rect 330 -2789 333 -2783
rect 337 -2789 340 -2783
rect 344 -2789 347 -2783
rect 351 -2789 354 -2783
rect 358 -2789 361 -2783
rect 365 -2789 368 -2783
rect 372 -2789 375 -2783
rect 379 -2789 382 -2783
rect 386 -2789 389 -2783
rect 393 -2789 396 -2783
rect 400 -2789 403 -2783
rect 407 -2789 410 -2783
rect 414 -2789 417 -2783
rect 421 -2789 424 -2783
rect 428 -2789 431 -2783
rect 435 -2789 438 -2783
rect 442 -2789 448 -2783
rect 449 -2789 452 -2783
rect 456 -2789 459 -2783
rect 463 -2789 466 -2783
rect 470 -2789 473 -2783
rect 477 -2789 483 -2783
rect 484 -2789 487 -2783
rect 491 -2789 494 -2783
rect 498 -2789 501 -2783
rect 505 -2789 508 -2783
rect 512 -2789 515 -2783
rect 519 -2789 522 -2783
rect 526 -2789 529 -2783
rect 533 -2789 536 -2783
rect 540 -2789 543 -2783
rect 547 -2789 550 -2783
rect 554 -2789 557 -2783
rect 561 -2789 567 -2783
rect 568 -2789 571 -2783
rect 575 -2789 578 -2783
rect 582 -2789 585 -2783
rect 589 -2789 595 -2783
rect 596 -2789 599 -2783
rect 603 -2789 606 -2783
rect 610 -2789 613 -2783
rect 617 -2789 620 -2783
rect 624 -2789 627 -2783
rect 631 -2789 634 -2783
rect 638 -2789 641 -2783
rect 645 -2789 648 -2783
rect 652 -2789 655 -2783
rect 659 -2789 665 -2783
rect 666 -2789 672 -2783
rect 673 -2789 679 -2783
rect 680 -2789 683 -2783
rect 687 -2789 693 -2783
rect 694 -2789 697 -2783
rect 701 -2789 704 -2783
rect 708 -2789 711 -2783
rect 715 -2789 718 -2783
rect 722 -2789 725 -2783
rect 729 -2789 732 -2783
rect 736 -2789 739 -2783
rect 743 -2789 749 -2783
rect 750 -2789 753 -2783
rect 757 -2789 763 -2783
rect 764 -2789 767 -2783
rect 771 -2789 774 -2783
rect 778 -2789 784 -2783
rect 785 -2789 791 -2783
rect 792 -2789 795 -2783
rect 799 -2789 802 -2783
rect 806 -2789 812 -2783
rect 813 -2789 819 -2783
rect 820 -2789 823 -2783
rect 827 -2789 830 -2783
rect 834 -2789 837 -2783
rect 841 -2789 847 -2783
rect 848 -2789 851 -2783
rect 855 -2789 858 -2783
rect 862 -2789 865 -2783
rect 869 -2789 872 -2783
rect 876 -2789 882 -2783
rect 883 -2789 886 -2783
rect 890 -2789 893 -2783
rect 897 -2789 900 -2783
rect 904 -2789 910 -2783
rect 911 -2789 914 -2783
rect 918 -2789 921 -2783
rect 925 -2789 928 -2783
rect 932 -2789 935 -2783
rect 939 -2789 942 -2783
rect 946 -2789 949 -2783
rect 953 -2789 956 -2783
rect 960 -2789 963 -2783
rect 967 -2789 970 -2783
rect 974 -2789 977 -2783
rect 981 -2789 984 -2783
rect 988 -2789 991 -2783
rect 995 -2789 998 -2783
rect 1002 -2789 1008 -2783
rect 1009 -2789 1012 -2783
rect 1016 -2789 1019 -2783
rect 1023 -2789 1026 -2783
rect 1030 -2789 1033 -2783
rect 1037 -2789 1040 -2783
rect 1044 -2789 1047 -2783
rect 1051 -2789 1054 -2783
rect 1058 -2789 1061 -2783
rect 1065 -2789 1068 -2783
rect 1072 -2789 1075 -2783
rect 1079 -2789 1082 -2783
rect 1086 -2789 1089 -2783
rect 1093 -2789 1096 -2783
rect 1100 -2789 1103 -2783
rect 1107 -2789 1110 -2783
rect 1114 -2789 1117 -2783
rect 1121 -2789 1124 -2783
rect 1128 -2789 1131 -2783
rect 1135 -2789 1138 -2783
rect 1142 -2789 1145 -2783
rect 1149 -2789 1152 -2783
rect 1156 -2789 1162 -2783
rect 1163 -2789 1166 -2783
rect 1170 -2789 1173 -2783
rect 1177 -2789 1180 -2783
rect 1184 -2789 1190 -2783
rect 1191 -2789 1194 -2783
rect 1198 -2789 1201 -2783
rect 1205 -2789 1208 -2783
rect 1212 -2789 1215 -2783
rect 1219 -2789 1222 -2783
rect 1226 -2789 1229 -2783
rect 1233 -2789 1236 -2783
rect 1240 -2789 1243 -2783
rect 1247 -2789 1250 -2783
rect 1254 -2789 1257 -2783
rect 1261 -2789 1264 -2783
rect 1268 -2789 1271 -2783
rect 1275 -2789 1278 -2783
rect 1282 -2789 1285 -2783
rect 1289 -2789 1292 -2783
rect 1296 -2789 1302 -2783
rect 1303 -2789 1306 -2783
rect 1310 -2789 1313 -2783
rect 1317 -2789 1320 -2783
rect 1324 -2789 1327 -2783
rect 1331 -2789 1334 -2783
rect 1338 -2789 1341 -2783
rect 1345 -2789 1348 -2783
rect 1352 -2789 1355 -2783
rect 1359 -2789 1362 -2783
rect 1366 -2789 1369 -2783
rect 1373 -2789 1376 -2783
rect 1380 -2789 1383 -2783
rect 1387 -2789 1390 -2783
rect 1394 -2789 1397 -2783
rect 1401 -2789 1404 -2783
rect 1408 -2789 1411 -2783
rect 1415 -2789 1418 -2783
rect 1422 -2789 1425 -2783
rect 1429 -2789 1432 -2783
rect 1436 -2789 1439 -2783
rect 1443 -2789 1446 -2783
rect 1450 -2789 1453 -2783
rect 1457 -2789 1460 -2783
rect 1464 -2789 1467 -2783
rect 1471 -2789 1474 -2783
rect 1478 -2789 1481 -2783
rect 1485 -2789 1488 -2783
rect 1492 -2789 1495 -2783
rect 1499 -2789 1502 -2783
rect 1506 -2789 1509 -2783
rect 1513 -2789 1516 -2783
rect 1520 -2789 1526 -2783
rect 1 -2914 7 -2908
rect 8 -2914 14 -2908
rect 15 -2914 21 -2908
rect 22 -2914 28 -2908
rect 29 -2914 35 -2908
rect 36 -2914 42 -2908
rect 43 -2914 49 -2908
rect 50 -2914 56 -2908
rect 57 -2914 63 -2908
rect 64 -2914 70 -2908
rect 71 -2914 74 -2908
rect 78 -2914 81 -2908
rect 85 -2914 88 -2908
rect 92 -2914 95 -2908
rect 99 -2914 105 -2908
rect 106 -2914 109 -2908
rect 113 -2914 116 -2908
rect 120 -2914 126 -2908
rect 127 -2914 130 -2908
rect 134 -2914 137 -2908
rect 141 -2914 147 -2908
rect 148 -2914 151 -2908
rect 155 -2914 158 -2908
rect 162 -2914 165 -2908
rect 169 -2914 172 -2908
rect 176 -2914 179 -2908
rect 183 -2914 186 -2908
rect 190 -2914 193 -2908
rect 197 -2914 200 -2908
rect 204 -2914 210 -2908
rect 211 -2914 214 -2908
rect 218 -2914 221 -2908
rect 225 -2914 231 -2908
rect 232 -2914 235 -2908
rect 239 -2914 242 -2908
rect 246 -2914 252 -2908
rect 253 -2914 256 -2908
rect 260 -2914 263 -2908
rect 267 -2914 270 -2908
rect 274 -2914 280 -2908
rect 281 -2914 287 -2908
rect 288 -2914 294 -2908
rect 295 -2914 298 -2908
rect 302 -2914 305 -2908
rect 309 -2914 312 -2908
rect 316 -2914 319 -2908
rect 323 -2914 326 -2908
rect 330 -2914 333 -2908
rect 337 -2914 340 -2908
rect 344 -2914 347 -2908
rect 351 -2914 354 -2908
rect 358 -2914 361 -2908
rect 365 -2914 368 -2908
rect 372 -2914 375 -2908
rect 379 -2914 382 -2908
rect 386 -2914 389 -2908
rect 393 -2914 396 -2908
rect 400 -2914 403 -2908
rect 407 -2914 410 -2908
rect 414 -2914 417 -2908
rect 421 -2914 424 -2908
rect 428 -2914 431 -2908
rect 435 -2914 438 -2908
rect 442 -2914 445 -2908
rect 449 -2914 452 -2908
rect 456 -2914 459 -2908
rect 463 -2914 466 -2908
rect 470 -2914 473 -2908
rect 477 -2914 480 -2908
rect 484 -2914 487 -2908
rect 491 -2914 497 -2908
rect 498 -2914 501 -2908
rect 505 -2914 508 -2908
rect 512 -2914 515 -2908
rect 519 -2914 522 -2908
rect 526 -2914 529 -2908
rect 533 -2914 536 -2908
rect 540 -2914 543 -2908
rect 547 -2914 550 -2908
rect 554 -2914 560 -2908
rect 561 -2914 564 -2908
rect 568 -2914 571 -2908
rect 575 -2914 578 -2908
rect 582 -2914 588 -2908
rect 589 -2914 592 -2908
rect 596 -2914 599 -2908
rect 603 -2914 606 -2908
rect 610 -2914 613 -2908
rect 617 -2914 620 -2908
rect 624 -2914 627 -2908
rect 631 -2914 634 -2908
rect 638 -2914 644 -2908
rect 645 -2914 648 -2908
rect 652 -2914 655 -2908
rect 659 -2914 665 -2908
rect 666 -2914 669 -2908
rect 673 -2914 676 -2908
rect 680 -2914 683 -2908
rect 687 -2914 690 -2908
rect 694 -2914 697 -2908
rect 701 -2914 707 -2908
rect 708 -2914 711 -2908
rect 715 -2914 718 -2908
rect 722 -2914 725 -2908
rect 729 -2914 732 -2908
rect 736 -2914 739 -2908
rect 743 -2914 749 -2908
rect 750 -2914 753 -2908
rect 757 -2914 763 -2908
rect 764 -2914 767 -2908
rect 771 -2914 774 -2908
rect 778 -2914 781 -2908
rect 785 -2914 788 -2908
rect 792 -2914 795 -2908
rect 799 -2914 802 -2908
rect 806 -2914 809 -2908
rect 813 -2914 816 -2908
rect 820 -2914 826 -2908
rect 827 -2914 830 -2908
rect 834 -2914 840 -2908
rect 841 -2914 847 -2908
rect 848 -2914 851 -2908
rect 855 -2914 858 -2908
rect 862 -2914 868 -2908
rect 869 -2914 872 -2908
rect 876 -2914 879 -2908
rect 883 -2914 886 -2908
rect 890 -2914 893 -2908
rect 897 -2914 900 -2908
rect 904 -2914 907 -2908
rect 911 -2914 917 -2908
rect 918 -2914 924 -2908
rect 925 -2914 928 -2908
rect 932 -2914 935 -2908
rect 939 -2914 942 -2908
rect 946 -2914 952 -2908
rect 953 -2914 959 -2908
rect 960 -2914 963 -2908
rect 967 -2914 970 -2908
rect 974 -2914 977 -2908
rect 981 -2914 984 -2908
rect 988 -2914 991 -2908
rect 995 -2914 998 -2908
rect 1002 -2914 1005 -2908
rect 1009 -2914 1012 -2908
rect 1016 -2914 1022 -2908
rect 1023 -2914 1026 -2908
rect 1030 -2914 1033 -2908
rect 1037 -2914 1040 -2908
rect 1044 -2914 1047 -2908
rect 1051 -2914 1054 -2908
rect 1058 -2914 1061 -2908
rect 1065 -2914 1068 -2908
rect 1072 -2914 1075 -2908
rect 1079 -2914 1082 -2908
rect 1086 -2914 1089 -2908
rect 1093 -2914 1099 -2908
rect 1100 -2914 1103 -2908
rect 1107 -2914 1110 -2908
rect 1114 -2914 1117 -2908
rect 1121 -2914 1124 -2908
rect 1128 -2914 1131 -2908
rect 1135 -2914 1138 -2908
rect 1142 -2914 1145 -2908
rect 1149 -2914 1152 -2908
rect 1156 -2914 1159 -2908
rect 1163 -2914 1166 -2908
rect 1170 -2914 1173 -2908
rect 1177 -2914 1180 -2908
rect 1184 -2914 1187 -2908
rect 1191 -2914 1194 -2908
rect 1198 -2914 1201 -2908
rect 1205 -2914 1208 -2908
rect 1212 -2914 1215 -2908
rect 1219 -2914 1222 -2908
rect 1226 -2914 1229 -2908
rect 1233 -2914 1236 -2908
rect 1240 -2914 1243 -2908
rect 1247 -2914 1250 -2908
rect 1254 -2914 1257 -2908
rect 1261 -2914 1264 -2908
rect 1268 -2914 1271 -2908
rect 1275 -2914 1278 -2908
rect 1282 -2914 1285 -2908
rect 1289 -2914 1292 -2908
rect 1296 -2914 1299 -2908
rect 1303 -2914 1306 -2908
rect 1310 -2914 1313 -2908
rect 1317 -2914 1320 -2908
rect 1324 -2914 1327 -2908
rect 1331 -2914 1334 -2908
rect 1338 -2914 1341 -2908
rect 1345 -2914 1348 -2908
rect 1352 -2914 1355 -2908
rect 1359 -2914 1365 -2908
rect 1366 -2914 1369 -2908
rect 1373 -2914 1376 -2908
rect 1380 -2914 1383 -2908
rect 1387 -2914 1390 -2908
rect 1394 -2914 1397 -2908
rect 1401 -2914 1404 -2908
rect 1408 -2914 1411 -2908
rect 1415 -2914 1418 -2908
rect 1422 -2914 1425 -2908
rect 1429 -2914 1432 -2908
rect 1 -3033 7 -3027
rect 8 -3033 14 -3027
rect 15 -3033 21 -3027
rect 22 -3033 28 -3027
rect 29 -3033 35 -3027
rect 36 -3033 42 -3027
rect 43 -3033 49 -3027
rect 50 -3033 56 -3027
rect 57 -3033 63 -3027
rect 64 -3033 70 -3027
rect 71 -3033 77 -3027
rect 78 -3033 84 -3027
rect 85 -3033 88 -3027
rect 92 -3033 95 -3027
rect 99 -3033 102 -3027
rect 106 -3033 109 -3027
rect 113 -3033 116 -3027
rect 120 -3033 123 -3027
rect 127 -3033 130 -3027
rect 134 -3033 137 -3027
rect 141 -3033 144 -3027
rect 148 -3033 154 -3027
rect 155 -3033 158 -3027
rect 162 -3033 168 -3027
rect 169 -3033 172 -3027
rect 176 -3033 179 -3027
rect 183 -3033 186 -3027
rect 190 -3033 193 -3027
rect 197 -3033 200 -3027
rect 204 -3033 210 -3027
rect 211 -3033 214 -3027
rect 218 -3033 224 -3027
rect 225 -3033 228 -3027
rect 232 -3033 235 -3027
rect 239 -3033 242 -3027
rect 246 -3033 252 -3027
rect 253 -3033 256 -3027
rect 260 -3033 266 -3027
rect 267 -3033 270 -3027
rect 274 -3033 277 -3027
rect 281 -3033 284 -3027
rect 288 -3033 291 -3027
rect 295 -3033 298 -3027
rect 302 -3033 305 -3027
rect 309 -3033 312 -3027
rect 316 -3033 319 -3027
rect 323 -3033 326 -3027
rect 330 -3033 333 -3027
rect 337 -3033 340 -3027
rect 344 -3033 347 -3027
rect 351 -3033 354 -3027
rect 358 -3033 361 -3027
rect 365 -3033 368 -3027
rect 372 -3033 375 -3027
rect 379 -3033 382 -3027
rect 386 -3033 389 -3027
rect 393 -3033 396 -3027
rect 400 -3033 403 -3027
rect 407 -3033 413 -3027
rect 414 -3033 417 -3027
rect 421 -3033 424 -3027
rect 428 -3033 431 -3027
rect 435 -3033 438 -3027
rect 442 -3033 445 -3027
rect 449 -3033 452 -3027
rect 456 -3033 459 -3027
rect 463 -3033 466 -3027
rect 470 -3033 473 -3027
rect 477 -3033 480 -3027
rect 484 -3033 487 -3027
rect 491 -3033 494 -3027
rect 498 -3033 501 -3027
rect 505 -3033 511 -3027
rect 512 -3033 515 -3027
rect 519 -3033 522 -3027
rect 526 -3033 529 -3027
rect 533 -3033 536 -3027
rect 540 -3033 543 -3027
rect 547 -3033 550 -3027
rect 554 -3033 557 -3027
rect 561 -3033 564 -3027
rect 568 -3033 571 -3027
rect 575 -3033 578 -3027
rect 582 -3033 585 -3027
rect 589 -3033 592 -3027
rect 596 -3033 599 -3027
rect 603 -3033 606 -3027
rect 610 -3033 613 -3027
rect 617 -3033 620 -3027
rect 624 -3033 627 -3027
rect 631 -3033 637 -3027
rect 638 -3033 641 -3027
rect 645 -3033 651 -3027
rect 652 -3033 655 -3027
rect 659 -3033 665 -3027
rect 666 -3033 669 -3027
rect 673 -3033 676 -3027
rect 680 -3033 683 -3027
rect 687 -3033 693 -3027
rect 694 -3033 700 -3027
rect 701 -3033 704 -3027
rect 708 -3033 711 -3027
rect 715 -3033 718 -3027
rect 722 -3033 725 -3027
rect 729 -3033 732 -3027
rect 736 -3033 739 -3027
rect 743 -3033 746 -3027
rect 750 -3033 756 -3027
rect 757 -3033 760 -3027
rect 764 -3033 770 -3027
rect 771 -3033 774 -3027
rect 778 -3033 781 -3027
rect 785 -3033 791 -3027
rect 792 -3033 795 -3027
rect 799 -3033 802 -3027
rect 806 -3033 809 -3027
rect 813 -3033 816 -3027
rect 820 -3033 823 -3027
rect 827 -3033 830 -3027
rect 834 -3033 840 -3027
rect 841 -3033 844 -3027
rect 848 -3033 851 -3027
rect 855 -3033 858 -3027
rect 862 -3033 868 -3027
rect 869 -3033 875 -3027
rect 876 -3033 879 -3027
rect 883 -3033 889 -3027
rect 890 -3033 893 -3027
rect 897 -3033 900 -3027
rect 904 -3033 907 -3027
rect 911 -3033 917 -3027
rect 918 -3033 924 -3027
rect 925 -3033 928 -3027
rect 932 -3033 935 -3027
rect 939 -3033 942 -3027
rect 946 -3033 949 -3027
rect 953 -3033 956 -3027
rect 960 -3033 963 -3027
rect 967 -3033 970 -3027
rect 974 -3033 977 -3027
rect 981 -3033 984 -3027
rect 988 -3033 991 -3027
rect 995 -3033 998 -3027
rect 1002 -3033 1005 -3027
rect 1009 -3033 1012 -3027
rect 1016 -3033 1022 -3027
rect 1023 -3033 1026 -3027
rect 1030 -3033 1033 -3027
rect 1037 -3033 1040 -3027
rect 1044 -3033 1047 -3027
rect 1051 -3033 1054 -3027
rect 1058 -3033 1061 -3027
rect 1065 -3033 1068 -3027
rect 1072 -3033 1078 -3027
rect 1079 -3033 1082 -3027
rect 1086 -3033 1089 -3027
rect 1093 -3033 1096 -3027
rect 1100 -3033 1103 -3027
rect 1107 -3033 1110 -3027
rect 1114 -3033 1117 -3027
rect 1121 -3033 1124 -3027
rect 1128 -3033 1131 -3027
rect 1135 -3033 1138 -3027
rect 1142 -3033 1145 -3027
rect 1149 -3033 1155 -3027
rect 1156 -3033 1159 -3027
rect 1163 -3033 1166 -3027
rect 1170 -3033 1173 -3027
rect 1177 -3033 1180 -3027
rect 1184 -3033 1187 -3027
rect 1191 -3033 1194 -3027
rect 1198 -3033 1201 -3027
rect 1205 -3033 1208 -3027
rect 1212 -3033 1215 -3027
rect 1219 -3033 1222 -3027
rect 1226 -3033 1229 -3027
rect 1233 -3033 1236 -3027
rect 1240 -3033 1243 -3027
rect 1247 -3033 1250 -3027
rect 1254 -3033 1257 -3027
rect 1261 -3033 1264 -3027
rect 1268 -3033 1271 -3027
rect 1275 -3033 1278 -3027
rect 1282 -3033 1285 -3027
rect 1289 -3033 1292 -3027
rect 1296 -3033 1299 -3027
rect 1303 -3033 1306 -3027
rect 1310 -3033 1313 -3027
rect 1317 -3033 1320 -3027
rect 1324 -3033 1327 -3027
rect 1331 -3033 1334 -3027
rect 1338 -3033 1341 -3027
rect 1345 -3033 1348 -3027
rect 1352 -3033 1355 -3027
rect 1359 -3033 1362 -3027
rect 1366 -3033 1369 -3027
rect 1373 -3033 1376 -3027
rect 1380 -3033 1383 -3027
rect 1387 -3033 1390 -3027
rect 1394 -3033 1397 -3027
rect 1401 -3033 1404 -3027
rect 1408 -3033 1411 -3027
rect 1 -3144 7 -3138
rect 8 -3144 14 -3138
rect 15 -3144 21 -3138
rect 22 -3144 28 -3138
rect 29 -3144 35 -3138
rect 36 -3144 42 -3138
rect 43 -3144 49 -3138
rect 50 -3144 56 -3138
rect 57 -3144 63 -3138
rect 64 -3144 70 -3138
rect 71 -3144 77 -3138
rect 78 -3144 84 -3138
rect 99 -3144 102 -3138
rect 106 -3144 109 -3138
rect 113 -3144 116 -3138
rect 120 -3144 123 -3138
rect 127 -3144 130 -3138
rect 134 -3144 137 -3138
rect 141 -3144 144 -3138
rect 148 -3144 151 -3138
rect 155 -3144 161 -3138
rect 162 -3144 165 -3138
rect 169 -3144 172 -3138
rect 176 -3144 179 -3138
rect 183 -3144 186 -3138
rect 190 -3144 193 -3138
rect 197 -3144 200 -3138
rect 204 -3144 207 -3138
rect 211 -3144 214 -3138
rect 218 -3144 224 -3138
rect 225 -3144 231 -3138
rect 232 -3144 235 -3138
rect 239 -3144 242 -3138
rect 246 -3144 252 -3138
rect 253 -3144 259 -3138
rect 260 -3144 263 -3138
rect 267 -3144 270 -3138
rect 274 -3144 277 -3138
rect 281 -3144 284 -3138
rect 288 -3144 291 -3138
rect 295 -3144 298 -3138
rect 302 -3144 305 -3138
rect 309 -3144 312 -3138
rect 316 -3144 319 -3138
rect 323 -3144 329 -3138
rect 330 -3144 333 -3138
rect 337 -3144 340 -3138
rect 344 -3144 347 -3138
rect 351 -3144 354 -3138
rect 358 -3144 361 -3138
rect 365 -3144 368 -3138
rect 372 -3144 375 -3138
rect 379 -3144 382 -3138
rect 386 -3144 392 -3138
rect 393 -3144 396 -3138
rect 400 -3144 403 -3138
rect 407 -3144 413 -3138
rect 414 -3144 417 -3138
rect 421 -3144 424 -3138
rect 428 -3144 431 -3138
rect 435 -3144 438 -3138
rect 442 -3144 445 -3138
rect 449 -3144 452 -3138
rect 456 -3144 459 -3138
rect 463 -3144 466 -3138
rect 470 -3144 473 -3138
rect 477 -3144 480 -3138
rect 484 -3144 487 -3138
rect 491 -3144 494 -3138
rect 498 -3144 501 -3138
rect 505 -3144 508 -3138
rect 512 -3144 518 -3138
rect 519 -3144 522 -3138
rect 526 -3144 529 -3138
rect 533 -3144 536 -3138
rect 540 -3144 543 -3138
rect 547 -3144 550 -3138
rect 554 -3144 557 -3138
rect 561 -3144 564 -3138
rect 568 -3144 571 -3138
rect 575 -3144 578 -3138
rect 582 -3144 585 -3138
rect 589 -3144 595 -3138
rect 596 -3144 599 -3138
rect 603 -3144 609 -3138
rect 610 -3144 613 -3138
rect 617 -3144 620 -3138
rect 624 -3144 627 -3138
rect 631 -3144 634 -3138
rect 638 -3144 641 -3138
rect 645 -3144 651 -3138
rect 652 -3144 655 -3138
rect 659 -3144 662 -3138
rect 666 -3144 669 -3138
rect 673 -3144 676 -3138
rect 680 -3144 683 -3138
rect 687 -3144 690 -3138
rect 694 -3144 700 -3138
rect 701 -3144 704 -3138
rect 708 -3144 711 -3138
rect 715 -3144 718 -3138
rect 722 -3144 725 -3138
rect 729 -3144 732 -3138
rect 736 -3144 742 -3138
rect 743 -3144 749 -3138
rect 750 -3144 753 -3138
rect 757 -3144 763 -3138
rect 764 -3144 767 -3138
rect 771 -3144 774 -3138
rect 778 -3144 781 -3138
rect 785 -3144 788 -3138
rect 792 -3144 798 -3138
rect 799 -3144 802 -3138
rect 806 -3144 812 -3138
rect 813 -3144 816 -3138
rect 820 -3144 823 -3138
rect 827 -3144 830 -3138
rect 834 -3144 837 -3138
rect 841 -3144 844 -3138
rect 848 -3144 851 -3138
rect 855 -3144 858 -3138
rect 862 -3144 865 -3138
rect 869 -3144 872 -3138
rect 876 -3144 879 -3138
rect 883 -3144 886 -3138
rect 890 -3144 893 -3138
rect 897 -3144 903 -3138
rect 904 -3144 907 -3138
rect 911 -3144 917 -3138
rect 918 -3144 921 -3138
rect 925 -3144 928 -3138
rect 932 -3144 935 -3138
rect 939 -3144 942 -3138
rect 946 -3144 949 -3138
rect 953 -3144 956 -3138
rect 960 -3144 963 -3138
rect 967 -3144 970 -3138
rect 974 -3144 977 -3138
rect 981 -3144 984 -3138
rect 988 -3144 991 -3138
rect 995 -3144 998 -3138
rect 1002 -3144 1005 -3138
rect 1009 -3144 1015 -3138
rect 1016 -3144 1019 -3138
rect 1023 -3144 1026 -3138
rect 1030 -3144 1033 -3138
rect 1037 -3144 1040 -3138
rect 1044 -3144 1047 -3138
rect 1051 -3144 1054 -3138
rect 1058 -3144 1061 -3138
rect 1065 -3144 1068 -3138
rect 1072 -3144 1075 -3138
rect 1079 -3144 1082 -3138
rect 1086 -3144 1089 -3138
rect 1093 -3144 1096 -3138
rect 1100 -3144 1103 -3138
rect 1107 -3144 1110 -3138
rect 1114 -3144 1117 -3138
rect 1121 -3144 1124 -3138
rect 1128 -3144 1131 -3138
rect 1135 -3144 1138 -3138
rect 1142 -3144 1145 -3138
rect 1149 -3144 1152 -3138
rect 1156 -3144 1159 -3138
rect 1163 -3144 1166 -3138
rect 1170 -3144 1173 -3138
rect 1177 -3144 1180 -3138
rect 1184 -3144 1187 -3138
rect 1191 -3144 1194 -3138
rect 1198 -3144 1204 -3138
rect 1205 -3144 1211 -3138
rect 1212 -3144 1215 -3138
rect 1219 -3144 1222 -3138
rect 1226 -3144 1229 -3138
rect 1233 -3144 1236 -3138
rect 1240 -3144 1243 -3138
rect 1247 -3144 1250 -3138
rect 1254 -3144 1257 -3138
rect 1261 -3144 1264 -3138
rect 1268 -3144 1271 -3138
rect 1275 -3144 1278 -3138
rect 1282 -3144 1285 -3138
rect 1289 -3144 1292 -3138
rect 1296 -3144 1299 -3138
rect 1303 -3144 1306 -3138
rect 1310 -3144 1313 -3138
rect 1317 -3144 1320 -3138
rect 1324 -3144 1327 -3138
rect 1331 -3144 1337 -3138
rect 1338 -3144 1341 -3138
rect 1352 -3144 1355 -3138
rect 1359 -3144 1362 -3138
rect 1366 -3144 1369 -3138
rect 1373 -3144 1376 -3138
rect 1 -3237 7 -3231
rect 8 -3237 14 -3231
rect 15 -3237 21 -3231
rect 22 -3237 28 -3231
rect 29 -3237 35 -3231
rect 36 -3237 42 -3231
rect 43 -3237 49 -3231
rect 50 -3237 56 -3231
rect 57 -3237 63 -3231
rect 64 -3237 70 -3231
rect 71 -3237 77 -3231
rect 78 -3237 84 -3231
rect 85 -3237 91 -3231
rect 92 -3237 98 -3231
rect 162 -3237 165 -3231
rect 169 -3237 172 -3231
rect 176 -3237 179 -3231
rect 183 -3237 189 -3231
rect 190 -3237 193 -3231
rect 197 -3237 200 -3231
rect 204 -3237 207 -3231
rect 211 -3237 214 -3231
rect 218 -3237 221 -3231
rect 225 -3237 228 -3231
rect 232 -3237 235 -3231
rect 239 -3237 242 -3231
rect 246 -3237 249 -3231
rect 253 -3237 256 -3231
rect 260 -3237 263 -3231
rect 267 -3237 270 -3231
rect 274 -3237 277 -3231
rect 281 -3237 287 -3231
rect 288 -3237 291 -3231
rect 295 -3237 298 -3231
rect 302 -3237 305 -3231
rect 309 -3237 312 -3231
rect 316 -3237 319 -3231
rect 323 -3237 326 -3231
rect 330 -3237 333 -3231
rect 337 -3237 340 -3231
rect 344 -3237 347 -3231
rect 351 -3237 354 -3231
rect 358 -3237 361 -3231
rect 365 -3237 368 -3231
rect 372 -3237 375 -3231
rect 379 -3237 382 -3231
rect 386 -3237 389 -3231
rect 393 -3237 396 -3231
rect 400 -3237 403 -3231
rect 407 -3237 410 -3231
rect 414 -3237 417 -3231
rect 421 -3237 424 -3231
rect 428 -3237 431 -3231
rect 435 -3237 438 -3231
rect 442 -3237 445 -3231
rect 449 -3237 452 -3231
rect 456 -3237 462 -3231
rect 463 -3237 466 -3231
rect 470 -3237 473 -3231
rect 477 -3237 483 -3231
rect 484 -3237 487 -3231
rect 491 -3237 494 -3231
rect 498 -3237 501 -3231
rect 505 -3237 508 -3231
rect 512 -3237 515 -3231
rect 519 -3237 522 -3231
rect 526 -3237 529 -3231
rect 533 -3237 536 -3231
rect 540 -3237 546 -3231
rect 547 -3237 550 -3231
rect 554 -3237 557 -3231
rect 561 -3237 564 -3231
rect 568 -3237 571 -3231
rect 575 -3237 581 -3231
rect 582 -3237 585 -3231
rect 589 -3237 592 -3231
rect 596 -3237 599 -3231
rect 603 -3237 606 -3231
rect 610 -3237 613 -3231
rect 617 -3237 620 -3231
rect 624 -3237 627 -3231
rect 631 -3237 637 -3231
rect 638 -3237 641 -3231
rect 645 -3237 648 -3231
rect 652 -3237 655 -3231
rect 659 -3237 662 -3231
rect 666 -3237 669 -3231
rect 673 -3237 676 -3231
rect 680 -3237 683 -3231
rect 687 -3237 690 -3231
rect 694 -3237 697 -3231
rect 701 -3237 704 -3231
rect 708 -3237 714 -3231
rect 715 -3237 718 -3231
rect 722 -3237 725 -3231
rect 729 -3237 732 -3231
rect 736 -3237 739 -3231
rect 743 -3237 749 -3231
rect 750 -3237 756 -3231
rect 757 -3237 760 -3231
rect 764 -3237 770 -3231
rect 771 -3237 774 -3231
rect 778 -3237 781 -3231
rect 785 -3237 788 -3231
rect 792 -3237 795 -3231
rect 799 -3237 802 -3231
rect 806 -3237 812 -3231
rect 813 -3237 816 -3231
rect 820 -3237 823 -3231
rect 827 -3237 830 -3231
rect 834 -3237 837 -3231
rect 841 -3237 844 -3231
rect 848 -3237 851 -3231
rect 855 -3237 858 -3231
rect 862 -3237 865 -3231
rect 869 -3237 872 -3231
rect 876 -3237 879 -3231
rect 883 -3237 886 -3231
rect 890 -3237 896 -3231
rect 897 -3237 900 -3231
rect 904 -3237 907 -3231
rect 911 -3237 914 -3231
rect 918 -3237 921 -3231
rect 925 -3237 928 -3231
rect 932 -3237 935 -3231
rect 939 -3237 945 -3231
rect 946 -3237 949 -3231
rect 953 -3237 956 -3231
rect 960 -3237 966 -3231
rect 967 -3237 970 -3231
rect 974 -3237 977 -3231
rect 981 -3237 984 -3231
rect 988 -3237 991 -3231
rect 995 -3237 998 -3231
rect 1002 -3237 1005 -3231
rect 1009 -3237 1012 -3231
rect 1016 -3237 1019 -3231
rect 1023 -3237 1026 -3231
rect 1030 -3237 1033 -3231
rect 1037 -3237 1040 -3231
rect 1044 -3237 1047 -3231
rect 1051 -3237 1054 -3231
rect 1058 -3237 1061 -3231
rect 1065 -3237 1068 -3231
rect 1072 -3237 1075 -3231
rect 1079 -3237 1082 -3231
rect 1086 -3237 1089 -3231
rect 1093 -3237 1096 -3231
rect 1100 -3237 1103 -3231
rect 1107 -3237 1110 -3231
rect 1114 -3237 1117 -3231
rect 1121 -3237 1124 -3231
rect 1128 -3237 1131 -3231
rect 1135 -3237 1138 -3231
rect 1142 -3237 1145 -3231
rect 1149 -3237 1152 -3231
rect 1156 -3237 1159 -3231
rect 1163 -3237 1169 -3231
rect 1170 -3237 1173 -3231
rect 1177 -3237 1180 -3231
rect 1184 -3237 1187 -3231
rect 1191 -3237 1194 -3231
rect 1198 -3237 1204 -3231
rect 1205 -3237 1208 -3231
rect 1212 -3237 1215 -3231
rect 1219 -3237 1222 -3231
rect 1226 -3237 1232 -3231
rect 1233 -3237 1236 -3231
rect 1240 -3237 1243 -3231
rect 1247 -3237 1250 -3231
rect 1254 -3237 1260 -3231
rect 1261 -3237 1264 -3231
rect 1268 -3237 1271 -3231
rect 1275 -3237 1278 -3231
rect 1282 -3237 1288 -3231
rect 1289 -3237 1295 -3231
rect 1296 -3237 1299 -3231
rect 1303 -3237 1306 -3231
rect 1345 -3237 1348 -3231
rect 1352 -3237 1355 -3231
rect 1359 -3237 1362 -3231
rect 1 -3314 7 -3308
rect 8 -3314 14 -3308
rect 15 -3314 21 -3308
rect 22 -3314 28 -3308
rect 29 -3314 35 -3308
rect 36 -3314 42 -3308
rect 43 -3314 49 -3308
rect 50 -3314 56 -3308
rect 57 -3314 63 -3308
rect 64 -3314 70 -3308
rect 71 -3314 77 -3308
rect 78 -3314 84 -3308
rect 85 -3314 91 -3308
rect 92 -3314 98 -3308
rect 155 -3314 158 -3308
rect 162 -3314 165 -3308
rect 169 -3314 172 -3308
rect 176 -3314 179 -3308
rect 183 -3314 186 -3308
rect 190 -3314 193 -3308
rect 197 -3314 203 -3308
rect 204 -3314 207 -3308
rect 211 -3314 214 -3308
rect 218 -3314 221 -3308
rect 225 -3314 228 -3308
rect 232 -3314 235 -3308
rect 239 -3314 245 -3308
rect 246 -3314 249 -3308
rect 253 -3314 256 -3308
rect 260 -3314 263 -3308
rect 267 -3314 270 -3308
rect 274 -3314 277 -3308
rect 281 -3314 284 -3308
rect 288 -3314 291 -3308
rect 295 -3314 298 -3308
rect 302 -3314 305 -3308
rect 309 -3314 312 -3308
rect 316 -3314 319 -3308
rect 323 -3314 326 -3308
rect 330 -3314 333 -3308
rect 337 -3314 340 -3308
rect 344 -3314 347 -3308
rect 351 -3314 354 -3308
rect 358 -3314 361 -3308
rect 365 -3314 368 -3308
rect 372 -3314 375 -3308
rect 379 -3314 382 -3308
rect 386 -3314 389 -3308
rect 393 -3314 399 -3308
rect 400 -3314 403 -3308
rect 407 -3314 410 -3308
rect 414 -3314 417 -3308
rect 421 -3314 424 -3308
rect 428 -3314 431 -3308
rect 435 -3314 438 -3308
rect 442 -3314 445 -3308
rect 449 -3314 452 -3308
rect 456 -3314 459 -3308
rect 463 -3314 466 -3308
rect 470 -3314 473 -3308
rect 477 -3314 480 -3308
rect 484 -3314 490 -3308
rect 491 -3314 494 -3308
rect 498 -3314 501 -3308
rect 505 -3314 508 -3308
rect 512 -3314 515 -3308
rect 519 -3314 522 -3308
rect 526 -3314 529 -3308
rect 533 -3314 539 -3308
rect 540 -3314 543 -3308
rect 547 -3314 550 -3308
rect 554 -3314 557 -3308
rect 561 -3314 564 -3308
rect 568 -3314 571 -3308
rect 575 -3314 578 -3308
rect 582 -3314 585 -3308
rect 589 -3314 592 -3308
rect 596 -3314 599 -3308
rect 603 -3314 606 -3308
rect 610 -3314 616 -3308
rect 617 -3314 620 -3308
rect 624 -3314 627 -3308
rect 631 -3314 634 -3308
rect 638 -3314 641 -3308
rect 645 -3314 648 -3308
rect 652 -3314 658 -3308
rect 659 -3314 665 -3308
rect 666 -3314 672 -3308
rect 673 -3314 676 -3308
rect 680 -3314 683 -3308
rect 687 -3314 693 -3308
rect 694 -3314 697 -3308
rect 701 -3314 704 -3308
rect 708 -3314 711 -3308
rect 715 -3314 718 -3308
rect 722 -3314 725 -3308
rect 729 -3314 735 -3308
rect 736 -3314 739 -3308
rect 743 -3314 746 -3308
rect 750 -3314 753 -3308
rect 757 -3314 763 -3308
rect 764 -3314 767 -3308
rect 771 -3314 774 -3308
rect 778 -3314 781 -3308
rect 785 -3314 788 -3308
rect 792 -3314 795 -3308
rect 799 -3314 802 -3308
rect 806 -3314 809 -3308
rect 813 -3314 816 -3308
rect 820 -3314 826 -3308
rect 827 -3314 830 -3308
rect 834 -3314 840 -3308
rect 841 -3314 844 -3308
rect 848 -3314 851 -3308
rect 855 -3314 861 -3308
rect 862 -3314 865 -3308
rect 869 -3314 875 -3308
rect 876 -3314 879 -3308
rect 883 -3314 886 -3308
rect 890 -3314 896 -3308
rect 897 -3314 900 -3308
rect 904 -3314 907 -3308
rect 911 -3314 914 -3308
rect 918 -3314 921 -3308
rect 925 -3314 928 -3308
rect 932 -3314 935 -3308
rect 939 -3314 942 -3308
rect 946 -3314 949 -3308
rect 953 -3314 956 -3308
rect 960 -3314 963 -3308
rect 967 -3314 970 -3308
rect 974 -3314 977 -3308
rect 981 -3314 984 -3308
rect 988 -3314 991 -3308
rect 995 -3314 998 -3308
rect 1002 -3314 1008 -3308
rect 1009 -3314 1012 -3308
rect 1016 -3314 1019 -3308
rect 1023 -3314 1029 -3308
rect 1030 -3314 1033 -3308
rect 1037 -3314 1040 -3308
rect 1044 -3314 1047 -3308
rect 1051 -3314 1054 -3308
rect 1058 -3314 1061 -3308
rect 1065 -3314 1068 -3308
rect 1072 -3314 1075 -3308
rect 1079 -3314 1082 -3308
rect 1086 -3314 1089 -3308
rect 1093 -3314 1096 -3308
rect 1100 -3314 1103 -3308
rect 1107 -3314 1110 -3308
rect 1114 -3314 1117 -3308
rect 1121 -3314 1124 -3308
rect 1128 -3314 1131 -3308
rect 1135 -3314 1141 -3308
rect 1142 -3314 1145 -3308
rect 1149 -3314 1152 -3308
rect 1156 -3314 1159 -3308
rect 1163 -3314 1166 -3308
rect 1170 -3314 1173 -3308
rect 1177 -3314 1180 -3308
rect 1184 -3314 1187 -3308
rect 1191 -3314 1194 -3308
rect 1198 -3314 1201 -3308
rect 1205 -3314 1208 -3308
rect 1212 -3314 1215 -3308
rect 1219 -3314 1222 -3308
rect 1226 -3314 1229 -3308
rect 1233 -3314 1236 -3308
rect 1240 -3314 1243 -3308
rect 1247 -3314 1250 -3308
rect 1254 -3314 1257 -3308
rect 1261 -3314 1264 -3308
rect 1268 -3314 1274 -3308
rect 1275 -3314 1278 -3308
rect 1289 -3314 1292 -3308
rect 1338 -3314 1341 -3308
rect 1345 -3314 1348 -3308
rect 1352 -3314 1355 -3308
rect 1 -3387 7 -3381
rect 8 -3387 14 -3381
rect 15 -3387 21 -3381
rect 22 -3387 28 -3381
rect 29 -3387 35 -3381
rect 36 -3387 42 -3381
rect 43 -3387 49 -3381
rect 50 -3387 56 -3381
rect 57 -3387 63 -3381
rect 64 -3387 70 -3381
rect 71 -3387 77 -3381
rect 78 -3387 84 -3381
rect 85 -3387 91 -3381
rect 92 -3387 98 -3381
rect 197 -3387 200 -3381
rect 204 -3387 207 -3381
rect 211 -3387 214 -3381
rect 218 -3387 221 -3381
rect 225 -3387 228 -3381
rect 232 -3387 235 -3381
rect 239 -3387 242 -3381
rect 246 -3387 249 -3381
rect 253 -3387 256 -3381
rect 260 -3387 266 -3381
rect 267 -3387 273 -3381
rect 274 -3387 280 -3381
rect 281 -3387 284 -3381
rect 288 -3387 291 -3381
rect 295 -3387 298 -3381
rect 302 -3387 305 -3381
rect 309 -3387 312 -3381
rect 316 -3387 319 -3381
rect 323 -3387 326 -3381
rect 330 -3387 333 -3381
rect 337 -3387 340 -3381
rect 344 -3387 347 -3381
rect 351 -3387 354 -3381
rect 358 -3387 361 -3381
rect 365 -3387 368 -3381
rect 372 -3387 375 -3381
rect 379 -3387 382 -3381
rect 386 -3387 389 -3381
rect 393 -3387 396 -3381
rect 400 -3387 406 -3381
rect 407 -3387 413 -3381
rect 414 -3387 417 -3381
rect 421 -3387 427 -3381
rect 428 -3387 431 -3381
rect 435 -3387 438 -3381
rect 442 -3387 445 -3381
rect 449 -3387 452 -3381
rect 456 -3387 459 -3381
rect 463 -3387 466 -3381
rect 470 -3387 476 -3381
rect 477 -3387 480 -3381
rect 484 -3387 487 -3381
rect 491 -3387 494 -3381
rect 498 -3387 501 -3381
rect 505 -3387 508 -3381
rect 512 -3387 515 -3381
rect 519 -3387 522 -3381
rect 526 -3387 529 -3381
rect 533 -3387 536 -3381
rect 540 -3387 546 -3381
rect 547 -3387 550 -3381
rect 554 -3387 560 -3381
rect 561 -3387 564 -3381
rect 568 -3387 574 -3381
rect 575 -3387 581 -3381
rect 582 -3387 585 -3381
rect 589 -3387 592 -3381
rect 596 -3387 599 -3381
rect 603 -3387 606 -3381
rect 610 -3387 613 -3381
rect 617 -3387 620 -3381
rect 624 -3387 627 -3381
rect 631 -3387 634 -3381
rect 638 -3387 641 -3381
rect 645 -3387 648 -3381
rect 652 -3387 658 -3381
rect 659 -3387 662 -3381
rect 666 -3387 669 -3381
rect 673 -3387 676 -3381
rect 680 -3387 683 -3381
rect 687 -3387 690 -3381
rect 694 -3387 697 -3381
rect 701 -3387 704 -3381
rect 708 -3387 711 -3381
rect 715 -3387 718 -3381
rect 722 -3387 725 -3381
rect 729 -3387 732 -3381
rect 736 -3387 739 -3381
rect 743 -3387 746 -3381
rect 750 -3387 753 -3381
rect 757 -3387 763 -3381
rect 764 -3387 767 -3381
rect 771 -3387 774 -3381
rect 778 -3387 781 -3381
rect 785 -3387 788 -3381
rect 792 -3387 798 -3381
rect 799 -3387 802 -3381
rect 806 -3387 809 -3381
rect 813 -3387 816 -3381
rect 820 -3387 823 -3381
rect 827 -3387 830 -3381
rect 834 -3387 837 -3381
rect 841 -3387 844 -3381
rect 848 -3387 851 -3381
rect 855 -3387 858 -3381
rect 862 -3387 865 -3381
rect 869 -3387 872 -3381
rect 876 -3387 879 -3381
rect 883 -3387 886 -3381
rect 890 -3387 893 -3381
rect 897 -3387 900 -3381
rect 904 -3387 907 -3381
rect 911 -3387 914 -3381
rect 918 -3387 921 -3381
rect 925 -3387 928 -3381
rect 932 -3387 935 -3381
rect 939 -3387 942 -3381
rect 946 -3387 949 -3381
rect 953 -3387 959 -3381
rect 960 -3387 963 -3381
rect 967 -3387 970 -3381
rect 974 -3387 977 -3381
rect 981 -3387 984 -3381
rect 988 -3387 991 -3381
rect 995 -3387 998 -3381
rect 1002 -3387 1005 -3381
rect 1009 -3387 1015 -3381
rect 1016 -3387 1019 -3381
rect 1023 -3387 1026 -3381
rect 1030 -3387 1033 -3381
rect 1037 -3387 1043 -3381
rect 1044 -3387 1047 -3381
rect 1051 -3387 1057 -3381
rect 1058 -3387 1061 -3381
rect 1065 -3387 1071 -3381
rect 1072 -3387 1075 -3381
rect 1079 -3387 1082 -3381
rect 1086 -3387 1089 -3381
rect 1093 -3387 1096 -3381
rect 1100 -3387 1103 -3381
rect 1121 -3387 1124 -3381
rect 1128 -3387 1131 -3381
rect 1177 -3387 1183 -3381
rect 1184 -3387 1187 -3381
rect 1191 -3387 1194 -3381
rect 1338 -3387 1341 -3381
rect 1345 -3387 1348 -3381
rect 1352 -3387 1355 -3381
rect 1 -3450 7 -3444
rect 8 -3450 14 -3444
rect 15 -3450 21 -3444
rect 22 -3450 28 -3444
rect 29 -3450 35 -3444
rect 36 -3450 42 -3444
rect 43 -3450 49 -3444
rect 50 -3450 56 -3444
rect 57 -3450 63 -3444
rect 64 -3450 70 -3444
rect 71 -3450 77 -3444
rect 78 -3450 84 -3444
rect 85 -3450 91 -3444
rect 92 -3450 98 -3444
rect 99 -3450 105 -3444
rect 106 -3450 112 -3444
rect 246 -3450 249 -3444
rect 260 -3450 263 -3444
rect 288 -3450 294 -3444
rect 309 -3450 312 -3444
rect 316 -3450 319 -3444
rect 323 -3450 326 -3444
rect 330 -3450 333 -3444
rect 337 -3450 340 -3444
rect 344 -3450 350 -3444
rect 351 -3450 354 -3444
rect 358 -3450 361 -3444
rect 365 -3450 371 -3444
rect 372 -3450 375 -3444
rect 379 -3450 382 -3444
rect 386 -3450 389 -3444
rect 393 -3450 396 -3444
rect 400 -3450 403 -3444
rect 407 -3450 410 -3444
rect 414 -3450 417 -3444
rect 421 -3450 424 -3444
rect 428 -3450 431 -3444
rect 435 -3450 438 -3444
rect 442 -3450 448 -3444
rect 449 -3450 452 -3444
rect 456 -3450 459 -3444
rect 463 -3450 466 -3444
rect 470 -3450 473 -3444
rect 477 -3450 480 -3444
rect 484 -3450 487 -3444
rect 491 -3450 494 -3444
rect 498 -3450 504 -3444
rect 505 -3450 508 -3444
rect 512 -3450 515 -3444
rect 519 -3450 522 -3444
rect 526 -3450 532 -3444
rect 533 -3450 536 -3444
rect 540 -3450 543 -3444
rect 547 -3450 553 -3444
rect 554 -3450 557 -3444
rect 561 -3450 564 -3444
rect 568 -3450 571 -3444
rect 575 -3450 578 -3444
rect 582 -3450 588 -3444
rect 589 -3450 592 -3444
rect 596 -3450 599 -3444
rect 603 -3450 606 -3444
rect 610 -3450 613 -3444
rect 617 -3450 620 -3444
rect 624 -3450 627 -3444
rect 631 -3450 634 -3444
rect 638 -3450 641 -3444
rect 645 -3450 651 -3444
rect 652 -3450 655 -3444
rect 659 -3450 662 -3444
rect 666 -3450 669 -3444
rect 673 -3450 676 -3444
rect 680 -3450 683 -3444
rect 687 -3450 693 -3444
rect 694 -3450 697 -3444
rect 701 -3450 704 -3444
rect 708 -3450 711 -3444
rect 715 -3450 718 -3444
rect 722 -3450 725 -3444
rect 729 -3450 732 -3444
rect 736 -3450 742 -3444
rect 743 -3450 746 -3444
rect 750 -3450 753 -3444
rect 757 -3450 760 -3444
rect 764 -3450 767 -3444
rect 771 -3450 774 -3444
rect 778 -3450 781 -3444
rect 785 -3450 788 -3444
rect 792 -3450 795 -3444
rect 799 -3450 802 -3444
rect 806 -3450 809 -3444
rect 813 -3450 816 -3444
rect 820 -3450 826 -3444
rect 827 -3450 830 -3444
rect 834 -3450 837 -3444
rect 841 -3450 844 -3444
rect 848 -3450 851 -3444
rect 855 -3450 861 -3444
rect 862 -3450 865 -3444
rect 869 -3450 875 -3444
rect 876 -3450 879 -3444
rect 883 -3450 889 -3444
rect 890 -3450 893 -3444
rect 897 -3450 903 -3444
rect 904 -3450 907 -3444
rect 911 -3450 914 -3444
rect 918 -3450 921 -3444
rect 925 -3450 928 -3444
rect 932 -3450 935 -3444
rect 939 -3450 942 -3444
rect 946 -3450 949 -3444
rect 953 -3450 956 -3444
rect 960 -3450 963 -3444
rect 967 -3450 970 -3444
rect 974 -3450 977 -3444
rect 981 -3450 984 -3444
rect 1002 -3450 1005 -3444
rect 1009 -3450 1012 -3444
rect 1023 -3450 1029 -3444
rect 1030 -3450 1033 -3444
rect 1037 -3450 1040 -3444
rect 1044 -3450 1047 -3444
rect 1086 -3450 1089 -3444
rect 1093 -3450 1096 -3444
rect 1114 -3450 1117 -3444
rect 1135 -3450 1138 -3444
rect 1177 -3450 1180 -3444
rect 1338 -3450 1341 -3444
rect 1345 -3450 1348 -3444
rect 1352 -3450 1355 -3444
rect 1 -3507 7 -3501
rect 8 -3507 14 -3501
rect 15 -3507 21 -3501
rect 22 -3507 28 -3501
rect 29 -3507 35 -3501
rect 36 -3507 42 -3501
rect 43 -3507 49 -3501
rect 50 -3507 56 -3501
rect 57 -3507 63 -3501
rect 64 -3507 70 -3501
rect 71 -3507 77 -3501
rect 78 -3507 84 -3501
rect 85 -3507 91 -3501
rect 92 -3507 98 -3501
rect 99 -3507 105 -3501
rect 106 -3507 112 -3501
rect 113 -3507 119 -3501
rect 246 -3507 249 -3501
rect 260 -3507 263 -3501
rect 274 -3507 277 -3501
rect 330 -3507 333 -3501
rect 337 -3507 340 -3501
rect 344 -3507 347 -3501
rect 351 -3507 354 -3501
rect 358 -3507 361 -3501
rect 365 -3507 368 -3501
rect 372 -3507 375 -3501
rect 379 -3507 382 -3501
rect 386 -3507 389 -3501
rect 393 -3507 396 -3501
rect 400 -3507 403 -3501
rect 407 -3507 410 -3501
rect 414 -3507 417 -3501
rect 421 -3507 427 -3501
rect 428 -3507 431 -3501
rect 435 -3507 438 -3501
rect 442 -3507 445 -3501
rect 449 -3507 452 -3501
rect 456 -3507 459 -3501
rect 463 -3507 469 -3501
rect 470 -3507 473 -3501
rect 477 -3507 480 -3501
rect 484 -3507 487 -3501
rect 491 -3507 497 -3501
rect 498 -3507 501 -3501
rect 505 -3507 508 -3501
rect 512 -3507 515 -3501
rect 519 -3507 522 -3501
rect 526 -3507 529 -3501
rect 533 -3507 539 -3501
rect 540 -3507 543 -3501
rect 547 -3507 550 -3501
rect 554 -3507 557 -3501
rect 561 -3507 567 -3501
rect 568 -3507 571 -3501
rect 575 -3507 581 -3501
rect 582 -3507 585 -3501
rect 589 -3507 592 -3501
rect 596 -3507 599 -3501
rect 603 -3507 606 -3501
rect 610 -3507 613 -3501
rect 617 -3507 620 -3501
rect 624 -3507 630 -3501
rect 631 -3507 634 -3501
rect 638 -3507 644 -3501
rect 645 -3507 648 -3501
rect 652 -3507 655 -3501
rect 659 -3507 662 -3501
rect 666 -3507 669 -3501
rect 673 -3507 679 -3501
rect 680 -3507 683 -3501
rect 687 -3507 690 -3501
rect 694 -3507 697 -3501
rect 701 -3507 704 -3501
rect 708 -3507 711 -3501
rect 715 -3507 718 -3501
rect 722 -3507 728 -3501
rect 729 -3507 732 -3501
rect 736 -3507 739 -3501
rect 743 -3507 746 -3501
rect 750 -3507 753 -3501
rect 757 -3507 760 -3501
rect 764 -3507 767 -3501
rect 771 -3507 774 -3501
rect 778 -3507 781 -3501
rect 799 -3507 802 -3501
rect 806 -3507 809 -3501
rect 813 -3507 819 -3501
rect 820 -3507 823 -3501
rect 834 -3507 837 -3501
rect 841 -3507 844 -3501
rect 848 -3507 851 -3501
rect 855 -3507 858 -3501
rect 862 -3507 865 -3501
rect 869 -3507 872 -3501
rect 876 -3507 879 -3501
rect 904 -3507 907 -3501
rect 911 -3507 914 -3501
rect 918 -3507 921 -3501
rect 925 -3507 928 -3501
rect 932 -3507 935 -3501
rect 939 -3507 942 -3501
rect 946 -3507 949 -3501
rect 953 -3507 959 -3501
rect 960 -3507 963 -3501
rect 967 -3507 970 -3501
rect 981 -3507 984 -3501
rect 988 -3507 991 -3501
rect 995 -3507 1001 -3501
rect 1002 -3507 1005 -3501
rect 1009 -3507 1012 -3501
rect 1051 -3507 1054 -3501
rect 1079 -3507 1082 -3501
rect 1086 -3507 1089 -3501
rect 1107 -3507 1110 -3501
rect 1121 -3507 1124 -3501
rect 1149 -3507 1152 -3501
rect 1170 -3507 1176 -3501
rect 1177 -3507 1180 -3501
rect 1338 -3507 1341 -3501
rect 1345 -3507 1351 -3501
rect 1352 -3507 1355 -3501
rect 1 -3548 7 -3542
rect 8 -3548 14 -3542
rect 15 -3548 21 -3542
rect 22 -3548 28 -3542
rect 29 -3548 35 -3542
rect 36 -3548 42 -3542
rect 43 -3548 49 -3542
rect 50 -3548 56 -3542
rect 57 -3548 63 -3542
rect 64 -3548 70 -3542
rect 71 -3548 77 -3542
rect 78 -3548 84 -3542
rect 85 -3548 91 -3542
rect 92 -3548 98 -3542
rect 99 -3548 105 -3542
rect 106 -3548 112 -3542
rect 113 -3548 119 -3542
rect 120 -3548 126 -3542
rect 246 -3548 249 -3542
rect 253 -3548 259 -3542
rect 260 -3548 263 -3542
rect 267 -3548 270 -3542
rect 295 -3548 298 -3542
rect 344 -3548 347 -3542
rect 358 -3548 361 -3542
rect 379 -3548 382 -3542
rect 393 -3548 396 -3542
rect 400 -3548 403 -3542
rect 407 -3548 410 -3542
rect 414 -3548 417 -3542
rect 421 -3548 424 -3542
rect 428 -3548 434 -3542
rect 435 -3548 438 -3542
rect 442 -3548 448 -3542
rect 449 -3548 455 -3542
rect 456 -3548 459 -3542
rect 463 -3548 466 -3542
rect 470 -3548 473 -3542
rect 477 -3548 480 -3542
rect 484 -3548 490 -3542
rect 491 -3548 494 -3542
rect 498 -3548 501 -3542
rect 505 -3548 508 -3542
rect 512 -3548 515 -3542
rect 519 -3548 522 -3542
rect 526 -3548 529 -3542
rect 533 -3548 536 -3542
rect 540 -3548 546 -3542
rect 547 -3548 550 -3542
rect 554 -3548 557 -3542
rect 561 -3548 564 -3542
rect 568 -3548 571 -3542
rect 575 -3548 578 -3542
rect 582 -3548 585 -3542
rect 589 -3548 592 -3542
rect 596 -3548 602 -3542
rect 603 -3548 606 -3542
rect 610 -3548 613 -3542
rect 624 -3548 630 -3542
rect 638 -3548 641 -3542
rect 666 -3548 669 -3542
rect 680 -3548 683 -3542
rect 687 -3548 693 -3542
rect 694 -3548 697 -3542
rect 701 -3548 704 -3542
rect 708 -3548 711 -3542
rect 715 -3548 718 -3542
rect 722 -3548 725 -3542
rect 729 -3548 732 -3542
rect 736 -3548 739 -3542
rect 743 -3548 746 -3542
rect 750 -3548 753 -3542
rect 757 -3548 760 -3542
rect 764 -3548 767 -3542
rect 834 -3548 837 -3542
rect 848 -3548 851 -3542
rect 862 -3548 865 -3542
rect 869 -3548 872 -3542
rect 876 -3548 879 -3542
rect 883 -3548 886 -3542
rect 890 -3548 893 -3542
rect 897 -3548 900 -3542
rect 904 -3548 907 -3542
rect 911 -3548 914 -3542
rect 918 -3548 924 -3542
rect 925 -3548 928 -3542
rect 932 -3548 938 -3542
rect 939 -3548 945 -3542
rect 946 -3548 949 -3542
rect 967 -3548 970 -3542
rect 974 -3548 977 -3542
rect 988 -3548 991 -3542
rect 1002 -3548 1008 -3542
rect 1009 -3548 1012 -3542
rect 1051 -3548 1054 -3542
rect 1058 -3548 1061 -3542
rect 1079 -3548 1082 -3542
rect 1107 -3548 1110 -3542
rect 1149 -3548 1152 -3542
rect 1156 -3548 1162 -3542
rect 1 -3585 7 -3579
rect 8 -3585 14 -3579
rect 15 -3585 21 -3579
rect 22 -3585 28 -3579
rect 29 -3585 35 -3579
rect 36 -3585 42 -3579
rect 43 -3585 49 -3579
rect 50 -3585 56 -3579
rect 57 -3585 63 -3579
rect 64 -3585 70 -3579
rect 71 -3585 77 -3579
rect 78 -3585 84 -3579
rect 85 -3585 91 -3579
rect 92 -3585 98 -3579
rect 99 -3585 105 -3579
rect 106 -3585 112 -3579
rect 113 -3585 119 -3579
rect 120 -3585 126 -3579
rect 260 -3585 266 -3579
rect 267 -3585 270 -3579
rect 309 -3585 312 -3579
rect 323 -3585 329 -3579
rect 351 -3585 354 -3579
rect 358 -3585 361 -3579
rect 365 -3585 368 -3579
rect 372 -3585 378 -3579
rect 393 -3585 396 -3579
rect 400 -3585 406 -3579
rect 407 -3585 410 -3579
rect 414 -3585 417 -3579
rect 435 -3585 438 -3579
rect 442 -3585 448 -3579
rect 449 -3585 455 -3579
rect 456 -3585 459 -3579
rect 463 -3585 466 -3579
rect 470 -3585 473 -3579
rect 477 -3585 480 -3579
rect 484 -3585 490 -3579
rect 491 -3585 494 -3579
rect 498 -3585 501 -3579
rect 505 -3585 508 -3579
rect 512 -3585 518 -3579
rect 519 -3585 522 -3579
rect 526 -3585 529 -3579
rect 533 -3585 536 -3579
rect 540 -3585 543 -3579
rect 547 -3585 550 -3579
rect 554 -3585 557 -3579
rect 561 -3585 564 -3579
rect 568 -3585 571 -3579
rect 596 -3585 599 -3579
rect 610 -3585 613 -3579
rect 617 -3585 620 -3579
rect 645 -3585 648 -3579
rect 659 -3585 662 -3579
rect 673 -3585 679 -3579
rect 687 -3585 690 -3579
rect 694 -3585 697 -3579
rect 701 -3585 704 -3579
rect 708 -3585 711 -3579
rect 715 -3585 718 -3579
rect 722 -3585 725 -3579
rect 729 -3585 732 -3579
rect 736 -3585 739 -3579
rect 743 -3585 746 -3579
rect 750 -3585 753 -3579
rect 757 -3585 760 -3579
rect 764 -3585 767 -3579
rect 848 -3585 851 -3579
rect 855 -3585 858 -3579
rect 890 -3585 893 -3579
rect 897 -3585 903 -3579
rect 904 -3585 907 -3579
rect 911 -3585 914 -3579
rect 918 -3585 924 -3579
rect 925 -3585 928 -3579
rect 939 -3585 942 -3579
rect 967 -3585 970 -3579
rect 974 -3585 977 -3579
rect 981 -3585 987 -3579
rect 988 -3585 991 -3579
rect 1037 -3585 1040 -3579
rect 1051 -3585 1054 -3579
rect 1079 -3585 1085 -3579
rect 1086 -3585 1089 -3579
rect 1107 -3585 1110 -3579
rect 1 -3608 7 -3602
rect 8 -3608 14 -3602
rect 15 -3608 21 -3602
rect 22 -3608 28 -3602
rect 29 -3608 35 -3602
rect 36 -3608 42 -3602
rect 43 -3608 49 -3602
rect 50 -3608 56 -3602
rect 57 -3608 63 -3602
rect 64 -3608 70 -3602
rect 71 -3608 77 -3602
rect 78 -3608 84 -3602
rect 85 -3608 91 -3602
rect 92 -3608 98 -3602
rect 99 -3608 105 -3602
rect 106 -3608 112 -3602
rect 113 -3608 119 -3602
rect 120 -3608 126 -3602
rect 127 -3608 133 -3602
rect 134 -3608 140 -3602
rect 141 -3608 147 -3602
rect 148 -3608 154 -3602
rect 155 -3608 161 -3602
rect 162 -3608 168 -3602
rect 169 -3608 175 -3602
rect 176 -3608 182 -3602
rect 183 -3608 189 -3602
rect 190 -3608 196 -3602
rect 197 -3608 203 -3602
rect 204 -3608 210 -3602
rect 211 -3608 217 -3602
rect 218 -3608 224 -3602
rect 225 -3608 231 -3602
rect 232 -3608 238 -3602
rect 323 -3608 329 -3602
rect 351 -3608 357 -3602
rect 400 -3608 403 -3602
rect 407 -3608 410 -3602
rect 456 -3608 459 -3602
rect 470 -3608 473 -3602
rect 491 -3608 494 -3602
rect 505 -3608 508 -3602
rect 512 -3608 518 -3602
rect 519 -3608 522 -3602
rect 540 -3608 546 -3602
rect 547 -3608 550 -3602
rect 554 -3608 557 -3602
rect 561 -3608 564 -3602
rect 568 -3608 571 -3602
rect 575 -3608 578 -3602
rect 596 -3608 599 -3602
rect 603 -3608 606 -3602
rect 610 -3608 616 -3602
rect 680 -3608 686 -3602
rect 694 -3608 697 -3602
rect 701 -3608 704 -3602
rect 708 -3608 711 -3602
rect 715 -3608 718 -3602
rect 722 -3608 725 -3602
rect 729 -3608 732 -3602
rect 736 -3608 739 -3602
rect 743 -3608 746 -3602
rect 750 -3608 753 -3602
rect 757 -3608 763 -3602
rect 764 -3608 767 -3602
rect 771 -3608 774 -3602
rect 855 -3608 858 -3602
rect 862 -3608 865 -3602
rect 904 -3608 910 -3602
rect 918 -3608 921 -3602
rect 925 -3608 928 -3602
rect 974 -3608 977 -3602
rect 981 -3608 984 -3602
rect 1030 -3608 1033 -3602
rect 1044 -3608 1047 -3602
rect 1051 -3608 1054 -3602
rect 1107 -3608 1110 -3602
rect 1 -3633 7 -3627
rect 8 -3633 14 -3627
rect 15 -3633 21 -3627
rect 22 -3633 28 -3627
rect 29 -3633 35 -3627
rect 36 -3633 42 -3627
rect 43 -3633 49 -3627
rect 50 -3633 56 -3627
rect 57 -3633 63 -3627
rect 64 -3633 70 -3627
rect 71 -3633 77 -3627
rect 78 -3633 84 -3627
rect 85 -3633 91 -3627
rect 92 -3633 98 -3627
rect 99 -3633 105 -3627
rect 106 -3633 112 -3627
rect 113 -3633 119 -3627
rect 120 -3633 126 -3627
rect 127 -3633 133 -3627
rect 134 -3633 140 -3627
rect 141 -3633 147 -3627
rect 148 -3633 154 -3627
rect 155 -3633 161 -3627
rect 162 -3633 168 -3627
rect 169 -3633 175 -3627
rect 176 -3633 182 -3627
rect 183 -3633 189 -3627
rect 190 -3633 196 -3627
rect 400 -3633 403 -3627
rect 407 -3633 410 -3627
rect 463 -3633 466 -3627
rect 470 -3633 473 -3627
rect 526 -3633 529 -3627
rect 561 -3633 564 -3627
rect 568 -3633 571 -3627
rect 575 -3633 578 -3627
rect 582 -3633 585 -3627
rect 589 -3633 592 -3627
rect 701 -3633 704 -3627
rect 708 -3633 711 -3627
rect 715 -3633 718 -3627
rect 722 -3633 725 -3627
rect 743 -3633 746 -3627
rect 750 -3633 753 -3627
rect 757 -3633 760 -3627
rect 764 -3633 767 -3627
rect 771 -3633 777 -3627
rect 799 -3633 802 -3627
rect 855 -3633 858 -3627
rect 862 -3633 865 -3627
rect 925 -3633 928 -3627
rect 932 -3633 935 -3627
rect 981 -3633 984 -3627
rect 1002 -3633 1005 -3627
rect 1030 -3633 1033 -3627
rect 1051 -3633 1057 -3627
rect 1058 -3633 1061 -3627
rect 1079 -3633 1082 -3627
rect 1107 -3633 1110 -3627
rect 1 -3648 7 -3642
rect 8 -3648 14 -3642
rect 15 -3648 21 -3642
rect 22 -3648 28 -3642
rect 29 -3648 35 -3642
rect 36 -3648 42 -3642
rect 43 -3648 49 -3642
rect 50 -3648 56 -3642
rect 57 -3648 63 -3642
rect 64 -3648 70 -3642
rect 71 -3648 77 -3642
rect 78 -3648 84 -3642
rect 85 -3648 91 -3642
rect 92 -3648 98 -3642
rect 99 -3648 105 -3642
rect 400 -3648 403 -3642
rect 407 -3648 410 -3642
rect 463 -3648 466 -3642
rect 470 -3648 476 -3642
rect 526 -3648 529 -3642
rect 568 -3648 574 -3642
rect 575 -3648 578 -3642
rect 582 -3648 588 -3642
rect 589 -3648 592 -3642
rect 596 -3648 599 -3642
rect 708 -3648 711 -3642
rect 715 -3648 721 -3642
rect 722 -3648 725 -3642
rect 750 -3648 753 -3642
rect 757 -3648 760 -3642
rect 764 -3648 767 -3642
rect 855 -3648 861 -3642
rect 862 -3648 865 -3642
rect 925 -3648 931 -3642
rect 932 -3648 935 -3642
rect 981 -3648 987 -3642
rect 988 -3648 991 -3642
rect 1030 -3648 1036 -3642
rect 1093 -3648 1096 -3642
rect 1107 -3648 1113 -3642
rect 1 -3663 7 -3657
rect 8 -3663 14 -3657
rect 15 -3663 21 -3657
rect 22 -3663 28 -3657
rect 29 -3663 35 -3657
rect 36 -3663 42 -3657
rect 43 -3663 49 -3657
rect 50 -3663 56 -3657
rect 57 -3663 63 -3657
rect 64 -3663 70 -3657
rect 71 -3663 77 -3657
rect 78 -3663 84 -3657
rect 85 -3663 91 -3657
rect 92 -3663 98 -3657
rect 99 -3663 105 -3657
rect 400 -3663 406 -3657
rect 407 -3663 410 -3657
rect 526 -3663 532 -3657
rect 533 -3663 536 -3657
rect 757 -3663 760 -3657
rect 764 -3663 770 -3657
rect 771 -3663 774 -3657
rect 1 -3674 7 -3668
rect 8 -3674 14 -3668
rect 15 -3674 21 -3668
rect 22 -3674 28 -3668
rect 29 -3674 35 -3668
rect 36 -3674 42 -3668
rect 43 -3674 49 -3668
rect 50 -3674 56 -3668
rect 57 -3674 63 -3668
rect 64 -3674 70 -3668
rect 71 -3674 77 -3668
rect 78 -3674 84 -3668
rect 85 -3674 91 -3668
rect 1 -3683 7 -3677
rect 8 -3683 14 -3677
rect 15 -3683 21 -3677
rect 22 -3683 28 -3677
rect 29 -3683 35 -3677
rect 36 -3683 42 -3677
rect 43 -3683 49 -3677
rect 50 -3683 56 -3677
rect 57 -3683 63 -3677
rect 64 -3683 70 -3677
rect 71 -3683 77 -3677
rect 78 -3683 84 -3677
rect 85 -3683 91 -3677
rect 1 -3692 7 -3686
rect 8 -3692 14 -3686
rect 15 -3692 21 -3686
rect 22 -3692 28 -3686
rect 29 -3692 35 -3686
rect 36 -3692 42 -3686
rect 43 -3692 49 -3686
rect 50 -3692 56 -3686
rect 57 -3692 63 -3686
rect 64 -3692 70 -3686
rect 71 -3692 77 -3686
rect 78 -3692 84 -3686
rect 85 -3692 91 -3686
rect 1 -3701 7 -3695
rect 8 -3701 14 -3695
rect 15 -3701 21 -3695
rect 22 -3701 28 -3695
rect 29 -3701 35 -3695
rect 36 -3701 42 -3695
rect 43 -3701 49 -3695
rect 50 -3701 56 -3695
rect 57 -3701 63 -3695
rect 64 -3701 70 -3695
<< polysilicon >>
rect 226 -9 227 -7
rect 226 -15 227 -13
rect 254 -9 255 -7
rect 254 -15 255 -13
rect 275 -9 276 -7
rect 275 -15 276 -13
rect 317 -9 318 -7
rect 317 -15 318 -13
rect 331 -9 332 -7
rect 331 -15 332 -13
rect 366 -9 367 -7
rect 366 -15 367 -13
rect 373 -9 374 -7
rect 376 -15 377 -13
rect 380 -9 381 -7
rect 383 -15 384 -13
rect 394 -15 395 -13
rect 401 -9 402 -7
rect 404 -9 405 -7
rect 415 -9 416 -7
rect 415 -15 416 -13
rect 429 -9 430 -7
rect 436 -9 437 -7
rect 436 -15 437 -13
rect 443 -15 444 -13
rect 446 -15 447 -13
rect 450 -9 451 -7
rect 450 -15 451 -13
rect 457 -9 458 -7
rect 460 -9 461 -7
rect 457 -15 458 -13
rect 471 -9 472 -7
rect 471 -15 472 -13
rect 492 -9 493 -7
rect 492 -15 493 -13
rect 506 -9 507 -7
rect 506 -15 507 -13
rect 513 -9 514 -7
rect 516 -9 517 -7
rect 527 -9 528 -7
rect 527 -15 528 -13
rect 534 -9 535 -7
rect 537 -9 538 -7
rect 541 -15 542 -13
rect 562 -9 563 -7
rect 565 -15 566 -13
rect 569 -9 570 -7
rect 569 -15 570 -13
rect 590 -9 591 -7
rect 590 -15 591 -13
rect 618 -15 619 -13
rect 642 -9 643 -7
rect 639 -15 640 -13
rect 667 -9 668 -7
rect 674 -9 675 -7
rect 674 -15 675 -13
rect 705 -9 706 -7
rect 705 -15 706 -13
rect 765 -9 766 -7
rect 765 -15 766 -13
rect 800 -9 801 -7
rect 803 -9 804 -7
rect 828 -9 829 -7
rect 828 -15 829 -13
rect 842 -9 843 -7
rect 842 -15 843 -13
rect 135 -38 136 -36
rect 135 -44 136 -42
rect 177 -44 178 -42
rect 180 -44 181 -42
rect 191 -38 192 -36
rect 191 -44 192 -42
rect 205 -38 206 -36
rect 205 -44 206 -42
rect 212 -38 213 -36
rect 212 -44 213 -42
rect 222 -38 223 -36
rect 222 -44 223 -42
rect 226 -38 227 -36
rect 226 -44 227 -42
rect 236 -44 237 -42
rect 254 -38 255 -36
rect 254 -44 255 -42
rect 296 -38 297 -36
rect 299 -38 300 -36
rect 296 -44 297 -42
rect 303 -38 304 -36
rect 303 -44 304 -42
rect 310 -38 311 -36
rect 310 -44 311 -42
rect 317 -38 318 -36
rect 317 -44 318 -42
rect 327 -38 328 -36
rect 327 -44 328 -42
rect 331 -38 332 -36
rect 331 -44 332 -42
rect 338 -38 339 -36
rect 338 -44 339 -42
rect 345 -38 346 -36
rect 345 -44 346 -42
rect 352 -38 353 -36
rect 352 -44 353 -42
rect 359 -38 360 -36
rect 359 -44 360 -42
rect 366 -38 367 -36
rect 366 -44 367 -42
rect 369 -44 370 -42
rect 373 -38 374 -36
rect 373 -44 374 -42
rect 380 -38 381 -36
rect 380 -44 381 -42
rect 387 -38 388 -36
rect 387 -44 388 -42
rect 394 -38 395 -36
rect 397 -44 398 -42
rect 401 -38 402 -36
rect 404 -38 405 -36
rect 408 -38 409 -36
rect 408 -44 409 -42
rect 415 -38 416 -36
rect 415 -44 416 -42
rect 422 -38 423 -36
rect 422 -44 423 -42
rect 443 -38 444 -36
rect 446 -38 447 -36
rect 450 -38 451 -36
rect 450 -44 451 -42
rect 453 -44 454 -42
rect 457 -38 458 -36
rect 457 -44 458 -42
rect 464 -38 465 -36
rect 464 -44 465 -42
rect 467 -44 468 -42
rect 471 -38 472 -36
rect 471 -44 472 -42
rect 478 -38 479 -36
rect 478 -44 479 -42
rect 488 -38 489 -36
rect 488 -44 489 -42
rect 492 -38 493 -36
rect 492 -44 493 -42
rect 513 -38 514 -36
rect 513 -44 514 -42
rect 520 -38 521 -36
rect 520 -44 521 -42
rect 527 -38 528 -36
rect 527 -44 528 -42
rect 534 -38 535 -36
rect 534 -44 535 -42
rect 541 -38 542 -36
rect 541 -44 542 -42
rect 548 -38 549 -36
rect 548 -44 549 -42
rect 555 -38 556 -36
rect 555 -44 556 -42
rect 569 -38 570 -36
rect 569 -44 570 -42
rect 576 -38 577 -36
rect 576 -44 577 -42
rect 583 -38 584 -36
rect 583 -44 584 -42
rect 590 -44 591 -42
rect 593 -44 594 -42
rect 618 -38 619 -36
rect 618 -44 619 -42
rect 621 -44 622 -42
rect 632 -38 633 -36
rect 635 -38 636 -36
rect 639 -38 640 -36
rect 639 -44 640 -42
rect 646 -38 647 -36
rect 646 -44 647 -42
rect 653 -38 654 -36
rect 653 -44 654 -42
rect 660 -38 661 -36
rect 660 -44 661 -42
rect 667 -38 668 -36
rect 667 -44 668 -42
rect 684 -38 685 -36
rect 681 -44 682 -42
rect 695 -38 696 -36
rect 695 -44 696 -42
rect 702 -38 703 -36
rect 702 -44 703 -42
rect 709 -38 710 -36
rect 709 -44 710 -42
rect 761 -38 762 -36
rect 761 -44 762 -42
rect 765 -38 766 -36
rect 765 -44 766 -42
rect 775 -38 776 -36
rect 782 -38 783 -36
rect 786 -38 787 -36
rect 786 -44 787 -42
rect 793 -38 794 -36
rect 793 -44 794 -42
rect 800 -38 801 -36
rect 800 -44 801 -42
rect 821 -38 822 -36
rect 824 -44 825 -42
rect 856 -38 857 -36
rect 856 -44 857 -42
rect 877 -38 878 -36
rect 877 -44 878 -42
rect 919 -38 920 -36
rect 919 -44 920 -42
rect 79 -87 80 -85
rect 79 -93 80 -91
rect 100 -87 101 -85
rect 100 -93 101 -91
rect 114 -93 115 -91
rect 117 -93 118 -91
rect 128 -87 129 -85
rect 128 -93 129 -91
rect 142 -87 143 -85
rect 142 -93 143 -91
rect 145 -93 146 -91
rect 149 -87 150 -85
rect 149 -93 150 -91
rect 156 -87 157 -85
rect 156 -93 157 -91
rect 163 -87 164 -85
rect 163 -93 164 -91
rect 170 -87 171 -85
rect 170 -93 171 -91
rect 177 -87 178 -85
rect 180 -87 181 -85
rect 177 -93 178 -91
rect 184 -87 185 -85
rect 184 -93 185 -91
rect 191 -87 192 -85
rect 191 -93 192 -91
rect 198 -87 199 -85
rect 198 -93 199 -91
rect 205 -87 206 -85
rect 205 -93 206 -91
rect 212 -93 213 -91
rect 215 -93 216 -91
rect 219 -87 220 -85
rect 219 -93 220 -91
rect 226 -87 227 -85
rect 229 -87 230 -85
rect 226 -93 227 -91
rect 236 -87 237 -85
rect 236 -93 237 -91
rect 243 -87 244 -85
rect 240 -93 241 -91
rect 254 -87 255 -85
rect 254 -93 255 -91
rect 261 -87 262 -85
rect 261 -93 262 -91
rect 268 -87 269 -85
rect 268 -93 269 -91
rect 278 -87 279 -85
rect 275 -93 276 -91
rect 278 -93 279 -91
rect 282 -93 283 -91
rect 285 -93 286 -91
rect 289 -87 290 -85
rect 289 -93 290 -91
rect 296 -87 297 -85
rect 296 -93 297 -91
rect 299 -93 300 -91
rect 303 -87 304 -85
rect 303 -93 304 -91
rect 310 -87 311 -85
rect 310 -93 311 -91
rect 317 -87 318 -85
rect 317 -93 318 -91
rect 324 -87 325 -85
rect 324 -93 325 -91
rect 331 -87 332 -85
rect 334 -93 335 -91
rect 338 -87 339 -85
rect 338 -93 339 -91
rect 345 -87 346 -85
rect 345 -93 346 -91
rect 352 -87 353 -85
rect 352 -93 353 -91
rect 359 -87 360 -85
rect 359 -93 360 -91
rect 366 -87 367 -85
rect 369 -87 370 -85
rect 366 -93 367 -91
rect 373 -87 374 -85
rect 373 -93 374 -91
rect 380 -87 381 -85
rect 401 -87 402 -85
rect 401 -93 402 -91
rect 408 -87 409 -85
rect 408 -93 409 -91
rect 415 -87 416 -85
rect 415 -93 416 -91
rect 422 -87 423 -85
rect 422 -93 423 -91
rect 429 -87 430 -85
rect 429 -93 430 -91
rect 436 -87 437 -85
rect 436 -93 437 -91
rect 446 -87 447 -85
rect 443 -93 444 -91
rect 446 -93 447 -91
rect 450 -87 451 -85
rect 450 -93 451 -91
rect 453 -93 454 -91
rect 457 -87 458 -85
rect 457 -93 458 -91
rect 464 -87 465 -85
rect 464 -93 465 -91
rect 474 -87 475 -85
rect 471 -93 472 -91
rect 478 -87 479 -85
rect 478 -93 479 -91
rect 485 -87 486 -85
rect 485 -93 486 -91
rect 492 -87 493 -85
rect 492 -93 493 -91
rect 499 -87 500 -85
rect 499 -93 500 -91
rect 506 -87 507 -85
rect 506 -93 507 -91
rect 513 -87 514 -85
rect 513 -93 514 -91
rect 520 -87 521 -85
rect 520 -93 521 -91
rect 527 -87 528 -85
rect 527 -93 528 -91
rect 534 -87 535 -85
rect 534 -93 535 -91
rect 541 -87 542 -85
rect 541 -93 542 -91
rect 548 -87 549 -85
rect 548 -93 549 -91
rect 555 -87 556 -85
rect 555 -93 556 -91
rect 562 -87 563 -85
rect 562 -93 563 -91
rect 569 -87 570 -85
rect 572 -87 573 -85
rect 569 -93 570 -91
rect 576 -87 577 -85
rect 576 -93 577 -91
rect 583 -87 584 -85
rect 583 -93 584 -91
rect 593 -87 594 -85
rect 590 -93 591 -91
rect 597 -87 598 -85
rect 597 -93 598 -91
rect 604 -87 605 -85
rect 604 -93 605 -91
rect 611 -87 612 -85
rect 611 -93 612 -91
rect 618 -87 619 -85
rect 618 -93 619 -91
rect 625 -87 626 -85
rect 628 -87 629 -85
rect 632 -87 633 -85
rect 632 -93 633 -91
rect 642 -87 643 -85
rect 642 -93 643 -91
rect 646 -87 647 -85
rect 646 -93 647 -91
rect 649 -93 650 -91
rect 653 -87 654 -85
rect 653 -93 654 -91
rect 660 -87 661 -85
rect 660 -93 661 -91
rect 667 -87 668 -85
rect 667 -93 668 -91
rect 674 -87 675 -85
rect 674 -93 675 -91
rect 681 -87 682 -85
rect 681 -93 682 -91
rect 688 -87 689 -85
rect 688 -93 689 -91
rect 695 -87 696 -85
rect 695 -93 696 -91
rect 702 -87 703 -85
rect 702 -93 703 -91
rect 709 -87 710 -85
rect 709 -93 710 -91
rect 716 -87 717 -85
rect 716 -93 717 -91
rect 723 -87 724 -85
rect 723 -93 724 -91
rect 733 -87 734 -85
rect 730 -93 731 -91
rect 740 -87 741 -85
rect 740 -93 741 -91
rect 744 -87 745 -85
rect 744 -93 745 -91
rect 751 -87 752 -85
rect 751 -93 752 -91
rect 758 -87 759 -85
rect 761 -93 762 -91
rect 765 -87 766 -85
rect 765 -93 766 -91
rect 772 -87 773 -85
rect 772 -93 773 -91
rect 779 -87 780 -85
rect 782 -87 783 -85
rect 786 -87 787 -85
rect 786 -93 787 -91
rect 793 -87 794 -85
rect 793 -93 794 -91
rect 800 -87 801 -85
rect 800 -93 801 -91
rect 807 -87 808 -85
rect 807 -93 808 -91
rect 814 -87 815 -85
rect 814 -93 815 -91
rect 821 -87 822 -85
rect 821 -93 822 -91
rect 856 -87 857 -85
rect 856 -93 857 -91
rect 863 -87 864 -85
rect 863 -93 864 -91
rect 870 -87 871 -85
rect 870 -93 871 -91
rect 891 -87 892 -85
rect 891 -93 892 -91
rect 905 -87 906 -85
rect 905 -93 906 -91
rect 968 -87 969 -85
rect 968 -93 969 -91
rect 100 -158 101 -156
rect 100 -164 101 -162
rect 114 -158 115 -156
rect 114 -164 115 -162
rect 149 -158 150 -156
rect 149 -164 150 -162
rect 156 -164 157 -162
rect 163 -158 164 -156
rect 163 -164 164 -162
rect 170 -158 171 -156
rect 170 -164 171 -162
rect 177 -158 178 -156
rect 177 -164 178 -162
rect 184 -158 185 -156
rect 184 -164 185 -162
rect 191 -158 192 -156
rect 191 -164 192 -162
rect 198 -158 199 -156
rect 198 -164 199 -162
rect 205 -158 206 -156
rect 205 -164 206 -162
rect 212 -158 213 -156
rect 212 -164 213 -162
rect 219 -158 220 -156
rect 219 -164 220 -162
rect 226 -158 227 -156
rect 226 -164 227 -162
rect 233 -158 234 -156
rect 233 -164 234 -162
rect 240 -158 241 -156
rect 240 -164 241 -162
rect 250 -158 251 -156
rect 247 -164 248 -162
rect 250 -164 251 -162
rect 254 -158 255 -156
rect 257 -164 258 -162
rect 261 -158 262 -156
rect 261 -164 262 -162
rect 268 -158 269 -156
rect 271 -158 272 -156
rect 271 -164 272 -162
rect 275 -158 276 -156
rect 275 -164 276 -162
rect 278 -164 279 -162
rect 282 -158 283 -156
rect 285 -158 286 -156
rect 282 -164 283 -162
rect 289 -158 290 -156
rect 292 -158 293 -156
rect 289 -164 290 -162
rect 292 -164 293 -162
rect 296 -158 297 -156
rect 299 -158 300 -156
rect 296 -164 297 -162
rect 303 -158 304 -156
rect 303 -164 304 -162
rect 310 -158 311 -156
rect 310 -164 311 -162
rect 317 -158 318 -156
rect 317 -164 318 -162
rect 324 -158 325 -156
rect 324 -164 325 -162
rect 331 -158 332 -156
rect 331 -164 332 -162
rect 338 -158 339 -156
rect 338 -164 339 -162
rect 345 -158 346 -156
rect 345 -164 346 -162
rect 352 -158 353 -156
rect 352 -164 353 -162
rect 359 -158 360 -156
rect 359 -164 360 -162
rect 366 -158 367 -156
rect 366 -164 367 -162
rect 373 -158 374 -156
rect 373 -164 374 -162
rect 380 -164 381 -162
rect 390 -158 391 -156
rect 387 -164 388 -162
rect 390 -164 391 -162
rect 394 -158 395 -156
rect 394 -164 395 -162
rect 401 -158 402 -156
rect 401 -164 402 -162
rect 408 -158 409 -156
rect 408 -164 409 -162
rect 415 -158 416 -156
rect 418 -158 419 -156
rect 418 -164 419 -162
rect 422 -158 423 -156
rect 422 -164 423 -162
rect 429 -158 430 -156
rect 432 -158 433 -156
rect 429 -164 430 -162
rect 432 -164 433 -162
rect 436 -158 437 -156
rect 436 -164 437 -162
rect 443 -158 444 -156
rect 443 -164 444 -162
rect 450 -158 451 -156
rect 450 -164 451 -162
rect 457 -158 458 -156
rect 457 -164 458 -162
rect 464 -158 465 -156
rect 467 -158 468 -156
rect 464 -164 465 -162
rect 467 -164 468 -162
rect 471 -158 472 -156
rect 474 -158 475 -156
rect 474 -164 475 -162
rect 478 -158 479 -156
rect 478 -164 479 -162
rect 488 -158 489 -156
rect 485 -164 486 -162
rect 488 -164 489 -162
rect 492 -158 493 -156
rect 492 -164 493 -162
rect 499 -158 500 -156
rect 499 -164 500 -162
rect 506 -158 507 -156
rect 509 -158 510 -156
rect 506 -164 507 -162
rect 509 -164 510 -162
rect 513 -158 514 -156
rect 513 -164 514 -162
rect 520 -158 521 -156
rect 520 -164 521 -162
rect 527 -158 528 -156
rect 527 -164 528 -162
rect 534 -158 535 -156
rect 534 -164 535 -162
rect 541 -158 542 -156
rect 541 -164 542 -162
rect 548 -158 549 -156
rect 548 -164 549 -162
rect 558 -158 559 -156
rect 558 -164 559 -162
rect 562 -158 563 -156
rect 562 -164 563 -162
rect 569 -158 570 -156
rect 569 -164 570 -162
rect 576 -158 577 -156
rect 576 -164 577 -162
rect 583 -158 584 -156
rect 583 -164 584 -162
rect 590 -158 591 -156
rect 590 -164 591 -162
rect 597 -158 598 -156
rect 597 -164 598 -162
rect 604 -158 605 -156
rect 604 -164 605 -162
rect 611 -158 612 -156
rect 611 -164 612 -162
rect 618 -158 619 -156
rect 618 -164 619 -162
rect 621 -164 622 -162
rect 625 -158 626 -156
rect 625 -164 626 -162
rect 632 -158 633 -156
rect 632 -164 633 -162
rect 639 -158 640 -156
rect 639 -164 640 -162
rect 646 -158 647 -156
rect 649 -158 650 -156
rect 646 -164 647 -162
rect 653 -158 654 -156
rect 653 -164 654 -162
rect 660 -158 661 -156
rect 660 -164 661 -162
rect 667 -158 668 -156
rect 667 -164 668 -162
rect 674 -158 675 -156
rect 674 -164 675 -162
rect 681 -158 682 -156
rect 684 -158 685 -156
rect 681 -164 682 -162
rect 688 -158 689 -156
rect 695 -164 696 -162
rect 698 -164 699 -162
rect 702 -158 703 -156
rect 702 -164 703 -162
rect 705 -164 706 -162
rect 709 -158 710 -156
rect 709 -164 710 -162
rect 712 -164 713 -162
rect 716 -158 717 -156
rect 716 -164 717 -162
rect 723 -158 724 -156
rect 723 -164 724 -162
rect 730 -158 731 -156
rect 730 -164 731 -162
rect 737 -158 738 -156
rect 737 -164 738 -162
rect 744 -158 745 -156
rect 744 -164 745 -162
rect 751 -158 752 -156
rect 754 -158 755 -156
rect 754 -164 755 -162
rect 758 -158 759 -156
rect 758 -164 759 -162
rect 765 -158 766 -156
rect 765 -164 766 -162
rect 772 -158 773 -156
rect 772 -164 773 -162
rect 779 -158 780 -156
rect 779 -164 780 -162
rect 786 -158 787 -156
rect 786 -164 787 -162
rect 793 -158 794 -156
rect 793 -164 794 -162
rect 800 -158 801 -156
rect 800 -164 801 -162
rect 807 -158 808 -156
rect 807 -164 808 -162
rect 814 -158 815 -156
rect 814 -164 815 -162
rect 821 -158 822 -156
rect 821 -164 822 -162
rect 828 -158 829 -156
rect 828 -164 829 -162
rect 835 -158 836 -156
rect 835 -164 836 -162
rect 842 -158 843 -156
rect 842 -164 843 -162
rect 849 -158 850 -156
rect 849 -164 850 -162
rect 856 -158 857 -156
rect 856 -164 857 -162
rect 863 -158 864 -156
rect 863 -164 864 -162
rect 870 -158 871 -156
rect 870 -164 871 -162
rect 877 -158 878 -156
rect 877 -164 878 -162
rect 884 -158 885 -156
rect 884 -164 885 -162
rect 891 -158 892 -156
rect 891 -164 892 -162
rect 898 -158 899 -156
rect 898 -164 899 -162
rect 905 -158 906 -156
rect 905 -164 906 -162
rect 912 -158 913 -156
rect 912 -164 913 -162
rect 919 -158 920 -156
rect 919 -164 920 -162
rect 926 -158 927 -156
rect 926 -164 927 -162
rect 933 -158 934 -156
rect 933 -164 934 -162
rect 940 -158 941 -156
rect 943 -164 944 -162
rect 947 -158 948 -156
rect 947 -164 948 -162
rect 954 -158 955 -156
rect 954 -164 955 -162
rect 961 -158 962 -156
rect 961 -164 962 -162
rect 968 -158 969 -156
rect 968 -164 969 -162
rect 975 -158 976 -156
rect 975 -164 976 -162
rect 982 -158 983 -156
rect 982 -164 983 -162
rect 989 -158 990 -156
rect 989 -164 990 -162
rect 996 -164 997 -162
rect 999 -164 1000 -162
rect 1003 -158 1004 -156
rect 1003 -164 1004 -162
rect 54 -259 55 -257
rect 72 -253 73 -251
rect 72 -259 73 -257
rect 100 -253 101 -251
rect 100 -259 101 -257
rect 107 -253 108 -251
rect 110 -253 111 -251
rect 107 -259 108 -257
rect 110 -259 111 -257
rect 114 -253 115 -251
rect 114 -259 115 -257
rect 121 -253 122 -251
rect 124 -253 125 -251
rect 124 -259 125 -257
rect 128 -253 129 -251
rect 128 -259 129 -257
rect 135 -253 136 -251
rect 135 -259 136 -257
rect 163 -253 164 -251
rect 166 -253 167 -251
rect 163 -259 164 -257
rect 173 -253 174 -251
rect 170 -259 171 -257
rect 173 -259 174 -257
rect 177 -253 178 -251
rect 177 -259 178 -257
rect 184 -253 185 -251
rect 184 -259 185 -257
rect 191 -253 192 -251
rect 191 -259 192 -257
rect 198 -253 199 -251
rect 198 -259 199 -257
rect 205 -253 206 -251
rect 208 -253 209 -251
rect 205 -259 206 -257
rect 208 -259 209 -257
rect 212 -253 213 -251
rect 212 -259 213 -257
rect 219 -253 220 -251
rect 222 -253 223 -251
rect 219 -259 220 -257
rect 226 -253 227 -251
rect 226 -259 227 -257
rect 233 -253 234 -251
rect 233 -259 234 -257
rect 247 -253 248 -251
rect 247 -259 248 -257
rect 254 -253 255 -251
rect 254 -259 255 -257
rect 261 -253 262 -251
rect 261 -259 262 -257
rect 268 -253 269 -251
rect 268 -259 269 -257
rect 275 -253 276 -251
rect 275 -259 276 -257
rect 282 -253 283 -251
rect 285 -253 286 -251
rect 282 -259 283 -257
rect 289 -253 290 -251
rect 289 -259 290 -257
rect 296 -253 297 -251
rect 296 -259 297 -257
rect 303 -253 304 -251
rect 303 -259 304 -257
rect 310 -253 311 -251
rect 310 -259 311 -257
rect 317 -259 318 -257
rect 320 -259 321 -257
rect 324 -253 325 -251
rect 324 -259 325 -257
rect 331 -253 332 -251
rect 331 -259 332 -257
rect 338 -253 339 -251
rect 341 -253 342 -251
rect 338 -259 339 -257
rect 341 -259 342 -257
rect 345 -253 346 -251
rect 345 -259 346 -257
rect 352 -253 353 -251
rect 352 -259 353 -257
rect 359 -253 360 -251
rect 359 -259 360 -257
rect 366 -253 367 -251
rect 366 -259 367 -257
rect 373 -253 374 -251
rect 373 -259 374 -257
rect 380 -253 381 -251
rect 380 -259 381 -257
rect 387 -253 388 -251
rect 387 -259 388 -257
rect 394 -253 395 -251
rect 394 -259 395 -257
rect 401 -253 402 -251
rect 404 -253 405 -251
rect 401 -259 402 -257
rect 404 -259 405 -257
rect 408 -253 409 -251
rect 408 -259 409 -257
rect 415 -253 416 -251
rect 415 -259 416 -257
rect 422 -253 423 -251
rect 422 -259 423 -257
rect 429 -253 430 -251
rect 432 -253 433 -251
rect 436 -253 437 -251
rect 436 -259 437 -257
rect 443 -253 444 -251
rect 446 -253 447 -251
rect 446 -259 447 -257
rect 450 -253 451 -251
rect 453 -253 454 -251
rect 450 -259 451 -257
rect 457 -253 458 -251
rect 457 -259 458 -257
rect 464 -253 465 -251
rect 464 -259 465 -257
rect 471 -253 472 -251
rect 471 -259 472 -257
rect 478 -253 479 -251
rect 481 -253 482 -251
rect 478 -259 479 -257
rect 481 -259 482 -257
rect 488 -253 489 -251
rect 485 -259 486 -257
rect 488 -259 489 -257
rect 492 -253 493 -251
rect 495 -253 496 -251
rect 492 -259 493 -257
rect 495 -259 496 -257
rect 499 -253 500 -251
rect 499 -259 500 -257
rect 506 -253 507 -251
rect 506 -259 507 -257
rect 513 -253 514 -251
rect 513 -259 514 -257
rect 516 -259 517 -257
rect 520 -253 521 -251
rect 520 -259 521 -257
rect 527 -253 528 -251
rect 527 -259 528 -257
rect 534 -253 535 -251
rect 534 -259 535 -257
rect 541 -253 542 -251
rect 541 -259 542 -257
rect 544 -259 545 -257
rect 548 -253 549 -251
rect 548 -259 549 -257
rect 555 -253 556 -251
rect 555 -259 556 -257
rect 562 -253 563 -251
rect 562 -259 563 -257
rect 569 -253 570 -251
rect 569 -259 570 -257
rect 576 -253 577 -251
rect 576 -259 577 -257
rect 583 -253 584 -251
rect 583 -259 584 -257
rect 586 -259 587 -257
rect 590 -253 591 -251
rect 590 -259 591 -257
rect 597 -253 598 -251
rect 597 -259 598 -257
rect 604 -253 605 -251
rect 604 -259 605 -257
rect 611 -253 612 -251
rect 611 -259 612 -257
rect 614 -259 615 -257
rect 618 -253 619 -251
rect 618 -259 619 -257
rect 625 -253 626 -251
rect 625 -259 626 -257
rect 632 -253 633 -251
rect 632 -259 633 -257
rect 639 -253 640 -251
rect 639 -259 640 -257
rect 646 -253 647 -251
rect 646 -259 647 -257
rect 653 -253 654 -251
rect 653 -259 654 -257
rect 660 -253 661 -251
rect 660 -259 661 -257
rect 667 -253 668 -251
rect 667 -259 668 -257
rect 674 -253 675 -251
rect 674 -259 675 -257
rect 681 -253 682 -251
rect 684 -253 685 -251
rect 688 -259 689 -257
rect 695 -253 696 -251
rect 695 -259 696 -257
rect 702 -253 703 -251
rect 702 -259 703 -257
rect 709 -253 710 -251
rect 712 -253 713 -251
rect 709 -259 710 -257
rect 716 -253 717 -251
rect 716 -259 717 -257
rect 723 -253 724 -251
rect 723 -259 724 -257
rect 730 -253 731 -251
rect 730 -259 731 -257
rect 737 -253 738 -251
rect 737 -259 738 -257
rect 744 -253 745 -251
rect 744 -259 745 -257
rect 751 -253 752 -251
rect 751 -259 752 -257
rect 758 -253 759 -251
rect 758 -259 759 -257
rect 765 -253 766 -251
rect 765 -259 766 -257
rect 768 -259 769 -257
rect 772 -253 773 -251
rect 772 -259 773 -257
rect 779 -253 780 -251
rect 779 -259 780 -257
rect 786 -253 787 -251
rect 786 -259 787 -257
rect 793 -253 794 -251
rect 793 -259 794 -257
rect 800 -253 801 -251
rect 800 -259 801 -257
rect 807 -253 808 -251
rect 807 -259 808 -257
rect 814 -253 815 -251
rect 814 -259 815 -257
rect 821 -253 822 -251
rect 821 -259 822 -257
rect 828 -253 829 -251
rect 831 -259 832 -257
rect 835 -253 836 -251
rect 835 -259 836 -257
rect 842 -259 843 -257
rect 845 -259 846 -257
rect 849 -253 850 -251
rect 849 -259 850 -257
rect 856 -253 857 -251
rect 856 -259 857 -257
rect 863 -253 864 -251
rect 863 -259 864 -257
rect 870 -253 871 -251
rect 870 -259 871 -257
rect 877 -253 878 -251
rect 877 -259 878 -257
rect 884 -253 885 -251
rect 884 -259 885 -257
rect 891 -253 892 -251
rect 891 -259 892 -257
rect 898 -253 899 -251
rect 898 -259 899 -257
rect 905 -253 906 -251
rect 905 -259 906 -257
rect 912 -253 913 -251
rect 912 -259 913 -257
rect 919 -253 920 -251
rect 919 -259 920 -257
rect 926 -253 927 -251
rect 926 -259 927 -257
rect 933 -253 934 -251
rect 933 -259 934 -257
rect 940 -253 941 -251
rect 940 -259 941 -257
rect 947 -253 948 -251
rect 947 -259 948 -257
rect 954 -253 955 -251
rect 954 -259 955 -257
rect 961 -253 962 -251
rect 961 -259 962 -257
rect 968 -253 969 -251
rect 968 -259 969 -257
rect 975 -253 976 -251
rect 975 -259 976 -257
rect 982 -253 983 -251
rect 982 -259 983 -257
rect 989 -253 990 -251
rect 989 -259 990 -257
rect 996 -253 997 -251
rect 996 -259 997 -257
rect 1003 -253 1004 -251
rect 1003 -259 1004 -257
rect 1010 -253 1011 -251
rect 1010 -259 1011 -257
rect 1017 -253 1018 -251
rect 1017 -259 1018 -257
rect 1024 -253 1025 -251
rect 1024 -259 1025 -257
rect 1031 -253 1032 -251
rect 1031 -259 1032 -257
rect 1038 -253 1039 -251
rect 1038 -259 1039 -257
rect 1045 -253 1046 -251
rect 1045 -259 1046 -257
rect 1052 -253 1053 -251
rect 1052 -259 1053 -257
rect 1059 -253 1060 -251
rect 1059 -259 1060 -257
rect 1066 -253 1067 -251
rect 1066 -259 1067 -257
rect 1073 -253 1074 -251
rect 1073 -259 1074 -257
rect 1080 -253 1081 -251
rect 1080 -259 1081 -257
rect 1087 -253 1088 -251
rect 1087 -259 1088 -257
rect 1094 -253 1095 -251
rect 1094 -259 1095 -257
rect 1101 -253 1102 -251
rect 1101 -259 1102 -257
rect 1108 -253 1109 -251
rect 1108 -259 1109 -257
rect 1115 -253 1116 -251
rect 1115 -259 1116 -257
rect 1122 -253 1123 -251
rect 1122 -259 1123 -257
rect 1129 -253 1130 -251
rect 1129 -259 1130 -257
rect 51 -356 52 -354
rect 51 -362 52 -360
rect 58 -356 59 -354
rect 58 -362 59 -360
rect 72 -356 73 -354
rect 72 -362 73 -360
rect 79 -356 80 -354
rect 82 -356 83 -354
rect 82 -362 83 -360
rect 86 -356 87 -354
rect 86 -362 87 -360
rect 93 -356 94 -354
rect 93 -362 94 -360
rect 100 -356 101 -354
rect 100 -362 101 -360
rect 107 -356 108 -354
rect 107 -362 108 -360
rect 114 -356 115 -354
rect 114 -362 115 -360
rect 121 -356 122 -354
rect 124 -356 125 -354
rect 124 -362 125 -360
rect 128 -356 129 -354
rect 128 -362 129 -360
rect 135 -356 136 -354
rect 135 -362 136 -360
rect 142 -356 143 -354
rect 142 -362 143 -360
rect 149 -356 150 -354
rect 149 -362 150 -360
rect 156 -356 157 -354
rect 156 -362 157 -360
rect 159 -362 160 -360
rect 163 -356 164 -354
rect 163 -362 164 -360
rect 170 -356 171 -354
rect 170 -362 171 -360
rect 173 -362 174 -360
rect 177 -356 178 -354
rect 177 -362 178 -360
rect 184 -356 185 -354
rect 184 -362 185 -360
rect 191 -356 192 -354
rect 191 -362 192 -360
rect 198 -356 199 -354
rect 198 -362 199 -360
rect 205 -356 206 -354
rect 205 -362 206 -360
rect 212 -356 213 -354
rect 212 -362 213 -360
rect 219 -356 220 -354
rect 219 -362 220 -360
rect 226 -356 227 -354
rect 226 -362 227 -360
rect 236 -356 237 -354
rect 233 -362 234 -360
rect 240 -356 241 -354
rect 240 -362 241 -360
rect 254 -356 255 -354
rect 254 -362 255 -360
rect 268 -356 269 -354
rect 268 -362 269 -360
rect 275 -356 276 -354
rect 275 -362 276 -360
rect 289 -356 290 -354
rect 289 -362 290 -360
rect 296 -356 297 -354
rect 296 -362 297 -360
rect 303 -356 304 -354
rect 303 -362 304 -360
rect 310 -356 311 -354
rect 310 -362 311 -360
rect 317 -356 318 -354
rect 317 -362 318 -360
rect 324 -356 325 -354
rect 324 -362 325 -360
rect 338 -356 339 -354
rect 338 -362 339 -360
rect 345 -356 346 -354
rect 345 -362 346 -360
rect 352 -356 353 -354
rect 352 -362 353 -360
rect 373 -356 374 -354
rect 373 -362 374 -360
rect 380 -356 381 -354
rect 380 -362 381 -360
rect 387 -356 388 -354
rect 387 -362 388 -360
rect 394 -356 395 -354
rect 394 -362 395 -360
rect 401 -356 402 -354
rect 401 -362 402 -360
rect 408 -356 409 -354
rect 408 -362 409 -360
rect 415 -356 416 -354
rect 415 -362 416 -360
rect 422 -356 423 -354
rect 422 -362 423 -360
rect 429 -356 430 -354
rect 429 -362 430 -360
rect 436 -356 437 -354
rect 436 -362 437 -360
rect 443 -356 444 -354
rect 443 -362 444 -360
rect 450 -356 451 -354
rect 450 -362 451 -360
rect 457 -356 458 -354
rect 457 -362 458 -360
rect 467 -356 468 -354
rect 467 -362 468 -360
rect 471 -356 472 -354
rect 471 -362 472 -360
rect 474 -362 475 -360
rect 478 -356 479 -354
rect 481 -356 482 -354
rect 478 -362 479 -360
rect 481 -362 482 -360
rect 485 -356 486 -354
rect 488 -356 489 -354
rect 485 -362 486 -360
rect 488 -362 489 -360
rect 499 -356 500 -354
rect 499 -362 500 -360
rect 506 -356 507 -354
rect 506 -362 507 -360
rect 513 -356 514 -354
rect 513 -362 514 -360
rect 516 -362 517 -360
rect 520 -356 521 -354
rect 520 -362 521 -360
rect 527 -356 528 -354
rect 530 -356 531 -354
rect 527 -362 528 -360
rect 530 -362 531 -360
rect 534 -356 535 -354
rect 534 -362 535 -360
rect 541 -356 542 -354
rect 541 -362 542 -360
rect 548 -356 549 -354
rect 548 -362 549 -360
rect 555 -356 556 -354
rect 555 -362 556 -360
rect 562 -356 563 -354
rect 562 -362 563 -360
rect 565 -362 566 -360
rect 569 -356 570 -354
rect 569 -362 570 -360
rect 572 -362 573 -360
rect 576 -356 577 -354
rect 579 -356 580 -354
rect 576 -362 577 -360
rect 579 -362 580 -360
rect 583 -356 584 -354
rect 586 -356 587 -354
rect 583 -362 584 -360
rect 586 -362 587 -360
rect 590 -356 591 -354
rect 593 -356 594 -354
rect 590 -362 591 -360
rect 597 -356 598 -354
rect 597 -362 598 -360
rect 604 -356 605 -354
rect 607 -356 608 -354
rect 604 -362 605 -360
rect 607 -362 608 -360
rect 611 -356 612 -354
rect 611 -362 612 -360
rect 618 -356 619 -354
rect 618 -362 619 -360
rect 625 -356 626 -354
rect 625 -362 626 -360
rect 632 -356 633 -354
rect 635 -356 636 -354
rect 632 -362 633 -360
rect 635 -362 636 -360
rect 639 -356 640 -354
rect 639 -362 640 -360
rect 646 -356 647 -354
rect 646 -362 647 -360
rect 653 -356 654 -354
rect 653 -362 654 -360
rect 663 -356 664 -354
rect 660 -362 661 -360
rect 663 -362 664 -360
rect 667 -356 668 -354
rect 667 -362 668 -360
rect 674 -356 675 -354
rect 674 -362 675 -360
rect 684 -356 685 -354
rect 681 -362 682 -360
rect 684 -362 685 -360
rect 688 -356 689 -354
rect 688 -362 689 -360
rect 695 -356 696 -354
rect 695 -362 696 -360
rect 702 -356 703 -354
rect 702 -362 703 -360
rect 709 -356 710 -354
rect 709 -362 710 -360
rect 719 -356 720 -354
rect 716 -362 717 -360
rect 726 -356 727 -354
rect 723 -362 724 -360
rect 726 -362 727 -360
rect 730 -356 731 -354
rect 730 -362 731 -360
rect 737 -356 738 -354
rect 737 -362 738 -360
rect 744 -356 745 -354
rect 744 -362 745 -360
rect 751 -356 752 -354
rect 751 -362 752 -360
rect 758 -356 759 -354
rect 758 -362 759 -360
rect 765 -356 766 -354
rect 765 -362 766 -360
rect 772 -362 773 -360
rect 775 -362 776 -360
rect 779 -356 780 -354
rect 779 -362 780 -360
rect 786 -356 787 -354
rect 789 -362 790 -360
rect 793 -356 794 -354
rect 793 -362 794 -360
rect 800 -356 801 -354
rect 800 -362 801 -360
rect 807 -356 808 -354
rect 807 -362 808 -360
rect 814 -356 815 -354
rect 814 -362 815 -360
rect 821 -356 822 -354
rect 821 -362 822 -360
rect 828 -356 829 -354
rect 828 -362 829 -360
rect 835 -356 836 -354
rect 835 -362 836 -360
rect 842 -356 843 -354
rect 842 -362 843 -360
rect 849 -356 850 -354
rect 849 -362 850 -360
rect 856 -356 857 -354
rect 856 -362 857 -360
rect 863 -356 864 -354
rect 863 -362 864 -360
rect 870 -356 871 -354
rect 870 -362 871 -360
rect 877 -356 878 -354
rect 877 -362 878 -360
rect 884 -356 885 -354
rect 884 -362 885 -360
rect 891 -356 892 -354
rect 891 -362 892 -360
rect 898 -356 899 -354
rect 898 -362 899 -360
rect 905 -356 906 -354
rect 905 -362 906 -360
rect 912 -356 913 -354
rect 912 -362 913 -360
rect 919 -356 920 -354
rect 919 -362 920 -360
rect 926 -356 927 -354
rect 926 -362 927 -360
rect 933 -356 934 -354
rect 933 -362 934 -360
rect 940 -356 941 -354
rect 940 -362 941 -360
rect 947 -356 948 -354
rect 947 -362 948 -360
rect 954 -356 955 -354
rect 954 -362 955 -360
rect 961 -356 962 -354
rect 961 -362 962 -360
rect 968 -356 969 -354
rect 968 -362 969 -360
rect 975 -356 976 -354
rect 975 -362 976 -360
rect 982 -356 983 -354
rect 982 -362 983 -360
rect 989 -356 990 -354
rect 989 -362 990 -360
rect 996 -356 997 -354
rect 996 -362 997 -360
rect 1003 -356 1004 -354
rect 1003 -362 1004 -360
rect 1010 -356 1011 -354
rect 1010 -362 1011 -360
rect 1017 -356 1018 -354
rect 1017 -362 1018 -360
rect 1024 -356 1025 -354
rect 1024 -362 1025 -360
rect 1031 -356 1032 -354
rect 1031 -362 1032 -360
rect 1038 -356 1039 -354
rect 1038 -362 1039 -360
rect 1045 -356 1046 -354
rect 1045 -362 1046 -360
rect 1052 -356 1053 -354
rect 1052 -362 1053 -360
rect 1059 -356 1060 -354
rect 1059 -362 1060 -360
rect 1066 -356 1067 -354
rect 1066 -362 1067 -360
rect 1073 -356 1074 -354
rect 1073 -362 1074 -360
rect 1080 -356 1081 -354
rect 1080 -362 1081 -360
rect 1087 -356 1088 -354
rect 1087 -362 1088 -360
rect 1094 -356 1095 -354
rect 1094 -362 1095 -360
rect 1101 -356 1102 -354
rect 1101 -362 1102 -360
rect 1108 -356 1109 -354
rect 1108 -362 1109 -360
rect 1115 -356 1116 -354
rect 1115 -362 1116 -360
rect 1122 -356 1123 -354
rect 1122 -362 1123 -360
rect 1129 -356 1130 -354
rect 1129 -362 1130 -360
rect 1136 -356 1137 -354
rect 1136 -362 1137 -360
rect 1143 -356 1144 -354
rect 1143 -362 1144 -360
rect 1150 -356 1151 -354
rect 1150 -362 1151 -360
rect 1157 -356 1158 -354
rect 1157 -362 1158 -360
rect 1164 -356 1165 -354
rect 1164 -362 1165 -360
rect 1171 -356 1172 -354
rect 1171 -362 1172 -360
rect 1178 -356 1179 -354
rect 1178 -362 1179 -360
rect 1185 -356 1186 -354
rect 1185 -362 1186 -360
rect 1192 -356 1193 -354
rect 1192 -362 1193 -360
rect 1199 -356 1200 -354
rect 1199 -362 1200 -360
rect 1206 -356 1207 -354
rect 1206 -362 1207 -360
rect 1213 -356 1214 -354
rect 1213 -362 1214 -360
rect 1220 -356 1221 -354
rect 1220 -362 1221 -360
rect 1227 -356 1228 -354
rect 1227 -362 1228 -360
rect 1234 -356 1235 -354
rect 1234 -362 1235 -360
rect 1241 -356 1242 -354
rect 1241 -362 1242 -360
rect 1248 -356 1249 -354
rect 1248 -362 1249 -360
rect 1255 -356 1256 -354
rect 1255 -362 1256 -360
rect 1262 -356 1263 -354
rect 1262 -362 1263 -360
rect 1269 -356 1270 -354
rect 1269 -362 1270 -360
rect 1276 -356 1277 -354
rect 1276 -362 1277 -360
rect 1283 -356 1284 -354
rect 1283 -362 1284 -360
rect 1290 -356 1291 -354
rect 1290 -362 1291 -360
rect 1300 -362 1301 -360
rect 40 -487 41 -485
rect 65 -481 66 -479
rect 65 -487 66 -485
rect 72 -481 73 -479
rect 72 -487 73 -485
rect 79 -481 80 -479
rect 79 -487 80 -485
rect 86 -481 87 -479
rect 86 -487 87 -485
rect 96 -481 97 -479
rect 93 -487 94 -485
rect 96 -487 97 -485
rect 100 -481 101 -479
rect 100 -487 101 -485
rect 107 -481 108 -479
rect 107 -487 108 -485
rect 124 -481 125 -479
rect 121 -487 122 -485
rect 124 -487 125 -485
rect 128 -481 129 -479
rect 131 -481 132 -479
rect 128 -487 129 -485
rect 131 -487 132 -485
rect 135 -481 136 -479
rect 135 -487 136 -485
rect 142 -481 143 -479
rect 142 -487 143 -485
rect 149 -481 150 -479
rect 152 -481 153 -479
rect 149 -487 150 -485
rect 152 -487 153 -485
rect 156 -481 157 -479
rect 156 -487 157 -485
rect 163 -481 164 -479
rect 163 -487 164 -485
rect 170 -481 171 -479
rect 170 -487 171 -485
rect 177 -481 178 -479
rect 177 -487 178 -485
rect 184 -481 185 -479
rect 184 -487 185 -485
rect 191 -481 192 -479
rect 191 -487 192 -485
rect 198 -481 199 -479
rect 198 -487 199 -485
rect 205 -481 206 -479
rect 205 -487 206 -485
rect 212 -481 213 -479
rect 215 -481 216 -479
rect 215 -487 216 -485
rect 219 -481 220 -479
rect 219 -487 220 -485
rect 226 -481 227 -479
rect 226 -487 227 -485
rect 233 -481 234 -479
rect 233 -487 234 -485
rect 240 -481 241 -479
rect 240 -487 241 -485
rect 247 -481 248 -479
rect 247 -487 248 -485
rect 254 -481 255 -479
rect 254 -487 255 -485
rect 261 -481 262 -479
rect 261 -487 262 -485
rect 268 -481 269 -479
rect 268 -487 269 -485
rect 296 -481 297 -479
rect 296 -487 297 -485
rect 303 -481 304 -479
rect 303 -487 304 -485
rect 310 -481 311 -479
rect 310 -487 311 -485
rect 317 -481 318 -479
rect 317 -487 318 -485
rect 324 -481 325 -479
rect 324 -487 325 -485
rect 331 -481 332 -479
rect 331 -487 332 -485
rect 338 -481 339 -479
rect 338 -487 339 -485
rect 345 -481 346 -479
rect 345 -487 346 -485
rect 352 -481 353 -479
rect 355 -481 356 -479
rect 355 -487 356 -485
rect 359 -481 360 -479
rect 359 -487 360 -485
rect 366 -481 367 -479
rect 366 -487 367 -485
rect 373 -481 374 -479
rect 373 -487 374 -485
rect 380 -481 381 -479
rect 380 -487 381 -485
rect 387 -481 388 -479
rect 387 -487 388 -485
rect 394 -481 395 -479
rect 394 -487 395 -485
rect 401 -481 402 -479
rect 401 -487 402 -485
rect 408 -481 409 -479
rect 408 -487 409 -485
rect 415 -481 416 -479
rect 415 -487 416 -485
rect 422 -481 423 -479
rect 422 -487 423 -485
rect 429 -481 430 -479
rect 429 -487 430 -485
rect 436 -481 437 -479
rect 436 -487 437 -485
rect 443 -481 444 -479
rect 443 -487 444 -485
rect 450 -481 451 -479
rect 450 -487 451 -485
rect 457 -481 458 -479
rect 460 -481 461 -479
rect 457 -487 458 -485
rect 460 -487 461 -485
rect 464 -481 465 -479
rect 464 -487 465 -485
rect 471 -481 472 -479
rect 471 -487 472 -485
rect 478 -481 479 -479
rect 478 -487 479 -485
rect 485 -481 486 -479
rect 485 -487 486 -485
rect 492 -481 493 -479
rect 492 -487 493 -485
rect 499 -481 500 -479
rect 502 -481 503 -479
rect 499 -487 500 -485
rect 502 -487 503 -485
rect 506 -481 507 -479
rect 506 -487 507 -485
rect 513 -481 514 -479
rect 516 -481 517 -479
rect 513 -487 514 -485
rect 520 -481 521 -479
rect 520 -487 521 -485
rect 527 -481 528 -479
rect 527 -487 528 -485
rect 534 -481 535 -479
rect 537 -481 538 -479
rect 534 -487 535 -485
rect 537 -487 538 -485
rect 541 -481 542 -479
rect 541 -487 542 -485
rect 548 -481 549 -479
rect 548 -487 549 -485
rect 555 -481 556 -479
rect 558 -481 559 -479
rect 555 -487 556 -485
rect 562 -481 563 -479
rect 562 -487 563 -485
rect 569 -481 570 -479
rect 569 -487 570 -485
rect 576 -481 577 -479
rect 579 -481 580 -479
rect 579 -487 580 -485
rect 583 -481 584 -479
rect 583 -487 584 -485
rect 590 -481 591 -479
rect 590 -487 591 -485
rect 597 -481 598 -479
rect 597 -487 598 -485
rect 600 -487 601 -485
rect 604 -481 605 -479
rect 604 -487 605 -485
rect 611 -481 612 -479
rect 614 -481 615 -479
rect 611 -487 612 -485
rect 614 -487 615 -485
rect 618 -481 619 -479
rect 618 -487 619 -485
rect 625 -481 626 -479
rect 625 -487 626 -485
rect 632 -481 633 -479
rect 635 -481 636 -479
rect 632 -487 633 -485
rect 635 -487 636 -485
rect 639 -481 640 -479
rect 642 -481 643 -479
rect 639 -487 640 -485
rect 646 -481 647 -479
rect 646 -487 647 -485
rect 653 -481 654 -479
rect 653 -487 654 -485
rect 660 -481 661 -479
rect 660 -487 661 -485
rect 667 -481 668 -479
rect 667 -487 668 -485
rect 674 -481 675 -479
rect 677 -481 678 -479
rect 674 -487 675 -485
rect 684 -481 685 -479
rect 684 -487 685 -485
rect 688 -481 689 -479
rect 688 -487 689 -485
rect 695 -481 696 -479
rect 695 -487 696 -485
rect 702 -481 703 -479
rect 702 -487 703 -485
rect 709 -481 710 -479
rect 709 -487 710 -485
rect 716 -481 717 -479
rect 719 -481 720 -479
rect 716 -487 717 -485
rect 719 -487 720 -485
rect 723 -481 724 -479
rect 723 -487 724 -485
rect 730 -481 731 -479
rect 730 -487 731 -485
rect 737 -481 738 -479
rect 737 -487 738 -485
rect 744 -481 745 -479
rect 744 -487 745 -485
rect 754 -481 755 -479
rect 751 -487 752 -485
rect 754 -487 755 -485
rect 758 -481 759 -479
rect 758 -487 759 -485
rect 761 -487 762 -485
rect 765 -481 766 -479
rect 765 -487 766 -485
rect 772 -487 773 -485
rect 779 -481 780 -479
rect 779 -487 780 -485
rect 786 -481 787 -479
rect 789 -481 790 -479
rect 786 -487 787 -485
rect 789 -487 790 -485
rect 793 -481 794 -479
rect 793 -487 794 -485
rect 800 -481 801 -479
rect 800 -487 801 -485
rect 807 -481 808 -479
rect 807 -487 808 -485
rect 814 -481 815 -479
rect 814 -487 815 -485
rect 821 -481 822 -479
rect 821 -487 822 -485
rect 831 -481 832 -479
rect 828 -487 829 -485
rect 831 -487 832 -485
rect 835 -481 836 -479
rect 835 -487 836 -485
rect 842 -481 843 -479
rect 842 -487 843 -485
rect 849 -481 850 -479
rect 849 -487 850 -485
rect 856 -481 857 -479
rect 856 -487 857 -485
rect 863 -481 864 -479
rect 863 -487 864 -485
rect 870 -481 871 -479
rect 870 -487 871 -485
rect 877 -481 878 -479
rect 877 -487 878 -485
rect 884 -481 885 -479
rect 887 -481 888 -479
rect 884 -487 885 -485
rect 887 -487 888 -485
rect 891 -481 892 -479
rect 891 -487 892 -485
rect 898 -481 899 -479
rect 898 -487 899 -485
rect 905 -481 906 -479
rect 905 -487 906 -485
rect 912 -481 913 -479
rect 912 -487 913 -485
rect 919 -481 920 -479
rect 919 -487 920 -485
rect 926 -481 927 -479
rect 926 -487 927 -485
rect 933 -481 934 -479
rect 933 -487 934 -485
rect 940 -481 941 -479
rect 940 -487 941 -485
rect 947 -481 948 -479
rect 947 -487 948 -485
rect 954 -481 955 -479
rect 954 -487 955 -485
rect 961 -481 962 -479
rect 961 -487 962 -485
rect 968 -481 969 -479
rect 968 -487 969 -485
rect 975 -481 976 -479
rect 975 -487 976 -485
rect 982 -481 983 -479
rect 982 -487 983 -485
rect 989 -481 990 -479
rect 989 -487 990 -485
rect 996 -481 997 -479
rect 996 -487 997 -485
rect 1003 -481 1004 -479
rect 1003 -487 1004 -485
rect 1010 -481 1011 -479
rect 1010 -487 1011 -485
rect 1017 -481 1018 -479
rect 1017 -487 1018 -485
rect 1024 -481 1025 -479
rect 1024 -487 1025 -485
rect 1031 -481 1032 -479
rect 1031 -487 1032 -485
rect 1038 -481 1039 -479
rect 1038 -487 1039 -485
rect 1045 -481 1046 -479
rect 1045 -487 1046 -485
rect 1052 -481 1053 -479
rect 1052 -487 1053 -485
rect 1059 -481 1060 -479
rect 1059 -487 1060 -485
rect 1066 -481 1067 -479
rect 1066 -487 1067 -485
rect 1073 -481 1074 -479
rect 1073 -487 1074 -485
rect 1080 -481 1081 -479
rect 1080 -487 1081 -485
rect 1087 -481 1088 -479
rect 1087 -487 1088 -485
rect 1094 -481 1095 -479
rect 1094 -487 1095 -485
rect 1101 -481 1102 -479
rect 1101 -487 1102 -485
rect 1108 -481 1109 -479
rect 1108 -487 1109 -485
rect 1115 -481 1116 -479
rect 1115 -487 1116 -485
rect 1122 -481 1123 -479
rect 1122 -487 1123 -485
rect 1129 -481 1130 -479
rect 1129 -487 1130 -485
rect 1136 -481 1137 -479
rect 1136 -487 1137 -485
rect 1143 -481 1144 -479
rect 1143 -487 1144 -485
rect 1150 -481 1151 -479
rect 1150 -487 1151 -485
rect 1157 -481 1158 -479
rect 1157 -487 1158 -485
rect 1164 -481 1165 -479
rect 1164 -487 1165 -485
rect 1171 -481 1172 -479
rect 1171 -487 1172 -485
rect 1178 -481 1179 -479
rect 1178 -487 1179 -485
rect 1185 -481 1186 -479
rect 1185 -487 1186 -485
rect 1192 -481 1193 -479
rect 1192 -487 1193 -485
rect 1199 -481 1200 -479
rect 1199 -487 1200 -485
rect 1206 -481 1207 -479
rect 1206 -487 1207 -485
rect 1213 -481 1214 -479
rect 1213 -487 1214 -485
rect 1220 -481 1221 -479
rect 1220 -487 1221 -485
rect 1227 -481 1228 -479
rect 1227 -487 1228 -485
rect 1234 -481 1235 -479
rect 1234 -487 1235 -485
rect 1241 -481 1242 -479
rect 1241 -487 1242 -485
rect 1248 -481 1249 -479
rect 1248 -487 1249 -485
rect 1255 -481 1256 -479
rect 1255 -487 1256 -485
rect 1262 -481 1263 -479
rect 1262 -487 1263 -485
rect 1269 -481 1270 -479
rect 1269 -487 1270 -485
rect 1276 -481 1277 -479
rect 1276 -487 1277 -485
rect 1283 -481 1284 -479
rect 1283 -487 1284 -485
rect 1290 -481 1291 -479
rect 1290 -487 1291 -485
rect 1297 -481 1298 -479
rect 1297 -487 1298 -485
rect 1304 -481 1305 -479
rect 1304 -487 1305 -485
rect 1311 -481 1312 -479
rect 1311 -487 1312 -485
rect 1318 -481 1319 -479
rect 1318 -487 1319 -485
rect 1325 -481 1326 -479
rect 1325 -487 1326 -485
rect 1332 -481 1333 -479
rect 1332 -487 1333 -485
rect 1339 -481 1340 -479
rect 1339 -487 1340 -485
rect 1346 -481 1347 -479
rect 1346 -487 1347 -485
rect 1353 -481 1354 -479
rect 1353 -487 1354 -485
rect 1360 -481 1361 -479
rect 1360 -487 1361 -485
rect 1367 -481 1368 -479
rect 1367 -487 1368 -485
rect 1374 -481 1375 -479
rect 1377 -487 1378 -485
rect 40 -614 41 -612
rect 51 -614 52 -612
rect 51 -620 52 -618
rect 58 -614 59 -612
rect 58 -620 59 -618
rect 65 -614 66 -612
rect 68 -614 69 -612
rect 65 -620 66 -618
rect 68 -620 69 -618
rect 72 -614 73 -612
rect 72 -620 73 -618
rect 79 -614 80 -612
rect 82 -620 83 -618
rect 86 -614 87 -612
rect 86 -620 87 -618
rect 100 -614 101 -612
rect 100 -620 101 -618
rect 107 -614 108 -612
rect 107 -620 108 -618
rect 114 -614 115 -612
rect 117 -620 118 -618
rect 121 -614 122 -612
rect 121 -620 122 -618
rect 128 -614 129 -612
rect 128 -620 129 -618
rect 135 -614 136 -612
rect 135 -620 136 -618
rect 138 -620 139 -618
rect 142 -614 143 -612
rect 142 -620 143 -618
rect 149 -614 150 -612
rect 152 -614 153 -612
rect 149 -620 150 -618
rect 152 -620 153 -618
rect 156 -614 157 -612
rect 159 -614 160 -612
rect 156 -620 157 -618
rect 159 -620 160 -618
rect 163 -614 164 -612
rect 163 -620 164 -618
rect 177 -614 178 -612
rect 177 -620 178 -618
rect 184 -614 185 -612
rect 184 -620 185 -618
rect 191 -614 192 -612
rect 191 -620 192 -618
rect 198 -614 199 -612
rect 198 -620 199 -618
rect 201 -620 202 -618
rect 205 -614 206 -612
rect 205 -620 206 -618
rect 212 -614 213 -612
rect 212 -620 213 -618
rect 219 -614 220 -612
rect 222 -614 223 -612
rect 219 -620 220 -618
rect 226 -614 227 -612
rect 226 -620 227 -618
rect 243 -614 244 -612
rect 243 -620 244 -618
rect 250 -614 251 -612
rect 247 -620 248 -618
rect 250 -620 251 -618
rect 261 -614 262 -612
rect 261 -620 262 -618
rect 268 -614 269 -612
rect 268 -620 269 -618
rect 275 -614 276 -612
rect 275 -620 276 -618
rect 282 -614 283 -612
rect 282 -620 283 -618
rect 289 -614 290 -612
rect 289 -620 290 -618
rect 296 -614 297 -612
rect 296 -620 297 -618
rect 303 -614 304 -612
rect 303 -620 304 -618
rect 310 -614 311 -612
rect 310 -620 311 -618
rect 317 -614 318 -612
rect 317 -620 318 -618
rect 324 -614 325 -612
rect 324 -620 325 -618
rect 331 -614 332 -612
rect 331 -620 332 -618
rect 338 -614 339 -612
rect 338 -620 339 -618
rect 345 -614 346 -612
rect 345 -620 346 -618
rect 352 -614 353 -612
rect 352 -620 353 -618
rect 359 -614 360 -612
rect 359 -620 360 -618
rect 373 -614 374 -612
rect 373 -620 374 -618
rect 380 -614 381 -612
rect 380 -620 381 -618
rect 387 -614 388 -612
rect 387 -620 388 -618
rect 394 -614 395 -612
rect 397 -614 398 -612
rect 394 -620 395 -618
rect 397 -620 398 -618
rect 401 -614 402 -612
rect 401 -620 402 -618
rect 408 -614 409 -612
rect 408 -620 409 -618
rect 415 -614 416 -612
rect 415 -620 416 -618
rect 422 -614 423 -612
rect 422 -620 423 -618
rect 429 -614 430 -612
rect 429 -620 430 -618
rect 436 -614 437 -612
rect 436 -620 437 -618
rect 443 -614 444 -612
rect 443 -620 444 -618
rect 450 -614 451 -612
rect 450 -620 451 -618
rect 457 -614 458 -612
rect 457 -620 458 -618
rect 464 -614 465 -612
rect 464 -620 465 -618
rect 471 -614 472 -612
rect 471 -620 472 -618
rect 478 -614 479 -612
rect 478 -620 479 -618
rect 485 -614 486 -612
rect 485 -620 486 -618
rect 492 -614 493 -612
rect 492 -620 493 -618
rect 499 -614 500 -612
rect 502 -614 503 -612
rect 502 -620 503 -618
rect 506 -614 507 -612
rect 506 -620 507 -618
rect 513 -614 514 -612
rect 513 -620 514 -618
rect 516 -620 517 -618
rect 520 -614 521 -612
rect 520 -620 521 -618
rect 527 -614 528 -612
rect 530 -614 531 -612
rect 527 -620 528 -618
rect 530 -620 531 -618
rect 534 -614 535 -612
rect 534 -620 535 -618
rect 541 -614 542 -612
rect 544 -614 545 -612
rect 541 -620 542 -618
rect 548 -614 549 -612
rect 548 -620 549 -618
rect 555 -614 556 -612
rect 555 -620 556 -618
rect 562 -614 563 -612
rect 562 -620 563 -618
rect 569 -614 570 -612
rect 569 -620 570 -618
rect 576 -614 577 -612
rect 576 -620 577 -618
rect 583 -614 584 -612
rect 586 -614 587 -612
rect 583 -620 584 -618
rect 586 -620 587 -618
rect 590 -614 591 -612
rect 590 -620 591 -618
rect 597 -614 598 -612
rect 597 -620 598 -618
rect 604 -614 605 -612
rect 604 -620 605 -618
rect 611 -614 612 -612
rect 611 -620 612 -618
rect 618 -614 619 -612
rect 618 -620 619 -618
rect 625 -614 626 -612
rect 625 -620 626 -618
rect 632 -614 633 -612
rect 632 -620 633 -618
rect 639 -614 640 -612
rect 639 -620 640 -618
rect 646 -614 647 -612
rect 646 -620 647 -618
rect 653 -614 654 -612
rect 653 -620 654 -618
rect 660 -614 661 -612
rect 660 -620 661 -618
rect 670 -614 671 -612
rect 667 -620 668 -618
rect 670 -620 671 -618
rect 674 -614 675 -612
rect 674 -620 675 -618
rect 681 -614 682 -612
rect 684 -614 685 -612
rect 684 -620 685 -618
rect 688 -614 689 -612
rect 688 -620 689 -618
rect 695 -614 696 -612
rect 698 -614 699 -612
rect 695 -620 696 -618
rect 698 -620 699 -618
rect 702 -614 703 -612
rect 705 -614 706 -612
rect 702 -620 703 -618
rect 705 -620 706 -618
rect 709 -614 710 -612
rect 709 -620 710 -618
rect 716 -614 717 -612
rect 716 -620 717 -618
rect 719 -620 720 -618
rect 723 -614 724 -612
rect 723 -620 724 -618
rect 730 -614 731 -612
rect 733 -614 734 -612
rect 733 -620 734 -618
rect 737 -614 738 -612
rect 737 -620 738 -618
rect 744 -614 745 -612
rect 744 -620 745 -618
rect 751 -614 752 -612
rect 751 -620 752 -618
rect 758 -614 759 -612
rect 758 -620 759 -618
rect 765 -614 766 -612
rect 768 -614 769 -612
rect 765 -620 766 -618
rect 768 -620 769 -618
rect 775 -614 776 -612
rect 772 -620 773 -618
rect 775 -620 776 -618
rect 779 -614 780 -612
rect 782 -614 783 -612
rect 779 -620 780 -618
rect 786 -614 787 -612
rect 786 -620 787 -618
rect 793 -614 794 -612
rect 793 -620 794 -618
rect 796 -620 797 -618
rect 800 -614 801 -612
rect 800 -620 801 -618
rect 807 -614 808 -612
rect 810 -614 811 -612
rect 807 -620 808 -618
rect 814 -614 815 -612
rect 814 -620 815 -618
rect 821 -614 822 -612
rect 821 -620 822 -618
rect 828 -614 829 -612
rect 828 -620 829 -618
rect 835 -614 836 -612
rect 835 -620 836 -618
rect 842 -614 843 -612
rect 842 -620 843 -618
rect 849 -614 850 -612
rect 849 -620 850 -618
rect 856 -614 857 -612
rect 856 -620 857 -618
rect 863 -614 864 -612
rect 863 -620 864 -618
rect 870 -614 871 -612
rect 870 -620 871 -618
rect 877 -614 878 -612
rect 877 -620 878 -618
rect 884 -614 885 -612
rect 884 -620 885 -618
rect 891 -614 892 -612
rect 891 -620 892 -618
rect 898 -614 899 -612
rect 901 -614 902 -612
rect 898 -620 899 -618
rect 901 -620 902 -618
rect 905 -614 906 -612
rect 905 -620 906 -618
rect 912 -614 913 -612
rect 912 -620 913 -618
rect 919 -614 920 -612
rect 919 -620 920 -618
rect 926 -614 927 -612
rect 926 -620 927 -618
rect 933 -614 934 -612
rect 933 -620 934 -618
rect 940 -614 941 -612
rect 940 -620 941 -618
rect 947 -614 948 -612
rect 947 -620 948 -618
rect 954 -614 955 -612
rect 954 -620 955 -618
rect 961 -614 962 -612
rect 961 -620 962 -618
rect 968 -614 969 -612
rect 968 -620 969 -618
rect 975 -614 976 -612
rect 978 -614 979 -612
rect 978 -620 979 -618
rect 982 -614 983 -612
rect 982 -620 983 -618
rect 989 -614 990 -612
rect 989 -620 990 -618
rect 996 -614 997 -612
rect 996 -620 997 -618
rect 1003 -614 1004 -612
rect 1003 -620 1004 -618
rect 1010 -614 1011 -612
rect 1010 -620 1011 -618
rect 1017 -614 1018 -612
rect 1017 -620 1018 -618
rect 1024 -614 1025 -612
rect 1024 -620 1025 -618
rect 1031 -614 1032 -612
rect 1031 -620 1032 -618
rect 1038 -614 1039 -612
rect 1038 -620 1039 -618
rect 1045 -614 1046 -612
rect 1045 -620 1046 -618
rect 1052 -614 1053 -612
rect 1052 -620 1053 -618
rect 1059 -614 1060 -612
rect 1059 -620 1060 -618
rect 1066 -614 1067 -612
rect 1066 -620 1067 -618
rect 1073 -614 1074 -612
rect 1073 -620 1074 -618
rect 1080 -614 1081 -612
rect 1080 -620 1081 -618
rect 1087 -614 1088 -612
rect 1087 -620 1088 -618
rect 1094 -614 1095 -612
rect 1094 -620 1095 -618
rect 1101 -614 1102 -612
rect 1101 -620 1102 -618
rect 1108 -614 1109 -612
rect 1108 -620 1109 -618
rect 1115 -614 1116 -612
rect 1115 -620 1116 -618
rect 1122 -614 1123 -612
rect 1122 -620 1123 -618
rect 1129 -614 1130 -612
rect 1129 -620 1130 -618
rect 1136 -614 1137 -612
rect 1136 -620 1137 -618
rect 1143 -614 1144 -612
rect 1143 -620 1144 -618
rect 1150 -614 1151 -612
rect 1150 -620 1151 -618
rect 1157 -614 1158 -612
rect 1157 -620 1158 -618
rect 1164 -614 1165 -612
rect 1164 -620 1165 -618
rect 1171 -614 1172 -612
rect 1171 -620 1172 -618
rect 1178 -614 1179 -612
rect 1178 -620 1179 -618
rect 1185 -614 1186 -612
rect 1185 -620 1186 -618
rect 1192 -614 1193 -612
rect 1192 -620 1193 -618
rect 1199 -614 1200 -612
rect 1199 -620 1200 -618
rect 1206 -614 1207 -612
rect 1206 -620 1207 -618
rect 1213 -614 1214 -612
rect 1213 -620 1214 -618
rect 1220 -614 1221 -612
rect 1220 -620 1221 -618
rect 1227 -614 1228 -612
rect 1227 -620 1228 -618
rect 1234 -614 1235 -612
rect 1234 -620 1235 -618
rect 1241 -614 1242 -612
rect 1241 -620 1242 -618
rect 1248 -614 1249 -612
rect 1248 -620 1249 -618
rect 1255 -614 1256 -612
rect 1255 -620 1256 -618
rect 1262 -614 1263 -612
rect 1262 -620 1263 -618
rect 1269 -614 1270 -612
rect 1269 -620 1270 -618
rect 1276 -614 1277 -612
rect 1276 -620 1277 -618
rect 1283 -614 1284 -612
rect 1283 -620 1284 -618
rect 1290 -614 1291 -612
rect 1290 -620 1291 -618
rect 1297 -614 1298 -612
rect 1297 -620 1298 -618
rect 1304 -614 1305 -612
rect 1304 -620 1305 -618
rect 1311 -614 1312 -612
rect 1311 -620 1312 -618
rect 1318 -614 1319 -612
rect 1318 -620 1319 -618
rect 1325 -614 1326 -612
rect 1325 -620 1326 -618
rect 1332 -614 1333 -612
rect 1332 -620 1333 -618
rect 1339 -614 1340 -612
rect 1339 -620 1340 -618
rect 1346 -614 1347 -612
rect 1346 -620 1347 -618
rect 1353 -614 1354 -612
rect 1353 -620 1354 -618
rect 1356 -620 1357 -618
rect 1360 -614 1361 -612
rect 1360 -620 1361 -618
rect 1367 -614 1368 -612
rect 1367 -620 1368 -618
rect 1374 -614 1375 -612
rect 1374 -620 1375 -618
rect 1381 -614 1382 -612
rect 1381 -620 1382 -618
rect 1388 -614 1389 -612
rect 1388 -620 1389 -618
rect 1472 -614 1473 -612
rect 1472 -620 1473 -618
rect 44 -737 45 -735
rect 44 -743 45 -741
rect 51 -737 52 -735
rect 51 -743 52 -741
rect 58 -737 59 -735
rect 58 -743 59 -741
rect 65 -737 66 -735
rect 65 -743 66 -741
rect 72 -737 73 -735
rect 72 -743 73 -741
rect 82 -737 83 -735
rect 79 -743 80 -741
rect 82 -743 83 -741
rect 86 -737 87 -735
rect 86 -743 87 -741
rect 93 -737 94 -735
rect 96 -737 97 -735
rect 93 -743 94 -741
rect 100 -737 101 -735
rect 100 -743 101 -741
rect 107 -737 108 -735
rect 107 -743 108 -741
rect 114 -737 115 -735
rect 114 -743 115 -741
rect 121 -737 122 -735
rect 124 -737 125 -735
rect 121 -743 122 -741
rect 124 -743 125 -741
rect 128 -737 129 -735
rect 128 -743 129 -741
rect 135 -737 136 -735
rect 135 -743 136 -741
rect 149 -737 150 -735
rect 149 -743 150 -741
rect 156 -737 157 -735
rect 156 -743 157 -741
rect 163 -737 164 -735
rect 163 -743 164 -741
rect 170 -737 171 -735
rect 170 -743 171 -741
rect 177 -737 178 -735
rect 177 -743 178 -741
rect 184 -737 185 -735
rect 187 -737 188 -735
rect 184 -743 185 -741
rect 187 -743 188 -741
rect 191 -737 192 -735
rect 191 -743 192 -741
rect 198 -737 199 -735
rect 198 -743 199 -741
rect 205 -737 206 -735
rect 205 -743 206 -741
rect 212 -737 213 -735
rect 212 -743 213 -741
rect 219 -737 220 -735
rect 219 -743 220 -741
rect 226 -737 227 -735
rect 226 -743 227 -741
rect 233 -737 234 -735
rect 233 -743 234 -741
rect 240 -737 241 -735
rect 240 -743 241 -741
rect 247 -737 248 -735
rect 250 -737 251 -735
rect 250 -743 251 -741
rect 254 -737 255 -735
rect 254 -743 255 -741
rect 261 -737 262 -735
rect 261 -743 262 -741
rect 268 -737 269 -735
rect 268 -743 269 -741
rect 275 -737 276 -735
rect 275 -743 276 -741
rect 282 -737 283 -735
rect 282 -743 283 -741
rect 292 -737 293 -735
rect 289 -743 290 -741
rect 292 -743 293 -741
rect 296 -737 297 -735
rect 296 -743 297 -741
rect 303 -737 304 -735
rect 303 -743 304 -741
rect 310 -737 311 -735
rect 310 -743 311 -741
rect 317 -737 318 -735
rect 317 -743 318 -741
rect 324 -737 325 -735
rect 324 -743 325 -741
rect 331 -737 332 -735
rect 331 -743 332 -741
rect 338 -737 339 -735
rect 338 -743 339 -741
rect 345 -737 346 -735
rect 345 -743 346 -741
rect 352 -737 353 -735
rect 352 -743 353 -741
rect 359 -737 360 -735
rect 359 -743 360 -741
rect 366 -737 367 -735
rect 366 -743 367 -741
rect 373 -737 374 -735
rect 373 -743 374 -741
rect 380 -737 381 -735
rect 380 -743 381 -741
rect 387 -737 388 -735
rect 387 -743 388 -741
rect 394 -737 395 -735
rect 394 -743 395 -741
rect 401 -737 402 -735
rect 401 -743 402 -741
rect 408 -737 409 -735
rect 408 -743 409 -741
rect 415 -737 416 -735
rect 415 -743 416 -741
rect 422 -737 423 -735
rect 422 -743 423 -741
rect 429 -737 430 -735
rect 432 -737 433 -735
rect 429 -743 430 -741
rect 432 -743 433 -741
rect 436 -737 437 -735
rect 439 -737 440 -735
rect 436 -743 437 -741
rect 439 -743 440 -741
rect 443 -737 444 -735
rect 443 -743 444 -741
rect 450 -737 451 -735
rect 450 -743 451 -741
rect 457 -737 458 -735
rect 457 -743 458 -741
rect 464 -737 465 -735
rect 464 -743 465 -741
rect 471 -737 472 -735
rect 471 -743 472 -741
rect 478 -737 479 -735
rect 478 -743 479 -741
rect 488 -737 489 -735
rect 488 -743 489 -741
rect 492 -737 493 -735
rect 492 -743 493 -741
rect 506 -737 507 -735
rect 506 -743 507 -741
rect 513 -737 514 -735
rect 513 -743 514 -741
rect 520 -737 521 -735
rect 520 -743 521 -741
rect 527 -737 528 -735
rect 527 -743 528 -741
rect 534 -737 535 -735
rect 537 -737 538 -735
rect 534 -743 535 -741
rect 537 -743 538 -741
rect 541 -737 542 -735
rect 541 -743 542 -741
rect 548 -737 549 -735
rect 548 -743 549 -741
rect 555 -737 556 -735
rect 558 -737 559 -735
rect 555 -743 556 -741
rect 558 -743 559 -741
rect 562 -737 563 -735
rect 565 -737 566 -735
rect 562 -743 563 -741
rect 565 -743 566 -741
rect 569 -737 570 -735
rect 569 -743 570 -741
rect 576 -737 577 -735
rect 579 -737 580 -735
rect 576 -743 577 -741
rect 579 -743 580 -741
rect 583 -737 584 -735
rect 583 -743 584 -741
rect 590 -737 591 -735
rect 593 -737 594 -735
rect 590 -743 591 -741
rect 593 -743 594 -741
rect 597 -737 598 -735
rect 597 -743 598 -741
rect 604 -737 605 -735
rect 607 -737 608 -735
rect 607 -743 608 -741
rect 611 -737 612 -735
rect 611 -743 612 -741
rect 618 -737 619 -735
rect 618 -743 619 -741
rect 625 -737 626 -735
rect 625 -743 626 -741
rect 639 -737 640 -735
rect 639 -743 640 -741
rect 646 -737 647 -735
rect 649 -737 650 -735
rect 649 -743 650 -741
rect 653 -737 654 -735
rect 656 -737 657 -735
rect 653 -743 654 -741
rect 656 -743 657 -741
rect 660 -737 661 -735
rect 660 -743 661 -741
rect 667 -737 668 -735
rect 667 -743 668 -741
rect 674 -737 675 -735
rect 674 -743 675 -741
rect 681 -737 682 -735
rect 681 -743 682 -741
rect 688 -737 689 -735
rect 688 -743 689 -741
rect 695 -737 696 -735
rect 695 -743 696 -741
rect 702 -737 703 -735
rect 702 -743 703 -741
rect 709 -737 710 -735
rect 712 -737 713 -735
rect 709 -743 710 -741
rect 712 -743 713 -741
rect 716 -737 717 -735
rect 716 -743 717 -741
rect 723 -737 724 -735
rect 726 -737 727 -735
rect 723 -743 724 -741
rect 726 -743 727 -741
rect 730 -737 731 -735
rect 733 -737 734 -735
rect 730 -743 731 -741
rect 733 -743 734 -741
rect 737 -737 738 -735
rect 737 -743 738 -741
rect 744 -737 745 -735
rect 744 -743 745 -741
rect 751 -737 752 -735
rect 751 -743 752 -741
rect 758 -737 759 -735
rect 758 -743 759 -741
rect 765 -737 766 -735
rect 765 -743 766 -741
rect 772 -737 773 -735
rect 772 -743 773 -741
rect 779 -737 780 -735
rect 779 -743 780 -741
rect 786 -737 787 -735
rect 786 -743 787 -741
rect 793 -737 794 -735
rect 796 -743 797 -741
rect 800 -737 801 -735
rect 800 -743 801 -741
rect 807 -737 808 -735
rect 807 -743 808 -741
rect 814 -737 815 -735
rect 814 -743 815 -741
rect 821 -737 822 -735
rect 821 -743 822 -741
rect 828 -737 829 -735
rect 831 -737 832 -735
rect 828 -743 829 -741
rect 831 -743 832 -741
rect 835 -737 836 -735
rect 835 -743 836 -741
rect 842 -737 843 -735
rect 842 -743 843 -741
rect 849 -737 850 -735
rect 849 -743 850 -741
rect 856 -737 857 -735
rect 859 -737 860 -735
rect 856 -743 857 -741
rect 859 -743 860 -741
rect 863 -737 864 -735
rect 863 -743 864 -741
rect 870 -743 871 -741
rect 873 -743 874 -741
rect 877 -737 878 -735
rect 877 -743 878 -741
rect 884 -737 885 -735
rect 887 -737 888 -735
rect 884 -743 885 -741
rect 887 -743 888 -741
rect 891 -737 892 -735
rect 891 -743 892 -741
rect 898 -737 899 -735
rect 898 -743 899 -741
rect 905 -737 906 -735
rect 908 -737 909 -735
rect 905 -743 906 -741
rect 912 -737 913 -735
rect 912 -743 913 -741
rect 919 -737 920 -735
rect 919 -743 920 -741
rect 922 -743 923 -741
rect 926 -737 927 -735
rect 926 -743 927 -741
rect 933 -737 934 -735
rect 933 -743 934 -741
rect 940 -737 941 -735
rect 940 -743 941 -741
rect 947 -737 948 -735
rect 947 -743 948 -741
rect 954 -737 955 -735
rect 954 -743 955 -741
rect 961 -737 962 -735
rect 961 -743 962 -741
rect 968 -737 969 -735
rect 968 -743 969 -741
rect 975 -737 976 -735
rect 975 -743 976 -741
rect 982 -737 983 -735
rect 982 -743 983 -741
rect 992 -737 993 -735
rect 989 -743 990 -741
rect 992 -743 993 -741
rect 996 -737 997 -735
rect 996 -743 997 -741
rect 1006 -737 1007 -735
rect 1003 -743 1004 -741
rect 1006 -743 1007 -741
rect 1010 -737 1011 -735
rect 1010 -743 1011 -741
rect 1017 -737 1018 -735
rect 1017 -743 1018 -741
rect 1024 -737 1025 -735
rect 1024 -743 1025 -741
rect 1031 -737 1032 -735
rect 1031 -743 1032 -741
rect 1038 -737 1039 -735
rect 1038 -743 1039 -741
rect 1045 -737 1046 -735
rect 1045 -743 1046 -741
rect 1052 -737 1053 -735
rect 1052 -743 1053 -741
rect 1059 -737 1060 -735
rect 1062 -737 1063 -735
rect 1066 -737 1067 -735
rect 1066 -743 1067 -741
rect 1073 -737 1074 -735
rect 1073 -743 1074 -741
rect 1080 -737 1081 -735
rect 1080 -743 1081 -741
rect 1087 -737 1088 -735
rect 1087 -743 1088 -741
rect 1094 -737 1095 -735
rect 1094 -743 1095 -741
rect 1101 -737 1102 -735
rect 1101 -743 1102 -741
rect 1108 -737 1109 -735
rect 1108 -743 1109 -741
rect 1115 -737 1116 -735
rect 1115 -743 1116 -741
rect 1122 -737 1123 -735
rect 1122 -743 1123 -741
rect 1129 -737 1130 -735
rect 1129 -743 1130 -741
rect 1136 -737 1137 -735
rect 1136 -743 1137 -741
rect 1143 -737 1144 -735
rect 1143 -743 1144 -741
rect 1150 -737 1151 -735
rect 1150 -743 1151 -741
rect 1157 -737 1158 -735
rect 1157 -743 1158 -741
rect 1164 -737 1165 -735
rect 1164 -743 1165 -741
rect 1171 -737 1172 -735
rect 1171 -743 1172 -741
rect 1178 -737 1179 -735
rect 1178 -743 1179 -741
rect 1185 -737 1186 -735
rect 1185 -743 1186 -741
rect 1192 -737 1193 -735
rect 1192 -743 1193 -741
rect 1199 -737 1200 -735
rect 1199 -743 1200 -741
rect 1206 -737 1207 -735
rect 1206 -743 1207 -741
rect 1213 -737 1214 -735
rect 1213 -743 1214 -741
rect 1220 -737 1221 -735
rect 1220 -743 1221 -741
rect 1227 -737 1228 -735
rect 1227 -743 1228 -741
rect 1234 -737 1235 -735
rect 1234 -743 1235 -741
rect 1241 -737 1242 -735
rect 1241 -743 1242 -741
rect 1248 -737 1249 -735
rect 1248 -743 1249 -741
rect 1255 -737 1256 -735
rect 1255 -743 1256 -741
rect 1262 -737 1263 -735
rect 1262 -743 1263 -741
rect 1269 -737 1270 -735
rect 1269 -743 1270 -741
rect 1276 -737 1277 -735
rect 1276 -743 1277 -741
rect 1283 -737 1284 -735
rect 1283 -743 1284 -741
rect 1290 -737 1291 -735
rect 1290 -743 1291 -741
rect 1297 -737 1298 -735
rect 1297 -743 1298 -741
rect 1304 -737 1305 -735
rect 1304 -743 1305 -741
rect 1311 -737 1312 -735
rect 1311 -743 1312 -741
rect 1318 -737 1319 -735
rect 1318 -743 1319 -741
rect 1325 -737 1326 -735
rect 1325 -743 1326 -741
rect 1332 -737 1333 -735
rect 1332 -743 1333 -741
rect 1339 -737 1340 -735
rect 1339 -743 1340 -741
rect 1346 -737 1347 -735
rect 1346 -743 1347 -741
rect 1353 -737 1354 -735
rect 1353 -743 1354 -741
rect 1360 -737 1361 -735
rect 1360 -743 1361 -741
rect 1367 -737 1368 -735
rect 1367 -743 1368 -741
rect 1374 -737 1375 -735
rect 1374 -743 1375 -741
rect 1381 -737 1382 -735
rect 1381 -743 1382 -741
rect 1388 -737 1389 -735
rect 1388 -743 1389 -741
rect 1395 -737 1396 -735
rect 1395 -743 1396 -741
rect 1402 -737 1403 -735
rect 1402 -743 1403 -741
rect 1409 -737 1410 -735
rect 1409 -743 1410 -741
rect 1416 -737 1417 -735
rect 1416 -743 1417 -741
rect 1426 -737 1427 -735
rect 1423 -743 1424 -741
rect 1426 -743 1427 -741
rect 1430 -737 1431 -735
rect 1430 -743 1431 -741
rect 1500 -737 1501 -735
rect 1500 -743 1501 -741
rect 1521 -737 1522 -735
rect 1521 -743 1522 -741
rect 1570 -737 1571 -735
rect 1570 -743 1571 -741
rect 1633 -737 1634 -735
rect 1633 -743 1634 -741
rect 23 -876 24 -874
rect 23 -882 24 -880
rect 33 -876 34 -874
rect 37 -876 38 -874
rect 37 -882 38 -880
rect 44 -876 45 -874
rect 44 -882 45 -880
rect 51 -876 52 -874
rect 54 -882 55 -880
rect 58 -876 59 -874
rect 58 -882 59 -880
rect 65 -876 66 -874
rect 65 -882 66 -880
rect 72 -876 73 -874
rect 72 -882 73 -880
rect 79 -876 80 -874
rect 79 -882 80 -880
rect 86 -882 87 -880
rect 89 -882 90 -880
rect 93 -876 94 -874
rect 93 -882 94 -880
rect 100 -876 101 -874
rect 103 -876 104 -874
rect 100 -882 101 -880
rect 103 -882 104 -880
rect 107 -876 108 -874
rect 110 -876 111 -874
rect 107 -882 108 -880
rect 114 -876 115 -874
rect 114 -882 115 -880
rect 121 -876 122 -874
rect 121 -882 122 -880
rect 128 -876 129 -874
rect 128 -882 129 -880
rect 135 -876 136 -874
rect 138 -876 139 -874
rect 135 -882 136 -880
rect 138 -882 139 -880
rect 142 -876 143 -874
rect 142 -882 143 -880
rect 149 -876 150 -874
rect 149 -882 150 -880
rect 156 -876 157 -874
rect 156 -882 157 -880
rect 166 -876 167 -874
rect 163 -882 164 -880
rect 166 -882 167 -880
rect 170 -876 171 -874
rect 170 -882 171 -880
rect 177 -876 178 -874
rect 177 -882 178 -880
rect 184 -876 185 -874
rect 184 -882 185 -880
rect 191 -876 192 -874
rect 191 -882 192 -880
rect 198 -876 199 -874
rect 198 -882 199 -880
rect 205 -876 206 -874
rect 208 -882 209 -880
rect 212 -876 213 -874
rect 212 -882 213 -880
rect 219 -876 220 -874
rect 219 -882 220 -880
rect 229 -876 230 -874
rect 226 -882 227 -880
rect 229 -882 230 -880
rect 233 -876 234 -874
rect 236 -876 237 -874
rect 233 -882 234 -880
rect 236 -882 237 -880
rect 240 -876 241 -874
rect 240 -882 241 -880
rect 247 -876 248 -874
rect 250 -876 251 -874
rect 250 -882 251 -880
rect 254 -876 255 -874
rect 254 -882 255 -880
rect 261 -876 262 -874
rect 261 -882 262 -880
rect 268 -876 269 -874
rect 268 -882 269 -880
rect 275 -876 276 -874
rect 275 -882 276 -880
rect 282 -876 283 -874
rect 282 -882 283 -880
rect 289 -876 290 -874
rect 289 -882 290 -880
rect 303 -876 304 -874
rect 303 -882 304 -880
rect 310 -876 311 -874
rect 310 -882 311 -880
rect 324 -876 325 -874
rect 324 -882 325 -880
rect 331 -876 332 -874
rect 331 -882 332 -880
rect 338 -876 339 -874
rect 338 -882 339 -880
rect 345 -876 346 -874
rect 345 -882 346 -880
rect 352 -876 353 -874
rect 352 -882 353 -880
rect 359 -876 360 -874
rect 359 -882 360 -880
rect 366 -876 367 -874
rect 366 -882 367 -880
rect 373 -876 374 -874
rect 373 -882 374 -880
rect 380 -876 381 -874
rect 380 -882 381 -880
rect 387 -876 388 -874
rect 387 -882 388 -880
rect 394 -876 395 -874
rect 394 -882 395 -880
rect 401 -876 402 -874
rect 401 -882 402 -880
rect 408 -876 409 -874
rect 408 -882 409 -880
rect 415 -876 416 -874
rect 415 -882 416 -880
rect 422 -876 423 -874
rect 422 -882 423 -880
rect 429 -876 430 -874
rect 429 -882 430 -880
rect 436 -876 437 -874
rect 436 -882 437 -880
rect 443 -876 444 -874
rect 443 -882 444 -880
rect 450 -876 451 -874
rect 450 -882 451 -880
rect 457 -876 458 -874
rect 457 -882 458 -880
rect 464 -876 465 -874
rect 467 -876 468 -874
rect 467 -882 468 -880
rect 471 -876 472 -874
rect 471 -882 472 -880
rect 478 -876 479 -874
rect 478 -882 479 -880
rect 481 -882 482 -880
rect 485 -876 486 -874
rect 485 -882 486 -880
rect 492 -876 493 -874
rect 492 -882 493 -880
rect 499 -876 500 -874
rect 499 -882 500 -880
rect 506 -876 507 -874
rect 506 -882 507 -880
rect 513 -876 514 -874
rect 513 -882 514 -880
rect 520 -876 521 -874
rect 520 -882 521 -880
rect 527 -876 528 -874
rect 527 -882 528 -880
rect 534 -876 535 -874
rect 534 -882 535 -880
rect 541 -876 542 -874
rect 541 -882 542 -880
rect 548 -876 549 -874
rect 548 -882 549 -880
rect 555 -876 556 -874
rect 555 -882 556 -880
rect 562 -876 563 -874
rect 565 -876 566 -874
rect 562 -882 563 -880
rect 569 -876 570 -874
rect 569 -882 570 -880
rect 576 -876 577 -874
rect 576 -882 577 -880
rect 579 -882 580 -880
rect 583 -876 584 -874
rect 586 -876 587 -874
rect 583 -882 584 -880
rect 586 -882 587 -880
rect 590 -876 591 -874
rect 590 -882 591 -880
rect 597 -876 598 -874
rect 597 -882 598 -880
rect 604 -876 605 -874
rect 604 -882 605 -880
rect 611 -876 612 -874
rect 611 -882 612 -880
rect 614 -882 615 -880
rect 618 -876 619 -874
rect 618 -882 619 -880
rect 625 -876 626 -874
rect 628 -876 629 -874
rect 625 -882 626 -880
rect 628 -882 629 -880
rect 632 -876 633 -874
rect 632 -882 633 -880
rect 639 -876 640 -874
rect 642 -876 643 -874
rect 639 -882 640 -880
rect 646 -876 647 -874
rect 646 -882 647 -880
rect 660 -876 661 -874
rect 660 -882 661 -880
rect 663 -882 664 -880
rect 667 -876 668 -874
rect 667 -882 668 -880
rect 674 -876 675 -874
rect 674 -882 675 -880
rect 681 -876 682 -874
rect 681 -882 682 -880
rect 688 -876 689 -874
rect 691 -876 692 -874
rect 691 -882 692 -880
rect 695 -876 696 -874
rect 695 -882 696 -880
rect 702 -876 703 -874
rect 705 -882 706 -880
rect 709 -876 710 -874
rect 709 -882 710 -880
rect 716 -876 717 -874
rect 716 -882 717 -880
rect 723 -876 724 -874
rect 723 -882 724 -880
rect 730 -876 731 -874
rect 730 -882 731 -880
rect 737 -876 738 -874
rect 740 -876 741 -874
rect 737 -882 738 -880
rect 740 -882 741 -880
rect 744 -876 745 -874
rect 744 -882 745 -880
rect 751 -876 752 -874
rect 751 -882 752 -880
rect 758 -876 759 -874
rect 758 -882 759 -880
rect 761 -882 762 -880
rect 765 -876 766 -874
rect 765 -882 766 -880
rect 772 -876 773 -874
rect 772 -882 773 -880
rect 782 -876 783 -874
rect 779 -882 780 -880
rect 786 -876 787 -874
rect 789 -876 790 -874
rect 786 -882 787 -880
rect 789 -882 790 -880
rect 793 -876 794 -874
rect 793 -882 794 -880
rect 796 -882 797 -880
rect 800 -876 801 -874
rect 800 -882 801 -880
rect 807 -876 808 -874
rect 807 -882 808 -880
rect 814 -876 815 -874
rect 814 -882 815 -880
rect 821 -876 822 -874
rect 821 -882 822 -880
rect 828 -876 829 -874
rect 831 -876 832 -874
rect 828 -882 829 -880
rect 835 -876 836 -874
rect 835 -882 836 -880
rect 842 -876 843 -874
rect 842 -882 843 -880
rect 849 -876 850 -874
rect 849 -882 850 -880
rect 856 -876 857 -874
rect 856 -882 857 -880
rect 863 -876 864 -874
rect 863 -882 864 -880
rect 870 -876 871 -874
rect 870 -882 871 -880
rect 877 -876 878 -874
rect 877 -882 878 -880
rect 880 -882 881 -880
rect 884 -876 885 -874
rect 884 -882 885 -880
rect 891 -876 892 -874
rect 891 -882 892 -880
rect 898 -876 899 -874
rect 898 -882 899 -880
rect 905 -876 906 -874
rect 908 -876 909 -874
rect 905 -882 906 -880
rect 908 -882 909 -880
rect 912 -876 913 -874
rect 912 -882 913 -880
rect 919 -876 920 -874
rect 919 -882 920 -880
rect 929 -876 930 -874
rect 926 -882 927 -880
rect 929 -882 930 -880
rect 933 -876 934 -874
rect 933 -882 934 -880
rect 940 -876 941 -874
rect 940 -882 941 -880
rect 947 -876 948 -874
rect 947 -882 948 -880
rect 954 -876 955 -874
rect 954 -882 955 -880
rect 961 -882 962 -880
rect 964 -882 965 -880
rect 968 -876 969 -874
rect 968 -882 969 -880
rect 975 -876 976 -874
rect 975 -882 976 -880
rect 982 -876 983 -874
rect 982 -882 983 -880
rect 989 -876 990 -874
rect 989 -882 990 -880
rect 996 -876 997 -874
rect 996 -882 997 -880
rect 1003 -876 1004 -874
rect 1003 -882 1004 -880
rect 1010 -876 1011 -874
rect 1010 -882 1011 -880
rect 1017 -876 1018 -874
rect 1017 -882 1018 -880
rect 1024 -876 1025 -874
rect 1024 -882 1025 -880
rect 1031 -876 1032 -874
rect 1031 -882 1032 -880
rect 1038 -876 1039 -874
rect 1038 -882 1039 -880
rect 1045 -876 1046 -874
rect 1045 -882 1046 -880
rect 1052 -876 1053 -874
rect 1052 -882 1053 -880
rect 1059 -876 1060 -874
rect 1059 -882 1060 -880
rect 1062 -882 1063 -880
rect 1066 -876 1067 -874
rect 1066 -882 1067 -880
rect 1073 -876 1074 -874
rect 1073 -882 1074 -880
rect 1080 -876 1081 -874
rect 1080 -882 1081 -880
rect 1087 -876 1088 -874
rect 1087 -882 1088 -880
rect 1094 -876 1095 -874
rect 1094 -882 1095 -880
rect 1101 -876 1102 -874
rect 1101 -882 1102 -880
rect 1108 -876 1109 -874
rect 1108 -882 1109 -880
rect 1115 -876 1116 -874
rect 1115 -882 1116 -880
rect 1122 -876 1123 -874
rect 1122 -882 1123 -880
rect 1129 -876 1130 -874
rect 1129 -882 1130 -880
rect 1136 -876 1137 -874
rect 1136 -882 1137 -880
rect 1143 -876 1144 -874
rect 1143 -882 1144 -880
rect 1150 -876 1151 -874
rect 1150 -882 1151 -880
rect 1157 -876 1158 -874
rect 1157 -882 1158 -880
rect 1164 -876 1165 -874
rect 1164 -882 1165 -880
rect 1171 -876 1172 -874
rect 1171 -882 1172 -880
rect 1178 -876 1179 -874
rect 1178 -882 1179 -880
rect 1185 -876 1186 -874
rect 1185 -882 1186 -880
rect 1192 -876 1193 -874
rect 1192 -882 1193 -880
rect 1199 -876 1200 -874
rect 1199 -882 1200 -880
rect 1206 -876 1207 -874
rect 1206 -882 1207 -880
rect 1213 -876 1214 -874
rect 1213 -882 1214 -880
rect 1220 -876 1221 -874
rect 1220 -882 1221 -880
rect 1227 -876 1228 -874
rect 1227 -882 1228 -880
rect 1234 -876 1235 -874
rect 1234 -882 1235 -880
rect 1241 -876 1242 -874
rect 1241 -882 1242 -880
rect 1248 -876 1249 -874
rect 1248 -882 1249 -880
rect 1255 -876 1256 -874
rect 1255 -882 1256 -880
rect 1262 -876 1263 -874
rect 1262 -882 1263 -880
rect 1269 -876 1270 -874
rect 1269 -882 1270 -880
rect 1276 -876 1277 -874
rect 1276 -882 1277 -880
rect 1283 -876 1284 -874
rect 1283 -882 1284 -880
rect 1290 -876 1291 -874
rect 1290 -882 1291 -880
rect 1297 -876 1298 -874
rect 1297 -882 1298 -880
rect 1304 -876 1305 -874
rect 1304 -882 1305 -880
rect 1311 -876 1312 -874
rect 1311 -882 1312 -880
rect 1318 -876 1319 -874
rect 1318 -882 1319 -880
rect 1325 -876 1326 -874
rect 1325 -882 1326 -880
rect 1332 -876 1333 -874
rect 1332 -882 1333 -880
rect 1339 -876 1340 -874
rect 1339 -882 1340 -880
rect 1346 -876 1347 -874
rect 1346 -882 1347 -880
rect 1353 -876 1354 -874
rect 1353 -882 1354 -880
rect 1360 -876 1361 -874
rect 1360 -882 1361 -880
rect 1367 -876 1368 -874
rect 1367 -882 1368 -880
rect 1374 -876 1375 -874
rect 1374 -882 1375 -880
rect 1381 -876 1382 -874
rect 1381 -882 1382 -880
rect 1388 -876 1389 -874
rect 1388 -882 1389 -880
rect 1395 -876 1396 -874
rect 1395 -882 1396 -880
rect 1402 -876 1403 -874
rect 1402 -882 1403 -880
rect 1409 -876 1410 -874
rect 1409 -882 1410 -880
rect 1416 -876 1417 -874
rect 1416 -882 1417 -880
rect 1423 -876 1424 -874
rect 1423 -882 1424 -880
rect 1430 -876 1431 -874
rect 1430 -882 1431 -880
rect 1437 -876 1438 -874
rect 1437 -882 1438 -880
rect 1444 -876 1445 -874
rect 1444 -882 1445 -880
rect 1451 -876 1452 -874
rect 1451 -882 1452 -880
rect 1458 -876 1459 -874
rect 1458 -882 1459 -880
rect 1465 -876 1466 -874
rect 1465 -882 1466 -880
rect 1472 -876 1473 -874
rect 1472 -882 1473 -880
rect 1479 -876 1480 -874
rect 1479 -882 1480 -880
rect 1486 -876 1487 -874
rect 1486 -882 1487 -880
rect 1493 -876 1494 -874
rect 1493 -882 1494 -880
rect 1500 -876 1501 -874
rect 1500 -882 1501 -880
rect 1507 -876 1508 -874
rect 1507 -882 1508 -880
rect 1514 -876 1515 -874
rect 1514 -882 1515 -880
rect 1521 -876 1522 -874
rect 1521 -882 1522 -880
rect 1528 -876 1529 -874
rect 1528 -882 1529 -880
rect 1535 -876 1536 -874
rect 1535 -882 1536 -880
rect 1542 -876 1543 -874
rect 1542 -882 1543 -880
rect 1549 -876 1550 -874
rect 1549 -882 1550 -880
rect 1556 -876 1557 -874
rect 1556 -882 1557 -880
rect 1563 -876 1564 -874
rect 1563 -882 1564 -880
rect 1570 -876 1571 -874
rect 1570 -882 1571 -880
rect 1577 -876 1578 -874
rect 1577 -882 1578 -880
rect 1584 -876 1585 -874
rect 1584 -882 1585 -880
rect 1591 -876 1592 -874
rect 1591 -882 1592 -880
rect 1601 -882 1602 -880
rect 1605 -876 1606 -874
rect 1608 -876 1609 -874
rect 1608 -882 1609 -880
rect 1612 -876 1613 -874
rect 1612 -882 1613 -880
rect 1619 -876 1620 -874
rect 1619 -882 1620 -880
rect 1626 -876 1627 -874
rect 1626 -882 1627 -880
rect 1633 -876 1634 -874
rect 1633 -882 1634 -880
rect 1696 -876 1697 -874
rect 1696 -882 1697 -880
rect 30 -1037 31 -1035
rect 30 -1043 31 -1041
rect 37 -1037 38 -1035
rect 37 -1043 38 -1041
rect 44 -1037 45 -1035
rect 47 -1043 48 -1041
rect 54 -1037 55 -1035
rect 51 -1043 52 -1041
rect 54 -1043 55 -1041
rect 58 -1037 59 -1035
rect 58 -1043 59 -1041
rect 65 -1037 66 -1035
rect 65 -1043 66 -1041
rect 72 -1037 73 -1035
rect 72 -1043 73 -1041
rect 79 -1037 80 -1035
rect 79 -1043 80 -1041
rect 86 -1037 87 -1035
rect 89 -1037 90 -1035
rect 86 -1043 87 -1041
rect 89 -1043 90 -1041
rect 93 -1037 94 -1035
rect 93 -1043 94 -1041
rect 100 -1037 101 -1035
rect 100 -1043 101 -1041
rect 107 -1037 108 -1035
rect 110 -1037 111 -1035
rect 107 -1043 108 -1041
rect 110 -1043 111 -1041
rect 114 -1037 115 -1035
rect 114 -1043 115 -1041
rect 121 -1037 122 -1035
rect 124 -1037 125 -1035
rect 121 -1043 122 -1041
rect 128 -1037 129 -1035
rect 128 -1043 129 -1041
rect 135 -1037 136 -1035
rect 135 -1043 136 -1041
rect 142 -1037 143 -1035
rect 142 -1043 143 -1041
rect 149 -1037 150 -1035
rect 149 -1043 150 -1041
rect 156 -1037 157 -1035
rect 156 -1043 157 -1041
rect 163 -1037 164 -1035
rect 163 -1043 164 -1041
rect 170 -1037 171 -1035
rect 170 -1043 171 -1041
rect 177 -1037 178 -1035
rect 177 -1043 178 -1041
rect 184 -1037 185 -1035
rect 184 -1043 185 -1041
rect 191 -1037 192 -1035
rect 191 -1043 192 -1041
rect 198 -1037 199 -1035
rect 201 -1037 202 -1035
rect 198 -1043 199 -1041
rect 201 -1043 202 -1041
rect 205 -1037 206 -1035
rect 205 -1043 206 -1041
rect 212 -1037 213 -1035
rect 212 -1043 213 -1041
rect 226 -1037 227 -1035
rect 226 -1043 227 -1041
rect 233 -1037 234 -1035
rect 233 -1043 234 -1041
rect 240 -1037 241 -1035
rect 240 -1043 241 -1041
rect 247 -1037 248 -1035
rect 247 -1043 248 -1041
rect 254 -1037 255 -1035
rect 254 -1043 255 -1041
rect 261 -1037 262 -1035
rect 261 -1043 262 -1041
rect 268 -1037 269 -1035
rect 268 -1043 269 -1041
rect 275 -1037 276 -1035
rect 275 -1043 276 -1041
rect 282 -1037 283 -1035
rect 282 -1043 283 -1041
rect 289 -1037 290 -1035
rect 292 -1037 293 -1035
rect 289 -1043 290 -1041
rect 292 -1043 293 -1041
rect 296 -1037 297 -1035
rect 296 -1043 297 -1041
rect 303 -1037 304 -1035
rect 303 -1043 304 -1041
rect 313 -1037 314 -1035
rect 317 -1037 318 -1035
rect 317 -1043 318 -1041
rect 324 -1037 325 -1035
rect 324 -1043 325 -1041
rect 331 -1037 332 -1035
rect 331 -1043 332 -1041
rect 338 -1037 339 -1035
rect 338 -1043 339 -1041
rect 345 -1037 346 -1035
rect 345 -1043 346 -1041
rect 352 -1037 353 -1035
rect 352 -1043 353 -1041
rect 359 -1037 360 -1035
rect 359 -1043 360 -1041
rect 366 -1037 367 -1035
rect 366 -1043 367 -1041
rect 373 -1037 374 -1035
rect 373 -1043 374 -1041
rect 380 -1037 381 -1035
rect 380 -1043 381 -1041
rect 387 -1037 388 -1035
rect 387 -1043 388 -1041
rect 394 -1037 395 -1035
rect 394 -1043 395 -1041
rect 401 -1037 402 -1035
rect 401 -1043 402 -1041
rect 408 -1037 409 -1035
rect 408 -1043 409 -1041
rect 415 -1037 416 -1035
rect 415 -1043 416 -1041
rect 422 -1037 423 -1035
rect 422 -1043 423 -1041
rect 429 -1037 430 -1035
rect 429 -1043 430 -1041
rect 436 -1037 437 -1035
rect 436 -1043 437 -1041
rect 443 -1037 444 -1035
rect 443 -1043 444 -1041
rect 450 -1037 451 -1035
rect 450 -1043 451 -1041
rect 457 -1037 458 -1035
rect 457 -1043 458 -1041
rect 467 -1037 468 -1035
rect 467 -1043 468 -1041
rect 471 -1037 472 -1035
rect 474 -1037 475 -1035
rect 471 -1043 472 -1041
rect 474 -1043 475 -1041
rect 478 -1037 479 -1035
rect 478 -1043 479 -1041
rect 485 -1037 486 -1035
rect 485 -1043 486 -1041
rect 492 -1037 493 -1035
rect 492 -1043 493 -1041
rect 499 -1037 500 -1035
rect 499 -1043 500 -1041
rect 506 -1037 507 -1035
rect 506 -1043 507 -1041
rect 513 -1037 514 -1035
rect 513 -1043 514 -1041
rect 520 -1037 521 -1035
rect 520 -1043 521 -1041
rect 527 -1037 528 -1035
rect 527 -1043 528 -1041
rect 534 -1037 535 -1035
rect 537 -1037 538 -1035
rect 534 -1043 535 -1041
rect 537 -1043 538 -1041
rect 541 -1037 542 -1035
rect 541 -1043 542 -1041
rect 548 -1037 549 -1035
rect 551 -1037 552 -1035
rect 548 -1043 549 -1041
rect 551 -1043 552 -1041
rect 555 -1037 556 -1035
rect 555 -1043 556 -1041
rect 562 -1037 563 -1035
rect 562 -1043 563 -1041
rect 569 -1037 570 -1035
rect 569 -1043 570 -1041
rect 576 -1037 577 -1035
rect 576 -1043 577 -1041
rect 583 -1037 584 -1035
rect 583 -1043 584 -1041
rect 593 -1037 594 -1035
rect 590 -1043 591 -1041
rect 593 -1043 594 -1041
rect 597 -1037 598 -1035
rect 600 -1037 601 -1035
rect 597 -1043 598 -1041
rect 600 -1043 601 -1041
rect 604 -1037 605 -1035
rect 607 -1037 608 -1035
rect 604 -1043 605 -1041
rect 607 -1043 608 -1041
rect 611 -1037 612 -1035
rect 611 -1043 612 -1041
rect 618 -1037 619 -1035
rect 621 -1037 622 -1035
rect 621 -1043 622 -1041
rect 625 -1037 626 -1035
rect 625 -1043 626 -1041
rect 628 -1043 629 -1041
rect 632 -1037 633 -1035
rect 635 -1037 636 -1035
rect 632 -1043 633 -1041
rect 635 -1043 636 -1041
rect 639 -1037 640 -1035
rect 639 -1043 640 -1041
rect 646 -1037 647 -1035
rect 646 -1043 647 -1041
rect 653 -1037 654 -1035
rect 653 -1043 654 -1041
rect 660 -1037 661 -1035
rect 660 -1043 661 -1041
rect 667 -1037 668 -1035
rect 667 -1043 668 -1041
rect 674 -1037 675 -1035
rect 674 -1043 675 -1041
rect 681 -1037 682 -1035
rect 681 -1043 682 -1041
rect 688 -1037 689 -1035
rect 688 -1043 689 -1041
rect 695 -1037 696 -1035
rect 695 -1043 696 -1041
rect 702 -1037 703 -1035
rect 702 -1043 703 -1041
rect 709 -1037 710 -1035
rect 709 -1043 710 -1041
rect 716 -1037 717 -1035
rect 716 -1043 717 -1041
rect 723 -1037 724 -1035
rect 723 -1043 724 -1041
rect 726 -1043 727 -1041
rect 730 -1037 731 -1035
rect 733 -1037 734 -1035
rect 730 -1043 731 -1041
rect 733 -1043 734 -1041
rect 737 -1037 738 -1035
rect 737 -1043 738 -1041
rect 744 -1037 745 -1035
rect 744 -1043 745 -1041
rect 751 -1037 752 -1035
rect 751 -1043 752 -1041
rect 761 -1037 762 -1035
rect 758 -1043 759 -1041
rect 761 -1043 762 -1041
rect 765 -1037 766 -1035
rect 768 -1037 769 -1035
rect 765 -1043 766 -1041
rect 768 -1043 769 -1041
rect 772 -1037 773 -1035
rect 772 -1043 773 -1041
rect 779 -1037 780 -1035
rect 779 -1043 780 -1041
rect 786 -1037 787 -1035
rect 786 -1043 787 -1041
rect 793 -1037 794 -1035
rect 796 -1037 797 -1035
rect 793 -1043 794 -1041
rect 800 -1037 801 -1035
rect 800 -1043 801 -1041
rect 807 -1037 808 -1035
rect 810 -1037 811 -1035
rect 807 -1043 808 -1041
rect 810 -1043 811 -1041
rect 814 -1037 815 -1035
rect 814 -1043 815 -1041
rect 821 -1037 822 -1035
rect 821 -1043 822 -1041
rect 828 -1037 829 -1035
rect 831 -1043 832 -1041
rect 835 -1037 836 -1035
rect 835 -1043 836 -1041
rect 842 -1037 843 -1035
rect 845 -1037 846 -1035
rect 842 -1043 843 -1041
rect 845 -1043 846 -1041
rect 849 -1037 850 -1035
rect 849 -1043 850 -1041
rect 856 -1037 857 -1035
rect 856 -1043 857 -1041
rect 859 -1043 860 -1041
rect 863 -1037 864 -1035
rect 863 -1043 864 -1041
rect 870 -1037 871 -1035
rect 873 -1037 874 -1035
rect 870 -1043 871 -1041
rect 873 -1043 874 -1041
rect 877 -1037 878 -1035
rect 880 -1037 881 -1035
rect 877 -1043 878 -1041
rect 880 -1043 881 -1041
rect 884 -1037 885 -1035
rect 884 -1043 885 -1041
rect 891 -1037 892 -1035
rect 891 -1043 892 -1041
rect 898 -1037 899 -1035
rect 901 -1037 902 -1035
rect 898 -1043 899 -1041
rect 905 -1037 906 -1035
rect 905 -1043 906 -1041
rect 912 -1037 913 -1035
rect 912 -1043 913 -1041
rect 919 -1037 920 -1035
rect 919 -1043 920 -1041
rect 926 -1037 927 -1035
rect 926 -1043 927 -1041
rect 933 -1037 934 -1035
rect 933 -1043 934 -1041
rect 940 -1037 941 -1035
rect 940 -1043 941 -1041
rect 947 -1037 948 -1035
rect 947 -1043 948 -1041
rect 954 -1037 955 -1035
rect 957 -1037 958 -1035
rect 954 -1043 955 -1041
rect 957 -1043 958 -1041
rect 961 -1037 962 -1035
rect 961 -1043 962 -1041
rect 968 -1037 969 -1035
rect 968 -1043 969 -1041
rect 975 -1037 976 -1035
rect 978 -1037 979 -1035
rect 978 -1043 979 -1041
rect 982 -1037 983 -1035
rect 982 -1043 983 -1041
rect 989 -1037 990 -1035
rect 992 -1037 993 -1035
rect 989 -1043 990 -1041
rect 992 -1043 993 -1041
rect 996 -1037 997 -1035
rect 996 -1043 997 -1041
rect 1003 -1037 1004 -1035
rect 1003 -1043 1004 -1041
rect 1010 -1037 1011 -1035
rect 1010 -1043 1011 -1041
rect 1017 -1037 1018 -1035
rect 1017 -1043 1018 -1041
rect 1024 -1037 1025 -1035
rect 1024 -1043 1025 -1041
rect 1031 -1037 1032 -1035
rect 1031 -1043 1032 -1041
rect 1038 -1037 1039 -1035
rect 1038 -1043 1039 -1041
rect 1045 -1037 1046 -1035
rect 1045 -1043 1046 -1041
rect 1052 -1037 1053 -1035
rect 1052 -1043 1053 -1041
rect 1062 -1037 1063 -1035
rect 1062 -1043 1063 -1041
rect 1066 -1037 1067 -1035
rect 1066 -1043 1067 -1041
rect 1069 -1043 1070 -1041
rect 1073 -1037 1074 -1035
rect 1073 -1043 1074 -1041
rect 1080 -1037 1081 -1035
rect 1080 -1043 1081 -1041
rect 1087 -1037 1088 -1035
rect 1087 -1043 1088 -1041
rect 1094 -1037 1095 -1035
rect 1094 -1043 1095 -1041
rect 1101 -1037 1102 -1035
rect 1101 -1043 1102 -1041
rect 1108 -1037 1109 -1035
rect 1108 -1043 1109 -1041
rect 1115 -1037 1116 -1035
rect 1115 -1043 1116 -1041
rect 1122 -1037 1123 -1035
rect 1122 -1043 1123 -1041
rect 1129 -1037 1130 -1035
rect 1129 -1043 1130 -1041
rect 1136 -1037 1137 -1035
rect 1136 -1043 1137 -1041
rect 1143 -1037 1144 -1035
rect 1143 -1043 1144 -1041
rect 1150 -1037 1151 -1035
rect 1150 -1043 1151 -1041
rect 1157 -1037 1158 -1035
rect 1157 -1043 1158 -1041
rect 1164 -1037 1165 -1035
rect 1164 -1043 1165 -1041
rect 1171 -1037 1172 -1035
rect 1171 -1043 1172 -1041
rect 1178 -1037 1179 -1035
rect 1178 -1043 1179 -1041
rect 1185 -1037 1186 -1035
rect 1185 -1043 1186 -1041
rect 1192 -1037 1193 -1035
rect 1192 -1043 1193 -1041
rect 1199 -1037 1200 -1035
rect 1199 -1043 1200 -1041
rect 1206 -1037 1207 -1035
rect 1206 -1043 1207 -1041
rect 1213 -1037 1214 -1035
rect 1213 -1043 1214 -1041
rect 1220 -1037 1221 -1035
rect 1220 -1043 1221 -1041
rect 1227 -1037 1228 -1035
rect 1227 -1043 1228 -1041
rect 1234 -1037 1235 -1035
rect 1234 -1043 1235 -1041
rect 1241 -1037 1242 -1035
rect 1241 -1043 1242 -1041
rect 1248 -1037 1249 -1035
rect 1248 -1043 1249 -1041
rect 1255 -1037 1256 -1035
rect 1255 -1043 1256 -1041
rect 1262 -1037 1263 -1035
rect 1262 -1043 1263 -1041
rect 1269 -1037 1270 -1035
rect 1269 -1043 1270 -1041
rect 1276 -1037 1277 -1035
rect 1276 -1043 1277 -1041
rect 1283 -1037 1284 -1035
rect 1283 -1043 1284 -1041
rect 1290 -1037 1291 -1035
rect 1290 -1043 1291 -1041
rect 1297 -1037 1298 -1035
rect 1297 -1043 1298 -1041
rect 1304 -1037 1305 -1035
rect 1304 -1043 1305 -1041
rect 1311 -1037 1312 -1035
rect 1311 -1043 1312 -1041
rect 1318 -1037 1319 -1035
rect 1318 -1043 1319 -1041
rect 1325 -1037 1326 -1035
rect 1325 -1043 1326 -1041
rect 1332 -1037 1333 -1035
rect 1332 -1043 1333 -1041
rect 1339 -1037 1340 -1035
rect 1339 -1043 1340 -1041
rect 1346 -1037 1347 -1035
rect 1346 -1043 1347 -1041
rect 1353 -1037 1354 -1035
rect 1353 -1043 1354 -1041
rect 1360 -1037 1361 -1035
rect 1360 -1043 1361 -1041
rect 1367 -1037 1368 -1035
rect 1367 -1043 1368 -1041
rect 1374 -1037 1375 -1035
rect 1374 -1043 1375 -1041
rect 1381 -1037 1382 -1035
rect 1381 -1043 1382 -1041
rect 1388 -1037 1389 -1035
rect 1388 -1043 1389 -1041
rect 1395 -1037 1396 -1035
rect 1395 -1043 1396 -1041
rect 1402 -1037 1403 -1035
rect 1402 -1043 1403 -1041
rect 1409 -1037 1410 -1035
rect 1409 -1043 1410 -1041
rect 1416 -1037 1417 -1035
rect 1416 -1043 1417 -1041
rect 1423 -1037 1424 -1035
rect 1423 -1043 1424 -1041
rect 1430 -1037 1431 -1035
rect 1430 -1043 1431 -1041
rect 1437 -1037 1438 -1035
rect 1437 -1043 1438 -1041
rect 1444 -1037 1445 -1035
rect 1444 -1043 1445 -1041
rect 1451 -1037 1452 -1035
rect 1451 -1043 1452 -1041
rect 1458 -1037 1459 -1035
rect 1458 -1043 1459 -1041
rect 1465 -1037 1466 -1035
rect 1465 -1043 1466 -1041
rect 1472 -1037 1473 -1035
rect 1472 -1043 1473 -1041
rect 1479 -1037 1480 -1035
rect 1479 -1043 1480 -1041
rect 1486 -1037 1487 -1035
rect 1486 -1043 1487 -1041
rect 1493 -1037 1494 -1035
rect 1493 -1043 1494 -1041
rect 1500 -1037 1501 -1035
rect 1500 -1043 1501 -1041
rect 1507 -1037 1508 -1035
rect 1507 -1043 1508 -1041
rect 1514 -1037 1515 -1035
rect 1514 -1043 1515 -1041
rect 1521 -1037 1522 -1035
rect 1521 -1043 1522 -1041
rect 1528 -1037 1529 -1035
rect 1528 -1043 1529 -1041
rect 1535 -1037 1536 -1035
rect 1535 -1043 1536 -1041
rect 1542 -1037 1543 -1035
rect 1542 -1043 1543 -1041
rect 1549 -1037 1550 -1035
rect 1549 -1043 1550 -1041
rect 1556 -1037 1557 -1035
rect 1556 -1043 1557 -1041
rect 1563 -1037 1564 -1035
rect 1563 -1043 1564 -1041
rect 1570 -1037 1571 -1035
rect 1570 -1043 1571 -1041
rect 1577 -1037 1578 -1035
rect 1577 -1043 1578 -1041
rect 1584 -1037 1585 -1035
rect 1584 -1043 1585 -1041
rect 1591 -1037 1592 -1035
rect 1591 -1043 1592 -1041
rect 1598 -1037 1599 -1035
rect 1598 -1043 1599 -1041
rect 1605 -1037 1606 -1035
rect 1605 -1043 1606 -1041
rect 1612 -1037 1613 -1035
rect 1612 -1043 1613 -1041
rect 1619 -1037 1620 -1035
rect 1619 -1043 1620 -1041
rect 1626 -1037 1627 -1035
rect 1626 -1043 1627 -1041
rect 1633 -1037 1634 -1035
rect 1633 -1043 1634 -1041
rect 1640 -1037 1641 -1035
rect 1640 -1043 1641 -1041
rect 1647 -1037 1648 -1035
rect 1647 -1043 1648 -1041
rect 1654 -1037 1655 -1035
rect 1654 -1043 1655 -1041
rect 1661 -1037 1662 -1035
rect 1661 -1043 1662 -1041
rect 1668 -1037 1669 -1035
rect 1668 -1043 1669 -1041
rect 1675 -1037 1676 -1035
rect 1675 -1043 1676 -1041
rect 1682 -1037 1683 -1035
rect 1682 -1043 1683 -1041
rect 1689 -1037 1690 -1035
rect 1689 -1043 1690 -1041
rect 1696 -1037 1697 -1035
rect 1696 -1043 1697 -1041
rect 1703 -1037 1704 -1035
rect 1703 -1043 1704 -1041
rect 1710 -1037 1711 -1035
rect 1710 -1043 1711 -1041
rect 1717 -1037 1718 -1035
rect 1717 -1043 1718 -1041
rect 1724 -1037 1725 -1035
rect 1724 -1043 1725 -1041
rect 30 -1188 31 -1186
rect 30 -1194 31 -1192
rect 37 -1188 38 -1186
rect 37 -1194 38 -1192
rect 44 -1188 45 -1186
rect 44 -1194 45 -1192
rect 51 -1188 52 -1186
rect 51 -1194 52 -1192
rect 58 -1188 59 -1186
rect 58 -1194 59 -1192
rect 65 -1188 66 -1186
rect 65 -1194 66 -1192
rect 75 -1188 76 -1186
rect 75 -1194 76 -1192
rect 79 -1188 80 -1186
rect 82 -1194 83 -1192
rect 89 -1188 90 -1186
rect 86 -1194 87 -1192
rect 89 -1194 90 -1192
rect 93 -1188 94 -1186
rect 93 -1194 94 -1192
rect 100 -1188 101 -1186
rect 103 -1188 104 -1186
rect 107 -1188 108 -1186
rect 107 -1194 108 -1192
rect 114 -1188 115 -1186
rect 114 -1194 115 -1192
rect 121 -1188 122 -1186
rect 124 -1188 125 -1186
rect 121 -1194 122 -1192
rect 124 -1194 125 -1192
rect 128 -1188 129 -1186
rect 128 -1194 129 -1192
rect 135 -1188 136 -1186
rect 135 -1194 136 -1192
rect 142 -1188 143 -1186
rect 142 -1194 143 -1192
rect 149 -1188 150 -1186
rect 149 -1194 150 -1192
rect 152 -1194 153 -1192
rect 156 -1188 157 -1186
rect 156 -1194 157 -1192
rect 163 -1188 164 -1186
rect 166 -1188 167 -1186
rect 163 -1194 164 -1192
rect 166 -1194 167 -1192
rect 170 -1188 171 -1186
rect 170 -1194 171 -1192
rect 177 -1188 178 -1186
rect 177 -1194 178 -1192
rect 184 -1188 185 -1186
rect 187 -1188 188 -1186
rect 184 -1194 185 -1192
rect 191 -1188 192 -1186
rect 191 -1194 192 -1192
rect 198 -1188 199 -1186
rect 201 -1188 202 -1186
rect 198 -1194 199 -1192
rect 201 -1194 202 -1192
rect 205 -1188 206 -1186
rect 208 -1188 209 -1186
rect 205 -1194 206 -1192
rect 208 -1194 209 -1192
rect 212 -1188 213 -1186
rect 212 -1194 213 -1192
rect 219 -1188 220 -1186
rect 219 -1194 220 -1192
rect 226 -1188 227 -1186
rect 226 -1194 227 -1192
rect 236 -1188 237 -1186
rect 233 -1194 234 -1192
rect 236 -1194 237 -1192
rect 240 -1188 241 -1186
rect 240 -1194 241 -1192
rect 247 -1188 248 -1186
rect 247 -1194 248 -1192
rect 254 -1188 255 -1186
rect 257 -1194 258 -1192
rect 261 -1188 262 -1186
rect 261 -1194 262 -1192
rect 268 -1188 269 -1186
rect 268 -1194 269 -1192
rect 275 -1188 276 -1186
rect 278 -1194 279 -1192
rect 282 -1188 283 -1186
rect 282 -1194 283 -1192
rect 289 -1188 290 -1186
rect 289 -1194 290 -1192
rect 296 -1188 297 -1186
rect 296 -1194 297 -1192
rect 303 -1188 304 -1186
rect 303 -1194 304 -1192
rect 310 -1188 311 -1186
rect 310 -1194 311 -1192
rect 317 -1188 318 -1186
rect 317 -1194 318 -1192
rect 324 -1188 325 -1186
rect 324 -1194 325 -1192
rect 331 -1188 332 -1186
rect 331 -1194 332 -1192
rect 338 -1188 339 -1186
rect 338 -1194 339 -1192
rect 345 -1188 346 -1186
rect 345 -1194 346 -1192
rect 352 -1188 353 -1186
rect 352 -1194 353 -1192
rect 359 -1188 360 -1186
rect 359 -1194 360 -1192
rect 366 -1188 367 -1186
rect 366 -1194 367 -1192
rect 373 -1188 374 -1186
rect 373 -1194 374 -1192
rect 380 -1188 381 -1186
rect 380 -1194 381 -1192
rect 387 -1188 388 -1186
rect 387 -1194 388 -1192
rect 394 -1188 395 -1186
rect 394 -1194 395 -1192
rect 401 -1188 402 -1186
rect 401 -1194 402 -1192
rect 408 -1188 409 -1186
rect 408 -1194 409 -1192
rect 415 -1188 416 -1186
rect 415 -1194 416 -1192
rect 422 -1188 423 -1186
rect 422 -1194 423 -1192
rect 429 -1188 430 -1186
rect 429 -1194 430 -1192
rect 436 -1188 437 -1186
rect 436 -1194 437 -1192
rect 443 -1188 444 -1186
rect 443 -1194 444 -1192
rect 450 -1188 451 -1186
rect 450 -1194 451 -1192
rect 457 -1188 458 -1186
rect 457 -1194 458 -1192
rect 464 -1188 465 -1186
rect 467 -1188 468 -1186
rect 464 -1194 465 -1192
rect 467 -1194 468 -1192
rect 471 -1188 472 -1186
rect 471 -1194 472 -1192
rect 478 -1188 479 -1186
rect 478 -1194 479 -1192
rect 485 -1188 486 -1186
rect 488 -1188 489 -1186
rect 488 -1194 489 -1192
rect 492 -1188 493 -1186
rect 492 -1194 493 -1192
rect 499 -1188 500 -1186
rect 499 -1194 500 -1192
rect 506 -1188 507 -1186
rect 509 -1194 510 -1192
rect 513 -1188 514 -1186
rect 516 -1188 517 -1186
rect 513 -1194 514 -1192
rect 516 -1194 517 -1192
rect 520 -1188 521 -1186
rect 527 -1188 528 -1186
rect 527 -1194 528 -1192
rect 534 -1188 535 -1186
rect 534 -1194 535 -1192
rect 541 -1188 542 -1186
rect 544 -1188 545 -1186
rect 544 -1194 545 -1192
rect 548 -1188 549 -1186
rect 548 -1194 549 -1192
rect 555 -1188 556 -1186
rect 555 -1194 556 -1192
rect 562 -1188 563 -1186
rect 562 -1194 563 -1192
rect 569 -1188 570 -1186
rect 569 -1194 570 -1192
rect 579 -1188 580 -1186
rect 576 -1194 577 -1192
rect 583 -1188 584 -1186
rect 583 -1194 584 -1192
rect 590 -1188 591 -1186
rect 590 -1194 591 -1192
rect 597 -1188 598 -1186
rect 600 -1188 601 -1186
rect 597 -1194 598 -1192
rect 604 -1188 605 -1186
rect 604 -1194 605 -1192
rect 611 -1188 612 -1186
rect 614 -1188 615 -1186
rect 611 -1194 612 -1192
rect 614 -1194 615 -1192
rect 621 -1188 622 -1186
rect 618 -1194 619 -1192
rect 621 -1194 622 -1192
rect 625 -1188 626 -1186
rect 625 -1194 626 -1192
rect 632 -1188 633 -1186
rect 632 -1194 633 -1192
rect 639 -1188 640 -1186
rect 639 -1194 640 -1192
rect 646 -1188 647 -1186
rect 646 -1194 647 -1192
rect 653 -1188 654 -1186
rect 653 -1194 654 -1192
rect 660 -1188 661 -1186
rect 663 -1188 664 -1186
rect 660 -1194 661 -1192
rect 663 -1194 664 -1192
rect 667 -1188 668 -1186
rect 667 -1194 668 -1192
rect 674 -1188 675 -1186
rect 674 -1194 675 -1192
rect 681 -1188 682 -1186
rect 681 -1194 682 -1192
rect 688 -1188 689 -1186
rect 688 -1194 689 -1192
rect 695 -1188 696 -1186
rect 695 -1194 696 -1192
rect 702 -1188 703 -1186
rect 702 -1194 703 -1192
rect 709 -1188 710 -1186
rect 709 -1194 710 -1192
rect 716 -1188 717 -1186
rect 719 -1188 720 -1186
rect 719 -1194 720 -1192
rect 723 -1188 724 -1186
rect 726 -1188 727 -1186
rect 723 -1194 724 -1192
rect 726 -1194 727 -1192
rect 730 -1188 731 -1186
rect 730 -1194 731 -1192
rect 737 -1188 738 -1186
rect 737 -1194 738 -1192
rect 744 -1188 745 -1186
rect 747 -1188 748 -1186
rect 744 -1194 745 -1192
rect 747 -1194 748 -1192
rect 751 -1188 752 -1186
rect 754 -1188 755 -1186
rect 751 -1194 752 -1192
rect 758 -1188 759 -1186
rect 758 -1194 759 -1192
rect 765 -1188 766 -1186
rect 765 -1194 766 -1192
rect 772 -1188 773 -1186
rect 772 -1194 773 -1192
rect 779 -1188 780 -1186
rect 779 -1194 780 -1192
rect 786 -1188 787 -1186
rect 786 -1194 787 -1192
rect 793 -1188 794 -1186
rect 793 -1194 794 -1192
rect 800 -1188 801 -1186
rect 800 -1194 801 -1192
rect 807 -1188 808 -1186
rect 807 -1194 808 -1192
rect 814 -1188 815 -1186
rect 814 -1194 815 -1192
rect 821 -1188 822 -1186
rect 821 -1194 822 -1192
rect 828 -1188 829 -1186
rect 828 -1194 829 -1192
rect 831 -1194 832 -1192
rect 835 -1188 836 -1186
rect 835 -1194 836 -1192
rect 842 -1188 843 -1186
rect 842 -1194 843 -1192
rect 849 -1188 850 -1186
rect 849 -1194 850 -1192
rect 856 -1188 857 -1186
rect 856 -1194 857 -1192
rect 863 -1188 864 -1186
rect 863 -1194 864 -1192
rect 870 -1188 871 -1186
rect 870 -1194 871 -1192
rect 873 -1194 874 -1192
rect 877 -1188 878 -1186
rect 877 -1194 878 -1192
rect 884 -1188 885 -1186
rect 884 -1194 885 -1192
rect 894 -1188 895 -1186
rect 891 -1194 892 -1192
rect 894 -1194 895 -1192
rect 898 -1188 899 -1186
rect 901 -1188 902 -1186
rect 898 -1194 899 -1192
rect 901 -1194 902 -1192
rect 905 -1188 906 -1186
rect 905 -1194 906 -1192
rect 912 -1188 913 -1186
rect 912 -1194 913 -1192
rect 919 -1188 920 -1186
rect 919 -1194 920 -1192
rect 926 -1188 927 -1186
rect 926 -1194 927 -1192
rect 933 -1188 934 -1186
rect 933 -1194 934 -1192
rect 940 -1188 941 -1186
rect 940 -1194 941 -1192
rect 947 -1188 948 -1186
rect 947 -1194 948 -1192
rect 954 -1188 955 -1186
rect 957 -1188 958 -1186
rect 954 -1194 955 -1192
rect 957 -1194 958 -1192
rect 961 -1188 962 -1186
rect 961 -1194 962 -1192
rect 968 -1188 969 -1186
rect 971 -1188 972 -1186
rect 968 -1194 969 -1192
rect 971 -1194 972 -1192
rect 975 -1188 976 -1186
rect 975 -1194 976 -1192
rect 982 -1188 983 -1186
rect 982 -1194 983 -1192
rect 989 -1188 990 -1186
rect 992 -1188 993 -1186
rect 989 -1194 990 -1192
rect 992 -1194 993 -1192
rect 996 -1188 997 -1186
rect 996 -1194 997 -1192
rect 999 -1194 1000 -1192
rect 1003 -1188 1004 -1186
rect 1003 -1194 1004 -1192
rect 1010 -1188 1011 -1186
rect 1010 -1194 1011 -1192
rect 1017 -1188 1018 -1186
rect 1017 -1194 1018 -1192
rect 1024 -1188 1025 -1186
rect 1024 -1194 1025 -1192
rect 1031 -1188 1032 -1186
rect 1031 -1194 1032 -1192
rect 1038 -1188 1039 -1186
rect 1038 -1194 1039 -1192
rect 1045 -1188 1046 -1186
rect 1048 -1188 1049 -1186
rect 1045 -1194 1046 -1192
rect 1048 -1194 1049 -1192
rect 1052 -1188 1053 -1186
rect 1052 -1194 1053 -1192
rect 1059 -1188 1060 -1186
rect 1059 -1194 1060 -1192
rect 1066 -1188 1067 -1186
rect 1066 -1194 1067 -1192
rect 1073 -1188 1074 -1186
rect 1073 -1194 1074 -1192
rect 1080 -1188 1081 -1186
rect 1080 -1194 1081 -1192
rect 1087 -1188 1088 -1186
rect 1087 -1194 1088 -1192
rect 1094 -1188 1095 -1186
rect 1094 -1194 1095 -1192
rect 1101 -1188 1102 -1186
rect 1101 -1194 1102 -1192
rect 1108 -1188 1109 -1186
rect 1108 -1194 1109 -1192
rect 1115 -1188 1116 -1186
rect 1115 -1194 1116 -1192
rect 1122 -1188 1123 -1186
rect 1122 -1194 1123 -1192
rect 1129 -1188 1130 -1186
rect 1129 -1194 1130 -1192
rect 1136 -1188 1137 -1186
rect 1136 -1194 1137 -1192
rect 1143 -1188 1144 -1186
rect 1143 -1194 1144 -1192
rect 1150 -1188 1151 -1186
rect 1150 -1194 1151 -1192
rect 1157 -1188 1158 -1186
rect 1157 -1194 1158 -1192
rect 1164 -1188 1165 -1186
rect 1164 -1194 1165 -1192
rect 1171 -1188 1172 -1186
rect 1171 -1194 1172 -1192
rect 1178 -1188 1179 -1186
rect 1178 -1194 1179 -1192
rect 1185 -1188 1186 -1186
rect 1185 -1194 1186 -1192
rect 1192 -1188 1193 -1186
rect 1192 -1194 1193 -1192
rect 1199 -1188 1200 -1186
rect 1199 -1194 1200 -1192
rect 1206 -1188 1207 -1186
rect 1206 -1194 1207 -1192
rect 1213 -1188 1214 -1186
rect 1213 -1194 1214 -1192
rect 1220 -1188 1221 -1186
rect 1220 -1194 1221 -1192
rect 1227 -1188 1228 -1186
rect 1227 -1194 1228 -1192
rect 1234 -1188 1235 -1186
rect 1234 -1194 1235 -1192
rect 1241 -1188 1242 -1186
rect 1241 -1194 1242 -1192
rect 1248 -1188 1249 -1186
rect 1248 -1194 1249 -1192
rect 1255 -1188 1256 -1186
rect 1255 -1194 1256 -1192
rect 1262 -1188 1263 -1186
rect 1262 -1194 1263 -1192
rect 1269 -1188 1270 -1186
rect 1269 -1194 1270 -1192
rect 1276 -1188 1277 -1186
rect 1276 -1194 1277 -1192
rect 1283 -1188 1284 -1186
rect 1283 -1194 1284 -1192
rect 1290 -1188 1291 -1186
rect 1290 -1194 1291 -1192
rect 1297 -1188 1298 -1186
rect 1297 -1194 1298 -1192
rect 1304 -1188 1305 -1186
rect 1304 -1194 1305 -1192
rect 1311 -1188 1312 -1186
rect 1311 -1194 1312 -1192
rect 1318 -1188 1319 -1186
rect 1318 -1194 1319 -1192
rect 1325 -1188 1326 -1186
rect 1325 -1194 1326 -1192
rect 1332 -1188 1333 -1186
rect 1332 -1194 1333 -1192
rect 1339 -1188 1340 -1186
rect 1339 -1194 1340 -1192
rect 1346 -1188 1347 -1186
rect 1346 -1194 1347 -1192
rect 1353 -1188 1354 -1186
rect 1353 -1194 1354 -1192
rect 1360 -1188 1361 -1186
rect 1360 -1194 1361 -1192
rect 1367 -1188 1368 -1186
rect 1367 -1194 1368 -1192
rect 1374 -1188 1375 -1186
rect 1374 -1194 1375 -1192
rect 1381 -1188 1382 -1186
rect 1381 -1194 1382 -1192
rect 1388 -1188 1389 -1186
rect 1388 -1194 1389 -1192
rect 1395 -1188 1396 -1186
rect 1395 -1194 1396 -1192
rect 1402 -1188 1403 -1186
rect 1402 -1194 1403 -1192
rect 1409 -1188 1410 -1186
rect 1409 -1194 1410 -1192
rect 1416 -1188 1417 -1186
rect 1416 -1194 1417 -1192
rect 1423 -1188 1424 -1186
rect 1423 -1194 1424 -1192
rect 1430 -1188 1431 -1186
rect 1430 -1194 1431 -1192
rect 1437 -1188 1438 -1186
rect 1437 -1194 1438 -1192
rect 1444 -1188 1445 -1186
rect 1444 -1194 1445 -1192
rect 1451 -1188 1452 -1186
rect 1451 -1194 1452 -1192
rect 1458 -1188 1459 -1186
rect 1458 -1194 1459 -1192
rect 1465 -1188 1466 -1186
rect 1465 -1194 1466 -1192
rect 1472 -1188 1473 -1186
rect 1472 -1194 1473 -1192
rect 1479 -1188 1480 -1186
rect 1479 -1194 1480 -1192
rect 1486 -1188 1487 -1186
rect 1486 -1194 1487 -1192
rect 1493 -1188 1494 -1186
rect 1493 -1194 1494 -1192
rect 1500 -1188 1501 -1186
rect 1500 -1194 1501 -1192
rect 1507 -1188 1508 -1186
rect 1507 -1194 1508 -1192
rect 1514 -1188 1515 -1186
rect 1514 -1194 1515 -1192
rect 1521 -1188 1522 -1186
rect 1521 -1194 1522 -1192
rect 1528 -1188 1529 -1186
rect 1528 -1194 1529 -1192
rect 1535 -1188 1536 -1186
rect 1535 -1194 1536 -1192
rect 1542 -1188 1543 -1186
rect 1542 -1194 1543 -1192
rect 1549 -1188 1550 -1186
rect 1549 -1194 1550 -1192
rect 1556 -1188 1557 -1186
rect 1556 -1194 1557 -1192
rect 1563 -1188 1564 -1186
rect 1563 -1194 1564 -1192
rect 1570 -1188 1571 -1186
rect 1570 -1194 1571 -1192
rect 1577 -1188 1578 -1186
rect 1577 -1194 1578 -1192
rect 1584 -1188 1585 -1186
rect 1584 -1194 1585 -1192
rect 1591 -1188 1592 -1186
rect 1591 -1194 1592 -1192
rect 1598 -1188 1599 -1186
rect 1598 -1194 1599 -1192
rect 1605 -1188 1606 -1186
rect 1605 -1194 1606 -1192
rect 1612 -1188 1613 -1186
rect 1612 -1194 1613 -1192
rect 1619 -1188 1620 -1186
rect 1619 -1194 1620 -1192
rect 1626 -1188 1627 -1186
rect 1626 -1194 1627 -1192
rect 1633 -1188 1634 -1186
rect 1633 -1194 1634 -1192
rect 1640 -1188 1641 -1186
rect 1640 -1194 1641 -1192
rect 1647 -1188 1648 -1186
rect 1650 -1188 1651 -1186
rect 1647 -1194 1648 -1192
rect 1654 -1188 1655 -1186
rect 1654 -1194 1655 -1192
rect 1664 -1188 1665 -1186
rect 1661 -1194 1662 -1192
rect 1664 -1194 1665 -1192
rect 1675 -1188 1676 -1186
rect 1675 -1194 1676 -1192
rect 1724 -1188 1725 -1186
rect 1724 -1194 1725 -1192
rect 1731 -1188 1732 -1186
rect 1731 -1194 1732 -1192
rect 23 -1319 24 -1317
rect 23 -1325 24 -1323
rect 30 -1319 31 -1317
rect 30 -1325 31 -1323
rect 37 -1319 38 -1317
rect 37 -1325 38 -1323
rect 44 -1319 45 -1317
rect 44 -1325 45 -1323
rect 51 -1319 52 -1317
rect 51 -1325 52 -1323
rect 58 -1319 59 -1317
rect 58 -1325 59 -1323
rect 65 -1319 66 -1317
rect 65 -1325 66 -1323
rect 75 -1319 76 -1317
rect 72 -1325 73 -1323
rect 79 -1319 80 -1317
rect 82 -1319 83 -1317
rect 82 -1325 83 -1323
rect 86 -1319 87 -1317
rect 86 -1325 87 -1323
rect 93 -1319 94 -1317
rect 96 -1319 97 -1317
rect 93 -1325 94 -1323
rect 96 -1325 97 -1323
rect 100 -1319 101 -1317
rect 100 -1325 101 -1323
rect 107 -1319 108 -1317
rect 107 -1325 108 -1323
rect 114 -1319 115 -1317
rect 114 -1325 115 -1323
rect 121 -1319 122 -1317
rect 124 -1319 125 -1317
rect 121 -1325 122 -1323
rect 124 -1325 125 -1323
rect 128 -1319 129 -1317
rect 128 -1325 129 -1323
rect 135 -1319 136 -1317
rect 135 -1325 136 -1323
rect 142 -1319 143 -1317
rect 145 -1319 146 -1317
rect 142 -1325 143 -1323
rect 145 -1325 146 -1323
rect 149 -1319 150 -1317
rect 149 -1325 150 -1323
rect 156 -1319 157 -1317
rect 156 -1325 157 -1323
rect 163 -1319 164 -1317
rect 166 -1319 167 -1317
rect 163 -1325 164 -1323
rect 170 -1319 171 -1317
rect 170 -1325 171 -1323
rect 177 -1319 178 -1317
rect 177 -1325 178 -1323
rect 184 -1319 185 -1317
rect 184 -1325 185 -1323
rect 191 -1319 192 -1317
rect 191 -1325 192 -1323
rect 198 -1319 199 -1317
rect 198 -1325 199 -1323
rect 205 -1319 206 -1317
rect 205 -1325 206 -1323
rect 212 -1319 213 -1317
rect 212 -1325 213 -1323
rect 219 -1319 220 -1317
rect 219 -1325 220 -1323
rect 226 -1319 227 -1317
rect 226 -1325 227 -1323
rect 233 -1319 234 -1317
rect 236 -1325 237 -1323
rect 240 -1319 241 -1317
rect 240 -1325 241 -1323
rect 250 -1319 251 -1317
rect 247 -1325 248 -1323
rect 250 -1325 251 -1323
rect 254 -1319 255 -1317
rect 254 -1325 255 -1323
rect 261 -1319 262 -1317
rect 261 -1325 262 -1323
rect 268 -1319 269 -1317
rect 268 -1325 269 -1323
rect 275 -1325 276 -1323
rect 278 -1325 279 -1323
rect 282 -1319 283 -1317
rect 282 -1325 283 -1323
rect 289 -1319 290 -1317
rect 289 -1325 290 -1323
rect 296 -1319 297 -1317
rect 296 -1325 297 -1323
rect 303 -1319 304 -1317
rect 303 -1325 304 -1323
rect 310 -1319 311 -1317
rect 310 -1325 311 -1323
rect 317 -1319 318 -1317
rect 317 -1325 318 -1323
rect 324 -1319 325 -1317
rect 324 -1325 325 -1323
rect 331 -1319 332 -1317
rect 331 -1325 332 -1323
rect 338 -1319 339 -1317
rect 338 -1325 339 -1323
rect 345 -1319 346 -1317
rect 345 -1325 346 -1323
rect 352 -1319 353 -1317
rect 352 -1325 353 -1323
rect 359 -1319 360 -1317
rect 359 -1325 360 -1323
rect 366 -1319 367 -1317
rect 366 -1325 367 -1323
rect 373 -1319 374 -1317
rect 373 -1325 374 -1323
rect 380 -1319 381 -1317
rect 380 -1325 381 -1323
rect 387 -1319 388 -1317
rect 387 -1325 388 -1323
rect 394 -1319 395 -1317
rect 394 -1325 395 -1323
rect 401 -1319 402 -1317
rect 401 -1325 402 -1323
rect 408 -1319 409 -1317
rect 408 -1325 409 -1323
rect 415 -1319 416 -1317
rect 415 -1325 416 -1323
rect 422 -1319 423 -1317
rect 425 -1319 426 -1317
rect 422 -1325 423 -1323
rect 429 -1319 430 -1317
rect 429 -1325 430 -1323
rect 436 -1319 437 -1317
rect 436 -1325 437 -1323
rect 443 -1319 444 -1317
rect 443 -1325 444 -1323
rect 450 -1319 451 -1317
rect 450 -1325 451 -1323
rect 460 -1319 461 -1317
rect 457 -1325 458 -1323
rect 460 -1325 461 -1323
rect 464 -1319 465 -1317
rect 464 -1325 465 -1323
rect 471 -1319 472 -1317
rect 471 -1325 472 -1323
rect 478 -1319 479 -1317
rect 481 -1319 482 -1317
rect 478 -1325 479 -1323
rect 485 -1319 486 -1317
rect 485 -1325 486 -1323
rect 492 -1319 493 -1317
rect 492 -1325 493 -1323
rect 499 -1319 500 -1317
rect 499 -1325 500 -1323
rect 506 -1319 507 -1317
rect 509 -1319 510 -1317
rect 506 -1325 507 -1323
rect 509 -1325 510 -1323
rect 513 -1319 514 -1317
rect 516 -1319 517 -1317
rect 520 -1325 521 -1323
rect 527 -1319 528 -1317
rect 530 -1319 531 -1317
rect 527 -1325 528 -1323
rect 530 -1325 531 -1323
rect 534 -1319 535 -1317
rect 534 -1325 535 -1323
rect 541 -1319 542 -1317
rect 541 -1325 542 -1323
rect 548 -1319 549 -1317
rect 548 -1325 549 -1323
rect 555 -1319 556 -1317
rect 555 -1325 556 -1323
rect 562 -1319 563 -1317
rect 562 -1325 563 -1323
rect 569 -1319 570 -1317
rect 569 -1325 570 -1323
rect 576 -1319 577 -1317
rect 576 -1325 577 -1323
rect 579 -1325 580 -1323
rect 583 -1319 584 -1317
rect 583 -1325 584 -1323
rect 593 -1319 594 -1317
rect 590 -1325 591 -1323
rect 597 -1319 598 -1317
rect 597 -1325 598 -1323
rect 604 -1319 605 -1317
rect 604 -1325 605 -1323
rect 614 -1319 615 -1317
rect 611 -1325 612 -1323
rect 614 -1325 615 -1323
rect 618 -1319 619 -1317
rect 618 -1325 619 -1323
rect 625 -1319 626 -1317
rect 628 -1319 629 -1317
rect 625 -1325 626 -1323
rect 628 -1325 629 -1323
rect 632 -1319 633 -1317
rect 632 -1325 633 -1323
rect 639 -1319 640 -1317
rect 639 -1325 640 -1323
rect 646 -1319 647 -1317
rect 646 -1325 647 -1323
rect 653 -1319 654 -1317
rect 653 -1325 654 -1323
rect 660 -1319 661 -1317
rect 660 -1325 661 -1323
rect 663 -1325 664 -1323
rect 667 -1319 668 -1317
rect 667 -1325 668 -1323
rect 674 -1319 675 -1317
rect 674 -1325 675 -1323
rect 681 -1319 682 -1317
rect 681 -1325 682 -1323
rect 688 -1319 689 -1317
rect 691 -1319 692 -1317
rect 688 -1325 689 -1323
rect 691 -1325 692 -1323
rect 695 -1319 696 -1317
rect 695 -1325 696 -1323
rect 702 -1319 703 -1317
rect 702 -1325 703 -1323
rect 709 -1319 710 -1317
rect 709 -1325 710 -1323
rect 716 -1319 717 -1317
rect 716 -1325 717 -1323
rect 723 -1319 724 -1317
rect 723 -1325 724 -1323
rect 730 -1319 731 -1317
rect 730 -1325 731 -1323
rect 737 -1319 738 -1317
rect 737 -1325 738 -1323
rect 744 -1319 745 -1317
rect 744 -1325 745 -1323
rect 751 -1319 752 -1317
rect 751 -1325 752 -1323
rect 758 -1319 759 -1317
rect 758 -1325 759 -1323
rect 765 -1319 766 -1317
rect 768 -1319 769 -1317
rect 765 -1325 766 -1323
rect 768 -1325 769 -1323
rect 772 -1319 773 -1317
rect 772 -1325 773 -1323
rect 779 -1319 780 -1317
rect 779 -1325 780 -1323
rect 786 -1319 787 -1317
rect 786 -1325 787 -1323
rect 789 -1325 790 -1323
rect 793 -1325 794 -1323
rect 796 -1325 797 -1323
rect 800 -1319 801 -1317
rect 800 -1325 801 -1323
rect 807 -1319 808 -1317
rect 810 -1319 811 -1317
rect 814 -1319 815 -1317
rect 817 -1319 818 -1317
rect 814 -1325 815 -1323
rect 817 -1325 818 -1323
rect 821 -1319 822 -1317
rect 821 -1325 822 -1323
rect 824 -1325 825 -1323
rect 828 -1319 829 -1317
rect 831 -1319 832 -1317
rect 828 -1325 829 -1323
rect 831 -1325 832 -1323
rect 835 -1319 836 -1317
rect 835 -1325 836 -1323
rect 842 -1319 843 -1317
rect 842 -1325 843 -1323
rect 849 -1319 850 -1317
rect 849 -1325 850 -1323
rect 856 -1319 857 -1317
rect 856 -1325 857 -1323
rect 863 -1319 864 -1317
rect 863 -1325 864 -1323
rect 870 -1319 871 -1317
rect 870 -1325 871 -1323
rect 877 -1319 878 -1317
rect 877 -1325 878 -1323
rect 884 -1319 885 -1317
rect 884 -1325 885 -1323
rect 891 -1319 892 -1317
rect 891 -1325 892 -1323
rect 898 -1319 899 -1317
rect 898 -1325 899 -1323
rect 905 -1319 906 -1317
rect 905 -1325 906 -1323
rect 912 -1319 913 -1317
rect 912 -1325 913 -1323
rect 919 -1319 920 -1317
rect 919 -1325 920 -1323
rect 926 -1319 927 -1317
rect 926 -1325 927 -1323
rect 933 -1319 934 -1317
rect 936 -1319 937 -1317
rect 933 -1325 934 -1323
rect 936 -1325 937 -1323
rect 940 -1319 941 -1317
rect 940 -1325 941 -1323
rect 947 -1319 948 -1317
rect 950 -1319 951 -1317
rect 947 -1325 948 -1323
rect 954 -1319 955 -1317
rect 954 -1325 955 -1323
rect 961 -1319 962 -1317
rect 961 -1325 962 -1323
rect 968 -1319 969 -1317
rect 968 -1325 969 -1323
rect 975 -1319 976 -1317
rect 978 -1319 979 -1317
rect 975 -1325 976 -1323
rect 978 -1325 979 -1323
rect 982 -1319 983 -1317
rect 985 -1319 986 -1317
rect 982 -1325 983 -1323
rect 985 -1325 986 -1323
rect 989 -1319 990 -1317
rect 989 -1325 990 -1323
rect 996 -1319 997 -1317
rect 999 -1319 1000 -1317
rect 996 -1325 997 -1323
rect 1003 -1319 1004 -1317
rect 1003 -1325 1004 -1323
rect 1010 -1319 1011 -1317
rect 1013 -1319 1014 -1317
rect 1010 -1325 1011 -1323
rect 1013 -1325 1014 -1323
rect 1017 -1319 1018 -1317
rect 1017 -1325 1018 -1323
rect 1024 -1319 1025 -1317
rect 1024 -1325 1025 -1323
rect 1031 -1319 1032 -1317
rect 1031 -1325 1032 -1323
rect 1038 -1319 1039 -1317
rect 1038 -1325 1039 -1323
rect 1045 -1319 1046 -1317
rect 1045 -1325 1046 -1323
rect 1052 -1319 1053 -1317
rect 1055 -1319 1056 -1317
rect 1052 -1325 1053 -1323
rect 1055 -1325 1056 -1323
rect 1059 -1319 1060 -1317
rect 1059 -1325 1060 -1323
rect 1066 -1319 1067 -1317
rect 1066 -1325 1067 -1323
rect 1073 -1319 1074 -1317
rect 1073 -1325 1074 -1323
rect 1080 -1319 1081 -1317
rect 1080 -1325 1081 -1323
rect 1087 -1319 1088 -1317
rect 1087 -1325 1088 -1323
rect 1094 -1319 1095 -1317
rect 1094 -1325 1095 -1323
rect 1101 -1319 1102 -1317
rect 1101 -1325 1102 -1323
rect 1108 -1319 1109 -1317
rect 1108 -1325 1109 -1323
rect 1115 -1319 1116 -1317
rect 1115 -1325 1116 -1323
rect 1122 -1319 1123 -1317
rect 1122 -1325 1123 -1323
rect 1129 -1319 1130 -1317
rect 1129 -1325 1130 -1323
rect 1136 -1319 1137 -1317
rect 1136 -1325 1137 -1323
rect 1143 -1319 1144 -1317
rect 1143 -1325 1144 -1323
rect 1150 -1319 1151 -1317
rect 1150 -1325 1151 -1323
rect 1157 -1319 1158 -1317
rect 1157 -1325 1158 -1323
rect 1164 -1319 1165 -1317
rect 1164 -1325 1165 -1323
rect 1171 -1319 1172 -1317
rect 1171 -1325 1172 -1323
rect 1178 -1319 1179 -1317
rect 1178 -1325 1179 -1323
rect 1185 -1319 1186 -1317
rect 1185 -1325 1186 -1323
rect 1192 -1319 1193 -1317
rect 1192 -1325 1193 -1323
rect 1199 -1319 1200 -1317
rect 1199 -1325 1200 -1323
rect 1206 -1319 1207 -1317
rect 1206 -1325 1207 -1323
rect 1213 -1319 1214 -1317
rect 1213 -1325 1214 -1323
rect 1220 -1319 1221 -1317
rect 1220 -1325 1221 -1323
rect 1227 -1319 1228 -1317
rect 1227 -1325 1228 -1323
rect 1234 -1319 1235 -1317
rect 1234 -1325 1235 -1323
rect 1241 -1319 1242 -1317
rect 1241 -1325 1242 -1323
rect 1248 -1319 1249 -1317
rect 1248 -1325 1249 -1323
rect 1255 -1319 1256 -1317
rect 1255 -1325 1256 -1323
rect 1262 -1319 1263 -1317
rect 1262 -1325 1263 -1323
rect 1269 -1319 1270 -1317
rect 1269 -1325 1270 -1323
rect 1276 -1319 1277 -1317
rect 1276 -1325 1277 -1323
rect 1283 -1319 1284 -1317
rect 1283 -1325 1284 -1323
rect 1290 -1319 1291 -1317
rect 1290 -1325 1291 -1323
rect 1297 -1319 1298 -1317
rect 1297 -1325 1298 -1323
rect 1304 -1319 1305 -1317
rect 1304 -1325 1305 -1323
rect 1311 -1319 1312 -1317
rect 1311 -1325 1312 -1323
rect 1318 -1319 1319 -1317
rect 1318 -1325 1319 -1323
rect 1325 -1319 1326 -1317
rect 1325 -1325 1326 -1323
rect 1332 -1319 1333 -1317
rect 1332 -1325 1333 -1323
rect 1339 -1319 1340 -1317
rect 1339 -1325 1340 -1323
rect 1346 -1319 1347 -1317
rect 1346 -1325 1347 -1323
rect 1353 -1319 1354 -1317
rect 1356 -1319 1357 -1317
rect 1353 -1325 1354 -1323
rect 1360 -1319 1361 -1317
rect 1360 -1325 1361 -1323
rect 1367 -1319 1368 -1317
rect 1367 -1325 1368 -1323
rect 1374 -1319 1375 -1317
rect 1374 -1325 1375 -1323
rect 1381 -1319 1382 -1317
rect 1381 -1325 1382 -1323
rect 1388 -1319 1389 -1317
rect 1388 -1325 1389 -1323
rect 1395 -1319 1396 -1317
rect 1395 -1325 1396 -1323
rect 1402 -1319 1403 -1317
rect 1402 -1325 1403 -1323
rect 1409 -1319 1410 -1317
rect 1409 -1325 1410 -1323
rect 1416 -1319 1417 -1317
rect 1416 -1325 1417 -1323
rect 1423 -1319 1424 -1317
rect 1423 -1325 1424 -1323
rect 1430 -1319 1431 -1317
rect 1430 -1325 1431 -1323
rect 1437 -1319 1438 -1317
rect 1437 -1325 1438 -1323
rect 1444 -1319 1445 -1317
rect 1444 -1325 1445 -1323
rect 1451 -1319 1452 -1317
rect 1451 -1325 1452 -1323
rect 1458 -1319 1459 -1317
rect 1458 -1325 1459 -1323
rect 1465 -1319 1466 -1317
rect 1465 -1325 1466 -1323
rect 1472 -1319 1473 -1317
rect 1472 -1325 1473 -1323
rect 1479 -1319 1480 -1317
rect 1479 -1325 1480 -1323
rect 1486 -1319 1487 -1317
rect 1486 -1325 1487 -1323
rect 1493 -1319 1494 -1317
rect 1493 -1325 1494 -1323
rect 1500 -1319 1501 -1317
rect 1500 -1325 1501 -1323
rect 1507 -1319 1508 -1317
rect 1507 -1325 1508 -1323
rect 1514 -1319 1515 -1317
rect 1514 -1325 1515 -1323
rect 1521 -1319 1522 -1317
rect 1521 -1325 1522 -1323
rect 1528 -1319 1529 -1317
rect 1528 -1325 1529 -1323
rect 1535 -1319 1536 -1317
rect 1535 -1325 1536 -1323
rect 1542 -1319 1543 -1317
rect 1542 -1325 1543 -1323
rect 1549 -1319 1550 -1317
rect 1549 -1325 1550 -1323
rect 1556 -1319 1557 -1317
rect 1556 -1325 1557 -1323
rect 1563 -1319 1564 -1317
rect 1563 -1325 1564 -1323
rect 1570 -1319 1571 -1317
rect 1570 -1325 1571 -1323
rect 1577 -1319 1578 -1317
rect 1577 -1325 1578 -1323
rect 1584 -1319 1585 -1317
rect 1584 -1325 1585 -1323
rect 1591 -1319 1592 -1317
rect 1591 -1325 1592 -1323
rect 1598 -1319 1599 -1317
rect 1598 -1325 1599 -1323
rect 1605 -1319 1606 -1317
rect 1605 -1325 1606 -1323
rect 1612 -1319 1613 -1317
rect 1612 -1325 1613 -1323
rect 1619 -1319 1620 -1317
rect 1619 -1325 1620 -1323
rect 1626 -1319 1627 -1317
rect 1626 -1325 1627 -1323
rect 1633 -1319 1634 -1317
rect 1633 -1325 1634 -1323
rect 1640 -1319 1641 -1317
rect 1640 -1325 1641 -1323
rect 1647 -1319 1648 -1317
rect 1647 -1325 1648 -1323
rect 1654 -1319 1655 -1317
rect 1654 -1325 1655 -1323
rect 1661 -1319 1662 -1317
rect 1661 -1325 1662 -1323
rect 1668 -1319 1669 -1317
rect 1668 -1325 1669 -1323
rect 1675 -1319 1676 -1317
rect 1675 -1325 1676 -1323
rect 1682 -1319 1683 -1317
rect 1682 -1325 1683 -1323
rect 1689 -1319 1690 -1317
rect 1689 -1325 1690 -1323
rect 1696 -1319 1697 -1317
rect 1696 -1325 1697 -1323
rect 1706 -1325 1707 -1323
rect 1713 -1319 1714 -1317
rect 1717 -1319 1718 -1317
rect 1717 -1325 1718 -1323
rect 1724 -1319 1725 -1317
rect 1724 -1325 1725 -1323
rect 1731 -1319 1732 -1317
rect 1734 -1319 1735 -1317
rect 1731 -1325 1732 -1323
rect 1734 -1325 1735 -1323
rect 1738 -1319 1739 -1317
rect 1738 -1325 1739 -1323
rect 16 -1474 17 -1472
rect 16 -1480 17 -1478
rect 26 -1474 27 -1472
rect 30 -1474 31 -1472
rect 30 -1480 31 -1478
rect 37 -1474 38 -1472
rect 37 -1480 38 -1478
rect 44 -1474 45 -1472
rect 44 -1480 45 -1478
rect 51 -1474 52 -1472
rect 51 -1480 52 -1478
rect 58 -1474 59 -1472
rect 61 -1474 62 -1472
rect 65 -1474 66 -1472
rect 65 -1480 66 -1478
rect 75 -1474 76 -1472
rect 72 -1480 73 -1478
rect 75 -1480 76 -1478
rect 79 -1474 80 -1472
rect 82 -1474 83 -1472
rect 79 -1480 80 -1478
rect 82 -1480 83 -1478
rect 86 -1474 87 -1472
rect 86 -1480 87 -1478
rect 93 -1474 94 -1472
rect 96 -1474 97 -1472
rect 93 -1480 94 -1478
rect 100 -1474 101 -1472
rect 100 -1480 101 -1478
rect 107 -1474 108 -1472
rect 110 -1474 111 -1472
rect 107 -1480 108 -1478
rect 117 -1474 118 -1472
rect 114 -1480 115 -1478
rect 117 -1480 118 -1478
rect 121 -1474 122 -1472
rect 121 -1480 122 -1478
rect 128 -1474 129 -1472
rect 128 -1480 129 -1478
rect 135 -1474 136 -1472
rect 135 -1480 136 -1478
rect 142 -1474 143 -1472
rect 142 -1480 143 -1478
rect 149 -1474 150 -1472
rect 149 -1480 150 -1478
rect 156 -1474 157 -1472
rect 156 -1480 157 -1478
rect 159 -1480 160 -1478
rect 163 -1474 164 -1472
rect 163 -1480 164 -1478
rect 170 -1474 171 -1472
rect 170 -1480 171 -1478
rect 177 -1474 178 -1472
rect 177 -1480 178 -1478
rect 184 -1474 185 -1472
rect 184 -1480 185 -1478
rect 191 -1474 192 -1472
rect 191 -1480 192 -1478
rect 198 -1474 199 -1472
rect 198 -1480 199 -1478
rect 205 -1474 206 -1472
rect 205 -1480 206 -1478
rect 212 -1474 213 -1472
rect 212 -1480 213 -1478
rect 219 -1474 220 -1472
rect 222 -1474 223 -1472
rect 219 -1480 220 -1478
rect 226 -1474 227 -1472
rect 229 -1474 230 -1472
rect 226 -1480 227 -1478
rect 229 -1480 230 -1478
rect 233 -1474 234 -1472
rect 233 -1480 234 -1478
rect 240 -1474 241 -1472
rect 240 -1480 241 -1478
rect 247 -1474 248 -1472
rect 247 -1480 248 -1478
rect 254 -1474 255 -1472
rect 254 -1480 255 -1478
rect 261 -1474 262 -1472
rect 264 -1474 265 -1472
rect 264 -1480 265 -1478
rect 268 -1474 269 -1472
rect 268 -1480 269 -1478
rect 275 -1474 276 -1472
rect 275 -1480 276 -1478
rect 282 -1474 283 -1472
rect 282 -1480 283 -1478
rect 289 -1474 290 -1472
rect 289 -1480 290 -1478
rect 299 -1480 300 -1478
rect 303 -1474 304 -1472
rect 303 -1480 304 -1478
rect 310 -1474 311 -1472
rect 310 -1480 311 -1478
rect 317 -1474 318 -1472
rect 317 -1480 318 -1478
rect 324 -1474 325 -1472
rect 324 -1480 325 -1478
rect 331 -1474 332 -1472
rect 331 -1480 332 -1478
rect 338 -1474 339 -1472
rect 338 -1480 339 -1478
rect 345 -1474 346 -1472
rect 345 -1480 346 -1478
rect 352 -1474 353 -1472
rect 352 -1480 353 -1478
rect 359 -1474 360 -1472
rect 359 -1480 360 -1478
rect 366 -1474 367 -1472
rect 366 -1480 367 -1478
rect 373 -1474 374 -1472
rect 373 -1480 374 -1478
rect 380 -1474 381 -1472
rect 380 -1480 381 -1478
rect 387 -1474 388 -1472
rect 387 -1480 388 -1478
rect 390 -1480 391 -1478
rect 394 -1474 395 -1472
rect 394 -1480 395 -1478
rect 401 -1474 402 -1472
rect 401 -1480 402 -1478
rect 408 -1474 409 -1472
rect 408 -1480 409 -1478
rect 411 -1480 412 -1478
rect 415 -1474 416 -1472
rect 418 -1474 419 -1472
rect 415 -1480 416 -1478
rect 418 -1480 419 -1478
rect 422 -1474 423 -1472
rect 422 -1480 423 -1478
rect 429 -1474 430 -1472
rect 429 -1480 430 -1478
rect 436 -1474 437 -1472
rect 436 -1480 437 -1478
rect 443 -1474 444 -1472
rect 443 -1480 444 -1478
rect 450 -1474 451 -1472
rect 450 -1480 451 -1478
rect 457 -1474 458 -1472
rect 457 -1480 458 -1478
rect 464 -1474 465 -1472
rect 464 -1480 465 -1478
rect 471 -1474 472 -1472
rect 471 -1480 472 -1478
rect 478 -1474 479 -1472
rect 478 -1480 479 -1478
rect 485 -1474 486 -1472
rect 485 -1480 486 -1478
rect 492 -1474 493 -1472
rect 492 -1480 493 -1478
rect 499 -1474 500 -1472
rect 502 -1474 503 -1472
rect 502 -1480 503 -1478
rect 506 -1474 507 -1472
rect 506 -1480 507 -1478
rect 513 -1474 514 -1472
rect 513 -1480 514 -1478
rect 520 -1474 521 -1472
rect 520 -1480 521 -1478
rect 527 -1474 528 -1472
rect 527 -1480 528 -1478
rect 534 -1474 535 -1472
rect 534 -1480 535 -1478
rect 541 -1474 542 -1472
rect 541 -1480 542 -1478
rect 548 -1474 549 -1472
rect 548 -1480 549 -1478
rect 555 -1474 556 -1472
rect 555 -1480 556 -1478
rect 558 -1480 559 -1478
rect 562 -1474 563 -1472
rect 562 -1480 563 -1478
rect 569 -1474 570 -1472
rect 569 -1480 570 -1478
rect 576 -1474 577 -1472
rect 576 -1480 577 -1478
rect 583 -1474 584 -1472
rect 583 -1480 584 -1478
rect 590 -1474 591 -1472
rect 593 -1474 594 -1472
rect 590 -1480 591 -1478
rect 593 -1480 594 -1478
rect 597 -1474 598 -1472
rect 600 -1474 601 -1472
rect 597 -1480 598 -1478
rect 604 -1474 605 -1472
rect 604 -1480 605 -1478
rect 611 -1474 612 -1472
rect 614 -1474 615 -1472
rect 614 -1480 615 -1478
rect 618 -1474 619 -1472
rect 618 -1480 619 -1478
rect 625 -1474 626 -1472
rect 625 -1480 626 -1478
rect 632 -1474 633 -1472
rect 635 -1474 636 -1472
rect 632 -1480 633 -1478
rect 635 -1480 636 -1478
rect 639 -1474 640 -1472
rect 642 -1474 643 -1472
rect 639 -1480 640 -1478
rect 642 -1480 643 -1478
rect 646 -1474 647 -1472
rect 646 -1480 647 -1478
rect 653 -1474 654 -1472
rect 653 -1480 654 -1478
rect 660 -1474 661 -1472
rect 660 -1480 661 -1478
rect 667 -1474 668 -1472
rect 667 -1480 668 -1478
rect 674 -1474 675 -1472
rect 677 -1474 678 -1472
rect 674 -1480 675 -1478
rect 677 -1480 678 -1478
rect 681 -1474 682 -1472
rect 681 -1480 682 -1478
rect 688 -1474 689 -1472
rect 688 -1480 689 -1478
rect 695 -1474 696 -1472
rect 695 -1480 696 -1478
rect 702 -1474 703 -1472
rect 702 -1480 703 -1478
rect 709 -1474 710 -1472
rect 709 -1480 710 -1478
rect 716 -1474 717 -1472
rect 719 -1474 720 -1472
rect 716 -1480 717 -1478
rect 719 -1480 720 -1478
rect 723 -1474 724 -1472
rect 726 -1474 727 -1472
rect 723 -1480 724 -1478
rect 726 -1480 727 -1478
rect 730 -1474 731 -1472
rect 733 -1474 734 -1472
rect 730 -1480 731 -1478
rect 733 -1480 734 -1478
rect 737 -1474 738 -1472
rect 737 -1480 738 -1478
rect 744 -1474 745 -1472
rect 744 -1480 745 -1478
rect 751 -1474 752 -1472
rect 751 -1480 752 -1478
rect 758 -1474 759 -1472
rect 758 -1480 759 -1478
rect 765 -1474 766 -1472
rect 765 -1480 766 -1478
rect 768 -1480 769 -1478
rect 772 -1474 773 -1472
rect 772 -1480 773 -1478
rect 779 -1474 780 -1472
rect 779 -1480 780 -1478
rect 786 -1474 787 -1472
rect 786 -1480 787 -1478
rect 793 -1474 794 -1472
rect 793 -1480 794 -1478
rect 800 -1474 801 -1472
rect 800 -1480 801 -1478
rect 807 -1474 808 -1472
rect 807 -1480 808 -1478
rect 814 -1474 815 -1472
rect 814 -1480 815 -1478
rect 821 -1474 822 -1472
rect 821 -1480 822 -1478
rect 828 -1474 829 -1472
rect 828 -1480 829 -1478
rect 835 -1474 836 -1472
rect 835 -1480 836 -1478
rect 842 -1474 843 -1472
rect 842 -1480 843 -1478
rect 849 -1474 850 -1472
rect 849 -1480 850 -1478
rect 856 -1474 857 -1472
rect 856 -1480 857 -1478
rect 863 -1474 864 -1472
rect 866 -1474 867 -1472
rect 863 -1480 864 -1478
rect 866 -1480 867 -1478
rect 870 -1474 871 -1472
rect 873 -1474 874 -1472
rect 870 -1480 871 -1478
rect 873 -1480 874 -1478
rect 877 -1474 878 -1472
rect 877 -1480 878 -1478
rect 884 -1474 885 -1472
rect 884 -1480 885 -1478
rect 891 -1474 892 -1472
rect 894 -1474 895 -1472
rect 891 -1480 892 -1478
rect 898 -1474 899 -1472
rect 901 -1474 902 -1472
rect 901 -1480 902 -1478
rect 905 -1474 906 -1472
rect 905 -1480 906 -1478
rect 912 -1474 913 -1472
rect 912 -1480 913 -1478
rect 919 -1474 920 -1472
rect 919 -1480 920 -1478
rect 926 -1474 927 -1472
rect 926 -1480 927 -1478
rect 933 -1474 934 -1472
rect 936 -1474 937 -1472
rect 933 -1480 934 -1478
rect 936 -1480 937 -1478
rect 940 -1474 941 -1472
rect 940 -1480 941 -1478
rect 947 -1474 948 -1472
rect 947 -1480 948 -1478
rect 954 -1474 955 -1472
rect 954 -1480 955 -1478
rect 961 -1474 962 -1472
rect 961 -1480 962 -1478
rect 968 -1474 969 -1472
rect 968 -1480 969 -1478
rect 975 -1474 976 -1472
rect 975 -1480 976 -1478
rect 982 -1474 983 -1472
rect 982 -1480 983 -1478
rect 989 -1474 990 -1472
rect 989 -1480 990 -1478
rect 996 -1474 997 -1472
rect 996 -1480 997 -1478
rect 1003 -1474 1004 -1472
rect 1003 -1480 1004 -1478
rect 1010 -1474 1011 -1472
rect 1010 -1480 1011 -1478
rect 1017 -1474 1018 -1472
rect 1017 -1480 1018 -1478
rect 1027 -1474 1028 -1472
rect 1024 -1480 1025 -1478
rect 1031 -1474 1032 -1472
rect 1031 -1480 1032 -1478
rect 1038 -1474 1039 -1472
rect 1038 -1480 1039 -1478
rect 1045 -1474 1046 -1472
rect 1045 -1480 1046 -1478
rect 1052 -1474 1053 -1472
rect 1052 -1480 1053 -1478
rect 1059 -1474 1060 -1472
rect 1059 -1480 1060 -1478
rect 1066 -1474 1067 -1472
rect 1069 -1474 1070 -1472
rect 1066 -1480 1067 -1478
rect 1073 -1474 1074 -1472
rect 1073 -1480 1074 -1478
rect 1080 -1474 1081 -1472
rect 1080 -1480 1081 -1478
rect 1087 -1474 1088 -1472
rect 1087 -1480 1088 -1478
rect 1094 -1474 1095 -1472
rect 1094 -1480 1095 -1478
rect 1101 -1474 1102 -1472
rect 1101 -1480 1102 -1478
rect 1108 -1474 1109 -1472
rect 1108 -1480 1109 -1478
rect 1115 -1474 1116 -1472
rect 1115 -1480 1116 -1478
rect 1122 -1474 1123 -1472
rect 1125 -1474 1126 -1472
rect 1122 -1480 1123 -1478
rect 1125 -1480 1126 -1478
rect 1129 -1474 1130 -1472
rect 1129 -1480 1130 -1478
rect 1139 -1474 1140 -1472
rect 1139 -1480 1140 -1478
rect 1143 -1474 1144 -1472
rect 1146 -1474 1147 -1472
rect 1143 -1480 1144 -1478
rect 1146 -1480 1147 -1478
rect 1150 -1474 1151 -1472
rect 1150 -1480 1151 -1478
rect 1157 -1474 1158 -1472
rect 1157 -1480 1158 -1478
rect 1164 -1474 1165 -1472
rect 1164 -1480 1165 -1478
rect 1171 -1474 1172 -1472
rect 1171 -1480 1172 -1478
rect 1178 -1474 1179 -1472
rect 1178 -1480 1179 -1478
rect 1185 -1474 1186 -1472
rect 1185 -1480 1186 -1478
rect 1192 -1474 1193 -1472
rect 1192 -1480 1193 -1478
rect 1199 -1474 1200 -1472
rect 1199 -1480 1200 -1478
rect 1206 -1474 1207 -1472
rect 1206 -1480 1207 -1478
rect 1213 -1474 1214 -1472
rect 1213 -1480 1214 -1478
rect 1220 -1474 1221 -1472
rect 1220 -1480 1221 -1478
rect 1227 -1474 1228 -1472
rect 1227 -1480 1228 -1478
rect 1234 -1474 1235 -1472
rect 1234 -1480 1235 -1478
rect 1241 -1474 1242 -1472
rect 1241 -1480 1242 -1478
rect 1248 -1474 1249 -1472
rect 1248 -1480 1249 -1478
rect 1255 -1474 1256 -1472
rect 1255 -1480 1256 -1478
rect 1262 -1474 1263 -1472
rect 1262 -1480 1263 -1478
rect 1269 -1474 1270 -1472
rect 1269 -1480 1270 -1478
rect 1276 -1474 1277 -1472
rect 1276 -1480 1277 -1478
rect 1283 -1474 1284 -1472
rect 1283 -1480 1284 -1478
rect 1290 -1474 1291 -1472
rect 1290 -1480 1291 -1478
rect 1297 -1474 1298 -1472
rect 1297 -1480 1298 -1478
rect 1304 -1474 1305 -1472
rect 1304 -1480 1305 -1478
rect 1311 -1474 1312 -1472
rect 1311 -1480 1312 -1478
rect 1318 -1474 1319 -1472
rect 1318 -1480 1319 -1478
rect 1325 -1474 1326 -1472
rect 1325 -1480 1326 -1478
rect 1332 -1474 1333 -1472
rect 1332 -1480 1333 -1478
rect 1339 -1474 1340 -1472
rect 1339 -1480 1340 -1478
rect 1346 -1474 1347 -1472
rect 1346 -1480 1347 -1478
rect 1353 -1474 1354 -1472
rect 1353 -1480 1354 -1478
rect 1360 -1474 1361 -1472
rect 1360 -1480 1361 -1478
rect 1367 -1474 1368 -1472
rect 1367 -1480 1368 -1478
rect 1374 -1474 1375 -1472
rect 1374 -1480 1375 -1478
rect 1381 -1474 1382 -1472
rect 1381 -1480 1382 -1478
rect 1388 -1474 1389 -1472
rect 1388 -1480 1389 -1478
rect 1395 -1474 1396 -1472
rect 1395 -1480 1396 -1478
rect 1402 -1474 1403 -1472
rect 1402 -1480 1403 -1478
rect 1409 -1474 1410 -1472
rect 1409 -1480 1410 -1478
rect 1416 -1474 1417 -1472
rect 1416 -1480 1417 -1478
rect 1423 -1474 1424 -1472
rect 1423 -1480 1424 -1478
rect 1430 -1474 1431 -1472
rect 1430 -1480 1431 -1478
rect 1437 -1474 1438 -1472
rect 1437 -1480 1438 -1478
rect 1444 -1474 1445 -1472
rect 1444 -1480 1445 -1478
rect 1451 -1474 1452 -1472
rect 1451 -1480 1452 -1478
rect 1458 -1474 1459 -1472
rect 1458 -1480 1459 -1478
rect 1465 -1474 1466 -1472
rect 1465 -1480 1466 -1478
rect 1472 -1474 1473 -1472
rect 1472 -1480 1473 -1478
rect 1479 -1474 1480 -1472
rect 1479 -1480 1480 -1478
rect 1486 -1474 1487 -1472
rect 1486 -1480 1487 -1478
rect 1493 -1474 1494 -1472
rect 1493 -1480 1494 -1478
rect 1500 -1474 1501 -1472
rect 1500 -1480 1501 -1478
rect 1507 -1474 1508 -1472
rect 1507 -1480 1508 -1478
rect 1514 -1474 1515 -1472
rect 1514 -1480 1515 -1478
rect 1521 -1474 1522 -1472
rect 1521 -1480 1522 -1478
rect 1528 -1474 1529 -1472
rect 1528 -1480 1529 -1478
rect 1535 -1474 1536 -1472
rect 1535 -1480 1536 -1478
rect 1542 -1474 1543 -1472
rect 1542 -1480 1543 -1478
rect 1549 -1474 1550 -1472
rect 1549 -1480 1550 -1478
rect 1556 -1474 1557 -1472
rect 1556 -1480 1557 -1478
rect 1563 -1474 1564 -1472
rect 1563 -1480 1564 -1478
rect 1570 -1474 1571 -1472
rect 1570 -1480 1571 -1478
rect 1577 -1474 1578 -1472
rect 1577 -1480 1578 -1478
rect 1584 -1474 1585 -1472
rect 1584 -1480 1585 -1478
rect 1591 -1474 1592 -1472
rect 1591 -1480 1592 -1478
rect 1598 -1474 1599 -1472
rect 1598 -1480 1599 -1478
rect 1605 -1474 1606 -1472
rect 1605 -1480 1606 -1478
rect 1612 -1474 1613 -1472
rect 1612 -1480 1613 -1478
rect 1619 -1474 1620 -1472
rect 1619 -1480 1620 -1478
rect 1626 -1474 1627 -1472
rect 1626 -1480 1627 -1478
rect 1633 -1474 1634 -1472
rect 1633 -1480 1634 -1478
rect 1640 -1474 1641 -1472
rect 1640 -1480 1641 -1478
rect 1647 -1474 1648 -1472
rect 1647 -1480 1648 -1478
rect 1654 -1474 1655 -1472
rect 1654 -1480 1655 -1478
rect 1661 -1474 1662 -1472
rect 1661 -1480 1662 -1478
rect 1668 -1474 1669 -1472
rect 1668 -1480 1669 -1478
rect 1675 -1474 1676 -1472
rect 1675 -1480 1676 -1478
rect 1682 -1474 1683 -1472
rect 1682 -1480 1683 -1478
rect 1689 -1474 1690 -1472
rect 1689 -1480 1690 -1478
rect 1699 -1474 1700 -1472
rect 1703 -1474 1704 -1472
rect 1703 -1480 1704 -1478
rect 1710 -1474 1711 -1472
rect 1710 -1480 1711 -1478
rect 1717 -1474 1718 -1472
rect 1720 -1474 1721 -1472
rect 1717 -1480 1718 -1478
rect 1720 -1480 1721 -1478
rect 1724 -1474 1725 -1472
rect 1724 -1480 1725 -1478
rect 1745 -1474 1746 -1472
rect 1745 -1480 1746 -1478
rect 23 -1611 24 -1609
rect 23 -1617 24 -1615
rect 30 -1611 31 -1609
rect 30 -1617 31 -1615
rect 44 -1611 45 -1609
rect 44 -1617 45 -1615
rect 51 -1611 52 -1609
rect 51 -1617 52 -1615
rect 58 -1611 59 -1609
rect 61 -1611 62 -1609
rect 65 -1611 66 -1609
rect 68 -1611 69 -1609
rect 72 -1611 73 -1609
rect 72 -1617 73 -1615
rect 79 -1611 80 -1609
rect 79 -1617 80 -1615
rect 86 -1611 87 -1609
rect 86 -1617 87 -1615
rect 93 -1611 94 -1609
rect 96 -1611 97 -1609
rect 93 -1617 94 -1615
rect 96 -1617 97 -1615
rect 100 -1611 101 -1609
rect 100 -1617 101 -1615
rect 107 -1611 108 -1609
rect 107 -1617 108 -1615
rect 114 -1611 115 -1609
rect 114 -1617 115 -1615
rect 121 -1611 122 -1609
rect 121 -1617 122 -1615
rect 128 -1611 129 -1609
rect 128 -1617 129 -1615
rect 135 -1611 136 -1609
rect 135 -1617 136 -1615
rect 142 -1611 143 -1609
rect 142 -1617 143 -1615
rect 149 -1611 150 -1609
rect 149 -1617 150 -1615
rect 156 -1611 157 -1609
rect 156 -1617 157 -1615
rect 163 -1611 164 -1609
rect 163 -1617 164 -1615
rect 170 -1611 171 -1609
rect 170 -1617 171 -1615
rect 177 -1611 178 -1609
rect 177 -1617 178 -1615
rect 184 -1611 185 -1609
rect 184 -1617 185 -1615
rect 191 -1611 192 -1609
rect 194 -1611 195 -1609
rect 191 -1617 192 -1615
rect 194 -1617 195 -1615
rect 198 -1611 199 -1609
rect 198 -1617 199 -1615
rect 205 -1611 206 -1609
rect 208 -1611 209 -1609
rect 205 -1617 206 -1615
rect 208 -1617 209 -1615
rect 212 -1611 213 -1609
rect 212 -1617 213 -1615
rect 219 -1611 220 -1609
rect 219 -1617 220 -1615
rect 226 -1611 227 -1609
rect 226 -1617 227 -1615
rect 233 -1611 234 -1609
rect 233 -1617 234 -1615
rect 240 -1611 241 -1609
rect 240 -1617 241 -1615
rect 247 -1611 248 -1609
rect 247 -1617 248 -1615
rect 257 -1611 258 -1609
rect 254 -1617 255 -1615
rect 261 -1611 262 -1609
rect 261 -1617 262 -1615
rect 268 -1617 269 -1615
rect 271 -1617 272 -1615
rect 275 -1611 276 -1609
rect 275 -1617 276 -1615
rect 282 -1611 283 -1609
rect 282 -1617 283 -1615
rect 289 -1611 290 -1609
rect 292 -1611 293 -1609
rect 289 -1617 290 -1615
rect 296 -1611 297 -1609
rect 296 -1617 297 -1615
rect 303 -1611 304 -1609
rect 303 -1617 304 -1615
rect 310 -1611 311 -1609
rect 310 -1617 311 -1615
rect 320 -1617 321 -1615
rect 324 -1611 325 -1609
rect 324 -1617 325 -1615
rect 331 -1611 332 -1609
rect 331 -1617 332 -1615
rect 338 -1611 339 -1609
rect 338 -1617 339 -1615
rect 345 -1611 346 -1609
rect 345 -1617 346 -1615
rect 352 -1611 353 -1609
rect 352 -1617 353 -1615
rect 359 -1611 360 -1609
rect 359 -1617 360 -1615
rect 366 -1611 367 -1609
rect 369 -1611 370 -1609
rect 366 -1617 367 -1615
rect 369 -1617 370 -1615
rect 373 -1611 374 -1609
rect 373 -1617 374 -1615
rect 380 -1611 381 -1609
rect 383 -1611 384 -1609
rect 380 -1617 381 -1615
rect 383 -1617 384 -1615
rect 387 -1611 388 -1609
rect 387 -1617 388 -1615
rect 394 -1611 395 -1609
rect 394 -1617 395 -1615
rect 401 -1611 402 -1609
rect 401 -1617 402 -1615
rect 408 -1611 409 -1609
rect 408 -1617 409 -1615
rect 415 -1611 416 -1609
rect 415 -1617 416 -1615
rect 422 -1611 423 -1609
rect 422 -1617 423 -1615
rect 429 -1611 430 -1609
rect 429 -1617 430 -1615
rect 436 -1611 437 -1609
rect 436 -1617 437 -1615
rect 443 -1611 444 -1609
rect 443 -1617 444 -1615
rect 450 -1611 451 -1609
rect 450 -1617 451 -1615
rect 457 -1611 458 -1609
rect 457 -1617 458 -1615
rect 464 -1611 465 -1609
rect 464 -1617 465 -1615
rect 471 -1611 472 -1609
rect 474 -1611 475 -1609
rect 471 -1617 472 -1615
rect 478 -1611 479 -1609
rect 478 -1617 479 -1615
rect 485 -1611 486 -1609
rect 485 -1617 486 -1615
rect 492 -1611 493 -1609
rect 492 -1617 493 -1615
rect 495 -1617 496 -1615
rect 499 -1611 500 -1609
rect 499 -1617 500 -1615
rect 506 -1611 507 -1609
rect 506 -1617 507 -1615
rect 513 -1611 514 -1609
rect 513 -1617 514 -1615
rect 520 -1611 521 -1609
rect 520 -1617 521 -1615
rect 527 -1611 528 -1609
rect 527 -1617 528 -1615
rect 530 -1617 531 -1615
rect 534 -1611 535 -1609
rect 534 -1617 535 -1615
rect 541 -1611 542 -1609
rect 544 -1611 545 -1609
rect 541 -1617 542 -1615
rect 544 -1617 545 -1615
rect 548 -1611 549 -1609
rect 548 -1617 549 -1615
rect 555 -1611 556 -1609
rect 555 -1617 556 -1615
rect 562 -1611 563 -1609
rect 562 -1617 563 -1615
rect 565 -1617 566 -1615
rect 569 -1611 570 -1609
rect 569 -1617 570 -1615
rect 576 -1611 577 -1609
rect 576 -1617 577 -1615
rect 583 -1611 584 -1609
rect 583 -1617 584 -1615
rect 590 -1611 591 -1609
rect 590 -1617 591 -1615
rect 597 -1611 598 -1609
rect 597 -1617 598 -1615
rect 604 -1611 605 -1609
rect 607 -1611 608 -1609
rect 604 -1617 605 -1615
rect 607 -1617 608 -1615
rect 611 -1611 612 -1609
rect 614 -1611 615 -1609
rect 611 -1617 612 -1615
rect 614 -1617 615 -1615
rect 618 -1611 619 -1609
rect 621 -1611 622 -1609
rect 618 -1617 619 -1615
rect 621 -1617 622 -1615
rect 625 -1611 626 -1609
rect 632 -1611 633 -1609
rect 632 -1617 633 -1615
rect 639 -1611 640 -1609
rect 639 -1617 640 -1615
rect 646 -1611 647 -1609
rect 646 -1617 647 -1615
rect 653 -1611 654 -1609
rect 653 -1617 654 -1615
rect 660 -1611 661 -1609
rect 660 -1617 661 -1615
rect 667 -1611 668 -1609
rect 670 -1611 671 -1609
rect 667 -1617 668 -1615
rect 670 -1617 671 -1615
rect 674 -1611 675 -1609
rect 674 -1617 675 -1615
rect 681 -1611 682 -1609
rect 681 -1617 682 -1615
rect 688 -1611 689 -1609
rect 688 -1617 689 -1615
rect 695 -1611 696 -1609
rect 695 -1617 696 -1615
rect 702 -1611 703 -1609
rect 702 -1617 703 -1615
rect 709 -1611 710 -1609
rect 712 -1611 713 -1609
rect 709 -1617 710 -1615
rect 712 -1617 713 -1615
rect 716 -1611 717 -1609
rect 719 -1611 720 -1609
rect 716 -1617 717 -1615
rect 719 -1617 720 -1615
rect 723 -1611 724 -1609
rect 726 -1611 727 -1609
rect 723 -1617 724 -1615
rect 726 -1617 727 -1615
rect 730 -1611 731 -1609
rect 730 -1617 731 -1615
rect 737 -1611 738 -1609
rect 740 -1611 741 -1609
rect 737 -1617 738 -1615
rect 740 -1617 741 -1615
rect 744 -1611 745 -1609
rect 747 -1611 748 -1609
rect 747 -1617 748 -1615
rect 751 -1611 752 -1609
rect 751 -1617 752 -1615
rect 758 -1611 759 -1609
rect 761 -1611 762 -1609
rect 758 -1617 759 -1615
rect 761 -1617 762 -1615
rect 765 -1611 766 -1609
rect 765 -1617 766 -1615
rect 772 -1611 773 -1609
rect 772 -1617 773 -1615
rect 779 -1611 780 -1609
rect 779 -1617 780 -1615
rect 786 -1611 787 -1609
rect 786 -1617 787 -1615
rect 793 -1611 794 -1609
rect 796 -1611 797 -1609
rect 793 -1617 794 -1615
rect 796 -1617 797 -1615
rect 800 -1611 801 -1609
rect 800 -1617 801 -1615
rect 807 -1611 808 -1609
rect 807 -1617 808 -1615
rect 814 -1611 815 -1609
rect 814 -1617 815 -1615
rect 821 -1611 822 -1609
rect 821 -1617 822 -1615
rect 828 -1611 829 -1609
rect 828 -1617 829 -1615
rect 835 -1611 836 -1609
rect 835 -1617 836 -1615
rect 842 -1611 843 -1609
rect 842 -1617 843 -1615
rect 849 -1611 850 -1609
rect 849 -1617 850 -1615
rect 856 -1611 857 -1609
rect 856 -1617 857 -1615
rect 863 -1611 864 -1609
rect 863 -1617 864 -1615
rect 870 -1611 871 -1609
rect 870 -1617 871 -1615
rect 877 -1611 878 -1609
rect 877 -1617 878 -1615
rect 884 -1611 885 -1609
rect 884 -1617 885 -1615
rect 891 -1611 892 -1609
rect 891 -1617 892 -1615
rect 898 -1611 899 -1609
rect 898 -1617 899 -1615
rect 905 -1611 906 -1609
rect 905 -1617 906 -1615
rect 912 -1611 913 -1609
rect 912 -1617 913 -1615
rect 919 -1611 920 -1609
rect 919 -1617 920 -1615
rect 926 -1611 927 -1609
rect 929 -1611 930 -1609
rect 926 -1617 927 -1615
rect 929 -1617 930 -1615
rect 933 -1611 934 -1609
rect 933 -1617 934 -1615
rect 940 -1611 941 -1609
rect 940 -1617 941 -1615
rect 947 -1611 948 -1609
rect 947 -1617 948 -1615
rect 954 -1611 955 -1609
rect 954 -1617 955 -1615
rect 961 -1611 962 -1609
rect 961 -1617 962 -1615
rect 968 -1611 969 -1609
rect 968 -1617 969 -1615
rect 975 -1611 976 -1609
rect 975 -1617 976 -1615
rect 982 -1611 983 -1609
rect 982 -1617 983 -1615
rect 989 -1611 990 -1609
rect 989 -1617 990 -1615
rect 996 -1611 997 -1609
rect 996 -1617 997 -1615
rect 1003 -1611 1004 -1609
rect 1003 -1617 1004 -1615
rect 1010 -1611 1011 -1609
rect 1010 -1617 1011 -1615
rect 1017 -1611 1018 -1609
rect 1020 -1611 1021 -1609
rect 1017 -1617 1018 -1615
rect 1020 -1617 1021 -1615
rect 1024 -1611 1025 -1609
rect 1024 -1617 1025 -1615
rect 1031 -1611 1032 -1609
rect 1031 -1617 1032 -1615
rect 1038 -1611 1039 -1609
rect 1038 -1617 1039 -1615
rect 1045 -1611 1046 -1609
rect 1048 -1611 1049 -1609
rect 1045 -1617 1046 -1615
rect 1048 -1617 1049 -1615
rect 1052 -1611 1053 -1609
rect 1052 -1617 1053 -1615
rect 1062 -1611 1063 -1609
rect 1059 -1617 1060 -1615
rect 1066 -1611 1067 -1609
rect 1066 -1617 1067 -1615
rect 1073 -1611 1074 -1609
rect 1073 -1617 1074 -1615
rect 1080 -1611 1081 -1609
rect 1080 -1617 1081 -1615
rect 1087 -1611 1088 -1609
rect 1087 -1617 1088 -1615
rect 1094 -1611 1095 -1609
rect 1094 -1617 1095 -1615
rect 1101 -1611 1102 -1609
rect 1104 -1611 1105 -1609
rect 1101 -1617 1102 -1615
rect 1104 -1617 1105 -1615
rect 1108 -1611 1109 -1609
rect 1108 -1617 1109 -1615
rect 1115 -1611 1116 -1609
rect 1118 -1611 1119 -1609
rect 1115 -1617 1116 -1615
rect 1118 -1617 1119 -1615
rect 1122 -1611 1123 -1609
rect 1122 -1617 1123 -1615
rect 1129 -1611 1130 -1609
rect 1129 -1617 1130 -1615
rect 1136 -1611 1137 -1609
rect 1136 -1617 1137 -1615
rect 1143 -1611 1144 -1609
rect 1143 -1617 1144 -1615
rect 1153 -1611 1154 -1609
rect 1150 -1617 1151 -1615
rect 1153 -1617 1154 -1615
rect 1157 -1611 1158 -1609
rect 1157 -1617 1158 -1615
rect 1164 -1611 1165 -1609
rect 1164 -1617 1165 -1615
rect 1171 -1611 1172 -1609
rect 1171 -1617 1172 -1615
rect 1178 -1611 1179 -1609
rect 1178 -1617 1179 -1615
rect 1185 -1611 1186 -1609
rect 1185 -1617 1186 -1615
rect 1192 -1611 1193 -1609
rect 1192 -1617 1193 -1615
rect 1199 -1611 1200 -1609
rect 1199 -1617 1200 -1615
rect 1206 -1611 1207 -1609
rect 1206 -1617 1207 -1615
rect 1213 -1611 1214 -1609
rect 1213 -1617 1214 -1615
rect 1220 -1611 1221 -1609
rect 1220 -1617 1221 -1615
rect 1227 -1611 1228 -1609
rect 1227 -1617 1228 -1615
rect 1234 -1611 1235 -1609
rect 1234 -1617 1235 -1615
rect 1241 -1611 1242 -1609
rect 1241 -1617 1242 -1615
rect 1248 -1611 1249 -1609
rect 1248 -1617 1249 -1615
rect 1255 -1611 1256 -1609
rect 1258 -1611 1259 -1609
rect 1255 -1617 1256 -1615
rect 1262 -1611 1263 -1609
rect 1262 -1617 1263 -1615
rect 1269 -1611 1270 -1609
rect 1269 -1617 1270 -1615
rect 1276 -1611 1277 -1609
rect 1276 -1617 1277 -1615
rect 1283 -1611 1284 -1609
rect 1283 -1617 1284 -1615
rect 1290 -1611 1291 -1609
rect 1290 -1617 1291 -1615
rect 1297 -1611 1298 -1609
rect 1297 -1617 1298 -1615
rect 1304 -1611 1305 -1609
rect 1304 -1617 1305 -1615
rect 1311 -1611 1312 -1609
rect 1311 -1617 1312 -1615
rect 1318 -1611 1319 -1609
rect 1318 -1617 1319 -1615
rect 1325 -1611 1326 -1609
rect 1325 -1617 1326 -1615
rect 1332 -1611 1333 -1609
rect 1332 -1617 1333 -1615
rect 1339 -1611 1340 -1609
rect 1339 -1617 1340 -1615
rect 1346 -1611 1347 -1609
rect 1346 -1617 1347 -1615
rect 1353 -1611 1354 -1609
rect 1353 -1617 1354 -1615
rect 1360 -1611 1361 -1609
rect 1360 -1617 1361 -1615
rect 1367 -1611 1368 -1609
rect 1367 -1617 1368 -1615
rect 1374 -1611 1375 -1609
rect 1374 -1617 1375 -1615
rect 1381 -1611 1382 -1609
rect 1381 -1617 1382 -1615
rect 1384 -1617 1385 -1615
rect 1388 -1611 1389 -1609
rect 1388 -1617 1389 -1615
rect 1395 -1611 1396 -1609
rect 1395 -1617 1396 -1615
rect 1402 -1611 1403 -1609
rect 1402 -1617 1403 -1615
rect 1409 -1611 1410 -1609
rect 1409 -1617 1410 -1615
rect 1416 -1611 1417 -1609
rect 1416 -1617 1417 -1615
rect 1423 -1611 1424 -1609
rect 1423 -1617 1424 -1615
rect 1430 -1611 1431 -1609
rect 1430 -1617 1431 -1615
rect 1437 -1611 1438 -1609
rect 1437 -1617 1438 -1615
rect 1444 -1611 1445 -1609
rect 1444 -1617 1445 -1615
rect 1451 -1611 1452 -1609
rect 1451 -1617 1452 -1615
rect 1458 -1611 1459 -1609
rect 1458 -1617 1459 -1615
rect 1465 -1611 1466 -1609
rect 1465 -1617 1466 -1615
rect 1472 -1611 1473 -1609
rect 1472 -1617 1473 -1615
rect 1479 -1611 1480 -1609
rect 1479 -1617 1480 -1615
rect 1486 -1611 1487 -1609
rect 1486 -1617 1487 -1615
rect 1493 -1611 1494 -1609
rect 1493 -1617 1494 -1615
rect 1500 -1611 1501 -1609
rect 1500 -1617 1501 -1615
rect 1507 -1611 1508 -1609
rect 1507 -1617 1508 -1615
rect 1514 -1611 1515 -1609
rect 1514 -1617 1515 -1615
rect 1521 -1611 1522 -1609
rect 1521 -1617 1522 -1615
rect 1528 -1611 1529 -1609
rect 1528 -1617 1529 -1615
rect 1535 -1611 1536 -1609
rect 1535 -1617 1536 -1615
rect 1542 -1611 1543 -1609
rect 1542 -1617 1543 -1615
rect 1549 -1611 1550 -1609
rect 1549 -1617 1550 -1615
rect 1556 -1611 1557 -1609
rect 1556 -1617 1557 -1615
rect 1563 -1611 1564 -1609
rect 1563 -1617 1564 -1615
rect 1570 -1611 1571 -1609
rect 1570 -1617 1571 -1615
rect 1577 -1611 1578 -1609
rect 1577 -1617 1578 -1615
rect 1584 -1611 1585 -1609
rect 1584 -1617 1585 -1615
rect 1591 -1611 1592 -1609
rect 1591 -1617 1592 -1615
rect 1598 -1611 1599 -1609
rect 1598 -1617 1599 -1615
rect 1605 -1611 1606 -1609
rect 1605 -1617 1606 -1615
rect 1612 -1611 1613 -1609
rect 1612 -1617 1613 -1615
rect 1619 -1611 1620 -1609
rect 1619 -1617 1620 -1615
rect 1626 -1611 1627 -1609
rect 1626 -1617 1627 -1615
rect 1633 -1611 1634 -1609
rect 1633 -1617 1634 -1615
rect 1640 -1611 1641 -1609
rect 1640 -1617 1641 -1615
rect 1647 -1611 1648 -1609
rect 1647 -1617 1648 -1615
rect 1654 -1611 1655 -1609
rect 1654 -1617 1655 -1615
rect 1661 -1611 1662 -1609
rect 1661 -1617 1662 -1615
rect 1668 -1611 1669 -1609
rect 1668 -1617 1669 -1615
rect 1675 -1611 1676 -1609
rect 1675 -1617 1676 -1615
rect 1682 -1611 1683 -1609
rect 1682 -1617 1683 -1615
rect 1689 -1611 1690 -1609
rect 1689 -1617 1690 -1615
rect 1696 -1611 1697 -1609
rect 1696 -1617 1697 -1615
rect 1703 -1611 1704 -1609
rect 1706 -1611 1707 -1609
rect 1703 -1617 1704 -1615
rect 1706 -1617 1707 -1615
rect 1710 -1611 1711 -1609
rect 1713 -1611 1714 -1609
rect 1710 -1617 1711 -1615
rect 1717 -1611 1718 -1609
rect 1717 -1617 1718 -1615
rect 1752 -1611 1753 -1609
rect 1752 -1617 1753 -1615
rect 16 -1738 17 -1736
rect 37 -1738 38 -1736
rect 37 -1744 38 -1742
rect 44 -1738 45 -1736
rect 44 -1744 45 -1742
rect 51 -1738 52 -1736
rect 51 -1744 52 -1742
rect 58 -1738 59 -1736
rect 61 -1738 62 -1736
rect 61 -1744 62 -1742
rect 65 -1738 66 -1736
rect 65 -1744 66 -1742
rect 72 -1738 73 -1736
rect 72 -1744 73 -1742
rect 79 -1738 80 -1736
rect 79 -1744 80 -1742
rect 86 -1738 87 -1736
rect 86 -1744 87 -1742
rect 93 -1738 94 -1736
rect 93 -1744 94 -1742
rect 100 -1738 101 -1736
rect 100 -1744 101 -1742
rect 107 -1738 108 -1736
rect 107 -1744 108 -1742
rect 114 -1738 115 -1736
rect 114 -1744 115 -1742
rect 121 -1738 122 -1736
rect 121 -1744 122 -1742
rect 128 -1738 129 -1736
rect 128 -1744 129 -1742
rect 135 -1738 136 -1736
rect 135 -1744 136 -1742
rect 142 -1738 143 -1736
rect 142 -1744 143 -1742
rect 149 -1738 150 -1736
rect 149 -1744 150 -1742
rect 156 -1738 157 -1736
rect 159 -1738 160 -1736
rect 156 -1744 157 -1742
rect 159 -1744 160 -1742
rect 163 -1738 164 -1736
rect 163 -1744 164 -1742
rect 170 -1738 171 -1736
rect 173 -1738 174 -1736
rect 170 -1744 171 -1742
rect 177 -1738 178 -1736
rect 177 -1744 178 -1742
rect 180 -1744 181 -1742
rect 184 -1738 185 -1736
rect 184 -1744 185 -1742
rect 191 -1738 192 -1736
rect 191 -1744 192 -1742
rect 194 -1744 195 -1742
rect 198 -1738 199 -1736
rect 198 -1744 199 -1742
rect 205 -1738 206 -1736
rect 205 -1744 206 -1742
rect 212 -1738 213 -1736
rect 212 -1744 213 -1742
rect 219 -1738 220 -1736
rect 219 -1744 220 -1742
rect 226 -1738 227 -1736
rect 226 -1744 227 -1742
rect 233 -1738 234 -1736
rect 233 -1744 234 -1742
rect 240 -1738 241 -1736
rect 240 -1744 241 -1742
rect 247 -1738 248 -1736
rect 247 -1744 248 -1742
rect 257 -1738 258 -1736
rect 254 -1744 255 -1742
rect 257 -1744 258 -1742
rect 264 -1738 265 -1736
rect 264 -1744 265 -1742
rect 268 -1738 269 -1736
rect 268 -1744 269 -1742
rect 275 -1738 276 -1736
rect 278 -1738 279 -1736
rect 275 -1744 276 -1742
rect 282 -1738 283 -1736
rect 282 -1744 283 -1742
rect 289 -1738 290 -1736
rect 289 -1744 290 -1742
rect 296 -1738 297 -1736
rect 296 -1744 297 -1742
rect 303 -1738 304 -1736
rect 303 -1744 304 -1742
rect 310 -1738 311 -1736
rect 310 -1744 311 -1742
rect 317 -1738 318 -1736
rect 317 -1744 318 -1742
rect 324 -1738 325 -1736
rect 324 -1744 325 -1742
rect 331 -1738 332 -1736
rect 331 -1744 332 -1742
rect 338 -1738 339 -1736
rect 338 -1744 339 -1742
rect 345 -1738 346 -1736
rect 348 -1738 349 -1736
rect 348 -1744 349 -1742
rect 352 -1738 353 -1736
rect 352 -1744 353 -1742
rect 359 -1738 360 -1736
rect 359 -1744 360 -1742
rect 366 -1738 367 -1736
rect 366 -1744 367 -1742
rect 373 -1738 374 -1736
rect 373 -1744 374 -1742
rect 380 -1738 381 -1736
rect 380 -1744 381 -1742
rect 387 -1738 388 -1736
rect 387 -1744 388 -1742
rect 394 -1738 395 -1736
rect 394 -1744 395 -1742
rect 401 -1738 402 -1736
rect 401 -1744 402 -1742
rect 411 -1738 412 -1736
rect 411 -1744 412 -1742
rect 415 -1738 416 -1736
rect 415 -1744 416 -1742
rect 422 -1738 423 -1736
rect 422 -1744 423 -1742
rect 429 -1738 430 -1736
rect 432 -1738 433 -1736
rect 432 -1744 433 -1742
rect 436 -1738 437 -1736
rect 436 -1744 437 -1742
rect 443 -1738 444 -1736
rect 443 -1744 444 -1742
rect 450 -1738 451 -1736
rect 450 -1744 451 -1742
rect 457 -1738 458 -1736
rect 457 -1744 458 -1742
rect 464 -1738 465 -1736
rect 464 -1744 465 -1742
rect 471 -1738 472 -1736
rect 471 -1744 472 -1742
rect 478 -1738 479 -1736
rect 481 -1738 482 -1736
rect 478 -1744 479 -1742
rect 481 -1744 482 -1742
rect 485 -1738 486 -1736
rect 485 -1744 486 -1742
rect 492 -1738 493 -1736
rect 492 -1744 493 -1742
rect 499 -1738 500 -1736
rect 499 -1744 500 -1742
rect 506 -1738 507 -1736
rect 506 -1744 507 -1742
rect 513 -1738 514 -1736
rect 513 -1744 514 -1742
rect 520 -1738 521 -1736
rect 520 -1744 521 -1742
rect 527 -1738 528 -1736
rect 530 -1738 531 -1736
rect 527 -1744 528 -1742
rect 530 -1744 531 -1742
rect 534 -1738 535 -1736
rect 534 -1744 535 -1742
rect 541 -1738 542 -1736
rect 544 -1738 545 -1736
rect 541 -1744 542 -1742
rect 548 -1738 549 -1736
rect 548 -1744 549 -1742
rect 555 -1738 556 -1736
rect 555 -1744 556 -1742
rect 562 -1738 563 -1736
rect 562 -1744 563 -1742
rect 569 -1738 570 -1736
rect 569 -1744 570 -1742
rect 576 -1738 577 -1736
rect 576 -1744 577 -1742
rect 583 -1738 584 -1736
rect 583 -1744 584 -1742
rect 590 -1738 591 -1736
rect 590 -1744 591 -1742
rect 597 -1738 598 -1736
rect 597 -1744 598 -1742
rect 604 -1738 605 -1736
rect 604 -1744 605 -1742
rect 611 -1738 612 -1736
rect 611 -1744 612 -1742
rect 618 -1738 619 -1736
rect 618 -1744 619 -1742
rect 625 -1744 626 -1742
rect 632 -1738 633 -1736
rect 632 -1744 633 -1742
rect 639 -1738 640 -1736
rect 639 -1744 640 -1742
rect 646 -1738 647 -1736
rect 646 -1744 647 -1742
rect 653 -1738 654 -1736
rect 653 -1744 654 -1742
rect 660 -1738 661 -1736
rect 660 -1744 661 -1742
rect 667 -1738 668 -1736
rect 667 -1744 668 -1742
rect 677 -1738 678 -1736
rect 674 -1744 675 -1742
rect 677 -1744 678 -1742
rect 681 -1738 682 -1736
rect 681 -1744 682 -1742
rect 688 -1738 689 -1736
rect 688 -1744 689 -1742
rect 691 -1744 692 -1742
rect 695 -1738 696 -1736
rect 695 -1744 696 -1742
rect 702 -1744 703 -1742
rect 709 -1738 710 -1736
rect 709 -1744 710 -1742
rect 716 -1738 717 -1736
rect 716 -1744 717 -1742
rect 723 -1738 724 -1736
rect 726 -1738 727 -1736
rect 723 -1744 724 -1742
rect 726 -1744 727 -1742
rect 730 -1738 731 -1736
rect 733 -1738 734 -1736
rect 733 -1744 734 -1742
rect 740 -1738 741 -1736
rect 737 -1744 738 -1742
rect 740 -1744 741 -1742
rect 744 -1738 745 -1736
rect 744 -1744 745 -1742
rect 751 -1738 752 -1736
rect 751 -1744 752 -1742
rect 758 -1738 759 -1736
rect 758 -1744 759 -1742
rect 765 -1738 766 -1736
rect 765 -1744 766 -1742
rect 772 -1738 773 -1736
rect 772 -1744 773 -1742
rect 779 -1738 780 -1736
rect 782 -1738 783 -1736
rect 779 -1744 780 -1742
rect 782 -1744 783 -1742
rect 789 -1738 790 -1736
rect 789 -1744 790 -1742
rect 793 -1738 794 -1736
rect 793 -1744 794 -1742
rect 800 -1738 801 -1736
rect 803 -1738 804 -1736
rect 800 -1744 801 -1742
rect 803 -1744 804 -1742
rect 807 -1738 808 -1736
rect 807 -1744 808 -1742
rect 810 -1744 811 -1742
rect 814 -1738 815 -1736
rect 814 -1744 815 -1742
rect 821 -1738 822 -1736
rect 821 -1744 822 -1742
rect 828 -1738 829 -1736
rect 828 -1744 829 -1742
rect 831 -1744 832 -1742
rect 835 -1738 836 -1736
rect 835 -1744 836 -1742
rect 842 -1738 843 -1736
rect 842 -1744 843 -1742
rect 849 -1738 850 -1736
rect 849 -1744 850 -1742
rect 856 -1738 857 -1736
rect 856 -1744 857 -1742
rect 863 -1738 864 -1736
rect 863 -1744 864 -1742
rect 870 -1738 871 -1736
rect 873 -1738 874 -1736
rect 870 -1744 871 -1742
rect 877 -1738 878 -1736
rect 877 -1744 878 -1742
rect 884 -1738 885 -1736
rect 887 -1738 888 -1736
rect 887 -1744 888 -1742
rect 894 -1738 895 -1736
rect 891 -1744 892 -1742
rect 894 -1744 895 -1742
rect 898 -1738 899 -1736
rect 898 -1744 899 -1742
rect 905 -1738 906 -1736
rect 905 -1744 906 -1742
rect 915 -1738 916 -1736
rect 912 -1744 913 -1742
rect 915 -1744 916 -1742
rect 919 -1738 920 -1736
rect 922 -1738 923 -1736
rect 919 -1744 920 -1742
rect 922 -1744 923 -1742
rect 926 -1738 927 -1736
rect 929 -1738 930 -1736
rect 926 -1744 927 -1742
rect 929 -1744 930 -1742
rect 933 -1738 934 -1736
rect 933 -1744 934 -1742
rect 940 -1738 941 -1736
rect 940 -1744 941 -1742
rect 947 -1738 948 -1736
rect 947 -1744 948 -1742
rect 954 -1738 955 -1736
rect 954 -1744 955 -1742
rect 961 -1738 962 -1736
rect 961 -1744 962 -1742
rect 968 -1738 969 -1736
rect 968 -1744 969 -1742
rect 975 -1738 976 -1736
rect 978 -1738 979 -1736
rect 978 -1744 979 -1742
rect 982 -1738 983 -1736
rect 982 -1744 983 -1742
rect 989 -1738 990 -1736
rect 992 -1738 993 -1736
rect 989 -1744 990 -1742
rect 996 -1738 997 -1736
rect 996 -1744 997 -1742
rect 1003 -1738 1004 -1736
rect 1003 -1744 1004 -1742
rect 1010 -1738 1011 -1736
rect 1010 -1744 1011 -1742
rect 1017 -1738 1018 -1736
rect 1017 -1744 1018 -1742
rect 1024 -1738 1025 -1736
rect 1024 -1744 1025 -1742
rect 1031 -1738 1032 -1736
rect 1031 -1744 1032 -1742
rect 1038 -1738 1039 -1736
rect 1038 -1744 1039 -1742
rect 1045 -1738 1046 -1736
rect 1045 -1744 1046 -1742
rect 1052 -1738 1053 -1736
rect 1052 -1744 1053 -1742
rect 1059 -1738 1060 -1736
rect 1059 -1744 1060 -1742
rect 1066 -1738 1067 -1736
rect 1066 -1744 1067 -1742
rect 1069 -1744 1070 -1742
rect 1073 -1738 1074 -1736
rect 1073 -1744 1074 -1742
rect 1080 -1738 1081 -1736
rect 1080 -1744 1081 -1742
rect 1087 -1738 1088 -1736
rect 1087 -1744 1088 -1742
rect 1094 -1738 1095 -1736
rect 1094 -1744 1095 -1742
rect 1101 -1738 1102 -1736
rect 1101 -1744 1102 -1742
rect 1108 -1738 1109 -1736
rect 1108 -1744 1109 -1742
rect 1115 -1738 1116 -1736
rect 1118 -1738 1119 -1736
rect 1115 -1744 1116 -1742
rect 1122 -1738 1123 -1736
rect 1122 -1744 1123 -1742
rect 1129 -1738 1130 -1736
rect 1129 -1744 1130 -1742
rect 1136 -1738 1137 -1736
rect 1136 -1744 1137 -1742
rect 1143 -1738 1144 -1736
rect 1143 -1744 1144 -1742
rect 1150 -1738 1151 -1736
rect 1150 -1744 1151 -1742
rect 1157 -1738 1158 -1736
rect 1157 -1744 1158 -1742
rect 1164 -1738 1165 -1736
rect 1164 -1744 1165 -1742
rect 1171 -1738 1172 -1736
rect 1171 -1744 1172 -1742
rect 1178 -1738 1179 -1736
rect 1178 -1744 1179 -1742
rect 1185 -1738 1186 -1736
rect 1185 -1744 1186 -1742
rect 1192 -1738 1193 -1736
rect 1192 -1744 1193 -1742
rect 1199 -1738 1200 -1736
rect 1199 -1744 1200 -1742
rect 1206 -1738 1207 -1736
rect 1206 -1744 1207 -1742
rect 1213 -1738 1214 -1736
rect 1213 -1744 1214 -1742
rect 1220 -1738 1221 -1736
rect 1220 -1744 1221 -1742
rect 1227 -1738 1228 -1736
rect 1227 -1744 1228 -1742
rect 1234 -1738 1235 -1736
rect 1234 -1744 1235 -1742
rect 1241 -1738 1242 -1736
rect 1241 -1744 1242 -1742
rect 1251 -1738 1252 -1736
rect 1248 -1744 1249 -1742
rect 1251 -1744 1252 -1742
rect 1255 -1738 1256 -1736
rect 1255 -1744 1256 -1742
rect 1262 -1738 1263 -1736
rect 1262 -1744 1263 -1742
rect 1269 -1738 1270 -1736
rect 1269 -1744 1270 -1742
rect 1276 -1738 1277 -1736
rect 1276 -1744 1277 -1742
rect 1283 -1738 1284 -1736
rect 1283 -1744 1284 -1742
rect 1290 -1738 1291 -1736
rect 1290 -1744 1291 -1742
rect 1297 -1738 1298 -1736
rect 1297 -1744 1298 -1742
rect 1304 -1738 1305 -1736
rect 1304 -1744 1305 -1742
rect 1311 -1738 1312 -1736
rect 1311 -1744 1312 -1742
rect 1318 -1738 1319 -1736
rect 1318 -1744 1319 -1742
rect 1325 -1738 1326 -1736
rect 1325 -1744 1326 -1742
rect 1332 -1738 1333 -1736
rect 1332 -1744 1333 -1742
rect 1339 -1738 1340 -1736
rect 1339 -1744 1340 -1742
rect 1346 -1738 1347 -1736
rect 1346 -1744 1347 -1742
rect 1353 -1738 1354 -1736
rect 1353 -1744 1354 -1742
rect 1360 -1738 1361 -1736
rect 1360 -1744 1361 -1742
rect 1367 -1738 1368 -1736
rect 1367 -1744 1368 -1742
rect 1374 -1738 1375 -1736
rect 1374 -1744 1375 -1742
rect 1381 -1738 1382 -1736
rect 1384 -1738 1385 -1736
rect 1381 -1744 1382 -1742
rect 1388 -1738 1389 -1736
rect 1388 -1744 1389 -1742
rect 1395 -1738 1396 -1736
rect 1395 -1744 1396 -1742
rect 1402 -1738 1403 -1736
rect 1402 -1744 1403 -1742
rect 1409 -1738 1410 -1736
rect 1409 -1744 1410 -1742
rect 1416 -1738 1417 -1736
rect 1416 -1744 1417 -1742
rect 1423 -1738 1424 -1736
rect 1423 -1744 1424 -1742
rect 1430 -1738 1431 -1736
rect 1430 -1744 1431 -1742
rect 1437 -1738 1438 -1736
rect 1437 -1744 1438 -1742
rect 1444 -1738 1445 -1736
rect 1444 -1744 1445 -1742
rect 1451 -1738 1452 -1736
rect 1451 -1744 1452 -1742
rect 1458 -1738 1459 -1736
rect 1458 -1744 1459 -1742
rect 1465 -1738 1466 -1736
rect 1465 -1744 1466 -1742
rect 1472 -1738 1473 -1736
rect 1472 -1744 1473 -1742
rect 1479 -1738 1480 -1736
rect 1479 -1744 1480 -1742
rect 1486 -1738 1487 -1736
rect 1486 -1744 1487 -1742
rect 1493 -1738 1494 -1736
rect 1493 -1744 1494 -1742
rect 1500 -1738 1501 -1736
rect 1500 -1744 1501 -1742
rect 1507 -1738 1508 -1736
rect 1507 -1744 1508 -1742
rect 1514 -1738 1515 -1736
rect 1514 -1744 1515 -1742
rect 1521 -1738 1522 -1736
rect 1521 -1744 1522 -1742
rect 1528 -1738 1529 -1736
rect 1528 -1744 1529 -1742
rect 1535 -1738 1536 -1736
rect 1535 -1744 1536 -1742
rect 1542 -1738 1543 -1736
rect 1542 -1744 1543 -1742
rect 1549 -1738 1550 -1736
rect 1549 -1744 1550 -1742
rect 1556 -1738 1557 -1736
rect 1556 -1744 1557 -1742
rect 1563 -1738 1564 -1736
rect 1563 -1744 1564 -1742
rect 1570 -1738 1571 -1736
rect 1570 -1744 1571 -1742
rect 1577 -1738 1578 -1736
rect 1577 -1744 1578 -1742
rect 1584 -1738 1585 -1736
rect 1584 -1744 1585 -1742
rect 1591 -1738 1592 -1736
rect 1591 -1744 1592 -1742
rect 1598 -1738 1599 -1736
rect 1598 -1744 1599 -1742
rect 1605 -1738 1606 -1736
rect 1605 -1744 1606 -1742
rect 1612 -1738 1613 -1736
rect 1612 -1744 1613 -1742
rect 1619 -1738 1620 -1736
rect 1619 -1744 1620 -1742
rect 1626 -1738 1627 -1736
rect 1626 -1744 1627 -1742
rect 1633 -1738 1634 -1736
rect 1633 -1744 1634 -1742
rect 1640 -1738 1641 -1736
rect 1640 -1744 1641 -1742
rect 1647 -1738 1648 -1736
rect 1647 -1744 1648 -1742
rect 1654 -1738 1655 -1736
rect 1654 -1744 1655 -1742
rect 1661 -1738 1662 -1736
rect 1661 -1744 1662 -1742
rect 1668 -1738 1669 -1736
rect 1668 -1744 1669 -1742
rect 1675 -1738 1676 -1736
rect 1675 -1744 1676 -1742
rect 1682 -1738 1683 -1736
rect 1682 -1744 1683 -1742
rect 1689 -1738 1690 -1736
rect 1689 -1744 1690 -1742
rect 1696 -1738 1697 -1736
rect 1696 -1744 1697 -1742
rect 1703 -1738 1704 -1736
rect 1703 -1744 1704 -1742
rect 1710 -1738 1711 -1736
rect 1710 -1744 1711 -1742
rect 1717 -1738 1718 -1736
rect 1717 -1744 1718 -1742
rect 1724 -1738 1725 -1736
rect 1724 -1744 1725 -1742
rect 1731 -1738 1732 -1736
rect 1731 -1744 1732 -1742
rect 1738 -1738 1739 -1736
rect 1738 -1744 1739 -1742
rect 1748 -1738 1749 -1736
rect 1745 -1744 1746 -1742
rect 1748 -1744 1749 -1742
rect 1752 -1738 1753 -1736
rect 1752 -1744 1753 -1742
rect 1759 -1738 1760 -1736
rect 1759 -1744 1760 -1742
rect 1766 -1738 1767 -1736
rect 1766 -1744 1767 -1742
rect 1773 -1738 1774 -1736
rect 1773 -1744 1774 -1742
rect 1780 -1738 1781 -1736
rect 1780 -1744 1781 -1742
rect 30 -1885 31 -1883
rect 30 -1891 31 -1889
rect 37 -1885 38 -1883
rect 37 -1891 38 -1889
rect 44 -1885 45 -1883
rect 44 -1891 45 -1889
rect 51 -1885 52 -1883
rect 51 -1891 52 -1889
rect 58 -1885 59 -1883
rect 58 -1891 59 -1889
rect 65 -1885 66 -1883
rect 65 -1891 66 -1889
rect 72 -1885 73 -1883
rect 72 -1891 73 -1889
rect 79 -1885 80 -1883
rect 79 -1891 80 -1889
rect 86 -1885 87 -1883
rect 86 -1891 87 -1889
rect 93 -1885 94 -1883
rect 93 -1891 94 -1889
rect 100 -1885 101 -1883
rect 100 -1891 101 -1889
rect 107 -1885 108 -1883
rect 110 -1885 111 -1883
rect 107 -1891 108 -1889
rect 110 -1891 111 -1889
rect 114 -1885 115 -1883
rect 114 -1891 115 -1889
rect 121 -1885 122 -1883
rect 121 -1891 122 -1889
rect 128 -1885 129 -1883
rect 128 -1891 129 -1889
rect 135 -1885 136 -1883
rect 135 -1891 136 -1889
rect 142 -1885 143 -1883
rect 142 -1891 143 -1889
rect 149 -1885 150 -1883
rect 149 -1891 150 -1889
rect 156 -1885 157 -1883
rect 159 -1885 160 -1883
rect 156 -1891 157 -1889
rect 159 -1891 160 -1889
rect 163 -1885 164 -1883
rect 163 -1891 164 -1889
rect 170 -1885 171 -1883
rect 170 -1891 171 -1889
rect 177 -1885 178 -1883
rect 180 -1885 181 -1883
rect 177 -1891 178 -1889
rect 180 -1891 181 -1889
rect 184 -1885 185 -1883
rect 184 -1891 185 -1889
rect 191 -1885 192 -1883
rect 191 -1891 192 -1889
rect 198 -1885 199 -1883
rect 198 -1891 199 -1889
rect 205 -1885 206 -1883
rect 208 -1885 209 -1883
rect 208 -1891 209 -1889
rect 212 -1885 213 -1883
rect 212 -1891 213 -1889
rect 219 -1885 220 -1883
rect 219 -1891 220 -1889
rect 226 -1885 227 -1883
rect 226 -1891 227 -1889
rect 233 -1885 234 -1883
rect 233 -1891 234 -1889
rect 240 -1885 241 -1883
rect 240 -1891 241 -1889
rect 247 -1885 248 -1883
rect 250 -1885 251 -1883
rect 247 -1891 248 -1889
rect 250 -1891 251 -1889
rect 254 -1885 255 -1883
rect 254 -1891 255 -1889
rect 264 -1885 265 -1883
rect 264 -1891 265 -1889
rect 268 -1885 269 -1883
rect 268 -1891 269 -1889
rect 275 -1885 276 -1883
rect 275 -1891 276 -1889
rect 282 -1885 283 -1883
rect 282 -1891 283 -1889
rect 289 -1885 290 -1883
rect 289 -1891 290 -1889
rect 296 -1885 297 -1883
rect 296 -1891 297 -1889
rect 303 -1885 304 -1883
rect 303 -1891 304 -1889
rect 310 -1885 311 -1883
rect 310 -1891 311 -1889
rect 317 -1885 318 -1883
rect 317 -1891 318 -1889
rect 324 -1885 325 -1883
rect 324 -1891 325 -1889
rect 331 -1885 332 -1883
rect 331 -1891 332 -1889
rect 338 -1885 339 -1883
rect 341 -1885 342 -1883
rect 341 -1891 342 -1889
rect 345 -1885 346 -1883
rect 345 -1891 346 -1889
rect 352 -1885 353 -1883
rect 352 -1891 353 -1889
rect 359 -1885 360 -1883
rect 359 -1891 360 -1889
rect 366 -1885 367 -1883
rect 366 -1891 367 -1889
rect 373 -1885 374 -1883
rect 373 -1891 374 -1889
rect 380 -1885 381 -1883
rect 380 -1891 381 -1889
rect 387 -1885 388 -1883
rect 387 -1891 388 -1889
rect 394 -1885 395 -1883
rect 394 -1891 395 -1889
rect 401 -1885 402 -1883
rect 401 -1891 402 -1889
rect 408 -1885 409 -1883
rect 408 -1891 409 -1889
rect 415 -1885 416 -1883
rect 415 -1891 416 -1889
rect 422 -1885 423 -1883
rect 422 -1891 423 -1889
rect 429 -1885 430 -1883
rect 429 -1891 430 -1889
rect 436 -1885 437 -1883
rect 436 -1891 437 -1889
rect 443 -1885 444 -1883
rect 446 -1885 447 -1883
rect 443 -1891 444 -1889
rect 446 -1891 447 -1889
rect 450 -1885 451 -1883
rect 450 -1891 451 -1889
rect 457 -1885 458 -1883
rect 457 -1891 458 -1889
rect 464 -1885 465 -1883
rect 467 -1885 468 -1883
rect 464 -1891 465 -1889
rect 467 -1891 468 -1889
rect 471 -1885 472 -1883
rect 474 -1885 475 -1883
rect 471 -1891 472 -1889
rect 474 -1891 475 -1889
rect 478 -1885 479 -1883
rect 478 -1891 479 -1889
rect 485 -1885 486 -1883
rect 492 -1885 493 -1883
rect 492 -1891 493 -1889
rect 502 -1885 503 -1883
rect 506 -1885 507 -1883
rect 506 -1891 507 -1889
rect 513 -1885 514 -1883
rect 513 -1891 514 -1889
rect 520 -1885 521 -1883
rect 520 -1891 521 -1889
rect 527 -1885 528 -1883
rect 527 -1891 528 -1889
rect 530 -1891 531 -1889
rect 534 -1885 535 -1883
rect 534 -1891 535 -1889
rect 541 -1885 542 -1883
rect 541 -1891 542 -1889
rect 548 -1885 549 -1883
rect 548 -1891 549 -1889
rect 555 -1885 556 -1883
rect 555 -1891 556 -1889
rect 562 -1885 563 -1883
rect 562 -1891 563 -1889
rect 569 -1885 570 -1883
rect 569 -1891 570 -1889
rect 572 -1891 573 -1889
rect 576 -1885 577 -1883
rect 576 -1891 577 -1889
rect 583 -1885 584 -1883
rect 583 -1891 584 -1889
rect 590 -1885 591 -1883
rect 590 -1891 591 -1889
rect 597 -1885 598 -1883
rect 597 -1891 598 -1889
rect 604 -1885 605 -1883
rect 604 -1891 605 -1889
rect 611 -1885 612 -1883
rect 611 -1891 612 -1889
rect 618 -1885 619 -1883
rect 618 -1891 619 -1889
rect 625 -1885 626 -1883
rect 625 -1891 626 -1889
rect 632 -1885 633 -1883
rect 632 -1891 633 -1889
rect 639 -1885 640 -1883
rect 639 -1891 640 -1889
rect 649 -1885 650 -1883
rect 646 -1891 647 -1889
rect 649 -1891 650 -1889
rect 653 -1885 654 -1883
rect 656 -1885 657 -1883
rect 653 -1891 654 -1889
rect 656 -1891 657 -1889
rect 660 -1885 661 -1883
rect 660 -1891 661 -1889
rect 667 -1885 668 -1883
rect 667 -1891 668 -1889
rect 674 -1885 675 -1883
rect 674 -1891 675 -1889
rect 681 -1885 682 -1883
rect 681 -1891 682 -1889
rect 688 -1885 689 -1883
rect 688 -1891 689 -1889
rect 695 -1885 696 -1883
rect 695 -1891 696 -1889
rect 702 -1885 703 -1883
rect 702 -1891 703 -1889
rect 709 -1885 710 -1883
rect 709 -1891 710 -1889
rect 716 -1885 717 -1883
rect 716 -1891 717 -1889
rect 723 -1885 724 -1883
rect 723 -1891 724 -1889
rect 730 -1885 731 -1883
rect 730 -1891 731 -1889
rect 737 -1885 738 -1883
rect 737 -1891 738 -1889
rect 744 -1885 745 -1883
rect 744 -1891 745 -1889
rect 751 -1885 752 -1883
rect 751 -1891 752 -1889
rect 758 -1885 759 -1883
rect 758 -1891 759 -1889
rect 765 -1885 766 -1883
rect 765 -1891 766 -1889
rect 772 -1885 773 -1883
rect 772 -1891 773 -1889
rect 779 -1885 780 -1883
rect 779 -1891 780 -1889
rect 786 -1885 787 -1883
rect 786 -1891 787 -1889
rect 793 -1885 794 -1883
rect 793 -1891 794 -1889
rect 800 -1885 801 -1883
rect 800 -1891 801 -1889
rect 810 -1885 811 -1883
rect 807 -1891 808 -1889
rect 810 -1891 811 -1889
rect 814 -1885 815 -1883
rect 814 -1891 815 -1889
rect 821 -1885 822 -1883
rect 824 -1885 825 -1883
rect 821 -1891 822 -1889
rect 824 -1891 825 -1889
rect 828 -1885 829 -1883
rect 831 -1885 832 -1883
rect 831 -1891 832 -1889
rect 835 -1885 836 -1883
rect 838 -1891 839 -1889
rect 842 -1885 843 -1883
rect 842 -1891 843 -1889
rect 849 -1885 850 -1883
rect 849 -1891 850 -1889
rect 856 -1885 857 -1883
rect 856 -1891 857 -1889
rect 863 -1885 864 -1883
rect 866 -1885 867 -1883
rect 866 -1891 867 -1889
rect 870 -1885 871 -1883
rect 870 -1891 871 -1889
rect 877 -1885 878 -1883
rect 877 -1891 878 -1889
rect 884 -1885 885 -1883
rect 884 -1891 885 -1889
rect 891 -1885 892 -1883
rect 891 -1891 892 -1889
rect 898 -1885 899 -1883
rect 898 -1891 899 -1889
rect 905 -1885 906 -1883
rect 905 -1891 906 -1889
rect 908 -1891 909 -1889
rect 912 -1885 913 -1883
rect 912 -1891 913 -1889
rect 919 -1885 920 -1883
rect 919 -1891 920 -1889
rect 926 -1885 927 -1883
rect 929 -1885 930 -1883
rect 926 -1891 927 -1889
rect 929 -1891 930 -1889
rect 933 -1885 934 -1883
rect 936 -1885 937 -1883
rect 936 -1891 937 -1889
rect 940 -1885 941 -1883
rect 940 -1891 941 -1889
rect 947 -1885 948 -1883
rect 947 -1891 948 -1889
rect 957 -1891 958 -1889
rect 961 -1885 962 -1883
rect 961 -1891 962 -1889
rect 968 -1885 969 -1883
rect 968 -1891 969 -1889
rect 975 -1885 976 -1883
rect 975 -1891 976 -1889
rect 982 -1885 983 -1883
rect 985 -1885 986 -1883
rect 985 -1891 986 -1889
rect 989 -1885 990 -1883
rect 989 -1891 990 -1889
rect 996 -1885 997 -1883
rect 996 -1891 997 -1889
rect 1003 -1885 1004 -1883
rect 1003 -1891 1004 -1889
rect 1010 -1885 1011 -1883
rect 1010 -1891 1011 -1889
rect 1017 -1885 1018 -1883
rect 1017 -1891 1018 -1889
rect 1020 -1891 1021 -1889
rect 1024 -1885 1025 -1883
rect 1027 -1885 1028 -1883
rect 1024 -1891 1025 -1889
rect 1027 -1891 1028 -1889
rect 1031 -1885 1032 -1883
rect 1031 -1891 1032 -1889
rect 1038 -1885 1039 -1883
rect 1041 -1885 1042 -1883
rect 1038 -1891 1039 -1889
rect 1045 -1885 1046 -1883
rect 1048 -1885 1049 -1883
rect 1045 -1891 1046 -1889
rect 1048 -1891 1049 -1889
rect 1052 -1885 1053 -1883
rect 1052 -1891 1053 -1889
rect 1059 -1885 1060 -1883
rect 1059 -1891 1060 -1889
rect 1066 -1885 1067 -1883
rect 1066 -1891 1067 -1889
rect 1073 -1885 1074 -1883
rect 1073 -1891 1074 -1889
rect 1080 -1885 1081 -1883
rect 1080 -1891 1081 -1889
rect 1087 -1885 1088 -1883
rect 1087 -1891 1088 -1889
rect 1094 -1885 1095 -1883
rect 1094 -1891 1095 -1889
rect 1101 -1885 1102 -1883
rect 1101 -1891 1102 -1889
rect 1108 -1885 1109 -1883
rect 1111 -1885 1112 -1883
rect 1108 -1891 1109 -1889
rect 1115 -1885 1116 -1883
rect 1115 -1891 1116 -1889
rect 1122 -1885 1123 -1883
rect 1122 -1891 1123 -1889
rect 1129 -1885 1130 -1883
rect 1129 -1891 1130 -1889
rect 1136 -1885 1137 -1883
rect 1136 -1891 1137 -1889
rect 1143 -1885 1144 -1883
rect 1143 -1891 1144 -1889
rect 1150 -1885 1151 -1883
rect 1153 -1885 1154 -1883
rect 1150 -1891 1151 -1889
rect 1153 -1891 1154 -1889
rect 1157 -1885 1158 -1883
rect 1160 -1885 1161 -1883
rect 1157 -1891 1158 -1889
rect 1160 -1891 1161 -1889
rect 1164 -1885 1165 -1883
rect 1164 -1891 1165 -1889
rect 1171 -1885 1172 -1883
rect 1171 -1891 1172 -1889
rect 1178 -1885 1179 -1883
rect 1178 -1891 1179 -1889
rect 1185 -1885 1186 -1883
rect 1185 -1891 1186 -1889
rect 1192 -1885 1193 -1883
rect 1192 -1891 1193 -1889
rect 1199 -1885 1200 -1883
rect 1199 -1891 1200 -1889
rect 1206 -1885 1207 -1883
rect 1206 -1891 1207 -1889
rect 1213 -1885 1214 -1883
rect 1213 -1891 1214 -1889
rect 1220 -1885 1221 -1883
rect 1220 -1891 1221 -1889
rect 1227 -1885 1228 -1883
rect 1227 -1891 1228 -1889
rect 1234 -1885 1235 -1883
rect 1234 -1891 1235 -1889
rect 1241 -1885 1242 -1883
rect 1241 -1891 1242 -1889
rect 1248 -1885 1249 -1883
rect 1248 -1891 1249 -1889
rect 1255 -1885 1256 -1883
rect 1255 -1891 1256 -1889
rect 1262 -1885 1263 -1883
rect 1262 -1891 1263 -1889
rect 1269 -1885 1270 -1883
rect 1269 -1891 1270 -1889
rect 1276 -1885 1277 -1883
rect 1279 -1885 1280 -1883
rect 1276 -1891 1277 -1889
rect 1279 -1891 1280 -1889
rect 1283 -1885 1284 -1883
rect 1283 -1891 1284 -1889
rect 1290 -1885 1291 -1883
rect 1290 -1891 1291 -1889
rect 1297 -1885 1298 -1883
rect 1297 -1891 1298 -1889
rect 1304 -1885 1305 -1883
rect 1304 -1891 1305 -1889
rect 1311 -1891 1312 -1889
rect 1314 -1891 1315 -1889
rect 1318 -1885 1319 -1883
rect 1318 -1891 1319 -1889
rect 1325 -1885 1326 -1883
rect 1325 -1891 1326 -1889
rect 1332 -1885 1333 -1883
rect 1332 -1891 1333 -1889
rect 1339 -1885 1340 -1883
rect 1339 -1891 1340 -1889
rect 1346 -1885 1347 -1883
rect 1346 -1891 1347 -1889
rect 1353 -1885 1354 -1883
rect 1353 -1891 1354 -1889
rect 1360 -1885 1361 -1883
rect 1360 -1891 1361 -1889
rect 1367 -1885 1368 -1883
rect 1367 -1891 1368 -1889
rect 1374 -1885 1375 -1883
rect 1374 -1891 1375 -1889
rect 1381 -1885 1382 -1883
rect 1381 -1891 1382 -1889
rect 1384 -1891 1385 -1889
rect 1388 -1885 1389 -1883
rect 1388 -1891 1389 -1889
rect 1395 -1885 1396 -1883
rect 1395 -1891 1396 -1889
rect 1402 -1885 1403 -1883
rect 1402 -1891 1403 -1889
rect 1409 -1885 1410 -1883
rect 1409 -1891 1410 -1889
rect 1416 -1885 1417 -1883
rect 1416 -1891 1417 -1889
rect 1423 -1885 1424 -1883
rect 1423 -1891 1424 -1889
rect 1430 -1885 1431 -1883
rect 1430 -1891 1431 -1889
rect 1437 -1885 1438 -1883
rect 1437 -1891 1438 -1889
rect 1444 -1885 1445 -1883
rect 1444 -1891 1445 -1889
rect 1451 -1885 1452 -1883
rect 1451 -1891 1452 -1889
rect 1458 -1885 1459 -1883
rect 1458 -1891 1459 -1889
rect 1465 -1885 1466 -1883
rect 1465 -1891 1466 -1889
rect 1472 -1885 1473 -1883
rect 1472 -1891 1473 -1889
rect 1479 -1885 1480 -1883
rect 1479 -1891 1480 -1889
rect 1486 -1885 1487 -1883
rect 1486 -1891 1487 -1889
rect 1493 -1885 1494 -1883
rect 1493 -1891 1494 -1889
rect 1500 -1885 1501 -1883
rect 1500 -1891 1501 -1889
rect 1507 -1885 1508 -1883
rect 1507 -1891 1508 -1889
rect 1514 -1885 1515 -1883
rect 1514 -1891 1515 -1889
rect 1521 -1885 1522 -1883
rect 1521 -1891 1522 -1889
rect 1528 -1885 1529 -1883
rect 1528 -1891 1529 -1889
rect 1535 -1885 1536 -1883
rect 1535 -1891 1536 -1889
rect 1542 -1885 1543 -1883
rect 1542 -1891 1543 -1889
rect 1549 -1885 1550 -1883
rect 1549 -1891 1550 -1889
rect 1556 -1885 1557 -1883
rect 1556 -1891 1557 -1889
rect 1563 -1885 1564 -1883
rect 1563 -1891 1564 -1889
rect 1570 -1885 1571 -1883
rect 1570 -1891 1571 -1889
rect 1577 -1885 1578 -1883
rect 1577 -1891 1578 -1889
rect 1584 -1885 1585 -1883
rect 1584 -1891 1585 -1889
rect 1591 -1885 1592 -1883
rect 1591 -1891 1592 -1889
rect 1598 -1885 1599 -1883
rect 1598 -1891 1599 -1889
rect 1605 -1885 1606 -1883
rect 1605 -1891 1606 -1889
rect 1612 -1885 1613 -1883
rect 1612 -1891 1613 -1889
rect 1619 -1885 1620 -1883
rect 1619 -1891 1620 -1889
rect 1626 -1885 1627 -1883
rect 1626 -1891 1627 -1889
rect 1633 -1885 1634 -1883
rect 1633 -1891 1634 -1889
rect 1640 -1885 1641 -1883
rect 1640 -1891 1641 -1889
rect 1647 -1885 1648 -1883
rect 1647 -1891 1648 -1889
rect 1654 -1885 1655 -1883
rect 1654 -1891 1655 -1889
rect 1661 -1885 1662 -1883
rect 1661 -1891 1662 -1889
rect 1668 -1885 1669 -1883
rect 1668 -1891 1669 -1889
rect 1675 -1885 1676 -1883
rect 1675 -1891 1676 -1889
rect 1682 -1885 1683 -1883
rect 1682 -1891 1683 -1889
rect 1689 -1885 1690 -1883
rect 1689 -1891 1690 -1889
rect 1696 -1885 1697 -1883
rect 1696 -1891 1697 -1889
rect 1703 -1885 1704 -1883
rect 1703 -1891 1704 -1889
rect 1710 -1885 1711 -1883
rect 1710 -1891 1711 -1889
rect 1717 -1885 1718 -1883
rect 1717 -1891 1718 -1889
rect 1724 -1885 1725 -1883
rect 1724 -1891 1725 -1889
rect 1731 -1885 1732 -1883
rect 1731 -1891 1732 -1889
rect 1738 -1885 1739 -1883
rect 1738 -1891 1739 -1889
rect 1745 -1885 1746 -1883
rect 1745 -1891 1746 -1889
rect 1752 -1885 1753 -1883
rect 1752 -1891 1753 -1889
rect 1759 -1885 1760 -1883
rect 1759 -1891 1760 -1889
rect 1766 -1885 1767 -1883
rect 1766 -1891 1767 -1889
rect 1773 -1885 1774 -1883
rect 1776 -1885 1777 -1883
rect 1773 -1891 1774 -1889
rect 1776 -1891 1777 -1889
rect 1780 -1885 1781 -1883
rect 1780 -1891 1781 -1889
rect 1787 -1885 1788 -1883
rect 1787 -1891 1788 -1889
rect 1794 -1885 1795 -1883
rect 1794 -1891 1795 -1889
rect 1801 -1885 1802 -1883
rect 1804 -1885 1805 -1883
rect 1801 -1891 1802 -1889
rect 1804 -1891 1805 -1889
rect 1808 -1885 1809 -1883
rect 1808 -1891 1809 -1889
rect 1815 -1885 1816 -1883
rect 1815 -1891 1816 -1889
rect 30 -2018 31 -2016
rect 30 -2024 31 -2022
rect 44 -2018 45 -2016
rect 44 -2024 45 -2022
rect 51 -2018 52 -2016
rect 51 -2024 52 -2022
rect 58 -2018 59 -2016
rect 58 -2024 59 -2022
rect 65 -2018 66 -2016
rect 68 -2018 69 -2016
rect 65 -2024 66 -2022
rect 72 -2018 73 -2016
rect 72 -2024 73 -2022
rect 79 -2018 80 -2016
rect 79 -2024 80 -2022
rect 86 -2018 87 -2016
rect 89 -2018 90 -2016
rect 86 -2024 87 -2022
rect 93 -2018 94 -2016
rect 93 -2024 94 -2022
rect 100 -2018 101 -2016
rect 103 -2018 104 -2016
rect 100 -2024 101 -2022
rect 103 -2024 104 -2022
rect 107 -2018 108 -2016
rect 110 -2018 111 -2016
rect 107 -2024 108 -2022
rect 114 -2018 115 -2016
rect 114 -2024 115 -2022
rect 121 -2018 122 -2016
rect 124 -2018 125 -2016
rect 121 -2024 122 -2022
rect 124 -2024 125 -2022
rect 131 -2018 132 -2016
rect 128 -2024 129 -2022
rect 131 -2024 132 -2022
rect 135 -2018 136 -2016
rect 135 -2024 136 -2022
rect 142 -2018 143 -2016
rect 145 -2018 146 -2016
rect 142 -2024 143 -2022
rect 145 -2024 146 -2022
rect 149 -2018 150 -2016
rect 152 -2018 153 -2016
rect 152 -2024 153 -2022
rect 156 -2018 157 -2016
rect 156 -2024 157 -2022
rect 163 -2018 164 -2016
rect 163 -2024 164 -2022
rect 170 -2018 171 -2016
rect 170 -2024 171 -2022
rect 177 -2018 178 -2016
rect 180 -2018 181 -2016
rect 177 -2024 178 -2022
rect 180 -2024 181 -2022
rect 184 -2018 185 -2016
rect 184 -2024 185 -2022
rect 191 -2018 192 -2016
rect 191 -2024 192 -2022
rect 198 -2018 199 -2016
rect 198 -2024 199 -2022
rect 205 -2018 206 -2016
rect 205 -2024 206 -2022
rect 212 -2018 213 -2016
rect 215 -2018 216 -2016
rect 212 -2024 213 -2022
rect 219 -2018 220 -2016
rect 219 -2024 220 -2022
rect 222 -2024 223 -2022
rect 226 -2018 227 -2016
rect 226 -2024 227 -2022
rect 233 -2018 234 -2016
rect 233 -2024 234 -2022
rect 240 -2018 241 -2016
rect 240 -2024 241 -2022
rect 247 -2018 248 -2016
rect 247 -2024 248 -2022
rect 254 -2018 255 -2016
rect 254 -2024 255 -2022
rect 261 -2018 262 -2016
rect 261 -2024 262 -2022
rect 268 -2018 269 -2016
rect 268 -2024 269 -2022
rect 275 -2018 276 -2016
rect 275 -2024 276 -2022
rect 282 -2018 283 -2016
rect 282 -2024 283 -2022
rect 289 -2018 290 -2016
rect 289 -2024 290 -2022
rect 296 -2018 297 -2016
rect 296 -2024 297 -2022
rect 303 -2018 304 -2016
rect 303 -2024 304 -2022
rect 310 -2018 311 -2016
rect 310 -2024 311 -2022
rect 317 -2018 318 -2016
rect 317 -2024 318 -2022
rect 324 -2018 325 -2016
rect 324 -2024 325 -2022
rect 331 -2018 332 -2016
rect 334 -2018 335 -2016
rect 331 -2024 332 -2022
rect 338 -2018 339 -2016
rect 338 -2024 339 -2022
rect 345 -2018 346 -2016
rect 345 -2024 346 -2022
rect 352 -2018 353 -2016
rect 352 -2024 353 -2022
rect 359 -2018 360 -2016
rect 359 -2024 360 -2022
rect 366 -2018 367 -2016
rect 366 -2024 367 -2022
rect 373 -2018 374 -2016
rect 373 -2024 374 -2022
rect 380 -2018 381 -2016
rect 380 -2024 381 -2022
rect 387 -2024 388 -2022
rect 394 -2018 395 -2016
rect 394 -2024 395 -2022
rect 401 -2018 402 -2016
rect 401 -2024 402 -2022
rect 408 -2018 409 -2016
rect 408 -2024 409 -2022
rect 415 -2018 416 -2016
rect 415 -2024 416 -2022
rect 422 -2018 423 -2016
rect 422 -2024 423 -2022
rect 429 -2018 430 -2016
rect 429 -2024 430 -2022
rect 436 -2018 437 -2016
rect 436 -2024 437 -2022
rect 443 -2018 444 -2016
rect 443 -2024 444 -2022
rect 450 -2018 451 -2016
rect 450 -2024 451 -2022
rect 457 -2018 458 -2016
rect 460 -2018 461 -2016
rect 457 -2024 458 -2022
rect 460 -2024 461 -2022
rect 464 -2018 465 -2016
rect 464 -2024 465 -2022
rect 471 -2018 472 -2016
rect 471 -2024 472 -2022
rect 478 -2018 479 -2016
rect 478 -2024 479 -2022
rect 485 -2024 486 -2022
rect 492 -2018 493 -2016
rect 492 -2024 493 -2022
rect 499 -2018 500 -2016
rect 499 -2024 500 -2022
rect 506 -2018 507 -2016
rect 509 -2018 510 -2016
rect 509 -2024 510 -2022
rect 513 -2018 514 -2016
rect 513 -2024 514 -2022
rect 520 -2018 521 -2016
rect 520 -2024 521 -2022
rect 527 -2018 528 -2016
rect 527 -2024 528 -2022
rect 534 -2018 535 -2016
rect 541 -2018 542 -2016
rect 541 -2024 542 -2022
rect 548 -2018 549 -2016
rect 548 -2024 549 -2022
rect 555 -2018 556 -2016
rect 555 -2024 556 -2022
rect 562 -2018 563 -2016
rect 562 -2024 563 -2022
rect 569 -2018 570 -2016
rect 569 -2024 570 -2022
rect 572 -2024 573 -2022
rect 576 -2018 577 -2016
rect 576 -2024 577 -2022
rect 583 -2018 584 -2016
rect 583 -2024 584 -2022
rect 593 -2018 594 -2016
rect 593 -2024 594 -2022
rect 597 -2018 598 -2016
rect 597 -2024 598 -2022
rect 604 -2018 605 -2016
rect 604 -2024 605 -2022
rect 611 -2018 612 -2016
rect 611 -2024 612 -2022
rect 618 -2018 619 -2016
rect 618 -2024 619 -2022
rect 625 -2018 626 -2016
rect 628 -2018 629 -2016
rect 625 -2024 626 -2022
rect 628 -2024 629 -2022
rect 632 -2018 633 -2016
rect 632 -2024 633 -2022
rect 639 -2018 640 -2016
rect 639 -2024 640 -2022
rect 646 -2018 647 -2016
rect 646 -2024 647 -2022
rect 653 -2018 654 -2016
rect 653 -2024 654 -2022
rect 660 -2018 661 -2016
rect 660 -2024 661 -2022
rect 667 -2018 668 -2016
rect 667 -2024 668 -2022
rect 674 -2018 675 -2016
rect 674 -2024 675 -2022
rect 681 -2018 682 -2016
rect 681 -2024 682 -2022
rect 688 -2018 689 -2016
rect 688 -2024 689 -2022
rect 695 -2018 696 -2016
rect 695 -2024 696 -2022
rect 702 -2018 703 -2016
rect 702 -2024 703 -2022
rect 709 -2018 710 -2016
rect 709 -2024 710 -2022
rect 716 -2018 717 -2016
rect 719 -2018 720 -2016
rect 716 -2024 717 -2022
rect 719 -2024 720 -2022
rect 723 -2018 724 -2016
rect 723 -2024 724 -2022
rect 730 -2018 731 -2016
rect 730 -2024 731 -2022
rect 737 -2018 738 -2016
rect 737 -2024 738 -2022
rect 744 -2018 745 -2016
rect 744 -2024 745 -2022
rect 751 -2018 752 -2016
rect 751 -2024 752 -2022
rect 758 -2018 759 -2016
rect 761 -2018 762 -2016
rect 758 -2024 759 -2022
rect 761 -2024 762 -2022
rect 765 -2018 766 -2016
rect 765 -2024 766 -2022
rect 772 -2018 773 -2016
rect 772 -2024 773 -2022
rect 779 -2018 780 -2016
rect 779 -2024 780 -2022
rect 786 -2018 787 -2016
rect 786 -2024 787 -2022
rect 793 -2018 794 -2016
rect 796 -2018 797 -2016
rect 796 -2024 797 -2022
rect 800 -2018 801 -2016
rect 800 -2024 801 -2022
rect 807 -2018 808 -2016
rect 807 -2024 808 -2022
rect 814 -2018 815 -2016
rect 814 -2024 815 -2022
rect 821 -2018 822 -2016
rect 821 -2024 822 -2022
rect 828 -2018 829 -2016
rect 828 -2024 829 -2022
rect 835 -2018 836 -2016
rect 835 -2024 836 -2022
rect 842 -2018 843 -2016
rect 842 -2024 843 -2022
rect 849 -2018 850 -2016
rect 849 -2024 850 -2022
rect 856 -2018 857 -2016
rect 856 -2024 857 -2022
rect 863 -2018 864 -2016
rect 863 -2024 864 -2022
rect 870 -2018 871 -2016
rect 870 -2024 871 -2022
rect 877 -2018 878 -2016
rect 877 -2024 878 -2022
rect 884 -2018 885 -2016
rect 887 -2018 888 -2016
rect 884 -2024 885 -2022
rect 887 -2024 888 -2022
rect 891 -2018 892 -2016
rect 894 -2018 895 -2016
rect 891 -2024 892 -2022
rect 894 -2024 895 -2022
rect 898 -2018 899 -2016
rect 901 -2018 902 -2016
rect 901 -2024 902 -2022
rect 905 -2018 906 -2016
rect 905 -2024 906 -2022
rect 912 -2018 913 -2016
rect 912 -2024 913 -2022
rect 919 -2018 920 -2016
rect 922 -2018 923 -2016
rect 919 -2024 920 -2022
rect 922 -2024 923 -2022
rect 926 -2018 927 -2016
rect 926 -2024 927 -2022
rect 933 -2018 934 -2016
rect 933 -2024 934 -2022
rect 940 -2018 941 -2016
rect 940 -2024 941 -2022
rect 947 -2018 948 -2016
rect 947 -2024 948 -2022
rect 954 -2018 955 -2016
rect 954 -2024 955 -2022
rect 957 -2024 958 -2022
rect 961 -2018 962 -2016
rect 964 -2024 965 -2022
rect 968 -2018 969 -2016
rect 968 -2024 969 -2022
rect 975 -2018 976 -2016
rect 975 -2024 976 -2022
rect 982 -2018 983 -2016
rect 982 -2024 983 -2022
rect 989 -2018 990 -2016
rect 989 -2024 990 -2022
rect 992 -2024 993 -2022
rect 999 -2018 1000 -2016
rect 996 -2024 997 -2022
rect 999 -2024 1000 -2022
rect 1003 -2018 1004 -2016
rect 1003 -2024 1004 -2022
rect 1010 -2018 1011 -2016
rect 1010 -2024 1011 -2022
rect 1017 -2018 1018 -2016
rect 1017 -2024 1018 -2022
rect 1024 -2018 1025 -2016
rect 1024 -2024 1025 -2022
rect 1031 -2018 1032 -2016
rect 1031 -2024 1032 -2022
rect 1038 -2018 1039 -2016
rect 1041 -2018 1042 -2016
rect 1045 -2018 1046 -2016
rect 1045 -2024 1046 -2022
rect 1052 -2018 1053 -2016
rect 1052 -2024 1053 -2022
rect 1059 -2018 1060 -2016
rect 1059 -2024 1060 -2022
rect 1066 -2018 1067 -2016
rect 1066 -2024 1067 -2022
rect 1073 -2018 1074 -2016
rect 1073 -2024 1074 -2022
rect 1080 -2018 1081 -2016
rect 1080 -2024 1081 -2022
rect 1087 -2018 1088 -2016
rect 1087 -2024 1088 -2022
rect 1094 -2018 1095 -2016
rect 1094 -2024 1095 -2022
rect 1101 -2018 1102 -2016
rect 1101 -2024 1102 -2022
rect 1108 -2018 1109 -2016
rect 1111 -2018 1112 -2016
rect 1108 -2024 1109 -2022
rect 1115 -2018 1116 -2016
rect 1115 -2024 1116 -2022
rect 1122 -2018 1123 -2016
rect 1122 -2024 1123 -2022
rect 1129 -2018 1130 -2016
rect 1129 -2024 1130 -2022
rect 1136 -2018 1137 -2016
rect 1139 -2018 1140 -2016
rect 1139 -2024 1140 -2022
rect 1143 -2018 1144 -2016
rect 1143 -2024 1144 -2022
rect 1150 -2018 1151 -2016
rect 1150 -2024 1151 -2022
rect 1157 -2018 1158 -2016
rect 1157 -2024 1158 -2022
rect 1164 -2018 1165 -2016
rect 1164 -2024 1165 -2022
rect 1171 -2018 1172 -2016
rect 1171 -2024 1172 -2022
rect 1178 -2018 1179 -2016
rect 1178 -2024 1179 -2022
rect 1185 -2018 1186 -2016
rect 1185 -2024 1186 -2022
rect 1192 -2018 1193 -2016
rect 1195 -2024 1196 -2022
rect 1199 -2018 1200 -2016
rect 1199 -2024 1200 -2022
rect 1206 -2018 1207 -2016
rect 1206 -2024 1207 -2022
rect 1216 -2018 1217 -2016
rect 1213 -2024 1214 -2022
rect 1220 -2018 1221 -2016
rect 1220 -2024 1221 -2022
rect 1227 -2018 1228 -2016
rect 1227 -2024 1228 -2022
rect 1234 -2018 1235 -2016
rect 1234 -2024 1235 -2022
rect 1241 -2018 1242 -2016
rect 1241 -2024 1242 -2022
rect 1248 -2018 1249 -2016
rect 1248 -2024 1249 -2022
rect 1255 -2018 1256 -2016
rect 1255 -2024 1256 -2022
rect 1262 -2018 1263 -2016
rect 1262 -2024 1263 -2022
rect 1269 -2018 1270 -2016
rect 1269 -2024 1270 -2022
rect 1276 -2018 1277 -2016
rect 1276 -2024 1277 -2022
rect 1283 -2018 1284 -2016
rect 1283 -2024 1284 -2022
rect 1293 -2018 1294 -2016
rect 1290 -2024 1291 -2022
rect 1293 -2024 1294 -2022
rect 1297 -2018 1298 -2016
rect 1297 -2024 1298 -2022
rect 1304 -2018 1305 -2016
rect 1304 -2024 1305 -2022
rect 1311 -2018 1312 -2016
rect 1311 -2024 1312 -2022
rect 1318 -2018 1319 -2016
rect 1318 -2024 1319 -2022
rect 1325 -2018 1326 -2016
rect 1325 -2024 1326 -2022
rect 1332 -2018 1333 -2016
rect 1332 -2024 1333 -2022
rect 1339 -2018 1340 -2016
rect 1339 -2024 1340 -2022
rect 1346 -2018 1347 -2016
rect 1346 -2024 1347 -2022
rect 1353 -2018 1354 -2016
rect 1353 -2024 1354 -2022
rect 1360 -2018 1361 -2016
rect 1360 -2024 1361 -2022
rect 1367 -2018 1368 -2016
rect 1367 -2024 1368 -2022
rect 1374 -2018 1375 -2016
rect 1374 -2024 1375 -2022
rect 1381 -2018 1382 -2016
rect 1384 -2018 1385 -2016
rect 1381 -2024 1382 -2022
rect 1388 -2018 1389 -2016
rect 1388 -2024 1389 -2022
rect 1395 -2018 1396 -2016
rect 1395 -2024 1396 -2022
rect 1402 -2018 1403 -2016
rect 1402 -2024 1403 -2022
rect 1409 -2018 1410 -2016
rect 1409 -2024 1410 -2022
rect 1416 -2018 1417 -2016
rect 1416 -2024 1417 -2022
rect 1423 -2018 1424 -2016
rect 1423 -2024 1424 -2022
rect 1430 -2018 1431 -2016
rect 1430 -2024 1431 -2022
rect 1437 -2018 1438 -2016
rect 1437 -2024 1438 -2022
rect 1444 -2018 1445 -2016
rect 1444 -2024 1445 -2022
rect 1451 -2018 1452 -2016
rect 1451 -2024 1452 -2022
rect 1458 -2018 1459 -2016
rect 1458 -2024 1459 -2022
rect 1465 -2018 1466 -2016
rect 1465 -2024 1466 -2022
rect 1472 -2018 1473 -2016
rect 1472 -2024 1473 -2022
rect 1479 -2018 1480 -2016
rect 1479 -2024 1480 -2022
rect 1486 -2018 1487 -2016
rect 1486 -2024 1487 -2022
rect 1493 -2018 1494 -2016
rect 1493 -2024 1494 -2022
rect 1500 -2018 1501 -2016
rect 1500 -2024 1501 -2022
rect 1507 -2018 1508 -2016
rect 1507 -2024 1508 -2022
rect 1514 -2018 1515 -2016
rect 1514 -2024 1515 -2022
rect 1521 -2018 1522 -2016
rect 1521 -2024 1522 -2022
rect 1528 -2018 1529 -2016
rect 1528 -2024 1529 -2022
rect 1535 -2018 1536 -2016
rect 1535 -2024 1536 -2022
rect 1542 -2018 1543 -2016
rect 1542 -2024 1543 -2022
rect 1549 -2018 1550 -2016
rect 1549 -2024 1550 -2022
rect 1556 -2018 1557 -2016
rect 1556 -2024 1557 -2022
rect 1563 -2018 1564 -2016
rect 1563 -2024 1564 -2022
rect 1570 -2018 1571 -2016
rect 1570 -2024 1571 -2022
rect 1577 -2018 1578 -2016
rect 1577 -2024 1578 -2022
rect 1584 -2018 1585 -2016
rect 1584 -2024 1585 -2022
rect 1591 -2018 1592 -2016
rect 1591 -2024 1592 -2022
rect 1594 -2024 1595 -2022
rect 1598 -2018 1599 -2016
rect 1598 -2024 1599 -2022
rect 1605 -2018 1606 -2016
rect 1605 -2024 1606 -2022
rect 1612 -2018 1613 -2016
rect 1612 -2024 1613 -2022
rect 1619 -2018 1620 -2016
rect 1619 -2024 1620 -2022
rect 1626 -2018 1627 -2016
rect 1626 -2024 1627 -2022
rect 1633 -2018 1634 -2016
rect 1633 -2024 1634 -2022
rect 1640 -2018 1641 -2016
rect 1640 -2024 1641 -2022
rect 1647 -2018 1648 -2016
rect 1647 -2024 1648 -2022
rect 1654 -2018 1655 -2016
rect 1654 -2024 1655 -2022
rect 1661 -2018 1662 -2016
rect 1661 -2024 1662 -2022
rect 1668 -2018 1669 -2016
rect 1668 -2024 1669 -2022
rect 1675 -2018 1676 -2016
rect 1675 -2024 1676 -2022
rect 1682 -2018 1683 -2016
rect 1682 -2024 1683 -2022
rect 1689 -2018 1690 -2016
rect 1689 -2024 1690 -2022
rect 1696 -2018 1697 -2016
rect 1696 -2024 1697 -2022
rect 1703 -2018 1704 -2016
rect 1703 -2024 1704 -2022
rect 1710 -2018 1711 -2016
rect 1710 -2024 1711 -2022
rect 1717 -2018 1718 -2016
rect 1717 -2024 1718 -2022
rect 1724 -2018 1725 -2016
rect 1724 -2024 1725 -2022
rect 1731 -2018 1732 -2016
rect 1731 -2024 1732 -2022
rect 1738 -2018 1739 -2016
rect 1738 -2024 1739 -2022
rect 1745 -2024 1746 -2022
rect 1748 -2024 1749 -2022
rect 1752 -2018 1753 -2016
rect 1752 -2024 1753 -2022
rect 1759 -2018 1760 -2016
rect 1759 -2024 1760 -2022
rect 1766 -2018 1767 -2016
rect 1766 -2024 1767 -2022
rect 1773 -2018 1774 -2016
rect 1773 -2024 1774 -2022
rect 1780 -2018 1781 -2016
rect 1780 -2024 1781 -2022
rect 1787 -2018 1788 -2016
rect 1787 -2024 1788 -2022
rect 1794 -2018 1795 -2016
rect 1794 -2024 1795 -2022
rect 1801 -2018 1802 -2016
rect 1801 -2024 1802 -2022
rect 1808 -2018 1809 -2016
rect 1808 -2024 1809 -2022
rect 30 -2173 31 -2171
rect 30 -2179 31 -2177
rect 37 -2173 38 -2171
rect 37 -2179 38 -2177
rect 44 -2173 45 -2171
rect 44 -2179 45 -2177
rect 51 -2173 52 -2171
rect 51 -2179 52 -2177
rect 61 -2173 62 -2171
rect 61 -2179 62 -2177
rect 65 -2173 66 -2171
rect 65 -2179 66 -2177
rect 72 -2173 73 -2171
rect 72 -2179 73 -2177
rect 79 -2173 80 -2171
rect 79 -2179 80 -2177
rect 86 -2173 87 -2171
rect 86 -2179 87 -2177
rect 93 -2173 94 -2171
rect 96 -2173 97 -2171
rect 93 -2179 94 -2177
rect 96 -2179 97 -2177
rect 103 -2173 104 -2171
rect 100 -2179 101 -2177
rect 103 -2179 104 -2177
rect 107 -2173 108 -2171
rect 110 -2173 111 -2171
rect 110 -2179 111 -2177
rect 114 -2173 115 -2171
rect 114 -2179 115 -2177
rect 121 -2173 122 -2171
rect 124 -2173 125 -2171
rect 124 -2179 125 -2177
rect 128 -2173 129 -2171
rect 131 -2173 132 -2171
rect 128 -2179 129 -2177
rect 131 -2179 132 -2177
rect 135 -2173 136 -2171
rect 135 -2179 136 -2177
rect 142 -2173 143 -2171
rect 142 -2179 143 -2177
rect 149 -2173 150 -2171
rect 149 -2179 150 -2177
rect 156 -2173 157 -2171
rect 156 -2179 157 -2177
rect 163 -2173 164 -2171
rect 163 -2179 164 -2177
rect 170 -2173 171 -2171
rect 170 -2179 171 -2177
rect 177 -2173 178 -2171
rect 177 -2179 178 -2177
rect 184 -2173 185 -2171
rect 184 -2179 185 -2177
rect 191 -2173 192 -2171
rect 191 -2179 192 -2177
rect 198 -2173 199 -2171
rect 201 -2173 202 -2171
rect 201 -2179 202 -2177
rect 205 -2173 206 -2171
rect 205 -2179 206 -2177
rect 212 -2173 213 -2171
rect 212 -2179 213 -2177
rect 219 -2173 220 -2171
rect 219 -2179 220 -2177
rect 226 -2173 227 -2171
rect 229 -2173 230 -2171
rect 226 -2179 227 -2177
rect 229 -2179 230 -2177
rect 233 -2173 234 -2171
rect 233 -2179 234 -2177
rect 240 -2173 241 -2171
rect 240 -2179 241 -2177
rect 247 -2173 248 -2171
rect 250 -2173 251 -2171
rect 250 -2179 251 -2177
rect 254 -2173 255 -2171
rect 257 -2179 258 -2177
rect 261 -2173 262 -2171
rect 261 -2179 262 -2177
rect 268 -2173 269 -2171
rect 268 -2179 269 -2177
rect 275 -2173 276 -2171
rect 278 -2173 279 -2171
rect 282 -2173 283 -2171
rect 282 -2179 283 -2177
rect 289 -2173 290 -2171
rect 292 -2173 293 -2171
rect 296 -2173 297 -2171
rect 296 -2179 297 -2177
rect 303 -2173 304 -2171
rect 303 -2179 304 -2177
rect 310 -2173 311 -2171
rect 310 -2179 311 -2177
rect 317 -2173 318 -2171
rect 317 -2179 318 -2177
rect 324 -2173 325 -2171
rect 324 -2179 325 -2177
rect 331 -2173 332 -2171
rect 331 -2179 332 -2177
rect 338 -2173 339 -2171
rect 338 -2179 339 -2177
rect 345 -2173 346 -2171
rect 345 -2179 346 -2177
rect 352 -2173 353 -2171
rect 352 -2179 353 -2177
rect 359 -2173 360 -2171
rect 359 -2179 360 -2177
rect 366 -2173 367 -2171
rect 366 -2179 367 -2177
rect 373 -2173 374 -2171
rect 376 -2179 377 -2177
rect 380 -2173 381 -2171
rect 380 -2179 381 -2177
rect 387 -2173 388 -2171
rect 387 -2179 388 -2177
rect 394 -2173 395 -2171
rect 394 -2179 395 -2177
rect 401 -2173 402 -2171
rect 401 -2179 402 -2177
rect 408 -2173 409 -2171
rect 408 -2179 409 -2177
rect 418 -2173 419 -2171
rect 415 -2179 416 -2177
rect 418 -2179 419 -2177
rect 422 -2173 423 -2171
rect 422 -2179 423 -2177
rect 429 -2173 430 -2171
rect 436 -2173 437 -2171
rect 436 -2179 437 -2177
rect 443 -2173 444 -2171
rect 443 -2179 444 -2177
rect 450 -2173 451 -2171
rect 450 -2179 451 -2177
rect 457 -2173 458 -2171
rect 457 -2179 458 -2177
rect 464 -2173 465 -2171
rect 464 -2179 465 -2177
rect 471 -2173 472 -2171
rect 471 -2179 472 -2177
rect 478 -2173 479 -2171
rect 478 -2179 479 -2177
rect 485 -2173 486 -2171
rect 485 -2179 486 -2177
rect 492 -2173 493 -2171
rect 492 -2179 493 -2177
rect 499 -2173 500 -2171
rect 499 -2179 500 -2177
rect 506 -2173 507 -2171
rect 506 -2179 507 -2177
rect 513 -2173 514 -2171
rect 516 -2173 517 -2171
rect 513 -2179 514 -2177
rect 516 -2179 517 -2177
rect 520 -2173 521 -2171
rect 520 -2179 521 -2177
rect 527 -2173 528 -2171
rect 527 -2179 528 -2177
rect 534 -2179 535 -2177
rect 541 -2173 542 -2171
rect 541 -2179 542 -2177
rect 548 -2173 549 -2171
rect 548 -2179 549 -2177
rect 555 -2173 556 -2171
rect 558 -2173 559 -2171
rect 555 -2179 556 -2177
rect 558 -2179 559 -2177
rect 562 -2173 563 -2171
rect 562 -2179 563 -2177
rect 569 -2173 570 -2171
rect 569 -2179 570 -2177
rect 576 -2173 577 -2171
rect 576 -2179 577 -2177
rect 583 -2173 584 -2171
rect 586 -2173 587 -2171
rect 583 -2179 584 -2177
rect 586 -2179 587 -2177
rect 590 -2173 591 -2171
rect 590 -2179 591 -2177
rect 597 -2173 598 -2171
rect 597 -2179 598 -2177
rect 604 -2173 605 -2171
rect 604 -2179 605 -2177
rect 611 -2173 612 -2171
rect 614 -2173 615 -2171
rect 614 -2179 615 -2177
rect 618 -2173 619 -2171
rect 618 -2179 619 -2177
rect 625 -2173 626 -2171
rect 628 -2173 629 -2171
rect 625 -2179 626 -2177
rect 628 -2179 629 -2177
rect 632 -2173 633 -2171
rect 632 -2179 633 -2177
rect 639 -2173 640 -2171
rect 639 -2179 640 -2177
rect 646 -2173 647 -2171
rect 646 -2179 647 -2177
rect 653 -2173 654 -2171
rect 653 -2179 654 -2177
rect 660 -2173 661 -2171
rect 660 -2179 661 -2177
rect 667 -2173 668 -2171
rect 667 -2179 668 -2177
rect 674 -2173 675 -2171
rect 674 -2179 675 -2177
rect 681 -2173 682 -2171
rect 681 -2179 682 -2177
rect 688 -2173 689 -2171
rect 688 -2179 689 -2177
rect 695 -2173 696 -2171
rect 695 -2179 696 -2177
rect 702 -2173 703 -2171
rect 705 -2173 706 -2171
rect 702 -2179 703 -2177
rect 712 -2173 713 -2171
rect 709 -2179 710 -2177
rect 716 -2173 717 -2171
rect 716 -2179 717 -2177
rect 723 -2173 724 -2171
rect 723 -2179 724 -2177
rect 730 -2173 731 -2171
rect 730 -2179 731 -2177
rect 737 -2173 738 -2171
rect 737 -2179 738 -2177
rect 744 -2173 745 -2171
rect 744 -2179 745 -2177
rect 751 -2173 752 -2171
rect 751 -2179 752 -2177
rect 758 -2173 759 -2171
rect 758 -2179 759 -2177
rect 765 -2173 766 -2171
rect 765 -2179 766 -2177
rect 772 -2173 773 -2171
rect 772 -2179 773 -2177
rect 779 -2173 780 -2171
rect 779 -2179 780 -2177
rect 786 -2173 787 -2171
rect 786 -2179 787 -2177
rect 793 -2173 794 -2171
rect 793 -2179 794 -2177
rect 803 -2173 804 -2171
rect 803 -2179 804 -2177
rect 807 -2173 808 -2171
rect 807 -2179 808 -2177
rect 814 -2173 815 -2171
rect 817 -2173 818 -2171
rect 814 -2179 815 -2177
rect 817 -2179 818 -2177
rect 821 -2173 822 -2171
rect 821 -2179 822 -2177
rect 824 -2179 825 -2177
rect 831 -2173 832 -2171
rect 831 -2179 832 -2177
rect 835 -2173 836 -2171
rect 835 -2179 836 -2177
rect 842 -2173 843 -2171
rect 842 -2179 843 -2177
rect 849 -2173 850 -2171
rect 849 -2179 850 -2177
rect 856 -2173 857 -2171
rect 856 -2179 857 -2177
rect 863 -2173 864 -2171
rect 863 -2179 864 -2177
rect 873 -2173 874 -2171
rect 873 -2179 874 -2177
rect 877 -2173 878 -2171
rect 877 -2179 878 -2177
rect 884 -2173 885 -2171
rect 884 -2179 885 -2177
rect 891 -2173 892 -2171
rect 891 -2179 892 -2177
rect 898 -2173 899 -2171
rect 898 -2179 899 -2177
rect 905 -2173 906 -2171
rect 905 -2179 906 -2177
rect 912 -2173 913 -2171
rect 912 -2179 913 -2177
rect 919 -2173 920 -2171
rect 919 -2179 920 -2177
rect 929 -2173 930 -2171
rect 926 -2179 927 -2177
rect 929 -2179 930 -2177
rect 933 -2173 934 -2171
rect 933 -2179 934 -2177
rect 940 -2173 941 -2171
rect 940 -2179 941 -2177
rect 947 -2173 948 -2171
rect 947 -2179 948 -2177
rect 954 -2173 955 -2171
rect 954 -2179 955 -2177
rect 961 -2173 962 -2171
rect 961 -2179 962 -2177
rect 968 -2173 969 -2171
rect 968 -2179 969 -2177
rect 975 -2173 976 -2171
rect 978 -2173 979 -2171
rect 975 -2179 976 -2177
rect 978 -2179 979 -2177
rect 982 -2173 983 -2171
rect 982 -2179 983 -2177
rect 989 -2173 990 -2171
rect 989 -2179 990 -2177
rect 996 -2173 997 -2171
rect 999 -2173 1000 -2171
rect 996 -2179 997 -2177
rect 999 -2179 1000 -2177
rect 1003 -2173 1004 -2171
rect 1003 -2179 1004 -2177
rect 1010 -2173 1011 -2171
rect 1010 -2179 1011 -2177
rect 1017 -2173 1018 -2171
rect 1017 -2179 1018 -2177
rect 1024 -2173 1025 -2171
rect 1027 -2173 1028 -2171
rect 1024 -2179 1025 -2177
rect 1027 -2179 1028 -2177
rect 1031 -2173 1032 -2171
rect 1031 -2179 1032 -2177
rect 1038 -2173 1039 -2171
rect 1038 -2179 1039 -2177
rect 1045 -2173 1046 -2171
rect 1045 -2179 1046 -2177
rect 1052 -2173 1053 -2171
rect 1052 -2179 1053 -2177
rect 1059 -2173 1060 -2171
rect 1062 -2173 1063 -2171
rect 1059 -2179 1060 -2177
rect 1062 -2179 1063 -2177
rect 1066 -2173 1067 -2171
rect 1066 -2179 1067 -2177
rect 1073 -2173 1074 -2171
rect 1073 -2179 1074 -2177
rect 1080 -2173 1081 -2171
rect 1080 -2179 1081 -2177
rect 1087 -2173 1088 -2171
rect 1087 -2179 1088 -2177
rect 1094 -2173 1095 -2171
rect 1094 -2179 1095 -2177
rect 1101 -2173 1102 -2171
rect 1101 -2179 1102 -2177
rect 1108 -2173 1109 -2171
rect 1108 -2179 1109 -2177
rect 1115 -2173 1116 -2171
rect 1115 -2179 1116 -2177
rect 1125 -2173 1126 -2171
rect 1122 -2179 1123 -2177
rect 1125 -2179 1126 -2177
rect 1129 -2173 1130 -2171
rect 1132 -2173 1133 -2171
rect 1129 -2179 1130 -2177
rect 1132 -2179 1133 -2177
rect 1136 -2173 1137 -2171
rect 1136 -2179 1137 -2177
rect 1143 -2173 1144 -2171
rect 1143 -2179 1144 -2177
rect 1150 -2173 1151 -2171
rect 1150 -2179 1151 -2177
rect 1157 -2173 1158 -2171
rect 1157 -2179 1158 -2177
rect 1164 -2173 1165 -2171
rect 1164 -2179 1165 -2177
rect 1171 -2173 1172 -2171
rect 1171 -2179 1172 -2177
rect 1178 -2173 1179 -2171
rect 1178 -2179 1179 -2177
rect 1185 -2173 1186 -2171
rect 1185 -2179 1186 -2177
rect 1192 -2173 1193 -2171
rect 1195 -2173 1196 -2171
rect 1192 -2179 1193 -2177
rect 1195 -2179 1196 -2177
rect 1199 -2173 1200 -2171
rect 1199 -2179 1200 -2177
rect 1206 -2173 1207 -2171
rect 1206 -2179 1207 -2177
rect 1213 -2173 1214 -2171
rect 1213 -2179 1214 -2177
rect 1220 -2173 1221 -2171
rect 1220 -2179 1221 -2177
rect 1227 -2173 1228 -2171
rect 1227 -2179 1228 -2177
rect 1234 -2173 1235 -2171
rect 1234 -2179 1235 -2177
rect 1241 -2173 1242 -2171
rect 1241 -2179 1242 -2177
rect 1248 -2173 1249 -2171
rect 1248 -2179 1249 -2177
rect 1255 -2173 1256 -2171
rect 1255 -2179 1256 -2177
rect 1262 -2173 1263 -2171
rect 1262 -2179 1263 -2177
rect 1269 -2173 1270 -2171
rect 1269 -2179 1270 -2177
rect 1276 -2173 1277 -2171
rect 1276 -2179 1277 -2177
rect 1283 -2173 1284 -2171
rect 1283 -2179 1284 -2177
rect 1290 -2173 1291 -2171
rect 1290 -2179 1291 -2177
rect 1297 -2173 1298 -2171
rect 1297 -2179 1298 -2177
rect 1304 -2173 1305 -2171
rect 1304 -2179 1305 -2177
rect 1311 -2173 1312 -2171
rect 1314 -2173 1315 -2171
rect 1311 -2179 1312 -2177
rect 1314 -2179 1315 -2177
rect 1318 -2173 1319 -2171
rect 1318 -2179 1319 -2177
rect 1325 -2173 1326 -2171
rect 1325 -2179 1326 -2177
rect 1332 -2173 1333 -2171
rect 1332 -2179 1333 -2177
rect 1339 -2173 1340 -2171
rect 1339 -2179 1340 -2177
rect 1346 -2173 1347 -2171
rect 1346 -2179 1347 -2177
rect 1353 -2173 1354 -2171
rect 1353 -2179 1354 -2177
rect 1360 -2173 1361 -2171
rect 1360 -2179 1361 -2177
rect 1367 -2173 1368 -2171
rect 1367 -2179 1368 -2177
rect 1374 -2173 1375 -2171
rect 1374 -2179 1375 -2177
rect 1381 -2173 1382 -2171
rect 1381 -2179 1382 -2177
rect 1388 -2173 1389 -2171
rect 1388 -2179 1389 -2177
rect 1395 -2173 1396 -2171
rect 1395 -2179 1396 -2177
rect 1402 -2173 1403 -2171
rect 1402 -2179 1403 -2177
rect 1409 -2173 1410 -2171
rect 1409 -2179 1410 -2177
rect 1412 -2179 1413 -2177
rect 1416 -2173 1417 -2171
rect 1416 -2179 1417 -2177
rect 1423 -2173 1424 -2171
rect 1423 -2179 1424 -2177
rect 1430 -2173 1431 -2171
rect 1430 -2179 1431 -2177
rect 1437 -2173 1438 -2171
rect 1437 -2179 1438 -2177
rect 1444 -2173 1445 -2171
rect 1444 -2179 1445 -2177
rect 1451 -2173 1452 -2171
rect 1451 -2179 1452 -2177
rect 1458 -2173 1459 -2171
rect 1458 -2179 1459 -2177
rect 1465 -2173 1466 -2171
rect 1465 -2179 1466 -2177
rect 1472 -2173 1473 -2171
rect 1472 -2179 1473 -2177
rect 1479 -2173 1480 -2171
rect 1479 -2179 1480 -2177
rect 1486 -2173 1487 -2171
rect 1486 -2179 1487 -2177
rect 1493 -2173 1494 -2171
rect 1493 -2179 1494 -2177
rect 1500 -2173 1501 -2171
rect 1500 -2179 1501 -2177
rect 1507 -2173 1508 -2171
rect 1507 -2179 1508 -2177
rect 1514 -2173 1515 -2171
rect 1514 -2179 1515 -2177
rect 1521 -2173 1522 -2171
rect 1521 -2179 1522 -2177
rect 1528 -2173 1529 -2171
rect 1528 -2179 1529 -2177
rect 1535 -2173 1536 -2171
rect 1535 -2179 1536 -2177
rect 1542 -2173 1543 -2171
rect 1542 -2179 1543 -2177
rect 1549 -2173 1550 -2171
rect 1549 -2179 1550 -2177
rect 1556 -2173 1557 -2171
rect 1556 -2179 1557 -2177
rect 1563 -2173 1564 -2171
rect 1563 -2179 1564 -2177
rect 1570 -2173 1571 -2171
rect 1570 -2179 1571 -2177
rect 1577 -2173 1578 -2171
rect 1577 -2179 1578 -2177
rect 1584 -2173 1585 -2171
rect 1584 -2179 1585 -2177
rect 1591 -2173 1592 -2171
rect 1594 -2173 1595 -2171
rect 1591 -2179 1592 -2177
rect 1598 -2173 1599 -2171
rect 1598 -2179 1599 -2177
rect 1605 -2173 1606 -2171
rect 1605 -2179 1606 -2177
rect 1612 -2173 1613 -2171
rect 1612 -2179 1613 -2177
rect 1619 -2173 1620 -2171
rect 1619 -2179 1620 -2177
rect 1626 -2173 1627 -2171
rect 1626 -2179 1627 -2177
rect 1633 -2173 1634 -2171
rect 1633 -2179 1634 -2177
rect 1640 -2173 1641 -2171
rect 1640 -2179 1641 -2177
rect 1647 -2173 1648 -2171
rect 1647 -2179 1648 -2177
rect 1654 -2173 1655 -2171
rect 1654 -2179 1655 -2177
rect 1661 -2173 1662 -2171
rect 1661 -2179 1662 -2177
rect 1668 -2173 1669 -2171
rect 1668 -2179 1669 -2177
rect 1675 -2173 1676 -2171
rect 1675 -2179 1676 -2177
rect 1682 -2173 1683 -2171
rect 1682 -2179 1683 -2177
rect 1689 -2173 1690 -2171
rect 1689 -2179 1690 -2177
rect 1696 -2173 1697 -2171
rect 1696 -2179 1697 -2177
rect 1703 -2173 1704 -2171
rect 1703 -2179 1704 -2177
rect 1710 -2173 1711 -2171
rect 1713 -2173 1714 -2171
rect 1710 -2179 1711 -2177
rect 1713 -2179 1714 -2177
rect 1717 -2179 1718 -2177
rect 1720 -2179 1721 -2177
rect 1724 -2173 1725 -2171
rect 1724 -2179 1725 -2177
rect 1731 -2173 1732 -2171
rect 1731 -2179 1732 -2177
rect 1738 -2173 1739 -2171
rect 1738 -2179 1739 -2177
rect 30 -2302 31 -2300
rect 30 -2308 31 -2306
rect 44 -2302 45 -2300
rect 44 -2308 45 -2306
rect 58 -2302 59 -2300
rect 58 -2308 59 -2306
rect 65 -2302 66 -2300
rect 65 -2308 66 -2306
rect 72 -2302 73 -2300
rect 72 -2308 73 -2306
rect 79 -2302 80 -2300
rect 79 -2308 80 -2306
rect 86 -2302 87 -2300
rect 86 -2308 87 -2306
rect 93 -2302 94 -2300
rect 93 -2308 94 -2306
rect 100 -2302 101 -2300
rect 100 -2308 101 -2306
rect 107 -2302 108 -2300
rect 107 -2308 108 -2306
rect 114 -2302 115 -2300
rect 114 -2308 115 -2306
rect 121 -2302 122 -2300
rect 121 -2308 122 -2306
rect 128 -2302 129 -2300
rect 128 -2308 129 -2306
rect 135 -2302 136 -2300
rect 138 -2302 139 -2300
rect 138 -2308 139 -2306
rect 142 -2302 143 -2300
rect 145 -2302 146 -2300
rect 142 -2308 143 -2306
rect 149 -2302 150 -2300
rect 152 -2302 153 -2300
rect 149 -2308 150 -2306
rect 152 -2308 153 -2306
rect 156 -2302 157 -2300
rect 156 -2308 157 -2306
rect 163 -2302 164 -2300
rect 163 -2308 164 -2306
rect 170 -2302 171 -2300
rect 170 -2308 171 -2306
rect 177 -2302 178 -2300
rect 177 -2308 178 -2306
rect 184 -2302 185 -2300
rect 184 -2308 185 -2306
rect 191 -2302 192 -2300
rect 191 -2308 192 -2306
rect 198 -2302 199 -2300
rect 198 -2308 199 -2306
rect 205 -2302 206 -2300
rect 208 -2302 209 -2300
rect 208 -2308 209 -2306
rect 215 -2302 216 -2300
rect 212 -2308 213 -2306
rect 215 -2308 216 -2306
rect 219 -2302 220 -2300
rect 219 -2308 220 -2306
rect 226 -2302 227 -2300
rect 226 -2308 227 -2306
rect 233 -2302 234 -2300
rect 233 -2308 234 -2306
rect 240 -2302 241 -2300
rect 240 -2308 241 -2306
rect 247 -2302 248 -2300
rect 247 -2308 248 -2306
rect 254 -2302 255 -2300
rect 254 -2308 255 -2306
rect 261 -2302 262 -2300
rect 261 -2308 262 -2306
rect 268 -2302 269 -2300
rect 268 -2308 269 -2306
rect 275 -2302 276 -2300
rect 275 -2308 276 -2306
rect 282 -2302 283 -2300
rect 285 -2302 286 -2300
rect 282 -2308 283 -2306
rect 289 -2302 290 -2300
rect 289 -2308 290 -2306
rect 296 -2302 297 -2300
rect 296 -2308 297 -2306
rect 303 -2302 304 -2300
rect 303 -2308 304 -2306
rect 310 -2302 311 -2300
rect 310 -2308 311 -2306
rect 317 -2302 318 -2300
rect 317 -2308 318 -2306
rect 324 -2302 325 -2300
rect 324 -2308 325 -2306
rect 331 -2302 332 -2300
rect 331 -2308 332 -2306
rect 338 -2302 339 -2300
rect 338 -2308 339 -2306
rect 345 -2302 346 -2300
rect 345 -2308 346 -2306
rect 352 -2302 353 -2300
rect 352 -2308 353 -2306
rect 359 -2302 360 -2300
rect 359 -2308 360 -2306
rect 366 -2302 367 -2300
rect 366 -2308 367 -2306
rect 373 -2302 374 -2300
rect 373 -2308 374 -2306
rect 380 -2302 381 -2300
rect 380 -2308 381 -2306
rect 387 -2302 388 -2300
rect 387 -2308 388 -2306
rect 394 -2302 395 -2300
rect 394 -2308 395 -2306
rect 401 -2302 402 -2300
rect 401 -2308 402 -2306
rect 408 -2302 409 -2300
rect 408 -2308 409 -2306
rect 415 -2302 416 -2300
rect 415 -2308 416 -2306
rect 422 -2302 423 -2300
rect 422 -2308 423 -2306
rect 429 -2308 430 -2306
rect 436 -2302 437 -2300
rect 436 -2308 437 -2306
rect 443 -2302 444 -2300
rect 443 -2308 444 -2306
rect 450 -2302 451 -2300
rect 450 -2308 451 -2306
rect 453 -2308 454 -2306
rect 457 -2302 458 -2300
rect 457 -2308 458 -2306
rect 464 -2302 465 -2300
rect 464 -2308 465 -2306
rect 471 -2302 472 -2300
rect 471 -2308 472 -2306
rect 478 -2302 479 -2300
rect 478 -2308 479 -2306
rect 485 -2302 486 -2300
rect 495 -2302 496 -2300
rect 492 -2308 493 -2306
rect 495 -2308 496 -2306
rect 499 -2302 500 -2300
rect 499 -2308 500 -2306
rect 506 -2302 507 -2300
rect 509 -2302 510 -2300
rect 506 -2308 507 -2306
rect 509 -2308 510 -2306
rect 513 -2302 514 -2300
rect 513 -2308 514 -2306
rect 520 -2302 521 -2300
rect 520 -2308 521 -2306
rect 527 -2302 528 -2300
rect 527 -2308 528 -2306
rect 534 -2302 535 -2300
rect 534 -2308 535 -2306
rect 541 -2302 542 -2300
rect 541 -2308 542 -2306
rect 548 -2302 549 -2300
rect 548 -2308 549 -2306
rect 555 -2302 556 -2300
rect 555 -2308 556 -2306
rect 562 -2302 563 -2300
rect 562 -2308 563 -2306
rect 569 -2302 570 -2300
rect 569 -2308 570 -2306
rect 579 -2302 580 -2300
rect 576 -2308 577 -2306
rect 579 -2308 580 -2306
rect 583 -2302 584 -2300
rect 583 -2308 584 -2306
rect 590 -2302 591 -2300
rect 590 -2308 591 -2306
rect 597 -2302 598 -2300
rect 600 -2302 601 -2300
rect 600 -2308 601 -2306
rect 604 -2302 605 -2300
rect 604 -2308 605 -2306
rect 611 -2302 612 -2300
rect 611 -2308 612 -2306
rect 618 -2302 619 -2300
rect 618 -2308 619 -2306
rect 628 -2302 629 -2300
rect 625 -2308 626 -2306
rect 632 -2302 633 -2300
rect 632 -2308 633 -2306
rect 642 -2302 643 -2300
rect 639 -2308 640 -2306
rect 642 -2308 643 -2306
rect 646 -2302 647 -2300
rect 646 -2308 647 -2306
rect 653 -2302 654 -2300
rect 653 -2308 654 -2306
rect 660 -2302 661 -2300
rect 660 -2308 661 -2306
rect 667 -2302 668 -2300
rect 670 -2302 671 -2300
rect 670 -2308 671 -2306
rect 677 -2302 678 -2300
rect 677 -2308 678 -2306
rect 681 -2302 682 -2300
rect 681 -2308 682 -2306
rect 688 -2302 689 -2300
rect 691 -2302 692 -2300
rect 688 -2308 689 -2306
rect 691 -2308 692 -2306
rect 698 -2302 699 -2300
rect 695 -2308 696 -2306
rect 702 -2302 703 -2300
rect 705 -2302 706 -2300
rect 702 -2308 703 -2306
rect 705 -2308 706 -2306
rect 709 -2302 710 -2300
rect 709 -2308 710 -2306
rect 716 -2302 717 -2300
rect 716 -2308 717 -2306
rect 723 -2302 724 -2300
rect 723 -2308 724 -2306
rect 730 -2302 731 -2300
rect 730 -2308 731 -2306
rect 737 -2302 738 -2300
rect 737 -2308 738 -2306
rect 744 -2302 745 -2300
rect 744 -2308 745 -2306
rect 751 -2302 752 -2300
rect 751 -2308 752 -2306
rect 758 -2302 759 -2300
rect 761 -2302 762 -2300
rect 758 -2308 759 -2306
rect 761 -2308 762 -2306
rect 765 -2302 766 -2300
rect 765 -2308 766 -2306
rect 772 -2302 773 -2300
rect 772 -2308 773 -2306
rect 779 -2302 780 -2300
rect 779 -2308 780 -2306
rect 782 -2308 783 -2306
rect 786 -2302 787 -2300
rect 786 -2308 787 -2306
rect 793 -2302 794 -2300
rect 793 -2308 794 -2306
rect 800 -2302 801 -2300
rect 800 -2308 801 -2306
rect 807 -2302 808 -2300
rect 807 -2308 808 -2306
rect 814 -2302 815 -2300
rect 814 -2308 815 -2306
rect 821 -2302 822 -2300
rect 821 -2308 822 -2306
rect 828 -2302 829 -2300
rect 828 -2308 829 -2306
rect 835 -2302 836 -2300
rect 838 -2302 839 -2300
rect 835 -2308 836 -2306
rect 838 -2308 839 -2306
rect 842 -2302 843 -2300
rect 842 -2308 843 -2306
rect 849 -2302 850 -2300
rect 849 -2308 850 -2306
rect 856 -2302 857 -2300
rect 856 -2308 857 -2306
rect 863 -2302 864 -2300
rect 866 -2302 867 -2300
rect 863 -2308 864 -2306
rect 866 -2308 867 -2306
rect 870 -2302 871 -2300
rect 873 -2302 874 -2300
rect 870 -2308 871 -2306
rect 873 -2308 874 -2306
rect 877 -2302 878 -2300
rect 877 -2308 878 -2306
rect 884 -2302 885 -2300
rect 884 -2308 885 -2306
rect 891 -2302 892 -2300
rect 891 -2308 892 -2306
rect 898 -2302 899 -2300
rect 898 -2308 899 -2306
rect 905 -2302 906 -2300
rect 905 -2308 906 -2306
rect 912 -2302 913 -2300
rect 912 -2308 913 -2306
rect 915 -2308 916 -2306
rect 919 -2302 920 -2300
rect 919 -2308 920 -2306
rect 926 -2302 927 -2300
rect 926 -2308 927 -2306
rect 933 -2302 934 -2300
rect 933 -2308 934 -2306
rect 943 -2302 944 -2300
rect 940 -2308 941 -2306
rect 943 -2308 944 -2306
rect 947 -2302 948 -2300
rect 947 -2308 948 -2306
rect 954 -2302 955 -2300
rect 954 -2308 955 -2306
rect 961 -2302 962 -2300
rect 961 -2308 962 -2306
rect 968 -2302 969 -2300
rect 968 -2308 969 -2306
rect 975 -2302 976 -2300
rect 975 -2308 976 -2306
rect 982 -2302 983 -2300
rect 982 -2308 983 -2306
rect 989 -2302 990 -2300
rect 989 -2308 990 -2306
rect 992 -2308 993 -2306
rect 996 -2302 997 -2300
rect 996 -2308 997 -2306
rect 1003 -2302 1004 -2300
rect 1003 -2308 1004 -2306
rect 1010 -2302 1011 -2300
rect 1010 -2308 1011 -2306
rect 1017 -2302 1018 -2300
rect 1020 -2302 1021 -2300
rect 1017 -2308 1018 -2306
rect 1020 -2308 1021 -2306
rect 1024 -2302 1025 -2300
rect 1027 -2302 1028 -2300
rect 1024 -2308 1025 -2306
rect 1031 -2302 1032 -2300
rect 1031 -2308 1032 -2306
rect 1038 -2302 1039 -2300
rect 1041 -2302 1042 -2300
rect 1038 -2308 1039 -2306
rect 1041 -2308 1042 -2306
rect 1045 -2302 1046 -2300
rect 1045 -2308 1046 -2306
rect 1052 -2302 1053 -2300
rect 1052 -2308 1053 -2306
rect 1059 -2302 1060 -2300
rect 1059 -2308 1060 -2306
rect 1066 -2302 1067 -2300
rect 1066 -2308 1067 -2306
rect 1073 -2302 1074 -2300
rect 1073 -2308 1074 -2306
rect 1080 -2302 1081 -2300
rect 1080 -2308 1081 -2306
rect 1087 -2302 1088 -2300
rect 1087 -2308 1088 -2306
rect 1094 -2302 1095 -2300
rect 1094 -2308 1095 -2306
rect 1101 -2302 1102 -2300
rect 1101 -2308 1102 -2306
rect 1108 -2302 1109 -2300
rect 1108 -2308 1109 -2306
rect 1115 -2302 1116 -2300
rect 1115 -2308 1116 -2306
rect 1122 -2302 1123 -2300
rect 1122 -2308 1123 -2306
rect 1129 -2302 1130 -2300
rect 1129 -2308 1130 -2306
rect 1136 -2302 1137 -2300
rect 1136 -2308 1137 -2306
rect 1143 -2302 1144 -2300
rect 1143 -2308 1144 -2306
rect 1150 -2302 1151 -2300
rect 1150 -2308 1151 -2306
rect 1157 -2302 1158 -2300
rect 1157 -2308 1158 -2306
rect 1164 -2302 1165 -2300
rect 1164 -2308 1165 -2306
rect 1174 -2302 1175 -2300
rect 1171 -2308 1172 -2306
rect 1174 -2308 1175 -2306
rect 1178 -2302 1179 -2300
rect 1178 -2308 1179 -2306
rect 1185 -2302 1186 -2300
rect 1185 -2308 1186 -2306
rect 1192 -2302 1193 -2300
rect 1192 -2308 1193 -2306
rect 1202 -2302 1203 -2300
rect 1202 -2308 1203 -2306
rect 1206 -2302 1207 -2300
rect 1206 -2308 1207 -2306
rect 1213 -2302 1214 -2300
rect 1213 -2308 1214 -2306
rect 1220 -2302 1221 -2300
rect 1220 -2308 1221 -2306
rect 1227 -2302 1228 -2300
rect 1227 -2308 1228 -2306
rect 1234 -2302 1235 -2300
rect 1234 -2308 1235 -2306
rect 1241 -2302 1242 -2300
rect 1241 -2308 1242 -2306
rect 1244 -2308 1245 -2306
rect 1248 -2302 1249 -2300
rect 1248 -2308 1249 -2306
rect 1255 -2302 1256 -2300
rect 1255 -2308 1256 -2306
rect 1262 -2302 1263 -2300
rect 1262 -2308 1263 -2306
rect 1269 -2302 1270 -2300
rect 1269 -2308 1270 -2306
rect 1276 -2302 1277 -2300
rect 1276 -2308 1277 -2306
rect 1283 -2302 1284 -2300
rect 1283 -2308 1284 -2306
rect 1290 -2302 1291 -2300
rect 1290 -2308 1291 -2306
rect 1297 -2302 1298 -2300
rect 1297 -2308 1298 -2306
rect 1304 -2302 1305 -2300
rect 1304 -2308 1305 -2306
rect 1311 -2302 1312 -2300
rect 1311 -2308 1312 -2306
rect 1318 -2302 1319 -2300
rect 1318 -2308 1319 -2306
rect 1325 -2302 1326 -2300
rect 1325 -2308 1326 -2306
rect 1332 -2302 1333 -2300
rect 1332 -2308 1333 -2306
rect 1339 -2302 1340 -2300
rect 1339 -2308 1340 -2306
rect 1346 -2302 1347 -2300
rect 1346 -2308 1347 -2306
rect 1353 -2302 1354 -2300
rect 1353 -2308 1354 -2306
rect 1360 -2302 1361 -2300
rect 1360 -2308 1361 -2306
rect 1367 -2302 1368 -2300
rect 1367 -2308 1368 -2306
rect 1374 -2302 1375 -2300
rect 1374 -2308 1375 -2306
rect 1381 -2302 1382 -2300
rect 1381 -2308 1382 -2306
rect 1388 -2302 1389 -2300
rect 1388 -2308 1389 -2306
rect 1395 -2302 1396 -2300
rect 1395 -2308 1396 -2306
rect 1402 -2302 1403 -2300
rect 1402 -2308 1403 -2306
rect 1409 -2302 1410 -2300
rect 1412 -2302 1413 -2300
rect 1409 -2308 1410 -2306
rect 1416 -2302 1417 -2300
rect 1416 -2308 1417 -2306
rect 1423 -2302 1424 -2300
rect 1423 -2308 1424 -2306
rect 1430 -2302 1431 -2300
rect 1430 -2308 1431 -2306
rect 1437 -2302 1438 -2300
rect 1437 -2308 1438 -2306
rect 1444 -2302 1445 -2300
rect 1444 -2308 1445 -2306
rect 1451 -2302 1452 -2300
rect 1451 -2308 1452 -2306
rect 1458 -2302 1459 -2300
rect 1458 -2308 1459 -2306
rect 1465 -2302 1466 -2300
rect 1465 -2308 1466 -2306
rect 1472 -2302 1473 -2300
rect 1472 -2308 1473 -2306
rect 1479 -2302 1480 -2300
rect 1479 -2308 1480 -2306
rect 1486 -2302 1487 -2300
rect 1486 -2308 1487 -2306
rect 1493 -2302 1494 -2300
rect 1493 -2308 1494 -2306
rect 1500 -2302 1501 -2300
rect 1500 -2308 1501 -2306
rect 1507 -2302 1508 -2300
rect 1507 -2308 1508 -2306
rect 1514 -2302 1515 -2300
rect 1514 -2308 1515 -2306
rect 1521 -2302 1522 -2300
rect 1521 -2308 1522 -2306
rect 1528 -2302 1529 -2300
rect 1528 -2308 1529 -2306
rect 1535 -2302 1536 -2300
rect 1535 -2308 1536 -2306
rect 1542 -2302 1543 -2300
rect 1542 -2308 1543 -2306
rect 1549 -2302 1550 -2300
rect 1549 -2308 1550 -2306
rect 1556 -2302 1557 -2300
rect 1556 -2308 1557 -2306
rect 1563 -2302 1564 -2300
rect 1563 -2308 1564 -2306
rect 1570 -2302 1571 -2300
rect 1570 -2308 1571 -2306
rect 1577 -2302 1578 -2300
rect 1577 -2308 1578 -2306
rect 1584 -2302 1585 -2300
rect 1584 -2308 1585 -2306
rect 1591 -2302 1592 -2300
rect 1591 -2308 1592 -2306
rect 1598 -2302 1599 -2300
rect 1598 -2308 1599 -2306
rect 1605 -2302 1606 -2300
rect 1605 -2308 1606 -2306
rect 1612 -2302 1613 -2300
rect 1612 -2308 1613 -2306
rect 1619 -2302 1620 -2300
rect 1619 -2308 1620 -2306
rect 1626 -2302 1627 -2300
rect 1626 -2308 1627 -2306
rect 1633 -2302 1634 -2300
rect 1633 -2308 1634 -2306
rect 1640 -2302 1641 -2300
rect 1640 -2308 1641 -2306
rect 1647 -2302 1648 -2300
rect 1650 -2302 1651 -2300
rect 1647 -2308 1648 -2306
rect 1650 -2308 1651 -2306
rect 1654 -2308 1655 -2306
rect 1661 -2302 1662 -2300
rect 1661 -2308 1662 -2306
rect 1668 -2302 1669 -2300
rect 1671 -2302 1672 -2300
rect 1668 -2308 1669 -2306
rect 1671 -2308 1672 -2306
rect 1675 -2302 1676 -2300
rect 1675 -2308 1676 -2306
rect 1682 -2302 1683 -2300
rect 1682 -2308 1683 -2306
rect 1689 -2302 1690 -2300
rect 1689 -2308 1690 -2306
rect 1696 -2302 1697 -2300
rect 1696 -2308 1697 -2306
rect 44 -2423 45 -2421
rect 44 -2429 45 -2427
rect 51 -2423 52 -2421
rect 51 -2429 52 -2427
rect 58 -2423 59 -2421
rect 58 -2429 59 -2427
rect 65 -2423 66 -2421
rect 65 -2429 66 -2427
rect 72 -2423 73 -2421
rect 72 -2429 73 -2427
rect 79 -2423 80 -2421
rect 79 -2429 80 -2427
rect 86 -2423 87 -2421
rect 86 -2429 87 -2427
rect 93 -2423 94 -2421
rect 93 -2429 94 -2427
rect 100 -2423 101 -2421
rect 100 -2429 101 -2427
rect 107 -2429 108 -2427
rect 110 -2429 111 -2427
rect 114 -2423 115 -2421
rect 117 -2423 118 -2421
rect 114 -2429 115 -2427
rect 117 -2429 118 -2427
rect 121 -2423 122 -2421
rect 121 -2429 122 -2427
rect 128 -2423 129 -2421
rect 128 -2429 129 -2427
rect 135 -2423 136 -2421
rect 135 -2429 136 -2427
rect 142 -2423 143 -2421
rect 142 -2429 143 -2427
rect 149 -2423 150 -2421
rect 149 -2429 150 -2427
rect 156 -2423 157 -2421
rect 156 -2429 157 -2427
rect 163 -2423 164 -2421
rect 163 -2429 164 -2427
rect 170 -2423 171 -2421
rect 170 -2429 171 -2427
rect 177 -2423 178 -2421
rect 177 -2429 178 -2427
rect 184 -2423 185 -2421
rect 184 -2429 185 -2427
rect 191 -2423 192 -2421
rect 191 -2429 192 -2427
rect 198 -2423 199 -2421
rect 198 -2429 199 -2427
rect 205 -2423 206 -2421
rect 205 -2429 206 -2427
rect 212 -2423 213 -2421
rect 212 -2429 213 -2427
rect 219 -2423 220 -2421
rect 219 -2429 220 -2427
rect 226 -2423 227 -2421
rect 229 -2423 230 -2421
rect 229 -2429 230 -2427
rect 233 -2423 234 -2421
rect 233 -2429 234 -2427
rect 240 -2423 241 -2421
rect 240 -2429 241 -2427
rect 247 -2423 248 -2421
rect 247 -2429 248 -2427
rect 254 -2423 255 -2421
rect 254 -2429 255 -2427
rect 261 -2423 262 -2421
rect 261 -2429 262 -2427
rect 268 -2423 269 -2421
rect 268 -2429 269 -2427
rect 275 -2423 276 -2421
rect 275 -2429 276 -2427
rect 282 -2423 283 -2421
rect 285 -2423 286 -2421
rect 282 -2429 283 -2427
rect 289 -2423 290 -2421
rect 289 -2429 290 -2427
rect 296 -2423 297 -2421
rect 296 -2429 297 -2427
rect 303 -2423 304 -2421
rect 303 -2429 304 -2427
rect 310 -2423 311 -2421
rect 310 -2429 311 -2427
rect 317 -2423 318 -2421
rect 317 -2429 318 -2427
rect 324 -2423 325 -2421
rect 324 -2429 325 -2427
rect 331 -2423 332 -2421
rect 331 -2429 332 -2427
rect 338 -2423 339 -2421
rect 338 -2429 339 -2427
rect 345 -2423 346 -2421
rect 345 -2429 346 -2427
rect 352 -2423 353 -2421
rect 352 -2429 353 -2427
rect 359 -2423 360 -2421
rect 359 -2429 360 -2427
rect 366 -2423 367 -2421
rect 366 -2429 367 -2427
rect 373 -2423 374 -2421
rect 373 -2429 374 -2427
rect 380 -2423 381 -2421
rect 380 -2429 381 -2427
rect 387 -2423 388 -2421
rect 387 -2429 388 -2427
rect 394 -2423 395 -2421
rect 394 -2429 395 -2427
rect 401 -2423 402 -2421
rect 404 -2423 405 -2421
rect 401 -2429 402 -2427
rect 404 -2429 405 -2427
rect 408 -2423 409 -2421
rect 408 -2429 409 -2427
rect 415 -2423 416 -2421
rect 415 -2429 416 -2427
rect 422 -2423 423 -2421
rect 422 -2429 423 -2427
rect 429 -2423 430 -2421
rect 429 -2429 430 -2427
rect 436 -2423 437 -2421
rect 436 -2429 437 -2427
rect 443 -2423 444 -2421
rect 443 -2429 444 -2427
rect 450 -2423 451 -2421
rect 450 -2429 451 -2427
rect 457 -2423 458 -2421
rect 457 -2429 458 -2427
rect 464 -2423 465 -2421
rect 464 -2429 465 -2427
rect 471 -2423 472 -2421
rect 471 -2429 472 -2427
rect 478 -2423 479 -2421
rect 478 -2429 479 -2427
rect 485 -2429 486 -2427
rect 492 -2423 493 -2421
rect 492 -2429 493 -2427
rect 499 -2423 500 -2421
rect 499 -2429 500 -2427
rect 506 -2423 507 -2421
rect 506 -2429 507 -2427
rect 513 -2423 514 -2421
rect 513 -2429 514 -2427
rect 520 -2423 521 -2421
rect 523 -2423 524 -2421
rect 520 -2429 521 -2427
rect 523 -2429 524 -2427
rect 527 -2423 528 -2421
rect 527 -2429 528 -2427
rect 534 -2423 535 -2421
rect 534 -2429 535 -2427
rect 541 -2423 542 -2421
rect 541 -2429 542 -2427
rect 548 -2423 549 -2421
rect 548 -2429 549 -2427
rect 555 -2423 556 -2421
rect 555 -2429 556 -2427
rect 562 -2423 563 -2421
rect 562 -2429 563 -2427
rect 565 -2429 566 -2427
rect 569 -2423 570 -2421
rect 569 -2429 570 -2427
rect 576 -2423 577 -2421
rect 576 -2429 577 -2427
rect 583 -2423 584 -2421
rect 586 -2423 587 -2421
rect 583 -2429 584 -2427
rect 586 -2429 587 -2427
rect 590 -2423 591 -2421
rect 590 -2429 591 -2427
rect 597 -2423 598 -2421
rect 597 -2429 598 -2427
rect 604 -2423 605 -2421
rect 604 -2429 605 -2427
rect 611 -2423 612 -2421
rect 611 -2429 612 -2427
rect 614 -2429 615 -2427
rect 618 -2423 619 -2421
rect 621 -2423 622 -2421
rect 618 -2429 619 -2427
rect 621 -2429 622 -2427
rect 625 -2423 626 -2421
rect 625 -2429 626 -2427
rect 632 -2423 633 -2421
rect 635 -2423 636 -2421
rect 632 -2429 633 -2427
rect 639 -2423 640 -2421
rect 639 -2429 640 -2427
rect 646 -2423 647 -2421
rect 649 -2423 650 -2421
rect 646 -2429 647 -2427
rect 649 -2429 650 -2427
rect 653 -2423 654 -2421
rect 653 -2429 654 -2427
rect 660 -2423 661 -2421
rect 660 -2429 661 -2427
rect 667 -2423 668 -2421
rect 667 -2429 668 -2427
rect 674 -2423 675 -2421
rect 674 -2429 675 -2427
rect 681 -2423 682 -2421
rect 684 -2423 685 -2421
rect 681 -2429 682 -2427
rect 684 -2429 685 -2427
rect 688 -2423 689 -2421
rect 688 -2429 689 -2427
rect 695 -2423 696 -2421
rect 695 -2429 696 -2427
rect 702 -2423 703 -2421
rect 702 -2429 703 -2427
rect 709 -2423 710 -2421
rect 709 -2429 710 -2427
rect 716 -2423 717 -2421
rect 716 -2429 717 -2427
rect 723 -2423 724 -2421
rect 723 -2429 724 -2427
rect 730 -2423 731 -2421
rect 733 -2423 734 -2421
rect 730 -2429 731 -2427
rect 733 -2429 734 -2427
rect 737 -2423 738 -2421
rect 740 -2423 741 -2421
rect 737 -2429 738 -2427
rect 740 -2429 741 -2427
rect 744 -2423 745 -2421
rect 747 -2423 748 -2421
rect 744 -2429 745 -2427
rect 747 -2429 748 -2427
rect 751 -2423 752 -2421
rect 751 -2429 752 -2427
rect 758 -2423 759 -2421
rect 758 -2429 759 -2427
rect 765 -2423 766 -2421
rect 765 -2429 766 -2427
rect 772 -2423 773 -2421
rect 775 -2423 776 -2421
rect 772 -2429 773 -2427
rect 775 -2429 776 -2427
rect 779 -2423 780 -2421
rect 779 -2429 780 -2427
rect 786 -2423 787 -2421
rect 786 -2429 787 -2427
rect 793 -2423 794 -2421
rect 793 -2429 794 -2427
rect 800 -2423 801 -2421
rect 800 -2429 801 -2427
rect 807 -2423 808 -2421
rect 807 -2429 808 -2427
rect 814 -2423 815 -2421
rect 814 -2429 815 -2427
rect 821 -2423 822 -2421
rect 821 -2429 822 -2427
rect 828 -2423 829 -2421
rect 828 -2429 829 -2427
rect 835 -2423 836 -2421
rect 835 -2429 836 -2427
rect 838 -2429 839 -2427
rect 842 -2423 843 -2421
rect 842 -2429 843 -2427
rect 849 -2429 850 -2427
rect 852 -2429 853 -2427
rect 859 -2423 860 -2421
rect 856 -2429 857 -2427
rect 859 -2429 860 -2427
rect 863 -2423 864 -2421
rect 863 -2429 864 -2427
rect 870 -2423 871 -2421
rect 870 -2429 871 -2427
rect 877 -2423 878 -2421
rect 877 -2429 878 -2427
rect 884 -2423 885 -2421
rect 884 -2429 885 -2427
rect 891 -2423 892 -2421
rect 891 -2429 892 -2427
rect 898 -2423 899 -2421
rect 898 -2429 899 -2427
rect 905 -2423 906 -2421
rect 905 -2429 906 -2427
rect 912 -2423 913 -2421
rect 912 -2429 913 -2427
rect 919 -2423 920 -2421
rect 919 -2429 920 -2427
rect 926 -2423 927 -2421
rect 929 -2423 930 -2421
rect 926 -2429 927 -2427
rect 929 -2429 930 -2427
rect 933 -2423 934 -2421
rect 933 -2429 934 -2427
rect 940 -2423 941 -2421
rect 940 -2429 941 -2427
rect 947 -2423 948 -2421
rect 947 -2429 948 -2427
rect 954 -2423 955 -2421
rect 954 -2429 955 -2427
rect 961 -2423 962 -2421
rect 961 -2429 962 -2427
rect 971 -2423 972 -2421
rect 968 -2429 969 -2427
rect 971 -2429 972 -2427
rect 975 -2423 976 -2421
rect 975 -2429 976 -2427
rect 982 -2423 983 -2421
rect 982 -2429 983 -2427
rect 989 -2423 990 -2421
rect 992 -2423 993 -2421
rect 989 -2429 990 -2427
rect 996 -2423 997 -2421
rect 996 -2429 997 -2427
rect 1003 -2423 1004 -2421
rect 1003 -2429 1004 -2427
rect 1010 -2423 1011 -2421
rect 1010 -2429 1011 -2427
rect 1017 -2423 1018 -2421
rect 1017 -2429 1018 -2427
rect 1024 -2423 1025 -2421
rect 1024 -2429 1025 -2427
rect 1031 -2423 1032 -2421
rect 1031 -2429 1032 -2427
rect 1038 -2423 1039 -2421
rect 1038 -2429 1039 -2427
rect 1045 -2423 1046 -2421
rect 1045 -2429 1046 -2427
rect 1052 -2423 1053 -2421
rect 1052 -2429 1053 -2427
rect 1059 -2423 1060 -2421
rect 1059 -2429 1060 -2427
rect 1066 -2423 1067 -2421
rect 1066 -2429 1067 -2427
rect 1073 -2423 1074 -2421
rect 1073 -2429 1074 -2427
rect 1080 -2423 1081 -2421
rect 1080 -2429 1081 -2427
rect 1087 -2423 1088 -2421
rect 1087 -2429 1088 -2427
rect 1094 -2423 1095 -2421
rect 1094 -2429 1095 -2427
rect 1104 -2423 1105 -2421
rect 1104 -2429 1105 -2427
rect 1108 -2423 1109 -2421
rect 1108 -2429 1109 -2427
rect 1115 -2423 1116 -2421
rect 1115 -2429 1116 -2427
rect 1122 -2423 1123 -2421
rect 1125 -2429 1126 -2427
rect 1129 -2423 1130 -2421
rect 1129 -2429 1130 -2427
rect 1136 -2423 1137 -2421
rect 1136 -2429 1137 -2427
rect 1143 -2423 1144 -2421
rect 1143 -2429 1144 -2427
rect 1150 -2423 1151 -2421
rect 1150 -2429 1151 -2427
rect 1157 -2423 1158 -2421
rect 1157 -2429 1158 -2427
rect 1164 -2423 1165 -2421
rect 1164 -2429 1165 -2427
rect 1171 -2423 1172 -2421
rect 1171 -2429 1172 -2427
rect 1178 -2423 1179 -2421
rect 1178 -2429 1179 -2427
rect 1185 -2423 1186 -2421
rect 1185 -2429 1186 -2427
rect 1188 -2429 1189 -2427
rect 1192 -2423 1193 -2421
rect 1192 -2429 1193 -2427
rect 1199 -2423 1200 -2421
rect 1202 -2423 1203 -2421
rect 1199 -2429 1200 -2427
rect 1202 -2429 1203 -2427
rect 1206 -2423 1207 -2421
rect 1206 -2429 1207 -2427
rect 1213 -2423 1214 -2421
rect 1213 -2429 1214 -2427
rect 1220 -2423 1221 -2421
rect 1220 -2429 1221 -2427
rect 1227 -2423 1228 -2421
rect 1227 -2429 1228 -2427
rect 1234 -2423 1235 -2421
rect 1237 -2423 1238 -2421
rect 1237 -2429 1238 -2427
rect 1241 -2423 1242 -2421
rect 1241 -2429 1242 -2427
rect 1248 -2423 1249 -2421
rect 1251 -2423 1252 -2421
rect 1251 -2429 1252 -2427
rect 1255 -2423 1256 -2421
rect 1255 -2429 1256 -2427
rect 1262 -2423 1263 -2421
rect 1262 -2429 1263 -2427
rect 1269 -2423 1270 -2421
rect 1269 -2429 1270 -2427
rect 1276 -2423 1277 -2421
rect 1276 -2429 1277 -2427
rect 1283 -2423 1284 -2421
rect 1283 -2429 1284 -2427
rect 1290 -2423 1291 -2421
rect 1293 -2423 1294 -2421
rect 1290 -2429 1291 -2427
rect 1297 -2423 1298 -2421
rect 1297 -2429 1298 -2427
rect 1304 -2423 1305 -2421
rect 1304 -2429 1305 -2427
rect 1311 -2423 1312 -2421
rect 1311 -2429 1312 -2427
rect 1318 -2423 1319 -2421
rect 1318 -2429 1319 -2427
rect 1325 -2423 1326 -2421
rect 1325 -2429 1326 -2427
rect 1332 -2423 1333 -2421
rect 1332 -2429 1333 -2427
rect 1339 -2423 1340 -2421
rect 1339 -2429 1340 -2427
rect 1346 -2423 1347 -2421
rect 1346 -2429 1347 -2427
rect 1353 -2423 1354 -2421
rect 1353 -2429 1354 -2427
rect 1363 -2423 1364 -2421
rect 1360 -2429 1361 -2427
rect 1363 -2429 1364 -2427
rect 1367 -2423 1368 -2421
rect 1367 -2429 1368 -2427
rect 1374 -2423 1375 -2421
rect 1374 -2429 1375 -2427
rect 1381 -2423 1382 -2421
rect 1381 -2429 1382 -2427
rect 1384 -2429 1385 -2427
rect 1388 -2423 1389 -2421
rect 1388 -2429 1389 -2427
rect 1395 -2423 1396 -2421
rect 1395 -2429 1396 -2427
rect 1402 -2423 1403 -2421
rect 1402 -2429 1403 -2427
rect 1409 -2423 1410 -2421
rect 1409 -2429 1410 -2427
rect 1416 -2423 1417 -2421
rect 1416 -2429 1417 -2427
rect 1423 -2423 1424 -2421
rect 1423 -2429 1424 -2427
rect 1430 -2423 1431 -2421
rect 1430 -2429 1431 -2427
rect 1437 -2423 1438 -2421
rect 1437 -2429 1438 -2427
rect 1444 -2423 1445 -2421
rect 1444 -2429 1445 -2427
rect 1451 -2423 1452 -2421
rect 1451 -2429 1452 -2427
rect 1458 -2423 1459 -2421
rect 1458 -2429 1459 -2427
rect 1465 -2423 1466 -2421
rect 1465 -2429 1466 -2427
rect 1472 -2423 1473 -2421
rect 1472 -2429 1473 -2427
rect 1479 -2423 1480 -2421
rect 1479 -2429 1480 -2427
rect 1486 -2423 1487 -2421
rect 1486 -2429 1487 -2427
rect 1493 -2423 1494 -2421
rect 1493 -2429 1494 -2427
rect 1500 -2423 1501 -2421
rect 1500 -2429 1501 -2427
rect 1507 -2423 1508 -2421
rect 1507 -2429 1508 -2427
rect 1514 -2423 1515 -2421
rect 1514 -2429 1515 -2427
rect 1521 -2423 1522 -2421
rect 1521 -2429 1522 -2427
rect 1528 -2423 1529 -2421
rect 1528 -2429 1529 -2427
rect 1535 -2423 1536 -2421
rect 1535 -2429 1536 -2427
rect 1542 -2423 1543 -2421
rect 1542 -2429 1543 -2427
rect 1549 -2423 1550 -2421
rect 1549 -2429 1550 -2427
rect 1556 -2423 1557 -2421
rect 1556 -2429 1557 -2427
rect 1563 -2423 1564 -2421
rect 1563 -2429 1564 -2427
rect 1570 -2423 1571 -2421
rect 1570 -2429 1571 -2427
rect 1577 -2423 1578 -2421
rect 1577 -2429 1578 -2427
rect 1584 -2423 1585 -2421
rect 1584 -2429 1585 -2427
rect 1591 -2423 1592 -2421
rect 1591 -2429 1592 -2427
rect 1598 -2423 1599 -2421
rect 1598 -2429 1599 -2427
rect 1605 -2423 1606 -2421
rect 1605 -2429 1606 -2427
rect 1612 -2423 1613 -2421
rect 1612 -2429 1613 -2427
rect 1619 -2423 1620 -2421
rect 1622 -2423 1623 -2421
rect 1619 -2429 1620 -2427
rect 1622 -2429 1623 -2427
rect 1626 -2423 1627 -2421
rect 1626 -2429 1627 -2427
rect 1633 -2423 1634 -2421
rect 1633 -2429 1634 -2427
rect 1640 -2429 1641 -2427
rect 1643 -2429 1644 -2427
rect 1650 -2423 1651 -2421
rect 1647 -2429 1648 -2427
rect 1650 -2429 1651 -2427
rect 1654 -2423 1655 -2421
rect 1654 -2429 1655 -2427
rect 1661 -2423 1662 -2421
rect 1661 -2429 1662 -2427
rect 51 -2542 52 -2540
rect 51 -2548 52 -2546
rect 58 -2542 59 -2540
rect 58 -2548 59 -2546
rect 65 -2542 66 -2540
rect 65 -2548 66 -2546
rect 72 -2542 73 -2540
rect 72 -2548 73 -2546
rect 79 -2542 80 -2540
rect 79 -2548 80 -2546
rect 86 -2542 87 -2540
rect 89 -2542 90 -2540
rect 86 -2548 87 -2546
rect 89 -2548 90 -2546
rect 93 -2542 94 -2540
rect 93 -2548 94 -2546
rect 100 -2542 101 -2540
rect 100 -2548 101 -2546
rect 107 -2542 108 -2540
rect 107 -2548 108 -2546
rect 114 -2542 115 -2540
rect 114 -2548 115 -2546
rect 121 -2542 122 -2540
rect 121 -2548 122 -2546
rect 128 -2542 129 -2540
rect 128 -2548 129 -2546
rect 135 -2542 136 -2540
rect 135 -2548 136 -2546
rect 142 -2542 143 -2540
rect 142 -2548 143 -2546
rect 149 -2542 150 -2540
rect 149 -2548 150 -2546
rect 156 -2542 157 -2540
rect 156 -2548 157 -2546
rect 163 -2542 164 -2540
rect 163 -2548 164 -2546
rect 170 -2542 171 -2540
rect 173 -2542 174 -2540
rect 170 -2548 171 -2546
rect 177 -2542 178 -2540
rect 177 -2548 178 -2546
rect 184 -2542 185 -2540
rect 184 -2548 185 -2546
rect 191 -2542 192 -2540
rect 191 -2548 192 -2546
rect 198 -2542 199 -2540
rect 198 -2548 199 -2546
rect 205 -2542 206 -2540
rect 205 -2548 206 -2546
rect 212 -2542 213 -2540
rect 215 -2542 216 -2540
rect 212 -2548 213 -2546
rect 215 -2548 216 -2546
rect 219 -2542 220 -2540
rect 219 -2548 220 -2546
rect 226 -2542 227 -2540
rect 226 -2548 227 -2546
rect 233 -2542 234 -2540
rect 233 -2548 234 -2546
rect 240 -2542 241 -2540
rect 240 -2548 241 -2546
rect 247 -2542 248 -2540
rect 247 -2548 248 -2546
rect 254 -2542 255 -2540
rect 257 -2542 258 -2540
rect 254 -2548 255 -2546
rect 257 -2548 258 -2546
rect 261 -2542 262 -2540
rect 261 -2548 262 -2546
rect 268 -2542 269 -2540
rect 268 -2548 269 -2546
rect 275 -2542 276 -2540
rect 278 -2542 279 -2540
rect 275 -2548 276 -2546
rect 278 -2548 279 -2546
rect 282 -2542 283 -2540
rect 285 -2542 286 -2540
rect 282 -2548 283 -2546
rect 289 -2542 290 -2540
rect 289 -2548 290 -2546
rect 292 -2548 293 -2546
rect 296 -2542 297 -2540
rect 303 -2542 304 -2540
rect 303 -2548 304 -2546
rect 310 -2542 311 -2540
rect 310 -2548 311 -2546
rect 317 -2542 318 -2540
rect 317 -2548 318 -2546
rect 324 -2542 325 -2540
rect 324 -2548 325 -2546
rect 331 -2542 332 -2540
rect 331 -2548 332 -2546
rect 338 -2542 339 -2540
rect 338 -2548 339 -2546
rect 345 -2542 346 -2540
rect 345 -2548 346 -2546
rect 352 -2542 353 -2540
rect 352 -2548 353 -2546
rect 359 -2542 360 -2540
rect 359 -2548 360 -2546
rect 366 -2542 367 -2540
rect 366 -2548 367 -2546
rect 373 -2542 374 -2540
rect 373 -2548 374 -2546
rect 380 -2542 381 -2540
rect 380 -2548 381 -2546
rect 387 -2542 388 -2540
rect 390 -2542 391 -2540
rect 390 -2548 391 -2546
rect 394 -2542 395 -2540
rect 394 -2548 395 -2546
rect 401 -2542 402 -2540
rect 401 -2548 402 -2546
rect 408 -2542 409 -2540
rect 408 -2548 409 -2546
rect 415 -2548 416 -2546
rect 418 -2548 419 -2546
rect 422 -2542 423 -2540
rect 422 -2548 423 -2546
rect 429 -2542 430 -2540
rect 429 -2548 430 -2546
rect 436 -2542 437 -2540
rect 436 -2548 437 -2546
rect 443 -2542 444 -2540
rect 443 -2548 444 -2546
rect 450 -2542 451 -2540
rect 450 -2548 451 -2546
rect 457 -2542 458 -2540
rect 457 -2548 458 -2546
rect 464 -2542 465 -2540
rect 464 -2548 465 -2546
rect 471 -2542 472 -2540
rect 471 -2548 472 -2546
rect 478 -2542 479 -2540
rect 481 -2542 482 -2540
rect 481 -2548 482 -2546
rect 485 -2542 486 -2540
rect 485 -2548 486 -2546
rect 492 -2542 493 -2540
rect 492 -2548 493 -2546
rect 499 -2542 500 -2540
rect 499 -2548 500 -2546
rect 506 -2542 507 -2540
rect 506 -2548 507 -2546
rect 513 -2542 514 -2540
rect 513 -2548 514 -2546
rect 520 -2542 521 -2540
rect 520 -2548 521 -2546
rect 527 -2542 528 -2540
rect 530 -2542 531 -2540
rect 530 -2548 531 -2546
rect 534 -2542 535 -2540
rect 534 -2548 535 -2546
rect 541 -2542 542 -2540
rect 541 -2548 542 -2546
rect 544 -2548 545 -2546
rect 548 -2542 549 -2540
rect 548 -2548 549 -2546
rect 555 -2542 556 -2540
rect 555 -2548 556 -2546
rect 562 -2542 563 -2540
rect 565 -2542 566 -2540
rect 562 -2548 563 -2546
rect 565 -2548 566 -2546
rect 569 -2542 570 -2540
rect 572 -2542 573 -2540
rect 569 -2548 570 -2546
rect 572 -2548 573 -2546
rect 576 -2542 577 -2540
rect 576 -2548 577 -2546
rect 583 -2542 584 -2540
rect 583 -2548 584 -2546
rect 590 -2542 591 -2540
rect 590 -2548 591 -2546
rect 597 -2542 598 -2540
rect 600 -2542 601 -2540
rect 597 -2548 598 -2546
rect 600 -2548 601 -2546
rect 604 -2542 605 -2540
rect 604 -2548 605 -2546
rect 611 -2542 612 -2540
rect 611 -2548 612 -2546
rect 618 -2542 619 -2540
rect 618 -2548 619 -2546
rect 625 -2542 626 -2540
rect 625 -2548 626 -2546
rect 632 -2542 633 -2540
rect 632 -2548 633 -2546
rect 639 -2542 640 -2540
rect 639 -2548 640 -2546
rect 646 -2542 647 -2540
rect 646 -2548 647 -2546
rect 653 -2542 654 -2540
rect 653 -2548 654 -2546
rect 660 -2542 661 -2540
rect 660 -2548 661 -2546
rect 667 -2548 668 -2546
rect 670 -2548 671 -2546
rect 674 -2542 675 -2540
rect 674 -2548 675 -2546
rect 681 -2542 682 -2540
rect 681 -2548 682 -2546
rect 688 -2542 689 -2540
rect 688 -2548 689 -2546
rect 695 -2542 696 -2540
rect 695 -2548 696 -2546
rect 702 -2542 703 -2540
rect 702 -2548 703 -2546
rect 709 -2542 710 -2540
rect 709 -2548 710 -2546
rect 716 -2542 717 -2540
rect 716 -2548 717 -2546
rect 723 -2542 724 -2540
rect 723 -2548 724 -2546
rect 730 -2542 731 -2540
rect 730 -2548 731 -2546
rect 733 -2548 734 -2546
rect 737 -2542 738 -2540
rect 740 -2542 741 -2540
rect 737 -2548 738 -2546
rect 740 -2548 741 -2546
rect 744 -2542 745 -2540
rect 744 -2548 745 -2546
rect 747 -2548 748 -2546
rect 751 -2548 752 -2546
rect 754 -2548 755 -2546
rect 758 -2542 759 -2540
rect 758 -2548 759 -2546
rect 765 -2542 766 -2540
rect 765 -2548 766 -2546
rect 772 -2542 773 -2540
rect 772 -2548 773 -2546
rect 779 -2542 780 -2540
rect 779 -2548 780 -2546
rect 786 -2542 787 -2540
rect 786 -2548 787 -2546
rect 789 -2548 790 -2546
rect 793 -2542 794 -2540
rect 793 -2548 794 -2546
rect 800 -2542 801 -2540
rect 803 -2542 804 -2540
rect 800 -2548 801 -2546
rect 803 -2548 804 -2546
rect 807 -2542 808 -2540
rect 810 -2542 811 -2540
rect 810 -2548 811 -2546
rect 814 -2542 815 -2540
rect 814 -2548 815 -2546
rect 821 -2542 822 -2540
rect 821 -2548 822 -2546
rect 828 -2542 829 -2540
rect 831 -2542 832 -2540
rect 828 -2548 829 -2546
rect 831 -2548 832 -2546
rect 835 -2542 836 -2540
rect 835 -2548 836 -2546
rect 842 -2542 843 -2540
rect 842 -2548 843 -2546
rect 849 -2542 850 -2540
rect 849 -2548 850 -2546
rect 856 -2542 857 -2540
rect 856 -2548 857 -2546
rect 863 -2542 864 -2540
rect 863 -2548 864 -2546
rect 870 -2542 871 -2540
rect 870 -2548 871 -2546
rect 877 -2542 878 -2540
rect 877 -2548 878 -2546
rect 884 -2542 885 -2540
rect 884 -2548 885 -2546
rect 891 -2542 892 -2540
rect 891 -2548 892 -2546
rect 901 -2542 902 -2540
rect 898 -2548 899 -2546
rect 901 -2548 902 -2546
rect 905 -2542 906 -2540
rect 905 -2548 906 -2546
rect 912 -2542 913 -2540
rect 912 -2548 913 -2546
rect 919 -2542 920 -2540
rect 919 -2548 920 -2546
rect 926 -2542 927 -2540
rect 926 -2548 927 -2546
rect 933 -2542 934 -2540
rect 933 -2548 934 -2546
rect 940 -2542 941 -2540
rect 940 -2548 941 -2546
rect 947 -2542 948 -2540
rect 947 -2548 948 -2546
rect 954 -2542 955 -2540
rect 954 -2548 955 -2546
rect 961 -2542 962 -2540
rect 961 -2548 962 -2546
rect 968 -2542 969 -2540
rect 968 -2548 969 -2546
rect 975 -2542 976 -2540
rect 975 -2548 976 -2546
rect 982 -2542 983 -2540
rect 982 -2548 983 -2546
rect 989 -2542 990 -2540
rect 989 -2548 990 -2546
rect 996 -2542 997 -2540
rect 996 -2548 997 -2546
rect 1003 -2542 1004 -2540
rect 1003 -2548 1004 -2546
rect 1010 -2542 1011 -2540
rect 1013 -2542 1014 -2540
rect 1010 -2548 1011 -2546
rect 1017 -2542 1018 -2540
rect 1017 -2548 1018 -2546
rect 1024 -2542 1025 -2540
rect 1027 -2542 1028 -2540
rect 1031 -2542 1032 -2540
rect 1031 -2548 1032 -2546
rect 1038 -2542 1039 -2540
rect 1038 -2548 1039 -2546
rect 1045 -2542 1046 -2540
rect 1045 -2548 1046 -2546
rect 1052 -2542 1053 -2540
rect 1052 -2548 1053 -2546
rect 1059 -2542 1060 -2540
rect 1059 -2548 1060 -2546
rect 1066 -2542 1067 -2540
rect 1066 -2548 1067 -2546
rect 1073 -2542 1074 -2540
rect 1073 -2548 1074 -2546
rect 1080 -2542 1081 -2540
rect 1080 -2548 1081 -2546
rect 1087 -2542 1088 -2540
rect 1087 -2548 1088 -2546
rect 1094 -2542 1095 -2540
rect 1094 -2548 1095 -2546
rect 1101 -2542 1102 -2540
rect 1101 -2548 1102 -2546
rect 1108 -2542 1109 -2540
rect 1108 -2548 1109 -2546
rect 1115 -2542 1116 -2540
rect 1115 -2548 1116 -2546
rect 1122 -2542 1123 -2540
rect 1122 -2548 1123 -2546
rect 1129 -2542 1130 -2540
rect 1129 -2548 1130 -2546
rect 1136 -2542 1137 -2540
rect 1136 -2548 1137 -2546
rect 1146 -2542 1147 -2540
rect 1143 -2548 1144 -2546
rect 1146 -2548 1147 -2546
rect 1150 -2542 1151 -2540
rect 1150 -2548 1151 -2546
rect 1157 -2542 1158 -2540
rect 1157 -2548 1158 -2546
rect 1164 -2542 1165 -2540
rect 1164 -2548 1165 -2546
rect 1171 -2542 1172 -2540
rect 1171 -2548 1172 -2546
rect 1178 -2542 1179 -2540
rect 1178 -2548 1179 -2546
rect 1185 -2542 1186 -2540
rect 1185 -2548 1186 -2546
rect 1192 -2542 1193 -2540
rect 1192 -2548 1193 -2546
rect 1199 -2542 1200 -2540
rect 1199 -2548 1200 -2546
rect 1206 -2542 1207 -2540
rect 1206 -2548 1207 -2546
rect 1213 -2542 1214 -2540
rect 1213 -2548 1214 -2546
rect 1220 -2542 1221 -2540
rect 1220 -2548 1221 -2546
rect 1227 -2542 1228 -2540
rect 1227 -2548 1228 -2546
rect 1234 -2542 1235 -2540
rect 1234 -2548 1235 -2546
rect 1241 -2542 1242 -2540
rect 1241 -2548 1242 -2546
rect 1248 -2542 1249 -2540
rect 1251 -2542 1252 -2540
rect 1248 -2548 1249 -2546
rect 1251 -2548 1252 -2546
rect 1255 -2542 1256 -2540
rect 1255 -2548 1256 -2546
rect 1262 -2542 1263 -2540
rect 1262 -2548 1263 -2546
rect 1269 -2542 1270 -2540
rect 1269 -2548 1270 -2546
rect 1276 -2542 1277 -2540
rect 1276 -2548 1277 -2546
rect 1283 -2542 1284 -2540
rect 1283 -2548 1284 -2546
rect 1290 -2542 1291 -2540
rect 1290 -2548 1291 -2546
rect 1297 -2542 1298 -2540
rect 1297 -2548 1298 -2546
rect 1304 -2542 1305 -2540
rect 1304 -2548 1305 -2546
rect 1311 -2542 1312 -2540
rect 1311 -2548 1312 -2546
rect 1318 -2542 1319 -2540
rect 1318 -2548 1319 -2546
rect 1325 -2542 1326 -2540
rect 1325 -2548 1326 -2546
rect 1332 -2542 1333 -2540
rect 1332 -2548 1333 -2546
rect 1339 -2542 1340 -2540
rect 1339 -2548 1340 -2546
rect 1346 -2542 1347 -2540
rect 1346 -2548 1347 -2546
rect 1353 -2542 1354 -2540
rect 1353 -2548 1354 -2546
rect 1360 -2542 1361 -2540
rect 1360 -2548 1361 -2546
rect 1367 -2542 1368 -2540
rect 1367 -2548 1368 -2546
rect 1374 -2542 1375 -2540
rect 1374 -2548 1375 -2546
rect 1381 -2542 1382 -2540
rect 1381 -2548 1382 -2546
rect 1388 -2542 1389 -2540
rect 1388 -2548 1389 -2546
rect 1395 -2542 1396 -2540
rect 1395 -2548 1396 -2546
rect 1405 -2542 1406 -2540
rect 1405 -2548 1406 -2546
rect 1409 -2542 1410 -2540
rect 1409 -2548 1410 -2546
rect 1416 -2542 1417 -2540
rect 1416 -2548 1417 -2546
rect 1423 -2542 1424 -2540
rect 1423 -2548 1424 -2546
rect 1430 -2542 1431 -2540
rect 1430 -2548 1431 -2546
rect 1437 -2542 1438 -2540
rect 1437 -2548 1438 -2546
rect 1444 -2542 1445 -2540
rect 1444 -2548 1445 -2546
rect 1451 -2542 1452 -2540
rect 1451 -2548 1452 -2546
rect 1458 -2542 1459 -2540
rect 1458 -2548 1459 -2546
rect 1465 -2542 1466 -2540
rect 1465 -2548 1466 -2546
rect 1472 -2542 1473 -2540
rect 1472 -2548 1473 -2546
rect 1479 -2542 1480 -2540
rect 1479 -2548 1480 -2546
rect 1486 -2542 1487 -2540
rect 1486 -2548 1487 -2546
rect 1493 -2542 1494 -2540
rect 1493 -2548 1494 -2546
rect 1500 -2542 1501 -2540
rect 1500 -2548 1501 -2546
rect 1507 -2542 1508 -2540
rect 1507 -2548 1508 -2546
rect 1514 -2542 1515 -2540
rect 1514 -2548 1515 -2546
rect 1521 -2542 1522 -2540
rect 1521 -2548 1522 -2546
rect 1528 -2542 1529 -2540
rect 1528 -2548 1529 -2546
rect 1535 -2542 1536 -2540
rect 1535 -2548 1536 -2546
rect 1542 -2542 1543 -2540
rect 1542 -2548 1543 -2546
rect 1549 -2542 1550 -2540
rect 1549 -2548 1550 -2546
rect 1556 -2542 1557 -2540
rect 1556 -2548 1557 -2546
rect 1563 -2542 1564 -2540
rect 1563 -2548 1564 -2546
rect 1570 -2542 1571 -2540
rect 1570 -2548 1571 -2546
rect 1577 -2542 1578 -2540
rect 1577 -2548 1578 -2546
rect 1587 -2542 1588 -2540
rect 1584 -2548 1585 -2546
rect 1587 -2548 1588 -2546
rect 1591 -2542 1592 -2540
rect 1591 -2548 1592 -2546
rect 1598 -2542 1599 -2540
rect 1598 -2548 1599 -2546
rect 1605 -2542 1606 -2540
rect 1605 -2548 1606 -2546
rect 1612 -2542 1613 -2540
rect 1615 -2542 1616 -2540
rect 1612 -2548 1613 -2546
rect 1615 -2548 1616 -2546
rect 1640 -2542 1641 -2540
rect 1640 -2548 1641 -2546
rect 44 -2671 45 -2669
rect 44 -2677 45 -2675
rect 51 -2671 52 -2669
rect 51 -2677 52 -2675
rect 58 -2671 59 -2669
rect 58 -2677 59 -2675
rect 65 -2671 66 -2669
rect 65 -2677 66 -2675
rect 72 -2671 73 -2669
rect 72 -2677 73 -2675
rect 79 -2671 80 -2669
rect 79 -2677 80 -2675
rect 86 -2671 87 -2669
rect 86 -2677 87 -2675
rect 93 -2671 94 -2669
rect 93 -2677 94 -2675
rect 100 -2671 101 -2669
rect 100 -2677 101 -2675
rect 107 -2671 108 -2669
rect 107 -2677 108 -2675
rect 114 -2671 115 -2669
rect 114 -2677 115 -2675
rect 121 -2671 122 -2669
rect 121 -2677 122 -2675
rect 131 -2671 132 -2669
rect 128 -2677 129 -2675
rect 131 -2677 132 -2675
rect 135 -2671 136 -2669
rect 135 -2677 136 -2675
rect 142 -2671 143 -2669
rect 142 -2677 143 -2675
rect 149 -2671 150 -2669
rect 152 -2671 153 -2669
rect 149 -2677 150 -2675
rect 152 -2677 153 -2675
rect 156 -2671 157 -2669
rect 156 -2677 157 -2675
rect 163 -2671 164 -2669
rect 163 -2677 164 -2675
rect 170 -2671 171 -2669
rect 170 -2677 171 -2675
rect 180 -2671 181 -2669
rect 177 -2677 178 -2675
rect 184 -2671 185 -2669
rect 184 -2677 185 -2675
rect 191 -2671 192 -2669
rect 191 -2677 192 -2675
rect 201 -2671 202 -2669
rect 198 -2677 199 -2675
rect 201 -2677 202 -2675
rect 205 -2671 206 -2669
rect 208 -2671 209 -2669
rect 205 -2677 206 -2675
rect 208 -2677 209 -2675
rect 212 -2671 213 -2669
rect 212 -2677 213 -2675
rect 219 -2671 220 -2669
rect 219 -2677 220 -2675
rect 226 -2671 227 -2669
rect 226 -2677 227 -2675
rect 233 -2671 234 -2669
rect 236 -2671 237 -2669
rect 233 -2677 234 -2675
rect 236 -2677 237 -2675
rect 240 -2671 241 -2669
rect 240 -2677 241 -2675
rect 247 -2671 248 -2669
rect 247 -2677 248 -2675
rect 254 -2671 255 -2669
rect 254 -2677 255 -2675
rect 261 -2671 262 -2669
rect 264 -2671 265 -2669
rect 264 -2677 265 -2675
rect 268 -2671 269 -2669
rect 268 -2677 269 -2675
rect 275 -2671 276 -2669
rect 275 -2677 276 -2675
rect 282 -2671 283 -2669
rect 282 -2677 283 -2675
rect 289 -2671 290 -2669
rect 289 -2677 290 -2675
rect 296 -2671 297 -2669
rect 296 -2677 297 -2675
rect 303 -2671 304 -2669
rect 303 -2677 304 -2675
rect 310 -2671 311 -2669
rect 310 -2677 311 -2675
rect 317 -2671 318 -2669
rect 317 -2677 318 -2675
rect 324 -2671 325 -2669
rect 324 -2677 325 -2675
rect 331 -2671 332 -2669
rect 331 -2677 332 -2675
rect 338 -2671 339 -2669
rect 338 -2677 339 -2675
rect 345 -2671 346 -2669
rect 345 -2677 346 -2675
rect 352 -2671 353 -2669
rect 352 -2677 353 -2675
rect 359 -2671 360 -2669
rect 359 -2677 360 -2675
rect 366 -2671 367 -2669
rect 366 -2677 367 -2675
rect 376 -2671 377 -2669
rect 373 -2677 374 -2675
rect 380 -2671 381 -2669
rect 380 -2677 381 -2675
rect 387 -2671 388 -2669
rect 387 -2677 388 -2675
rect 394 -2677 395 -2675
rect 397 -2677 398 -2675
rect 401 -2671 402 -2669
rect 401 -2677 402 -2675
rect 408 -2671 409 -2669
rect 408 -2677 409 -2675
rect 415 -2671 416 -2669
rect 415 -2677 416 -2675
rect 422 -2671 423 -2669
rect 425 -2671 426 -2669
rect 422 -2677 423 -2675
rect 425 -2677 426 -2675
rect 429 -2671 430 -2669
rect 429 -2677 430 -2675
rect 436 -2671 437 -2669
rect 436 -2677 437 -2675
rect 443 -2671 444 -2669
rect 443 -2677 444 -2675
rect 450 -2671 451 -2669
rect 450 -2677 451 -2675
rect 457 -2671 458 -2669
rect 457 -2677 458 -2675
rect 464 -2671 465 -2669
rect 464 -2677 465 -2675
rect 471 -2671 472 -2669
rect 471 -2677 472 -2675
rect 478 -2671 479 -2669
rect 478 -2677 479 -2675
rect 485 -2671 486 -2669
rect 485 -2677 486 -2675
rect 492 -2671 493 -2669
rect 492 -2677 493 -2675
rect 499 -2671 500 -2669
rect 502 -2671 503 -2669
rect 499 -2677 500 -2675
rect 506 -2671 507 -2669
rect 506 -2677 507 -2675
rect 513 -2671 514 -2669
rect 513 -2677 514 -2675
rect 520 -2671 521 -2669
rect 520 -2677 521 -2675
rect 527 -2671 528 -2669
rect 527 -2677 528 -2675
rect 534 -2671 535 -2669
rect 534 -2677 535 -2675
rect 541 -2671 542 -2669
rect 541 -2677 542 -2675
rect 548 -2671 549 -2669
rect 548 -2677 549 -2675
rect 555 -2671 556 -2669
rect 555 -2677 556 -2675
rect 562 -2671 563 -2669
rect 562 -2677 563 -2675
rect 569 -2671 570 -2669
rect 569 -2677 570 -2675
rect 576 -2671 577 -2669
rect 576 -2677 577 -2675
rect 583 -2671 584 -2669
rect 583 -2677 584 -2675
rect 590 -2671 591 -2669
rect 590 -2677 591 -2675
rect 597 -2671 598 -2669
rect 597 -2677 598 -2675
rect 604 -2671 605 -2669
rect 604 -2677 605 -2675
rect 611 -2671 612 -2669
rect 614 -2671 615 -2669
rect 611 -2677 612 -2675
rect 614 -2677 615 -2675
rect 618 -2671 619 -2669
rect 618 -2677 619 -2675
rect 625 -2671 626 -2669
rect 625 -2677 626 -2675
rect 632 -2671 633 -2669
rect 632 -2677 633 -2675
rect 639 -2671 640 -2669
rect 639 -2677 640 -2675
rect 646 -2671 647 -2669
rect 649 -2677 650 -2675
rect 653 -2671 654 -2669
rect 656 -2671 657 -2669
rect 653 -2677 654 -2675
rect 656 -2677 657 -2675
rect 660 -2671 661 -2669
rect 660 -2677 661 -2675
rect 667 -2671 668 -2669
rect 667 -2677 668 -2675
rect 674 -2671 675 -2669
rect 674 -2677 675 -2675
rect 681 -2671 682 -2669
rect 681 -2677 682 -2675
rect 688 -2671 689 -2669
rect 688 -2677 689 -2675
rect 695 -2671 696 -2669
rect 695 -2677 696 -2675
rect 702 -2671 703 -2669
rect 702 -2677 703 -2675
rect 709 -2671 710 -2669
rect 709 -2677 710 -2675
rect 719 -2671 720 -2669
rect 723 -2671 724 -2669
rect 723 -2677 724 -2675
rect 730 -2671 731 -2669
rect 733 -2671 734 -2669
rect 733 -2677 734 -2675
rect 737 -2671 738 -2669
rect 737 -2677 738 -2675
rect 744 -2671 745 -2669
rect 744 -2677 745 -2675
rect 751 -2671 752 -2669
rect 751 -2677 752 -2675
rect 758 -2671 759 -2669
rect 758 -2677 759 -2675
rect 765 -2671 766 -2669
rect 765 -2677 766 -2675
rect 772 -2671 773 -2669
rect 772 -2677 773 -2675
rect 779 -2671 780 -2669
rect 779 -2677 780 -2675
rect 786 -2671 787 -2669
rect 786 -2677 787 -2675
rect 793 -2671 794 -2669
rect 793 -2677 794 -2675
rect 803 -2671 804 -2669
rect 800 -2677 801 -2675
rect 803 -2677 804 -2675
rect 807 -2671 808 -2669
rect 807 -2677 808 -2675
rect 814 -2671 815 -2669
rect 814 -2677 815 -2675
rect 821 -2671 822 -2669
rect 821 -2677 822 -2675
rect 828 -2671 829 -2669
rect 828 -2677 829 -2675
rect 835 -2671 836 -2669
rect 835 -2677 836 -2675
rect 842 -2671 843 -2669
rect 842 -2677 843 -2675
rect 849 -2671 850 -2669
rect 849 -2677 850 -2675
rect 859 -2671 860 -2669
rect 856 -2677 857 -2675
rect 859 -2677 860 -2675
rect 863 -2671 864 -2669
rect 863 -2677 864 -2675
rect 870 -2671 871 -2669
rect 870 -2677 871 -2675
rect 877 -2671 878 -2669
rect 880 -2671 881 -2669
rect 877 -2677 878 -2675
rect 880 -2677 881 -2675
rect 884 -2671 885 -2669
rect 887 -2671 888 -2669
rect 884 -2677 885 -2675
rect 887 -2677 888 -2675
rect 891 -2671 892 -2669
rect 891 -2677 892 -2675
rect 898 -2671 899 -2669
rect 901 -2671 902 -2669
rect 898 -2677 899 -2675
rect 901 -2677 902 -2675
rect 905 -2671 906 -2669
rect 905 -2677 906 -2675
rect 912 -2671 913 -2669
rect 912 -2677 913 -2675
rect 919 -2671 920 -2669
rect 919 -2677 920 -2675
rect 926 -2671 927 -2669
rect 926 -2677 927 -2675
rect 933 -2671 934 -2669
rect 933 -2677 934 -2675
rect 940 -2671 941 -2669
rect 940 -2677 941 -2675
rect 947 -2671 948 -2669
rect 950 -2671 951 -2669
rect 947 -2677 948 -2675
rect 950 -2677 951 -2675
rect 954 -2671 955 -2669
rect 957 -2671 958 -2669
rect 954 -2677 955 -2675
rect 957 -2677 958 -2675
rect 961 -2671 962 -2669
rect 961 -2677 962 -2675
rect 968 -2671 969 -2669
rect 971 -2671 972 -2669
rect 971 -2677 972 -2675
rect 975 -2671 976 -2669
rect 978 -2671 979 -2669
rect 975 -2677 976 -2675
rect 978 -2677 979 -2675
rect 982 -2671 983 -2669
rect 982 -2677 983 -2675
rect 989 -2671 990 -2669
rect 989 -2677 990 -2675
rect 996 -2671 997 -2669
rect 996 -2677 997 -2675
rect 1003 -2671 1004 -2669
rect 1003 -2677 1004 -2675
rect 1010 -2671 1011 -2669
rect 1010 -2677 1011 -2675
rect 1017 -2671 1018 -2669
rect 1017 -2677 1018 -2675
rect 1024 -2671 1025 -2669
rect 1027 -2671 1028 -2669
rect 1024 -2677 1025 -2675
rect 1031 -2671 1032 -2669
rect 1031 -2677 1032 -2675
rect 1038 -2671 1039 -2669
rect 1038 -2677 1039 -2675
rect 1045 -2671 1046 -2669
rect 1045 -2677 1046 -2675
rect 1052 -2671 1053 -2669
rect 1052 -2677 1053 -2675
rect 1059 -2671 1060 -2669
rect 1059 -2677 1060 -2675
rect 1066 -2671 1067 -2669
rect 1066 -2677 1067 -2675
rect 1073 -2671 1074 -2669
rect 1073 -2677 1074 -2675
rect 1080 -2671 1081 -2669
rect 1080 -2677 1081 -2675
rect 1087 -2671 1088 -2669
rect 1090 -2671 1091 -2669
rect 1090 -2677 1091 -2675
rect 1094 -2671 1095 -2669
rect 1094 -2677 1095 -2675
rect 1101 -2671 1102 -2669
rect 1101 -2677 1102 -2675
rect 1108 -2671 1109 -2669
rect 1108 -2677 1109 -2675
rect 1115 -2671 1116 -2669
rect 1115 -2677 1116 -2675
rect 1122 -2671 1123 -2669
rect 1122 -2677 1123 -2675
rect 1129 -2671 1130 -2669
rect 1129 -2677 1130 -2675
rect 1136 -2671 1137 -2669
rect 1136 -2677 1137 -2675
rect 1143 -2671 1144 -2669
rect 1143 -2677 1144 -2675
rect 1150 -2671 1151 -2669
rect 1153 -2671 1154 -2669
rect 1150 -2677 1151 -2675
rect 1153 -2677 1154 -2675
rect 1157 -2671 1158 -2669
rect 1157 -2677 1158 -2675
rect 1164 -2671 1165 -2669
rect 1164 -2677 1165 -2675
rect 1171 -2671 1172 -2669
rect 1171 -2677 1172 -2675
rect 1178 -2671 1179 -2669
rect 1178 -2677 1179 -2675
rect 1185 -2671 1186 -2669
rect 1188 -2671 1189 -2669
rect 1185 -2677 1186 -2675
rect 1188 -2677 1189 -2675
rect 1192 -2671 1193 -2669
rect 1192 -2677 1193 -2675
rect 1199 -2671 1200 -2669
rect 1199 -2677 1200 -2675
rect 1206 -2671 1207 -2669
rect 1206 -2677 1207 -2675
rect 1213 -2671 1214 -2669
rect 1213 -2677 1214 -2675
rect 1220 -2671 1221 -2669
rect 1220 -2677 1221 -2675
rect 1227 -2671 1228 -2669
rect 1227 -2677 1228 -2675
rect 1234 -2671 1235 -2669
rect 1234 -2677 1235 -2675
rect 1241 -2671 1242 -2669
rect 1241 -2677 1242 -2675
rect 1248 -2671 1249 -2669
rect 1248 -2677 1249 -2675
rect 1255 -2671 1256 -2669
rect 1255 -2677 1256 -2675
rect 1262 -2671 1263 -2669
rect 1262 -2677 1263 -2675
rect 1269 -2671 1270 -2669
rect 1269 -2677 1270 -2675
rect 1276 -2671 1277 -2669
rect 1276 -2677 1277 -2675
rect 1283 -2671 1284 -2669
rect 1283 -2677 1284 -2675
rect 1290 -2671 1291 -2669
rect 1290 -2677 1291 -2675
rect 1297 -2671 1298 -2669
rect 1297 -2677 1298 -2675
rect 1304 -2671 1305 -2669
rect 1304 -2677 1305 -2675
rect 1311 -2671 1312 -2669
rect 1311 -2677 1312 -2675
rect 1318 -2671 1319 -2669
rect 1318 -2677 1319 -2675
rect 1325 -2671 1326 -2669
rect 1325 -2677 1326 -2675
rect 1332 -2671 1333 -2669
rect 1332 -2677 1333 -2675
rect 1339 -2671 1340 -2669
rect 1339 -2677 1340 -2675
rect 1346 -2671 1347 -2669
rect 1346 -2677 1347 -2675
rect 1353 -2671 1354 -2669
rect 1353 -2677 1354 -2675
rect 1360 -2671 1361 -2669
rect 1360 -2677 1361 -2675
rect 1367 -2671 1368 -2669
rect 1367 -2677 1368 -2675
rect 1374 -2671 1375 -2669
rect 1374 -2677 1375 -2675
rect 1381 -2671 1382 -2669
rect 1381 -2677 1382 -2675
rect 1388 -2671 1389 -2669
rect 1388 -2677 1389 -2675
rect 1395 -2671 1396 -2669
rect 1395 -2677 1396 -2675
rect 1402 -2671 1403 -2669
rect 1402 -2677 1403 -2675
rect 1409 -2671 1410 -2669
rect 1409 -2677 1410 -2675
rect 1416 -2671 1417 -2669
rect 1416 -2677 1417 -2675
rect 1423 -2671 1424 -2669
rect 1423 -2677 1424 -2675
rect 1430 -2671 1431 -2669
rect 1430 -2677 1431 -2675
rect 1437 -2671 1438 -2669
rect 1437 -2677 1438 -2675
rect 1444 -2671 1445 -2669
rect 1444 -2677 1445 -2675
rect 1451 -2671 1452 -2669
rect 1451 -2677 1452 -2675
rect 1458 -2671 1459 -2669
rect 1458 -2677 1459 -2675
rect 1465 -2671 1466 -2669
rect 1465 -2677 1466 -2675
rect 1472 -2671 1473 -2669
rect 1472 -2677 1473 -2675
rect 1479 -2671 1480 -2669
rect 1479 -2677 1480 -2675
rect 1486 -2671 1487 -2669
rect 1486 -2677 1487 -2675
rect 1493 -2671 1494 -2669
rect 1493 -2677 1494 -2675
rect 1500 -2671 1501 -2669
rect 1500 -2677 1501 -2675
rect 1507 -2671 1508 -2669
rect 1507 -2677 1508 -2675
rect 1514 -2671 1515 -2669
rect 1514 -2677 1515 -2675
rect 1521 -2671 1522 -2669
rect 1521 -2677 1522 -2675
rect 1528 -2671 1529 -2669
rect 1528 -2677 1529 -2675
rect 1535 -2671 1536 -2669
rect 1535 -2677 1536 -2675
rect 1542 -2671 1543 -2669
rect 1542 -2677 1543 -2675
rect 1549 -2671 1550 -2669
rect 1549 -2677 1550 -2675
rect 1556 -2671 1557 -2669
rect 1556 -2677 1557 -2675
rect 1563 -2671 1564 -2669
rect 1563 -2677 1564 -2675
rect 1570 -2671 1571 -2669
rect 1570 -2677 1571 -2675
rect 1577 -2671 1578 -2669
rect 1577 -2677 1578 -2675
rect 1584 -2671 1585 -2669
rect 1584 -2677 1585 -2675
rect 1591 -2671 1592 -2669
rect 1591 -2677 1592 -2675
rect 1598 -2671 1599 -2669
rect 1598 -2677 1599 -2675
rect 1605 -2671 1606 -2669
rect 1605 -2677 1606 -2675
rect 1612 -2671 1613 -2669
rect 1612 -2677 1613 -2675
rect 1619 -2671 1620 -2669
rect 1619 -2677 1620 -2675
rect 1626 -2671 1627 -2669
rect 1629 -2671 1630 -2669
rect 1626 -2677 1627 -2675
rect 1629 -2677 1630 -2675
rect 1636 -2671 1637 -2669
rect 1633 -2677 1634 -2675
rect 1636 -2677 1637 -2675
rect 44 -2784 45 -2782
rect 44 -2790 45 -2788
rect 58 -2784 59 -2782
rect 58 -2790 59 -2788
rect 65 -2784 66 -2782
rect 65 -2790 66 -2788
rect 72 -2784 73 -2782
rect 72 -2790 73 -2788
rect 79 -2784 80 -2782
rect 79 -2790 80 -2788
rect 86 -2784 87 -2782
rect 86 -2790 87 -2788
rect 93 -2784 94 -2782
rect 93 -2790 94 -2788
rect 100 -2784 101 -2782
rect 100 -2790 101 -2788
rect 107 -2784 108 -2782
rect 107 -2790 108 -2788
rect 110 -2790 111 -2788
rect 114 -2784 115 -2782
rect 114 -2790 115 -2788
rect 121 -2784 122 -2782
rect 124 -2784 125 -2782
rect 121 -2790 122 -2788
rect 124 -2790 125 -2788
rect 128 -2784 129 -2782
rect 131 -2784 132 -2782
rect 128 -2790 129 -2788
rect 135 -2784 136 -2782
rect 138 -2784 139 -2782
rect 135 -2790 136 -2788
rect 138 -2790 139 -2788
rect 142 -2784 143 -2782
rect 142 -2790 143 -2788
rect 149 -2784 150 -2782
rect 149 -2790 150 -2788
rect 156 -2784 157 -2782
rect 159 -2784 160 -2782
rect 159 -2790 160 -2788
rect 163 -2784 164 -2782
rect 163 -2790 164 -2788
rect 170 -2784 171 -2782
rect 170 -2790 171 -2788
rect 177 -2784 178 -2782
rect 177 -2790 178 -2788
rect 184 -2784 185 -2782
rect 184 -2790 185 -2788
rect 191 -2784 192 -2782
rect 191 -2790 192 -2788
rect 198 -2784 199 -2782
rect 198 -2790 199 -2788
rect 205 -2784 206 -2782
rect 205 -2790 206 -2788
rect 212 -2784 213 -2782
rect 215 -2784 216 -2782
rect 212 -2790 213 -2788
rect 215 -2790 216 -2788
rect 219 -2784 220 -2782
rect 219 -2790 220 -2788
rect 226 -2784 227 -2782
rect 226 -2790 227 -2788
rect 233 -2790 234 -2788
rect 236 -2790 237 -2788
rect 240 -2784 241 -2782
rect 240 -2790 241 -2788
rect 247 -2784 248 -2782
rect 247 -2790 248 -2788
rect 254 -2784 255 -2782
rect 254 -2790 255 -2788
rect 261 -2784 262 -2782
rect 264 -2784 265 -2782
rect 264 -2790 265 -2788
rect 268 -2784 269 -2782
rect 268 -2790 269 -2788
rect 275 -2784 276 -2782
rect 275 -2790 276 -2788
rect 282 -2790 283 -2788
rect 289 -2784 290 -2782
rect 292 -2784 293 -2782
rect 292 -2790 293 -2788
rect 296 -2784 297 -2782
rect 296 -2790 297 -2788
rect 303 -2784 304 -2782
rect 303 -2790 304 -2788
rect 310 -2784 311 -2782
rect 310 -2790 311 -2788
rect 317 -2784 318 -2782
rect 317 -2790 318 -2788
rect 324 -2784 325 -2782
rect 324 -2790 325 -2788
rect 331 -2784 332 -2782
rect 331 -2790 332 -2788
rect 338 -2784 339 -2782
rect 338 -2790 339 -2788
rect 345 -2784 346 -2782
rect 345 -2790 346 -2788
rect 352 -2784 353 -2782
rect 352 -2790 353 -2788
rect 359 -2784 360 -2782
rect 359 -2790 360 -2788
rect 366 -2784 367 -2782
rect 366 -2790 367 -2788
rect 373 -2784 374 -2782
rect 373 -2790 374 -2788
rect 380 -2784 381 -2782
rect 380 -2790 381 -2788
rect 387 -2784 388 -2782
rect 387 -2790 388 -2788
rect 394 -2784 395 -2782
rect 394 -2790 395 -2788
rect 401 -2784 402 -2782
rect 401 -2790 402 -2788
rect 408 -2784 409 -2782
rect 408 -2790 409 -2788
rect 415 -2784 416 -2782
rect 415 -2790 416 -2788
rect 422 -2784 423 -2782
rect 422 -2790 423 -2788
rect 429 -2784 430 -2782
rect 429 -2790 430 -2788
rect 436 -2784 437 -2782
rect 436 -2790 437 -2788
rect 446 -2784 447 -2782
rect 443 -2790 444 -2788
rect 446 -2790 447 -2788
rect 450 -2784 451 -2782
rect 450 -2790 451 -2788
rect 457 -2784 458 -2782
rect 457 -2790 458 -2788
rect 464 -2784 465 -2782
rect 464 -2790 465 -2788
rect 471 -2784 472 -2782
rect 471 -2790 472 -2788
rect 478 -2784 479 -2782
rect 485 -2784 486 -2782
rect 485 -2790 486 -2788
rect 492 -2784 493 -2782
rect 492 -2790 493 -2788
rect 499 -2784 500 -2782
rect 499 -2790 500 -2788
rect 506 -2784 507 -2782
rect 506 -2790 507 -2788
rect 513 -2784 514 -2782
rect 513 -2790 514 -2788
rect 520 -2784 521 -2782
rect 520 -2790 521 -2788
rect 527 -2784 528 -2782
rect 527 -2790 528 -2788
rect 534 -2784 535 -2782
rect 534 -2790 535 -2788
rect 541 -2784 542 -2782
rect 541 -2790 542 -2788
rect 548 -2784 549 -2782
rect 548 -2790 549 -2788
rect 555 -2784 556 -2782
rect 555 -2790 556 -2788
rect 562 -2784 563 -2782
rect 565 -2784 566 -2782
rect 562 -2790 563 -2788
rect 565 -2790 566 -2788
rect 569 -2784 570 -2782
rect 569 -2790 570 -2788
rect 576 -2784 577 -2782
rect 576 -2790 577 -2788
rect 583 -2784 584 -2782
rect 583 -2790 584 -2788
rect 590 -2790 591 -2788
rect 593 -2790 594 -2788
rect 597 -2784 598 -2782
rect 597 -2790 598 -2788
rect 604 -2784 605 -2782
rect 604 -2790 605 -2788
rect 611 -2784 612 -2782
rect 611 -2790 612 -2788
rect 618 -2784 619 -2782
rect 618 -2790 619 -2788
rect 625 -2784 626 -2782
rect 625 -2790 626 -2788
rect 632 -2784 633 -2782
rect 632 -2790 633 -2788
rect 639 -2784 640 -2782
rect 639 -2790 640 -2788
rect 646 -2784 647 -2782
rect 646 -2790 647 -2788
rect 653 -2784 654 -2782
rect 653 -2790 654 -2788
rect 660 -2784 661 -2782
rect 663 -2784 664 -2782
rect 660 -2790 661 -2788
rect 663 -2790 664 -2788
rect 667 -2784 668 -2782
rect 667 -2790 668 -2788
rect 670 -2790 671 -2788
rect 674 -2784 675 -2782
rect 677 -2784 678 -2782
rect 677 -2790 678 -2788
rect 681 -2784 682 -2782
rect 681 -2790 682 -2788
rect 691 -2784 692 -2782
rect 688 -2790 689 -2788
rect 695 -2784 696 -2782
rect 695 -2790 696 -2788
rect 702 -2784 703 -2782
rect 702 -2790 703 -2788
rect 709 -2784 710 -2782
rect 709 -2790 710 -2788
rect 716 -2784 717 -2782
rect 716 -2790 717 -2788
rect 723 -2784 724 -2782
rect 723 -2790 724 -2788
rect 730 -2784 731 -2782
rect 730 -2790 731 -2788
rect 737 -2784 738 -2782
rect 737 -2790 738 -2788
rect 744 -2784 745 -2782
rect 747 -2784 748 -2782
rect 744 -2790 745 -2788
rect 747 -2790 748 -2788
rect 751 -2784 752 -2782
rect 751 -2790 752 -2788
rect 758 -2784 759 -2782
rect 761 -2784 762 -2782
rect 761 -2790 762 -2788
rect 765 -2784 766 -2782
rect 765 -2790 766 -2788
rect 772 -2784 773 -2782
rect 772 -2790 773 -2788
rect 779 -2784 780 -2782
rect 782 -2784 783 -2782
rect 779 -2790 780 -2788
rect 786 -2784 787 -2782
rect 786 -2790 787 -2788
rect 789 -2790 790 -2788
rect 793 -2784 794 -2782
rect 793 -2790 794 -2788
rect 800 -2784 801 -2782
rect 800 -2790 801 -2788
rect 807 -2790 808 -2788
rect 810 -2790 811 -2788
rect 814 -2784 815 -2782
rect 817 -2784 818 -2782
rect 814 -2790 815 -2788
rect 817 -2790 818 -2788
rect 821 -2784 822 -2782
rect 821 -2790 822 -2788
rect 828 -2784 829 -2782
rect 828 -2790 829 -2788
rect 835 -2784 836 -2782
rect 835 -2790 836 -2788
rect 842 -2784 843 -2782
rect 845 -2784 846 -2782
rect 842 -2790 843 -2788
rect 845 -2790 846 -2788
rect 849 -2784 850 -2782
rect 849 -2790 850 -2788
rect 856 -2784 857 -2782
rect 856 -2790 857 -2788
rect 863 -2784 864 -2782
rect 863 -2790 864 -2788
rect 870 -2784 871 -2782
rect 870 -2790 871 -2788
rect 877 -2784 878 -2782
rect 880 -2784 881 -2782
rect 877 -2790 878 -2788
rect 880 -2790 881 -2788
rect 884 -2784 885 -2782
rect 884 -2790 885 -2788
rect 891 -2784 892 -2782
rect 891 -2790 892 -2788
rect 898 -2784 899 -2782
rect 898 -2790 899 -2788
rect 905 -2784 906 -2782
rect 908 -2784 909 -2782
rect 905 -2790 906 -2788
rect 908 -2790 909 -2788
rect 912 -2784 913 -2782
rect 912 -2790 913 -2788
rect 919 -2784 920 -2782
rect 919 -2790 920 -2788
rect 926 -2784 927 -2782
rect 926 -2790 927 -2788
rect 933 -2784 934 -2782
rect 933 -2790 934 -2788
rect 940 -2784 941 -2782
rect 940 -2790 941 -2788
rect 947 -2784 948 -2782
rect 947 -2790 948 -2788
rect 954 -2784 955 -2782
rect 954 -2790 955 -2788
rect 961 -2784 962 -2782
rect 961 -2790 962 -2788
rect 968 -2784 969 -2782
rect 968 -2790 969 -2788
rect 975 -2784 976 -2782
rect 975 -2790 976 -2788
rect 982 -2784 983 -2782
rect 982 -2790 983 -2788
rect 989 -2784 990 -2782
rect 989 -2790 990 -2788
rect 996 -2784 997 -2782
rect 996 -2790 997 -2788
rect 1003 -2790 1004 -2788
rect 1006 -2790 1007 -2788
rect 1010 -2784 1011 -2782
rect 1010 -2790 1011 -2788
rect 1017 -2784 1018 -2782
rect 1017 -2790 1018 -2788
rect 1024 -2784 1025 -2782
rect 1024 -2790 1025 -2788
rect 1031 -2784 1032 -2782
rect 1031 -2790 1032 -2788
rect 1038 -2784 1039 -2782
rect 1038 -2790 1039 -2788
rect 1045 -2784 1046 -2782
rect 1045 -2790 1046 -2788
rect 1052 -2784 1053 -2782
rect 1052 -2790 1053 -2788
rect 1059 -2784 1060 -2782
rect 1059 -2790 1060 -2788
rect 1066 -2784 1067 -2782
rect 1066 -2790 1067 -2788
rect 1073 -2784 1074 -2782
rect 1073 -2790 1074 -2788
rect 1080 -2784 1081 -2782
rect 1080 -2790 1081 -2788
rect 1087 -2784 1088 -2782
rect 1087 -2790 1088 -2788
rect 1094 -2784 1095 -2782
rect 1094 -2790 1095 -2788
rect 1101 -2784 1102 -2782
rect 1101 -2790 1102 -2788
rect 1108 -2784 1109 -2782
rect 1108 -2790 1109 -2788
rect 1115 -2784 1116 -2782
rect 1115 -2790 1116 -2788
rect 1122 -2784 1123 -2782
rect 1122 -2790 1123 -2788
rect 1129 -2784 1130 -2782
rect 1129 -2790 1130 -2788
rect 1136 -2784 1137 -2782
rect 1136 -2790 1137 -2788
rect 1143 -2784 1144 -2782
rect 1143 -2790 1144 -2788
rect 1150 -2784 1151 -2782
rect 1150 -2790 1151 -2788
rect 1157 -2784 1158 -2782
rect 1160 -2784 1161 -2782
rect 1157 -2790 1158 -2788
rect 1160 -2790 1161 -2788
rect 1164 -2784 1165 -2782
rect 1164 -2790 1165 -2788
rect 1171 -2784 1172 -2782
rect 1171 -2790 1172 -2788
rect 1178 -2784 1179 -2782
rect 1178 -2790 1179 -2788
rect 1185 -2784 1186 -2782
rect 1188 -2784 1189 -2782
rect 1185 -2790 1186 -2788
rect 1192 -2784 1193 -2782
rect 1192 -2790 1193 -2788
rect 1199 -2784 1200 -2782
rect 1199 -2790 1200 -2788
rect 1206 -2784 1207 -2782
rect 1206 -2790 1207 -2788
rect 1213 -2784 1214 -2782
rect 1213 -2790 1214 -2788
rect 1220 -2784 1221 -2782
rect 1220 -2790 1221 -2788
rect 1227 -2784 1228 -2782
rect 1227 -2790 1228 -2788
rect 1234 -2784 1235 -2782
rect 1234 -2790 1235 -2788
rect 1241 -2784 1242 -2782
rect 1241 -2790 1242 -2788
rect 1248 -2784 1249 -2782
rect 1248 -2790 1249 -2788
rect 1255 -2784 1256 -2782
rect 1255 -2790 1256 -2788
rect 1262 -2784 1263 -2782
rect 1262 -2790 1263 -2788
rect 1269 -2784 1270 -2782
rect 1269 -2790 1270 -2788
rect 1276 -2784 1277 -2782
rect 1276 -2790 1277 -2788
rect 1283 -2784 1284 -2782
rect 1283 -2790 1284 -2788
rect 1290 -2784 1291 -2782
rect 1290 -2790 1291 -2788
rect 1300 -2784 1301 -2782
rect 1297 -2790 1298 -2788
rect 1300 -2790 1301 -2788
rect 1304 -2784 1305 -2782
rect 1304 -2790 1305 -2788
rect 1311 -2784 1312 -2782
rect 1311 -2790 1312 -2788
rect 1318 -2784 1319 -2782
rect 1318 -2790 1319 -2788
rect 1325 -2784 1326 -2782
rect 1325 -2790 1326 -2788
rect 1332 -2784 1333 -2782
rect 1332 -2790 1333 -2788
rect 1339 -2784 1340 -2782
rect 1339 -2790 1340 -2788
rect 1346 -2784 1347 -2782
rect 1346 -2790 1347 -2788
rect 1353 -2784 1354 -2782
rect 1353 -2790 1354 -2788
rect 1360 -2784 1361 -2782
rect 1360 -2790 1361 -2788
rect 1367 -2784 1368 -2782
rect 1367 -2790 1368 -2788
rect 1374 -2784 1375 -2782
rect 1374 -2790 1375 -2788
rect 1381 -2784 1382 -2782
rect 1381 -2790 1382 -2788
rect 1388 -2784 1389 -2782
rect 1388 -2790 1389 -2788
rect 1395 -2784 1396 -2782
rect 1395 -2790 1396 -2788
rect 1402 -2784 1403 -2782
rect 1402 -2790 1403 -2788
rect 1409 -2784 1410 -2782
rect 1409 -2790 1410 -2788
rect 1416 -2784 1417 -2782
rect 1416 -2790 1417 -2788
rect 1423 -2784 1424 -2782
rect 1423 -2790 1424 -2788
rect 1430 -2784 1431 -2782
rect 1430 -2790 1431 -2788
rect 1437 -2784 1438 -2782
rect 1437 -2790 1438 -2788
rect 1444 -2784 1445 -2782
rect 1444 -2790 1445 -2788
rect 1451 -2784 1452 -2782
rect 1451 -2790 1452 -2788
rect 1458 -2784 1459 -2782
rect 1458 -2790 1459 -2788
rect 1465 -2784 1466 -2782
rect 1465 -2790 1466 -2788
rect 1472 -2784 1473 -2782
rect 1472 -2790 1473 -2788
rect 1479 -2784 1480 -2782
rect 1479 -2790 1480 -2788
rect 1486 -2784 1487 -2782
rect 1486 -2790 1487 -2788
rect 1493 -2784 1494 -2782
rect 1493 -2790 1494 -2788
rect 1500 -2784 1501 -2782
rect 1500 -2790 1501 -2788
rect 1507 -2784 1508 -2782
rect 1507 -2790 1508 -2788
rect 1514 -2784 1515 -2782
rect 1514 -2790 1515 -2788
rect 1521 -2784 1522 -2782
rect 1524 -2784 1525 -2782
rect 1521 -2790 1522 -2788
rect 72 -2909 73 -2907
rect 72 -2915 73 -2913
rect 79 -2909 80 -2907
rect 79 -2915 80 -2913
rect 86 -2909 87 -2907
rect 86 -2915 87 -2913
rect 93 -2909 94 -2907
rect 93 -2915 94 -2913
rect 103 -2909 104 -2907
rect 103 -2915 104 -2913
rect 107 -2909 108 -2907
rect 107 -2915 108 -2913
rect 114 -2909 115 -2907
rect 114 -2915 115 -2913
rect 121 -2909 122 -2907
rect 124 -2909 125 -2907
rect 121 -2915 122 -2913
rect 124 -2915 125 -2913
rect 128 -2909 129 -2907
rect 128 -2915 129 -2913
rect 135 -2909 136 -2907
rect 135 -2915 136 -2913
rect 142 -2909 143 -2907
rect 145 -2909 146 -2907
rect 142 -2915 143 -2913
rect 145 -2915 146 -2913
rect 149 -2909 150 -2907
rect 149 -2915 150 -2913
rect 156 -2909 157 -2907
rect 156 -2915 157 -2913
rect 163 -2909 164 -2907
rect 163 -2915 164 -2913
rect 170 -2909 171 -2907
rect 170 -2915 171 -2913
rect 177 -2909 178 -2907
rect 177 -2915 178 -2913
rect 184 -2909 185 -2907
rect 184 -2915 185 -2913
rect 191 -2909 192 -2907
rect 191 -2915 192 -2913
rect 198 -2909 199 -2907
rect 198 -2915 199 -2913
rect 205 -2909 206 -2907
rect 208 -2909 209 -2907
rect 205 -2915 206 -2913
rect 208 -2915 209 -2913
rect 212 -2909 213 -2907
rect 212 -2915 213 -2913
rect 219 -2909 220 -2907
rect 219 -2915 220 -2913
rect 226 -2909 227 -2907
rect 229 -2909 230 -2907
rect 229 -2915 230 -2913
rect 233 -2909 234 -2907
rect 233 -2915 234 -2913
rect 240 -2909 241 -2907
rect 240 -2915 241 -2913
rect 247 -2909 248 -2907
rect 250 -2909 251 -2907
rect 247 -2915 248 -2913
rect 250 -2915 251 -2913
rect 254 -2909 255 -2907
rect 254 -2915 255 -2913
rect 261 -2909 262 -2907
rect 261 -2915 262 -2913
rect 268 -2909 269 -2907
rect 268 -2915 269 -2913
rect 275 -2909 276 -2907
rect 278 -2909 279 -2907
rect 275 -2915 276 -2913
rect 278 -2915 279 -2913
rect 282 -2909 283 -2907
rect 285 -2909 286 -2907
rect 282 -2915 283 -2913
rect 285 -2915 286 -2913
rect 292 -2909 293 -2907
rect 289 -2915 290 -2913
rect 292 -2915 293 -2913
rect 296 -2909 297 -2907
rect 296 -2915 297 -2913
rect 303 -2909 304 -2907
rect 303 -2915 304 -2913
rect 310 -2909 311 -2907
rect 310 -2915 311 -2913
rect 317 -2909 318 -2907
rect 317 -2915 318 -2913
rect 324 -2909 325 -2907
rect 324 -2915 325 -2913
rect 331 -2909 332 -2907
rect 331 -2915 332 -2913
rect 338 -2909 339 -2907
rect 338 -2915 339 -2913
rect 345 -2909 346 -2907
rect 345 -2915 346 -2913
rect 352 -2909 353 -2907
rect 352 -2915 353 -2913
rect 359 -2909 360 -2907
rect 359 -2915 360 -2913
rect 366 -2909 367 -2907
rect 366 -2915 367 -2913
rect 373 -2909 374 -2907
rect 373 -2915 374 -2913
rect 380 -2909 381 -2907
rect 380 -2915 381 -2913
rect 387 -2909 388 -2907
rect 387 -2915 388 -2913
rect 394 -2909 395 -2907
rect 394 -2915 395 -2913
rect 401 -2909 402 -2907
rect 401 -2915 402 -2913
rect 408 -2909 409 -2907
rect 408 -2915 409 -2913
rect 415 -2909 416 -2907
rect 415 -2915 416 -2913
rect 422 -2909 423 -2907
rect 422 -2915 423 -2913
rect 429 -2909 430 -2907
rect 429 -2915 430 -2913
rect 436 -2909 437 -2907
rect 436 -2915 437 -2913
rect 443 -2909 444 -2907
rect 443 -2915 444 -2913
rect 450 -2909 451 -2907
rect 450 -2915 451 -2913
rect 457 -2909 458 -2907
rect 457 -2915 458 -2913
rect 464 -2909 465 -2907
rect 464 -2915 465 -2913
rect 471 -2909 472 -2907
rect 471 -2915 472 -2913
rect 478 -2909 479 -2907
rect 478 -2915 479 -2913
rect 485 -2909 486 -2907
rect 485 -2915 486 -2913
rect 495 -2909 496 -2907
rect 492 -2915 493 -2913
rect 495 -2915 496 -2913
rect 499 -2909 500 -2907
rect 499 -2915 500 -2913
rect 506 -2909 507 -2907
rect 506 -2915 507 -2913
rect 513 -2909 514 -2907
rect 513 -2915 514 -2913
rect 520 -2909 521 -2907
rect 520 -2915 521 -2913
rect 527 -2909 528 -2907
rect 527 -2915 528 -2913
rect 534 -2909 535 -2907
rect 534 -2915 535 -2913
rect 541 -2909 542 -2907
rect 541 -2915 542 -2913
rect 548 -2909 549 -2907
rect 548 -2915 549 -2913
rect 555 -2909 556 -2907
rect 558 -2909 559 -2907
rect 562 -2909 563 -2907
rect 562 -2915 563 -2913
rect 569 -2909 570 -2907
rect 569 -2915 570 -2913
rect 576 -2909 577 -2907
rect 576 -2915 577 -2913
rect 583 -2915 584 -2913
rect 586 -2915 587 -2913
rect 590 -2909 591 -2907
rect 590 -2915 591 -2913
rect 597 -2909 598 -2907
rect 597 -2915 598 -2913
rect 604 -2909 605 -2907
rect 604 -2915 605 -2913
rect 611 -2909 612 -2907
rect 611 -2915 612 -2913
rect 618 -2909 619 -2907
rect 618 -2915 619 -2913
rect 625 -2909 626 -2907
rect 625 -2915 626 -2913
rect 632 -2909 633 -2907
rect 632 -2915 633 -2913
rect 639 -2909 640 -2907
rect 642 -2909 643 -2907
rect 639 -2915 640 -2913
rect 642 -2915 643 -2913
rect 646 -2909 647 -2907
rect 646 -2915 647 -2913
rect 653 -2909 654 -2907
rect 653 -2915 654 -2913
rect 660 -2909 661 -2907
rect 663 -2909 664 -2907
rect 660 -2915 661 -2913
rect 663 -2915 664 -2913
rect 667 -2909 668 -2907
rect 667 -2915 668 -2913
rect 674 -2909 675 -2907
rect 674 -2915 675 -2913
rect 681 -2909 682 -2907
rect 681 -2915 682 -2913
rect 688 -2909 689 -2907
rect 688 -2915 689 -2913
rect 695 -2909 696 -2907
rect 695 -2915 696 -2913
rect 702 -2909 703 -2907
rect 705 -2909 706 -2907
rect 702 -2915 703 -2913
rect 705 -2915 706 -2913
rect 709 -2909 710 -2907
rect 709 -2915 710 -2913
rect 716 -2909 717 -2907
rect 716 -2915 717 -2913
rect 723 -2909 724 -2907
rect 723 -2915 724 -2913
rect 730 -2909 731 -2907
rect 730 -2915 731 -2913
rect 737 -2909 738 -2907
rect 737 -2915 738 -2913
rect 744 -2909 745 -2907
rect 744 -2915 745 -2913
rect 747 -2915 748 -2913
rect 751 -2909 752 -2907
rect 751 -2915 752 -2913
rect 758 -2909 759 -2907
rect 761 -2909 762 -2907
rect 758 -2915 759 -2913
rect 761 -2915 762 -2913
rect 765 -2909 766 -2907
rect 765 -2915 766 -2913
rect 772 -2909 773 -2907
rect 772 -2915 773 -2913
rect 779 -2909 780 -2907
rect 779 -2915 780 -2913
rect 786 -2909 787 -2907
rect 786 -2915 787 -2913
rect 793 -2909 794 -2907
rect 793 -2915 794 -2913
rect 800 -2909 801 -2907
rect 800 -2915 801 -2913
rect 807 -2909 808 -2907
rect 807 -2915 808 -2913
rect 814 -2909 815 -2907
rect 814 -2915 815 -2913
rect 821 -2909 822 -2907
rect 824 -2909 825 -2907
rect 821 -2915 822 -2913
rect 824 -2915 825 -2913
rect 828 -2909 829 -2907
rect 828 -2915 829 -2913
rect 835 -2909 836 -2907
rect 838 -2909 839 -2907
rect 835 -2915 836 -2913
rect 838 -2915 839 -2913
rect 842 -2909 843 -2907
rect 845 -2909 846 -2907
rect 842 -2915 843 -2913
rect 849 -2909 850 -2907
rect 849 -2915 850 -2913
rect 856 -2909 857 -2907
rect 856 -2915 857 -2913
rect 866 -2909 867 -2907
rect 863 -2915 864 -2913
rect 866 -2915 867 -2913
rect 870 -2909 871 -2907
rect 870 -2915 871 -2913
rect 877 -2909 878 -2907
rect 877 -2915 878 -2913
rect 884 -2909 885 -2907
rect 884 -2915 885 -2913
rect 891 -2909 892 -2907
rect 891 -2915 892 -2913
rect 898 -2909 899 -2907
rect 898 -2915 899 -2913
rect 905 -2909 906 -2907
rect 912 -2909 913 -2907
rect 915 -2909 916 -2907
rect 912 -2915 913 -2913
rect 915 -2915 916 -2913
rect 919 -2909 920 -2907
rect 922 -2909 923 -2907
rect 919 -2915 920 -2913
rect 922 -2915 923 -2913
rect 926 -2909 927 -2907
rect 926 -2915 927 -2913
rect 933 -2909 934 -2907
rect 933 -2915 934 -2913
rect 940 -2909 941 -2907
rect 940 -2915 941 -2913
rect 947 -2909 948 -2907
rect 947 -2915 948 -2913
rect 950 -2915 951 -2913
rect 954 -2909 955 -2907
rect 957 -2909 958 -2907
rect 954 -2915 955 -2913
rect 957 -2915 958 -2913
rect 961 -2909 962 -2907
rect 961 -2915 962 -2913
rect 968 -2909 969 -2907
rect 968 -2915 969 -2913
rect 975 -2909 976 -2907
rect 975 -2915 976 -2913
rect 982 -2909 983 -2907
rect 982 -2915 983 -2913
rect 989 -2909 990 -2907
rect 989 -2915 990 -2913
rect 996 -2909 997 -2907
rect 996 -2915 997 -2913
rect 1003 -2909 1004 -2907
rect 1003 -2915 1004 -2913
rect 1010 -2909 1011 -2907
rect 1010 -2915 1011 -2913
rect 1017 -2909 1018 -2907
rect 1020 -2909 1021 -2907
rect 1017 -2915 1018 -2913
rect 1020 -2915 1021 -2913
rect 1024 -2909 1025 -2907
rect 1024 -2915 1025 -2913
rect 1031 -2909 1032 -2907
rect 1031 -2915 1032 -2913
rect 1038 -2909 1039 -2907
rect 1038 -2915 1039 -2913
rect 1045 -2909 1046 -2907
rect 1045 -2915 1046 -2913
rect 1052 -2909 1053 -2907
rect 1052 -2915 1053 -2913
rect 1059 -2909 1060 -2907
rect 1059 -2915 1060 -2913
rect 1066 -2909 1067 -2907
rect 1066 -2915 1067 -2913
rect 1073 -2909 1074 -2907
rect 1073 -2915 1074 -2913
rect 1080 -2909 1081 -2907
rect 1080 -2915 1081 -2913
rect 1087 -2909 1088 -2907
rect 1087 -2915 1088 -2913
rect 1094 -2909 1095 -2907
rect 1097 -2909 1098 -2907
rect 1094 -2915 1095 -2913
rect 1097 -2915 1098 -2913
rect 1101 -2909 1102 -2907
rect 1101 -2915 1102 -2913
rect 1108 -2909 1109 -2907
rect 1108 -2915 1109 -2913
rect 1115 -2909 1116 -2907
rect 1115 -2915 1116 -2913
rect 1122 -2909 1123 -2907
rect 1122 -2915 1123 -2913
rect 1129 -2909 1130 -2907
rect 1129 -2915 1130 -2913
rect 1136 -2909 1137 -2907
rect 1136 -2915 1137 -2913
rect 1143 -2909 1144 -2907
rect 1143 -2915 1144 -2913
rect 1150 -2909 1151 -2907
rect 1150 -2915 1151 -2913
rect 1157 -2909 1158 -2907
rect 1157 -2915 1158 -2913
rect 1164 -2909 1165 -2907
rect 1164 -2915 1165 -2913
rect 1171 -2909 1172 -2907
rect 1171 -2915 1172 -2913
rect 1178 -2909 1179 -2907
rect 1178 -2915 1179 -2913
rect 1185 -2909 1186 -2907
rect 1185 -2915 1186 -2913
rect 1192 -2909 1193 -2907
rect 1192 -2915 1193 -2913
rect 1199 -2909 1200 -2907
rect 1199 -2915 1200 -2913
rect 1206 -2909 1207 -2907
rect 1206 -2915 1207 -2913
rect 1213 -2909 1214 -2907
rect 1213 -2915 1214 -2913
rect 1220 -2909 1221 -2907
rect 1220 -2915 1221 -2913
rect 1227 -2909 1228 -2907
rect 1227 -2915 1228 -2913
rect 1230 -2915 1231 -2913
rect 1234 -2909 1235 -2907
rect 1234 -2915 1235 -2913
rect 1241 -2909 1242 -2907
rect 1241 -2915 1242 -2913
rect 1248 -2909 1249 -2907
rect 1248 -2915 1249 -2913
rect 1255 -2909 1256 -2907
rect 1255 -2915 1256 -2913
rect 1262 -2909 1263 -2907
rect 1262 -2915 1263 -2913
rect 1269 -2909 1270 -2907
rect 1269 -2915 1270 -2913
rect 1276 -2909 1277 -2907
rect 1276 -2915 1277 -2913
rect 1283 -2909 1284 -2907
rect 1283 -2915 1284 -2913
rect 1290 -2909 1291 -2907
rect 1290 -2915 1291 -2913
rect 1297 -2909 1298 -2907
rect 1297 -2915 1298 -2913
rect 1304 -2909 1305 -2907
rect 1304 -2915 1305 -2913
rect 1311 -2909 1312 -2907
rect 1311 -2915 1312 -2913
rect 1318 -2909 1319 -2907
rect 1318 -2915 1319 -2913
rect 1325 -2909 1326 -2907
rect 1325 -2915 1326 -2913
rect 1332 -2909 1333 -2907
rect 1332 -2915 1333 -2913
rect 1339 -2909 1340 -2907
rect 1339 -2915 1340 -2913
rect 1346 -2909 1347 -2907
rect 1346 -2915 1347 -2913
rect 1353 -2909 1354 -2907
rect 1353 -2915 1354 -2913
rect 1363 -2909 1364 -2907
rect 1360 -2915 1361 -2913
rect 1367 -2909 1368 -2907
rect 1367 -2915 1368 -2913
rect 1374 -2909 1375 -2907
rect 1374 -2915 1375 -2913
rect 1381 -2909 1382 -2907
rect 1381 -2915 1382 -2913
rect 1388 -2909 1389 -2907
rect 1388 -2915 1389 -2913
rect 1395 -2909 1396 -2907
rect 1395 -2915 1396 -2913
rect 1402 -2909 1403 -2907
rect 1402 -2915 1403 -2913
rect 1409 -2909 1410 -2907
rect 1409 -2915 1410 -2913
rect 1416 -2909 1417 -2907
rect 1416 -2915 1417 -2913
rect 1423 -2909 1424 -2907
rect 1423 -2915 1424 -2913
rect 1430 -2909 1431 -2907
rect 1430 -2915 1431 -2913
rect 86 -3028 87 -3026
rect 86 -3034 87 -3032
rect 93 -3028 94 -3026
rect 93 -3034 94 -3032
rect 100 -3028 101 -3026
rect 100 -3034 101 -3032
rect 107 -3028 108 -3026
rect 107 -3034 108 -3032
rect 114 -3028 115 -3026
rect 114 -3034 115 -3032
rect 121 -3028 122 -3026
rect 121 -3034 122 -3032
rect 128 -3028 129 -3026
rect 128 -3034 129 -3032
rect 135 -3028 136 -3026
rect 135 -3034 136 -3032
rect 142 -3028 143 -3026
rect 142 -3034 143 -3032
rect 149 -3028 150 -3026
rect 149 -3034 150 -3032
rect 152 -3034 153 -3032
rect 156 -3028 157 -3026
rect 156 -3034 157 -3032
rect 163 -3028 164 -3026
rect 166 -3028 167 -3026
rect 163 -3034 164 -3032
rect 166 -3034 167 -3032
rect 170 -3028 171 -3026
rect 170 -3034 171 -3032
rect 177 -3028 178 -3026
rect 177 -3034 178 -3032
rect 184 -3028 185 -3026
rect 184 -3034 185 -3032
rect 191 -3028 192 -3026
rect 191 -3034 192 -3032
rect 198 -3028 199 -3026
rect 198 -3034 199 -3032
rect 208 -3028 209 -3026
rect 208 -3034 209 -3032
rect 212 -3028 213 -3026
rect 212 -3034 213 -3032
rect 219 -3028 220 -3026
rect 222 -3028 223 -3026
rect 219 -3034 220 -3032
rect 226 -3028 227 -3026
rect 226 -3034 227 -3032
rect 233 -3028 234 -3026
rect 233 -3034 234 -3032
rect 240 -3028 241 -3026
rect 240 -3034 241 -3032
rect 247 -3028 248 -3026
rect 254 -3028 255 -3026
rect 254 -3034 255 -3032
rect 261 -3028 262 -3026
rect 264 -3028 265 -3026
rect 261 -3034 262 -3032
rect 268 -3028 269 -3026
rect 268 -3034 269 -3032
rect 275 -3028 276 -3026
rect 275 -3034 276 -3032
rect 282 -3028 283 -3026
rect 289 -3028 290 -3026
rect 289 -3034 290 -3032
rect 296 -3028 297 -3026
rect 296 -3034 297 -3032
rect 303 -3028 304 -3026
rect 303 -3034 304 -3032
rect 310 -3028 311 -3026
rect 310 -3034 311 -3032
rect 317 -3028 318 -3026
rect 317 -3034 318 -3032
rect 324 -3028 325 -3026
rect 324 -3034 325 -3032
rect 331 -3028 332 -3026
rect 331 -3034 332 -3032
rect 338 -3028 339 -3026
rect 338 -3034 339 -3032
rect 345 -3028 346 -3026
rect 345 -3034 346 -3032
rect 352 -3028 353 -3026
rect 352 -3034 353 -3032
rect 359 -3028 360 -3026
rect 359 -3034 360 -3032
rect 366 -3028 367 -3026
rect 366 -3034 367 -3032
rect 373 -3028 374 -3026
rect 373 -3034 374 -3032
rect 380 -3028 381 -3026
rect 380 -3034 381 -3032
rect 387 -3028 388 -3026
rect 387 -3034 388 -3032
rect 394 -3028 395 -3026
rect 394 -3034 395 -3032
rect 401 -3028 402 -3026
rect 401 -3034 402 -3032
rect 408 -3028 409 -3026
rect 411 -3028 412 -3026
rect 408 -3034 409 -3032
rect 411 -3034 412 -3032
rect 415 -3028 416 -3026
rect 415 -3034 416 -3032
rect 422 -3028 423 -3026
rect 422 -3034 423 -3032
rect 429 -3028 430 -3026
rect 429 -3034 430 -3032
rect 436 -3028 437 -3026
rect 436 -3034 437 -3032
rect 443 -3028 444 -3026
rect 443 -3034 444 -3032
rect 450 -3028 451 -3026
rect 450 -3034 451 -3032
rect 457 -3028 458 -3026
rect 457 -3034 458 -3032
rect 464 -3028 465 -3026
rect 464 -3034 465 -3032
rect 471 -3028 472 -3026
rect 471 -3034 472 -3032
rect 478 -3028 479 -3026
rect 478 -3034 479 -3032
rect 485 -3028 486 -3026
rect 485 -3034 486 -3032
rect 492 -3028 493 -3026
rect 492 -3034 493 -3032
rect 499 -3028 500 -3026
rect 499 -3034 500 -3032
rect 509 -3034 510 -3032
rect 513 -3028 514 -3026
rect 513 -3034 514 -3032
rect 520 -3028 521 -3026
rect 520 -3034 521 -3032
rect 527 -3028 528 -3026
rect 527 -3034 528 -3032
rect 534 -3028 535 -3026
rect 534 -3034 535 -3032
rect 541 -3028 542 -3026
rect 541 -3034 542 -3032
rect 548 -3028 549 -3026
rect 548 -3034 549 -3032
rect 555 -3028 556 -3026
rect 555 -3034 556 -3032
rect 562 -3028 563 -3026
rect 562 -3034 563 -3032
rect 569 -3028 570 -3026
rect 569 -3034 570 -3032
rect 576 -3028 577 -3026
rect 576 -3034 577 -3032
rect 583 -3028 584 -3026
rect 583 -3034 584 -3032
rect 590 -3028 591 -3026
rect 590 -3034 591 -3032
rect 597 -3028 598 -3026
rect 597 -3034 598 -3032
rect 604 -3028 605 -3026
rect 604 -3034 605 -3032
rect 611 -3028 612 -3026
rect 611 -3034 612 -3032
rect 618 -3028 619 -3026
rect 618 -3034 619 -3032
rect 625 -3028 626 -3026
rect 625 -3034 626 -3032
rect 632 -3028 633 -3026
rect 635 -3028 636 -3026
rect 635 -3034 636 -3032
rect 639 -3028 640 -3026
rect 639 -3034 640 -3032
rect 646 -3028 647 -3026
rect 649 -3028 650 -3026
rect 649 -3034 650 -3032
rect 653 -3028 654 -3026
rect 653 -3034 654 -3032
rect 660 -3028 661 -3026
rect 663 -3028 664 -3026
rect 660 -3034 661 -3032
rect 667 -3028 668 -3026
rect 667 -3034 668 -3032
rect 674 -3028 675 -3026
rect 674 -3034 675 -3032
rect 681 -3028 682 -3026
rect 681 -3034 682 -3032
rect 688 -3028 689 -3026
rect 691 -3028 692 -3026
rect 688 -3034 689 -3032
rect 691 -3034 692 -3032
rect 695 -3028 696 -3026
rect 698 -3028 699 -3026
rect 695 -3034 696 -3032
rect 698 -3034 699 -3032
rect 702 -3028 703 -3026
rect 702 -3034 703 -3032
rect 709 -3028 710 -3026
rect 709 -3034 710 -3032
rect 716 -3028 717 -3026
rect 716 -3034 717 -3032
rect 723 -3028 724 -3026
rect 723 -3034 724 -3032
rect 730 -3028 731 -3026
rect 730 -3034 731 -3032
rect 733 -3034 734 -3032
rect 737 -3028 738 -3026
rect 737 -3034 738 -3032
rect 744 -3028 745 -3026
rect 744 -3034 745 -3032
rect 751 -3028 752 -3026
rect 754 -3028 755 -3026
rect 754 -3034 755 -3032
rect 758 -3028 759 -3026
rect 758 -3034 759 -3032
rect 768 -3028 769 -3026
rect 765 -3034 766 -3032
rect 772 -3028 773 -3026
rect 772 -3034 773 -3032
rect 779 -3028 780 -3026
rect 779 -3034 780 -3032
rect 786 -3028 787 -3026
rect 789 -3028 790 -3026
rect 786 -3034 787 -3032
rect 789 -3034 790 -3032
rect 793 -3028 794 -3026
rect 793 -3034 794 -3032
rect 800 -3028 801 -3026
rect 800 -3034 801 -3032
rect 807 -3028 808 -3026
rect 807 -3034 808 -3032
rect 814 -3028 815 -3026
rect 814 -3034 815 -3032
rect 821 -3028 822 -3026
rect 821 -3034 822 -3032
rect 828 -3028 829 -3026
rect 828 -3034 829 -3032
rect 835 -3028 836 -3026
rect 838 -3028 839 -3026
rect 835 -3034 836 -3032
rect 838 -3034 839 -3032
rect 842 -3028 843 -3026
rect 842 -3034 843 -3032
rect 849 -3028 850 -3026
rect 849 -3034 850 -3032
rect 856 -3028 857 -3026
rect 856 -3034 857 -3032
rect 863 -3028 864 -3026
rect 866 -3028 867 -3026
rect 863 -3034 864 -3032
rect 866 -3034 867 -3032
rect 870 -3028 871 -3026
rect 873 -3028 874 -3026
rect 873 -3034 874 -3032
rect 877 -3028 878 -3026
rect 877 -3034 878 -3032
rect 884 -3028 885 -3026
rect 884 -3034 885 -3032
rect 887 -3034 888 -3032
rect 891 -3028 892 -3026
rect 891 -3034 892 -3032
rect 898 -3028 899 -3026
rect 898 -3034 899 -3032
rect 905 -3034 906 -3032
rect 912 -3028 913 -3026
rect 915 -3028 916 -3026
rect 912 -3034 913 -3032
rect 919 -3028 920 -3026
rect 922 -3028 923 -3026
rect 919 -3034 920 -3032
rect 922 -3034 923 -3032
rect 926 -3028 927 -3026
rect 926 -3034 927 -3032
rect 933 -3028 934 -3026
rect 933 -3034 934 -3032
rect 940 -3028 941 -3026
rect 940 -3034 941 -3032
rect 947 -3028 948 -3026
rect 947 -3034 948 -3032
rect 954 -3028 955 -3026
rect 954 -3034 955 -3032
rect 961 -3028 962 -3026
rect 961 -3034 962 -3032
rect 968 -3028 969 -3026
rect 968 -3034 969 -3032
rect 975 -3028 976 -3026
rect 975 -3034 976 -3032
rect 982 -3028 983 -3026
rect 982 -3034 983 -3032
rect 989 -3028 990 -3026
rect 989 -3034 990 -3032
rect 996 -3028 997 -3026
rect 996 -3034 997 -3032
rect 1003 -3028 1004 -3026
rect 1003 -3034 1004 -3032
rect 1010 -3028 1011 -3026
rect 1010 -3034 1011 -3032
rect 1017 -3028 1018 -3026
rect 1020 -3034 1021 -3032
rect 1024 -3028 1025 -3026
rect 1024 -3034 1025 -3032
rect 1031 -3028 1032 -3026
rect 1031 -3034 1032 -3032
rect 1038 -3028 1039 -3026
rect 1038 -3034 1039 -3032
rect 1045 -3028 1046 -3026
rect 1045 -3034 1046 -3032
rect 1052 -3028 1053 -3026
rect 1052 -3034 1053 -3032
rect 1059 -3028 1060 -3026
rect 1059 -3034 1060 -3032
rect 1066 -3028 1067 -3026
rect 1066 -3034 1067 -3032
rect 1073 -3028 1074 -3026
rect 1076 -3028 1077 -3026
rect 1073 -3034 1074 -3032
rect 1080 -3028 1081 -3026
rect 1080 -3034 1081 -3032
rect 1087 -3028 1088 -3026
rect 1087 -3034 1088 -3032
rect 1094 -3028 1095 -3026
rect 1094 -3034 1095 -3032
rect 1101 -3028 1102 -3026
rect 1101 -3034 1102 -3032
rect 1108 -3028 1109 -3026
rect 1108 -3034 1109 -3032
rect 1115 -3028 1116 -3026
rect 1115 -3034 1116 -3032
rect 1122 -3028 1123 -3026
rect 1122 -3034 1123 -3032
rect 1129 -3028 1130 -3026
rect 1129 -3034 1130 -3032
rect 1136 -3028 1137 -3026
rect 1136 -3034 1137 -3032
rect 1143 -3028 1144 -3026
rect 1143 -3034 1144 -3032
rect 1150 -3034 1151 -3032
rect 1153 -3034 1154 -3032
rect 1157 -3028 1158 -3026
rect 1157 -3034 1158 -3032
rect 1164 -3028 1165 -3026
rect 1164 -3034 1165 -3032
rect 1171 -3028 1172 -3026
rect 1171 -3034 1172 -3032
rect 1178 -3028 1179 -3026
rect 1178 -3034 1179 -3032
rect 1185 -3028 1186 -3026
rect 1185 -3034 1186 -3032
rect 1192 -3028 1193 -3026
rect 1192 -3034 1193 -3032
rect 1199 -3028 1200 -3026
rect 1199 -3034 1200 -3032
rect 1206 -3028 1207 -3026
rect 1206 -3034 1207 -3032
rect 1213 -3028 1214 -3026
rect 1213 -3034 1214 -3032
rect 1220 -3028 1221 -3026
rect 1220 -3034 1221 -3032
rect 1227 -3028 1228 -3026
rect 1230 -3028 1231 -3026
rect 1227 -3034 1228 -3032
rect 1234 -3028 1235 -3026
rect 1234 -3034 1235 -3032
rect 1241 -3028 1242 -3026
rect 1241 -3034 1242 -3032
rect 1248 -3028 1249 -3026
rect 1248 -3034 1249 -3032
rect 1255 -3028 1256 -3026
rect 1255 -3034 1256 -3032
rect 1262 -3028 1263 -3026
rect 1262 -3034 1263 -3032
rect 1269 -3028 1270 -3026
rect 1269 -3034 1270 -3032
rect 1276 -3028 1277 -3026
rect 1276 -3034 1277 -3032
rect 1283 -3028 1284 -3026
rect 1283 -3034 1284 -3032
rect 1290 -3028 1291 -3026
rect 1290 -3034 1291 -3032
rect 1297 -3028 1298 -3026
rect 1297 -3034 1298 -3032
rect 1304 -3028 1305 -3026
rect 1304 -3034 1305 -3032
rect 1311 -3028 1312 -3026
rect 1311 -3034 1312 -3032
rect 1318 -3028 1319 -3026
rect 1318 -3034 1319 -3032
rect 1325 -3028 1326 -3026
rect 1325 -3034 1326 -3032
rect 1332 -3028 1333 -3026
rect 1332 -3034 1333 -3032
rect 1339 -3028 1340 -3026
rect 1339 -3034 1340 -3032
rect 1346 -3028 1347 -3026
rect 1346 -3034 1347 -3032
rect 1353 -3028 1354 -3026
rect 1353 -3034 1354 -3032
rect 1360 -3028 1361 -3026
rect 1360 -3034 1361 -3032
rect 1367 -3028 1368 -3026
rect 1367 -3034 1368 -3032
rect 1374 -3028 1375 -3026
rect 1374 -3034 1375 -3032
rect 1381 -3028 1382 -3026
rect 1381 -3034 1382 -3032
rect 1388 -3028 1389 -3026
rect 1388 -3034 1389 -3032
rect 1395 -3028 1396 -3026
rect 1395 -3034 1396 -3032
rect 1402 -3028 1403 -3026
rect 1402 -3034 1403 -3032
rect 1409 -3028 1410 -3026
rect 1409 -3034 1410 -3032
rect 100 -3139 101 -3137
rect 100 -3145 101 -3143
rect 107 -3139 108 -3137
rect 107 -3145 108 -3143
rect 114 -3139 115 -3137
rect 114 -3145 115 -3143
rect 121 -3139 122 -3137
rect 121 -3145 122 -3143
rect 128 -3139 129 -3137
rect 128 -3145 129 -3143
rect 135 -3139 136 -3137
rect 135 -3145 136 -3143
rect 142 -3139 143 -3137
rect 142 -3145 143 -3143
rect 149 -3139 150 -3137
rect 149 -3145 150 -3143
rect 156 -3139 157 -3137
rect 156 -3145 157 -3143
rect 159 -3145 160 -3143
rect 163 -3139 164 -3137
rect 163 -3145 164 -3143
rect 170 -3139 171 -3137
rect 170 -3145 171 -3143
rect 177 -3139 178 -3137
rect 177 -3145 178 -3143
rect 184 -3139 185 -3137
rect 184 -3145 185 -3143
rect 191 -3139 192 -3137
rect 191 -3145 192 -3143
rect 198 -3139 199 -3137
rect 198 -3145 199 -3143
rect 205 -3139 206 -3137
rect 205 -3145 206 -3143
rect 212 -3139 213 -3137
rect 212 -3145 213 -3143
rect 222 -3139 223 -3137
rect 222 -3145 223 -3143
rect 226 -3139 227 -3137
rect 229 -3139 230 -3137
rect 229 -3145 230 -3143
rect 233 -3139 234 -3137
rect 233 -3145 234 -3143
rect 240 -3139 241 -3137
rect 240 -3145 241 -3143
rect 247 -3139 248 -3137
rect 247 -3145 248 -3143
rect 250 -3145 251 -3143
rect 254 -3139 255 -3137
rect 257 -3139 258 -3137
rect 261 -3139 262 -3137
rect 261 -3145 262 -3143
rect 268 -3139 269 -3137
rect 268 -3145 269 -3143
rect 275 -3139 276 -3137
rect 275 -3145 276 -3143
rect 282 -3145 283 -3143
rect 289 -3139 290 -3137
rect 289 -3145 290 -3143
rect 296 -3139 297 -3137
rect 296 -3145 297 -3143
rect 303 -3139 304 -3137
rect 303 -3145 304 -3143
rect 310 -3139 311 -3137
rect 310 -3145 311 -3143
rect 317 -3139 318 -3137
rect 317 -3145 318 -3143
rect 324 -3139 325 -3137
rect 327 -3139 328 -3137
rect 324 -3145 325 -3143
rect 327 -3145 328 -3143
rect 331 -3139 332 -3137
rect 331 -3145 332 -3143
rect 338 -3139 339 -3137
rect 338 -3145 339 -3143
rect 345 -3139 346 -3137
rect 345 -3145 346 -3143
rect 352 -3139 353 -3137
rect 352 -3145 353 -3143
rect 359 -3139 360 -3137
rect 359 -3145 360 -3143
rect 366 -3139 367 -3137
rect 366 -3145 367 -3143
rect 373 -3139 374 -3137
rect 373 -3145 374 -3143
rect 380 -3139 381 -3137
rect 380 -3145 381 -3143
rect 387 -3145 388 -3143
rect 390 -3145 391 -3143
rect 394 -3139 395 -3137
rect 394 -3145 395 -3143
rect 401 -3139 402 -3137
rect 401 -3145 402 -3143
rect 411 -3139 412 -3137
rect 408 -3145 409 -3143
rect 411 -3145 412 -3143
rect 415 -3139 416 -3137
rect 415 -3145 416 -3143
rect 422 -3139 423 -3137
rect 422 -3145 423 -3143
rect 429 -3139 430 -3137
rect 429 -3145 430 -3143
rect 436 -3139 437 -3137
rect 436 -3145 437 -3143
rect 443 -3139 444 -3137
rect 443 -3145 444 -3143
rect 450 -3139 451 -3137
rect 450 -3145 451 -3143
rect 457 -3139 458 -3137
rect 457 -3145 458 -3143
rect 464 -3139 465 -3137
rect 464 -3145 465 -3143
rect 471 -3139 472 -3137
rect 471 -3145 472 -3143
rect 478 -3139 479 -3137
rect 478 -3145 479 -3143
rect 485 -3139 486 -3137
rect 485 -3145 486 -3143
rect 492 -3139 493 -3137
rect 492 -3145 493 -3143
rect 499 -3139 500 -3137
rect 499 -3145 500 -3143
rect 506 -3139 507 -3137
rect 506 -3145 507 -3143
rect 513 -3139 514 -3137
rect 516 -3139 517 -3137
rect 513 -3145 514 -3143
rect 516 -3145 517 -3143
rect 520 -3139 521 -3137
rect 520 -3145 521 -3143
rect 527 -3139 528 -3137
rect 527 -3145 528 -3143
rect 534 -3139 535 -3137
rect 534 -3145 535 -3143
rect 541 -3139 542 -3137
rect 541 -3145 542 -3143
rect 548 -3139 549 -3137
rect 548 -3145 549 -3143
rect 555 -3139 556 -3137
rect 555 -3145 556 -3143
rect 562 -3139 563 -3137
rect 562 -3145 563 -3143
rect 569 -3139 570 -3137
rect 569 -3145 570 -3143
rect 576 -3139 577 -3137
rect 576 -3145 577 -3143
rect 583 -3139 584 -3137
rect 583 -3145 584 -3143
rect 590 -3139 591 -3137
rect 590 -3145 591 -3143
rect 593 -3145 594 -3143
rect 597 -3139 598 -3137
rect 597 -3145 598 -3143
rect 607 -3139 608 -3137
rect 604 -3145 605 -3143
rect 607 -3145 608 -3143
rect 611 -3139 612 -3137
rect 611 -3145 612 -3143
rect 618 -3139 619 -3137
rect 618 -3145 619 -3143
rect 625 -3139 626 -3137
rect 625 -3145 626 -3143
rect 632 -3139 633 -3137
rect 632 -3145 633 -3143
rect 639 -3139 640 -3137
rect 639 -3145 640 -3143
rect 646 -3139 647 -3137
rect 649 -3139 650 -3137
rect 646 -3145 647 -3143
rect 653 -3139 654 -3137
rect 653 -3145 654 -3143
rect 660 -3139 661 -3137
rect 660 -3145 661 -3143
rect 667 -3139 668 -3137
rect 667 -3145 668 -3143
rect 674 -3139 675 -3137
rect 674 -3145 675 -3143
rect 681 -3139 682 -3137
rect 681 -3145 682 -3143
rect 688 -3139 689 -3137
rect 688 -3145 689 -3143
rect 695 -3139 696 -3137
rect 698 -3139 699 -3137
rect 695 -3145 696 -3143
rect 698 -3145 699 -3143
rect 702 -3139 703 -3137
rect 702 -3145 703 -3143
rect 709 -3139 710 -3137
rect 709 -3145 710 -3143
rect 716 -3139 717 -3137
rect 716 -3145 717 -3143
rect 723 -3139 724 -3137
rect 723 -3145 724 -3143
rect 730 -3139 731 -3137
rect 733 -3139 734 -3137
rect 730 -3145 731 -3143
rect 737 -3139 738 -3137
rect 740 -3139 741 -3137
rect 737 -3145 738 -3143
rect 740 -3145 741 -3143
rect 744 -3139 745 -3137
rect 747 -3139 748 -3137
rect 744 -3145 745 -3143
rect 747 -3145 748 -3143
rect 751 -3139 752 -3137
rect 751 -3145 752 -3143
rect 761 -3139 762 -3137
rect 758 -3145 759 -3143
rect 761 -3145 762 -3143
rect 765 -3139 766 -3137
rect 765 -3145 766 -3143
rect 772 -3139 773 -3137
rect 772 -3145 773 -3143
rect 779 -3139 780 -3137
rect 779 -3145 780 -3143
rect 786 -3139 787 -3137
rect 786 -3145 787 -3143
rect 793 -3139 794 -3137
rect 796 -3139 797 -3137
rect 793 -3145 794 -3143
rect 796 -3145 797 -3143
rect 800 -3139 801 -3137
rect 800 -3145 801 -3143
rect 807 -3139 808 -3137
rect 810 -3139 811 -3137
rect 807 -3145 808 -3143
rect 810 -3145 811 -3143
rect 814 -3139 815 -3137
rect 814 -3145 815 -3143
rect 821 -3139 822 -3137
rect 821 -3145 822 -3143
rect 828 -3139 829 -3137
rect 828 -3145 829 -3143
rect 835 -3139 836 -3137
rect 835 -3145 836 -3143
rect 842 -3139 843 -3137
rect 842 -3145 843 -3143
rect 849 -3139 850 -3137
rect 849 -3145 850 -3143
rect 856 -3139 857 -3137
rect 856 -3145 857 -3143
rect 863 -3139 864 -3137
rect 863 -3145 864 -3143
rect 870 -3139 871 -3137
rect 870 -3145 871 -3143
rect 877 -3139 878 -3137
rect 877 -3145 878 -3143
rect 884 -3139 885 -3137
rect 884 -3145 885 -3143
rect 891 -3139 892 -3137
rect 891 -3145 892 -3143
rect 898 -3139 899 -3137
rect 901 -3139 902 -3137
rect 898 -3145 899 -3143
rect 901 -3145 902 -3143
rect 905 -3139 906 -3137
rect 905 -3145 906 -3143
rect 912 -3139 913 -3137
rect 915 -3139 916 -3137
rect 915 -3145 916 -3143
rect 919 -3139 920 -3137
rect 919 -3145 920 -3143
rect 926 -3139 927 -3137
rect 926 -3145 927 -3143
rect 933 -3139 934 -3137
rect 933 -3145 934 -3143
rect 940 -3139 941 -3137
rect 940 -3145 941 -3143
rect 947 -3139 948 -3137
rect 947 -3145 948 -3143
rect 954 -3139 955 -3137
rect 954 -3145 955 -3143
rect 961 -3139 962 -3137
rect 961 -3145 962 -3143
rect 968 -3139 969 -3137
rect 968 -3145 969 -3143
rect 975 -3139 976 -3137
rect 975 -3145 976 -3143
rect 982 -3139 983 -3137
rect 982 -3145 983 -3143
rect 989 -3139 990 -3137
rect 989 -3145 990 -3143
rect 996 -3139 997 -3137
rect 996 -3145 997 -3143
rect 1003 -3139 1004 -3137
rect 1003 -3145 1004 -3143
rect 1010 -3139 1011 -3137
rect 1010 -3145 1011 -3143
rect 1017 -3139 1018 -3137
rect 1017 -3145 1018 -3143
rect 1024 -3139 1025 -3137
rect 1024 -3145 1025 -3143
rect 1031 -3139 1032 -3137
rect 1031 -3145 1032 -3143
rect 1038 -3139 1039 -3137
rect 1038 -3145 1039 -3143
rect 1045 -3139 1046 -3137
rect 1045 -3145 1046 -3143
rect 1052 -3139 1053 -3137
rect 1052 -3145 1053 -3143
rect 1059 -3139 1060 -3137
rect 1059 -3145 1060 -3143
rect 1066 -3139 1067 -3137
rect 1066 -3145 1067 -3143
rect 1073 -3139 1074 -3137
rect 1073 -3145 1074 -3143
rect 1080 -3139 1081 -3137
rect 1080 -3145 1081 -3143
rect 1087 -3139 1088 -3137
rect 1087 -3145 1088 -3143
rect 1094 -3139 1095 -3137
rect 1094 -3145 1095 -3143
rect 1101 -3139 1102 -3137
rect 1101 -3145 1102 -3143
rect 1108 -3139 1109 -3137
rect 1108 -3145 1109 -3143
rect 1115 -3139 1116 -3137
rect 1115 -3145 1116 -3143
rect 1122 -3139 1123 -3137
rect 1122 -3145 1123 -3143
rect 1129 -3139 1130 -3137
rect 1129 -3145 1130 -3143
rect 1136 -3139 1137 -3137
rect 1136 -3145 1137 -3143
rect 1143 -3139 1144 -3137
rect 1143 -3145 1144 -3143
rect 1150 -3139 1151 -3137
rect 1150 -3145 1151 -3143
rect 1157 -3139 1158 -3137
rect 1157 -3145 1158 -3143
rect 1164 -3139 1165 -3137
rect 1164 -3145 1165 -3143
rect 1171 -3139 1172 -3137
rect 1171 -3145 1172 -3143
rect 1178 -3139 1179 -3137
rect 1178 -3145 1179 -3143
rect 1185 -3139 1186 -3137
rect 1185 -3145 1186 -3143
rect 1192 -3139 1193 -3137
rect 1192 -3145 1193 -3143
rect 1202 -3139 1203 -3137
rect 1199 -3145 1200 -3143
rect 1202 -3145 1203 -3143
rect 1209 -3139 1210 -3137
rect 1206 -3145 1207 -3143
rect 1209 -3145 1210 -3143
rect 1213 -3139 1214 -3137
rect 1213 -3145 1214 -3143
rect 1220 -3139 1221 -3137
rect 1220 -3145 1221 -3143
rect 1227 -3139 1228 -3137
rect 1227 -3145 1228 -3143
rect 1234 -3139 1235 -3137
rect 1234 -3145 1235 -3143
rect 1241 -3139 1242 -3137
rect 1241 -3145 1242 -3143
rect 1248 -3139 1249 -3137
rect 1248 -3145 1249 -3143
rect 1255 -3139 1256 -3137
rect 1255 -3145 1256 -3143
rect 1262 -3139 1263 -3137
rect 1262 -3145 1263 -3143
rect 1269 -3139 1270 -3137
rect 1269 -3145 1270 -3143
rect 1276 -3139 1277 -3137
rect 1276 -3145 1277 -3143
rect 1283 -3139 1284 -3137
rect 1283 -3145 1284 -3143
rect 1290 -3139 1291 -3137
rect 1290 -3145 1291 -3143
rect 1297 -3139 1298 -3137
rect 1297 -3145 1298 -3143
rect 1304 -3139 1305 -3137
rect 1304 -3145 1305 -3143
rect 1311 -3139 1312 -3137
rect 1311 -3145 1312 -3143
rect 1318 -3139 1319 -3137
rect 1318 -3145 1319 -3143
rect 1325 -3139 1326 -3137
rect 1325 -3145 1326 -3143
rect 1332 -3139 1333 -3137
rect 1335 -3139 1336 -3137
rect 1332 -3145 1333 -3143
rect 1335 -3145 1336 -3143
rect 1339 -3139 1340 -3137
rect 1339 -3145 1340 -3143
rect 1353 -3139 1354 -3137
rect 1353 -3145 1354 -3143
rect 1360 -3139 1361 -3137
rect 1360 -3145 1361 -3143
rect 1367 -3139 1368 -3137
rect 1367 -3145 1368 -3143
rect 1374 -3139 1375 -3137
rect 1374 -3145 1375 -3143
rect 163 -3232 164 -3230
rect 163 -3238 164 -3236
rect 170 -3232 171 -3230
rect 170 -3238 171 -3236
rect 177 -3232 178 -3230
rect 177 -3238 178 -3236
rect 184 -3232 185 -3230
rect 187 -3232 188 -3230
rect 184 -3238 185 -3236
rect 187 -3238 188 -3236
rect 191 -3232 192 -3230
rect 191 -3238 192 -3236
rect 198 -3232 199 -3230
rect 198 -3238 199 -3236
rect 205 -3232 206 -3230
rect 205 -3238 206 -3236
rect 212 -3232 213 -3230
rect 212 -3238 213 -3236
rect 219 -3232 220 -3230
rect 219 -3238 220 -3236
rect 226 -3232 227 -3230
rect 226 -3238 227 -3236
rect 233 -3232 234 -3230
rect 233 -3238 234 -3236
rect 240 -3232 241 -3230
rect 240 -3238 241 -3236
rect 247 -3232 248 -3230
rect 247 -3238 248 -3236
rect 254 -3232 255 -3230
rect 254 -3238 255 -3236
rect 261 -3232 262 -3230
rect 261 -3238 262 -3236
rect 268 -3232 269 -3230
rect 268 -3238 269 -3236
rect 275 -3232 276 -3230
rect 275 -3238 276 -3236
rect 282 -3232 283 -3230
rect 285 -3232 286 -3230
rect 282 -3238 283 -3236
rect 289 -3232 290 -3230
rect 289 -3238 290 -3236
rect 296 -3232 297 -3230
rect 296 -3238 297 -3236
rect 303 -3232 304 -3230
rect 303 -3238 304 -3236
rect 310 -3232 311 -3230
rect 310 -3238 311 -3236
rect 317 -3232 318 -3230
rect 317 -3238 318 -3236
rect 324 -3232 325 -3230
rect 324 -3238 325 -3236
rect 331 -3232 332 -3230
rect 331 -3238 332 -3236
rect 338 -3232 339 -3230
rect 338 -3238 339 -3236
rect 345 -3232 346 -3230
rect 345 -3238 346 -3236
rect 352 -3232 353 -3230
rect 352 -3238 353 -3236
rect 359 -3232 360 -3230
rect 359 -3238 360 -3236
rect 366 -3232 367 -3230
rect 366 -3238 367 -3236
rect 373 -3232 374 -3230
rect 373 -3238 374 -3236
rect 380 -3232 381 -3230
rect 380 -3238 381 -3236
rect 387 -3232 388 -3230
rect 387 -3238 388 -3236
rect 394 -3232 395 -3230
rect 394 -3238 395 -3236
rect 401 -3232 402 -3230
rect 401 -3238 402 -3236
rect 408 -3232 409 -3230
rect 408 -3238 409 -3236
rect 415 -3232 416 -3230
rect 415 -3238 416 -3236
rect 422 -3232 423 -3230
rect 422 -3238 423 -3236
rect 429 -3232 430 -3230
rect 429 -3238 430 -3236
rect 436 -3232 437 -3230
rect 436 -3238 437 -3236
rect 443 -3232 444 -3230
rect 443 -3238 444 -3236
rect 450 -3232 451 -3230
rect 450 -3238 451 -3236
rect 457 -3232 458 -3230
rect 460 -3232 461 -3230
rect 457 -3238 458 -3236
rect 460 -3238 461 -3236
rect 464 -3232 465 -3230
rect 464 -3238 465 -3236
rect 471 -3232 472 -3230
rect 471 -3238 472 -3236
rect 478 -3232 479 -3230
rect 478 -3238 479 -3236
rect 481 -3238 482 -3236
rect 485 -3232 486 -3230
rect 485 -3238 486 -3236
rect 492 -3232 493 -3230
rect 492 -3238 493 -3236
rect 499 -3232 500 -3230
rect 499 -3238 500 -3236
rect 506 -3232 507 -3230
rect 506 -3238 507 -3236
rect 513 -3232 514 -3230
rect 513 -3238 514 -3236
rect 520 -3232 521 -3230
rect 520 -3238 521 -3236
rect 527 -3232 528 -3230
rect 527 -3238 528 -3236
rect 534 -3232 535 -3230
rect 534 -3238 535 -3236
rect 544 -3232 545 -3230
rect 541 -3238 542 -3236
rect 544 -3238 545 -3236
rect 548 -3232 549 -3230
rect 548 -3238 549 -3236
rect 555 -3232 556 -3230
rect 555 -3238 556 -3236
rect 562 -3232 563 -3230
rect 562 -3238 563 -3236
rect 569 -3232 570 -3230
rect 569 -3238 570 -3236
rect 576 -3232 577 -3230
rect 579 -3238 580 -3236
rect 583 -3232 584 -3230
rect 583 -3238 584 -3236
rect 590 -3232 591 -3230
rect 590 -3238 591 -3236
rect 597 -3232 598 -3230
rect 597 -3238 598 -3236
rect 604 -3232 605 -3230
rect 604 -3238 605 -3236
rect 611 -3232 612 -3230
rect 611 -3238 612 -3236
rect 618 -3232 619 -3230
rect 618 -3238 619 -3236
rect 625 -3232 626 -3230
rect 625 -3238 626 -3236
rect 632 -3232 633 -3230
rect 635 -3232 636 -3230
rect 639 -3232 640 -3230
rect 639 -3238 640 -3236
rect 646 -3232 647 -3230
rect 646 -3238 647 -3236
rect 653 -3232 654 -3230
rect 653 -3238 654 -3236
rect 660 -3232 661 -3230
rect 660 -3238 661 -3236
rect 667 -3232 668 -3230
rect 667 -3238 668 -3236
rect 674 -3232 675 -3230
rect 674 -3238 675 -3236
rect 681 -3232 682 -3230
rect 681 -3238 682 -3236
rect 688 -3232 689 -3230
rect 688 -3238 689 -3236
rect 695 -3232 696 -3230
rect 695 -3238 696 -3236
rect 702 -3232 703 -3230
rect 702 -3238 703 -3236
rect 709 -3232 710 -3230
rect 709 -3238 710 -3236
rect 712 -3238 713 -3236
rect 716 -3232 717 -3230
rect 716 -3238 717 -3236
rect 723 -3232 724 -3230
rect 723 -3238 724 -3236
rect 730 -3232 731 -3230
rect 730 -3238 731 -3236
rect 737 -3232 738 -3230
rect 737 -3238 738 -3236
rect 744 -3232 745 -3230
rect 747 -3232 748 -3230
rect 744 -3238 745 -3236
rect 747 -3238 748 -3236
rect 751 -3232 752 -3230
rect 754 -3232 755 -3230
rect 751 -3238 752 -3236
rect 754 -3238 755 -3236
rect 758 -3232 759 -3230
rect 758 -3238 759 -3236
rect 765 -3232 766 -3230
rect 768 -3232 769 -3230
rect 768 -3238 769 -3236
rect 772 -3232 773 -3230
rect 772 -3238 773 -3236
rect 779 -3232 780 -3230
rect 779 -3238 780 -3236
rect 786 -3232 787 -3230
rect 786 -3238 787 -3236
rect 793 -3232 794 -3230
rect 793 -3238 794 -3236
rect 800 -3232 801 -3230
rect 800 -3238 801 -3236
rect 807 -3232 808 -3230
rect 810 -3232 811 -3230
rect 807 -3238 808 -3236
rect 810 -3238 811 -3236
rect 814 -3232 815 -3230
rect 814 -3238 815 -3236
rect 821 -3232 822 -3230
rect 821 -3238 822 -3236
rect 828 -3232 829 -3230
rect 828 -3238 829 -3236
rect 835 -3232 836 -3230
rect 835 -3238 836 -3236
rect 842 -3232 843 -3230
rect 842 -3238 843 -3236
rect 849 -3232 850 -3230
rect 849 -3238 850 -3236
rect 856 -3232 857 -3230
rect 856 -3238 857 -3236
rect 863 -3232 864 -3230
rect 863 -3238 864 -3236
rect 870 -3232 871 -3230
rect 870 -3238 871 -3236
rect 877 -3232 878 -3230
rect 877 -3238 878 -3236
rect 884 -3232 885 -3230
rect 884 -3238 885 -3236
rect 891 -3232 892 -3230
rect 894 -3232 895 -3230
rect 891 -3238 892 -3236
rect 898 -3232 899 -3230
rect 898 -3238 899 -3236
rect 905 -3232 906 -3230
rect 905 -3238 906 -3236
rect 912 -3232 913 -3230
rect 912 -3238 913 -3236
rect 919 -3232 920 -3230
rect 919 -3238 920 -3236
rect 926 -3232 927 -3230
rect 926 -3238 927 -3236
rect 933 -3232 934 -3230
rect 933 -3238 934 -3236
rect 940 -3232 941 -3230
rect 943 -3232 944 -3230
rect 940 -3238 941 -3236
rect 947 -3232 948 -3230
rect 947 -3238 948 -3236
rect 954 -3232 955 -3230
rect 954 -3238 955 -3236
rect 961 -3232 962 -3230
rect 961 -3238 962 -3236
rect 964 -3238 965 -3236
rect 968 -3232 969 -3230
rect 968 -3238 969 -3236
rect 975 -3232 976 -3230
rect 975 -3238 976 -3236
rect 982 -3232 983 -3230
rect 982 -3238 983 -3236
rect 989 -3232 990 -3230
rect 989 -3238 990 -3236
rect 996 -3232 997 -3230
rect 996 -3238 997 -3236
rect 1003 -3232 1004 -3230
rect 1003 -3238 1004 -3236
rect 1010 -3232 1011 -3230
rect 1010 -3238 1011 -3236
rect 1017 -3232 1018 -3230
rect 1017 -3238 1018 -3236
rect 1024 -3232 1025 -3230
rect 1024 -3238 1025 -3236
rect 1031 -3232 1032 -3230
rect 1031 -3238 1032 -3236
rect 1038 -3232 1039 -3230
rect 1038 -3238 1039 -3236
rect 1045 -3232 1046 -3230
rect 1045 -3238 1046 -3236
rect 1052 -3232 1053 -3230
rect 1052 -3238 1053 -3236
rect 1059 -3232 1060 -3230
rect 1059 -3238 1060 -3236
rect 1066 -3232 1067 -3230
rect 1066 -3238 1067 -3236
rect 1073 -3232 1074 -3230
rect 1073 -3238 1074 -3236
rect 1080 -3232 1081 -3230
rect 1080 -3238 1081 -3236
rect 1087 -3232 1088 -3230
rect 1087 -3238 1088 -3236
rect 1094 -3232 1095 -3230
rect 1094 -3238 1095 -3236
rect 1101 -3232 1102 -3230
rect 1101 -3238 1102 -3236
rect 1108 -3232 1109 -3230
rect 1108 -3238 1109 -3236
rect 1115 -3232 1116 -3230
rect 1115 -3238 1116 -3236
rect 1122 -3232 1123 -3230
rect 1122 -3238 1123 -3236
rect 1129 -3232 1130 -3230
rect 1129 -3238 1130 -3236
rect 1136 -3232 1137 -3230
rect 1136 -3238 1137 -3236
rect 1143 -3232 1144 -3230
rect 1143 -3238 1144 -3236
rect 1150 -3232 1151 -3230
rect 1150 -3238 1151 -3236
rect 1157 -3232 1158 -3230
rect 1157 -3238 1158 -3236
rect 1164 -3232 1165 -3230
rect 1167 -3232 1168 -3230
rect 1164 -3238 1165 -3236
rect 1171 -3232 1172 -3230
rect 1171 -3238 1172 -3236
rect 1178 -3232 1179 -3230
rect 1178 -3238 1179 -3236
rect 1185 -3232 1186 -3230
rect 1185 -3238 1186 -3236
rect 1192 -3232 1193 -3230
rect 1192 -3238 1193 -3236
rect 1199 -3232 1200 -3230
rect 1202 -3232 1203 -3230
rect 1202 -3238 1203 -3236
rect 1206 -3232 1207 -3230
rect 1206 -3238 1207 -3236
rect 1213 -3232 1214 -3230
rect 1213 -3238 1214 -3236
rect 1220 -3232 1221 -3230
rect 1220 -3238 1221 -3236
rect 1230 -3232 1231 -3230
rect 1227 -3238 1228 -3236
rect 1234 -3232 1235 -3230
rect 1234 -3238 1235 -3236
rect 1241 -3232 1242 -3230
rect 1241 -3238 1242 -3236
rect 1248 -3232 1249 -3230
rect 1248 -3238 1249 -3236
rect 1255 -3232 1256 -3230
rect 1255 -3238 1256 -3236
rect 1258 -3238 1259 -3236
rect 1262 -3232 1263 -3230
rect 1262 -3238 1263 -3236
rect 1269 -3232 1270 -3230
rect 1269 -3238 1270 -3236
rect 1276 -3232 1277 -3230
rect 1276 -3238 1277 -3236
rect 1283 -3232 1284 -3230
rect 1286 -3232 1287 -3230
rect 1283 -3238 1284 -3236
rect 1290 -3232 1291 -3230
rect 1293 -3232 1294 -3230
rect 1293 -3238 1294 -3236
rect 1297 -3232 1298 -3230
rect 1297 -3238 1298 -3236
rect 1304 -3232 1305 -3230
rect 1304 -3238 1305 -3236
rect 1346 -3232 1347 -3230
rect 1346 -3238 1347 -3236
rect 1353 -3232 1354 -3230
rect 1353 -3238 1354 -3236
rect 1360 -3232 1361 -3230
rect 1360 -3238 1361 -3236
rect 156 -3309 157 -3307
rect 156 -3315 157 -3313
rect 163 -3309 164 -3307
rect 163 -3315 164 -3313
rect 170 -3309 171 -3307
rect 170 -3315 171 -3313
rect 177 -3309 178 -3307
rect 177 -3315 178 -3313
rect 184 -3309 185 -3307
rect 184 -3315 185 -3313
rect 191 -3309 192 -3307
rect 191 -3315 192 -3313
rect 198 -3309 199 -3307
rect 201 -3309 202 -3307
rect 205 -3309 206 -3307
rect 205 -3315 206 -3313
rect 212 -3309 213 -3307
rect 212 -3315 213 -3313
rect 219 -3309 220 -3307
rect 219 -3315 220 -3313
rect 226 -3309 227 -3307
rect 226 -3315 227 -3313
rect 233 -3309 234 -3307
rect 233 -3315 234 -3313
rect 243 -3309 244 -3307
rect 243 -3315 244 -3313
rect 247 -3309 248 -3307
rect 247 -3315 248 -3313
rect 254 -3309 255 -3307
rect 254 -3315 255 -3313
rect 261 -3309 262 -3307
rect 261 -3315 262 -3313
rect 268 -3309 269 -3307
rect 268 -3315 269 -3313
rect 275 -3309 276 -3307
rect 275 -3315 276 -3313
rect 282 -3309 283 -3307
rect 282 -3315 283 -3313
rect 289 -3309 290 -3307
rect 289 -3315 290 -3313
rect 296 -3309 297 -3307
rect 296 -3315 297 -3313
rect 303 -3309 304 -3307
rect 303 -3315 304 -3313
rect 310 -3309 311 -3307
rect 310 -3315 311 -3313
rect 317 -3309 318 -3307
rect 317 -3315 318 -3313
rect 324 -3309 325 -3307
rect 324 -3315 325 -3313
rect 331 -3309 332 -3307
rect 331 -3315 332 -3313
rect 338 -3309 339 -3307
rect 338 -3315 339 -3313
rect 345 -3309 346 -3307
rect 345 -3315 346 -3313
rect 352 -3309 353 -3307
rect 352 -3315 353 -3313
rect 359 -3309 360 -3307
rect 359 -3315 360 -3313
rect 366 -3309 367 -3307
rect 366 -3315 367 -3313
rect 373 -3309 374 -3307
rect 373 -3315 374 -3313
rect 380 -3309 381 -3307
rect 380 -3315 381 -3313
rect 387 -3309 388 -3307
rect 387 -3315 388 -3313
rect 394 -3309 395 -3307
rect 394 -3315 395 -3313
rect 401 -3309 402 -3307
rect 401 -3315 402 -3313
rect 408 -3309 409 -3307
rect 408 -3315 409 -3313
rect 415 -3309 416 -3307
rect 415 -3315 416 -3313
rect 422 -3309 423 -3307
rect 422 -3315 423 -3313
rect 429 -3309 430 -3307
rect 429 -3315 430 -3313
rect 436 -3309 437 -3307
rect 436 -3315 437 -3313
rect 443 -3309 444 -3307
rect 443 -3315 444 -3313
rect 450 -3309 451 -3307
rect 450 -3315 451 -3313
rect 457 -3309 458 -3307
rect 457 -3315 458 -3313
rect 464 -3309 465 -3307
rect 464 -3315 465 -3313
rect 471 -3309 472 -3307
rect 471 -3315 472 -3313
rect 478 -3309 479 -3307
rect 478 -3315 479 -3313
rect 485 -3309 486 -3307
rect 488 -3309 489 -3307
rect 485 -3315 486 -3313
rect 492 -3309 493 -3307
rect 492 -3315 493 -3313
rect 499 -3309 500 -3307
rect 499 -3315 500 -3313
rect 506 -3309 507 -3307
rect 506 -3315 507 -3313
rect 513 -3309 514 -3307
rect 513 -3315 514 -3313
rect 520 -3309 521 -3307
rect 520 -3315 521 -3313
rect 527 -3309 528 -3307
rect 527 -3315 528 -3313
rect 537 -3309 538 -3307
rect 534 -3315 535 -3313
rect 537 -3315 538 -3313
rect 541 -3309 542 -3307
rect 541 -3315 542 -3313
rect 548 -3309 549 -3307
rect 548 -3315 549 -3313
rect 555 -3309 556 -3307
rect 555 -3315 556 -3313
rect 562 -3309 563 -3307
rect 562 -3315 563 -3313
rect 569 -3309 570 -3307
rect 569 -3315 570 -3313
rect 576 -3309 577 -3307
rect 576 -3315 577 -3313
rect 583 -3309 584 -3307
rect 583 -3315 584 -3313
rect 590 -3309 591 -3307
rect 590 -3315 591 -3313
rect 597 -3309 598 -3307
rect 597 -3315 598 -3313
rect 604 -3309 605 -3307
rect 604 -3315 605 -3313
rect 611 -3309 612 -3307
rect 614 -3309 615 -3307
rect 614 -3315 615 -3313
rect 618 -3309 619 -3307
rect 618 -3315 619 -3313
rect 625 -3309 626 -3307
rect 625 -3315 626 -3313
rect 632 -3309 633 -3307
rect 632 -3315 633 -3313
rect 639 -3309 640 -3307
rect 639 -3315 640 -3313
rect 646 -3309 647 -3307
rect 646 -3315 647 -3313
rect 653 -3309 654 -3307
rect 656 -3309 657 -3307
rect 653 -3315 654 -3313
rect 656 -3315 657 -3313
rect 660 -3309 661 -3307
rect 663 -3309 664 -3307
rect 660 -3315 661 -3313
rect 663 -3315 664 -3313
rect 667 -3309 668 -3307
rect 670 -3309 671 -3307
rect 667 -3315 668 -3313
rect 670 -3315 671 -3313
rect 674 -3309 675 -3307
rect 674 -3315 675 -3313
rect 681 -3309 682 -3307
rect 681 -3315 682 -3313
rect 688 -3309 689 -3307
rect 691 -3309 692 -3307
rect 688 -3315 689 -3313
rect 691 -3315 692 -3313
rect 695 -3309 696 -3307
rect 695 -3315 696 -3313
rect 702 -3309 703 -3307
rect 702 -3315 703 -3313
rect 709 -3309 710 -3307
rect 709 -3315 710 -3313
rect 716 -3309 717 -3307
rect 716 -3315 717 -3313
rect 723 -3309 724 -3307
rect 723 -3315 724 -3313
rect 733 -3309 734 -3307
rect 730 -3315 731 -3313
rect 737 -3309 738 -3307
rect 737 -3315 738 -3313
rect 744 -3309 745 -3307
rect 744 -3315 745 -3313
rect 751 -3309 752 -3307
rect 751 -3315 752 -3313
rect 758 -3309 759 -3307
rect 758 -3315 759 -3313
rect 761 -3315 762 -3313
rect 765 -3309 766 -3307
rect 765 -3315 766 -3313
rect 772 -3309 773 -3307
rect 772 -3315 773 -3313
rect 779 -3309 780 -3307
rect 779 -3315 780 -3313
rect 786 -3309 787 -3307
rect 786 -3315 787 -3313
rect 793 -3309 794 -3307
rect 793 -3315 794 -3313
rect 800 -3309 801 -3307
rect 800 -3315 801 -3313
rect 807 -3309 808 -3307
rect 807 -3315 808 -3313
rect 814 -3309 815 -3307
rect 814 -3315 815 -3313
rect 821 -3309 822 -3307
rect 824 -3309 825 -3307
rect 824 -3315 825 -3313
rect 828 -3309 829 -3307
rect 828 -3315 829 -3313
rect 838 -3309 839 -3307
rect 835 -3315 836 -3313
rect 838 -3315 839 -3313
rect 842 -3309 843 -3307
rect 842 -3315 843 -3313
rect 849 -3309 850 -3307
rect 849 -3315 850 -3313
rect 859 -3309 860 -3307
rect 856 -3315 857 -3313
rect 859 -3315 860 -3313
rect 863 -3309 864 -3307
rect 863 -3315 864 -3313
rect 873 -3309 874 -3307
rect 870 -3315 871 -3313
rect 873 -3315 874 -3313
rect 877 -3309 878 -3307
rect 877 -3315 878 -3313
rect 884 -3309 885 -3307
rect 884 -3315 885 -3313
rect 891 -3309 892 -3307
rect 894 -3309 895 -3307
rect 891 -3315 892 -3313
rect 894 -3315 895 -3313
rect 898 -3309 899 -3307
rect 898 -3315 899 -3313
rect 905 -3309 906 -3307
rect 905 -3315 906 -3313
rect 912 -3309 913 -3307
rect 912 -3315 913 -3313
rect 919 -3309 920 -3307
rect 919 -3315 920 -3313
rect 926 -3309 927 -3307
rect 926 -3315 927 -3313
rect 933 -3309 934 -3307
rect 933 -3315 934 -3313
rect 940 -3309 941 -3307
rect 940 -3315 941 -3313
rect 947 -3309 948 -3307
rect 947 -3315 948 -3313
rect 954 -3309 955 -3307
rect 954 -3315 955 -3313
rect 961 -3309 962 -3307
rect 961 -3315 962 -3313
rect 968 -3309 969 -3307
rect 968 -3315 969 -3313
rect 975 -3309 976 -3307
rect 975 -3315 976 -3313
rect 982 -3309 983 -3307
rect 982 -3315 983 -3313
rect 989 -3309 990 -3307
rect 989 -3315 990 -3313
rect 996 -3309 997 -3307
rect 996 -3315 997 -3313
rect 1003 -3309 1004 -3307
rect 1006 -3309 1007 -3307
rect 1003 -3315 1004 -3313
rect 1010 -3309 1011 -3307
rect 1010 -3315 1011 -3313
rect 1017 -3309 1018 -3307
rect 1017 -3315 1018 -3313
rect 1024 -3309 1025 -3307
rect 1027 -3309 1028 -3307
rect 1027 -3315 1028 -3313
rect 1031 -3309 1032 -3307
rect 1031 -3315 1032 -3313
rect 1038 -3309 1039 -3307
rect 1038 -3315 1039 -3313
rect 1045 -3309 1046 -3307
rect 1045 -3315 1046 -3313
rect 1052 -3309 1053 -3307
rect 1052 -3315 1053 -3313
rect 1059 -3309 1060 -3307
rect 1059 -3315 1060 -3313
rect 1066 -3309 1067 -3307
rect 1066 -3315 1067 -3313
rect 1073 -3309 1074 -3307
rect 1073 -3315 1074 -3313
rect 1080 -3309 1081 -3307
rect 1080 -3315 1081 -3313
rect 1087 -3309 1088 -3307
rect 1087 -3315 1088 -3313
rect 1094 -3309 1095 -3307
rect 1094 -3315 1095 -3313
rect 1101 -3309 1102 -3307
rect 1101 -3315 1102 -3313
rect 1108 -3309 1109 -3307
rect 1108 -3315 1109 -3313
rect 1115 -3309 1116 -3307
rect 1115 -3315 1116 -3313
rect 1122 -3309 1123 -3307
rect 1122 -3315 1123 -3313
rect 1129 -3309 1130 -3307
rect 1129 -3315 1130 -3313
rect 1136 -3309 1137 -3307
rect 1136 -3315 1137 -3313
rect 1139 -3315 1140 -3313
rect 1143 -3309 1144 -3307
rect 1143 -3315 1144 -3313
rect 1150 -3309 1151 -3307
rect 1150 -3315 1151 -3313
rect 1157 -3309 1158 -3307
rect 1157 -3315 1158 -3313
rect 1164 -3309 1165 -3307
rect 1164 -3315 1165 -3313
rect 1171 -3309 1172 -3307
rect 1171 -3315 1172 -3313
rect 1178 -3309 1179 -3307
rect 1178 -3315 1179 -3313
rect 1185 -3309 1186 -3307
rect 1185 -3315 1186 -3313
rect 1192 -3309 1193 -3307
rect 1192 -3315 1193 -3313
rect 1199 -3309 1200 -3307
rect 1199 -3315 1200 -3313
rect 1206 -3309 1207 -3307
rect 1206 -3315 1207 -3313
rect 1213 -3309 1214 -3307
rect 1213 -3315 1214 -3313
rect 1220 -3309 1221 -3307
rect 1220 -3315 1221 -3313
rect 1227 -3309 1228 -3307
rect 1227 -3315 1228 -3313
rect 1234 -3309 1235 -3307
rect 1234 -3315 1235 -3313
rect 1241 -3309 1242 -3307
rect 1241 -3315 1242 -3313
rect 1248 -3309 1249 -3307
rect 1248 -3315 1249 -3313
rect 1255 -3309 1256 -3307
rect 1255 -3315 1256 -3313
rect 1262 -3309 1263 -3307
rect 1262 -3315 1263 -3313
rect 1272 -3309 1273 -3307
rect 1269 -3315 1270 -3313
rect 1272 -3315 1273 -3313
rect 1276 -3309 1277 -3307
rect 1276 -3315 1277 -3313
rect 1290 -3309 1291 -3307
rect 1290 -3315 1291 -3313
rect 1339 -3309 1340 -3307
rect 1339 -3315 1340 -3313
rect 1346 -3309 1347 -3307
rect 1346 -3315 1347 -3313
rect 1353 -3309 1354 -3307
rect 1353 -3315 1354 -3313
rect 198 -3382 199 -3380
rect 198 -3388 199 -3386
rect 205 -3382 206 -3380
rect 205 -3388 206 -3386
rect 212 -3382 213 -3380
rect 212 -3388 213 -3386
rect 219 -3382 220 -3380
rect 219 -3388 220 -3386
rect 226 -3382 227 -3380
rect 226 -3388 227 -3386
rect 233 -3382 234 -3380
rect 233 -3388 234 -3386
rect 240 -3382 241 -3380
rect 240 -3388 241 -3386
rect 247 -3382 248 -3380
rect 247 -3388 248 -3386
rect 254 -3382 255 -3380
rect 254 -3388 255 -3386
rect 261 -3388 262 -3386
rect 271 -3382 272 -3380
rect 268 -3388 269 -3386
rect 271 -3388 272 -3386
rect 275 -3382 276 -3380
rect 278 -3388 279 -3386
rect 282 -3382 283 -3380
rect 282 -3388 283 -3386
rect 289 -3382 290 -3380
rect 289 -3388 290 -3386
rect 296 -3382 297 -3380
rect 296 -3388 297 -3386
rect 303 -3382 304 -3380
rect 303 -3388 304 -3386
rect 310 -3382 311 -3380
rect 310 -3388 311 -3386
rect 317 -3382 318 -3380
rect 317 -3388 318 -3386
rect 324 -3382 325 -3380
rect 324 -3388 325 -3386
rect 331 -3382 332 -3380
rect 331 -3388 332 -3386
rect 338 -3382 339 -3380
rect 338 -3388 339 -3386
rect 345 -3382 346 -3380
rect 345 -3388 346 -3386
rect 352 -3382 353 -3380
rect 352 -3388 353 -3386
rect 359 -3382 360 -3380
rect 359 -3388 360 -3386
rect 366 -3382 367 -3380
rect 366 -3388 367 -3386
rect 373 -3382 374 -3380
rect 373 -3388 374 -3386
rect 380 -3382 381 -3380
rect 380 -3388 381 -3386
rect 387 -3382 388 -3380
rect 387 -3388 388 -3386
rect 394 -3382 395 -3380
rect 394 -3388 395 -3386
rect 401 -3382 402 -3380
rect 404 -3382 405 -3380
rect 404 -3388 405 -3386
rect 408 -3382 409 -3380
rect 411 -3382 412 -3380
rect 408 -3388 409 -3386
rect 411 -3388 412 -3386
rect 415 -3382 416 -3380
rect 415 -3388 416 -3386
rect 422 -3382 423 -3380
rect 425 -3382 426 -3380
rect 422 -3388 423 -3386
rect 429 -3382 430 -3380
rect 429 -3388 430 -3386
rect 436 -3382 437 -3380
rect 436 -3388 437 -3386
rect 443 -3382 444 -3380
rect 443 -3388 444 -3386
rect 450 -3382 451 -3380
rect 450 -3388 451 -3386
rect 457 -3382 458 -3380
rect 457 -3388 458 -3386
rect 464 -3382 465 -3380
rect 464 -3388 465 -3386
rect 471 -3382 472 -3380
rect 471 -3388 472 -3386
rect 474 -3388 475 -3386
rect 478 -3382 479 -3380
rect 478 -3388 479 -3386
rect 485 -3382 486 -3380
rect 485 -3388 486 -3386
rect 492 -3382 493 -3380
rect 492 -3388 493 -3386
rect 499 -3382 500 -3380
rect 499 -3388 500 -3386
rect 506 -3382 507 -3380
rect 506 -3388 507 -3386
rect 513 -3382 514 -3380
rect 513 -3388 514 -3386
rect 520 -3382 521 -3380
rect 520 -3388 521 -3386
rect 527 -3382 528 -3380
rect 534 -3382 535 -3380
rect 534 -3388 535 -3386
rect 541 -3382 542 -3380
rect 544 -3382 545 -3380
rect 541 -3388 542 -3386
rect 548 -3382 549 -3380
rect 548 -3388 549 -3386
rect 555 -3382 556 -3380
rect 558 -3382 559 -3380
rect 558 -3388 559 -3386
rect 562 -3382 563 -3380
rect 562 -3388 563 -3386
rect 569 -3382 570 -3380
rect 572 -3382 573 -3380
rect 569 -3388 570 -3386
rect 572 -3388 573 -3386
rect 576 -3382 577 -3380
rect 579 -3382 580 -3380
rect 576 -3388 577 -3386
rect 579 -3388 580 -3386
rect 583 -3382 584 -3380
rect 583 -3388 584 -3386
rect 590 -3382 591 -3380
rect 590 -3388 591 -3386
rect 597 -3382 598 -3380
rect 597 -3388 598 -3386
rect 604 -3382 605 -3380
rect 604 -3388 605 -3386
rect 611 -3382 612 -3380
rect 611 -3388 612 -3386
rect 618 -3382 619 -3380
rect 618 -3388 619 -3386
rect 625 -3382 626 -3380
rect 625 -3388 626 -3386
rect 632 -3382 633 -3380
rect 632 -3388 633 -3386
rect 639 -3382 640 -3380
rect 639 -3388 640 -3386
rect 646 -3382 647 -3380
rect 646 -3388 647 -3386
rect 653 -3382 654 -3380
rect 656 -3382 657 -3380
rect 656 -3388 657 -3386
rect 660 -3382 661 -3380
rect 660 -3388 661 -3386
rect 667 -3382 668 -3380
rect 667 -3388 668 -3386
rect 674 -3382 675 -3380
rect 674 -3388 675 -3386
rect 681 -3382 682 -3380
rect 681 -3388 682 -3386
rect 688 -3382 689 -3380
rect 688 -3388 689 -3386
rect 695 -3382 696 -3380
rect 695 -3388 696 -3386
rect 702 -3382 703 -3380
rect 702 -3388 703 -3386
rect 709 -3382 710 -3380
rect 709 -3388 710 -3386
rect 716 -3382 717 -3380
rect 716 -3388 717 -3386
rect 723 -3382 724 -3380
rect 723 -3388 724 -3386
rect 730 -3382 731 -3380
rect 730 -3388 731 -3386
rect 737 -3382 738 -3380
rect 737 -3388 738 -3386
rect 744 -3382 745 -3380
rect 744 -3388 745 -3386
rect 751 -3382 752 -3380
rect 751 -3388 752 -3386
rect 761 -3382 762 -3380
rect 758 -3388 759 -3386
rect 765 -3382 766 -3380
rect 765 -3388 766 -3386
rect 772 -3382 773 -3380
rect 772 -3388 773 -3386
rect 779 -3382 780 -3380
rect 779 -3388 780 -3386
rect 786 -3382 787 -3380
rect 786 -3388 787 -3386
rect 793 -3382 794 -3380
rect 793 -3388 794 -3386
rect 796 -3388 797 -3386
rect 800 -3382 801 -3380
rect 800 -3388 801 -3386
rect 807 -3382 808 -3380
rect 807 -3388 808 -3386
rect 814 -3382 815 -3380
rect 814 -3388 815 -3386
rect 821 -3382 822 -3380
rect 821 -3388 822 -3386
rect 828 -3382 829 -3380
rect 828 -3388 829 -3386
rect 835 -3382 836 -3380
rect 835 -3388 836 -3386
rect 842 -3382 843 -3380
rect 842 -3388 843 -3386
rect 849 -3382 850 -3380
rect 849 -3388 850 -3386
rect 856 -3382 857 -3380
rect 856 -3388 857 -3386
rect 863 -3382 864 -3380
rect 863 -3388 864 -3386
rect 870 -3382 871 -3380
rect 870 -3388 871 -3386
rect 877 -3382 878 -3380
rect 877 -3388 878 -3386
rect 884 -3382 885 -3380
rect 884 -3388 885 -3386
rect 891 -3382 892 -3380
rect 891 -3388 892 -3386
rect 898 -3382 899 -3380
rect 898 -3388 899 -3386
rect 905 -3382 906 -3380
rect 905 -3388 906 -3386
rect 912 -3382 913 -3380
rect 912 -3388 913 -3386
rect 919 -3382 920 -3380
rect 919 -3388 920 -3386
rect 926 -3382 927 -3380
rect 926 -3388 927 -3386
rect 933 -3382 934 -3380
rect 933 -3388 934 -3386
rect 940 -3382 941 -3380
rect 940 -3388 941 -3386
rect 947 -3382 948 -3380
rect 947 -3388 948 -3386
rect 954 -3382 955 -3380
rect 957 -3388 958 -3386
rect 961 -3382 962 -3380
rect 961 -3388 962 -3386
rect 968 -3382 969 -3380
rect 968 -3388 969 -3386
rect 975 -3382 976 -3380
rect 975 -3388 976 -3386
rect 982 -3382 983 -3380
rect 982 -3388 983 -3386
rect 989 -3382 990 -3380
rect 989 -3388 990 -3386
rect 996 -3382 997 -3380
rect 996 -3388 997 -3386
rect 1003 -3382 1004 -3380
rect 1003 -3388 1004 -3386
rect 1010 -3382 1011 -3380
rect 1013 -3382 1014 -3380
rect 1010 -3388 1011 -3386
rect 1013 -3388 1014 -3386
rect 1017 -3382 1018 -3380
rect 1017 -3388 1018 -3386
rect 1024 -3382 1025 -3380
rect 1024 -3388 1025 -3386
rect 1031 -3382 1032 -3380
rect 1031 -3388 1032 -3386
rect 1041 -3382 1042 -3380
rect 1038 -3388 1039 -3386
rect 1045 -3382 1046 -3380
rect 1045 -3388 1046 -3386
rect 1052 -3382 1053 -3380
rect 1055 -3382 1056 -3380
rect 1059 -3382 1060 -3380
rect 1059 -3388 1060 -3386
rect 1066 -3382 1067 -3380
rect 1069 -3382 1070 -3380
rect 1066 -3388 1067 -3386
rect 1073 -3382 1074 -3380
rect 1073 -3388 1074 -3386
rect 1080 -3382 1081 -3380
rect 1080 -3388 1081 -3386
rect 1087 -3382 1088 -3380
rect 1087 -3388 1088 -3386
rect 1094 -3382 1095 -3380
rect 1094 -3388 1095 -3386
rect 1101 -3382 1102 -3380
rect 1101 -3388 1102 -3386
rect 1122 -3382 1123 -3380
rect 1122 -3388 1123 -3386
rect 1129 -3382 1130 -3380
rect 1129 -3388 1130 -3386
rect 1181 -3382 1182 -3380
rect 1181 -3388 1182 -3386
rect 1185 -3382 1186 -3380
rect 1185 -3388 1186 -3386
rect 1192 -3382 1193 -3380
rect 1192 -3388 1193 -3386
rect 1339 -3382 1340 -3380
rect 1339 -3388 1340 -3386
rect 1346 -3382 1347 -3380
rect 1346 -3388 1347 -3386
rect 1349 -3388 1350 -3386
rect 1353 -3382 1354 -3380
rect 1353 -3388 1354 -3386
rect 247 -3445 248 -3443
rect 247 -3451 248 -3449
rect 261 -3445 262 -3443
rect 261 -3451 262 -3449
rect 292 -3445 293 -3443
rect 289 -3451 290 -3449
rect 292 -3451 293 -3449
rect 310 -3445 311 -3443
rect 310 -3451 311 -3449
rect 317 -3445 318 -3443
rect 317 -3451 318 -3449
rect 324 -3445 325 -3443
rect 324 -3451 325 -3449
rect 331 -3445 332 -3443
rect 331 -3451 332 -3449
rect 338 -3445 339 -3443
rect 338 -3451 339 -3449
rect 345 -3445 346 -3443
rect 348 -3445 349 -3443
rect 352 -3445 353 -3443
rect 352 -3451 353 -3449
rect 359 -3445 360 -3443
rect 359 -3451 360 -3449
rect 366 -3445 367 -3443
rect 373 -3445 374 -3443
rect 373 -3451 374 -3449
rect 380 -3445 381 -3443
rect 380 -3451 381 -3449
rect 387 -3445 388 -3443
rect 394 -3445 395 -3443
rect 394 -3451 395 -3449
rect 401 -3445 402 -3443
rect 408 -3445 409 -3443
rect 408 -3451 409 -3449
rect 415 -3445 416 -3443
rect 415 -3451 416 -3449
rect 422 -3445 423 -3443
rect 422 -3451 423 -3449
rect 429 -3445 430 -3443
rect 429 -3451 430 -3449
rect 436 -3445 437 -3443
rect 436 -3451 437 -3449
rect 446 -3445 447 -3443
rect 443 -3451 444 -3449
rect 446 -3451 447 -3449
rect 450 -3445 451 -3443
rect 450 -3451 451 -3449
rect 457 -3445 458 -3443
rect 457 -3451 458 -3449
rect 464 -3445 465 -3443
rect 464 -3451 465 -3449
rect 471 -3445 472 -3443
rect 471 -3451 472 -3449
rect 478 -3445 479 -3443
rect 478 -3451 479 -3449
rect 485 -3445 486 -3443
rect 485 -3451 486 -3449
rect 492 -3445 493 -3443
rect 492 -3451 493 -3449
rect 499 -3445 500 -3443
rect 502 -3445 503 -3443
rect 499 -3451 500 -3449
rect 506 -3445 507 -3443
rect 506 -3451 507 -3449
rect 513 -3445 514 -3443
rect 513 -3451 514 -3449
rect 520 -3445 521 -3443
rect 520 -3451 521 -3449
rect 530 -3445 531 -3443
rect 527 -3451 528 -3449
rect 530 -3451 531 -3449
rect 534 -3445 535 -3443
rect 534 -3451 535 -3449
rect 541 -3445 542 -3443
rect 541 -3451 542 -3449
rect 548 -3445 549 -3443
rect 548 -3451 549 -3449
rect 555 -3445 556 -3443
rect 555 -3451 556 -3449
rect 562 -3445 563 -3443
rect 562 -3451 563 -3449
rect 569 -3445 570 -3443
rect 569 -3451 570 -3449
rect 576 -3445 577 -3443
rect 576 -3451 577 -3449
rect 583 -3445 584 -3443
rect 583 -3451 584 -3449
rect 590 -3445 591 -3443
rect 590 -3451 591 -3449
rect 597 -3445 598 -3443
rect 597 -3451 598 -3449
rect 604 -3445 605 -3443
rect 604 -3451 605 -3449
rect 611 -3445 612 -3443
rect 611 -3451 612 -3449
rect 618 -3445 619 -3443
rect 618 -3451 619 -3449
rect 625 -3445 626 -3443
rect 625 -3451 626 -3449
rect 632 -3445 633 -3443
rect 632 -3451 633 -3449
rect 639 -3445 640 -3443
rect 639 -3451 640 -3449
rect 646 -3445 647 -3443
rect 649 -3445 650 -3443
rect 649 -3451 650 -3449
rect 653 -3445 654 -3443
rect 653 -3451 654 -3449
rect 660 -3445 661 -3443
rect 660 -3451 661 -3449
rect 667 -3445 668 -3443
rect 667 -3451 668 -3449
rect 674 -3445 675 -3443
rect 674 -3451 675 -3449
rect 681 -3445 682 -3443
rect 681 -3451 682 -3449
rect 691 -3445 692 -3443
rect 688 -3451 689 -3449
rect 691 -3451 692 -3449
rect 695 -3445 696 -3443
rect 695 -3451 696 -3449
rect 702 -3445 703 -3443
rect 702 -3451 703 -3449
rect 709 -3445 710 -3443
rect 709 -3451 710 -3449
rect 716 -3445 717 -3443
rect 716 -3451 717 -3449
rect 723 -3445 724 -3443
rect 723 -3451 724 -3449
rect 730 -3445 731 -3443
rect 730 -3451 731 -3449
rect 737 -3445 738 -3443
rect 740 -3445 741 -3443
rect 737 -3451 738 -3449
rect 740 -3451 741 -3449
rect 744 -3445 745 -3443
rect 744 -3451 745 -3449
rect 751 -3445 752 -3443
rect 751 -3451 752 -3449
rect 758 -3445 759 -3443
rect 765 -3445 766 -3443
rect 765 -3451 766 -3449
rect 772 -3445 773 -3443
rect 772 -3451 773 -3449
rect 779 -3445 780 -3443
rect 779 -3451 780 -3449
rect 786 -3445 787 -3443
rect 786 -3451 787 -3449
rect 793 -3445 794 -3443
rect 793 -3451 794 -3449
rect 800 -3445 801 -3443
rect 800 -3451 801 -3449
rect 807 -3445 808 -3443
rect 807 -3451 808 -3449
rect 814 -3445 815 -3443
rect 814 -3451 815 -3449
rect 824 -3445 825 -3443
rect 821 -3451 822 -3449
rect 824 -3451 825 -3449
rect 828 -3445 829 -3443
rect 828 -3451 829 -3449
rect 835 -3445 836 -3443
rect 835 -3451 836 -3449
rect 842 -3445 843 -3443
rect 842 -3451 843 -3449
rect 849 -3445 850 -3443
rect 849 -3451 850 -3449
rect 859 -3445 860 -3443
rect 856 -3451 857 -3449
rect 859 -3451 860 -3449
rect 863 -3445 864 -3443
rect 863 -3451 864 -3449
rect 873 -3445 874 -3443
rect 870 -3451 871 -3449
rect 877 -3445 878 -3443
rect 877 -3451 878 -3449
rect 884 -3445 885 -3443
rect 887 -3445 888 -3443
rect 884 -3451 885 -3449
rect 887 -3451 888 -3449
rect 891 -3445 892 -3443
rect 891 -3451 892 -3449
rect 898 -3451 899 -3449
rect 901 -3451 902 -3449
rect 905 -3445 906 -3443
rect 905 -3451 906 -3449
rect 912 -3445 913 -3443
rect 912 -3451 913 -3449
rect 919 -3445 920 -3443
rect 919 -3451 920 -3449
rect 926 -3445 927 -3443
rect 926 -3451 927 -3449
rect 933 -3445 934 -3443
rect 933 -3451 934 -3449
rect 936 -3451 937 -3449
rect 940 -3445 941 -3443
rect 940 -3451 941 -3449
rect 943 -3451 944 -3449
rect 947 -3445 948 -3443
rect 947 -3451 948 -3449
rect 954 -3445 955 -3443
rect 954 -3451 955 -3449
rect 961 -3445 962 -3443
rect 961 -3451 962 -3449
rect 968 -3445 969 -3443
rect 968 -3451 969 -3449
rect 975 -3445 976 -3443
rect 975 -3451 976 -3449
rect 982 -3445 983 -3443
rect 982 -3451 983 -3449
rect 1003 -3445 1004 -3443
rect 1003 -3451 1004 -3449
rect 1010 -3445 1011 -3443
rect 1010 -3451 1011 -3449
rect 1024 -3445 1025 -3443
rect 1027 -3445 1028 -3443
rect 1027 -3451 1028 -3449
rect 1031 -3445 1032 -3443
rect 1031 -3451 1032 -3449
rect 1038 -3445 1039 -3443
rect 1038 -3451 1039 -3449
rect 1045 -3445 1046 -3443
rect 1045 -3451 1046 -3449
rect 1087 -3445 1088 -3443
rect 1087 -3451 1088 -3449
rect 1094 -3445 1095 -3443
rect 1094 -3451 1095 -3449
rect 1115 -3445 1116 -3443
rect 1115 -3451 1116 -3449
rect 1136 -3445 1137 -3443
rect 1136 -3451 1137 -3449
rect 1178 -3445 1179 -3443
rect 1178 -3451 1179 -3449
rect 1339 -3445 1340 -3443
rect 1339 -3451 1340 -3449
rect 1342 -3451 1343 -3449
rect 1346 -3445 1347 -3443
rect 1349 -3445 1350 -3443
rect 1346 -3451 1347 -3449
rect 1353 -3445 1354 -3443
rect 1353 -3451 1354 -3449
rect 247 -3502 248 -3500
rect 247 -3508 248 -3506
rect 261 -3502 262 -3500
rect 261 -3508 262 -3506
rect 275 -3502 276 -3500
rect 275 -3508 276 -3506
rect 331 -3502 332 -3500
rect 331 -3508 332 -3506
rect 338 -3502 339 -3500
rect 338 -3508 339 -3506
rect 345 -3502 346 -3500
rect 345 -3508 346 -3506
rect 352 -3502 353 -3500
rect 352 -3508 353 -3506
rect 359 -3502 360 -3500
rect 359 -3508 360 -3506
rect 366 -3502 367 -3500
rect 366 -3508 367 -3506
rect 373 -3502 374 -3500
rect 373 -3508 374 -3506
rect 380 -3502 381 -3500
rect 380 -3508 381 -3506
rect 387 -3508 388 -3506
rect 394 -3502 395 -3500
rect 394 -3508 395 -3506
rect 401 -3508 402 -3506
rect 408 -3502 409 -3500
rect 408 -3508 409 -3506
rect 415 -3502 416 -3500
rect 415 -3508 416 -3506
rect 422 -3502 423 -3500
rect 425 -3502 426 -3500
rect 422 -3508 423 -3506
rect 425 -3508 426 -3506
rect 429 -3502 430 -3500
rect 429 -3508 430 -3506
rect 436 -3502 437 -3500
rect 436 -3508 437 -3506
rect 443 -3502 444 -3500
rect 443 -3508 444 -3506
rect 450 -3502 451 -3500
rect 450 -3508 451 -3506
rect 457 -3502 458 -3500
rect 457 -3508 458 -3506
rect 464 -3502 465 -3500
rect 467 -3502 468 -3500
rect 464 -3508 465 -3506
rect 467 -3508 468 -3506
rect 471 -3502 472 -3500
rect 471 -3508 472 -3506
rect 478 -3502 479 -3500
rect 478 -3508 479 -3506
rect 485 -3502 486 -3500
rect 485 -3508 486 -3506
rect 492 -3502 493 -3500
rect 492 -3508 493 -3506
rect 495 -3508 496 -3506
rect 499 -3502 500 -3500
rect 499 -3508 500 -3506
rect 506 -3502 507 -3500
rect 506 -3508 507 -3506
rect 513 -3502 514 -3500
rect 513 -3508 514 -3506
rect 520 -3502 521 -3500
rect 520 -3508 521 -3506
rect 527 -3502 528 -3500
rect 527 -3508 528 -3506
rect 534 -3502 535 -3500
rect 537 -3502 538 -3500
rect 534 -3508 535 -3506
rect 541 -3502 542 -3500
rect 541 -3508 542 -3506
rect 548 -3502 549 -3500
rect 548 -3508 549 -3506
rect 555 -3502 556 -3500
rect 555 -3508 556 -3506
rect 562 -3502 563 -3500
rect 562 -3508 563 -3506
rect 565 -3508 566 -3506
rect 569 -3502 570 -3500
rect 569 -3508 570 -3506
rect 579 -3502 580 -3500
rect 576 -3508 577 -3506
rect 579 -3508 580 -3506
rect 583 -3502 584 -3500
rect 583 -3508 584 -3506
rect 590 -3502 591 -3500
rect 590 -3508 591 -3506
rect 597 -3502 598 -3500
rect 597 -3508 598 -3506
rect 604 -3502 605 -3500
rect 604 -3508 605 -3506
rect 611 -3502 612 -3500
rect 611 -3508 612 -3506
rect 618 -3502 619 -3500
rect 618 -3508 619 -3506
rect 625 -3502 626 -3500
rect 628 -3502 629 -3500
rect 625 -3508 626 -3506
rect 632 -3502 633 -3500
rect 632 -3508 633 -3506
rect 639 -3502 640 -3500
rect 639 -3508 640 -3506
rect 642 -3508 643 -3506
rect 646 -3502 647 -3500
rect 646 -3508 647 -3506
rect 653 -3502 654 -3500
rect 653 -3508 654 -3506
rect 660 -3502 661 -3500
rect 660 -3508 661 -3506
rect 667 -3502 668 -3500
rect 667 -3508 668 -3506
rect 677 -3502 678 -3500
rect 674 -3508 675 -3506
rect 677 -3508 678 -3506
rect 681 -3502 682 -3500
rect 681 -3508 682 -3506
rect 688 -3502 689 -3500
rect 688 -3508 689 -3506
rect 695 -3502 696 -3500
rect 695 -3508 696 -3506
rect 702 -3502 703 -3500
rect 702 -3508 703 -3506
rect 709 -3502 710 -3500
rect 709 -3508 710 -3506
rect 716 -3502 717 -3500
rect 716 -3508 717 -3506
rect 726 -3502 727 -3500
rect 726 -3508 727 -3506
rect 730 -3502 731 -3500
rect 730 -3508 731 -3506
rect 737 -3502 738 -3500
rect 737 -3508 738 -3506
rect 744 -3502 745 -3500
rect 744 -3508 745 -3506
rect 751 -3502 752 -3500
rect 751 -3508 752 -3506
rect 758 -3508 759 -3506
rect 765 -3502 766 -3500
rect 765 -3508 766 -3506
rect 772 -3502 773 -3500
rect 772 -3508 773 -3506
rect 779 -3502 780 -3500
rect 779 -3508 780 -3506
rect 800 -3502 801 -3500
rect 800 -3508 801 -3506
rect 807 -3502 808 -3500
rect 807 -3508 808 -3506
rect 814 -3502 815 -3500
rect 817 -3502 818 -3500
rect 821 -3502 822 -3500
rect 821 -3508 822 -3506
rect 835 -3502 836 -3500
rect 835 -3508 836 -3506
rect 842 -3502 843 -3500
rect 842 -3508 843 -3506
rect 849 -3502 850 -3500
rect 849 -3508 850 -3506
rect 856 -3502 857 -3500
rect 856 -3508 857 -3506
rect 863 -3502 864 -3500
rect 863 -3508 864 -3506
rect 870 -3502 871 -3500
rect 870 -3508 871 -3506
rect 877 -3502 878 -3500
rect 877 -3508 878 -3506
rect 905 -3502 906 -3500
rect 905 -3508 906 -3506
rect 912 -3502 913 -3500
rect 912 -3508 913 -3506
rect 919 -3502 920 -3500
rect 919 -3508 920 -3506
rect 926 -3502 927 -3500
rect 926 -3508 927 -3506
rect 933 -3502 934 -3500
rect 936 -3502 937 -3500
rect 933 -3508 934 -3506
rect 940 -3502 941 -3500
rect 943 -3502 944 -3500
rect 940 -3508 941 -3506
rect 947 -3502 948 -3500
rect 947 -3508 948 -3506
rect 954 -3502 955 -3500
rect 957 -3502 958 -3500
rect 954 -3508 955 -3506
rect 961 -3502 962 -3500
rect 961 -3508 962 -3506
rect 968 -3502 969 -3500
rect 968 -3508 969 -3506
rect 982 -3502 983 -3500
rect 982 -3508 983 -3506
rect 989 -3502 990 -3500
rect 989 -3508 990 -3506
rect 996 -3502 997 -3500
rect 999 -3502 1000 -3500
rect 996 -3508 997 -3506
rect 1003 -3502 1004 -3500
rect 1003 -3508 1004 -3506
rect 1010 -3502 1011 -3500
rect 1010 -3508 1011 -3506
rect 1052 -3502 1053 -3500
rect 1052 -3508 1053 -3506
rect 1080 -3502 1081 -3500
rect 1080 -3508 1081 -3506
rect 1087 -3502 1088 -3500
rect 1087 -3508 1088 -3506
rect 1108 -3502 1109 -3500
rect 1108 -3508 1109 -3506
rect 1122 -3502 1123 -3500
rect 1122 -3508 1123 -3506
rect 1150 -3502 1151 -3500
rect 1150 -3508 1151 -3506
rect 1171 -3502 1172 -3500
rect 1174 -3502 1175 -3500
rect 1171 -3508 1172 -3506
rect 1178 -3502 1179 -3500
rect 1178 -3508 1179 -3506
rect 1339 -3502 1340 -3500
rect 1342 -3502 1343 -3500
rect 1339 -3508 1340 -3506
rect 1346 -3502 1347 -3500
rect 1346 -3508 1347 -3506
rect 1349 -3508 1350 -3506
rect 1353 -3502 1354 -3500
rect 1353 -3508 1354 -3506
rect 247 -3543 248 -3541
rect 247 -3549 248 -3547
rect 254 -3543 255 -3541
rect 257 -3549 258 -3547
rect 261 -3543 262 -3541
rect 261 -3549 262 -3547
rect 268 -3543 269 -3541
rect 268 -3549 269 -3547
rect 296 -3543 297 -3541
rect 296 -3549 297 -3547
rect 345 -3543 346 -3541
rect 345 -3549 346 -3547
rect 359 -3543 360 -3541
rect 359 -3549 360 -3547
rect 380 -3543 381 -3541
rect 380 -3549 381 -3547
rect 394 -3543 395 -3541
rect 394 -3549 395 -3547
rect 401 -3543 402 -3541
rect 401 -3549 402 -3547
rect 408 -3543 409 -3541
rect 408 -3549 409 -3547
rect 415 -3543 416 -3541
rect 415 -3549 416 -3547
rect 422 -3543 423 -3541
rect 422 -3549 423 -3547
rect 429 -3543 430 -3541
rect 432 -3549 433 -3547
rect 436 -3543 437 -3541
rect 436 -3549 437 -3547
rect 443 -3543 444 -3541
rect 450 -3543 451 -3541
rect 453 -3543 454 -3541
rect 450 -3549 451 -3547
rect 453 -3549 454 -3547
rect 457 -3543 458 -3541
rect 457 -3549 458 -3547
rect 464 -3543 465 -3541
rect 464 -3549 465 -3547
rect 471 -3543 472 -3541
rect 471 -3549 472 -3547
rect 478 -3543 479 -3541
rect 478 -3549 479 -3547
rect 488 -3549 489 -3547
rect 492 -3543 493 -3541
rect 492 -3549 493 -3547
rect 499 -3543 500 -3541
rect 499 -3549 500 -3547
rect 506 -3543 507 -3541
rect 506 -3549 507 -3547
rect 513 -3543 514 -3541
rect 513 -3549 514 -3547
rect 520 -3543 521 -3541
rect 520 -3549 521 -3547
rect 527 -3543 528 -3541
rect 527 -3549 528 -3547
rect 534 -3543 535 -3541
rect 534 -3549 535 -3547
rect 541 -3543 542 -3541
rect 544 -3543 545 -3541
rect 541 -3549 542 -3547
rect 544 -3549 545 -3547
rect 548 -3543 549 -3541
rect 548 -3549 549 -3547
rect 555 -3543 556 -3541
rect 555 -3549 556 -3547
rect 562 -3543 563 -3541
rect 562 -3549 563 -3547
rect 569 -3543 570 -3541
rect 569 -3549 570 -3547
rect 576 -3543 577 -3541
rect 576 -3549 577 -3547
rect 583 -3543 584 -3541
rect 583 -3549 584 -3547
rect 590 -3543 591 -3541
rect 590 -3549 591 -3547
rect 600 -3543 601 -3541
rect 600 -3549 601 -3547
rect 604 -3543 605 -3541
rect 604 -3549 605 -3547
rect 611 -3543 612 -3541
rect 611 -3549 612 -3547
rect 625 -3543 626 -3541
rect 628 -3543 629 -3541
rect 628 -3549 629 -3547
rect 639 -3543 640 -3541
rect 639 -3549 640 -3547
rect 667 -3543 668 -3541
rect 667 -3549 668 -3547
rect 681 -3543 682 -3541
rect 681 -3549 682 -3547
rect 688 -3543 689 -3541
rect 691 -3543 692 -3541
rect 695 -3543 696 -3541
rect 695 -3549 696 -3547
rect 702 -3543 703 -3541
rect 702 -3549 703 -3547
rect 709 -3543 710 -3541
rect 716 -3543 717 -3541
rect 716 -3549 717 -3547
rect 723 -3543 724 -3541
rect 723 -3549 724 -3547
rect 726 -3549 727 -3547
rect 730 -3543 731 -3541
rect 730 -3549 731 -3547
rect 737 -3543 738 -3541
rect 737 -3549 738 -3547
rect 744 -3543 745 -3541
rect 744 -3549 745 -3547
rect 751 -3543 752 -3541
rect 751 -3549 752 -3547
rect 758 -3543 759 -3541
rect 758 -3549 759 -3547
rect 765 -3543 766 -3541
rect 765 -3549 766 -3547
rect 835 -3543 836 -3541
rect 835 -3549 836 -3547
rect 849 -3543 850 -3541
rect 849 -3549 850 -3547
rect 863 -3543 864 -3541
rect 863 -3549 864 -3547
rect 870 -3543 871 -3541
rect 870 -3549 871 -3547
rect 877 -3543 878 -3541
rect 877 -3549 878 -3547
rect 884 -3543 885 -3541
rect 884 -3549 885 -3547
rect 891 -3543 892 -3541
rect 891 -3549 892 -3547
rect 898 -3543 899 -3541
rect 898 -3549 899 -3547
rect 905 -3543 906 -3541
rect 905 -3549 906 -3547
rect 912 -3543 913 -3541
rect 912 -3549 913 -3547
rect 922 -3543 923 -3541
rect 919 -3549 920 -3547
rect 926 -3543 927 -3541
rect 926 -3549 927 -3547
rect 933 -3543 934 -3541
rect 933 -3549 934 -3547
rect 940 -3543 941 -3541
rect 943 -3543 944 -3541
rect 947 -3543 948 -3541
rect 947 -3549 948 -3547
rect 968 -3543 969 -3541
rect 968 -3549 969 -3547
rect 975 -3543 976 -3541
rect 975 -3549 976 -3547
rect 989 -3543 990 -3541
rect 989 -3549 990 -3547
rect 1006 -3543 1007 -3541
rect 1006 -3549 1007 -3547
rect 1010 -3543 1011 -3541
rect 1010 -3549 1011 -3547
rect 1052 -3543 1053 -3541
rect 1052 -3549 1053 -3547
rect 1059 -3543 1060 -3541
rect 1059 -3549 1060 -3547
rect 1080 -3543 1081 -3541
rect 1080 -3549 1081 -3547
rect 1108 -3543 1109 -3541
rect 1108 -3549 1109 -3547
rect 1150 -3543 1151 -3541
rect 1150 -3549 1151 -3547
rect 1160 -3543 1161 -3541
rect 1157 -3549 1158 -3547
rect 261 -3580 262 -3578
rect 264 -3586 265 -3584
rect 268 -3580 269 -3578
rect 268 -3586 269 -3584
rect 310 -3580 311 -3578
rect 310 -3586 311 -3584
rect 327 -3580 328 -3578
rect 324 -3586 325 -3584
rect 327 -3586 328 -3584
rect 352 -3580 353 -3578
rect 352 -3586 353 -3584
rect 359 -3580 360 -3578
rect 359 -3586 360 -3584
rect 366 -3580 367 -3578
rect 366 -3586 367 -3584
rect 376 -3580 377 -3578
rect 376 -3586 377 -3584
rect 394 -3580 395 -3578
rect 394 -3586 395 -3584
rect 401 -3580 402 -3578
rect 404 -3586 405 -3584
rect 408 -3580 409 -3578
rect 408 -3586 409 -3584
rect 415 -3580 416 -3578
rect 415 -3586 416 -3584
rect 436 -3580 437 -3578
rect 436 -3586 437 -3584
rect 443 -3580 444 -3578
rect 443 -3586 444 -3584
rect 446 -3586 447 -3584
rect 450 -3580 451 -3578
rect 450 -3586 451 -3584
rect 457 -3580 458 -3578
rect 457 -3586 458 -3584
rect 464 -3580 465 -3578
rect 464 -3586 465 -3584
rect 471 -3580 472 -3578
rect 471 -3586 472 -3584
rect 478 -3580 479 -3578
rect 478 -3586 479 -3584
rect 485 -3580 486 -3578
rect 488 -3580 489 -3578
rect 492 -3580 493 -3578
rect 492 -3586 493 -3584
rect 499 -3580 500 -3578
rect 499 -3586 500 -3584
rect 506 -3580 507 -3578
rect 506 -3586 507 -3584
rect 513 -3580 514 -3578
rect 516 -3586 517 -3584
rect 520 -3580 521 -3578
rect 520 -3586 521 -3584
rect 527 -3580 528 -3578
rect 527 -3586 528 -3584
rect 534 -3580 535 -3578
rect 534 -3586 535 -3584
rect 541 -3580 542 -3578
rect 541 -3586 542 -3584
rect 548 -3580 549 -3578
rect 548 -3586 549 -3584
rect 555 -3580 556 -3578
rect 555 -3586 556 -3584
rect 562 -3580 563 -3578
rect 562 -3586 563 -3584
rect 569 -3580 570 -3578
rect 569 -3586 570 -3584
rect 597 -3580 598 -3578
rect 597 -3586 598 -3584
rect 611 -3580 612 -3578
rect 611 -3586 612 -3584
rect 618 -3580 619 -3578
rect 618 -3586 619 -3584
rect 646 -3580 647 -3578
rect 646 -3586 647 -3584
rect 660 -3580 661 -3578
rect 660 -3586 661 -3584
rect 677 -3580 678 -3578
rect 674 -3586 675 -3584
rect 677 -3586 678 -3584
rect 688 -3580 689 -3578
rect 688 -3586 689 -3584
rect 695 -3580 696 -3578
rect 695 -3586 696 -3584
rect 702 -3580 703 -3578
rect 702 -3586 703 -3584
rect 709 -3586 710 -3584
rect 716 -3580 717 -3578
rect 716 -3586 717 -3584
rect 723 -3580 724 -3578
rect 726 -3580 727 -3578
rect 723 -3586 724 -3584
rect 730 -3580 731 -3578
rect 730 -3586 731 -3584
rect 737 -3580 738 -3578
rect 737 -3586 738 -3584
rect 744 -3580 745 -3578
rect 744 -3586 745 -3584
rect 751 -3580 752 -3578
rect 751 -3586 752 -3584
rect 758 -3580 759 -3578
rect 758 -3586 759 -3584
rect 765 -3580 766 -3578
rect 765 -3586 766 -3584
rect 849 -3580 850 -3578
rect 849 -3586 850 -3584
rect 856 -3580 857 -3578
rect 856 -3586 857 -3584
rect 891 -3580 892 -3578
rect 891 -3586 892 -3584
rect 901 -3580 902 -3578
rect 901 -3586 902 -3584
rect 905 -3580 906 -3578
rect 905 -3586 906 -3584
rect 912 -3580 913 -3578
rect 912 -3586 913 -3584
rect 919 -3580 920 -3578
rect 922 -3580 923 -3578
rect 926 -3580 927 -3578
rect 926 -3586 927 -3584
rect 940 -3580 941 -3578
rect 940 -3586 941 -3584
rect 968 -3580 969 -3578
rect 968 -3586 969 -3584
rect 975 -3580 976 -3578
rect 975 -3586 976 -3584
rect 982 -3580 983 -3578
rect 982 -3586 983 -3584
rect 985 -3586 986 -3584
rect 989 -3580 990 -3578
rect 989 -3586 990 -3584
rect 1038 -3580 1039 -3578
rect 1038 -3586 1039 -3584
rect 1052 -3580 1053 -3578
rect 1052 -3586 1053 -3584
rect 1083 -3586 1084 -3584
rect 1087 -3580 1088 -3578
rect 1087 -3586 1088 -3584
rect 1108 -3580 1109 -3578
rect 1108 -3586 1109 -3584
rect 327 -3603 328 -3601
rect 352 -3603 353 -3601
rect 401 -3603 402 -3601
rect 401 -3609 402 -3607
rect 408 -3603 409 -3601
rect 457 -3603 458 -3601
rect 457 -3609 458 -3607
rect 471 -3603 472 -3601
rect 471 -3609 472 -3607
rect 492 -3603 493 -3601
rect 492 -3609 493 -3607
rect 506 -3603 507 -3601
rect 506 -3609 507 -3607
rect 516 -3603 517 -3601
rect 513 -3609 514 -3607
rect 516 -3609 517 -3607
rect 520 -3603 521 -3601
rect 520 -3609 521 -3607
rect 544 -3603 545 -3601
rect 541 -3609 542 -3607
rect 548 -3603 549 -3601
rect 548 -3609 549 -3607
rect 555 -3603 556 -3601
rect 555 -3609 556 -3607
rect 562 -3603 563 -3601
rect 562 -3609 563 -3607
rect 569 -3603 570 -3601
rect 569 -3609 570 -3607
rect 576 -3603 577 -3601
rect 576 -3609 577 -3607
rect 597 -3603 598 -3601
rect 597 -3609 598 -3607
rect 604 -3603 605 -3601
rect 604 -3609 605 -3607
rect 614 -3603 615 -3601
rect 611 -3609 612 -3607
rect 681 -3603 682 -3601
rect 684 -3609 685 -3607
rect 695 -3603 696 -3601
rect 695 -3609 696 -3607
rect 702 -3603 703 -3601
rect 702 -3609 703 -3607
rect 709 -3603 710 -3601
rect 709 -3609 710 -3607
rect 712 -3609 713 -3607
rect 716 -3603 717 -3601
rect 716 -3609 717 -3607
rect 723 -3603 724 -3601
rect 723 -3609 724 -3607
rect 730 -3603 731 -3601
rect 730 -3609 731 -3607
rect 737 -3603 738 -3601
rect 737 -3609 738 -3607
rect 744 -3603 745 -3601
rect 744 -3609 745 -3607
rect 751 -3603 752 -3601
rect 751 -3609 752 -3607
rect 758 -3603 759 -3601
rect 758 -3609 759 -3607
rect 761 -3609 762 -3607
rect 765 -3603 766 -3601
rect 765 -3609 766 -3607
rect 772 -3603 773 -3601
rect 772 -3609 773 -3607
rect 856 -3603 857 -3601
rect 856 -3609 857 -3607
rect 863 -3603 864 -3601
rect 863 -3609 864 -3607
rect 905 -3603 906 -3601
rect 908 -3603 909 -3601
rect 919 -3603 920 -3601
rect 919 -3609 920 -3607
rect 926 -3603 927 -3601
rect 926 -3609 927 -3607
rect 975 -3603 976 -3601
rect 975 -3609 976 -3607
rect 982 -3603 983 -3601
rect 982 -3609 983 -3607
rect 1031 -3603 1032 -3601
rect 1031 -3609 1032 -3607
rect 1045 -3603 1046 -3601
rect 1045 -3609 1046 -3607
rect 1052 -3603 1053 -3601
rect 1052 -3609 1053 -3607
rect 1108 -3603 1109 -3601
rect 1108 -3609 1109 -3607
rect 401 -3628 402 -3626
rect 401 -3634 402 -3632
rect 408 -3634 409 -3632
rect 464 -3628 465 -3626
rect 464 -3634 465 -3632
rect 471 -3628 472 -3626
rect 471 -3634 472 -3632
rect 527 -3628 528 -3626
rect 527 -3634 528 -3632
rect 562 -3628 563 -3626
rect 562 -3634 563 -3632
rect 569 -3628 570 -3626
rect 569 -3634 570 -3632
rect 576 -3628 577 -3626
rect 576 -3634 577 -3632
rect 583 -3628 584 -3626
rect 583 -3634 584 -3632
rect 590 -3628 591 -3626
rect 590 -3634 591 -3632
rect 702 -3628 703 -3626
rect 702 -3634 703 -3632
rect 709 -3628 710 -3626
rect 712 -3628 713 -3626
rect 709 -3634 710 -3632
rect 716 -3628 717 -3626
rect 716 -3634 717 -3632
rect 723 -3628 724 -3626
rect 723 -3634 724 -3632
rect 744 -3628 745 -3626
rect 744 -3634 745 -3632
rect 751 -3628 752 -3626
rect 751 -3634 752 -3632
rect 758 -3628 759 -3626
rect 758 -3634 759 -3632
rect 765 -3628 766 -3626
rect 765 -3634 766 -3632
rect 775 -3628 776 -3626
rect 772 -3634 773 -3632
rect 800 -3628 801 -3626
rect 800 -3634 801 -3632
rect 856 -3628 857 -3626
rect 856 -3634 857 -3632
rect 863 -3628 864 -3626
rect 863 -3634 864 -3632
rect 926 -3628 927 -3626
rect 926 -3634 927 -3632
rect 933 -3628 934 -3626
rect 933 -3634 934 -3632
rect 982 -3628 983 -3626
rect 982 -3634 983 -3632
rect 1003 -3628 1004 -3626
rect 1003 -3634 1004 -3632
rect 1031 -3628 1032 -3626
rect 1031 -3634 1032 -3632
rect 1052 -3634 1053 -3632
rect 1055 -3634 1056 -3632
rect 1059 -3628 1060 -3626
rect 1059 -3634 1060 -3632
rect 1080 -3628 1081 -3626
rect 1080 -3634 1081 -3632
rect 1108 -3628 1109 -3626
rect 1108 -3634 1109 -3632
rect 401 -3643 402 -3641
rect 401 -3649 402 -3647
rect 408 -3643 409 -3641
rect 408 -3649 409 -3647
rect 464 -3643 465 -3641
rect 464 -3649 465 -3647
rect 474 -3643 475 -3641
rect 474 -3649 475 -3647
rect 527 -3643 528 -3641
rect 527 -3649 528 -3647
rect 572 -3643 573 -3641
rect 569 -3649 570 -3647
rect 576 -3643 577 -3641
rect 576 -3649 577 -3647
rect 583 -3643 584 -3641
rect 583 -3649 584 -3647
rect 586 -3649 587 -3647
rect 590 -3643 591 -3641
rect 590 -3649 591 -3647
rect 597 -3643 598 -3641
rect 597 -3649 598 -3647
rect 709 -3643 710 -3641
rect 709 -3649 710 -3647
rect 716 -3643 717 -3641
rect 719 -3643 720 -3641
rect 716 -3649 717 -3647
rect 719 -3649 720 -3647
rect 723 -3643 724 -3641
rect 723 -3649 724 -3647
rect 751 -3643 752 -3641
rect 751 -3649 752 -3647
rect 758 -3643 759 -3641
rect 758 -3649 759 -3647
rect 765 -3643 766 -3641
rect 765 -3649 766 -3647
rect 859 -3643 860 -3641
rect 856 -3649 857 -3647
rect 863 -3643 864 -3641
rect 863 -3649 864 -3647
rect 926 -3643 927 -3641
rect 929 -3643 930 -3641
rect 929 -3649 930 -3647
rect 933 -3643 934 -3641
rect 933 -3649 934 -3647
rect 985 -3643 986 -3641
rect 985 -3649 986 -3647
rect 989 -3643 990 -3641
rect 989 -3649 990 -3647
rect 1031 -3643 1032 -3641
rect 1034 -3643 1035 -3641
rect 1094 -3643 1095 -3641
rect 1094 -3649 1095 -3647
rect 1111 -3643 1112 -3641
rect 1108 -3649 1109 -3647
rect 401 -3658 402 -3656
rect 404 -3664 405 -3662
rect 408 -3658 409 -3656
rect 408 -3664 409 -3662
rect 527 -3664 528 -3662
rect 534 -3658 535 -3656
rect 534 -3664 535 -3662
rect 758 -3658 759 -3656
rect 758 -3664 759 -3662
rect 765 -3658 766 -3656
rect 765 -3664 766 -3662
rect 768 -3664 769 -3662
rect 772 -3658 773 -3656
rect 772 -3664 773 -3662
<< metal1 >>
rect 226 0 332 1
rect 366 0 405 1
rect 415 0 563 1
rect 590 0 643 1
rect 667 0 675 1
rect 705 0 829 1
rect 254 -2 381 -1
rect 401 -2 451 -1
rect 457 -2 472 -1
rect 492 -2 538 -1
rect 765 -2 801 -1
rect 803 -2 843 -1
rect 275 -4 461 -3
rect 506 -4 514 -3
rect 516 -4 528 -3
rect 534 -4 570 -3
rect 317 -6 374 -5
rect 429 -6 437 -5
rect 135 -17 223 -16
rect 303 -17 318 -16
rect 327 -17 381 -16
rect 383 -17 535 -16
rect 541 -17 549 -16
rect 565 -17 710 -16
rect 775 -17 801 -16
rect 821 -17 920 -16
rect 191 -19 227 -18
rect 310 -19 339 -18
rect 345 -19 367 -18
rect 373 -19 444 -18
rect 450 -19 521 -18
rect 527 -19 542 -18
rect 569 -19 584 -18
rect 632 -19 668 -18
rect 674 -19 696 -18
rect 782 -19 794 -18
rect 828 -19 878 -18
rect 205 -21 255 -20
rect 331 -21 479 -20
rect 488 -21 556 -20
rect 569 -21 706 -20
rect 842 -21 857 -20
rect 212 -23 276 -22
rect 331 -23 405 -22
rect 408 -23 465 -22
rect 506 -23 514 -22
rect 576 -23 591 -22
rect 635 -23 654 -22
rect 660 -23 762 -22
rect 226 -25 297 -24
rect 352 -25 416 -24
rect 436 -25 447 -24
rect 450 -25 528 -24
rect 639 -25 703 -24
rect 254 -27 367 -26
rect 376 -27 423 -26
rect 443 -27 685 -26
rect 299 -29 416 -28
rect 457 -29 647 -28
rect 317 -31 447 -30
rect 618 -31 640 -30
rect 387 -33 395 -32
rect 401 -33 458 -32
rect 618 -33 787 -32
rect 359 -35 395 -34
rect 79 -46 237 -45
rect 268 -46 332 -45
rect 380 -46 447 -45
rect 450 -46 605 -45
rect 618 -46 808 -45
rect 856 -46 864 -45
rect 877 -46 906 -45
rect 919 -46 969 -45
rect 100 -48 136 -47
rect 142 -48 328 -47
rect 380 -48 573 -47
rect 576 -48 598 -47
rect 632 -48 654 -47
rect 667 -48 724 -47
rect 758 -48 871 -47
rect 128 -50 237 -49
rect 278 -50 304 -49
rect 324 -50 475 -49
rect 478 -50 612 -49
rect 639 -50 689 -49
rect 695 -50 752 -49
rect 761 -50 892 -49
rect 149 -52 318 -51
rect 397 -52 402 -51
rect 408 -52 507 -51
rect 541 -52 563 -51
rect 576 -52 584 -51
rect 590 -52 654 -51
rect 660 -52 668 -51
rect 702 -52 745 -51
rect 765 -52 773 -51
rect 786 -52 857 -51
rect 156 -54 255 -53
rect 289 -54 367 -53
rect 422 -54 468 -53
rect 485 -54 643 -53
rect 702 -54 825 -53
rect 163 -56 181 -55
rect 184 -56 192 -55
rect 219 -56 454 -55
rect 464 -56 696 -55
rect 709 -56 787 -55
rect 793 -56 815 -55
rect 170 -58 297 -57
rect 303 -58 360 -57
rect 366 -58 479 -57
rect 499 -58 570 -57
rect 625 -58 766 -57
rect 800 -58 822 -57
rect 177 -60 199 -59
rect 222 -60 360 -59
rect 415 -60 423 -59
rect 436 -60 472 -59
rect 520 -60 710 -59
rect 177 -62 465 -61
rect 527 -62 542 -61
rect 555 -62 717 -61
rect 180 -64 206 -63
rect 226 -64 255 -63
rect 261 -64 297 -63
rect 317 -64 353 -63
rect 369 -64 521 -63
rect 527 -64 741 -63
rect 191 -66 213 -65
rect 226 -66 584 -65
rect 646 -66 801 -65
rect 205 -68 374 -67
rect 415 -68 458 -67
rect 534 -68 661 -67
rect 681 -68 794 -67
rect 229 -70 430 -69
rect 450 -70 489 -69
rect 513 -70 535 -69
rect 548 -70 556 -69
rect 569 -70 619 -69
rect 646 -70 783 -69
rect 243 -72 353 -71
rect 369 -72 780 -71
rect 331 -74 682 -73
rect 338 -76 409 -75
rect 457 -76 629 -75
rect 338 -78 622 -77
rect 373 -80 388 -79
rect 492 -80 514 -79
rect 548 -80 594 -79
rect 492 -82 734 -81
rect 593 -84 675 -83
rect 79 -95 391 -94
rect 418 -95 759 -94
rect 814 -95 850 -94
rect 856 -95 920 -94
rect 940 -95 976 -94
rect 114 -97 339 -96
rect 352 -97 395 -96
rect 432 -97 710 -96
rect 730 -97 773 -96
rect 842 -97 948 -96
rect 968 -97 1004 -96
rect 100 -99 115 -98
rect 128 -99 227 -98
rect 250 -99 731 -98
rect 744 -99 836 -98
rect 870 -99 955 -98
rect 100 -101 118 -100
rect 149 -101 335 -100
rect 352 -101 416 -100
rect 443 -101 710 -100
rect 744 -101 787 -100
rect 863 -101 871 -100
rect 891 -101 962 -100
rect 156 -103 237 -102
rect 240 -103 444 -102
rect 446 -103 549 -102
rect 558 -103 969 -102
rect 205 -105 339 -104
rect 453 -105 717 -104
rect 723 -105 864 -104
rect 905 -105 927 -104
rect 205 -107 276 -106
rect 282 -107 311 -106
rect 324 -107 328 -106
rect 506 -107 780 -106
rect 793 -107 906 -106
rect 149 -109 276 -108
rect 292 -109 409 -108
rect 499 -109 507 -108
rect 513 -109 626 -108
rect 642 -109 829 -108
rect 145 -111 409 -110
rect 513 -111 685 -110
rect 688 -111 815 -110
rect 821 -111 892 -110
rect 170 -113 283 -112
rect 296 -113 416 -112
rect 562 -113 640 -112
rect 646 -113 650 -112
rect 660 -113 983 -112
rect 170 -115 468 -114
rect 485 -115 563 -114
rect 569 -115 934 -114
rect 215 -117 227 -116
rect 268 -117 300 -116
rect 303 -117 367 -116
rect 569 -117 633 -116
rect 646 -117 654 -116
rect 660 -117 741 -116
rect 751 -117 899 -116
rect 177 -119 300 -118
rect 310 -119 318 -118
rect 324 -119 381 -118
rect 471 -119 633 -118
rect 653 -119 808 -118
rect 177 -121 262 -120
rect 268 -121 304 -120
rect 359 -121 500 -120
rect 548 -121 752 -120
rect 754 -121 822 -120
rect 191 -123 262 -122
rect 278 -123 297 -122
rect 345 -123 360 -122
rect 471 -123 612 -122
rect 618 -123 885 -122
rect 142 -125 346 -124
rect 450 -125 619 -124
rect 649 -125 808 -124
rect 184 -127 192 -126
rect 212 -127 367 -126
rect 436 -127 451 -126
rect 534 -127 612 -126
rect 667 -127 990 -126
rect 184 -129 475 -128
rect 555 -129 668 -128
rect 674 -129 773 -128
rect 198 -131 213 -130
rect 254 -131 318 -130
rect 457 -131 535 -130
rect 583 -131 878 -130
rect 198 -133 220 -132
rect 240 -133 255 -132
rect 285 -133 437 -132
rect 457 -133 510 -132
rect 583 -133 605 -132
rect 674 -133 762 -132
rect 765 -133 787 -132
rect 219 -135 272 -134
rect 285 -135 332 -134
rect 492 -135 605 -134
rect 688 -135 703 -134
rect 716 -135 801 -134
rect 422 -137 493 -136
rect 520 -137 801 -136
rect 401 -139 423 -138
rect 520 -139 528 -138
rect 590 -139 682 -138
rect 695 -139 913 -138
rect 373 -141 402 -140
rect 429 -141 528 -140
rect 597 -141 724 -140
rect 289 -143 374 -142
rect 429 -143 794 -142
rect 233 -145 290 -144
rect 478 -145 591 -144
rect 681 -145 766 -144
rect 478 -147 577 -146
rect 702 -147 738 -146
rect 464 -149 577 -148
rect 464 -151 857 -150
rect 541 -153 598 -152
rect 488 -155 542 -154
rect 72 -166 433 -165
rect 450 -166 482 -165
rect 495 -166 591 -165
rect 618 -166 864 -165
rect 870 -166 941 -165
rect 954 -166 1088 -165
rect 100 -168 129 -167
rect 135 -168 353 -167
rect 390 -168 437 -167
rect 453 -168 528 -167
rect 541 -168 556 -167
rect 618 -168 717 -167
rect 730 -168 1123 -167
rect 100 -170 115 -169
rect 124 -170 1053 -169
rect 107 -172 871 -171
rect 877 -172 1032 -171
rect 110 -174 419 -173
rect 457 -174 591 -173
rect 621 -174 1130 -173
rect 114 -176 493 -175
rect 509 -176 1081 -175
rect 149 -178 248 -177
rect 254 -178 430 -177
rect 467 -178 675 -177
rect 695 -178 713 -177
rect 730 -178 983 -177
rect 1003 -178 1060 -177
rect 156 -180 493 -179
rect 506 -180 675 -179
rect 695 -180 990 -179
rect 996 -180 1004 -179
rect 170 -182 290 -181
rect 310 -182 342 -181
rect 352 -182 489 -181
rect 506 -182 521 -181
rect 632 -182 717 -181
rect 786 -182 864 -181
rect 884 -182 1074 -181
rect 166 -184 521 -183
rect 562 -184 633 -183
rect 667 -184 671 -183
rect 828 -184 1046 -183
rect 173 -186 293 -185
rect 310 -186 475 -185
rect 488 -186 699 -185
rect 835 -186 885 -185
rect 891 -186 1018 -185
rect 184 -188 451 -187
rect 471 -188 542 -187
rect 562 -188 703 -187
rect 814 -188 892 -187
rect 898 -188 1067 -187
rect 163 -190 185 -189
rect 208 -190 213 -189
rect 219 -190 248 -189
rect 261 -190 437 -189
rect 639 -190 703 -189
rect 814 -190 829 -189
rect 856 -190 983 -189
rect 163 -192 836 -191
rect 905 -192 990 -191
rect 177 -194 640 -193
rect 667 -194 745 -193
rect 758 -194 857 -193
rect 912 -194 1109 -193
rect 177 -196 304 -195
rect 324 -196 458 -195
rect 653 -196 759 -195
rect 779 -196 913 -195
rect 919 -196 1025 -195
rect 121 -198 325 -197
rect 380 -198 528 -197
rect 597 -198 654 -197
rect 688 -198 745 -197
rect 793 -198 906 -197
rect 926 -198 1011 -197
rect 212 -200 367 -199
rect 380 -200 423 -199
rect 432 -200 598 -199
rect 712 -200 794 -199
rect 821 -200 899 -199
rect 933 -200 1095 -199
rect 219 -202 269 -201
rect 282 -202 374 -201
rect 394 -202 465 -201
rect 737 -202 780 -201
rect 842 -202 927 -201
rect 943 -202 955 -201
rect 961 -202 1039 -201
rect 222 -204 304 -203
rect 331 -204 423 -203
rect 464 -204 479 -203
rect 611 -204 738 -203
rect 754 -204 934 -203
rect 947 -204 997 -203
rect 226 -206 276 -205
rect 285 -206 559 -205
rect 681 -206 962 -205
rect 968 -206 1116 -205
rect 226 -208 549 -207
rect 681 -208 948 -207
rect 975 -208 1000 -207
rect 240 -210 276 -209
rect 289 -210 612 -209
rect 705 -210 969 -209
rect 250 -212 283 -211
rect 317 -212 976 -211
rect 261 -214 430 -213
rect 478 -214 878 -213
rect 271 -216 332 -215
rect 359 -216 374 -215
rect 394 -216 409 -215
rect 415 -216 514 -215
rect 548 -216 584 -215
rect 772 -216 822 -215
rect 849 -216 920 -215
rect 205 -218 360 -217
rect 366 -218 685 -217
rect 723 -218 773 -217
rect 205 -220 486 -219
rect 513 -220 661 -219
rect 765 -220 850 -219
rect 257 -222 409 -221
rect 604 -222 661 -221
rect 765 -222 787 -221
rect 345 -224 584 -223
rect 646 -224 724 -223
rect 278 -226 346 -225
rect 401 -226 405 -225
rect 569 -226 605 -225
rect 401 -228 752 -227
rect 534 -230 570 -229
rect 576 -230 647 -229
rect 233 -232 577 -231
rect 191 -234 234 -233
rect 534 -234 808 -233
rect 191 -236 447 -235
rect 800 -236 808 -235
rect 709 -238 801 -237
rect 387 -240 710 -239
rect 387 -242 500 -241
rect 443 -244 500 -243
rect 296 -246 444 -245
rect 296 -248 339 -247
rect 338 -250 1102 -249
rect 54 -261 283 -260
rect 296 -261 444 -260
rect 481 -261 577 -260
rect 614 -261 1032 -260
rect 1038 -261 1207 -260
rect 72 -263 122 -262
rect 124 -263 209 -262
rect 219 -263 913 -262
rect 947 -263 1032 -262
rect 1052 -263 1263 -262
rect 79 -265 1186 -264
rect 86 -267 101 -266
rect 110 -267 339 -266
rect 345 -267 430 -266
rect 481 -267 857 -266
rect 898 -267 948 -266
rect 954 -267 1137 -266
rect 93 -269 580 -268
rect 635 -269 1179 -268
rect 100 -271 374 -270
rect 401 -271 472 -270
rect 485 -271 507 -270
rect 516 -271 717 -270
rect 726 -271 1144 -270
rect 124 -273 1053 -272
rect 1059 -273 1228 -272
rect 128 -275 132 -274
rect 142 -275 192 -274
rect 219 -275 605 -274
rect 663 -275 1067 -274
rect 1073 -275 1242 -274
rect 128 -277 206 -276
rect 240 -277 262 -276
rect 289 -277 346 -276
rect 359 -277 402 -276
rect 457 -277 507 -276
rect 530 -277 843 -276
rect 849 -277 899 -276
rect 954 -277 1130 -276
rect 149 -279 234 -278
rect 254 -279 584 -278
rect 604 -279 1046 -278
rect 1080 -279 1270 -278
rect 156 -281 339 -280
rect 488 -281 1039 -280
rect 1087 -281 1291 -280
rect 163 -283 437 -282
rect 467 -283 1088 -282
rect 1094 -283 1284 -282
rect 82 -285 437 -284
rect 492 -285 738 -284
rect 744 -285 857 -284
rect 877 -285 1067 -284
rect 163 -287 416 -286
rect 541 -287 731 -286
rect 765 -287 1277 -286
rect 184 -289 192 -288
rect 198 -289 206 -288
rect 212 -289 458 -288
rect 513 -289 542 -288
rect 544 -289 1151 -288
rect 58 -291 213 -290
rect 254 -291 388 -290
rect 408 -291 731 -290
rect 768 -291 906 -290
rect 933 -291 1081 -290
rect 107 -293 185 -292
rect 268 -293 290 -292
rect 296 -293 318 -292
rect 320 -293 640 -292
rect 646 -293 766 -292
rect 779 -293 878 -292
rect 884 -293 1095 -292
rect 107 -295 276 -294
rect 303 -295 374 -294
rect 387 -295 535 -294
rect 548 -295 594 -294
rect 597 -295 745 -294
rect 751 -295 885 -294
rect 891 -295 1046 -294
rect 114 -297 549 -296
rect 562 -297 598 -296
rect 625 -297 647 -296
rect 702 -297 829 -296
rect 831 -297 997 -296
rect 1003 -297 1172 -296
rect 135 -299 199 -298
rect 247 -299 269 -298
rect 275 -299 423 -298
rect 471 -299 780 -298
rect 786 -299 1060 -298
rect 131 -301 136 -300
rect 177 -301 409 -300
rect 415 -301 563 -300
rect 569 -301 626 -300
rect 632 -301 738 -300
rect 772 -301 892 -300
rect 940 -301 997 -300
rect 1010 -301 1200 -300
rect 177 -303 496 -302
rect 499 -303 535 -302
rect 569 -303 801 -302
rect 807 -303 1074 -302
rect 236 -305 941 -304
rect 968 -305 1158 -304
rect 303 -307 479 -306
rect 513 -307 1011 -306
rect 1017 -307 1235 -306
rect 114 -309 479 -308
rect 520 -309 752 -308
rect 793 -309 913 -308
rect 968 -309 1123 -308
rect 317 -311 353 -310
rect 366 -311 423 -310
rect 464 -311 500 -310
rect 520 -311 528 -310
rect 576 -311 794 -310
rect 814 -311 906 -310
rect 961 -311 1123 -310
rect 310 -313 353 -312
rect 404 -313 962 -312
rect 975 -313 1165 -312
rect 310 -315 325 -314
rect 485 -315 815 -314
rect 821 -315 850 -314
rect 863 -315 934 -314
rect 982 -315 1193 -314
rect 324 -317 332 -316
rect 527 -317 1221 -316
rect 583 -319 1102 -318
rect 632 -321 1109 -320
rect 586 -323 1109 -322
rect 586 -325 976 -324
rect 989 -325 1256 -324
rect 639 -327 668 -326
rect 674 -327 822 -326
rect 835 -327 1130 -326
rect 607 -329 836 -328
rect 842 -329 1116 -328
rect 611 -331 675 -330
rect 684 -331 808 -330
rect 870 -331 1004 -330
rect 1024 -331 1249 -330
rect 72 -333 612 -332
rect 618 -333 668 -332
rect 688 -333 871 -332
rect 919 -333 1116 -332
rect 450 -335 619 -334
rect 653 -335 689 -334
rect 695 -335 864 -334
rect 926 -335 1102 -334
rect 226 -337 696 -336
rect 709 -337 1018 -336
rect 226 -339 342 -338
rect 446 -339 451 -338
rect 488 -339 920 -338
rect 555 -341 654 -340
rect 660 -341 703 -340
rect 719 -341 983 -340
rect 394 -343 556 -342
rect 590 -343 710 -342
rect 723 -343 801 -342
rect 845 -343 1025 -342
rect 173 -345 395 -344
rect 590 -345 1214 -344
rect 758 -347 990 -346
rect 380 -349 759 -348
rect 786 -349 927 -348
rect 170 -351 381 -350
rect 51 -353 171 -352
rect 58 -364 1060 -363
rect 1227 -364 1312 -363
rect 1332 -364 1375 -363
rect 65 -366 339 -365
rect 366 -366 542 -365
rect 558 -366 892 -365
rect 919 -366 1319 -365
rect 79 -368 83 -367
rect 96 -368 976 -367
rect 1038 -368 1298 -367
rect 1300 -368 1305 -367
rect 114 -370 475 -369
rect 485 -370 759 -369
rect 786 -370 1172 -369
rect 1234 -370 1326 -369
rect 124 -372 129 -371
rect 149 -372 160 -371
rect 163 -372 262 -371
rect 296 -372 517 -371
rect 530 -372 864 -371
rect 891 -372 955 -371
rect 996 -372 1172 -371
rect 1248 -372 1340 -371
rect 128 -374 304 -373
rect 310 -374 538 -373
rect 565 -374 1144 -373
rect 1157 -374 1249 -373
rect 1255 -374 1347 -373
rect 152 -376 174 -375
rect 184 -376 360 -375
rect 380 -376 465 -375
rect 488 -376 1088 -375
rect 1136 -376 1235 -375
rect 1262 -376 1354 -375
rect 163 -378 626 -377
rect 677 -378 1074 -377
rect 1087 -378 1214 -377
rect 1276 -378 1361 -377
rect 170 -380 1242 -379
rect 1290 -380 1368 -379
rect 170 -382 192 -381
rect 198 -382 486 -381
rect 513 -382 794 -381
rect 800 -382 804 -381
rect 831 -382 1004 -381
rect 1024 -382 1074 -381
rect 1115 -382 1214 -381
rect 184 -384 227 -383
rect 247 -384 503 -383
rect 516 -384 1228 -383
rect 191 -386 563 -385
rect 579 -386 1284 -385
rect 198 -388 206 -387
rect 219 -388 493 -387
rect 534 -388 542 -387
rect 562 -388 598 -387
rect 604 -388 724 -387
rect 726 -388 1123 -387
rect 1150 -388 1242 -387
rect 124 -390 605 -389
rect 607 -390 1060 -389
rect 1066 -390 1137 -389
rect 1164 -390 1263 -389
rect 135 -392 206 -391
rect 219 -392 636 -391
rect 684 -392 1081 -391
rect 1122 -392 1179 -391
rect 1185 -392 1277 -391
rect 135 -394 731 -393
rect 754 -394 1221 -393
rect 226 -396 409 -395
rect 457 -396 615 -395
rect 632 -396 794 -395
rect 800 -396 843 -395
rect 849 -396 1067 -395
rect 1094 -396 1186 -395
rect 1192 -396 1284 -395
rect 296 -398 514 -397
rect 576 -398 1165 -397
rect 1206 -398 1291 -397
rect 303 -400 346 -399
rect 373 -400 409 -399
rect 481 -400 1081 -399
rect 1101 -400 1193 -399
rect 310 -402 664 -401
rect 716 -402 864 -401
rect 898 -402 1256 -401
rect 324 -404 479 -403
rect 576 -404 815 -403
rect 828 -404 899 -403
rect 905 -404 1151 -403
rect 107 -406 479 -405
rect 579 -406 1207 -405
rect 107 -408 234 -407
rect 289 -408 325 -407
rect 331 -408 528 -407
rect 583 -408 776 -407
rect 803 -408 843 -407
rect 849 -408 990 -407
rect 1031 -408 1039 -407
rect 1052 -408 1095 -407
rect 1101 -408 1200 -407
rect 177 -410 528 -409
rect 583 -410 717 -409
rect 719 -410 955 -409
rect 968 -410 1004 -409
rect 1010 -410 1053 -409
rect 1108 -410 1200 -409
rect 156 -412 1109 -411
rect 131 -414 157 -413
rect 177 -414 468 -413
rect 586 -414 885 -413
rect 912 -414 1144 -413
rect 233 -416 710 -415
rect 723 -416 885 -415
rect 926 -416 990 -415
rect 338 -418 458 -417
rect 520 -418 913 -417
rect 940 -418 997 -417
rect 345 -420 444 -419
rect 506 -420 521 -419
rect 597 -420 1046 -419
rect 149 -422 1046 -421
rect 373 -424 682 -423
rect 702 -424 815 -423
rect 835 -424 906 -423
rect 982 -424 1025 -423
rect 380 -426 437 -425
rect 611 -426 626 -425
rect 632 -426 1018 -425
rect 387 -428 507 -427
rect 635 -428 1270 -427
rect 352 -430 388 -429
rect 394 -430 573 -429
rect 642 -430 1011 -429
rect 72 -432 395 -431
rect 401 -432 976 -431
rect 72 -434 87 -433
rect 100 -434 353 -433
rect 401 -434 500 -433
rect 660 -434 1179 -433
rect 86 -436 213 -435
rect 422 -436 437 -435
rect 499 -436 556 -435
rect 660 -436 675 -435
rect 684 -436 1270 -435
rect 100 -438 276 -437
rect 415 -438 423 -437
rect 429 -438 444 -437
rect 555 -438 1116 -437
rect 212 -440 962 -439
rect 254 -442 430 -441
rect 667 -442 710 -441
rect 730 -442 766 -441
rect 772 -442 941 -441
rect 947 -442 962 -441
rect 254 -444 472 -443
rect 534 -444 948 -443
rect 317 -446 416 -445
rect 667 -446 822 -445
rect 870 -446 927 -445
rect 933 -446 983 -445
rect 268 -448 318 -447
rect 355 -448 472 -447
rect 590 -448 871 -447
rect 877 -448 934 -447
rect 93 -450 269 -449
rect 590 -450 654 -449
rect 688 -450 878 -449
rect 887 -450 1018 -449
rect 51 -452 689 -451
rect 702 -452 738 -451
rect 744 -452 766 -451
rect 789 -452 836 -451
rect 569 -454 654 -453
rect 674 -454 738 -453
rect 751 -454 1032 -453
rect 142 -456 570 -455
rect 695 -456 745 -455
rect 758 -456 969 -455
rect 142 -458 216 -457
rect 695 -458 1158 -457
rect 789 -460 920 -459
rect 807 -462 1221 -461
rect 779 -464 808 -463
rect 821 -464 857 -463
rect 639 -466 780 -465
rect 639 -468 1130 -467
rect 611 -470 1130 -469
rect 646 -472 857 -471
rect 618 -474 647 -473
rect 450 -476 619 -475
rect 450 -478 461 -477
rect 58 -489 591 -488
rect 611 -489 1298 -488
rect 1377 -489 1382 -488
rect 65 -491 276 -490
rect 310 -491 356 -490
rect 373 -491 601 -490
rect 625 -491 696 -490
rect 698 -491 1319 -490
rect 51 -493 66 -492
rect 68 -493 206 -492
rect 212 -493 220 -492
rect 233 -493 762 -492
rect 768 -493 1326 -492
rect 72 -495 97 -494
rect 114 -495 129 -494
rect 131 -495 283 -494
rect 338 -495 790 -494
rect 831 -495 1284 -494
rect 1325 -495 1354 -494
rect 72 -497 80 -496
rect 124 -497 507 -496
rect 513 -497 976 -496
rect 978 -497 1284 -496
rect 128 -499 248 -498
rect 254 -499 545 -498
rect 569 -499 811 -498
rect 884 -499 1368 -498
rect 152 -501 171 -500
rect 177 -501 339 -500
rect 373 -501 776 -500
rect 782 -501 1144 -500
rect 152 -503 185 -502
rect 198 -503 206 -502
rect 215 -503 913 -502
rect 954 -503 1144 -502
rect 156 -505 580 -504
rect 586 -505 878 -504
rect 887 -505 1389 -504
rect 163 -507 626 -506
rect 646 -507 671 -506
rect 688 -507 885 -506
rect 891 -507 1375 -506
rect 163 -509 409 -508
rect 460 -509 857 -508
rect 870 -509 1368 -508
rect 156 -511 871 -510
rect 912 -511 927 -510
rect 968 -511 1319 -510
rect 177 -513 640 -512
rect 688 -513 780 -512
rect 786 -513 1214 -512
rect 184 -515 654 -514
rect 705 -515 1032 -514
rect 1045 -515 1473 -514
rect 219 -517 479 -516
rect 499 -517 990 -516
rect 1045 -517 1354 -516
rect 222 -519 969 -518
rect 989 -519 1004 -518
rect 1087 -519 1298 -518
rect 240 -521 290 -520
rect 296 -521 647 -520
rect 653 -521 738 -520
rect 754 -521 1060 -520
rect 1178 -521 1214 -520
rect 243 -523 612 -522
rect 614 -523 1060 -522
rect 1178 -523 1235 -522
rect 268 -525 311 -524
rect 380 -525 507 -524
rect 513 -525 668 -524
rect 716 -525 1256 -524
rect 268 -527 332 -526
rect 359 -527 717 -526
rect 719 -527 1151 -526
rect 1248 -527 1256 -526
rect 107 -529 360 -528
rect 397 -529 682 -528
rect 737 -529 745 -528
rect 751 -529 1235 -528
rect 1241 -529 1249 -528
rect 107 -531 829 -530
rect 835 -531 878 -530
rect 901 -531 1032 -530
rect 1150 -531 1165 -530
rect 159 -533 1242 -532
rect 296 -535 402 -534
rect 408 -535 416 -534
rect 499 -535 892 -534
rect 926 -535 1081 -534
rect 1164 -535 1172 -534
rect 317 -537 381 -536
rect 401 -537 633 -536
rect 733 -537 752 -536
rect 772 -537 1018 -536
rect 1073 -537 1081 -536
rect 1171 -537 1186 -536
rect 303 -539 318 -538
rect 324 -539 332 -538
rect 366 -539 745 -538
rect 786 -539 801 -538
rect 814 -539 829 -538
rect 835 -539 843 -538
rect 856 -539 1053 -538
rect 1073 -539 1109 -538
rect 1185 -539 1200 -538
rect 261 -541 304 -540
rect 324 -541 388 -540
rect 415 -541 444 -540
rect 502 -541 794 -540
rect 821 -541 843 -540
rect 919 -541 1018 -540
rect 1108 -541 1193 -540
rect 387 -543 458 -542
rect 502 -543 1277 -542
rect 443 -545 619 -544
rect 674 -545 1053 -544
rect 1101 -545 1193 -544
rect 1276 -545 1305 -544
rect 450 -547 458 -546
rect 492 -547 619 -546
rect 660 -547 675 -546
rect 730 -547 801 -546
rect 807 -547 822 -546
rect 919 -547 997 -546
rect 1003 -547 1025 -546
rect 1094 -547 1102 -546
rect 1115 -547 1200 -546
rect 1304 -547 1312 -546
rect 121 -549 1116 -548
rect 1311 -549 1340 -548
rect 121 -551 531 -550
rect 534 -551 563 -550
rect 590 -551 598 -550
rect 604 -551 955 -550
rect 975 -551 1088 -550
rect 1094 -551 1130 -550
rect 1332 -551 1340 -550
rect 93 -553 1333 -552
rect 142 -555 598 -554
rect 635 -555 1130 -554
rect 135 -557 143 -556
rect 394 -557 535 -556
rect 537 -557 899 -556
rect 940 -557 997 -556
rect 135 -559 1263 -558
rect 149 -561 941 -560
rect 149 -563 696 -562
rect 779 -563 1263 -562
rect 191 -565 395 -564
rect 429 -565 605 -564
rect 639 -565 731 -564
rect 793 -565 1270 -564
rect 191 -567 486 -566
rect 492 -567 584 -566
rect 660 -567 685 -566
rect 1269 -567 1291 -566
rect 345 -569 430 -568
rect 436 -569 451 -568
rect 471 -569 563 -568
rect 583 -569 633 -568
rect 1290 -569 1361 -568
rect 198 -571 1361 -570
rect 250 -573 346 -572
rect 352 -573 685 -572
rect 422 -575 437 -574
rect 464 -575 472 -574
rect 485 -575 703 -574
rect 100 -577 465 -576
rect 478 -577 703 -576
rect 86 -579 101 -578
rect 422 -579 521 -578
rect 527 -579 577 -578
rect 79 -581 87 -580
rect 520 -581 724 -580
rect 527 -583 815 -582
rect 548 -585 570 -584
rect 723 -585 906 -584
rect 226 -587 549 -586
rect 555 -587 899 -586
rect 905 -587 948 -586
rect 40 -589 227 -588
rect 541 -589 556 -588
rect 947 -589 1011 -588
rect 40 -591 262 -590
rect 541 -591 1221 -590
rect 1010 -593 1123 -592
rect 1220 -593 1228 -592
rect 807 -595 1228 -594
rect 961 -597 1123 -596
rect 961 -599 1067 -598
rect 1066 -601 1137 -600
rect 1136 -603 1158 -602
rect 1038 -605 1158 -604
rect 758 -607 1039 -606
rect 758 -609 766 -608
rect 765 -611 1025 -610
rect 44 -622 293 -621
rect 387 -622 584 -621
rect 649 -622 1116 -621
rect 1185 -622 1396 -621
rect 1472 -622 1634 -621
rect 51 -624 517 -623
rect 527 -624 913 -623
rect 975 -624 1046 -623
rect 1059 -624 1186 -623
rect 1234 -624 1501 -623
rect 51 -626 311 -625
rect 397 -626 671 -625
rect 684 -626 1256 -625
rect 1311 -626 1410 -625
rect 72 -628 83 -627
rect 107 -628 559 -627
rect 698 -628 843 -627
rect 887 -628 1102 -627
rect 1136 -628 1235 -627
rect 1353 -628 1382 -627
rect 1388 -628 1571 -627
rect 65 -630 1102 -629
rect 1157 -630 1312 -629
rect 1332 -630 1382 -629
rect 65 -632 227 -631
rect 233 -632 489 -631
rect 537 -632 724 -631
rect 730 -632 1214 -631
rect 1227 -632 1256 -631
rect 1276 -632 1354 -631
rect 1356 -632 1368 -631
rect 72 -634 374 -633
rect 429 -634 503 -633
rect 541 -634 626 -633
rect 702 -634 1375 -633
rect 82 -636 101 -635
rect 114 -636 118 -635
rect 128 -636 227 -635
rect 243 -636 388 -635
rect 432 -636 752 -635
rect 772 -636 1340 -635
rect 1360 -636 1522 -635
rect 86 -638 101 -637
rect 128 -638 556 -637
rect 702 -638 759 -637
rect 768 -638 1361 -637
rect 86 -640 675 -639
rect 705 -640 843 -639
rect 898 -640 1011 -639
rect 1017 -640 1116 -639
rect 1129 -640 1228 -639
rect 1269 -640 1340 -639
rect 138 -642 220 -641
rect 247 -642 857 -641
rect 863 -642 899 -641
rect 940 -642 1011 -641
rect 1080 -642 1137 -641
rect 1157 -642 1165 -641
rect 1171 -642 1277 -641
rect 1290 -642 1389 -641
rect 107 -644 248 -643
rect 250 -644 528 -643
rect 555 -644 766 -643
rect 772 -644 909 -643
rect 954 -644 1046 -643
rect 1052 -644 1165 -643
rect 1192 -644 1333 -643
rect 142 -646 157 -645
rect 159 -646 1403 -645
rect 149 -648 241 -647
rect 250 -648 479 -647
rect 485 -648 594 -647
rect 674 -648 822 -647
rect 831 -648 1179 -647
rect 1206 -648 1270 -647
rect 1290 -648 1305 -647
rect 1325 -648 1375 -647
rect 152 -650 1200 -649
rect 1241 -650 1305 -649
rect 156 -652 797 -651
rect 807 -652 1347 -651
rect 163 -654 430 -653
rect 443 -654 584 -653
rect 586 -654 1200 -653
rect 1248 -654 1347 -653
rect 163 -656 657 -655
rect 695 -656 1130 -655
rect 1248 -656 1427 -655
rect 58 -658 696 -657
rect 709 -658 759 -657
rect 775 -658 979 -657
rect 982 -658 1053 -657
rect 1122 -658 1207 -657
rect 58 -660 94 -659
rect 170 -660 381 -659
rect 415 -660 444 -659
rect 471 -660 479 -659
rect 565 -660 1193 -659
rect 187 -662 206 -661
rect 219 -662 325 -661
rect 345 -662 626 -661
rect 716 -662 1326 -661
rect 124 -664 346 -663
rect 373 -664 465 -663
rect 471 -664 591 -663
rect 607 -664 1242 -663
rect 149 -666 591 -665
rect 716 -666 829 -665
rect 856 -666 1368 -665
rect 201 -668 213 -667
rect 268 -668 367 -667
rect 380 -668 493 -667
rect 719 -668 1095 -667
rect 205 -670 633 -669
rect 723 -670 1298 -669
rect 212 -672 353 -671
rect 401 -672 416 -671
rect 464 -672 713 -671
rect 726 -672 1018 -671
rect 1024 -672 1123 -671
rect 268 -674 531 -673
rect 733 -674 955 -673
rect 961 -674 1179 -673
rect 275 -676 752 -675
rect 779 -676 997 -675
rect 1003 -676 1214 -675
rect 254 -678 276 -677
rect 282 -678 440 -677
rect 611 -678 997 -677
rect 1006 -678 1144 -677
rect 282 -680 580 -679
rect 737 -680 766 -679
rect 786 -680 864 -679
rect 877 -680 962 -679
rect 968 -680 1081 -679
rect 121 -682 738 -681
rect 744 -682 780 -681
rect 793 -682 1417 -681
rect 121 -684 1074 -683
rect 296 -686 542 -685
rect 646 -686 787 -685
rect 793 -686 1319 -685
rect 289 -688 297 -687
rect 310 -688 892 -687
rect 905 -688 1025 -687
rect 1031 -688 1144 -687
rect 1262 -688 1319 -687
rect 317 -690 325 -689
rect 352 -690 605 -689
rect 618 -690 647 -689
rect 733 -690 1074 -689
rect 1108 -690 1263 -689
rect 317 -692 423 -691
rect 513 -692 745 -691
rect 800 -692 878 -691
rect 884 -692 969 -691
rect 989 -692 1095 -691
rect 401 -694 605 -693
rect 660 -694 801 -693
rect 807 -694 913 -693
rect 933 -694 983 -693
rect 992 -694 1151 -693
rect 408 -696 493 -695
rect 513 -696 535 -695
rect 576 -696 619 -695
rect 660 -696 689 -695
rect 814 -696 892 -695
rect 905 -696 1284 -695
rect 68 -698 689 -697
rect 821 -698 836 -697
rect 884 -698 927 -697
rect 1031 -698 1060 -697
rect 1062 -698 1298 -697
rect 96 -700 815 -699
rect 828 -700 941 -699
rect 1038 -700 1172 -699
rect 1220 -700 1284 -699
rect 135 -702 1039 -701
rect 1066 -702 1109 -701
rect 135 -704 262 -703
rect 359 -704 409 -703
rect 422 -704 437 -703
rect 520 -704 612 -703
rect 667 -704 934 -703
rect 1087 -704 1221 -703
rect 184 -706 262 -705
rect 359 -706 654 -705
rect 667 -706 860 -705
rect 870 -706 927 -705
rect 947 -706 1088 -705
rect 436 -708 1151 -707
rect 520 -710 598 -709
rect 653 -710 682 -709
rect 835 -710 902 -709
rect 919 -710 1067 -709
rect 534 -712 570 -711
rect 849 -712 948 -711
rect 548 -714 570 -713
rect 709 -714 850 -713
rect 919 -714 1431 -713
rect 548 -716 640 -715
rect 394 -718 640 -717
rect 177 -720 395 -719
rect 562 -720 598 -719
rect 177 -722 507 -721
rect 191 -724 507 -723
rect 191 -726 339 -725
rect 303 -728 563 -727
rect 303 -730 577 -729
rect 331 -732 339 -731
rect 184 -734 332 -733
rect 37 -745 59 -744
rect 79 -745 920 -744
rect 922 -745 1403 -744
rect 1416 -745 1609 -744
rect 1633 -745 1697 -744
rect 44 -747 1557 -746
rect 1570 -747 1627 -746
rect 44 -749 451 -748
rect 467 -749 1438 -748
rect 1500 -749 1620 -748
rect 58 -751 150 -750
rect 166 -751 1459 -750
rect 1521 -751 1592 -750
rect 1605 -751 1613 -750
rect 82 -753 605 -752
rect 607 -753 878 -752
rect 884 -753 1522 -752
rect 93 -755 801 -754
rect 821 -755 885 -754
rect 905 -755 1347 -754
rect 1353 -755 1550 -754
rect 93 -757 528 -756
rect 537 -757 724 -756
rect 730 -757 780 -756
rect 782 -757 1221 -756
rect 1241 -757 1417 -756
rect 1430 -757 1634 -756
rect 33 -759 528 -758
rect 558 -759 1508 -758
rect 103 -761 367 -760
rect 485 -761 563 -760
rect 565 -761 1095 -760
rect 1122 -761 1543 -760
rect 124 -763 1571 -762
rect 128 -765 132 -764
rect 138 -765 1361 -764
rect 1367 -765 1578 -764
rect 128 -767 619 -766
rect 632 -767 640 -766
rect 649 -767 1368 -766
rect 1374 -767 1585 -766
rect 142 -769 727 -768
rect 730 -769 759 -768
rect 765 -769 822 -768
rect 828 -769 962 -768
rect 1003 -769 1427 -768
rect 149 -771 626 -770
rect 628 -771 1375 -770
rect 1388 -771 1515 -770
rect 184 -773 1494 -772
rect 184 -775 199 -774
rect 205 -775 451 -774
rect 488 -775 556 -774
rect 576 -775 717 -774
rect 733 -775 1424 -774
rect 187 -777 1214 -776
rect 1227 -777 1389 -776
rect 191 -779 237 -778
rect 240 -779 367 -778
rect 471 -779 556 -778
rect 576 -779 864 -778
rect 870 -779 1445 -778
rect 191 -781 430 -780
rect 471 -781 479 -780
rect 499 -781 598 -780
rect 625 -781 703 -780
rect 709 -781 1277 -780
rect 1283 -781 1473 -780
rect 198 -783 563 -782
rect 579 -783 997 -782
rect 1038 -783 1095 -782
rect 1136 -783 1228 -782
rect 1269 -783 1466 -782
rect 205 -785 241 -784
rect 247 -785 1200 -784
rect 1206 -785 1347 -784
rect 1381 -785 1424 -784
rect 233 -787 997 -786
rect 1080 -787 1123 -786
rect 1157 -787 1354 -786
rect 23 -789 234 -788
rect 250 -789 1487 -788
rect 79 -791 251 -790
rect 275 -791 381 -790
rect 429 -791 493 -790
rect 534 -791 1081 -790
rect 1171 -791 1403 -790
rect 135 -793 535 -792
rect 583 -793 598 -792
rect 642 -793 1207 -792
rect 1248 -793 1270 -792
rect 1290 -793 1480 -792
rect 65 -795 584 -794
rect 590 -795 1564 -794
rect 65 -797 829 -796
rect 842 -797 864 -796
rect 877 -797 1200 -796
rect 1262 -797 1382 -796
rect 170 -799 381 -798
rect 408 -799 493 -798
rect 569 -799 591 -798
rect 593 -799 1137 -798
rect 1185 -799 1263 -798
rect 1304 -799 1501 -798
rect 275 -801 797 -800
rect 814 -801 1221 -800
rect 1318 -801 1431 -800
rect 289 -803 353 -802
rect 359 -803 874 -802
rect 908 -803 1284 -802
rect 1325 -803 1452 -802
rect 163 -805 290 -804
rect 310 -805 759 -804
rect 765 -805 836 -804
rect 842 -805 850 -804
rect 856 -805 1277 -804
rect 1332 -805 1529 -804
rect 261 -807 1326 -806
rect 1339 -807 1536 -806
rect 261 -809 283 -808
rect 310 -809 388 -808
rect 408 -809 458 -808
rect 541 -809 570 -808
rect 586 -809 1319 -808
rect 268 -811 360 -810
rect 387 -811 423 -810
rect 432 -811 857 -810
rect 859 -811 1410 -810
rect 177 -813 423 -812
rect 457 -813 640 -812
rect 646 -813 703 -812
rect 716 -813 794 -812
rect 912 -813 1396 -812
rect 177 -815 213 -814
rect 254 -815 269 -814
rect 282 -815 437 -814
rect 513 -815 542 -814
rect 565 -815 1186 -814
rect 1192 -815 1291 -814
rect 1297 -815 1410 -814
rect 110 -817 1298 -816
rect 156 -819 255 -818
rect 317 -819 440 -818
rect 653 -819 1242 -818
rect 1255 -819 1396 -818
rect 156 -821 293 -820
rect 345 -821 619 -820
rect 656 -821 1179 -820
rect 1234 -821 1340 -820
rect 135 -823 1235 -822
rect 212 -825 220 -824
rect 226 -825 437 -824
rect 660 -825 790 -824
rect 887 -825 1179 -824
rect 121 -827 220 -826
rect 345 -827 549 -826
rect 667 -827 801 -826
rect 912 -827 1165 -826
rect 114 -829 122 -828
rect 131 -829 549 -828
rect 667 -829 692 -828
rect 695 -829 713 -828
rect 740 -829 1361 -828
rect 51 -831 696 -830
rect 751 -831 815 -830
rect 919 -831 1151 -830
rect 100 -833 115 -832
rect 170 -833 661 -832
rect 681 -833 724 -832
rect 772 -833 836 -832
rect 929 -833 1312 -832
rect 51 -835 1312 -834
rect 100 -837 1249 -836
rect 352 -839 465 -838
rect 681 -839 738 -838
rect 744 -839 773 -838
rect 786 -839 850 -838
rect 954 -839 1004 -838
rect 1006 -839 1305 -838
rect 72 -841 745 -840
rect 786 -841 1214 -840
rect 72 -843 332 -842
rect 415 -843 514 -842
rect 688 -843 752 -842
rect 933 -843 955 -842
rect 982 -843 1039 -842
rect 1052 -843 1151 -842
rect 296 -845 332 -844
rect 401 -845 416 -844
rect 688 -845 710 -844
rect 831 -845 1053 -844
rect 1066 -845 1158 -844
rect 324 -847 465 -846
rect 831 -847 1256 -846
rect 324 -849 521 -848
rect 891 -849 934 -848
rect 1017 -849 1067 -848
rect 1101 -849 1193 -848
rect 401 -851 444 -850
rect 506 -851 521 -850
rect 611 -851 892 -850
rect 926 -851 983 -850
rect 989 -851 1102 -850
rect 1108 -851 1333 -850
rect 86 -853 444 -852
rect 611 -853 1144 -852
rect 107 -855 1144 -854
rect 107 -857 871 -856
rect 989 -857 993 -856
rect 1017 -857 1060 -856
rect 1115 -857 1165 -856
rect 373 -859 507 -858
rect 1045 -859 1109 -858
rect 1129 -859 1172 -858
rect 373 -861 395 -860
rect 1010 -861 1046 -860
rect 1073 -861 1116 -860
rect 229 -863 395 -862
rect 968 -863 1011 -862
rect 1024 -863 1074 -862
rect 1087 -863 1130 -862
rect 478 -865 1025 -864
rect 1031 -865 1088 -864
rect 940 -867 969 -866
rect 975 -867 1032 -866
rect 674 -869 941 -868
rect 674 -871 738 -870
rect 898 -871 976 -870
rect 898 -873 906 -872
rect 30 -884 73 -883
rect 89 -884 115 -883
rect 135 -884 283 -883
rect 292 -884 339 -883
rect 450 -884 601 -883
rect 618 -884 738 -883
rect 740 -884 1501 -883
rect 1521 -884 1676 -883
rect 1696 -884 1725 -883
rect 65 -886 654 -885
rect 663 -886 1578 -885
rect 1591 -886 1609 -885
rect 1619 -886 1718 -885
rect 65 -888 402 -887
rect 422 -888 451 -887
rect 457 -888 930 -887
rect 957 -888 1536 -887
rect 1598 -888 1627 -887
rect 1633 -888 1711 -887
rect 72 -890 591 -889
rect 597 -890 612 -889
rect 635 -890 1550 -889
rect 86 -892 1592 -891
rect 103 -894 143 -893
rect 149 -894 738 -893
rect 761 -894 892 -893
rect 905 -894 1529 -893
rect 107 -896 122 -895
rect 135 -896 388 -895
rect 422 -896 759 -895
rect 761 -896 892 -895
rect 898 -896 906 -895
rect 908 -896 1333 -895
rect 1374 -896 1522 -895
rect 110 -898 339 -897
rect 387 -898 815 -897
rect 873 -898 1655 -897
rect 114 -900 416 -899
rect 457 -900 668 -899
rect 691 -900 1158 -899
rect 1206 -900 1501 -899
rect 1514 -900 1697 -899
rect 142 -902 479 -901
rect 499 -902 689 -901
rect 705 -902 1193 -901
rect 1220 -902 1550 -901
rect 149 -904 178 -903
rect 184 -904 209 -903
rect 226 -904 269 -903
rect 296 -904 846 -903
rect 877 -904 1151 -903
rect 1234 -904 1627 -903
rect 128 -906 178 -905
rect 184 -906 251 -905
rect 261 -906 283 -905
rect 303 -906 608 -905
rect 611 -906 962 -905
rect 964 -906 1648 -905
rect 128 -908 794 -907
rect 796 -908 1347 -907
rect 1395 -908 1529 -907
rect 138 -910 269 -909
rect 303 -910 584 -909
rect 586 -910 1543 -909
rect 163 -912 997 -911
rect 1038 -912 1158 -911
rect 1248 -912 1375 -911
rect 1430 -912 1536 -911
rect 163 -914 325 -913
rect 331 -914 402 -913
rect 415 -914 717 -913
rect 768 -914 1634 -913
rect 93 -916 325 -915
rect 373 -916 500 -915
rect 548 -916 668 -915
rect 786 -916 1585 -915
rect 86 -918 94 -917
rect 166 -918 514 -917
rect 548 -918 1683 -917
rect 170 -920 482 -919
rect 513 -920 902 -919
rect 912 -920 927 -919
rect 933 -920 997 -919
rect 1059 -920 1466 -919
rect 1486 -920 1606 -919
rect 170 -922 241 -921
rect 247 -922 290 -921
rect 310 -922 594 -921
rect 646 -922 650 -921
rect 733 -922 1487 -921
rect 1493 -922 1669 -921
rect 191 -924 661 -923
rect 765 -924 787 -923
rect 810 -924 1704 -923
rect 79 -926 192 -925
rect 198 -926 661 -925
rect 765 -926 1326 -925
rect 1339 -926 1466 -925
rect 79 -928 563 -927
rect 576 -928 703 -927
rect 856 -928 913 -927
rect 919 -928 962 -927
rect 968 -928 972 -927
rect 975 -928 1039 -927
rect 1062 -928 1389 -927
rect 1437 -928 1585 -927
rect 124 -930 199 -929
rect 205 -930 622 -929
rect 646 -930 1095 -929
rect 1101 -930 1235 -929
rect 1262 -930 1396 -929
rect 1444 -930 1662 -929
rect 226 -932 580 -931
rect 583 -932 696 -931
rect 772 -932 1389 -931
rect 1458 -932 1620 -931
rect 229 -934 1144 -933
rect 1150 -934 1382 -933
rect 1458 -934 1508 -933
rect 121 -936 1508 -935
rect 233 -938 1571 -937
rect 89 -940 234 -939
rect 236 -940 1641 -939
rect 240 -942 353 -941
rect 373 -942 409 -941
rect 436 -942 1221 -941
rect 1255 -942 1571 -941
rect 261 -944 430 -943
rect 436 -944 724 -943
rect 730 -944 773 -943
rect 856 -944 1515 -943
rect 289 -946 1249 -945
rect 1255 -946 1270 -945
rect 1297 -946 1690 -945
rect 37 -948 1298 -947
rect 1304 -948 1445 -947
rect 313 -950 332 -949
rect 345 -950 563 -949
rect 576 -950 633 -949
rect 709 -950 731 -949
rect 863 -950 927 -949
rect 940 -950 1144 -949
rect 1178 -950 1305 -949
rect 1346 -950 1368 -949
rect 1381 -950 1613 -949
rect 317 -952 468 -951
rect 474 -952 675 -951
rect 800 -952 941 -951
rect 968 -952 1018 -951
rect 1031 -952 1340 -951
rect 1353 -952 1494 -951
rect 345 -954 367 -953
rect 394 -954 409 -953
rect 429 -954 626 -953
rect 632 -954 815 -953
rect 849 -954 864 -953
rect 870 -954 1438 -953
rect 107 -956 850 -955
rect 870 -956 1179 -955
rect 1199 -956 1326 -955
rect 1353 -956 1410 -955
rect 352 -958 381 -957
rect 394 -958 724 -957
rect 800 -958 822 -957
rect 877 -958 1417 -957
rect 366 -960 472 -959
rect 478 -960 556 -959
rect 604 -960 710 -959
rect 751 -960 822 -959
rect 884 -960 888 -959
rect 898 -960 1242 -959
rect 1283 -960 1410 -959
rect 37 -962 472 -961
rect 520 -962 556 -961
rect 604 -962 1578 -961
rect 380 -964 486 -963
rect 492 -964 521 -963
rect 527 -964 752 -963
rect 884 -964 983 -963
rect 1003 -964 1095 -963
rect 1115 -964 1263 -963
rect 1290 -964 1417 -963
rect 44 -966 486 -965
rect 534 -966 920 -965
rect 947 -966 1032 -965
rect 1052 -966 1200 -965
rect 1213 -966 1613 -965
rect 44 -968 55 -967
rect 58 -968 493 -967
rect 537 -968 934 -967
rect 975 -968 1431 -967
rect 54 -970 1557 -969
rect 58 -972 1137 -971
rect 1164 -972 1291 -971
rect 100 -974 1557 -973
rect 23 -976 101 -975
rect 219 -976 948 -975
rect 978 -976 1602 -975
rect 359 -978 528 -977
rect 551 -978 745 -977
rect 880 -978 1116 -977
rect 1129 -978 1270 -977
rect 212 -980 360 -979
rect 443 -980 717 -979
rect 744 -980 993 -979
rect 1003 -980 1109 -979
rect 1122 -980 1130 -979
rect 1164 -980 1172 -979
rect 156 -982 444 -981
rect 467 -982 1242 -981
rect 156 -984 794 -983
rect 835 -984 1123 -983
rect 212 -986 542 -985
rect 614 -986 675 -985
rect 835 -986 843 -985
rect 971 -986 1018 -985
rect 1024 -986 1137 -985
rect 541 -988 598 -987
rect 618 -988 696 -987
rect 796 -988 1025 -987
rect 1045 -988 1172 -987
rect 625 -990 682 -989
rect 842 -990 1333 -989
rect 639 -992 1368 -991
rect 639 -994 881 -993
rect 954 -994 1046 -993
rect 1062 -994 1473 -993
rect 681 -996 1284 -995
rect 789 -998 1473 -997
rect 954 -1000 1564 -999
rect 989 -1002 1053 -1001
rect 1066 -1002 1193 -1001
rect 1451 -1002 1564 -1001
rect 989 -1004 1543 -1003
rect 1010 -1006 1102 -1005
rect 1311 -1006 1452 -1005
rect 534 -1008 1312 -1007
rect 1066 -1010 1403 -1009
rect 1073 -1012 1207 -1011
rect 1402 -1012 1424 -1011
rect 628 -1014 1074 -1013
rect 1080 -1014 1214 -1013
rect 779 -1016 1081 -1015
rect 779 -1018 808 -1017
rect 828 -1018 1424 -1017
rect 807 -1020 1011 -1019
rect 828 -1022 1361 -1021
rect 1360 -1024 1480 -1023
rect 1318 -1026 1480 -1025
rect 1185 -1028 1319 -1027
rect 1185 -1030 1228 -1029
rect 1087 -1032 1228 -1031
rect 201 -1034 1088 -1033
rect 44 -1045 241 -1044
rect 261 -1045 633 -1044
rect 681 -1045 1144 -1044
rect 1710 -1045 1732 -1044
rect 65 -1047 489 -1046
rect 499 -1047 633 -1046
rect 681 -1047 696 -1046
rect 719 -1047 1522 -1046
rect 65 -1049 545 -1048
rect 579 -1049 1368 -1048
rect 86 -1051 941 -1050
rect 957 -1051 1627 -1050
rect 89 -1053 1515 -1052
rect 1626 -1053 1669 -1052
rect 93 -1055 188 -1054
rect 198 -1055 402 -1054
rect 408 -1055 535 -1054
rect 590 -1055 1501 -1054
rect 51 -1057 591 -1056
rect 597 -1057 717 -1056
rect 723 -1057 1550 -1056
rect 51 -1059 556 -1058
rect 600 -1059 1011 -1058
rect 1062 -1059 1522 -1058
rect 93 -1061 444 -1060
rect 450 -1061 500 -1060
rect 513 -1061 556 -1060
rect 569 -1061 601 -1060
rect 614 -1061 920 -1060
rect 940 -1061 1039 -1060
rect 1069 -1061 1697 -1060
rect 54 -1063 444 -1062
rect 450 -1063 521 -1062
rect 527 -1063 717 -1062
rect 726 -1063 731 -1062
rect 751 -1063 808 -1062
rect 810 -1063 1046 -1062
rect 1143 -1063 1235 -1062
rect 1360 -1063 1550 -1062
rect 100 -1065 290 -1064
rect 292 -1065 605 -1064
rect 702 -1065 731 -1064
rect 751 -1065 1382 -1064
rect 1500 -1065 1613 -1064
rect 103 -1067 1389 -1066
rect 1612 -1067 1655 -1066
rect 107 -1069 416 -1068
rect 464 -1069 948 -1068
rect 971 -1069 1049 -1068
rect 1234 -1069 1651 -1068
rect 107 -1071 748 -1070
rect 758 -1071 1228 -1070
rect 1276 -1071 1361 -1070
rect 1367 -1071 1466 -1070
rect 89 -1073 1466 -1072
rect 110 -1075 1480 -1074
rect 121 -1077 1221 -1076
rect 1227 -1077 1291 -1076
rect 1381 -1077 1536 -1076
rect 121 -1079 437 -1078
rect 478 -1079 535 -1078
rect 621 -1079 1277 -1078
rect 1290 -1079 1410 -1078
rect 1479 -1079 1641 -1078
rect 128 -1081 437 -1080
rect 506 -1081 528 -1080
rect 621 -1081 1123 -1080
rect 1388 -1081 1431 -1080
rect 1640 -1081 1676 -1080
rect 128 -1083 745 -1082
rect 768 -1083 1340 -1082
rect 1402 -1083 1655 -1082
rect 135 -1085 468 -1084
rect 506 -1085 1242 -1084
rect 1255 -1085 1431 -1084
rect 1619 -1085 1676 -1084
rect 135 -1087 206 -1086
rect 208 -1087 1312 -1086
rect 1339 -1087 1375 -1086
rect 1409 -1087 1452 -1086
rect 142 -1089 570 -1088
rect 628 -1089 1452 -1088
rect 142 -1091 150 -1090
rect 166 -1091 199 -1090
rect 219 -1091 248 -1090
rect 261 -1091 829 -1090
rect 845 -1091 1151 -1090
rect 1241 -1091 1298 -1090
rect 1311 -1091 1438 -1090
rect 149 -1093 304 -1092
rect 310 -1093 332 -1092
rect 359 -1093 416 -1092
rect 513 -1093 577 -1092
rect 702 -1093 1424 -1092
rect 1437 -1093 1459 -1092
rect 170 -1095 409 -1094
rect 516 -1095 759 -1094
rect 786 -1095 843 -1094
rect 859 -1095 1515 -1094
rect 170 -1097 192 -1096
rect 212 -1097 304 -1096
rect 331 -1097 346 -1096
rect 359 -1097 486 -1096
rect 520 -1097 542 -1096
rect 733 -1097 1221 -1096
rect 1297 -1097 1417 -1096
rect 1458 -1097 1473 -1096
rect 47 -1099 542 -1098
rect 744 -1099 997 -1098
rect 1010 -1099 1095 -1098
rect 1122 -1099 1179 -1098
rect 1346 -1099 1424 -1098
rect 1472 -1099 1529 -1098
rect 79 -1101 192 -1100
rect 212 -1101 255 -1100
rect 282 -1101 346 -1100
rect 366 -1101 475 -1100
rect 485 -1101 1536 -1100
rect 79 -1103 1557 -1102
rect 163 -1105 255 -1104
rect 275 -1105 283 -1104
rect 289 -1105 318 -1104
rect 366 -1105 552 -1104
rect 793 -1105 1585 -1104
rect 114 -1107 318 -1106
rect 380 -1107 696 -1106
rect 807 -1107 1074 -1106
rect 1115 -1107 1585 -1106
rect 114 -1109 780 -1108
rect 842 -1109 1046 -1108
rect 1073 -1109 1088 -1108
rect 1115 -1109 1172 -1108
rect 1178 -1109 1214 -1108
rect 1332 -1109 1347 -1108
rect 1374 -1109 1606 -1108
rect 156 -1111 276 -1110
rect 380 -1111 468 -1110
rect 723 -1111 1214 -1110
rect 1528 -1111 1543 -1110
rect 1556 -1111 1578 -1110
rect 156 -1113 647 -1112
rect 772 -1113 780 -1112
rect 849 -1113 1333 -1112
rect 1542 -1113 1662 -1112
rect 75 -1115 850 -1114
rect 856 -1115 1095 -1114
rect 1150 -1115 1249 -1114
rect 177 -1117 626 -1116
rect 646 -1117 668 -1116
rect 674 -1117 773 -1116
rect 835 -1117 857 -1116
rect 870 -1117 1060 -1116
rect 1164 -1117 1172 -1116
rect 1248 -1117 1326 -1116
rect 177 -1119 1665 -1118
rect 201 -1121 1088 -1120
rect 1164 -1121 1263 -1120
rect 201 -1123 458 -1122
rect 537 -1123 675 -1122
rect 821 -1123 871 -1122
rect 873 -1123 1494 -1122
rect 205 -1125 1606 -1124
rect 236 -1127 1256 -1126
rect 1353 -1127 1494 -1126
rect 240 -1129 640 -1128
rect 667 -1129 689 -1128
rect 821 -1129 1102 -1128
rect 1185 -1129 1263 -1128
rect 1353 -1129 1396 -1128
rect 58 -1131 689 -1130
rect 835 -1131 969 -1130
rect 975 -1131 1032 -1130
rect 1038 -1131 1207 -1130
rect 1395 -1131 1445 -1130
rect 58 -1133 664 -1132
rect 877 -1133 1620 -1132
rect 247 -1135 269 -1134
rect 387 -1135 605 -1134
rect 625 -1135 955 -1134
rect 978 -1135 1578 -1134
rect 163 -1137 269 -1136
rect 394 -1137 881 -1136
rect 894 -1137 1417 -1136
rect 1444 -1137 1508 -1136
rect 226 -1139 388 -1138
rect 394 -1139 755 -1138
rect 877 -1139 885 -1138
rect 898 -1139 1634 -1138
rect 30 -1141 227 -1140
rect 401 -1141 594 -1140
rect 639 -1141 738 -1140
rect 898 -1141 1508 -1140
rect 1598 -1141 1634 -1140
rect 30 -1143 584 -1142
rect 709 -1143 738 -1142
rect 912 -1143 969 -1142
rect 989 -1143 1690 -1142
rect 233 -1145 584 -1144
rect 709 -1145 1067 -1144
rect 1101 -1145 1158 -1144
rect 1563 -1145 1599 -1144
rect 422 -1147 787 -1146
rect 912 -1147 927 -1146
rect 933 -1147 1326 -1146
rect 1563 -1147 1592 -1146
rect 422 -1149 549 -1148
rect 726 -1149 927 -1148
rect 947 -1149 983 -1148
rect 989 -1149 1403 -1148
rect 1591 -1149 1648 -1148
rect 324 -1151 549 -1150
rect 765 -1151 934 -1150
rect 954 -1151 1571 -1150
rect 1647 -1151 1718 -1150
rect 100 -1153 325 -1152
rect 429 -1153 794 -1152
rect 814 -1153 983 -1152
rect 992 -1153 1207 -1152
rect 1570 -1153 1683 -1152
rect 373 -1155 430 -1154
rect 457 -1155 612 -1154
rect 814 -1155 864 -1154
rect 919 -1155 962 -1154
rect 992 -1155 1487 -1154
rect 373 -1157 661 -1156
rect 800 -1157 864 -1156
rect 996 -1157 1025 -1156
rect 1031 -1157 1109 -1156
rect 1157 -1157 1284 -1156
rect 1486 -1157 1704 -1156
rect 338 -1159 801 -1158
rect 831 -1159 962 -1158
rect 1003 -1159 1186 -1158
rect 1283 -1159 1319 -1158
rect 184 -1161 339 -1160
rect 471 -1161 885 -1160
rect 957 -1161 1319 -1160
rect 37 -1163 472 -1162
rect 562 -1163 766 -1162
rect 1003 -1163 1053 -1162
rect 37 -1165 73 -1164
rect 124 -1165 1053 -1164
rect 184 -1167 479 -1166
rect 492 -1167 563 -1166
rect 611 -1167 892 -1166
rect 1017 -1167 1067 -1166
rect 492 -1169 762 -1168
rect 1017 -1169 1081 -1168
rect 635 -1171 1109 -1170
rect 660 -1173 1200 -1172
rect 901 -1175 1200 -1174
rect 1024 -1177 1137 -1176
rect 1080 -1179 1270 -1178
rect 1136 -1181 1193 -1180
rect 1269 -1181 1305 -1180
rect 597 -1183 1193 -1182
rect 607 -1185 1305 -1184
rect 23 -1196 66 -1195
rect 79 -1196 101 -1195
rect 124 -1196 1116 -1195
rect 1486 -1196 1690 -1195
rect 1717 -1196 1725 -1195
rect 1731 -1196 1739 -1195
rect 30 -1198 90 -1197
rect 93 -1198 146 -1197
rect 149 -1198 206 -1197
rect 208 -1198 794 -1197
rect 810 -1198 836 -1197
rect 873 -1198 1599 -1197
rect 1605 -1198 1683 -1197
rect 30 -1200 489 -1199
rect 506 -1200 696 -1199
rect 723 -1200 1186 -1199
rect 1451 -1200 1487 -1199
rect 1500 -1200 1599 -1199
rect 1619 -1200 1669 -1199
rect 1675 -1200 1732 -1199
rect 58 -1202 122 -1201
rect 135 -1202 514 -1201
rect 541 -1202 710 -1201
rect 744 -1202 1137 -1201
rect 1185 -1202 1326 -1201
rect 1465 -1202 1620 -1201
rect 1654 -1202 1676 -1201
rect 58 -1204 248 -1203
rect 250 -1204 353 -1203
rect 380 -1204 724 -1203
rect 744 -1204 780 -1203
rect 814 -1204 899 -1203
rect 901 -1204 1445 -1203
rect 1591 -1204 1606 -1203
rect 1661 -1204 1725 -1203
rect 65 -1206 202 -1205
rect 205 -1206 577 -1205
rect 593 -1206 1403 -1205
rect 1416 -1206 1466 -1205
rect 1542 -1206 1662 -1205
rect 96 -1208 1515 -1207
rect 1528 -1208 1543 -1207
rect 121 -1210 1522 -1209
rect 135 -1212 360 -1211
rect 380 -1212 388 -1211
rect 422 -1212 517 -1211
rect 530 -1212 1137 -1211
rect 1206 -1212 1445 -1211
rect 1521 -1212 1571 -1211
rect 142 -1214 150 -1213
rect 163 -1214 1298 -1213
rect 1325 -1214 1396 -1213
rect 1416 -1214 1480 -1213
rect 142 -1216 1123 -1215
rect 1129 -1216 1207 -1215
rect 1241 -1216 1298 -1215
rect 1339 -1216 1403 -1215
rect 1409 -1216 1480 -1215
rect 124 -1218 1410 -1217
rect 1437 -1218 1655 -1217
rect 163 -1220 1193 -1219
rect 1213 -1220 1242 -1219
rect 1290 -1220 1438 -1219
rect 166 -1222 486 -1221
rect 492 -1222 780 -1221
rect 814 -1222 1641 -1221
rect 166 -1224 465 -1223
rect 492 -1224 640 -1223
rect 674 -1224 717 -1223
rect 768 -1224 1697 -1223
rect 184 -1226 689 -1225
rect 695 -1226 979 -1225
rect 982 -1226 1000 -1225
rect 1013 -1226 1368 -1225
rect 1374 -1226 1641 -1225
rect 82 -1228 185 -1227
rect 198 -1228 468 -1227
rect 513 -1228 1501 -1227
rect 198 -1230 626 -1229
rect 639 -1230 654 -1229
rect 709 -1230 720 -1229
rect 772 -1230 836 -1229
rect 894 -1230 913 -1229
rect 936 -1230 1627 -1229
rect 156 -1232 626 -1231
rect 646 -1232 675 -1231
rect 828 -1232 1515 -1231
rect 1535 -1232 1627 -1231
rect 156 -1234 619 -1233
rect 646 -1234 664 -1233
rect 831 -1234 941 -1233
rect 957 -1234 1578 -1233
rect 233 -1236 332 -1235
rect 352 -1236 451 -1235
rect 478 -1236 773 -1235
rect 884 -1236 941 -1235
rect 971 -1236 1585 -1235
rect 212 -1238 332 -1237
rect 387 -1238 500 -1237
rect 576 -1238 1529 -1237
rect 191 -1240 213 -1239
rect 233 -1240 500 -1239
rect 597 -1240 1578 -1239
rect 177 -1242 192 -1241
rect 236 -1242 1452 -1241
rect 1472 -1242 1536 -1241
rect 177 -1244 220 -1243
rect 240 -1244 619 -1243
rect 653 -1244 951 -1243
rect 975 -1244 1193 -1243
rect 1276 -1244 1291 -1243
rect 1356 -1244 1585 -1243
rect 219 -1246 818 -1245
rect 821 -1246 885 -1245
rect 898 -1246 906 -1245
rect 975 -1246 993 -1245
rect 1045 -1246 1557 -1245
rect 152 -1248 906 -1247
rect 982 -1248 1263 -1247
rect 1381 -1248 1571 -1247
rect 240 -1250 622 -1249
rect 821 -1250 1011 -1249
rect 1031 -1250 1263 -1249
rect 1395 -1250 1735 -1249
rect 254 -1252 346 -1251
rect 394 -1252 465 -1251
rect 478 -1252 528 -1251
rect 544 -1252 1382 -1251
rect 1423 -1252 1473 -1251
rect 1556 -1252 1648 -1251
rect 37 -1254 528 -1253
rect 562 -1254 598 -1253
rect 611 -1254 692 -1253
rect 989 -1254 1060 -1253
rect 1080 -1254 1368 -1253
rect 1388 -1254 1424 -1253
rect 1612 -1254 1648 -1253
rect 37 -1256 549 -1255
rect 614 -1256 1592 -1255
rect 278 -1258 808 -1257
rect 989 -1258 1088 -1257
rect 1108 -1258 1340 -1257
rect 1549 -1258 1613 -1257
rect 310 -1260 510 -1259
rect 548 -1260 556 -1259
rect 751 -1260 1389 -1259
rect 1493 -1260 1550 -1259
rect 310 -1262 461 -1261
rect 471 -1262 563 -1261
rect 751 -1262 759 -1261
rect 807 -1262 1116 -1261
rect 1129 -1262 1228 -1261
rect 1255 -1262 1494 -1261
rect 317 -1264 727 -1263
rect 1003 -1264 1060 -1263
rect 1108 -1264 1354 -1263
rect 282 -1266 318 -1265
rect 324 -1266 360 -1265
rect 394 -1266 871 -1265
rect 1003 -1266 1235 -1265
rect 1353 -1266 1375 -1265
rect 170 -1268 325 -1267
rect 345 -1268 409 -1267
rect 429 -1268 517 -1267
rect 555 -1268 832 -1267
rect 870 -1268 1018 -1267
rect 1024 -1268 1088 -1267
rect 1143 -1268 1214 -1267
rect 1220 -1268 1277 -1267
rect 170 -1270 605 -1269
rect 877 -1270 1221 -1269
rect 282 -1272 986 -1271
rect 996 -1272 1025 -1271
rect 1045 -1272 1165 -1271
rect 1171 -1272 1256 -1271
rect 338 -1274 430 -1273
rect 443 -1274 447 -1273
rect 450 -1274 584 -1273
rect 590 -1274 878 -1273
rect 933 -1274 997 -1273
rect 1010 -1274 1081 -1273
rect 1094 -1274 1172 -1273
rect 1199 -1274 1228 -1273
rect 86 -1276 584 -1275
rect 933 -1276 1067 -1275
rect 1094 -1276 1158 -1275
rect 1164 -1276 1179 -1275
rect 261 -1278 339 -1277
rect 408 -1278 416 -1277
rect 443 -1278 521 -1277
rect 534 -1278 605 -1277
rect 947 -1278 1018 -1277
rect 1048 -1278 1431 -1277
rect 44 -1280 535 -1279
rect 569 -1280 759 -1279
rect 947 -1280 1714 -1279
rect 44 -1282 76 -1281
rect 226 -1282 570 -1281
rect 954 -1282 1235 -1281
rect 1360 -1282 1431 -1281
rect 75 -1284 87 -1283
rect 226 -1284 458 -1283
rect 471 -1284 748 -1283
rect 863 -1284 955 -1283
rect 961 -1284 1067 -1283
rect 1101 -1284 1144 -1283
rect 1150 -1284 1200 -1283
rect 1304 -1284 1361 -1283
rect 261 -1286 423 -1285
rect 425 -1286 1305 -1285
rect 415 -1288 682 -1287
rect 702 -1288 962 -1287
rect 968 -1288 1179 -1287
rect 366 -1290 682 -1289
rect 800 -1290 864 -1289
rect 919 -1290 969 -1289
rect 999 -1290 1032 -1289
rect 1038 -1290 1151 -1289
rect 1157 -1290 1284 -1289
rect 128 -1292 801 -1291
rect 842 -1292 1102 -1291
rect 107 -1294 129 -1293
rect 303 -1294 367 -1293
rect 509 -1294 668 -1293
rect 842 -1294 857 -1293
rect 1052 -1294 1123 -1293
rect 107 -1296 269 -1295
rect 303 -1296 402 -1295
rect 628 -1296 668 -1295
rect 828 -1296 857 -1295
rect 1052 -1296 1564 -1295
rect 114 -1298 402 -1297
rect 632 -1298 703 -1297
rect 849 -1298 920 -1297
rect 1055 -1298 1312 -1297
rect 1507 -1298 1564 -1297
rect 114 -1300 689 -1299
rect 765 -1300 850 -1299
rect 1073 -1300 1284 -1299
rect 1311 -1300 1347 -1299
rect 1458 -1300 1508 -1299
rect 268 -1302 290 -1301
rect 373 -1302 633 -1301
rect 660 -1302 1039 -1301
rect 1458 -1302 1665 -1301
rect 51 -1304 290 -1303
rect 373 -1304 437 -1303
rect 660 -1304 738 -1303
rect 765 -1304 913 -1303
rect 51 -1306 615 -1305
rect 730 -1306 738 -1305
rect 786 -1306 1074 -1305
rect 257 -1308 437 -1307
rect 481 -1308 731 -1307
rect 786 -1308 1249 -1307
rect 891 -1310 1347 -1309
rect 891 -1312 927 -1311
rect 1248 -1312 1333 -1311
rect 82 -1314 927 -1313
rect 1269 -1314 1333 -1313
rect 93 -1316 1270 -1315
rect 16 -1327 52 -1326
rect 58 -1327 423 -1326
rect 478 -1327 1375 -1326
rect 1493 -1327 1732 -1326
rect 1738 -1327 1746 -1326
rect 37 -1329 423 -1328
rect 478 -1329 521 -1328
rect 579 -1329 1277 -1328
rect 1346 -1329 1707 -1328
rect 1717 -1329 1735 -1328
rect 37 -1331 230 -1330
rect 233 -1331 283 -1330
rect 289 -1331 528 -1330
rect 597 -1331 766 -1330
rect 768 -1331 1172 -1330
rect 1276 -1331 1361 -1330
rect 1493 -1331 1522 -1330
rect 1626 -1331 1721 -1330
rect 44 -1333 73 -1332
rect 82 -1333 1298 -1332
rect 1521 -1333 1592 -1332
rect 1675 -1333 1704 -1332
rect 44 -1335 199 -1334
rect 240 -1335 832 -1334
rect 873 -1335 1424 -1334
rect 1584 -1335 1627 -1334
rect 1682 -1335 1718 -1334
rect 51 -1337 626 -1336
rect 628 -1337 780 -1336
rect 786 -1337 843 -1336
rect 901 -1337 1095 -1336
rect 1125 -1337 1592 -1336
rect 1696 -1337 1711 -1336
rect 75 -1339 241 -1338
rect 250 -1339 1305 -1338
rect 1699 -1339 1725 -1338
rect 82 -1341 1340 -1340
rect 86 -1343 97 -1342
rect 124 -1343 150 -1342
rect 170 -1343 734 -1342
rect 765 -1343 1375 -1342
rect 93 -1345 1263 -1344
rect 1283 -1345 1676 -1344
rect 96 -1347 325 -1346
rect 366 -1347 577 -1346
rect 590 -1347 626 -1346
rect 632 -1347 787 -1346
rect 796 -1347 1361 -1346
rect 107 -1349 171 -1348
rect 177 -1349 237 -1348
rect 264 -1349 318 -1348
rect 324 -1349 542 -1348
rect 548 -1349 577 -1348
rect 597 -1349 1102 -1348
rect 1136 -1349 1725 -1348
rect 107 -1351 1508 -1350
rect 135 -1353 458 -1352
rect 460 -1353 1347 -1352
rect 135 -1355 503 -1354
rect 506 -1355 633 -1354
rect 653 -1355 818 -1354
rect 821 -1355 1193 -1354
rect 1262 -1355 1319 -1354
rect 1339 -1355 1550 -1354
rect 142 -1357 808 -1356
rect 828 -1357 1641 -1356
rect 30 -1359 143 -1358
rect 149 -1359 563 -1358
rect 593 -1359 1641 -1358
rect 26 -1361 31 -1360
rect 177 -1361 185 -1360
rect 191 -1361 199 -1360
rect 219 -1361 507 -1360
rect 520 -1361 892 -1360
rect 947 -1361 1543 -1360
rect 117 -1363 1543 -1362
rect 163 -1365 185 -1364
rect 219 -1365 255 -1364
rect 275 -1365 451 -1364
rect 457 -1365 731 -1364
rect 779 -1365 836 -1364
rect 891 -1365 990 -1364
rect 1010 -1365 1214 -1364
rect 1297 -1365 1312 -1364
rect 114 -1367 255 -1366
rect 275 -1367 332 -1366
rect 366 -1367 692 -1366
rect 695 -1367 895 -1366
rect 947 -1367 969 -1366
rect 978 -1367 1613 -1366
rect 156 -1369 164 -1368
rect 247 -1369 1319 -1368
rect 1612 -1369 1634 -1368
rect 156 -1371 192 -1370
rect 247 -1371 279 -1370
rect 282 -1371 346 -1370
rect 373 -1371 1508 -1370
rect 1605 -1371 1634 -1370
rect 289 -1373 419 -1372
rect 436 -1373 542 -1372
rect 548 -1373 556 -1372
rect 562 -1373 605 -1372
rect 614 -1373 822 -1372
rect 828 -1373 864 -1372
rect 968 -1373 1025 -1372
rect 1027 -1373 1585 -1372
rect 296 -1375 612 -1374
rect 618 -1375 664 -1374
rect 667 -1375 990 -1374
rect 1045 -1375 1049 -1374
rect 1055 -1375 1333 -1374
rect 1416 -1375 1606 -1374
rect 303 -1377 346 -1376
rect 352 -1377 615 -1376
rect 639 -1377 668 -1376
rect 688 -1377 1480 -1376
rect 317 -1379 790 -1378
rect 835 -1379 937 -1378
rect 982 -1379 1417 -1378
rect 1479 -1379 1515 -1378
rect 331 -1381 500 -1380
rect 590 -1381 1515 -1380
rect 352 -1383 409 -1382
rect 415 -1383 437 -1382
rect 450 -1383 773 -1382
rect 863 -1383 1109 -1382
rect 1129 -1383 1193 -1382
rect 1213 -1383 1256 -1382
rect 1304 -1383 1410 -1382
rect 338 -1385 409 -1384
rect 415 -1385 535 -1384
rect 604 -1385 636 -1384
rect 639 -1385 1074 -1384
rect 1094 -1385 1207 -1384
rect 1255 -1385 1403 -1384
rect 261 -1387 339 -1386
rect 373 -1387 584 -1386
rect 611 -1387 1424 -1386
rect 261 -1389 1102 -1388
rect 1146 -1389 1655 -1388
rect 387 -1391 528 -1390
rect 534 -1391 857 -1390
rect 877 -1391 937 -1390
rect 940 -1391 983 -1390
rect 985 -1391 1690 -1390
rect 303 -1393 388 -1392
rect 394 -1393 1011 -1392
rect 1017 -1393 1109 -1392
rect 1171 -1393 1242 -1392
rect 1311 -1393 1445 -1392
rect 1654 -1393 1662 -1392
rect 205 -1395 395 -1394
rect 401 -1395 843 -1394
rect 877 -1395 899 -1394
rect 905 -1395 1074 -1394
rect 1139 -1395 1242 -1394
rect 1325 -1395 1410 -1394
rect 79 -1397 899 -1396
rect 940 -1397 962 -1396
rect 1017 -1397 1067 -1396
rect 1069 -1397 1648 -1396
rect 110 -1399 206 -1398
rect 401 -1399 444 -1398
rect 464 -1399 619 -1398
rect 653 -1399 710 -1398
rect 719 -1399 955 -1398
rect 1045 -1399 1088 -1398
rect 1185 -1399 1284 -1398
rect 1332 -1399 1389 -1398
rect 1402 -1399 1459 -1398
rect 1619 -1399 1648 -1398
rect 121 -1401 1389 -1400
rect 1458 -1401 1487 -1400
rect 121 -1403 381 -1402
rect 464 -1403 647 -1402
rect 660 -1403 1221 -1402
rect 1353 -1403 1662 -1402
rect 128 -1405 647 -1404
rect 660 -1405 976 -1404
rect 1087 -1405 1151 -1404
rect 1185 -1405 1382 -1404
rect 1486 -1405 1529 -1404
rect 128 -1407 360 -1406
rect 380 -1407 430 -1406
rect 485 -1407 727 -1406
rect 730 -1407 1550 -1406
rect 23 -1409 486 -1408
rect 499 -1409 1620 -1408
rect 65 -1411 430 -1410
rect 513 -1411 1067 -1410
rect 1206 -1411 1291 -1410
rect 1353 -1411 1438 -1410
rect 1528 -1411 1571 -1410
rect 65 -1413 223 -1412
rect 226 -1413 444 -1412
rect 555 -1413 1690 -1412
rect 310 -1415 360 -1414
rect 583 -1415 1014 -1414
rect 1048 -1415 1151 -1414
rect 1157 -1415 1291 -1414
rect 310 -1417 472 -1416
rect 677 -1417 1221 -1416
rect 1248 -1417 1382 -1416
rect 58 -1419 472 -1418
rect 688 -1419 703 -1418
rect 709 -1419 717 -1418
rect 723 -1419 794 -1418
rect 800 -1419 1130 -1418
rect 1248 -1419 1396 -1418
rect 695 -1421 759 -1420
rect 800 -1421 850 -1420
rect 866 -1421 1571 -1420
rect 702 -1423 1032 -1422
rect 1395 -1423 1452 -1422
rect 61 -1425 1032 -1424
rect 1430 -1425 1452 -1424
rect 716 -1427 1158 -1426
rect 1430 -1427 1466 -1426
rect 226 -1429 1466 -1428
rect 723 -1431 1368 -1430
rect 744 -1433 794 -1432
rect 814 -1433 906 -1432
rect 919 -1433 962 -1432
rect 975 -1433 997 -1432
rect 1367 -1433 1473 -1432
rect 737 -1435 745 -1434
rect 751 -1435 773 -1434
rect 814 -1435 885 -1434
rect 919 -1435 1060 -1434
rect 1472 -1435 1501 -1434
rect 145 -1437 752 -1436
rect 758 -1437 871 -1436
rect 933 -1437 1438 -1436
rect 1500 -1437 1536 -1436
rect 569 -1439 738 -1438
rect 824 -1439 1445 -1438
rect 1535 -1439 1578 -1438
rect 509 -1441 570 -1440
rect 681 -1441 885 -1440
rect 933 -1441 1683 -1440
rect 674 -1443 682 -1442
rect 849 -1443 927 -1442
rect 954 -1443 1144 -1442
rect 1577 -1443 1599 -1442
rect 492 -1445 675 -1444
rect 856 -1445 871 -1444
rect 926 -1445 1004 -1444
rect 1059 -1445 1123 -1444
rect 1143 -1445 1326 -1444
rect 1563 -1445 1599 -1444
rect 86 -1447 1123 -1446
rect 1227 -1447 1564 -1446
rect 93 -1449 493 -1448
rect 530 -1449 1228 -1448
rect 996 -1451 1039 -1450
rect 1003 -1453 1200 -1452
rect 600 -1455 1200 -1454
rect 1038 -1457 1116 -1456
rect 1115 -1459 1165 -1458
rect 1164 -1461 1235 -1460
rect 1080 -1463 1235 -1462
rect 1080 -1465 1179 -1464
rect 1052 -1467 1179 -1466
rect 912 -1469 1053 -1468
rect 642 -1471 913 -1470
rect 16 -1482 766 -1481
rect 786 -1482 864 -1481
rect 870 -1482 920 -1481
rect 1024 -1482 1095 -1481
rect 1104 -1482 1340 -1481
rect 1745 -1482 1753 -1481
rect 23 -1484 76 -1483
rect 96 -1484 1641 -1483
rect 30 -1486 83 -1485
rect 107 -1486 416 -1485
rect 418 -1486 766 -1485
rect 786 -1486 906 -1485
rect 1024 -1486 1088 -1485
rect 1118 -1486 1711 -1485
rect 58 -1488 1690 -1487
rect 61 -1490 118 -1489
rect 142 -1490 209 -1489
rect 226 -1490 360 -1489
rect 373 -1490 762 -1489
rect 863 -1490 941 -1489
rect 1073 -1490 1714 -1489
rect 68 -1492 549 -1491
rect 555 -1492 612 -1491
rect 621 -1492 710 -1491
rect 719 -1492 1564 -1491
rect 1640 -1492 1669 -1491
rect 72 -1494 367 -1493
rect 390 -1494 430 -1493
rect 443 -1494 545 -1493
rect 562 -1494 710 -1493
rect 733 -1494 920 -1493
rect 1073 -1494 1144 -1493
rect 1153 -1494 1333 -1493
rect 1339 -1494 1417 -1493
rect 1493 -1494 1690 -1493
rect 44 -1496 73 -1495
rect 107 -1496 367 -1495
rect 394 -1496 769 -1495
rect 866 -1496 1095 -1495
rect 1122 -1496 1263 -1495
rect 1311 -1496 1333 -1495
rect 1416 -1496 1487 -1495
rect 1493 -1496 1536 -1495
rect 1563 -1496 1592 -1495
rect 1612 -1496 1669 -1495
rect 44 -1498 370 -1497
rect 394 -1498 472 -1497
rect 474 -1498 962 -1497
rect 989 -1498 1123 -1497
rect 1125 -1498 1704 -1497
rect 30 -1500 472 -1499
rect 492 -1500 902 -1499
rect 905 -1500 927 -1499
rect 961 -1500 969 -1499
rect 975 -1500 990 -1499
rect 1087 -1500 1172 -1499
rect 1311 -1500 1326 -1499
rect 1486 -1500 1606 -1499
rect 114 -1502 437 -1501
rect 443 -1502 1704 -1501
rect 114 -1504 671 -1503
rect 677 -1504 1550 -1503
rect 1556 -1504 1606 -1503
rect 142 -1506 402 -1505
rect 422 -1506 594 -1505
rect 607 -1506 668 -1505
rect 730 -1506 1263 -1505
rect 1325 -1506 1403 -1505
rect 1500 -1506 1613 -1505
rect 51 -1508 402 -1507
rect 436 -1508 930 -1507
rect 975 -1508 1347 -1507
rect 1402 -1508 1473 -1507
rect 1535 -1508 1578 -1507
rect 1584 -1508 1592 -1507
rect 156 -1510 1557 -1509
rect 1570 -1510 1578 -1509
rect 1584 -1510 1599 -1509
rect 156 -1512 213 -1511
rect 226 -1512 258 -1511
rect 261 -1512 283 -1511
rect 296 -1512 619 -1511
rect 632 -1512 1046 -1511
rect 1048 -1512 1571 -1511
rect 1598 -1512 1620 -1511
rect 159 -1514 584 -1513
rect 635 -1514 1508 -1513
rect 1549 -1514 1721 -1513
rect 149 -1516 584 -1515
rect 639 -1516 1707 -1515
rect 149 -1518 559 -1517
rect 562 -1518 682 -1517
rect 712 -1518 1501 -1517
rect 1619 -1518 1634 -1517
rect 191 -1520 220 -1519
rect 229 -1520 983 -1519
rect 1045 -1520 1130 -1519
rect 1139 -1520 1452 -1519
rect 1472 -1520 1655 -1519
rect 194 -1522 535 -1521
rect 541 -1522 556 -1521
rect 576 -1522 598 -1521
rect 604 -1522 682 -1521
rect 730 -1522 780 -1521
rect 796 -1522 1634 -1521
rect 79 -1524 577 -1523
rect 604 -1524 1683 -1523
rect 79 -1526 164 -1525
rect 212 -1526 241 -1525
rect 268 -1526 283 -1525
rect 310 -1526 416 -1525
rect 450 -1526 493 -1525
rect 499 -1526 619 -1525
rect 639 -1526 661 -1525
rect 747 -1526 815 -1525
rect 870 -1526 1018 -1525
rect 1020 -1526 1655 -1525
rect 121 -1528 241 -1527
rect 299 -1528 311 -1527
rect 331 -1528 423 -1527
rect 450 -1528 675 -1527
rect 779 -1528 801 -1527
rect 891 -1528 1137 -1527
rect 1143 -1528 1207 -1527
rect 1283 -1528 1683 -1527
rect 93 -1530 122 -1529
rect 163 -1530 591 -1529
rect 660 -1530 696 -1529
rect 719 -1530 1284 -1529
rect 1346 -1530 1424 -1529
rect 1451 -1530 1543 -1529
rect 93 -1532 626 -1531
rect 674 -1532 738 -1531
rect 793 -1532 815 -1531
rect 891 -1532 997 -1531
rect 1017 -1532 1676 -1531
rect 51 -1534 794 -1533
rect 800 -1534 843 -1533
rect 898 -1534 948 -1533
rect 982 -1534 1158 -1533
rect 1171 -1534 1235 -1533
rect 1258 -1534 1424 -1533
rect 1521 -1534 1543 -1533
rect 1626 -1534 1676 -1533
rect 205 -1536 332 -1535
rect 338 -1536 374 -1535
rect 464 -1536 633 -1535
rect 737 -1536 969 -1535
rect 996 -1536 1060 -1535
rect 1062 -1536 1158 -1535
rect 1199 -1536 1508 -1535
rect 1521 -1536 1662 -1535
rect 191 -1538 1200 -1537
rect 1206 -1538 1361 -1537
rect 1661 -1538 1711 -1537
rect 205 -1540 913 -1539
rect 926 -1540 1291 -1539
rect 219 -1542 248 -1541
rect 303 -1542 465 -1541
rect 502 -1542 689 -1541
rect 758 -1542 913 -1541
rect 933 -1542 1627 -1541
rect 184 -1544 248 -1543
rect 324 -1544 696 -1543
rect 758 -1544 1186 -1543
rect 1227 -1544 1361 -1543
rect 135 -1546 185 -1545
rect 233 -1546 304 -1545
rect 338 -1546 384 -1545
rect 506 -1546 717 -1545
rect 842 -1546 1067 -1545
rect 1129 -1546 1214 -1545
rect 1227 -1546 1725 -1545
rect 37 -1548 136 -1547
rect 233 -1548 388 -1547
rect 457 -1548 507 -1547
rect 520 -1548 1147 -1547
rect 1185 -1548 1242 -1547
rect 1290 -1548 1298 -1547
rect 86 -1550 388 -1549
rect 457 -1550 486 -1549
rect 527 -1550 535 -1549
rect 569 -1550 598 -1549
rect 625 -1550 741 -1549
rect 933 -1550 937 -1549
rect 947 -1550 1032 -1549
rect 1213 -1550 1354 -1549
rect 65 -1552 570 -1551
rect 590 -1552 808 -1551
rect 1031 -1552 1116 -1551
rect 1234 -1552 1256 -1551
rect 1297 -1552 1396 -1551
rect 65 -1554 941 -1553
rect 1241 -1554 1319 -1553
rect 1353 -1554 1438 -1553
rect 86 -1556 836 -1555
rect 873 -1556 1256 -1555
rect 1318 -1556 1375 -1555
rect 1437 -1556 1529 -1555
rect 128 -1558 521 -1557
rect 527 -1558 1718 -1557
rect 128 -1560 276 -1559
rect 345 -1560 430 -1559
rect 485 -1560 752 -1559
rect 807 -1560 1697 -1559
rect 170 -1562 836 -1561
rect 1115 -1562 1529 -1561
rect 170 -1564 353 -1563
rect 359 -1564 479 -1563
rect 667 -1564 1067 -1563
rect 1367 -1564 1375 -1563
rect 254 -1566 325 -1565
rect 352 -1566 381 -1565
rect 478 -1566 829 -1565
rect 1367 -1566 1445 -1565
rect 275 -1568 318 -1567
rect 380 -1568 727 -1567
rect 751 -1568 773 -1567
rect 821 -1568 1396 -1567
rect 1430 -1568 1445 -1567
rect 289 -1570 346 -1569
rect 688 -1570 1011 -1569
rect 1430 -1570 1466 -1569
rect 177 -1572 290 -1571
rect 614 -1572 1466 -1571
rect 177 -1574 412 -1573
rect 716 -1574 1109 -1573
rect 723 -1576 1718 -1575
rect 723 -1578 745 -1577
rect 772 -1578 857 -1577
rect 1010 -1578 1053 -1577
rect 1108 -1578 1193 -1577
rect 548 -1580 745 -1579
rect 821 -1580 1165 -1579
rect 1192 -1580 1270 -1579
rect 614 -1582 1270 -1581
rect 726 -1584 955 -1583
rect 1052 -1584 1081 -1583
rect 1164 -1584 1221 -1583
rect 828 -1586 878 -1585
rect 954 -1586 1102 -1585
rect 1220 -1586 1249 -1585
rect 849 -1588 857 -1587
rect 877 -1588 885 -1587
rect 1080 -1588 1151 -1587
rect 1248 -1588 1305 -1587
rect 702 -1590 885 -1589
rect 1101 -1590 1382 -1589
rect 292 -1592 703 -1591
rect 849 -1592 1004 -1591
rect 1304 -1592 1410 -1591
rect 541 -1594 1410 -1593
rect 1003 -1596 1039 -1595
rect 1381 -1596 1459 -1595
rect 1038 -1598 1179 -1597
rect 1458 -1598 1480 -1597
rect 1178 -1600 1277 -1599
rect 1479 -1600 1648 -1599
rect 264 -1602 1648 -1601
rect 1276 -1604 1389 -1603
rect 1388 -1606 1515 -1605
rect 642 -1608 1515 -1607
rect 16 -1619 31 -1618
rect 37 -1619 290 -1618
rect 296 -1619 384 -1618
rect 411 -1619 745 -1618
rect 758 -1619 1105 -1618
rect 1115 -1619 1319 -1618
rect 1381 -1619 1385 -1618
rect 1479 -1619 1725 -1618
rect 1752 -1619 1767 -1618
rect 44 -1621 255 -1620
rect 268 -1621 311 -1620
rect 317 -1621 916 -1620
rect 929 -1621 1683 -1620
rect 1717 -1621 1781 -1620
rect 44 -1623 346 -1622
rect 348 -1623 920 -1622
rect 996 -1623 1774 -1622
rect 58 -1625 1543 -1624
rect 1626 -1625 1732 -1624
rect 65 -1627 496 -1626
rect 513 -1627 727 -1626
rect 730 -1627 759 -1626
rect 761 -1627 1662 -1626
rect 1668 -1627 1704 -1626
rect 79 -1629 265 -1628
rect 268 -1629 321 -1628
rect 324 -1629 367 -1628
rect 369 -1629 416 -1628
rect 432 -1629 458 -1628
rect 478 -1629 615 -1628
rect 667 -1629 815 -1628
rect 828 -1629 895 -1628
rect 919 -1629 923 -1628
rect 975 -1629 1662 -1628
rect 23 -1631 367 -1630
rect 387 -1631 458 -1630
rect 513 -1631 608 -1630
rect 667 -1631 696 -1630
rect 712 -1631 1025 -1630
rect 1048 -1631 1613 -1630
rect 1640 -1631 1739 -1630
rect 61 -1633 388 -1632
rect 450 -1633 790 -1632
rect 793 -1633 1396 -1632
rect 1486 -1633 1669 -1632
rect 79 -1635 549 -1634
rect 562 -1635 1319 -1634
rect 1381 -1635 1403 -1634
rect 1500 -1635 1627 -1634
rect 1640 -1635 1676 -1634
rect 121 -1637 545 -1636
rect 548 -1637 556 -1636
rect 576 -1637 927 -1636
rect 975 -1637 1459 -1636
rect 1514 -1637 1683 -1636
rect 121 -1639 717 -1638
rect 726 -1639 899 -1638
rect 996 -1639 1039 -1638
rect 1059 -1639 1445 -1638
rect 1521 -1639 1718 -1638
rect 135 -1641 619 -1640
rect 674 -1641 741 -1640
rect 803 -1641 815 -1640
rect 863 -1641 1060 -1640
rect 1115 -1641 1459 -1640
rect 1591 -1641 1676 -1640
rect 135 -1643 682 -1642
rect 702 -1643 794 -1642
rect 807 -1643 1025 -1642
rect 1118 -1643 1235 -1642
rect 1241 -1643 1487 -1642
rect 1598 -1643 1704 -1642
rect 156 -1645 416 -1644
rect 450 -1645 748 -1644
rect 807 -1645 899 -1644
rect 992 -1645 1592 -1644
rect 1647 -1645 1753 -1644
rect 156 -1647 983 -1646
rect 1052 -1647 1242 -1646
rect 1251 -1647 1690 -1646
rect 170 -1649 325 -1648
rect 338 -1649 717 -1648
rect 733 -1649 969 -1648
rect 982 -1649 1018 -1648
rect 1101 -1649 1648 -1648
rect 1654 -1649 1760 -1648
rect 170 -1651 332 -1650
rect 338 -1651 647 -1650
rect 709 -1651 1039 -1650
rect 1101 -1651 1172 -1650
rect 1213 -1651 1501 -1650
rect 1689 -1651 1711 -1650
rect 191 -1653 272 -1652
rect 289 -1653 850 -1652
rect 863 -1653 885 -1652
rect 887 -1653 1431 -1652
rect 1437 -1653 1522 -1652
rect 1619 -1653 1711 -1652
rect 191 -1655 871 -1654
rect 968 -1655 990 -1654
rect 1010 -1655 1053 -1654
rect 1153 -1655 1333 -1654
rect 1367 -1655 1431 -1654
rect 1465 -1655 1599 -1654
rect 194 -1657 1557 -1656
rect 205 -1659 1235 -1658
rect 1255 -1659 1473 -1658
rect 1493 -1659 1557 -1658
rect 51 -1661 206 -1660
rect 208 -1661 1697 -1660
rect 51 -1663 409 -1662
rect 422 -1663 710 -1662
rect 737 -1663 1606 -1662
rect 177 -1665 1256 -1664
rect 1262 -1665 1445 -1664
rect 1507 -1665 1620 -1664
rect 212 -1667 311 -1666
rect 331 -1667 979 -1666
rect 1066 -1667 1473 -1666
rect 1563 -1667 1697 -1666
rect 86 -1669 213 -1668
rect 226 -1669 577 -1668
rect 597 -1669 601 -1668
rect 604 -1669 1123 -1668
rect 1206 -1669 1333 -1668
rect 1367 -1669 1550 -1668
rect 1563 -1669 1707 -1668
rect 86 -1671 143 -1670
rect 184 -1671 227 -1670
rect 233 -1671 1018 -1670
rect 1066 -1671 1438 -1670
rect 1535 -1671 1550 -1670
rect 1584 -1671 1606 -1670
rect 142 -1673 164 -1672
rect 184 -1673 199 -1672
rect 233 -1673 262 -1672
rect 278 -1673 1011 -1672
rect 1073 -1673 1123 -1672
rect 1157 -1673 1207 -1672
rect 1269 -1673 1543 -1672
rect 107 -1675 164 -1674
rect 240 -1675 423 -1674
rect 436 -1675 990 -1674
rect 1073 -1675 1228 -1674
rect 1276 -1675 1480 -1674
rect 100 -1677 108 -1676
rect 149 -1677 199 -1676
rect 240 -1677 283 -1676
rect 296 -1677 430 -1676
rect 436 -1677 661 -1676
rect 772 -1677 850 -1676
rect 870 -1677 878 -1676
rect 905 -1677 1263 -1676
rect 1304 -1677 1396 -1676
rect 1416 -1677 1494 -1676
rect 100 -1679 430 -1678
rect 478 -1679 682 -1678
rect 751 -1679 773 -1678
rect 782 -1679 1585 -1678
rect 149 -1681 678 -1680
rect 751 -1681 843 -1680
rect 877 -1681 892 -1680
rect 905 -1681 955 -1680
rect 1020 -1681 1277 -1680
rect 1339 -1681 1417 -1680
rect 1423 -1681 1515 -1680
rect 282 -1683 465 -1682
rect 492 -1683 1655 -1682
rect 359 -1685 465 -1684
rect 471 -1685 493 -1684
rect 499 -1685 696 -1684
rect 796 -1685 1214 -1684
rect 1339 -1685 1347 -1684
rect 1353 -1685 1424 -1684
rect 352 -1687 472 -1686
rect 499 -1687 521 -1686
rect 527 -1687 1634 -1686
rect 219 -1689 353 -1688
rect 359 -1689 1046 -1688
rect 1118 -1689 1508 -1688
rect 1570 -1689 1634 -1688
rect 219 -1691 276 -1690
rect 380 -1691 528 -1690
rect 534 -1691 556 -1690
rect 562 -1691 741 -1690
rect 884 -1691 955 -1690
rect 1150 -1691 1354 -1690
rect 1374 -1691 1466 -1690
rect 1528 -1691 1571 -1690
rect 173 -1693 276 -1692
rect 380 -1693 482 -1692
rect 520 -1693 724 -1692
rect 912 -1693 1158 -1692
rect 1164 -1693 1228 -1692
rect 1283 -1693 1347 -1692
rect 1374 -1693 1410 -1692
rect 177 -1695 1529 -1694
rect 443 -1697 843 -1696
rect 873 -1697 1410 -1696
rect 443 -1699 531 -1698
rect 534 -1699 566 -1698
rect 569 -1699 661 -1698
rect 723 -1699 857 -1698
rect 940 -1699 1046 -1698
rect 1087 -1699 1151 -1698
rect 1178 -1699 1305 -1698
rect 1388 -1699 1536 -1698
rect 530 -1701 836 -1700
rect 929 -1701 1088 -1700
rect 1108 -1701 1165 -1700
rect 1185 -1701 1270 -1700
rect 1297 -1701 1389 -1700
rect 128 -1703 836 -1702
rect 940 -1703 948 -1702
rect 1094 -1703 1186 -1702
rect 1199 -1703 1284 -1702
rect 1290 -1703 1298 -1702
rect 93 -1705 129 -1704
rect 541 -1705 1578 -1704
rect 93 -1707 731 -1706
rect 765 -1707 857 -1706
rect 1108 -1707 1144 -1706
rect 1192 -1707 1291 -1706
rect 1451 -1707 1578 -1706
rect 96 -1709 948 -1708
rect 1129 -1709 1144 -1708
rect 1360 -1709 1452 -1708
rect 159 -1711 1130 -1710
rect 1136 -1711 1200 -1710
rect 1325 -1711 1361 -1710
rect 247 -1713 1137 -1712
rect 1311 -1713 1326 -1712
rect 247 -1715 258 -1714
rect 506 -1715 766 -1714
rect 821 -1715 1193 -1714
rect 1248 -1715 1312 -1714
rect 394 -1717 507 -1716
rect 544 -1717 619 -1716
rect 621 -1717 1172 -1716
rect 394 -1719 402 -1718
rect 569 -1719 720 -1718
rect 800 -1719 822 -1718
rect 828 -1719 1095 -1718
rect 401 -1721 542 -1720
rect 583 -1721 605 -1720
rect 611 -1721 1613 -1720
rect 114 -1723 612 -1722
rect 646 -1723 654 -1722
rect 670 -1723 1179 -1722
rect 114 -1725 591 -1724
rect 597 -1725 626 -1724
rect 653 -1725 787 -1724
rect 800 -1725 1081 -1724
rect 303 -1727 584 -1726
rect 590 -1727 689 -1726
rect 1031 -1727 1081 -1726
rect 1384 -1727 1403 -1726
rect 303 -1729 1749 -1728
rect 688 -1731 780 -1730
rect 926 -1731 1032 -1730
rect 485 -1733 780 -1732
rect 345 -1735 486 -1734
rect 30 -1746 129 -1745
rect 159 -1746 531 -1745
rect 541 -1746 766 -1745
rect 810 -1746 878 -1745
rect 884 -1746 941 -1745
rect 978 -1746 1599 -1745
rect 1682 -1746 1795 -1745
rect 58 -1748 500 -1747
rect 502 -1748 843 -1747
rect 866 -1748 1809 -1747
rect 61 -1750 353 -1749
rect 401 -1750 941 -1749
rect 989 -1750 1648 -1749
rect 1748 -1750 1767 -1749
rect 1780 -1750 1816 -1749
rect 65 -1752 255 -1751
rect 275 -1752 416 -1751
rect 450 -1752 1249 -1751
rect 1367 -1752 1683 -1751
rect 1752 -1752 1767 -1751
rect 65 -1754 171 -1753
rect 177 -1754 1627 -1753
rect 1738 -1754 1753 -1753
rect 107 -1756 129 -1755
rect 159 -1756 297 -1755
rect 324 -1756 482 -1755
rect 618 -1756 731 -1755
rect 740 -1756 1060 -1755
rect 1069 -1756 1536 -1755
rect 1612 -1756 1648 -1755
rect 1710 -1756 1739 -1755
rect 107 -1758 1193 -1757
rect 1199 -1758 1249 -1757
rect 1332 -1758 1368 -1757
rect 1374 -1758 1536 -1757
rect 1605 -1758 1613 -1757
rect 1626 -1758 1641 -1757
rect 1696 -1758 1711 -1757
rect 110 -1760 255 -1759
rect 275 -1760 801 -1759
rect 814 -1760 843 -1759
rect 870 -1760 1060 -1759
rect 1080 -1760 1116 -1759
rect 1160 -1760 1214 -1759
rect 1374 -1760 1494 -1759
rect 1528 -1760 1641 -1759
rect 114 -1762 619 -1761
rect 667 -1762 766 -1761
rect 793 -1762 878 -1761
rect 887 -1762 1319 -1761
rect 1444 -1762 1494 -1761
rect 1528 -1762 1620 -1761
rect 1633 -1762 1697 -1761
rect 114 -1764 367 -1763
rect 408 -1764 486 -1763
rect 625 -1764 668 -1763
rect 677 -1764 773 -1763
rect 800 -1764 1046 -1763
rect 1073 -1764 1081 -1763
rect 1108 -1764 1200 -1763
rect 1276 -1764 1319 -1763
rect 1430 -1764 1445 -1763
rect 1563 -1764 1606 -1763
rect 149 -1766 1074 -1765
rect 1111 -1766 1669 -1765
rect 149 -1768 185 -1767
rect 191 -1768 437 -1767
rect 478 -1768 1781 -1767
rect 170 -1770 811 -1769
rect 821 -1770 871 -1769
rect 891 -1770 1480 -1769
rect 1549 -1770 1669 -1769
rect 180 -1772 423 -1771
rect 436 -1772 444 -1771
rect 625 -1772 727 -1771
rect 733 -1772 1480 -1771
rect 1584 -1772 1620 -1771
rect 180 -1774 1662 -1773
rect 184 -1776 549 -1775
rect 688 -1776 983 -1775
rect 989 -1776 1032 -1775
rect 1041 -1776 1270 -1775
rect 1279 -1776 1550 -1775
rect 1570 -1776 1662 -1775
rect 191 -1778 1655 -1777
rect 208 -1780 542 -1779
rect 548 -1780 1011 -1779
rect 1017 -1780 1214 -1779
rect 1234 -1780 1431 -1779
rect 1521 -1780 1585 -1779
rect 1591 -1780 1655 -1779
rect 233 -1782 342 -1781
rect 348 -1782 836 -1781
rect 849 -1782 892 -1781
rect 915 -1782 1389 -1781
rect 1507 -1782 1592 -1781
rect 233 -1784 433 -1783
rect 576 -1784 689 -1783
rect 695 -1784 787 -1783
rect 821 -1784 1284 -1783
rect 1381 -1784 1522 -1783
rect 1556 -1784 1571 -1783
rect 268 -1786 367 -1785
rect 411 -1786 804 -1785
rect 824 -1786 1634 -1785
rect 268 -1788 570 -1787
rect 576 -1788 895 -1787
rect 919 -1788 1725 -1787
rect 282 -1790 297 -1789
rect 317 -1790 479 -1789
rect 632 -1790 696 -1789
rect 702 -1790 1172 -1789
rect 1220 -1790 1235 -1789
rect 1269 -1790 1312 -1789
rect 1465 -1790 1508 -1789
rect 1703 -1790 1725 -1789
rect 156 -1792 1466 -1791
rect 1675 -1792 1704 -1791
rect 156 -1794 633 -1793
rect 639 -1794 703 -1793
rect 709 -1794 794 -1793
rect 828 -1794 1158 -1793
rect 1171 -1794 1805 -1793
rect 198 -1796 318 -1795
rect 324 -1796 395 -1795
rect 415 -1796 923 -1795
rect 926 -1796 1137 -1795
rect 1157 -1796 1417 -1795
rect 1675 -1796 1690 -1795
rect 198 -1798 514 -1797
rect 639 -1798 647 -1797
rect 709 -1798 1067 -1797
rect 1115 -1798 1165 -1797
rect 1178 -1798 1221 -1797
rect 1276 -1798 1690 -1797
rect 247 -1800 283 -1799
rect 289 -1800 1137 -1799
rect 1283 -1800 1291 -1799
rect 1416 -1800 1746 -1799
rect 121 -1802 290 -1801
rect 310 -1802 395 -1801
rect 422 -1802 675 -1801
rect 716 -1802 1011 -1801
rect 1017 -1802 1487 -1801
rect 1731 -1802 1746 -1801
rect 93 -1804 717 -1803
rect 737 -1804 1382 -1803
rect 1717 -1804 1732 -1803
rect 93 -1806 258 -1805
rect 303 -1806 738 -1805
rect 744 -1806 913 -1805
rect 919 -1806 1777 -1805
rect 79 -1808 304 -1807
rect 331 -1808 353 -1807
rect 359 -1808 486 -1807
rect 674 -1808 1109 -1807
rect 1153 -1808 1487 -1807
rect 79 -1810 381 -1809
rect 446 -1810 1557 -1809
rect 121 -1812 507 -1811
rect 744 -1812 752 -1811
rect 758 -1812 815 -1811
rect 828 -1812 1788 -1811
rect 135 -1814 759 -1813
rect 772 -1814 1802 -1813
rect 100 -1816 136 -1815
rect 205 -1816 311 -1815
rect 331 -1816 444 -1815
rect 464 -1816 514 -1815
rect 611 -1816 752 -1815
rect 789 -1816 1718 -1815
rect 100 -1818 227 -1817
rect 338 -1818 475 -1817
rect 506 -1818 556 -1817
rect 597 -1818 612 -1817
rect 849 -1818 1088 -1817
rect 1101 -1818 1179 -1817
rect 1290 -1818 1774 -1817
rect 86 -1820 556 -1819
rect 597 -1820 780 -1819
rect 863 -1820 1102 -1819
rect 1542 -1820 1774 -1819
rect 72 -1822 87 -1821
rect 205 -1822 1256 -1821
rect 1458 -1822 1543 -1821
rect 44 -1824 73 -1823
rect 212 -1824 780 -1823
rect 863 -1824 1263 -1823
rect 1423 -1824 1459 -1823
rect 44 -1826 164 -1825
rect 212 -1826 493 -1825
rect 912 -1826 955 -1825
rect 982 -1826 1242 -1825
rect 1339 -1826 1424 -1825
rect 163 -1828 832 -1827
rect 926 -1828 1578 -1827
rect 219 -1830 227 -1829
rect 338 -1830 468 -1829
rect 471 -1830 570 -1829
rect 831 -1830 1333 -1829
rect 1402 -1830 1578 -1829
rect 219 -1832 692 -1831
rect 929 -1832 1501 -1831
rect 359 -1834 374 -1833
rect 380 -1834 458 -1833
rect 492 -1834 528 -1833
rect 936 -1834 1151 -1833
rect 1206 -1834 1256 -1833
rect 1395 -1834 1403 -1833
rect 37 -1836 528 -1835
rect 947 -1836 1389 -1835
rect 37 -1838 52 -1837
rect 247 -1838 458 -1837
rect 898 -1838 948 -1837
rect 975 -1838 1151 -1837
rect 1206 -1838 1305 -1837
rect 1346 -1838 1396 -1837
rect 51 -1840 143 -1839
rect 373 -1840 563 -1839
rect 898 -1840 930 -1839
rect 933 -1840 1347 -1839
rect 142 -1842 178 -1841
rect 401 -1842 472 -1841
rect 562 -1842 650 -1841
rect 856 -1842 934 -1841
rect 996 -1842 1193 -1841
rect 1227 -1842 1263 -1841
rect 1297 -1842 1305 -1841
rect 429 -1844 465 -1843
rect 656 -1844 1228 -1843
rect 1251 -1844 1340 -1843
rect 681 -1846 857 -1845
rect 961 -1846 997 -1845
rect 1003 -1846 1032 -1845
rect 1038 -1846 1088 -1845
rect 1143 -1846 1242 -1845
rect 1297 -1846 1515 -1845
rect 345 -1848 1039 -1847
rect 1045 -1848 1564 -1847
rect 583 -1850 682 -1849
rect 835 -1850 1004 -1849
rect 1024 -1850 1165 -1849
rect 1353 -1850 1515 -1849
rect 583 -1852 591 -1851
rect 653 -1852 962 -1851
rect 968 -1852 1025 -1851
rect 1027 -1852 1599 -1851
rect 450 -1854 654 -1853
rect 968 -1854 986 -1853
rect 1048 -1854 1501 -1853
rect 590 -1856 661 -1855
rect 1066 -1856 1130 -1855
rect 1353 -1856 1473 -1855
rect 660 -1858 783 -1857
rect 905 -1858 1130 -1857
rect 1451 -1858 1473 -1857
rect 807 -1860 1452 -1859
rect 905 -1862 1438 -1861
rect 1094 -1864 1144 -1863
rect 1409 -1864 1438 -1863
rect 194 -1866 1410 -1865
rect 1094 -1868 1123 -1867
rect 1122 -1870 1186 -1869
rect 1185 -1872 1361 -1871
rect 1325 -1874 1361 -1873
rect 723 -1876 1326 -1875
rect 387 -1878 724 -1877
rect 387 -1880 521 -1879
rect 250 -1882 521 -1881
rect 51 -1893 216 -1892
rect 233 -1893 888 -1892
rect 905 -1893 1200 -1892
rect 1216 -1893 1228 -1892
rect 1276 -1893 1578 -1892
rect 1654 -1893 1805 -1892
rect 51 -1895 269 -1894
rect 303 -1895 475 -1894
rect 478 -1895 906 -1894
rect 919 -1895 983 -1894
rect 1017 -1895 1165 -1894
rect 1276 -1895 1417 -1894
rect 1773 -1895 1795 -1894
rect 68 -1897 549 -1896
rect 572 -1897 1347 -1896
rect 1381 -1897 1385 -1896
rect 1409 -1897 1777 -1896
rect 1794 -1897 1809 -1896
rect 72 -1899 108 -1898
rect 135 -1899 262 -1898
rect 303 -1899 563 -1898
rect 593 -1899 1452 -1898
rect 1493 -1899 1809 -1898
rect 72 -1901 150 -1900
rect 156 -1901 234 -1900
rect 250 -1901 549 -1900
rect 562 -1901 948 -1900
rect 954 -1901 969 -1900
rect 1024 -1901 1760 -1900
rect 79 -1903 339 -1902
rect 345 -1903 829 -1902
rect 831 -1903 1102 -1902
rect 1111 -1903 1725 -1902
rect 79 -1905 612 -1904
rect 646 -1905 780 -1904
rect 796 -1905 843 -1904
rect 849 -1905 1200 -1904
rect 1279 -1905 1725 -1904
rect 86 -1907 108 -1906
rect 135 -1907 402 -1906
rect 436 -1907 1000 -1906
rect 1024 -1907 1144 -1906
rect 1153 -1907 1732 -1906
rect 86 -1909 311 -1908
rect 324 -1909 468 -1908
rect 499 -1909 867 -1908
rect 922 -1909 986 -1908
rect 1031 -1909 1102 -1908
rect 1115 -1909 1228 -1908
rect 1314 -1909 1634 -1908
rect 1731 -1909 1753 -1908
rect 89 -1911 1165 -1910
rect 1353 -1911 1494 -1910
rect 1633 -1911 1648 -1910
rect 1752 -1911 1781 -1910
rect 100 -1913 447 -1912
rect 464 -1913 878 -1912
rect 926 -1913 997 -1912
rect 1003 -1913 1116 -1912
rect 1139 -1913 1774 -1912
rect 1780 -1913 1802 -1912
rect 100 -1915 1578 -1914
rect 1801 -1915 1816 -1914
rect 110 -1917 437 -1916
rect 509 -1917 1347 -1916
rect 1381 -1917 1508 -1916
rect 142 -1919 1655 -1918
rect 142 -1921 1557 -1920
rect 145 -1923 311 -1922
rect 324 -1923 395 -1922
rect 527 -1923 1690 -1922
rect 149 -1925 209 -1924
rect 212 -1925 444 -1924
rect 527 -1925 675 -1924
rect 723 -1925 948 -1924
rect 957 -1925 1319 -1924
rect 1409 -1925 1522 -1924
rect 1626 -1925 1690 -1924
rect 156 -1927 185 -1926
rect 191 -1927 269 -1926
rect 334 -1927 444 -1926
rect 541 -1927 612 -1926
rect 618 -1927 927 -1926
rect 929 -1927 1004 -1926
rect 1027 -1927 1648 -1926
rect 128 -1929 185 -1928
rect 191 -1929 416 -1928
rect 506 -1929 542 -1928
rect 597 -1929 780 -1928
rect 800 -1929 976 -1928
rect 1031 -1929 1081 -1928
rect 1143 -1929 1249 -1928
rect 1318 -1929 1361 -1928
rect 1374 -1929 1522 -1928
rect 1626 -1929 1676 -1928
rect 152 -1931 416 -1930
rect 457 -1931 598 -1930
rect 618 -1931 640 -1930
rect 653 -1931 1214 -1930
rect 1248 -1931 1263 -1930
rect 1360 -1931 1445 -1930
rect 1675 -1931 1711 -1930
rect 37 -1933 458 -1932
rect 506 -1933 1760 -1932
rect 159 -1935 864 -1934
rect 901 -1935 1557 -1934
rect 1710 -1935 1746 -1934
rect 163 -1937 248 -1936
rect 254 -1937 1049 -1936
rect 1059 -1937 1354 -1936
rect 1374 -1937 1396 -1936
rect 1423 -1937 1445 -1936
rect 163 -1939 342 -1938
rect 345 -1939 430 -1938
rect 632 -1939 647 -1938
rect 653 -1939 1042 -1938
rect 1045 -1939 1298 -1938
rect 1395 -1939 1501 -1938
rect 93 -1941 1501 -1940
rect 93 -1943 178 -1942
rect 198 -1943 430 -1942
rect 632 -1943 703 -1942
rect 793 -1943 801 -1942
rect 807 -1943 962 -1942
rect 968 -1943 1333 -1942
rect 1423 -1943 1515 -1942
rect 103 -1945 1333 -1944
rect 1437 -1945 1452 -1944
rect 1514 -1945 1536 -1944
rect 170 -1947 402 -1946
rect 460 -1947 703 -1946
rect 807 -1947 892 -1946
rect 933 -1947 941 -1946
rect 975 -1947 1340 -1946
rect 1402 -1947 1438 -1946
rect 1535 -1947 1564 -1946
rect 110 -1949 1403 -1948
rect 1563 -1949 1571 -1948
rect 170 -1951 227 -1950
rect 247 -1951 276 -1950
rect 373 -1951 377 -1950
rect 380 -1951 479 -1950
rect 639 -1951 822 -1950
rect 824 -1951 885 -1950
rect 891 -1951 1459 -1950
rect 114 -1953 822 -1952
rect 835 -1953 909 -1952
rect 1010 -1953 1046 -1952
rect 1080 -1953 1109 -1952
rect 1157 -1953 1186 -1952
rect 1206 -1953 1340 -1952
rect 1430 -1953 1459 -1952
rect 114 -1955 283 -1954
rect 373 -1955 493 -1954
rect 667 -1955 675 -1954
rect 719 -1955 1109 -1954
rect 1122 -1955 1431 -1954
rect 131 -1957 227 -1956
rect 254 -1957 535 -1956
rect 667 -1957 759 -1956
rect 786 -1957 941 -1956
rect 989 -1957 1011 -1956
rect 1020 -1957 1060 -1956
rect 1087 -1957 1123 -1956
rect 1129 -1957 1158 -1956
rect 1206 -1957 1242 -1956
rect 1262 -1957 1487 -1956
rect 177 -1959 895 -1958
rect 989 -1959 1585 -1958
rect 180 -1961 794 -1960
rect 814 -1961 843 -1960
rect 877 -1961 885 -1960
rect 1052 -1961 1186 -1960
rect 1241 -1961 1256 -1960
rect 1297 -1961 1326 -1960
rect 1486 -1961 1620 -1960
rect 180 -1963 423 -1962
rect 485 -1963 493 -1962
rect 534 -1963 556 -1962
rect 590 -1963 787 -1962
rect 810 -1963 1326 -1962
rect 1528 -1963 1585 -1962
rect 1619 -1963 1641 -1962
rect 58 -1965 556 -1964
rect 758 -1965 1067 -1964
rect 1073 -1965 1130 -1964
rect 1220 -1965 1256 -1964
rect 1311 -1965 1571 -1964
rect 1640 -1965 1683 -1964
rect 58 -1967 710 -1966
rect 814 -1967 857 -1966
rect 1052 -1967 1137 -1966
rect 1192 -1967 1221 -1966
rect 1269 -1967 1312 -1966
rect 1384 -1967 1508 -1966
rect 1528 -1967 1550 -1966
rect 1682 -1967 1718 -1966
rect 198 -1969 762 -1968
rect 838 -1969 1389 -1968
rect 1542 -1969 1550 -1968
rect 205 -1971 290 -1970
rect 387 -1971 465 -1970
rect 649 -1971 1718 -1970
rect 212 -1973 1599 -1972
rect 219 -1975 1088 -1974
rect 1178 -1975 1270 -1974
rect 1388 -1975 1473 -1974
rect 1598 -1975 1613 -1974
rect 219 -1977 381 -1976
rect 394 -1977 717 -1976
rect 856 -1977 871 -1976
rect 1017 -1977 1137 -1976
rect 1178 -1977 1368 -1976
rect 1465 -1977 1473 -1976
rect 1612 -1977 1662 -1976
rect 264 -1979 290 -1978
rect 422 -1979 731 -1978
rect 870 -1979 937 -1978
rect 1038 -1979 1543 -1978
rect 1661 -1979 1704 -1978
rect 275 -1981 360 -1980
rect 709 -1981 899 -1980
rect 1038 -1981 1697 -1980
rect 1703 -1981 1739 -1980
rect 282 -1983 472 -1982
rect 716 -1983 850 -1982
rect 1066 -1983 1291 -1982
rect 1293 -1983 1697 -1982
rect 1738 -1983 1767 -1982
rect 359 -1985 689 -1984
rect 723 -1985 899 -1984
rect 1073 -1985 1095 -1984
rect 1192 -1985 1417 -1984
rect 1465 -1985 1606 -1984
rect 1766 -1985 1788 -1984
rect 366 -1987 472 -1986
rect 583 -1987 1095 -1986
rect 1304 -1987 1368 -1986
rect 1591 -1987 1606 -1986
rect 317 -1989 367 -1988
rect 583 -1989 626 -1988
rect 628 -1989 1305 -1988
rect 317 -1991 409 -1990
rect 625 -1991 696 -1990
rect 730 -1991 1151 -1990
rect 1160 -1991 1592 -1990
rect 352 -1993 409 -1992
rect 576 -1993 696 -1992
rect 919 -1993 1788 -1992
rect 30 -1995 577 -1994
rect 681 -1995 689 -1994
rect 961 -1995 1151 -1994
rect 30 -1997 332 -1996
rect 681 -1997 766 -1996
rect 44 -1999 332 -1998
rect 744 -1999 766 -1998
rect 44 -2001 531 -2000
rect 660 -2001 745 -2000
rect 124 -2003 353 -2002
rect 520 -2003 661 -2002
rect 513 -2005 521 -2004
rect 450 -2007 514 -2006
rect 450 -2009 570 -2008
rect 121 -2011 570 -2010
rect 121 -2013 1480 -2012
rect 656 -2015 1480 -2014
rect 37 -2026 626 -2025
rect 667 -2026 671 -2025
rect 702 -2026 958 -2025
rect 964 -2026 1053 -2025
rect 1062 -2026 1081 -2025
rect 1139 -2026 1438 -2025
rect 1479 -2026 1749 -2025
rect 44 -2028 713 -2027
rect 719 -2028 927 -2027
rect 929 -2028 1431 -2027
rect 1591 -2028 1595 -2027
rect 1713 -2028 1795 -2027
rect 44 -2030 181 -2029
rect 222 -2030 248 -2029
rect 278 -2030 1165 -2029
rect 1195 -2030 1445 -2029
rect 1591 -2030 1606 -2029
rect 1745 -2030 1781 -2029
rect 51 -2032 178 -2031
rect 229 -2032 1200 -2031
rect 1213 -2032 1683 -2031
rect 51 -2034 276 -2033
rect 331 -2034 472 -2033
rect 516 -2034 941 -2033
rect 954 -2034 1340 -2033
rect 1423 -2034 1438 -2033
rect 1444 -2034 1522 -2033
rect 1682 -2034 1711 -2033
rect 61 -2036 1095 -2035
rect 1157 -2036 1480 -2035
rect 72 -2038 202 -2037
rect 240 -2038 251 -2037
rect 331 -2038 461 -2037
rect 464 -2038 507 -2037
rect 520 -2038 524 -2037
rect 555 -2038 587 -2037
rect 590 -2038 598 -2037
rect 614 -2038 976 -2037
rect 996 -2038 1340 -2037
rect 1395 -2038 1424 -2037
rect 1430 -2038 1515 -2037
rect 72 -2040 262 -2039
rect 338 -2040 594 -2039
rect 667 -2040 731 -2039
rect 751 -2040 895 -2039
rect 898 -2040 1298 -2039
rect 1314 -2040 1704 -2039
rect 100 -2042 423 -2041
rect 520 -2042 535 -2041
rect 558 -2042 1522 -2041
rect 1703 -2042 1725 -2041
rect 103 -2044 864 -2043
rect 877 -2044 962 -2043
rect 996 -2044 1179 -2043
rect 1195 -2044 1669 -2043
rect 1724 -2044 1788 -2043
rect 103 -2046 192 -2045
rect 205 -2046 465 -2045
rect 702 -2046 1452 -2045
rect 1514 -2046 1571 -2045
rect 1594 -2046 1606 -2045
rect 1626 -2046 1669 -2045
rect 110 -2048 150 -2047
rect 177 -2048 584 -2047
rect 751 -2048 773 -2047
rect 786 -2048 993 -2047
rect 999 -2048 1739 -2047
rect 114 -2050 598 -2049
rect 761 -2050 836 -2049
rect 856 -2050 864 -2049
rect 887 -2050 1620 -2049
rect 1626 -2050 1662 -2049
rect 1738 -2050 1809 -2049
rect 114 -2052 654 -2051
rect 786 -2052 885 -2051
rect 905 -2052 955 -2051
rect 999 -2052 1116 -2051
rect 1157 -2052 1172 -2051
rect 1199 -2052 1333 -2051
rect 1395 -2052 1410 -2051
rect 1451 -2052 1459 -2051
rect 1570 -2052 1578 -2051
rect 1619 -2052 1641 -2051
rect 1661 -2052 1760 -2051
rect 121 -2054 1501 -2053
rect 1507 -2054 1641 -2053
rect 121 -2056 458 -2055
rect 572 -2056 654 -2055
rect 695 -2056 885 -2055
rect 912 -2056 941 -2055
rect 1017 -2056 1039 -2055
rect 1052 -2056 1102 -2055
rect 1164 -2056 1249 -2055
rect 1293 -2056 1368 -2055
rect 1409 -2056 1417 -2055
rect 1458 -2056 1529 -2055
rect 1577 -2056 1599 -2055
rect 124 -2058 206 -2057
rect 219 -2058 1298 -2057
rect 1332 -2058 1389 -2057
rect 1500 -2058 1697 -2057
rect 124 -2060 311 -2059
rect 338 -2060 1109 -2059
rect 1171 -2060 1242 -2059
rect 1283 -2060 1368 -2059
rect 1507 -2060 1564 -2059
rect 1584 -2060 1599 -2059
rect 1689 -2060 1697 -2059
rect 131 -2062 563 -2061
rect 569 -2062 1249 -2061
rect 1283 -2062 1319 -2061
rect 1563 -2062 1613 -2061
rect 1689 -2062 1718 -2061
rect 131 -2064 1655 -2063
rect 135 -2066 276 -2065
rect 359 -2066 388 -2065
rect 394 -2066 804 -2065
rect 817 -2066 871 -2065
rect 873 -2066 1529 -2065
rect 1612 -2066 1648 -2065
rect 1654 -2066 1753 -2065
rect 30 -2068 136 -2067
rect 142 -2068 906 -2067
rect 912 -2068 948 -2067
rect 968 -2068 1109 -2067
rect 1241 -2068 1277 -2067
rect 1318 -2068 1382 -2067
rect 1647 -2068 1732 -2067
rect 30 -2070 97 -2069
rect 142 -2070 724 -2069
rect 793 -2070 829 -2069
rect 831 -2070 1256 -2069
rect 1381 -2070 1543 -2069
rect 1731 -2070 1802 -2069
rect 145 -2072 1004 -2071
rect 1024 -2072 1116 -2071
rect 1255 -2072 1312 -2071
rect 184 -2074 311 -2073
rect 317 -2074 360 -2073
rect 366 -2074 510 -2073
rect 548 -2074 1585 -2073
rect 184 -2076 213 -2075
rect 233 -2076 878 -2075
rect 922 -2076 1186 -2075
rect 1290 -2076 1543 -2075
rect 65 -2078 213 -2077
rect 240 -2078 293 -2077
rect 317 -2078 325 -2077
rect 366 -2078 486 -2077
rect 541 -2078 549 -2077
rect 628 -2078 724 -2077
rect 796 -2078 1214 -2077
rect 65 -2080 706 -2079
rect 709 -2080 1018 -2079
rect 1024 -2080 1144 -2079
rect 1185 -2080 1270 -2079
rect 86 -2082 234 -2081
rect 247 -2082 472 -2081
rect 541 -2082 822 -2081
rect 835 -2082 1028 -2081
rect 1073 -2082 1137 -2081
rect 1143 -2082 1305 -2081
rect 86 -2084 626 -2083
rect 695 -2084 738 -2083
rect 821 -2084 1473 -2083
rect 191 -2086 451 -2085
rect 457 -2086 605 -2085
rect 681 -2086 738 -2085
rect 856 -2086 892 -2085
rect 919 -2086 1291 -2085
rect 1304 -2086 1361 -2085
rect 1472 -2086 1494 -2085
rect 93 -2088 920 -2087
rect 933 -2088 969 -2087
rect 989 -2088 1277 -2087
rect 1493 -2088 1557 -2087
rect 93 -2090 1634 -2089
rect 163 -2092 605 -2091
rect 660 -2092 682 -2091
rect 807 -2092 934 -2091
rect 947 -2092 983 -2091
rect 1031 -2092 1074 -2091
rect 1080 -2092 1130 -2091
rect 1262 -2092 1361 -2091
rect 1486 -2092 1557 -2091
rect 1633 -2092 1676 -2091
rect 163 -2094 976 -2093
rect 978 -2094 1263 -2093
rect 1269 -2094 1326 -2093
rect 1675 -2094 1767 -2093
rect 198 -2096 388 -2095
rect 394 -2096 514 -2095
rect 555 -2096 990 -2095
rect 1010 -2096 1032 -2095
rect 1087 -2096 1417 -2095
rect 198 -2098 220 -2097
rect 254 -2098 563 -2097
rect 583 -2098 1487 -2097
rect 254 -2100 577 -2099
rect 807 -2100 850 -2099
rect 891 -2100 1133 -2099
rect 1325 -2100 1354 -2099
rect 156 -2102 577 -2101
rect 716 -2102 1354 -2101
rect 58 -2104 157 -2103
rect 268 -2104 423 -2103
rect 429 -2104 570 -2103
rect 716 -2104 1193 -2103
rect 226 -2106 269 -2105
rect 282 -2106 486 -2105
rect 814 -2106 850 -2105
rect 982 -2106 1060 -2105
rect 1087 -2106 1228 -2105
rect 226 -2108 1179 -2107
rect 1227 -2108 1711 -2107
rect 282 -2110 528 -2109
rect 1010 -2110 1375 -2109
rect 289 -2112 661 -2111
rect 1059 -2112 1389 -2111
rect 170 -2114 290 -2113
rect 324 -2114 374 -2113
rect 380 -2114 815 -2113
rect 1094 -2114 1123 -2113
rect 1129 -2114 1774 -2113
rect 170 -2116 479 -2115
rect 527 -2116 780 -2115
rect 1101 -2116 1151 -2115
rect 1374 -2116 1466 -2115
rect 107 -2118 1466 -2117
rect 107 -2120 689 -2119
rect 758 -2120 1151 -2119
rect 345 -2122 479 -2121
rect 499 -2122 689 -2121
rect 765 -2122 780 -2121
rect 345 -2124 444 -2123
rect 499 -2124 612 -2123
rect 765 -2124 801 -2123
rect 303 -2126 444 -2125
rect 492 -2126 612 -2125
rect 303 -2128 902 -2127
rect 352 -2130 759 -2129
rect 352 -2132 514 -2131
rect 373 -2134 1347 -2133
rect 128 -2136 1347 -2135
rect 128 -2138 262 -2137
rect 380 -2138 647 -2137
rect 401 -2140 493 -2139
rect 646 -2140 675 -2139
rect 79 -2142 402 -2141
rect 408 -2142 451 -2141
rect 674 -2142 1126 -2141
rect 79 -2144 416 -2143
rect 418 -2144 1004 -2143
rect 408 -2146 629 -2145
rect 429 -2148 1312 -2147
rect 436 -2150 773 -2149
rect 436 -2152 640 -2151
rect 618 -2154 640 -2153
rect 618 -2156 1046 -2155
rect 1045 -2158 1221 -2157
rect 1206 -2160 1221 -2159
rect 1206 -2162 1235 -2161
rect 1234 -2164 1403 -2163
rect 1402 -2166 1536 -2165
rect 1535 -2168 1550 -2167
rect 152 -2170 1550 -2169
rect 51 -2181 416 -2180
rect 418 -2181 801 -2180
rect 803 -2181 1690 -2180
rect 1696 -2181 1711 -2180
rect 58 -2183 136 -2182
rect 145 -2183 906 -2182
rect 940 -2183 1060 -2182
rect 1125 -2183 1424 -2182
rect 1640 -2183 1718 -2182
rect 72 -2185 629 -2184
rect 660 -2185 829 -2184
rect 866 -2185 1340 -2184
rect 1409 -2185 1413 -2184
rect 1650 -2185 1669 -2184
rect 1671 -2185 1739 -2184
rect 93 -2187 311 -2186
rect 317 -2187 377 -2186
rect 380 -2187 927 -2186
rect 943 -2187 1088 -2186
rect 1132 -2187 1683 -2186
rect 1689 -2187 1725 -2186
rect 93 -2189 1203 -2188
rect 1262 -2189 1683 -2188
rect 1696 -2189 1732 -2188
rect 100 -2191 1042 -2190
rect 1059 -2191 1067 -2190
rect 1087 -2191 1123 -2190
rect 1150 -2191 1340 -2190
rect 1388 -2191 1669 -2190
rect 61 -2193 101 -2192
rect 107 -2193 409 -2192
rect 492 -2193 584 -2192
rect 586 -2193 934 -2192
rect 975 -2193 1368 -2192
rect 1388 -2193 1445 -2192
rect 110 -2195 199 -2194
rect 201 -2195 423 -2194
rect 499 -2195 825 -2194
rect 873 -2195 1298 -2194
rect 1311 -2195 1508 -2194
rect 72 -2197 874 -2196
rect 877 -2197 927 -2196
rect 933 -2197 983 -2196
rect 999 -2197 1081 -2196
rect 1150 -2197 1721 -2196
rect 114 -2199 423 -2198
rect 499 -2199 507 -2198
rect 513 -2199 1123 -2198
rect 1174 -2199 1249 -2198
rect 1262 -2199 1354 -2198
rect 1409 -2199 1487 -2198
rect 1507 -2199 1543 -2198
rect 114 -2201 615 -2200
rect 618 -2201 671 -2200
rect 688 -2201 871 -2200
rect 877 -2201 1228 -2200
rect 1248 -2201 1270 -2200
rect 1311 -2201 1333 -2200
rect 1353 -2201 1466 -2200
rect 1542 -2201 1599 -2200
rect 121 -2203 458 -2202
rect 506 -2203 577 -2202
rect 583 -2203 591 -2202
rect 604 -2203 839 -2202
rect 905 -2203 962 -2202
rect 975 -2203 1039 -2202
rect 1066 -2203 1109 -2202
rect 1227 -2203 1417 -2202
rect 1444 -2203 1452 -2202
rect 1598 -2203 1634 -2202
rect 44 -2205 458 -2204
rect 495 -2205 591 -2204
rect 611 -2205 633 -2204
rect 660 -2205 913 -2204
rect 961 -2205 1004 -2204
rect 1020 -2205 1298 -2204
rect 1318 -2205 1368 -2204
rect 1374 -2205 1466 -2204
rect 44 -2207 97 -2206
rect 128 -2207 136 -2206
rect 156 -2207 409 -2206
rect 513 -2207 521 -2206
rect 534 -2207 559 -2206
rect 618 -2207 647 -2206
rect 688 -2207 808 -2206
rect 817 -2207 1641 -2206
rect 128 -2209 654 -2208
rect 691 -2209 724 -2208
rect 761 -2209 1018 -2208
rect 1027 -2209 1221 -2208
rect 1314 -2209 1375 -2208
rect 1381 -2209 1417 -2208
rect 131 -2211 150 -2210
rect 156 -2211 465 -2210
rect 520 -2211 570 -2210
rect 597 -2211 647 -2210
rect 698 -2211 787 -2210
rect 807 -2211 864 -2210
rect 978 -2211 1704 -2210
rect 65 -2213 864 -2212
rect 982 -2213 1053 -2212
rect 1062 -2213 1319 -2212
rect 1332 -2213 1431 -2212
rect 65 -2215 283 -2214
rect 285 -2215 1529 -2214
rect 124 -2217 1431 -2216
rect 1528 -2217 1627 -2216
rect 138 -2219 654 -2218
rect 709 -2219 1452 -2218
rect 1626 -2219 1676 -2218
rect 163 -2221 248 -2220
rect 254 -2221 339 -2220
rect 359 -2221 381 -2220
rect 394 -2221 580 -2220
rect 600 -2221 1053 -2220
rect 1080 -2221 1137 -2220
rect 1381 -2221 1396 -2220
rect 163 -2223 738 -2222
rect 786 -2223 850 -2222
rect 1003 -2223 1074 -2222
rect 1108 -2223 1196 -2222
rect 1395 -2223 1438 -2222
rect 170 -2225 416 -2224
rect 464 -2225 668 -2224
rect 674 -2225 850 -2224
rect 1017 -2225 1473 -2224
rect 30 -2227 171 -2226
rect 177 -2227 643 -2226
rect 667 -2227 920 -2226
rect 1024 -2227 1221 -2226
rect 1437 -2227 1557 -2226
rect 30 -2229 209 -2228
rect 212 -2229 290 -2228
rect 296 -2229 300 -2228
rect 303 -2229 703 -2228
rect 709 -2229 899 -2228
rect 1027 -2229 1165 -2228
rect 1556 -2229 1578 -2228
rect 177 -2231 696 -2230
rect 716 -2231 920 -2230
rect 1073 -2231 1179 -2230
rect 1577 -2231 1662 -2230
rect 215 -2233 1011 -2232
rect 1115 -2233 1634 -2232
rect 226 -2235 542 -2234
rect 555 -2235 640 -2234
rect 681 -2235 703 -2234
rect 737 -2235 1025 -2234
rect 1115 -2235 1158 -2234
rect 1178 -2235 1291 -2234
rect 1535 -2235 1662 -2234
rect 226 -2237 241 -2236
rect 261 -2237 374 -2236
rect 394 -2237 451 -2236
rect 509 -2237 717 -2236
rect 821 -2237 1424 -2236
rect 229 -2239 1473 -2238
rect 233 -2241 1137 -2240
rect 1143 -2241 1165 -2240
rect 1199 -2241 1291 -2240
rect 233 -2243 913 -2242
rect 989 -2243 1158 -2242
rect 1206 -2243 1536 -2242
rect 240 -2245 598 -2244
rect 625 -2245 1480 -2244
rect 261 -2247 1193 -2246
rect 1206 -2247 1242 -2246
rect 1479 -2247 1494 -2246
rect 268 -2249 276 -2248
rect 282 -2249 955 -2248
rect 989 -2249 1095 -2248
rect 1143 -2249 1186 -2248
rect 1241 -2249 1277 -2248
rect 1493 -2249 1571 -2248
rect 268 -2251 346 -2250
rect 359 -2251 832 -2250
rect 898 -2251 969 -2250
rect 996 -2251 1186 -2250
rect 1276 -2251 1459 -2250
rect 1570 -2251 1592 -2250
rect 79 -2253 346 -2252
rect 401 -2253 570 -2252
rect 628 -2253 1270 -2252
rect 1591 -2253 1613 -2252
rect 79 -2255 1522 -2254
rect 1605 -2255 1613 -2254
rect 103 -2257 1459 -2256
rect 1521 -2257 1585 -2256
rect 1605 -2257 1648 -2256
rect 250 -2259 402 -2258
rect 471 -2259 969 -2258
rect 996 -2259 1102 -2258
rect 1584 -2259 1620 -2258
rect 1647 -2259 1676 -2258
rect 296 -2261 430 -2260
rect 471 -2261 773 -2260
rect 821 -2261 857 -2260
rect 929 -2261 1193 -2260
rect 1619 -2261 1655 -2260
rect 257 -2263 773 -2262
rect 856 -2263 948 -2262
rect 954 -2263 1214 -2262
rect 1412 -2263 1487 -2262
rect 303 -2265 444 -2264
rect 534 -2265 731 -2264
rect 814 -2265 948 -2264
rect 1010 -2265 1714 -2264
rect 191 -2267 444 -2266
rect 541 -2267 843 -2266
rect 1094 -2267 1172 -2266
rect 1213 -2267 1256 -2266
rect 149 -2269 192 -2268
rect 310 -2269 332 -2268
rect 338 -2269 353 -2268
rect 548 -2269 556 -2268
rect 632 -2269 892 -2268
rect 1255 -2269 1347 -2268
rect 86 -2271 353 -2270
rect 681 -2271 752 -2270
rect 758 -2271 843 -2270
rect 1234 -2271 1347 -2270
rect 86 -2273 678 -2272
rect 705 -2273 1102 -2272
rect 1234 -2273 1326 -2272
rect 152 -2275 549 -2274
rect 730 -2275 780 -2274
rect 793 -2275 892 -2274
rect 1283 -2275 1326 -2274
rect 205 -2277 752 -2276
rect 814 -2277 885 -2276
rect 1283 -2277 1305 -2276
rect 317 -2279 367 -2278
rect 527 -2279 759 -2278
rect 884 -2279 1046 -2278
rect 1304 -2279 1361 -2278
rect 142 -2281 528 -2280
rect 604 -2281 780 -2280
rect 1031 -2281 1046 -2280
rect 1360 -2281 1403 -2280
rect 142 -2283 724 -2282
rect 744 -2283 794 -2282
rect 1031 -2283 1130 -2282
rect 1402 -2283 1501 -2282
rect 205 -2285 1130 -2284
rect 1500 -2285 1515 -2284
rect 324 -2287 517 -2286
rect 744 -2287 766 -2286
rect 324 -2289 486 -2288
rect 765 -2289 836 -2288
rect 331 -2291 437 -2290
rect 485 -2291 1039 -2290
rect 366 -2293 388 -2292
rect 436 -2293 563 -2292
rect 835 -2293 1515 -2292
rect 37 -2295 563 -2294
rect 387 -2297 479 -2296
rect 450 -2299 479 -2298
rect 30 -2310 150 -2309
rect 205 -2310 220 -2309
rect 254 -2310 524 -2309
rect 548 -2310 944 -2309
rect 971 -2310 1095 -2309
rect 1174 -2310 1494 -2309
rect 1622 -2310 1697 -2309
rect 51 -2312 360 -2311
rect 387 -2312 549 -2311
rect 576 -2312 829 -2311
rect 835 -2312 1452 -2311
rect 1493 -2312 1543 -2311
rect 1647 -2312 1690 -2311
rect 65 -2314 69 -2313
rect 79 -2314 563 -2313
rect 597 -2314 762 -2313
rect 779 -2314 1347 -2313
rect 1451 -2314 1655 -2313
rect 65 -2316 262 -2315
rect 285 -2316 311 -2315
rect 317 -2316 587 -2315
rect 625 -2316 752 -2315
rect 821 -2316 829 -2315
rect 859 -2316 1431 -2315
rect 1542 -2316 1585 -2315
rect 79 -2318 402 -2317
rect 415 -2318 601 -2317
rect 635 -2318 675 -2317
rect 677 -2318 731 -2317
rect 740 -2318 1634 -2317
rect 128 -2320 703 -2319
rect 705 -2320 808 -2319
rect 866 -2320 1249 -2319
rect 1251 -2320 1326 -2319
rect 1346 -2320 1375 -2319
rect 1430 -2320 1459 -2319
rect 1612 -2320 1634 -2319
rect 114 -2322 808 -2321
rect 873 -2322 1305 -2321
rect 1374 -2322 1396 -2321
rect 1444 -2322 1459 -2321
rect 1612 -2322 1641 -2321
rect 114 -2324 409 -2323
rect 450 -2324 1137 -2323
rect 1171 -2324 1655 -2323
rect 135 -2326 542 -2325
rect 562 -2326 892 -2325
rect 912 -2326 1291 -2325
rect 1444 -2326 1473 -2325
rect 149 -2328 1067 -2327
rect 1073 -2328 1137 -2327
rect 1164 -2328 1172 -2327
rect 1199 -2328 1536 -2327
rect 208 -2330 465 -2329
rect 492 -2330 1042 -2329
rect 1052 -2330 1095 -2329
rect 1129 -2330 1585 -2329
rect 215 -2332 325 -2331
rect 359 -2332 535 -2331
rect 541 -2332 570 -2331
rect 579 -2332 1053 -2331
rect 1073 -2332 1081 -2331
rect 1122 -2332 1130 -2331
rect 1157 -2332 1165 -2331
rect 1202 -2332 1382 -2331
rect 1472 -2332 1508 -2331
rect 1535 -2332 1592 -2331
rect 86 -2334 570 -2333
rect 590 -2334 626 -2333
rect 639 -2334 843 -2333
rect 891 -2334 899 -2333
rect 912 -2334 1294 -2333
rect 1591 -2334 1606 -2333
rect 72 -2336 591 -2335
rect 639 -2336 682 -2335
rect 684 -2336 822 -2335
rect 842 -2336 906 -2335
rect 915 -2336 1417 -2335
rect 1605 -2336 1672 -2335
rect 72 -2338 633 -2337
rect 667 -2338 857 -2337
rect 989 -2338 993 -2337
rect 1017 -2338 1109 -2337
rect 1122 -2338 1578 -2337
rect 86 -2340 230 -2339
rect 233 -2340 255 -2339
rect 261 -2340 276 -2339
rect 289 -2340 409 -2339
rect 436 -2340 493 -2339
rect 495 -2340 647 -2339
rect 681 -2340 1158 -2339
rect 1185 -2340 1508 -2339
rect 117 -2342 290 -2341
rect 296 -2342 577 -2341
rect 632 -2342 955 -2341
rect 975 -2342 1109 -2341
rect 1185 -2342 1368 -2341
rect 142 -2344 234 -2343
rect 247 -2344 325 -2343
rect 373 -2344 465 -2343
rect 478 -2344 906 -2343
rect 975 -2344 983 -2343
rect 989 -2344 1004 -2343
rect 1020 -2344 1060 -2343
rect 1206 -2344 1245 -2343
rect 1248 -2344 1627 -2343
rect 142 -2346 241 -2345
rect 247 -2346 332 -2345
rect 373 -2346 605 -2345
rect 688 -2346 787 -2345
rect 849 -2346 983 -2345
rect 1003 -2346 1032 -2345
rect 1038 -2346 1389 -2345
rect 1570 -2346 1627 -2345
rect 170 -2348 276 -2347
rect 282 -2348 955 -2347
rect 996 -2348 1032 -2347
rect 1045 -2348 1081 -2347
rect 1206 -2348 1364 -2347
rect 1367 -2348 1501 -2347
rect 170 -2350 192 -2349
rect 219 -2350 227 -2349
rect 240 -2350 367 -2349
rect 380 -2350 402 -2349
rect 422 -2350 647 -2349
rect 691 -2350 780 -2349
rect 786 -2350 1669 -2349
rect 184 -2352 192 -2351
rect 226 -2352 969 -2351
rect 1059 -2352 1228 -2351
rect 1237 -2352 1487 -2351
rect 184 -2354 486 -2353
rect 506 -2354 703 -2353
rect 709 -2354 1046 -2353
rect 1150 -2354 1228 -2353
rect 1241 -2354 1480 -2353
rect 1486 -2354 1651 -2353
rect 268 -2356 416 -2355
rect 422 -2356 458 -2355
rect 506 -2356 556 -2355
rect 604 -2356 612 -2355
rect 621 -2356 1501 -2355
rect 1650 -2356 1662 -2355
rect 268 -2358 836 -2357
rect 838 -2358 1571 -2357
rect 1661 -2358 1683 -2357
rect 282 -2360 1480 -2359
rect 296 -2362 339 -2361
rect 345 -2362 689 -2361
rect 695 -2362 878 -2361
rect 947 -2362 1039 -2361
rect 1150 -2362 1382 -2361
rect 1388 -2362 1410 -2361
rect 100 -2364 696 -2363
rect 709 -2364 794 -2363
rect 800 -2364 878 -2363
rect 947 -2364 962 -2363
rect 992 -2364 997 -2363
rect 1241 -2364 1298 -2363
rect 1318 -2364 1417 -2363
rect 100 -2366 815 -2365
rect 870 -2366 1298 -2365
rect 1318 -2366 1333 -2365
rect 1339 -2366 1410 -2365
rect 310 -2368 472 -2367
rect 509 -2368 514 -2367
rect 534 -2368 930 -2367
rect 1269 -2368 1326 -2367
rect 1332 -2368 1354 -2367
rect 58 -2370 514 -2369
rect 611 -2370 794 -2369
rect 870 -2370 1025 -2369
rect 1255 -2370 1270 -2369
rect 1283 -2370 1305 -2369
rect 1339 -2370 1361 -2369
rect 44 -2372 59 -2371
rect 317 -2372 671 -2371
rect 716 -2372 801 -2371
rect 926 -2372 962 -2371
rect 1234 -2372 1256 -2371
rect 1262 -2372 1284 -2371
rect 1290 -2372 1529 -2371
rect 44 -2374 783 -2373
rect 898 -2374 927 -2373
rect 1017 -2374 1235 -2373
rect 1353 -2374 1424 -2373
rect 1528 -2374 1550 -2373
rect 331 -2376 650 -2375
rect 653 -2376 1025 -2375
rect 1192 -2376 1424 -2375
rect 1549 -2376 1557 -2375
rect 107 -2378 654 -2377
rect 660 -2378 815 -2377
rect 1178 -2378 1193 -2377
rect 1213 -2378 1263 -2377
rect 1402 -2378 1557 -2377
rect 138 -2380 1179 -2379
rect 1213 -2380 1522 -2379
rect 163 -2382 661 -2381
rect 723 -2382 1067 -2381
rect 1276 -2382 1403 -2381
rect 1521 -2382 1564 -2381
rect 163 -2384 430 -2383
rect 436 -2384 521 -2383
rect 583 -2384 717 -2383
rect 723 -2384 1676 -2383
rect 338 -2386 353 -2385
rect 366 -2386 528 -2385
rect 730 -2386 885 -2385
rect 1202 -2386 1277 -2385
rect 1563 -2386 1599 -2385
rect 156 -2388 353 -2387
rect 380 -2388 1105 -2387
rect 1598 -2388 1620 -2387
rect 156 -2390 734 -2389
rect 747 -2390 1396 -2389
rect 345 -2392 584 -2391
rect 751 -2392 864 -2391
rect 387 -2394 395 -2393
rect 404 -2394 430 -2393
rect 443 -2394 479 -2393
rect 520 -2394 556 -2393
rect 744 -2394 864 -2393
rect 128 -2396 745 -2395
rect 758 -2396 885 -2395
rect 443 -2398 941 -2397
rect 450 -2400 1620 -2399
rect 453 -2402 738 -2401
rect 758 -2402 766 -2401
rect 775 -2402 1578 -2401
rect 394 -2404 738 -2403
rect 765 -2404 773 -2403
rect 933 -2404 941 -2403
rect 457 -2406 1011 -2405
rect 471 -2408 619 -2407
rect 642 -2408 934 -2407
rect 1010 -2408 1102 -2407
rect 121 -2410 619 -2409
rect 121 -2412 213 -2411
rect 527 -2412 773 -2411
rect 198 -2414 213 -2413
rect 93 -2416 199 -2415
rect 93 -2418 178 -2417
rect 152 -2420 178 -2419
rect 44 -2431 531 -2430
rect 562 -2431 1396 -2430
rect 1615 -2431 1634 -2430
rect 93 -2433 118 -2432
rect 121 -2433 776 -2432
rect 831 -2433 1214 -2432
rect 1234 -2433 1588 -2432
rect 1622 -2433 1662 -2432
rect 93 -2435 444 -2434
rect 471 -2435 615 -2434
rect 674 -2435 741 -2434
rect 747 -2435 1578 -2434
rect 1626 -2435 1644 -2434
rect 107 -2437 1515 -2436
rect 1577 -2437 1585 -2436
rect 107 -2439 111 -2438
rect 121 -2439 724 -2438
rect 737 -2439 1228 -2438
rect 1248 -2439 1606 -2438
rect 135 -2441 647 -2440
rect 674 -2441 1028 -2440
rect 1066 -2441 1123 -2440
rect 1185 -2441 1214 -2440
rect 1251 -2441 1410 -2440
rect 1549 -2441 1606 -2440
rect 135 -2443 458 -2442
rect 520 -2443 661 -2442
rect 681 -2443 864 -2442
rect 901 -2443 976 -2442
rect 989 -2443 1067 -2442
rect 1104 -2443 1263 -2442
rect 1290 -2443 1417 -2442
rect 1549 -2443 1571 -2442
rect 142 -2445 482 -2444
rect 572 -2445 717 -2444
rect 723 -2445 1189 -2444
rect 1199 -2445 1438 -2444
rect 142 -2447 388 -2446
rect 394 -2447 472 -2446
rect 569 -2447 717 -2446
rect 733 -2447 1571 -2446
rect 163 -2449 811 -2448
rect 821 -2449 990 -2448
rect 1013 -2449 1529 -2448
rect 163 -2451 391 -2450
rect 394 -2451 633 -2450
rect 639 -2451 647 -2450
rect 681 -2451 685 -2450
rect 688 -2451 804 -2450
rect 821 -2451 1406 -2450
rect 1493 -2451 1529 -2450
rect 170 -2453 258 -2452
rect 282 -2453 773 -2452
rect 835 -2453 1046 -2452
rect 1164 -2453 1200 -2452
rect 1220 -2453 1291 -2452
rect 1332 -2453 1396 -2452
rect 1486 -2453 1494 -2452
rect 51 -2455 171 -2454
rect 219 -2455 227 -2454
rect 229 -2455 1651 -2454
rect 51 -2457 402 -2456
rect 404 -2457 430 -2456
rect 583 -2457 1487 -2456
rect 114 -2459 220 -2458
rect 240 -2459 430 -2458
rect 583 -2459 710 -2458
rect 740 -2459 843 -2458
rect 849 -2459 1298 -2458
rect 1339 -2459 1410 -2458
rect 58 -2461 115 -2460
rect 128 -2461 836 -2460
rect 849 -2461 878 -2460
rect 919 -2461 1326 -2460
rect 1346 -2461 1417 -2460
rect 58 -2463 286 -2462
rect 303 -2463 731 -2462
rect 758 -2463 773 -2462
rect 828 -2463 843 -2462
rect 852 -2463 1109 -2462
rect 1192 -2463 1298 -2462
rect 1318 -2463 1326 -2462
rect 1353 -2463 1438 -2462
rect 79 -2465 759 -2464
rect 856 -2465 1515 -2464
rect 79 -2467 248 -2466
rect 254 -2467 283 -2466
rect 303 -2467 1126 -2466
rect 1143 -2467 1193 -2466
rect 1206 -2467 1340 -2466
rect 1360 -2467 1564 -2466
rect 247 -2469 479 -2468
rect 576 -2469 731 -2468
rect 793 -2469 857 -2468
rect 929 -2469 1403 -2468
rect 1563 -2469 1613 -2468
rect 254 -2471 860 -2470
rect 933 -2471 1109 -2470
rect 1171 -2471 1361 -2470
rect 1374 -2471 1382 -2470
rect 1384 -2471 1592 -2470
rect 338 -2473 458 -2472
rect 523 -2473 577 -2472
rect 586 -2473 1228 -2472
rect 1241 -2473 1347 -2472
rect 324 -2475 339 -2474
rect 359 -2475 479 -2474
rect 600 -2475 962 -2474
rect 1024 -2475 1102 -2474
rect 1150 -2475 1172 -2474
rect 1202 -2475 1242 -2474
rect 1251 -2475 1263 -2474
rect 1269 -2475 1319 -2474
rect 233 -2477 325 -2476
rect 359 -2477 465 -2476
rect 604 -2477 661 -2476
rect 667 -2477 878 -2476
rect 905 -2477 962 -2476
rect 1024 -2477 1508 -2476
rect 233 -2479 374 -2478
rect 380 -2479 864 -2478
rect 898 -2479 906 -2478
rect 947 -2479 976 -2478
rect 1038 -2479 1186 -2478
rect 1206 -2479 1641 -2478
rect 296 -2481 374 -2480
rect 380 -2481 703 -2480
rect 709 -2481 766 -2480
rect 793 -2481 801 -2480
rect 828 -2481 1382 -2480
rect 1507 -2481 1536 -2480
rect 1640 -2481 1655 -2480
rect 173 -2483 297 -2482
rect 366 -2483 563 -2482
rect 618 -2483 920 -2482
rect 947 -2483 1095 -2482
rect 1178 -2483 1270 -2482
rect 1276 -2483 1592 -2482
rect 366 -2485 500 -2484
rect 618 -2485 626 -2484
rect 639 -2485 839 -2484
rect 891 -2485 1277 -2484
rect 1283 -2485 1333 -2484
rect 1535 -2485 1557 -2484
rect 401 -2487 437 -2486
rect 464 -2487 654 -2486
rect 695 -2487 934 -2486
rect 996 -2487 1039 -2486
rect 1045 -2487 1088 -2486
rect 1129 -2487 1179 -2486
rect 1220 -2487 1238 -2486
rect 1304 -2487 1354 -2486
rect 1556 -2487 1599 -2486
rect 128 -2489 997 -2488
rect 1052 -2489 1151 -2488
rect 1304 -2489 1312 -2488
rect 1458 -2489 1599 -2488
rect 408 -2491 444 -2490
rect 485 -2491 605 -2490
rect 621 -2491 689 -2490
rect 702 -2491 808 -2490
rect 870 -2491 892 -2490
rect 926 -2491 1095 -2490
rect 1146 -2491 1459 -2490
rect 65 -2493 486 -2492
rect 499 -2493 542 -2492
rect 569 -2493 1130 -2492
rect 1255 -2493 1312 -2492
rect 65 -2495 1620 -2494
rect 310 -2497 409 -2496
rect 436 -2497 451 -2496
rect 513 -2497 696 -2496
rect 737 -2497 1613 -2496
rect 198 -2499 311 -2498
rect 352 -2499 542 -2498
rect 611 -2499 1256 -2498
rect 89 -2501 353 -2500
rect 450 -2501 566 -2500
rect 625 -2501 913 -2500
rect 1052 -2501 1081 -2500
rect 198 -2503 206 -2502
rect 492 -2503 514 -2502
rect 527 -2503 1284 -2502
rect 205 -2505 213 -2504
rect 345 -2505 528 -2504
rect 548 -2505 612 -2504
rect 649 -2505 1375 -2504
rect 212 -2507 276 -2506
rect 289 -2507 346 -2506
rect 492 -2507 787 -2506
rect 800 -2507 1452 -2506
rect 240 -2509 290 -2508
rect 548 -2509 598 -2508
rect 653 -2509 780 -2508
rect 807 -2509 1543 -2508
rect 275 -2511 423 -2510
rect 506 -2511 598 -2510
rect 744 -2511 1088 -2510
rect 1367 -2511 1452 -2510
rect 1521 -2511 1543 -2510
rect 86 -2513 507 -2512
rect 565 -2513 633 -2512
rect 765 -2513 1648 -2512
rect 86 -2515 521 -2514
rect 779 -2515 1364 -2514
rect 1479 -2515 1522 -2514
rect 156 -2517 423 -2516
rect 814 -2517 871 -2516
rect 884 -2517 927 -2516
rect 1010 -2517 1081 -2516
rect 1157 -2517 1368 -2516
rect 1472 -2517 1480 -2516
rect 100 -2519 157 -2518
rect 268 -2519 815 -2518
rect 884 -2519 1004 -2518
rect 1073 -2519 1165 -2518
rect 1465 -2519 1473 -2518
rect 100 -2521 332 -2520
rect 534 -2521 1011 -2520
rect 1073 -2521 1137 -2520
rect 1430 -2521 1466 -2520
rect 72 -2523 535 -2522
rect 786 -2523 1158 -2522
rect 1423 -2523 1431 -2522
rect 72 -2525 262 -2524
rect 331 -2525 416 -2524
rect 912 -2525 955 -2524
rect 968 -2525 1004 -2524
rect 1388 -2525 1424 -2524
rect 149 -2527 1137 -2526
rect 149 -2529 192 -2528
rect 261 -2529 318 -2528
rect 555 -2529 1389 -2528
rect 184 -2531 269 -2530
rect 278 -2531 556 -2530
rect 751 -2531 955 -2530
rect 968 -2531 983 -2530
rect 177 -2533 185 -2532
rect 191 -2533 745 -2532
rect 982 -2533 1018 -2532
rect 177 -2535 216 -2534
rect 317 -2535 388 -2534
rect 1017 -2535 1060 -2534
rect 1031 -2537 1060 -2536
rect 971 -2539 1032 -2538
rect 44 -2550 304 -2549
rect 387 -2550 640 -2549
rect 656 -2550 1550 -2549
rect 1556 -2550 1560 -2549
rect 1584 -2550 1606 -2549
rect 1629 -2550 1641 -2549
rect 72 -2552 293 -2551
rect 303 -2552 426 -2551
rect 457 -2552 479 -2551
rect 527 -2552 682 -2551
rect 730 -2552 1466 -2551
rect 1472 -2552 1550 -2551
rect 1556 -2552 1613 -2551
rect 72 -2554 619 -2553
rect 625 -2554 808 -2553
rect 849 -2554 899 -2553
rect 950 -2554 1480 -2553
rect 1514 -2554 1585 -2553
rect 1591 -2554 1620 -2553
rect 86 -2556 181 -2555
rect 212 -2556 297 -2555
rect 352 -2556 682 -2555
rect 737 -2556 1487 -2555
rect 1559 -2556 1613 -2555
rect 86 -2558 647 -2557
rect 737 -2558 902 -2557
rect 971 -2558 1123 -2557
rect 1143 -2558 1326 -2557
rect 1405 -2558 1543 -2557
rect 1598 -2558 1627 -2557
rect 93 -2560 213 -2559
rect 233 -2560 668 -2559
rect 744 -2560 1102 -2559
rect 1136 -2560 1144 -2559
rect 1188 -2560 1431 -2559
rect 1444 -2560 1480 -2559
rect 1507 -2560 1543 -2559
rect 1577 -2560 1599 -2559
rect 93 -2562 531 -2561
rect 534 -2562 748 -2561
rect 789 -2562 1277 -2561
rect 1304 -2562 1403 -2561
rect 1409 -2562 1487 -2561
rect 121 -2564 832 -2563
rect 835 -2564 850 -2563
rect 887 -2564 1298 -2563
rect 1304 -2564 1438 -2563
rect 1458 -2564 1515 -2563
rect 65 -2566 122 -2565
rect 135 -2566 829 -2565
rect 901 -2566 1067 -2565
rect 1073 -2566 1466 -2565
rect 65 -2568 101 -2567
rect 135 -2568 178 -2567
rect 201 -2568 1445 -2567
rect 100 -2570 108 -2569
rect 142 -2570 416 -2569
rect 422 -2570 647 -2569
rect 667 -2570 717 -2569
rect 730 -2570 745 -2569
rect 758 -2570 836 -2569
rect 954 -2570 1326 -2569
rect 1388 -2570 1438 -2569
rect 107 -2572 132 -2571
rect 142 -2572 206 -2571
rect 215 -2572 423 -2571
rect 450 -2572 1123 -2571
rect 1129 -2572 1137 -2571
rect 1234 -2572 1592 -2571
rect 152 -2574 1508 -2573
rect 163 -2576 237 -2575
rect 254 -2576 962 -2575
rect 978 -2576 1284 -2575
rect 1346 -2576 1389 -2575
rect 1409 -2576 1571 -2575
rect 226 -2578 255 -2577
rect 275 -2578 759 -2577
rect 803 -2578 1361 -2577
rect 1423 -2578 1459 -2577
rect 198 -2580 227 -2579
rect 268 -2580 276 -2579
rect 278 -2580 689 -2579
rect 828 -2580 878 -2579
rect 926 -2580 955 -2579
rect 961 -2580 1060 -2579
rect 1066 -2580 1088 -2579
rect 1090 -2580 1536 -2579
rect 268 -2582 377 -2581
rect 380 -2582 535 -2581
rect 562 -2582 591 -2581
rect 597 -2582 1578 -2581
rect 247 -2584 591 -2583
rect 600 -2584 1473 -2583
rect 247 -2586 311 -2585
rect 317 -2586 353 -2585
rect 390 -2586 409 -2585
rect 450 -2586 958 -2585
rect 996 -2586 1564 -2585
rect 89 -2588 1564 -2587
rect 191 -2590 311 -2589
rect 345 -2590 381 -2589
rect 394 -2590 416 -2589
rect 457 -2590 486 -2589
rect 492 -2590 619 -2589
rect 625 -2590 710 -2589
rect 880 -2590 997 -2589
rect 1017 -2590 1298 -2589
rect 1318 -2590 1361 -2589
rect 1374 -2590 1424 -2589
rect 58 -2592 192 -2591
rect 282 -2592 444 -2591
rect 464 -2592 563 -2591
rect 565 -2592 1536 -2591
rect 58 -2594 325 -2593
rect 345 -2594 374 -2593
rect 401 -2594 409 -2593
rect 464 -2594 822 -2593
rect 905 -2594 1060 -2593
rect 1073 -2594 1228 -2593
rect 1251 -2594 1529 -2593
rect 233 -2596 325 -2595
rect 401 -2596 542 -2595
rect 555 -2596 710 -2595
rect 786 -2596 1018 -2595
rect 1024 -2596 1522 -2595
rect 257 -2598 444 -2597
rect 481 -2598 493 -2597
rect 502 -2598 598 -2597
rect 611 -2598 640 -2597
rect 688 -2598 815 -2597
rect 821 -2598 892 -2597
rect 905 -2598 976 -2597
rect 1027 -2598 1340 -2597
rect 1493 -2598 1522 -2597
rect 156 -2600 612 -2599
rect 614 -2600 1284 -2599
rect 1339 -2600 1616 -2599
rect 156 -2602 206 -2601
rect 261 -2602 283 -2601
rect 289 -2602 318 -2601
rect 485 -2602 675 -2601
rect 786 -2602 794 -2601
rect 814 -2602 843 -2601
rect 877 -2602 892 -2601
rect 912 -2602 927 -2601
rect 1038 -2602 1102 -2601
rect 1129 -2602 1263 -2601
rect 1269 -2602 1319 -2601
rect 1416 -2602 1494 -2601
rect 1500 -2602 1529 -2601
rect 163 -2604 976 -2603
rect 1038 -2604 1116 -2603
rect 1178 -2604 1375 -2603
rect 1451 -2604 1501 -2603
rect 240 -2606 843 -2605
rect 912 -2606 934 -2605
rect 1045 -2606 1431 -2605
rect 219 -2608 241 -2607
rect 261 -2608 605 -2607
rect 733 -2608 1179 -2607
rect 1220 -2608 1263 -2607
rect 1269 -2608 1637 -2607
rect 219 -2610 265 -2609
rect 289 -2610 339 -2609
rect 520 -2610 675 -2609
rect 733 -2610 1242 -2609
rect 1255 -2610 1347 -2609
rect 1367 -2610 1417 -2609
rect 338 -2612 500 -2611
rect 520 -2612 545 -2611
rect 555 -2612 570 -2611
rect 572 -2612 661 -2611
rect 793 -2612 1011 -2611
rect 1052 -2612 1147 -2611
rect 1171 -2612 1221 -2611
rect 1227 -2612 1249 -2611
rect 1276 -2612 1588 -2611
rect 499 -2614 542 -2613
rect 569 -2614 724 -2613
rect 800 -2614 1046 -2613
rect 1087 -2614 1235 -2613
rect 1241 -2614 1382 -2613
rect 1395 -2614 1452 -2613
rect 471 -2616 724 -2615
rect 863 -2616 1249 -2615
rect 1332 -2616 1368 -2615
rect 359 -2618 472 -2617
rect 583 -2618 755 -2617
rect 863 -2618 871 -2617
rect 884 -2618 934 -2617
rect 940 -2618 1011 -2617
rect 1031 -2618 1053 -2617
rect 1108 -2618 1172 -2617
rect 1213 -2618 1256 -2617
rect 1290 -2618 1333 -2617
rect 1353 -2618 1396 -2617
rect 208 -2620 1109 -2619
rect 1115 -2620 1200 -2619
rect 1311 -2620 1354 -2619
rect 359 -2622 419 -2621
rect 583 -2622 654 -2621
rect 660 -2622 948 -2621
rect 1031 -2622 1207 -2621
rect 331 -2624 654 -2623
rect 670 -2624 1382 -2623
rect 79 -2626 332 -2625
rect 604 -2626 703 -2625
rect 740 -2626 1207 -2625
rect 79 -2628 129 -2627
rect 702 -2628 990 -2627
rect 1080 -2628 1214 -2627
rect 803 -2630 1291 -2629
rect 810 -2632 948 -2631
rect 989 -2632 1004 -2631
rect 1164 -2632 1200 -2631
rect 856 -2634 871 -2633
rect 884 -2634 1095 -2633
rect 1157 -2634 1165 -2633
rect 1192 -2634 1312 -2633
rect 170 -2636 1095 -2635
rect 1150 -2636 1158 -2635
rect 170 -2638 185 -2637
rect 751 -2638 1193 -2637
rect 184 -2640 720 -2639
rect 859 -2640 1081 -2639
rect 1150 -2640 1606 -2639
rect 506 -2642 752 -2641
rect 919 -2642 941 -2641
rect 982 -2642 1004 -2641
rect 506 -2644 549 -2643
rect 919 -2644 1154 -2643
rect 436 -2646 549 -2645
rect 968 -2646 983 -2645
rect 436 -2648 514 -2647
rect 968 -2648 1186 -2647
rect 513 -2650 577 -2649
rect 1185 -2650 1571 -2649
rect 576 -2652 766 -2651
rect 765 -2654 773 -2653
rect 695 -2656 773 -2655
rect 695 -2658 780 -2657
rect 51 -2660 780 -2659
rect 51 -2662 150 -2661
rect 114 -2664 150 -2663
rect 114 -2666 367 -2665
rect 366 -2668 899 -2667
rect 44 -2679 748 -2678
rect 782 -2679 1585 -2678
rect 44 -2681 395 -2680
rect 397 -2681 430 -2680
rect 436 -2681 500 -2680
rect 534 -2681 647 -2680
rect 649 -2681 773 -2680
rect 786 -2681 885 -2680
rect 908 -2681 1298 -2680
rect 1524 -2681 1599 -2680
rect 51 -2683 202 -2682
rect 205 -2683 346 -2682
rect 394 -2683 1189 -2682
rect 1262 -2683 1301 -2682
rect 58 -2685 237 -2684
rect 264 -2685 1284 -2684
rect 58 -2687 129 -2686
rect 135 -2687 178 -2686
rect 198 -2687 311 -2686
rect 331 -2687 430 -2686
rect 446 -2687 1508 -2686
rect 72 -2689 678 -2688
rect 681 -2689 773 -2688
rect 786 -2689 1466 -2688
rect 1507 -2689 1606 -2688
rect 72 -2691 171 -2690
rect 177 -2691 444 -2690
rect 499 -2691 794 -2690
rect 800 -2691 1172 -2690
rect 1185 -2691 1550 -2690
rect 79 -2693 374 -2692
rect 408 -2693 423 -2692
rect 534 -2693 808 -2692
rect 817 -2693 1487 -2692
rect 79 -2695 766 -2694
rect 793 -2695 815 -2694
rect 877 -2695 1011 -2694
rect 1024 -2695 1466 -2694
rect 1486 -2695 1578 -2694
rect 86 -2697 566 -2696
rect 576 -2697 717 -2696
rect 730 -2697 1154 -2696
rect 1185 -2697 1340 -2696
rect 86 -2699 101 -2698
rect 114 -2699 332 -2698
rect 345 -2699 353 -2698
rect 373 -2699 416 -2698
rect 422 -2699 542 -2698
rect 576 -2699 696 -2698
rect 709 -2699 734 -2698
rect 737 -2699 899 -2698
rect 940 -2699 951 -2698
rect 957 -2699 1312 -2698
rect 65 -2701 115 -2700
rect 124 -2701 199 -2700
rect 205 -2701 241 -2700
rect 264 -2701 297 -2700
rect 310 -2701 612 -2700
rect 653 -2701 801 -2700
rect 845 -2701 899 -2700
rect 933 -2701 941 -2700
rect 968 -2701 997 -2700
rect 1010 -2701 1627 -2700
rect 65 -2703 153 -2702
rect 156 -2703 619 -2702
rect 653 -2703 1144 -2702
rect 1150 -2703 1613 -2702
rect 93 -2705 160 -2704
rect 170 -2705 451 -2704
rect 464 -2705 542 -2704
rect 569 -2705 619 -2704
rect 656 -2705 1053 -2704
rect 1073 -2705 1172 -2704
rect 1241 -2705 1340 -2704
rect 93 -2707 248 -2706
rect 296 -2707 472 -2706
rect 520 -2707 878 -2706
rect 880 -2707 1375 -2706
rect 100 -2709 209 -2708
rect 212 -2709 248 -2708
rect 352 -2709 402 -2708
rect 415 -2709 556 -2708
rect 569 -2709 591 -2708
rect 604 -2709 738 -2708
rect 744 -2709 762 -2708
rect 765 -2709 822 -2708
rect 880 -2709 1102 -2708
rect 1150 -2709 1382 -2708
rect 128 -2711 437 -2710
rect 450 -2711 507 -2710
rect 555 -2711 724 -2710
rect 744 -2711 1431 -2710
rect 135 -2713 640 -2712
rect 660 -2713 1091 -2712
rect 1101 -2713 1207 -2712
rect 1241 -2713 1354 -2712
rect 1381 -2713 1543 -2712
rect 142 -2715 262 -2714
rect 401 -2715 493 -2714
rect 506 -2715 668 -2714
rect 674 -2715 815 -2714
rect 821 -2715 850 -2714
rect 884 -2715 948 -2714
rect 954 -2715 1144 -2714
rect 1188 -2715 1375 -2714
rect 1430 -2715 1515 -2714
rect 142 -2717 290 -2716
rect 425 -2717 605 -2716
rect 611 -2717 920 -2716
rect 926 -2717 1053 -2716
rect 1087 -2717 1179 -2716
rect 1262 -2717 1368 -2716
rect 1514 -2717 1620 -2716
rect 149 -2719 857 -2718
rect 870 -2719 920 -2718
rect 933 -2719 983 -2718
rect 996 -2719 1004 -2718
rect 1024 -2719 1109 -2718
rect 1129 -2719 1207 -2718
rect 1283 -2719 1452 -2718
rect 149 -2721 269 -2720
rect 464 -2721 598 -2720
rect 625 -2721 724 -2720
rect 779 -2721 1074 -2720
rect 1108 -2721 1193 -2720
rect 1311 -2721 1396 -2720
rect 1451 -2721 1529 -2720
rect 156 -2723 1270 -2722
rect 1353 -2723 1445 -2722
rect 163 -2725 269 -2724
rect 387 -2725 598 -2724
rect 660 -2725 1592 -2724
rect 163 -2727 220 -2726
rect 226 -2727 241 -2726
rect 387 -2727 549 -2726
rect 562 -2727 640 -2726
rect 663 -2727 871 -2726
rect 901 -2727 1270 -2726
rect 1367 -2727 1459 -2726
rect 138 -2729 1459 -2728
rect 215 -2731 255 -2730
rect 408 -2731 563 -2730
rect 681 -2731 752 -2730
rect 849 -2731 990 -2730
rect 1115 -2731 1130 -2730
rect 1192 -2731 1424 -2730
rect 1444 -2731 1630 -2730
rect 219 -2733 304 -2732
rect 366 -2733 752 -2732
rect 856 -2733 864 -2732
rect 905 -2733 1179 -2732
rect 1395 -2733 1473 -2732
rect 226 -2735 234 -2734
rect 254 -2735 283 -2734
rect 303 -2735 339 -2734
rect 471 -2735 486 -2734
rect 492 -2735 615 -2734
rect 691 -2735 1081 -2734
rect 1115 -2735 1228 -2734
rect 1472 -2735 1557 -2734
rect 212 -2737 486 -2736
rect 527 -2737 626 -2736
rect 695 -2737 1095 -2736
rect 1227 -2737 1326 -2736
rect 324 -2739 367 -2738
rect 478 -2739 521 -2738
rect 527 -2739 633 -2738
rect 702 -2739 927 -2738
rect 954 -2739 1137 -2738
rect 1255 -2739 1326 -2738
rect 292 -2741 479 -2740
rect 548 -2741 843 -2740
rect 859 -2741 1424 -2740
rect 324 -2743 514 -2742
rect 583 -2743 633 -2742
rect 702 -2743 759 -2742
rect 842 -2743 1060 -2742
rect 1080 -2743 1158 -2742
rect 1255 -2743 1361 -2742
rect 338 -2745 360 -2744
rect 457 -2745 514 -2744
rect 583 -2745 689 -2744
rect 709 -2745 836 -2744
rect 863 -2745 1158 -2744
rect 1160 -2745 1361 -2744
rect 184 -2747 360 -2746
rect 380 -2747 458 -2746
rect 758 -2747 1347 -2746
rect 184 -2749 804 -2748
rect 828 -2749 836 -2748
rect 891 -2749 906 -2748
rect 961 -2749 983 -2748
rect 989 -2749 1018 -2748
rect 1059 -2749 1221 -2748
rect 1346 -2749 1438 -2748
rect 121 -2751 892 -2750
rect 971 -2751 1039 -2750
rect 1094 -2751 1165 -2750
rect 1220 -2751 1637 -2750
rect 121 -2753 132 -2752
rect 317 -2753 381 -2752
rect 779 -2753 962 -2752
rect 975 -2753 1046 -2752
rect 1136 -2753 1235 -2752
rect 1437 -2753 1522 -2752
rect 107 -2755 132 -2754
rect 191 -2755 318 -2754
rect 828 -2755 913 -2754
rect 947 -2755 1522 -2754
rect 107 -2757 192 -2756
rect 289 -2757 976 -2756
rect 978 -2757 1494 -2756
rect 667 -2759 913 -2758
rect 1017 -2759 1032 -2758
rect 1038 -2759 1123 -2758
rect 1164 -2759 1249 -2758
rect 1493 -2759 1571 -2758
rect 1031 -2761 1067 -2760
rect 1122 -2761 1277 -2760
rect 1045 -2763 1214 -2762
rect 1234 -2763 1333 -2762
rect 1066 -2765 1200 -2764
rect 1213 -2765 1319 -2764
rect 1332 -2765 1410 -2764
rect 1199 -2767 1291 -2766
rect 1318 -2767 1417 -2766
rect 887 -2769 1417 -2768
rect 1248 -2771 1634 -2770
rect 1276 -2773 1389 -2772
rect 1409 -2773 1501 -2772
rect 1290 -2775 1536 -2774
rect 1304 -2777 1389 -2776
rect 1402 -2777 1501 -2776
rect 674 -2779 1305 -2778
rect 1402 -2779 1480 -2778
rect 1479 -2781 1564 -2780
rect 58 -2792 237 -2791
rect 247 -2792 293 -2791
rect 303 -2792 559 -2791
rect 593 -2792 731 -2791
rect 747 -2792 1144 -2791
rect 1160 -2792 1501 -2791
rect 65 -2794 139 -2793
rect 149 -2794 283 -2793
rect 285 -2794 367 -2793
rect 380 -2794 447 -2793
rect 499 -2794 790 -2793
rect 810 -2794 1480 -2793
rect 86 -2796 108 -2795
rect 110 -2796 829 -2795
rect 845 -2796 997 -2795
rect 1006 -2796 1326 -2795
rect 86 -2798 318 -2797
rect 324 -2798 706 -2797
rect 730 -2798 738 -2797
rect 772 -2798 923 -2797
rect 996 -2798 1137 -2797
rect 1297 -2798 1382 -2797
rect 93 -2800 839 -2799
rect 866 -2800 1487 -2799
rect 93 -2802 185 -2801
rect 198 -2802 293 -2801
rect 310 -2802 325 -2801
rect 331 -2802 496 -2801
rect 499 -2802 671 -2801
rect 688 -2802 724 -2801
rect 737 -2802 752 -2801
rect 772 -2802 885 -2801
rect 898 -2802 1186 -2801
rect 1297 -2802 1396 -2801
rect 107 -2804 353 -2803
rect 366 -2804 423 -2803
rect 429 -2804 661 -2803
rect 688 -2804 1151 -2803
rect 1185 -2804 1256 -2803
rect 1325 -2804 1438 -2803
rect 100 -2806 430 -2805
rect 443 -2806 909 -2805
rect 912 -2806 1158 -2805
rect 1255 -2806 1312 -2805
rect 1363 -2806 1396 -2805
rect 114 -2808 118 -2807
rect 121 -2808 654 -2807
rect 723 -2808 1011 -2807
rect 1020 -2808 1508 -2807
rect 114 -2810 276 -2809
rect 310 -2810 409 -2809
rect 443 -2810 493 -2809
rect 506 -2810 780 -2809
rect 828 -2810 850 -2809
rect 898 -2810 955 -2809
rect 1010 -2810 1165 -2809
rect 1311 -2810 1431 -2809
rect 117 -2812 276 -2811
rect 338 -2812 423 -2811
rect 506 -2812 626 -2811
rect 653 -2812 1004 -2811
rect 1097 -2812 1284 -2811
rect 1381 -2812 1522 -2811
rect 124 -2814 332 -2813
rect 345 -2814 591 -2813
rect 597 -2814 808 -2813
rect 842 -2814 885 -2813
rect 1003 -2814 1102 -2813
rect 1129 -2814 1144 -2813
rect 1150 -2814 1270 -2813
rect 1283 -2814 1375 -2813
rect 1430 -2814 1494 -2813
rect 44 -2816 125 -2815
rect 128 -2816 514 -2815
rect 520 -2816 563 -2815
rect 565 -2816 1270 -2815
rect 1374 -2816 1466 -2815
rect 103 -2818 129 -2817
rect 135 -2818 661 -2817
rect 744 -2818 1158 -2817
rect 1164 -2818 1277 -2817
rect 135 -2820 570 -2819
rect 590 -2820 605 -2819
rect 625 -2820 948 -2819
rect 1101 -2820 1263 -2819
rect 1276 -2820 1368 -2819
rect 142 -2822 339 -2821
rect 345 -2822 402 -2821
rect 408 -2822 486 -2821
rect 513 -2822 710 -2821
rect 744 -2822 1095 -2821
rect 1129 -2822 1214 -2821
rect 1262 -2822 1361 -2821
rect 1367 -2822 1459 -2821
rect 142 -2824 150 -2823
rect 156 -2824 556 -2823
rect 597 -2824 682 -2823
rect 709 -2824 881 -2823
rect 1136 -2824 1301 -2823
rect 159 -2826 857 -2825
rect 1213 -2826 1340 -2825
rect 170 -2828 304 -2827
rect 317 -2828 1095 -2827
rect 170 -2830 251 -2829
rect 261 -2830 542 -2829
rect 548 -2830 668 -2829
rect 681 -2830 948 -2829
rect 177 -2832 479 -2831
rect 520 -2832 766 -2831
rect 779 -2832 892 -2831
rect 177 -2834 451 -2833
rect 471 -2834 486 -2833
rect 527 -2834 563 -2833
rect 632 -2834 668 -2833
rect 765 -2834 864 -2833
rect 891 -2834 990 -2833
rect 184 -2836 206 -2835
rect 212 -2836 1291 -2835
rect 72 -2838 206 -2837
rect 212 -2838 283 -2837
rect 352 -2838 458 -2837
rect 527 -2838 958 -2837
rect 989 -2838 1088 -2837
rect 72 -2840 164 -2839
rect 191 -2840 199 -2839
rect 215 -2840 678 -2839
rect 800 -2840 808 -2839
rect 842 -2840 983 -2839
rect 163 -2842 269 -2841
rect 380 -2842 643 -2841
rect 663 -2842 1340 -2841
rect 191 -2844 209 -2843
rect 233 -2844 752 -2843
rect 800 -2844 941 -2843
rect 954 -2844 1088 -2843
rect 226 -2846 234 -2845
rect 247 -2846 696 -2845
rect 845 -2846 941 -2845
rect 982 -2846 1067 -2845
rect 226 -2848 619 -2847
rect 632 -2848 1025 -2847
rect 1066 -2848 1221 -2847
rect 254 -2850 269 -2849
rect 387 -2850 815 -2849
rect 849 -2850 1074 -2849
rect 219 -2852 388 -2851
rect 401 -2852 465 -2851
rect 534 -2852 825 -2851
rect 856 -2852 962 -2851
rect 1073 -2852 1242 -2851
rect 219 -2854 818 -2853
rect 912 -2854 1291 -2853
rect 229 -2856 465 -2855
rect 534 -2856 703 -2855
rect 761 -2856 1221 -2855
rect 1241 -2856 1354 -2855
rect 240 -2858 255 -2857
rect 264 -2858 360 -2857
rect 436 -2858 472 -2857
rect 541 -2858 647 -2857
rect 674 -2858 703 -2857
rect 761 -2858 1053 -2857
rect 1353 -2858 1473 -2857
rect 79 -2860 437 -2859
rect 450 -2860 577 -2859
rect 618 -2860 640 -2859
rect 695 -2860 794 -2859
rect 814 -2860 920 -2859
rect 961 -2860 1046 -2859
rect 1052 -2860 1228 -2859
rect 79 -2862 279 -2861
rect 359 -2862 416 -2861
rect 457 -2862 916 -2861
rect 919 -2862 1123 -2861
rect 121 -2864 647 -2863
rect 793 -2864 836 -2863
rect 877 -2864 1228 -2863
rect 240 -2866 871 -2865
rect 1045 -2866 1200 -2865
rect 394 -2868 416 -2867
rect 548 -2868 717 -2867
rect 786 -2868 878 -2867
rect 1122 -2868 1319 -2867
rect 145 -2870 395 -2869
rect 555 -2870 605 -2869
rect 611 -2870 640 -2869
rect 716 -2870 759 -2869
rect 786 -2870 822 -2869
rect 870 -2870 927 -2869
rect 1192 -2870 1200 -2869
rect 1318 -2870 1389 -2869
rect 569 -2872 836 -2871
rect 926 -2872 934 -2871
rect 1017 -2872 1193 -2871
rect 1332 -2872 1389 -2871
rect 576 -2874 1039 -2873
rect 1332 -2874 1445 -2873
rect 583 -2876 612 -2875
rect 821 -2876 1109 -2875
rect 933 -2878 976 -2877
rect 1017 -2878 1025 -2877
rect 1038 -2878 1207 -2877
rect 975 -2880 1060 -2879
rect 1108 -2880 1235 -2879
rect 1059 -2882 1081 -2881
rect 1206 -2882 1403 -2881
rect 1080 -2884 1172 -2883
rect 1234 -2884 1347 -2883
rect 1402 -2884 1515 -2883
rect 1171 -2886 1249 -2885
rect 1346 -2886 1452 -2885
rect 1248 -2888 1410 -2887
rect 905 -2890 1410 -2889
rect 905 -2892 969 -2891
rect 968 -2894 1116 -2893
rect 1115 -2896 1179 -2895
rect 1178 -2898 1305 -2897
rect 1304 -2900 1424 -2899
rect 1416 -2902 1424 -2901
rect 1031 -2904 1417 -2903
rect 663 -2906 1032 -2905
rect 72 -2917 248 -2916
rect 250 -2917 570 -2916
rect 583 -2917 955 -2916
rect 957 -2917 1186 -2916
rect 1227 -2917 1231 -2916
rect 1360 -2917 1431 -2916
rect 93 -2919 125 -2918
rect 166 -2919 577 -2918
rect 586 -2919 619 -2918
rect 754 -2919 794 -2918
rect 800 -2919 1095 -2918
rect 1097 -2919 1249 -2918
rect 1360 -2919 1410 -2918
rect 93 -2921 206 -2920
rect 208 -2921 311 -2920
rect 436 -2921 703 -2920
rect 765 -2921 794 -2920
rect 838 -2921 1193 -2920
rect 1227 -2921 1256 -2920
rect 1409 -2921 1424 -2920
rect 100 -2923 150 -2922
rect 184 -2923 286 -2922
rect 289 -2923 297 -2922
rect 310 -2923 325 -2922
rect 457 -2923 825 -2922
rect 838 -2923 885 -2922
rect 891 -2923 895 -2922
rect 912 -2923 1172 -2922
rect 1185 -2923 1214 -2922
rect 1248 -2923 1298 -2922
rect 103 -2925 745 -2924
rect 768 -2925 1116 -2924
rect 1192 -2925 1235 -2924
rect 1276 -2925 1298 -2924
rect 121 -2927 850 -2926
rect 884 -2927 927 -2926
rect 947 -2927 983 -2926
rect 1017 -2927 1060 -2926
rect 1076 -2927 1221 -2926
rect 1234 -2927 1291 -2926
rect 121 -2929 213 -2928
rect 219 -2929 577 -2928
rect 604 -2929 619 -2928
rect 667 -2929 703 -2928
rect 744 -2929 752 -2928
rect 789 -2929 1081 -2928
rect 1087 -2929 1116 -2928
rect 1213 -2929 1242 -2928
rect 1269 -2929 1277 -2928
rect 142 -2931 437 -2930
rect 457 -2931 591 -2930
rect 604 -2931 738 -2930
rect 821 -2931 983 -2930
rect 1024 -2931 1060 -2930
rect 1080 -2931 1130 -2930
rect 1220 -2931 1263 -2930
rect 1269 -2931 1326 -2930
rect 107 -2933 591 -2932
rect 611 -2933 643 -2932
rect 646 -2933 668 -2932
rect 681 -2933 850 -2932
rect 891 -2933 906 -2932
rect 912 -2933 990 -2932
rect 1094 -2933 1158 -2932
rect 1206 -2933 1326 -2932
rect 107 -2935 549 -2934
rect 597 -2935 612 -2934
rect 691 -2935 1088 -2934
rect 1101 -2935 1172 -2934
rect 1230 -2935 1256 -2934
rect 1262 -2935 1312 -2934
rect 142 -2937 647 -2936
rect 709 -2937 738 -2936
rect 807 -2937 1025 -2936
rect 1052 -2937 1158 -2936
rect 1241 -2937 1333 -2936
rect 184 -2939 640 -2938
rect 772 -2939 808 -2938
rect 821 -2939 871 -2938
rect 898 -2939 948 -2938
rect 954 -2939 962 -2938
rect 989 -2939 1046 -2938
rect 1066 -2939 1102 -2938
rect 1129 -2939 1165 -2938
rect 1304 -2939 1333 -2938
rect 208 -2941 234 -2940
rect 240 -2941 801 -2940
rect 835 -2941 1053 -2940
rect 1108 -2941 1165 -2940
rect 1311 -2941 1389 -2940
rect 212 -2943 367 -2942
rect 411 -2943 1291 -2942
rect 1388 -2943 1417 -2942
rect 222 -2945 451 -2944
rect 495 -2945 927 -2944
rect 950 -2945 1046 -2944
rect 1143 -2945 1207 -2944
rect 226 -2947 269 -2946
rect 275 -2947 584 -2946
rect 597 -2947 626 -2946
rect 639 -2947 661 -2946
rect 688 -2947 836 -2946
rect 842 -2947 1396 -2946
rect 163 -2949 269 -2948
rect 275 -2949 423 -2948
rect 443 -2949 682 -2948
rect 751 -2949 1067 -2948
rect 1143 -2949 1151 -2948
rect 163 -2951 381 -2950
rect 443 -2951 472 -2950
rect 513 -2951 626 -2950
rect 660 -2951 1396 -2950
rect 135 -2953 472 -2952
rect 520 -2953 650 -2952
rect 772 -2953 787 -2952
rect 842 -2953 857 -2952
rect 870 -2953 1123 -2952
rect 135 -2955 654 -2954
rect 898 -2955 934 -2954
rect 961 -2955 976 -2954
rect 1017 -2955 1123 -2954
rect 149 -2957 857 -2956
rect 915 -2957 1039 -2956
rect 191 -2959 423 -2958
rect 464 -2959 934 -2958
rect 1031 -2959 1305 -2958
rect 191 -2961 199 -2960
rect 229 -2961 633 -2960
rect 786 -2961 976 -2960
rect 1038 -2961 1074 -2960
rect 86 -2963 199 -2962
rect 233 -2963 293 -2962
rect 296 -2963 689 -2962
rect 919 -2963 1004 -2962
rect 1073 -2963 1319 -2962
rect 79 -2965 87 -2964
rect 219 -2965 920 -2964
rect 940 -2965 1032 -2964
rect 1283 -2965 1319 -2964
rect 240 -2967 374 -2966
rect 387 -2967 654 -2966
rect 674 -2967 941 -2966
rect 1003 -2967 1011 -2966
rect 1283 -2967 1340 -2966
rect 170 -2969 388 -2968
rect 401 -2969 514 -2968
rect 520 -2969 867 -2968
rect 1339 -2969 1347 -2968
rect 170 -2971 874 -2970
rect 1346 -2971 1382 -2970
rect 247 -2973 762 -2972
rect 282 -2975 748 -2974
rect 254 -2977 283 -2976
rect 289 -2977 664 -2976
rect 674 -2977 916 -2976
rect 254 -2979 279 -2978
rect 303 -2979 367 -2978
rect 373 -2979 395 -2978
rect 464 -2979 486 -2978
rect 534 -2979 570 -2978
rect 632 -2979 1109 -2978
rect 261 -2981 535 -2980
rect 548 -2981 878 -2980
rect 261 -2983 381 -2982
rect 394 -2983 409 -2982
rect 485 -2983 717 -2982
rect 303 -2985 318 -2984
rect 324 -2985 507 -2984
rect 555 -2985 867 -2984
rect 317 -2987 339 -2986
rect 345 -2987 451 -2986
rect 562 -2987 710 -2986
rect 716 -2987 864 -2986
rect 145 -2989 339 -2988
rect 345 -2989 500 -2988
rect 695 -2989 864 -2988
rect 264 -2991 563 -2990
rect 698 -2991 1011 -2990
rect 359 -2993 402 -2992
rect 408 -2993 878 -2992
rect 359 -2995 479 -2994
rect 499 -2995 636 -2994
rect 705 -2995 1382 -2994
rect 429 -2997 696 -2996
rect 177 -2999 430 -2998
rect 478 -2999 542 -2998
rect 156 -3001 178 -3000
rect 541 -3001 724 -3000
rect 156 -3003 353 -3002
rect 723 -3003 731 -3002
rect 352 -3005 416 -3004
rect 730 -3005 815 -3004
rect 331 -3007 416 -3006
rect 779 -3007 815 -3006
rect 114 -3009 332 -3008
rect 779 -3009 923 -3008
rect 114 -3011 1021 -3010
rect 922 -3013 1354 -3012
rect 1353 -3015 1368 -3014
rect 1367 -3017 1375 -3016
rect 1374 -3019 1403 -3018
rect 758 -3021 1403 -3020
rect 527 -3023 759 -3022
rect 527 -3025 664 -3024
rect 86 -3036 150 -3035
rect 156 -3036 409 -3035
rect 411 -3036 654 -3035
rect 660 -3036 983 -3035
rect 1017 -3036 1046 -3035
rect 1073 -3036 1403 -3035
rect 93 -3038 811 -3037
rect 835 -3038 1172 -3037
rect 100 -3040 153 -3039
rect 198 -3040 209 -3039
rect 275 -3040 279 -3039
rect 289 -3040 507 -3039
rect 516 -3040 542 -3039
rect 555 -3040 654 -3039
rect 660 -3040 878 -3039
rect 919 -3040 1333 -3039
rect 100 -3042 129 -3041
rect 135 -3042 206 -3041
rect 275 -3042 367 -3041
rect 422 -3042 916 -3041
rect 926 -3042 1336 -3041
rect 107 -3044 223 -3043
rect 310 -3044 412 -3043
rect 471 -3044 542 -3043
rect 576 -3044 633 -3043
rect 681 -3044 696 -3043
rect 698 -3044 990 -3043
rect 1020 -3044 1277 -3043
rect 107 -3046 262 -3045
rect 310 -3046 867 -3045
rect 873 -3046 1396 -3045
rect 128 -3048 234 -3047
rect 324 -3048 839 -3047
rect 863 -3048 1326 -3047
rect 135 -3050 1210 -3049
rect 1241 -3050 1277 -3049
rect 1325 -3050 1382 -3049
rect 149 -3052 923 -3051
rect 926 -3052 997 -3051
rect 1038 -3052 1074 -3051
rect 1136 -3052 1172 -3051
rect 1241 -3052 1270 -3051
rect 170 -3054 199 -3053
rect 229 -3054 262 -3053
rect 327 -3054 647 -3053
rect 691 -3054 1256 -3053
rect 170 -3056 248 -3055
rect 338 -3056 472 -3055
rect 513 -3056 556 -3055
rect 583 -3056 990 -3055
rect 1038 -3056 1067 -3055
rect 1115 -3056 1137 -3055
rect 1150 -3056 1298 -3055
rect 184 -3058 290 -3057
rect 338 -3058 528 -3057
rect 534 -3058 608 -3057
rect 618 -3058 650 -3057
rect 698 -3058 1179 -3057
rect 1234 -3058 1256 -3057
rect 1297 -3058 1333 -3057
rect 184 -3060 227 -3059
rect 233 -3060 255 -3059
rect 345 -3060 510 -3059
rect 527 -3060 591 -3059
rect 618 -3060 766 -3059
rect 789 -3060 871 -3059
rect 877 -3060 1221 -3059
rect 121 -3062 227 -3061
rect 345 -3062 437 -3061
rect 443 -3062 577 -3061
rect 590 -3062 1088 -3061
rect 1150 -3062 1207 -3061
rect 1220 -3062 1228 -3061
rect 121 -3064 220 -3063
rect 331 -3064 437 -3063
rect 464 -3064 514 -3063
rect 534 -3064 598 -3063
rect 635 -3064 682 -3063
rect 730 -3064 734 -3063
rect 740 -3064 948 -3063
rect 982 -3064 1203 -3063
rect 1213 -3064 1228 -3063
rect 166 -3066 332 -3065
rect 352 -3066 367 -3065
rect 380 -3066 465 -3065
rect 478 -3066 584 -3065
rect 597 -3066 668 -3065
rect 730 -3066 794 -3065
rect 796 -3066 1235 -3065
rect 177 -3068 255 -3067
rect 257 -3068 479 -3067
rect 520 -3068 668 -3067
rect 744 -3068 766 -3067
rect 835 -3068 843 -3067
rect 863 -3068 892 -3067
rect 898 -3068 920 -3067
rect 1045 -3068 1102 -3067
rect 1178 -3068 1368 -3067
rect 177 -3070 500 -3069
rect 520 -3070 640 -3069
rect 649 -3070 1088 -3069
rect 1101 -3070 1123 -3069
rect 1213 -3070 1305 -3069
rect 1367 -3070 1389 -3069
rect 282 -3072 353 -3071
rect 380 -3072 458 -3071
rect 499 -3072 605 -3071
rect 611 -3072 640 -3071
rect 744 -3072 1158 -3071
rect 1304 -3072 1354 -3071
rect 394 -3074 423 -3073
rect 429 -3074 458 -3073
rect 548 -3074 612 -3073
rect 733 -3074 794 -3073
rect 842 -3074 906 -3073
rect 933 -3074 1158 -3073
rect 1353 -3074 1361 -3073
rect 303 -3076 549 -3075
rect 747 -3076 1270 -3075
rect 1360 -3076 1375 -3075
rect 303 -3078 388 -3077
rect 394 -3078 762 -3077
rect 887 -3078 948 -3077
rect 1059 -3078 1067 -3077
rect 1122 -3078 1130 -3077
rect 1374 -3078 1410 -3077
rect 401 -3080 430 -3079
rect 751 -3080 780 -3079
rect 891 -3080 955 -3079
rect 1059 -3080 1081 -3079
rect 1108 -3080 1130 -3079
rect 296 -3082 402 -3081
rect 415 -3082 444 -3081
rect 772 -3082 780 -3081
rect 898 -3082 1200 -3081
rect 296 -3084 374 -3083
rect 415 -3084 755 -3083
rect 758 -3084 773 -3083
rect 901 -3084 1116 -3083
rect 373 -3086 689 -3085
rect 905 -3086 1025 -3085
rect 1080 -3086 1144 -3085
rect 688 -3088 724 -3087
rect 933 -3088 962 -3087
rect 1024 -3088 1053 -3087
rect 1108 -3088 1193 -3087
rect 674 -3090 1053 -3089
rect 1143 -3090 1186 -3089
rect 1192 -3090 1291 -3089
rect 674 -3092 703 -3091
rect 716 -3092 724 -3091
rect 940 -3092 962 -3091
rect 1003 -3092 1186 -3091
rect 1290 -3092 1340 -3091
rect 485 -3094 717 -3093
rect 940 -3094 969 -3093
rect 1003 -3094 1032 -3093
rect 1339 -3094 1347 -3093
rect 317 -3096 486 -3095
rect 702 -3096 710 -3095
rect 912 -3096 969 -3095
rect 1031 -3096 1095 -3095
rect 163 -3098 1095 -3097
rect 163 -3100 269 -3099
rect 317 -3100 360 -3099
rect 562 -3100 710 -3099
rect 912 -3100 1165 -3099
rect 212 -3102 269 -3101
rect 324 -3102 563 -3101
rect 954 -3102 976 -3101
rect 1164 -3102 1263 -3101
rect 191 -3104 213 -3103
rect 240 -3104 360 -3103
rect 975 -3104 1011 -3103
rect 1248 -3104 1263 -3103
rect 156 -3106 192 -3105
rect 240 -3106 1154 -3105
rect 695 -3108 1249 -3107
rect 1010 -3110 1319 -3109
rect 1311 -3112 1319 -3111
rect 884 -3114 1312 -3113
rect 856 -3116 885 -3115
rect 849 -3118 857 -3117
rect 828 -3120 850 -3119
rect 814 -3122 829 -3121
rect 814 -3124 822 -3123
rect 737 -3126 822 -3125
rect 492 -3128 738 -3127
rect 492 -3130 787 -3129
rect 786 -3132 801 -3131
rect 800 -3134 808 -3133
rect 807 -3136 997 -3135
rect 100 -3147 160 -3146
rect 184 -3147 325 -3146
rect 331 -3147 391 -3146
rect 394 -3147 755 -3146
rect 758 -3147 815 -3146
rect 898 -3147 1172 -3146
rect 1199 -3147 1221 -3146
rect 1293 -3147 1340 -3146
rect 1346 -3147 1361 -3146
rect 107 -3149 286 -3148
rect 296 -3149 696 -3148
rect 698 -3149 969 -3148
rect 1171 -3149 1214 -3148
rect 1335 -3149 1368 -3148
rect 114 -3151 188 -3150
rect 191 -3151 251 -3150
rect 254 -3151 374 -3150
rect 387 -3151 486 -3150
rect 492 -3151 811 -3150
rect 870 -3151 899 -3150
rect 912 -3151 1200 -3150
rect 1206 -3151 1242 -3150
rect 1360 -3151 1375 -3150
rect 121 -3153 223 -3152
rect 247 -3153 353 -3152
rect 373 -3153 430 -3152
rect 460 -3153 528 -3152
rect 593 -3153 1287 -3152
rect 177 -3155 388 -3154
rect 394 -3155 458 -3154
rect 464 -3155 545 -3154
rect 607 -3155 1158 -3154
rect 1206 -3155 1277 -3154
rect 177 -3157 769 -3156
rect 807 -3157 895 -3156
rect 915 -3157 1231 -3156
rect 1241 -3157 1319 -3156
rect 191 -3159 748 -3158
rect 758 -3159 850 -3158
rect 870 -3159 885 -3158
rect 943 -3159 1137 -3158
rect 1209 -3159 1221 -3158
rect 1276 -3159 1326 -3158
rect 198 -3161 227 -3160
rect 233 -3161 248 -3160
rect 275 -3161 297 -3160
rect 327 -3161 486 -3160
rect 492 -3161 612 -3160
rect 618 -3161 1011 -3160
rect 1059 -3161 1137 -3160
rect 1213 -3161 1305 -3160
rect 128 -3163 199 -3162
rect 219 -3163 290 -3162
rect 331 -3163 381 -3162
rect 401 -3163 619 -3162
rect 635 -3163 829 -3162
rect 849 -3163 976 -3162
rect 1234 -3163 1305 -3162
rect 135 -3165 276 -3164
rect 338 -3165 591 -3164
rect 611 -3165 682 -3164
rect 695 -3165 773 -3164
rect 810 -3165 1186 -3164
rect 1234 -3165 1291 -3164
rect 184 -3167 290 -3166
rect 338 -3167 367 -3166
rect 401 -3167 437 -3166
rect 464 -3167 1333 -3166
rect 233 -3169 283 -3168
rect 345 -3169 748 -3168
rect 772 -3169 787 -3168
rect 877 -3169 1060 -3168
rect 1108 -3169 1186 -3168
rect 282 -3171 325 -3170
rect 345 -3171 451 -3170
rect 506 -3171 745 -3170
rect 761 -3171 787 -3170
rect 877 -3171 955 -3170
rect 968 -3171 983 -3170
rect 1108 -3171 1228 -3170
rect 205 -3173 451 -3172
rect 471 -3173 507 -3172
rect 520 -3173 738 -3172
rect 740 -3173 1158 -3172
rect 205 -3175 262 -3174
rect 352 -3175 535 -3174
rect 590 -3175 745 -3174
rect 884 -3175 892 -3174
rect 905 -3175 955 -3174
rect 975 -3175 1025 -3174
rect 142 -3177 262 -3176
rect 317 -3177 892 -3176
rect 905 -3177 934 -3176
rect 982 -3177 1018 -3176
rect 1024 -3177 1102 -3176
rect 240 -3179 318 -3178
rect 359 -3179 381 -3178
rect 415 -3179 430 -3178
rect 471 -3179 556 -3178
rect 625 -3179 738 -3178
rect 919 -3179 1011 -3178
rect 1101 -3179 1144 -3178
rect 240 -3181 605 -3180
rect 646 -3181 766 -3180
rect 919 -3181 1203 -3180
rect 359 -3183 412 -3182
rect 422 -3183 437 -3182
rect 443 -3183 605 -3182
rect 646 -3183 710 -3182
rect 716 -3183 902 -3182
rect 926 -3183 934 -3182
rect 996 -3183 1018 -3182
rect 1143 -3183 1263 -3182
rect 366 -3185 640 -3184
rect 667 -3185 829 -3184
rect 926 -3185 1004 -3184
rect 1150 -3185 1203 -3184
rect 408 -3187 416 -3186
rect 422 -3187 500 -3186
rect 513 -3187 626 -3186
rect 667 -3187 794 -3186
rect 961 -3187 1263 -3186
rect 163 -3189 409 -3188
rect 443 -3189 458 -3188
rect 513 -3189 654 -3188
rect 681 -3189 752 -3188
rect 765 -3189 1312 -3188
rect 156 -3191 164 -3190
rect 303 -3191 500 -3190
rect 520 -3191 549 -3190
rect 555 -3191 570 -3190
rect 597 -3191 640 -3190
rect 709 -3191 1179 -3190
rect 303 -3193 311 -3192
rect 527 -3193 542 -3192
rect 548 -3193 577 -3192
rect 597 -3193 808 -3192
rect 996 -3193 1095 -3192
rect 1150 -3193 1270 -3192
rect 149 -3195 311 -3194
rect 534 -3195 822 -3194
rect 947 -3195 1095 -3194
rect 562 -3197 654 -3196
rect 716 -3197 731 -3196
rect 751 -3197 1179 -3196
rect 562 -3199 584 -3198
rect 730 -3199 780 -3198
rect 793 -3199 801 -3198
rect 821 -3199 836 -3198
rect 940 -3199 948 -3198
rect 1003 -3199 1074 -3198
rect 170 -3201 801 -3200
rect 835 -3201 857 -3200
rect 940 -3201 1067 -3200
rect 170 -3203 724 -3202
rect 856 -3203 990 -3202
rect 1031 -3203 1074 -3202
rect 478 -3205 780 -3204
rect 989 -3205 1039 -3204
rect 1066 -3205 1256 -3204
rect 478 -3207 1130 -3206
rect 516 -3209 584 -3208
rect 723 -3209 1088 -3208
rect 1129 -3209 1249 -3208
rect 569 -3211 633 -3210
rect 814 -3211 1256 -3210
rect 229 -3213 633 -3212
rect 1031 -3213 1116 -3212
rect 1248 -3213 1284 -3212
rect 576 -3215 703 -3214
rect 961 -3215 1116 -3214
rect 1269 -3215 1284 -3214
rect 688 -3217 703 -3216
rect 1038 -3217 1053 -3216
rect 1087 -3217 1291 -3216
rect 660 -3219 689 -3218
rect 1052 -3219 1081 -3218
rect 660 -3221 675 -3220
rect 1080 -3221 1123 -3220
rect 674 -3223 1168 -3222
rect 1122 -3225 1165 -3224
rect 1164 -3227 1193 -3226
rect 796 -3229 1193 -3228
rect 156 -3240 213 -3239
rect 219 -3240 461 -3239
rect 499 -3240 710 -3239
rect 712 -3240 1256 -3239
rect 1290 -3240 1305 -3239
rect 1339 -3240 1361 -3239
rect 163 -3242 202 -3241
rect 212 -3242 241 -3241
rect 243 -3242 325 -3241
rect 352 -3242 664 -3241
rect 733 -3242 815 -3241
rect 838 -3242 1193 -3241
rect 1199 -3242 1207 -3241
rect 1227 -3242 1284 -3241
rect 1293 -3242 1298 -3241
rect 1346 -3242 1350 -3241
rect 163 -3244 367 -3243
rect 394 -3244 545 -3243
rect 548 -3244 577 -3243
rect 632 -3244 682 -3243
rect 744 -3244 1067 -3243
rect 1136 -3244 1256 -3243
rect 1346 -3244 1354 -3243
rect 170 -3246 482 -3245
rect 499 -3246 748 -3245
rect 751 -3246 773 -3245
rect 807 -3246 1228 -3245
rect 1349 -3246 1354 -3245
rect 170 -3248 657 -3247
rect 667 -3248 752 -3247
rect 758 -3248 773 -3247
rect 807 -3248 895 -3247
rect 933 -3248 1067 -3247
rect 1164 -3248 1235 -3247
rect 177 -3250 395 -3249
rect 408 -3250 479 -3249
rect 541 -3250 738 -3249
rect 758 -3250 794 -3249
rect 810 -3250 1039 -3249
rect 1045 -3250 1259 -3249
rect 177 -3252 283 -3251
rect 289 -3252 815 -3251
rect 863 -3252 934 -3251
rect 947 -3252 1039 -3251
rect 1143 -3252 1165 -3251
rect 1178 -3252 1207 -3251
rect 1220 -3252 1235 -3251
rect 187 -3254 255 -3253
rect 282 -3254 297 -3253
rect 317 -3254 367 -3253
rect 408 -3254 437 -3253
rect 450 -3254 580 -3253
rect 618 -3254 745 -3253
rect 765 -3254 787 -3253
rect 793 -3254 829 -3253
rect 863 -3254 885 -3253
rect 891 -3254 1004 -3253
rect 1024 -3254 1193 -3253
rect 1213 -3254 1221 -3253
rect 198 -3256 220 -3255
rect 247 -3256 255 -3255
rect 296 -3256 444 -3255
rect 450 -3256 521 -3255
rect 541 -3256 570 -3255
rect 618 -3256 913 -3255
rect 947 -3256 1088 -3255
rect 1108 -3256 1144 -3255
rect 1213 -3256 1249 -3255
rect 205 -3258 290 -3257
rect 303 -3258 318 -3257
rect 324 -3258 346 -3257
rect 352 -3258 514 -3257
rect 548 -3258 563 -3257
rect 709 -3258 1025 -3257
rect 1059 -3258 1109 -3257
rect 205 -3260 227 -3259
rect 247 -3260 647 -3259
rect 737 -3260 1273 -3259
rect 198 -3262 227 -3261
rect 303 -3262 381 -3261
rect 387 -3262 521 -3261
rect 562 -3262 755 -3261
rect 768 -3262 899 -3261
rect 912 -3262 927 -3261
rect 954 -3262 1179 -3261
rect 191 -3264 381 -3263
rect 387 -3264 780 -3263
rect 786 -3264 920 -3263
rect 954 -3264 1137 -3263
rect 191 -3266 276 -3265
rect 331 -3266 346 -3265
rect 415 -3266 671 -3265
rect 779 -3266 843 -3265
rect 870 -3266 962 -3265
rect 964 -3266 1186 -3265
rect 275 -3268 360 -3267
rect 415 -3268 661 -3267
rect 800 -3268 927 -3267
rect 996 -3268 1046 -3267
rect 1059 -3268 1074 -3267
rect 1171 -3268 1186 -3267
rect 331 -3270 465 -3269
rect 478 -3270 640 -3269
rect 646 -3270 696 -3269
rect 828 -3270 850 -3269
rect 856 -3270 962 -3269
rect 996 -3270 1032 -3269
rect 1052 -3270 1074 -3269
rect 1157 -3270 1172 -3269
rect 184 -3272 696 -3271
rect 842 -3272 969 -3271
rect 982 -3272 1032 -3271
rect 1052 -3272 1151 -3271
rect 184 -3274 234 -3273
rect 310 -3274 465 -3273
rect 485 -3274 570 -3273
rect 614 -3274 899 -3273
rect 919 -3274 976 -3273
rect 982 -3274 990 -3273
rect 1010 -3274 1249 -3273
rect 233 -3276 941 -3275
rect 968 -3276 1123 -3275
rect 1129 -3276 1151 -3275
rect 310 -3278 598 -3277
rect 625 -3278 640 -3277
rect 660 -3278 1130 -3277
rect 359 -3280 591 -3279
rect 625 -3280 692 -3279
rect 821 -3280 976 -3279
rect 989 -3280 1203 -3279
rect 422 -3282 489 -3281
rect 513 -3282 654 -3281
rect 667 -3282 801 -3281
rect 884 -3282 906 -3281
rect 940 -3282 1004 -3281
rect 1017 -3282 1088 -3281
rect 1115 -3282 1123 -3281
rect 422 -3284 556 -3283
rect 583 -3284 598 -3283
rect 653 -3284 860 -3283
rect 877 -3284 906 -3283
rect 1017 -3284 1081 -3283
rect 1094 -3284 1116 -3283
rect 429 -3286 556 -3285
rect 583 -3286 612 -3285
rect 681 -3286 822 -3285
rect 877 -3286 1263 -3285
rect 429 -3288 825 -3287
rect 1006 -3288 1081 -3287
rect 1262 -3288 1277 -3287
rect 436 -3290 493 -3289
rect 534 -3290 591 -3289
rect 611 -3290 892 -3289
rect 1027 -3290 1158 -3289
rect 1269 -3290 1277 -3289
rect 261 -3292 493 -3291
rect 688 -3292 850 -3291
rect 261 -3294 402 -3293
rect 443 -3294 507 -3293
rect 688 -3294 1011 -3293
rect 338 -3296 402 -3295
rect 457 -3296 1095 -3295
rect 338 -3298 472 -3297
rect 485 -3298 724 -3297
rect 457 -3300 605 -3299
rect 716 -3300 724 -3299
rect 471 -3302 538 -3301
rect 604 -3302 836 -3301
rect 506 -3304 675 -3303
rect 716 -3304 731 -3303
rect 674 -3306 874 -3305
rect 156 -3317 272 -3316
rect 303 -3317 486 -3316
rect 520 -3317 559 -3316
rect 576 -3317 615 -3316
rect 653 -3317 850 -3316
rect 856 -3317 1144 -3316
rect 1181 -3317 1263 -3316
rect 1269 -3317 1291 -3316
rect 163 -3319 426 -3318
rect 436 -3319 486 -3318
rect 544 -3319 752 -3318
rect 761 -3319 906 -3318
rect 1003 -3319 1074 -3318
rect 1136 -3319 1242 -3318
rect 1272 -3319 1277 -3318
rect 177 -3321 580 -3320
rect 611 -3321 640 -3320
rect 660 -3321 780 -3320
rect 786 -3321 822 -3320
rect 824 -3321 1067 -3320
rect 1073 -3321 1151 -3320
rect 184 -3323 244 -3322
rect 261 -3323 395 -3322
rect 411 -3323 874 -3322
rect 891 -3323 1032 -3322
rect 1038 -3323 1042 -3322
rect 1055 -3323 1088 -3322
rect 1139 -3323 1158 -3322
rect 198 -3325 220 -3324
rect 226 -3325 241 -3324
rect 282 -3325 304 -3324
rect 359 -3325 668 -3324
rect 670 -3325 1179 -3324
rect 226 -3327 311 -3326
rect 387 -3327 860 -3326
rect 870 -3327 1193 -3326
rect 275 -3329 360 -3328
rect 387 -3329 479 -3328
rect 513 -3329 640 -3328
rect 660 -3329 738 -3328
rect 751 -3329 773 -3328
rect 779 -3329 815 -3328
rect 835 -3329 1249 -3328
rect 275 -3331 346 -3330
rect 394 -3331 507 -3330
rect 513 -3331 654 -3330
rect 667 -3331 724 -3330
rect 737 -3331 766 -3330
rect 807 -3331 815 -3330
rect 835 -3331 927 -3330
rect 947 -3331 1088 -3330
rect 1192 -3331 1214 -3330
rect 282 -3333 297 -3332
rect 310 -3333 318 -3332
rect 345 -3333 374 -3332
rect 422 -3333 538 -3332
rect 569 -3333 773 -3332
rect 838 -3333 1116 -3332
rect 219 -3335 570 -3334
rect 572 -3335 724 -3334
rect 761 -3335 1046 -3334
rect 296 -3337 325 -3336
rect 373 -3337 402 -3336
rect 436 -3337 465 -3336
rect 478 -3337 542 -3336
rect 632 -3337 808 -3336
rect 849 -3337 962 -3336
rect 1003 -3337 1053 -3336
rect 317 -3339 409 -3338
rect 506 -3339 542 -3338
rect 632 -3339 731 -3338
rect 765 -3339 794 -3338
rect 856 -3339 941 -3338
rect 947 -3339 969 -3338
rect 1024 -3339 1235 -3338
rect 324 -3341 472 -3340
rect 534 -3341 787 -3340
rect 870 -3341 1095 -3340
rect 170 -3343 472 -3342
rect 534 -3343 549 -3342
rect 681 -3343 969 -3342
rect 1027 -3343 1186 -3342
rect 331 -3345 794 -3344
rect 884 -3345 1032 -3344
rect 1045 -3345 1109 -3344
rect 1185 -3345 1200 -3344
rect 331 -3347 444 -3346
rect 548 -3347 626 -3346
rect 688 -3347 703 -3346
rect 730 -3347 745 -3346
rect 884 -3347 1011 -3346
rect 1052 -3347 1256 -3346
rect 380 -3349 402 -3348
rect 408 -3349 465 -3348
rect 492 -3349 626 -3348
rect 702 -3349 717 -3348
rect 744 -3349 878 -3348
rect 891 -3349 913 -3348
rect 926 -3349 1228 -3348
rect 380 -3351 500 -3350
rect 597 -3351 682 -3350
rect 691 -3351 717 -3350
rect 877 -3351 983 -3350
rect 1094 -3351 1123 -3350
rect 443 -3353 528 -3352
rect 618 -3353 689 -3352
rect 894 -3353 934 -3352
rect 940 -3353 1081 -3352
rect 1122 -3353 1221 -3352
rect 450 -3355 500 -3354
rect 527 -3355 664 -3354
rect 898 -3355 1070 -3354
rect 1080 -3355 1102 -3354
rect 233 -3357 451 -3356
rect 457 -3357 598 -3356
rect 898 -3357 955 -3356
rect 961 -3357 1207 -3356
rect 233 -3359 339 -3358
rect 422 -3359 458 -3358
rect 492 -3359 605 -3358
rect 758 -3359 955 -3358
rect 975 -3359 1011 -3358
rect 1017 -3359 1102 -3358
rect 338 -3361 563 -3360
rect 576 -3361 605 -3360
rect 674 -3361 976 -3360
rect 982 -3361 1172 -3360
rect 247 -3363 675 -3362
rect 905 -3363 920 -3362
rect 933 -3363 990 -3362
rect 1013 -3363 1018 -3362
rect 191 -3365 248 -3364
rect 352 -3365 563 -3364
rect 583 -3365 619 -3364
rect 912 -3365 997 -3364
rect 352 -3367 556 -3366
rect 583 -3367 710 -3366
rect 800 -3367 997 -3366
rect 415 -3369 556 -3368
rect 590 -3369 710 -3368
rect 800 -3369 864 -3368
rect 919 -3369 1067 -3368
rect 404 -3371 591 -3370
rect 695 -3371 864 -3370
rect 989 -3371 1060 -3370
rect 415 -3373 430 -3372
rect 656 -3373 696 -3372
rect 1059 -3373 1130 -3372
rect 366 -3375 430 -3374
rect 520 -3375 657 -3374
rect 1129 -3375 1165 -3374
rect 289 -3377 367 -3376
rect 268 -3379 290 -3378
rect 198 -3390 293 -3389
rect 296 -3390 447 -3389
rect 457 -3390 461 -3389
rect 492 -3390 657 -3389
rect 723 -3390 759 -3389
rect 793 -3390 871 -3389
rect 1013 -3390 1088 -3389
rect 1101 -3390 1137 -3389
rect 1178 -3390 1186 -3389
rect 1346 -3390 1350 -3389
rect 205 -3392 279 -3391
rect 317 -3392 409 -3391
rect 422 -3392 724 -3391
rect 737 -3392 794 -3391
rect 807 -3392 811 -3391
rect 824 -3392 899 -3391
rect 1027 -3392 1123 -3391
rect 1181 -3392 1193 -3391
rect 1346 -3392 1354 -3391
rect 212 -3394 269 -3393
rect 271 -3394 692 -3393
rect 737 -3394 976 -3393
rect 1066 -3394 1081 -3393
rect 1087 -3394 1095 -3393
rect 1115 -3394 1130 -3393
rect 219 -3396 503 -3395
rect 530 -3396 577 -3395
rect 579 -3396 647 -3395
rect 649 -3396 962 -3395
rect 1010 -3396 1095 -3395
rect 247 -3398 475 -3397
rect 555 -3398 591 -3397
rect 597 -3398 647 -3397
rect 653 -3398 997 -3397
rect 1010 -3398 1046 -3397
rect 240 -3400 248 -3399
rect 261 -3400 290 -3399
rect 324 -3400 349 -3399
rect 366 -3400 405 -3399
rect 408 -3400 430 -3399
rect 450 -3400 493 -3399
rect 558 -3400 591 -3399
rect 667 -3400 759 -3399
rect 807 -3400 878 -3399
rect 933 -3400 976 -3399
rect 1031 -3400 1046 -3399
rect 226 -3402 367 -3401
rect 387 -3402 430 -3401
rect 450 -3402 612 -3401
rect 667 -3402 787 -3401
rect 859 -3402 874 -3401
rect 877 -3402 892 -3401
rect 961 -3402 1025 -3401
rect 1031 -3402 1060 -3401
rect 254 -3404 262 -3403
rect 282 -3404 318 -3403
rect 359 -3404 388 -3403
rect 401 -3404 479 -3403
rect 485 -3404 598 -3403
rect 716 -3404 934 -3403
rect 968 -3404 1025 -3403
rect 303 -3406 325 -3405
rect 345 -3406 360 -3405
rect 415 -3406 423 -3405
rect 457 -3406 528 -3405
rect 548 -3406 612 -3405
rect 716 -3406 773 -3405
rect 786 -3406 801 -3405
rect 863 -3406 888 -3405
rect 968 -3406 990 -3405
rect 233 -3408 346 -3407
rect 373 -3408 416 -3407
rect 478 -3408 507 -3407
rect 541 -3408 549 -3407
rect 569 -3408 619 -3407
rect 660 -3408 773 -3407
rect 800 -3408 815 -3407
rect 863 -3408 920 -3407
rect 1349 -3408 1354 -3407
rect 373 -3410 797 -3409
rect 919 -3410 948 -3409
rect 394 -3412 570 -3411
rect 572 -3412 958 -3411
rect 338 -3414 395 -3413
rect 485 -3414 500 -3413
rect 506 -3414 605 -3413
rect 618 -3414 696 -3413
rect 940 -3414 948 -3413
rect 310 -3416 339 -3415
rect 436 -3416 605 -3415
rect 632 -3416 696 -3415
rect 905 -3416 941 -3415
rect 310 -3418 332 -3417
rect 380 -3418 437 -3417
rect 499 -3418 780 -3417
rect 856 -3418 906 -3417
rect 331 -3420 514 -3419
rect 541 -3420 640 -3419
rect 674 -3420 815 -3419
rect 380 -3422 465 -3421
rect 513 -3422 521 -3421
rect 562 -3422 661 -3421
rect 674 -3422 752 -3421
rect 352 -3424 563 -3423
rect 576 -3424 626 -3423
rect 632 -3424 836 -3423
rect 352 -3426 412 -3425
rect 443 -3426 521 -3425
rect 625 -3426 710 -3425
rect 835 -3426 843 -3425
rect 464 -3428 472 -3427
rect 639 -3428 766 -3427
rect 842 -3428 927 -3427
rect 471 -3430 535 -3429
rect 688 -3430 780 -3429
rect 912 -3430 927 -3429
rect 534 -3432 584 -3431
rect 702 -3432 752 -3431
rect 765 -3432 829 -3431
rect 912 -3432 983 -3431
rect 583 -3434 745 -3433
rect 828 -3434 885 -3433
rect 982 -3434 1039 -3433
rect 702 -3436 731 -3435
rect 744 -3436 1018 -3435
rect 1038 -3436 1074 -3435
rect 709 -3438 822 -3437
rect 884 -3438 955 -3437
rect 730 -3440 850 -3439
rect 740 -3442 850 -3441
rect 275 -3453 290 -3452
rect 292 -3453 311 -3452
rect 331 -3453 367 -3452
rect 380 -3453 384 -3452
rect 464 -3453 468 -3452
rect 513 -3453 580 -3452
rect 611 -3453 650 -3452
rect 677 -3453 958 -3452
rect 989 -3453 1011 -3452
rect 1045 -3453 1053 -3452
rect 1080 -3453 1088 -3452
rect 1094 -3453 1123 -3452
rect 1136 -3453 1151 -3452
rect 1339 -3453 1343 -3452
rect 317 -3455 332 -3454
rect 338 -3455 346 -3454
rect 359 -3455 363 -3454
rect 380 -3455 437 -3454
rect 513 -3455 535 -3454
rect 611 -3455 668 -3454
rect 688 -3455 703 -3454
rect 726 -3455 808 -3454
rect 817 -3455 864 -3454
rect 870 -3455 885 -3454
rect 898 -3455 983 -3454
rect 996 -3455 1039 -3454
rect 1087 -3455 1172 -3454
rect 1339 -3455 1347 -3454
rect 324 -3457 339 -3456
rect 359 -3457 388 -3456
rect 408 -3457 465 -3456
rect 478 -3457 535 -3456
rect 604 -3457 668 -3456
rect 681 -3457 689 -3456
rect 691 -3457 843 -3456
rect 849 -3457 902 -3456
rect 905 -3457 1000 -3456
rect 1010 -3457 1032 -3456
rect 1108 -3457 1116 -3456
rect 1346 -3457 1354 -3456
rect 408 -3459 451 -3458
rect 478 -3459 549 -3458
rect 597 -3459 605 -3458
rect 628 -3459 1028 -3458
rect 422 -3461 451 -3460
rect 499 -3461 549 -3460
rect 562 -3461 598 -3460
rect 646 -3461 738 -3460
rect 751 -3461 755 -3460
rect 779 -3461 864 -3460
rect 877 -3461 888 -3460
rect 905 -3461 913 -3460
rect 926 -3461 930 -3460
rect 933 -3461 937 -3460
rect 940 -3461 944 -3460
rect 954 -3461 983 -3460
rect 436 -3463 472 -3462
rect 520 -3463 584 -3462
rect 653 -3463 703 -3462
rect 751 -3463 759 -3462
rect 779 -3463 825 -3462
rect 835 -3463 857 -3462
rect 891 -3463 913 -3462
rect 926 -3463 969 -3462
rect 401 -3465 472 -3464
rect 527 -3465 577 -3464
rect 590 -3465 654 -3464
rect 660 -3465 682 -3464
rect 695 -3465 741 -3464
rect 772 -3465 836 -3464
rect 933 -3465 962 -3464
rect 425 -3467 521 -3466
rect 530 -3467 661 -3466
rect 674 -3467 738 -3466
rect 772 -3467 860 -3466
rect 940 -3467 948 -3466
rect 954 -3467 976 -3466
rect 443 -3469 591 -3468
rect 786 -3469 871 -3468
rect 1342 -3469 1354 -3468
rect 443 -3471 458 -3470
rect 506 -3471 528 -3470
rect 562 -3471 619 -3470
rect 793 -3471 822 -3470
rect 828 -3471 857 -3470
rect 422 -3473 507 -3472
rect 618 -3473 626 -3472
rect 723 -3473 822 -3472
rect 446 -3475 500 -3474
rect 583 -3475 626 -3474
rect 800 -3475 843 -3474
rect 457 -3477 486 -3476
rect 709 -3477 801 -3476
rect 807 -3477 1175 -3476
rect 485 -3479 542 -3478
rect 709 -3479 731 -3478
rect 814 -3479 878 -3478
rect 541 -3481 570 -3480
rect 695 -3481 815 -3480
rect 569 -3483 633 -3482
rect 716 -3483 731 -3482
rect 555 -3485 633 -3484
rect 639 -3485 717 -3484
rect 492 -3487 556 -3486
rect 639 -3487 850 -3486
rect 429 -3489 493 -3488
rect 394 -3491 430 -3490
rect 352 -3493 395 -3492
rect 352 -3495 374 -3494
rect 373 -3497 416 -3496
rect 415 -3499 538 -3498
rect 254 -3510 297 -3509
rect 352 -3510 535 -3509
rect 555 -3510 626 -3509
rect 639 -3510 689 -3509
rect 691 -3510 773 -3509
rect 821 -3510 923 -3509
rect 947 -3510 955 -3509
rect 968 -3510 976 -3509
rect 982 -3510 1007 -3509
rect 1059 -3510 1088 -3509
rect 1122 -3510 1161 -3509
rect 1171 -3510 1179 -3509
rect 1339 -3510 1350 -3509
rect 268 -3512 276 -3511
rect 401 -3512 426 -3511
rect 429 -3512 563 -3511
rect 576 -3512 605 -3511
rect 618 -3512 626 -3511
rect 653 -3512 689 -3511
rect 730 -3512 734 -3511
rect 849 -3512 899 -3511
rect 933 -3512 948 -3511
rect 961 -3512 969 -3511
rect 996 -3512 1011 -3511
rect 1346 -3512 1354 -3511
rect 387 -3514 402 -3513
rect 422 -3514 479 -3513
rect 495 -3514 643 -3513
rect 660 -3514 724 -3513
rect 730 -3514 745 -3513
rect 842 -3514 850 -3513
rect 870 -3514 885 -3513
rect 912 -3514 934 -3513
rect 1003 -3514 1011 -3513
rect 373 -3516 423 -3515
rect 429 -3516 605 -3515
rect 667 -3516 727 -3515
rect 737 -3516 745 -3515
rect 856 -3516 871 -3515
rect 877 -3516 892 -3515
rect 912 -3516 927 -3515
rect 450 -3518 493 -3517
rect 499 -3518 535 -3517
rect 548 -3518 577 -3517
rect 590 -3518 640 -3517
rect 667 -3518 808 -3517
rect 863 -3518 878 -3517
rect 919 -3518 927 -3517
rect 394 -3520 451 -3519
rect 453 -3520 479 -3519
rect 485 -3520 493 -3519
rect 499 -3520 566 -3519
rect 597 -3520 629 -3519
rect 674 -3520 682 -3519
rect 733 -3520 738 -3519
rect 835 -3520 864 -3519
rect 359 -3522 395 -3521
rect 457 -3522 549 -3521
rect 555 -3522 570 -3521
rect 600 -3522 647 -3521
rect 677 -3522 944 -3521
rect 338 -3524 360 -3523
rect 408 -3524 458 -3523
rect 513 -3524 563 -3523
rect 569 -3524 584 -3523
rect 632 -3524 682 -3523
rect 800 -3524 836 -3523
rect 408 -3526 465 -3525
rect 467 -3526 584 -3525
rect 443 -3528 514 -3527
rect 520 -3528 580 -3527
rect 366 -3530 444 -3529
rect 464 -3530 545 -3529
rect 436 -3532 521 -3531
rect 527 -3532 591 -3531
rect 415 -3534 437 -3533
rect 527 -3534 542 -3533
rect 380 -3536 416 -3535
rect 541 -3536 696 -3535
rect 345 -3538 381 -3537
rect 695 -3538 717 -3537
rect 331 -3540 346 -3539
rect 716 -3540 780 -3539
rect 247 -3551 258 -3550
rect 296 -3551 311 -3550
rect 327 -3551 367 -3550
rect 394 -3551 433 -3550
rect 457 -3551 601 -3550
rect 604 -3551 647 -3550
rect 677 -3551 941 -3550
rect 1006 -3551 1011 -3550
rect 1038 -3551 1060 -3550
rect 1080 -3551 1088 -3550
rect 1150 -3551 1158 -3550
rect 345 -3553 353 -3552
rect 380 -3553 395 -3552
rect 443 -3553 458 -3552
rect 485 -3553 507 -3552
rect 544 -3553 577 -3552
rect 583 -3553 598 -3552
rect 618 -3553 668 -3552
rect 681 -3553 689 -3552
rect 695 -3553 699 -3552
rect 723 -3553 727 -3552
rect 849 -3553 857 -3552
rect 870 -3553 902 -3552
rect 912 -3553 920 -3552
rect 933 -3553 948 -3552
rect 488 -3555 535 -3554
rect 562 -3555 629 -3554
rect 639 -3555 661 -3554
rect 695 -3555 703 -3554
rect 723 -3555 731 -3554
rect 835 -3555 850 -3554
rect 863 -3555 920 -3554
rect 450 -3557 563 -3556
rect 702 -3557 717 -3556
rect 730 -3557 738 -3556
rect 884 -3557 923 -3556
rect 450 -3559 454 -3558
rect 464 -3559 489 -3558
rect 492 -3559 535 -3558
rect 709 -3559 717 -3558
rect 737 -3559 752 -3558
rect 891 -3559 913 -3558
rect 436 -3561 465 -3560
rect 478 -3561 493 -3560
rect 499 -3561 507 -3560
rect 751 -3561 759 -3560
rect 877 -3561 892 -3560
rect 898 -3561 983 -3560
rect 415 -3563 437 -3562
rect 471 -3563 500 -3562
rect 744 -3563 759 -3562
rect 408 -3565 416 -3564
rect 422 -3565 472 -3564
rect 478 -3565 542 -3564
rect 726 -3565 745 -3564
rect 376 -3567 409 -3566
rect 541 -3567 556 -3566
rect 555 -3569 570 -3568
rect 548 -3571 570 -3570
rect 527 -3573 549 -3572
rect 513 -3575 528 -3574
rect 513 -3577 591 -3576
rect 264 -3588 269 -3587
rect 310 -3588 328 -3587
rect 359 -3588 377 -3587
rect 394 -3588 402 -3587
rect 408 -3588 447 -3587
rect 450 -3588 458 -3587
rect 492 -3588 517 -3587
rect 520 -3588 545 -3587
rect 562 -3588 678 -3587
rect 751 -3588 755 -3587
rect 758 -3588 773 -3587
rect 849 -3588 864 -3587
rect 905 -3588 909 -3587
rect 912 -3588 920 -3587
rect 940 -3588 1046 -3587
rect 1083 -3588 1088 -3587
rect 324 -3590 328 -3589
rect 366 -3590 405 -3589
rect 408 -3590 416 -3589
rect 436 -3590 458 -3589
rect 471 -3590 493 -3589
rect 506 -3590 521 -3589
rect 534 -3590 563 -3589
rect 569 -3590 577 -3589
rect 597 -3590 605 -3589
rect 611 -3590 615 -3589
rect 646 -3590 682 -3589
rect 744 -3590 759 -3589
rect 891 -3590 906 -3589
rect 968 -3590 983 -3589
rect 985 -3590 990 -3589
rect 1031 -3590 1039 -3589
rect 443 -3592 479 -3591
rect 499 -3592 507 -3591
rect 516 -3592 542 -3591
rect 548 -3592 570 -3591
rect 597 -3592 619 -3591
rect 660 -3592 675 -3591
rect 737 -3592 745 -3591
rect 751 -3592 766 -3591
rect 975 -3592 983 -3591
rect 464 -3594 472 -3593
rect 548 -3594 556 -3593
rect 730 -3594 738 -3593
rect 754 -3594 766 -3593
rect 901 -3594 976 -3593
rect 527 -3596 556 -3595
rect 723 -3596 731 -3595
rect 709 -3598 724 -3597
rect 688 -3600 710 -3599
rect 401 -3611 405 -3610
rect 457 -3611 465 -3610
rect 492 -3611 514 -3610
rect 520 -3611 528 -3610
rect 541 -3611 549 -3610
rect 555 -3611 584 -3610
rect 590 -3611 598 -3610
rect 604 -3611 612 -3610
rect 684 -3611 801 -3610
rect 926 -3611 934 -3610
rect 975 -3611 1004 -3610
rect 1045 -3611 1081 -3610
rect 401 -3613 409 -3612
rect 506 -3613 517 -3612
rect 709 -3613 713 -3612
rect 730 -3613 776 -3612
rect 919 -3613 927 -3612
rect 1052 -3613 1060 -3612
rect 709 -3615 717 -3614
rect 751 -3615 762 -3614
rect 712 -3617 717 -3616
rect 737 -3617 752 -3616
rect 758 -3617 766 -3616
rect 744 -3619 759 -3618
rect 765 -3619 773 -3618
rect 723 -3621 745 -3620
rect 702 -3623 724 -3622
rect 695 -3625 703 -3624
rect 471 -3636 475 -3635
rect 562 -3636 573 -3635
rect 583 -3636 598 -3635
rect 719 -3636 724 -3635
rect 744 -3636 773 -3635
rect 856 -3636 860 -3635
rect 926 -3636 930 -3635
rect 982 -3636 990 -3635
rect 1031 -3636 1035 -3635
rect 1055 -3636 1060 -3635
rect 1080 -3636 1095 -3635
rect 1108 -3636 1112 -3635
rect 576 -3638 584 -3637
rect 709 -3638 724 -3637
rect 800 -3638 927 -3637
rect 985 -3638 1053 -3637
rect 569 -3640 577 -3639
rect 702 -3640 710 -3639
rect 1003 -3640 1032 -3639
rect 464 -3651 475 -3650
rect 527 -3651 535 -3650
rect 569 -3651 577 -3650
rect 583 -3651 591 -3650
rect 709 -3651 720 -3650
rect 765 -3651 773 -3650
rect 856 -3651 864 -3650
rect 929 -3651 934 -3650
rect 985 -3651 990 -3650
rect 1094 -3651 1109 -3650
rect 586 -3653 598 -3652
rect 716 -3653 724 -3652
rect 758 -3653 766 -3652
rect 751 -3655 759 -3654
rect 404 -3666 409 -3665
rect 527 -3666 535 -3665
rect 758 -3666 766 -3665
rect 768 -3666 773 -3665
<< m2contact >>
rect 226 0 227 1
rect 331 0 332 1
rect 366 0 367 1
rect 404 0 405 1
rect 415 0 416 1
rect 562 0 563 1
rect 590 0 591 1
rect 642 0 643 1
rect 667 0 668 1
rect 674 0 675 1
rect 705 0 706 1
rect 828 0 829 1
rect 254 -2 255 -1
rect 380 -2 381 -1
rect 401 -2 402 -1
rect 450 -2 451 -1
rect 457 -2 458 -1
rect 471 -2 472 -1
rect 492 -2 493 -1
rect 537 -2 538 -1
rect 765 -2 766 -1
rect 800 -2 801 -1
rect 803 -2 804 -1
rect 842 -2 843 -1
rect 275 -4 276 -3
rect 460 -4 461 -3
rect 506 -4 507 -3
rect 513 -4 514 -3
rect 516 -4 517 -3
rect 527 -4 528 -3
rect 534 -4 535 -3
rect 569 -4 570 -3
rect 317 -6 318 -5
rect 373 -6 374 -5
rect 429 -6 430 -5
rect 436 -6 437 -5
rect 135 -17 136 -16
rect 222 -17 223 -16
rect 303 -17 304 -16
rect 317 -17 318 -16
rect 327 -17 328 -16
rect 380 -17 381 -16
rect 383 -17 384 -16
rect 534 -17 535 -16
rect 541 -17 542 -16
rect 548 -17 549 -16
rect 565 -17 566 -16
rect 709 -17 710 -16
rect 775 -17 776 -16
rect 800 -17 801 -16
rect 821 -17 822 -16
rect 919 -17 920 -16
rect 191 -19 192 -18
rect 226 -19 227 -18
rect 310 -19 311 -18
rect 338 -19 339 -18
rect 345 -19 346 -18
rect 366 -19 367 -18
rect 373 -19 374 -18
rect 443 -19 444 -18
rect 450 -19 451 -18
rect 520 -19 521 -18
rect 527 -19 528 -18
rect 541 -19 542 -18
rect 569 -19 570 -18
rect 583 -19 584 -18
rect 632 -19 633 -18
rect 667 -19 668 -18
rect 674 -19 675 -18
rect 695 -19 696 -18
rect 782 -19 783 -18
rect 793 -19 794 -18
rect 828 -19 829 -18
rect 877 -19 878 -18
rect 205 -21 206 -20
rect 254 -21 255 -20
rect 331 -21 332 -20
rect 478 -21 479 -20
rect 488 -21 489 -20
rect 555 -21 556 -20
rect 569 -21 570 -20
rect 705 -21 706 -20
rect 842 -21 843 -20
rect 856 -21 857 -20
rect 212 -23 213 -22
rect 275 -23 276 -22
rect 331 -23 332 -22
rect 404 -23 405 -22
rect 408 -23 409 -22
rect 464 -23 465 -22
rect 506 -23 507 -22
rect 513 -23 514 -22
rect 576 -23 577 -22
rect 590 -23 591 -22
rect 635 -23 636 -22
rect 653 -23 654 -22
rect 660 -23 661 -22
rect 761 -23 762 -22
rect 226 -25 227 -24
rect 296 -25 297 -24
rect 352 -25 353 -24
rect 415 -25 416 -24
rect 436 -25 437 -24
rect 446 -25 447 -24
rect 450 -25 451 -24
rect 527 -25 528 -24
rect 639 -25 640 -24
rect 702 -25 703 -24
rect 254 -27 255 -26
rect 366 -27 367 -26
rect 376 -27 377 -26
rect 422 -27 423 -26
rect 443 -27 444 -26
rect 684 -27 685 -26
rect 299 -29 300 -28
rect 415 -29 416 -28
rect 457 -29 458 -28
rect 646 -29 647 -28
rect 317 -31 318 -30
rect 446 -31 447 -30
rect 618 -31 619 -30
rect 639 -31 640 -30
rect 387 -33 388 -32
rect 394 -33 395 -32
rect 401 -33 402 -32
rect 457 -33 458 -32
rect 618 -33 619 -32
rect 786 -33 787 -32
rect 359 -35 360 -34
rect 394 -35 395 -34
rect 79 -46 80 -45
rect 236 -46 237 -45
rect 268 -46 269 -45
rect 331 -46 332 -45
rect 380 -46 381 -45
rect 446 -46 447 -45
rect 450 -46 451 -45
rect 604 -46 605 -45
rect 618 -46 619 -45
rect 807 -46 808 -45
rect 856 -46 857 -45
rect 863 -46 864 -45
rect 877 -46 878 -45
rect 905 -46 906 -45
rect 919 -46 920 -45
rect 968 -46 969 -45
rect 100 -48 101 -47
rect 135 -48 136 -47
rect 142 -48 143 -47
rect 327 -48 328 -47
rect 380 -48 381 -47
rect 572 -48 573 -47
rect 576 -48 577 -47
rect 597 -48 598 -47
rect 632 -48 633 -47
rect 653 -48 654 -47
rect 667 -48 668 -47
rect 723 -48 724 -47
rect 758 -48 759 -47
rect 870 -48 871 -47
rect 128 -50 129 -49
rect 236 -50 237 -49
rect 278 -50 279 -49
rect 303 -50 304 -49
rect 324 -50 325 -49
rect 474 -50 475 -49
rect 478 -50 479 -49
rect 611 -50 612 -49
rect 639 -50 640 -49
rect 688 -50 689 -49
rect 695 -50 696 -49
rect 751 -50 752 -49
rect 761 -50 762 -49
rect 891 -50 892 -49
rect 149 -52 150 -51
rect 317 -52 318 -51
rect 397 -52 398 -51
rect 401 -52 402 -51
rect 408 -52 409 -51
rect 506 -52 507 -51
rect 541 -52 542 -51
rect 562 -52 563 -51
rect 576 -52 577 -51
rect 583 -52 584 -51
rect 590 -52 591 -51
rect 653 -52 654 -51
rect 660 -52 661 -51
rect 667 -52 668 -51
rect 702 -52 703 -51
rect 744 -52 745 -51
rect 765 -52 766 -51
rect 772 -52 773 -51
rect 786 -52 787 -51
rect 856 -52 857 -51
rect 156 -54 157 -53
rect 254 -54 255 -53
rect 289 -54 290 -53
rect 366 -54 367 -53
rect 422 -54 423 -53
rect 467 -54 468 -53
rect 485 -54 486 -53
rect 642 -54 643 -53
rect 702 -54 703 -53
rect 824 -54 825 -53
rect 163 -56 164 -55
rect 180 -56 181 -55
rect 184 -56 185 -55
rect 191 -56 192 -55
rect 219 -56 220 -55
rect 453 -56 454 -55
rect 464 -56 465 -55
rect 695 -56 696 -55
rect 709 -56 710 -55
rect 786 -56 787 -55
rect 793 -56 794 -55
rect 814 -56 815 -55
rect 170 -58 171 -57
rect 296 -58 297 -57
rect 303 -58 304 -57
rect 359 -58 360 -57
rect 366 -58 367 -57
rect 478 -58 479 -57
rect 499 -58 500 -57
rect 569 -58 570 -57
rect 625 -58 626 -57
rect 765 -58 766 -57
rect 800 -58 801 -57
rect 821 -58 822 -57
rect 177 -60 178 -59
rect 198 -60 199 -59
rect 222 -60 223 -59
rect 359 -60 360 -59
rect 415 -60 416 -59
rect 422 -60 423 -59
rect 436 -60 437 -59
rect 471 -60 472 -59
rect 520 -60 521 -59
rect 709 -60 710 -59
rect 177 -62 178 -61
rect 464 -62 465 -61
rect 527 -62 528 -61
rect 541 -62 542 -61
rect 555 -62 556 -61
rect 716 -62 717 -61
rect 180 -64 181 -63
rect 205 -64 206 -63
rect 226 -64 227 -63
rect 254 -64 255 -63
rect 261 -64 262 -63
rect 296 -64 297 -63
rect 317 -64 318 -63
rect 352 -64 353 -63
rect 369 -64 370 -63
rect 520 -64 521 -63
rect 527 -64 528 -63
rect 740 -64 741 -63
rect 191 -66 192 -65
rect 212 -66 213 -65
rect 226 -66 227 -65
rect 583 -66 584 -65
rect 646 -66 647 -65
rect 800 -66 801 -65
rect 205 -68 206 -67
rect 373 -68 374 -67
rect 415 -68 416 -67
rect 457 -68 458 -67
rect 534 -68 535 -67
rect 660 -68 661 -67
rect 681 -68 682 -67
rect 793 -68 794 -67
rect 229 -70 230 -69
rect 429 -70 430 -69
rect 450 -70 451 -69
rect 488 -70 489 -69
rect 513 -70 514 -69
rect 534 -70 535 -69
rect 548 -70 549 -69
rect 555 -70 556 -69
rect 569 -70 570 -69
rect 618 -70 619 -69
rect 646 -70 647 -69
rect 782 -70 783 -69
rect 243 -72 244 -71
rect 352 -72 353 -71
rect 369 -72 370 -71
rect 779 -72 780 -71
rect 331 -74 332 -73
rect 681 -74 682 -73
rect 338 -76 339 -75
rect 408 -76 409 -75
rect 457 -76 458 -75
rect 628 -76 629 -75
rect 338 -78 339 -77
rect 621 -78 622 -77
rect 373 -80 374 -79
rect 387 -80 388 -79
rect 492 -80 493 -79
rect 513 -80 514 -79
rect 548 -80 549 -79
rect 593 -80 594 -79
rect 492 -82 493 -81
rect 733 -82 734 -81
rect 593 -84 594 -83
rect 674 -84 675 -83
rect 79 -95 80 -94
rect 390 -95 391 -94
rect 418 -95 419 -94
rect 758 -95 759 -94
rect 814 -95 815 -94
rect 849 -95 850 -94
rect 856 -95 857 -94
rect 919 -95 920 -94
rect 940 -95 941 -94
rect 975 -95 976 -94
rect 114 -97 115 -96
rect 338 -97 339 -96
rect 352 -97 353 -96
rect 394 -97 395 -96
rect 432 -97 433 -96
rect 709 -97 710 -96
rect 730 -97 731 -96
rect 772 -97 773 -96
rect 842 -97 843 -96
rect 947 -97 948 -96
rect 968 -97 969 -96
rect 1003 -97 1004 -96
rect 100 -99 101 -98
rect 114 -99 115 -98
rect 128 -99 129 -98
rect 226 -99 227 -98
rect 250 -99 251 -98
rect 730 -99 731 -98
rect 744 -99 745 -98
rect 835 -99 836 -98
rect 870 -99 871 -98
rect 954 -99 955 -98
rect 100 -101 101 -100
rect 117 -101 118 -100
rect 149 -101 150 -100
rect 334 -101 335 -100
rect 352 -101 353 -100
rect 415 -101 416 -100
rect 443 -101 444 -100
rect 709 -101 710 -100
rect 744 -101 745 -100
rect 786 -101 787 -100
rect 863 -101 864 -100
rect 870 -101 871 -100
rect 891 -101 892 -100
rect 961 -101 962 -100
rect 156 -103 157 -102
rect 236 -103 237 -102
rect 240 -103 241 -102
rect 443 -103 444 -102
rect 446 -103 447 -102
rect 548 -103 549 -102
rect 558 -103 559 -102
rect 968 -103 969 -102
rect 205 -105 206 -104
rect 338 -105 339 -104
rect 453 -105 454 -104
rect 716 -105 717 -104
rect 723 -105 724 -104
rect 863 -105 864 -104
rect 905 -105 906 -104
rect 926 -105 927 -104
rect 205 -107 206 -106
rect 275 -107 276 -106
rect 282 -107 283 -106
rect 310 -107 311 -106
rect 324 -107 325 -106
rect 327 -107 328 -106
rect 506 -107 507 -106
rect 779 -107 780 -106
rect 793 -107 794 -106
rect 905 -107 906 -106
rect 149 -109 150 -108
rect 275 -109 276 -108
rect 292 -109 293 -108
rect 408 -109 409 -108
rect 499 -109 500 -108
rect 506 -109 507 -108
rect 513 -109 514 -108
rect 625 -109 626 -108
rect 642 -109 643 -108
rect 828 -109 829 -108
rect 145 -111 146 -110
rect 408 -111 409 -110
rect 513 -111 514 -110
rect 684 -111 685 -110
rect 688 -111 689 -110
rect 814 -111 815 -110
rect 821 -111 822 -110
rect 891 -111 892 -110
rect 170 -113 171 -112
rect 282 -113 283 -112
rect 296 -113 297 -112
rect 415 -113 416 -112
rect 562 -113 563 -112
rect 639 -113 640 -112
rect 646 -113 647 -112
rect 649 -113 650 -112
rect 660 -113 661 -112
rect 982 -113 983 -112
rect 170 -115 171 -114
rect 467 -115 468 -114
rect 485 -115 486 -114
rect 562 -115 563 -114
rect 569 -115 570 -114
rect 933 -115 934 -114
rect 215 -117 216 -116
rect 226 -117 227 -116
rect 268 -117 269 -116
rect 299 -117 300 -116
rect 303 -117 304 -116
rect 366 -117 367 -116
rect 569 -117 570 -116
rect 632 -117 633 -116
rect 646 -117 647 -116
rect 653 -117 654 -116
rect 660 -117 661 -116
rect 740 -117 741 -116
rect 751 -117 752 -116
rect 898 -117 899 -116
rect 177 -119 178 -118
rect 299 -119 300 -118
rect 310 -119 311 -118
rect 317 -119 318 -118
rect 324 -119 325 -118
rect 380 -119 381 -118
rect 471 -119 472 -118
rect 632 -119 633 -118
rect 653 -119 654 -118
rect 807 -119 808 -118
rect 177 -121 178 -120
rect 261 -121 262 -120
rect 268 -121 269 -120
rect 303 -121 304 -120
rect 359 -121 360 -120
rect 499 -121 500 -120
rect 548 -121 549 -120
rect 751 -121 752 -120
rect 754 -121 755 -120
rect 821 -121 822 -120
rect 191 -123 192 -122
rect 261 -123 262 -122
rect 278 -123 279 -122
rect 296 -123 297 -122
rect 345 -123 346 -122
rect 359 -123 360 -122
rect 471 -123 472 -122
rect 611 -123 612 -122
rect 618 -123 619 -122
rect 884 -123 885 -122
rect 142 -125 143 -124
rect 345 -125 346 -124
rect 450 -125 451 -124
rect 618 -125 619 -124
rect 649 -125 650 -124
rect 807 -125 808 -124
rect 184 -127 185 -126
rect 191 -127 192 -126
rect 212 -127 213 -126
rect 366 -127 367 -126
rect 436 -127 437 -126
rect 450 -127 451 -126
rect 534 -127 535 -126
rect 611 -127 612 -126
rect 667 -127 668 -126
rect 989 -127 990 -126
rect 184 -129 185 -128
rect 474 -129 475 -128
rect 555 -129 556 -128
rect 667 -129 668 -128
rect 674 -129 675 -128
rect 772 -129 773 -128
rect 198 -131 199 -130
rect 212 -131 213 -130
rect 254 -131 255 -130
rect 317 -131 318 -130
rect 457 -131 458 -130
rect 534 -131 535 -130
rect 583 -131 584 -130
rect 877 -131 878 -130
rect 198 -133 199 -132
rect 219 -133 220 -132
rect 240 -133 241 -132
rect 254 -133 255 -132
rect 285 -133 286 -132
rect 436 -133 437 -132
rect 457 -133 458 -132
rect 509 -133 510 -132
rect 583 -133 584 -132
rect 604 -133 605 -132
rect 674 -133 675 -132
rect 761 -133 762 -132
rect 765 -133 766 -132
rect 786 -133 787 -132
rect 219 -135 220 -134
rect 271 -135 272 -134
rect 285 -135 286 -134
rect 331 -135 332 -134
rect 492 -135 493 -134
rect 604 -135 605 -134
rect 688 -135 689 -134
rect 702 -135 703 -134
rect 716 -135 717 -134
rect 800 -135 801 -134
rect 422 -137 423 -136
rect 492 -137 493 -136
rect 520 -137 521 -136
rect 800 -137 801 -136
rect 401 -139 402 -138
rect 422 -139 423 -138
rect 520 -139 521 -138
rect 527 -139 528 -138
rect 590 -139 591 -138
rect 681 -139 682 -138
rect 695 -139 696 -138
rect 912 -139 913 -138
rect 373 -141 374 -140
rect 401 -141 402 -140
rect 429 -141 430 -140
rect 527 -141 528 -140
rect 597 -141 598 -140
rect 723 -141 724 -140
rect 289 -143 290 -142
rect 373 -143 374 -142
rect 429 -143 430 -142
rect 793 -143 794 -142
rect 233 -145 234 -144
rect 289 -145 290 -144
rect 478 -145 479 -144
rect 590 -145 591 -144
rect 681 -145 682 -144
rect 765 -145 766 -144
rect 478 -147 479 -146
rect 576 -147 577 -146
rect 702 -147 703 -146
rect 737 -147 738 -146
rect 464 -149 465 -148
rect 576 -149 577 -148
rect 464 -151 465 -150
rect 856 -151 857 -150
rect 541 -153 542 -152
rect 597 -153 598 -152
rect 488 -155 489 -154
rect 541 -155 542 -154
rect 72 -166 73 -165
rect 432 -166 433 -165
rect 450 -166 451 -165
rect 481 -166 482 -165
rect 495 -166 496 -165
rect 590 -166 591 -165
rect 618 -166 619 -165
rect 863 -166 864 -165
rect 870 -166 871 -165
rect 940 -166 941 -165
rect 954 -166 955 -165
rect 1087 -166 1088 -165
rect 100 -168 101 -167
rect 128 -168 129 -167
rect 135 -168 136 -167
rect 352 -168 353 -167
rect 390 -168 391 -167
rect 436 -168 437 -167
rect 453 -168 454 -167
rect 527 -168 528 -167
rect 541 -168 542 -167
rect 555 -168 556 -167
rect 618 -168 619 -167
rect 716 -168 717 -167
rect 730 -168 731 -167
rect 1122 -168 1123 -167
rect 100 -170 101 -169
rect 114 -170 115 -169
rect 124 -170 125 -169
rect 1052 -170 1053 -169
rect 107 -172 108 -171
rect 870 -172 871 -171
rect 877 -172 878 -171
rect 1031 -172 1032 -171
rect 110 -174 111 -173
rect 418 -174 419 -173
rect 457 -174 458 -173
rect 590 -174 591 -173
rect 621 -174 622 -173
rect 1129 -174 1130 -173
rect 114 -176 115 -175
rect 492 -176 493 -175
rect 509 -176 510 -175
rect 1080 -176 1081 -175
rect 149 -178 150 -177
rect 247 -178 248 -177
rect 254 -178 255 -177
rect 429 -178 430 -177
rect 467 -178 468 -177
rect 674 -178 675 -177
rect 695 -178 696 -177
rect 712 -178 713 -177
rect 730 -178 731 -177
rect 982 -178 983 -177
rect 1003 -178 1004 -177
rect 1059 -178 1060 -177
rect 156 -180 157 -179
rect 492 -180 493 -179
rect 506 -180 507 -179
rect 674 -180 675 -179
rect 695 -180 696 -179
rect 989 -180 990 -179
rect 996 -180 997 -179
rect 1003 -180 1004 -179
rect 170 -182 171 -181
rect 289 -182 290 -181
rect 310 -182 311 -181
rect 341 -182 342 -181
rect 352 -182 353 -181
rect 488 -182 489 -181
rect 506 -182 507 -181
rect 520 -182 521 -181
rect 632 -182 633 -181
rect 716 -182 717 -181
rect 786 -182 787 -181
rect 863 -182 864 -181
rect 884 -182 885 -181
rect 1073 -182 1074 -181
rect 166 -184 167 -183
rect 520 -184 521 -183
rect 562 -184 563 -183
rect 632 -184 633 -183
rect 667 -184 668 -183
rect 670 -184 671 -183
rect 828 -184 829 -183
rect 1045 -184 1046 -183
rect 173 -186 174 -185
rect 292 -186 293 -185
rect 310 -186 311 -185
rect 474 -186 475 -185
rect 488 -186 489 -185
rect 698 -186 699 -185
rect 835 -186 836 -185
rect 884 -186 885 -185
rect 891 -186 892 -185
rect 1017 -186 1018 -185
rect 184 -188 185 -187
rect 450 -188 451 -187
rect 471 -188 472 -187
rect 541 -188 542 -187
rect 562 -188 563 -187
rect 702 -188 703 -187
rect 814 -188 815 -187
rect 891 -188 892 -187
rect 898 -188 899 -187
rect 1066 -188 1067 -187
rect 163 -190 164 -189
rect 184 -190 185 -189
rect 208 -190 209 -189
rect 212 -190 213 -189
rect 219 -190 220 -189
rect 247 -190 248 -189
rect 261 -190 262 -189
rect 436 -190 437 -189
rect 639 -190 640 -189
rect 702 -190 703 -189
rect 814 -190 815 -189
rect 828 -190 829 -189
rect 856 -190 857 -189
rect 982 -190 983 -189
rect 163 -192 164 -191
rect 835 -192 836 -191
rect 905 -192 906 -191
rect 989 -192 990 -191
rect 177 -194 178 -193
rect 639 -194 640 -193
rect 667 -194 668 -193
rect 744 -194 745 -193
rect 758 -194 759 -193
rect 856 -194 857 -193
rect 912 -194 913 -193
rect 1108 -194 1109 -193
rect 177 -196 178 -195
rect 303 -196 304 -195
rect 324 -196 325 -195
rect 457 -196 458 -195
rect 653 -196 654 -195
rect 758 -196 759 -195
rect 779 -196 780 -195
rect 912 -196 913 -195
rect 919 -196 920 -195
rect 1024 -196 1025 -195
rect 121 -198 122 -197
rect 324 -198 325 -197
rect 380 -198 381 -197
rect 527 -198 528 -197
rect 597 -198 598 -197
rect 653 -198 654 -197
rect 688 -198 689 -197
rect 744 -198 745 -197
rect 793 -198 794 -197
rect 905 -198 906 -197
rect 926 -198 927 -197
rect 1010 -198 1011 -197
rect 212 -200 213 -199
rect 366 -200 367 -199
rect 380 -200 381 -199
rect 422 -200 423 -199
rect 432 -200 433 -199
rect 597 -200 598 -199
rect 712 -200 713 -199
rect 793 -200 794 -199
rect 821 -200 822 -199
rect 898 -200 899 -199
rect 933 -200 934 -199
rect 1094 -200 1095 -199
rect 219 -202 220 -201
rect 268 -202 269 -201
rect 282 -202 283 -201
rect 373 -202 374 -201
rect 394 -202 395 -201
rect 464 -202 465 -201
rect 737 -202 738 -201
rect 779 -202 780 -201
rect 842 -202 843 -201
rect 926 -202 927 -201
rect 943 -202 944 -201
rect 954 -202 955 -201
rect 961 -202 962 -201
rect 1038 -202 1039 -201
rect 222 -204 223 -203
rect 303 -204 304 -203
rect 331 -204 332 -203
rect 422 -204 423 -203
rect 464 -204 465 -203
rect 478 -204 479 -203
rect 611 -204 612 -203
rect 737 -204 738 -203
rect 754 -204 755 -203
rect 933 -204 934 -203
rect 947 -204 948 -203
rect 996 -204 997 -203
rect 226 -206 227 -205
rect 275 -206 276 -205
rect 285 -206 286 -205
rect 558 -206 559 -205
rect 681 -206 682 -205
rect 961 -206 962 -205
rect 968 -206 969 -205
rect 1115 -206 1116 -205
rect 226 -208 227 -207
rect 548 -208 549 -207
rect 681 -208 682 -207
rect 947 -208 948 -207
rect 975 -208 976 -207
rect 999 -208 1000 -207
rect 240 -210 241 -209
rect 275 -210 276 -209
rect 289 -210 290 -209
rect 611 -210 612 -209
rect 705 -210 706 -209
rect 968 -210 969 -209
rect 250 -212 251 -211
rect 282 -212 283 -211
rect 317 -212 318 -211
rect 975 -212 976 -211
rect 261 -214 262 -213
rect 429 -214 430 -213
rect 478 -214 479 -213
rect 877 -214 878 -213
rect 271 -216 272 -215
rect 331 -216 332 -215
rect 359 -216 360 -215
rect 373 -216 374 -215
rect 394 -216 395 -215
rect 408 -216 409 -215
rect 415 -216 416 -215
rect 513 -216 514 -215
rect 548 -216 549 -215
rect 583 -216 584 -215
rect 772 -216 773 -215
rect 821 -216 822 -215
rect 849 -216 850 -215
rect 919 -216 920 -215
rect 205 -218 206 -217
rect 359 -218 360 -217
rect 366 -218 367 -217
rect 684 -218 685 -217
rect 723 -218 724 -217
rect 772 -218 773 -217
rect 205 -220 206 -219
rect 485 -220 486 -219
rect 513 -220 514 -219
rect 660 -220 661 -219
rect 765 -220 766 -219
rect 849 -220 850 -219
rect 257 -222 258 -221
rect 408 -222 409 -221
rect 604 -222 605 -221
rect 660 -222 661 -221
rect 765 -222 766 -221
rect 786 -222 787 -221
rect 345 -224 346 -223
rect 583 -224 584 -223
rect 646 -224 647 -223
rect 723 -224 724 -223
rect 278 -226 279 -225
rect 345 -226 346 -225
rect 401 -226 402 -225
rect 404 -226 405 -225
rect 569 -226 570 -225
rect 604 -226 605 -225
rect 401 -228 402 -227
rect 751 -228 752 -227
rect 534 -230 535 -229
rect 569 -230 570 -229
rect 576 -230 577 -229
rect 646 -230 647 -229
rect 233 -232 234 -231
rect 576 -232 577 -231
rect 191 -234 192 -233
rect 233 -234 234 -233
rect 534 -234 535 -233
rect 807 -234 808 -233
rect 191 -236 192 -235
rect 446 -236 447 -235
rect 800 -236 801 -235
rect 807 -236 808 -235
rect 709 -238 710 -237
rect 800 -238 801 -237
rect 387 -240 388 -239
rect 709 -240 710 -239
rect 387 -242 388 -241
rect 499 -242 500 -241
rect 443 -244 444 -243
rect 499 -244 500 -243
rect 296 -246 297 -245
rect 443 -246 444 -245
rect 296 -248 297 -247
rect 338 -248 339 -247
rect 338 -250 339 -249
rect 1101 -250 1102 -249
rect 54 -261 55 -260
rect 282 -261 283 -260
rect 296 -261 297 -260
rect 443 -261 444 -260
rect 481 -261 482 -260
rect 576 -261 577 -260
rect 614 -261 615 -260
rect 1031 -261 1032 -260
rect 1038 -261 1039 -260
rect 1206 -261 1207 -260
rect 72 -263 73 -262
rect 121 -263 122 -262
rect 124 -263 125 -262
rect 208 -263 209 -262
rect 219 -263 220 -262
rect 912 -263 913 -262
rect 947 -263 948 -262
rect 1031 -263 1032 -262
rect 1052 -263 1053 -262
rect 1262 -263 1263 -262
rect 79 -265 80 -264
rect 1185 -265 1186 -264
rect 86 -267 87 -266
rect 100 -267 101 -266
rect 110 -267 111 -266
rect 338 -267 339 -266
rect 345 -267 346 -266
rect 429 -267 430 -266
rect 481 -267 482 -266
rect 856 -267 857 -266
rect 898 -267 899 -266
rect 947 -267 948 -266
rect 954 -267 955 -266
rect 1136 -267 1137 -266
rect 93 -269 94 -268
rect 579 -269 580 -268
rect 635 -269 636 -268
rect 1178 -269 1179 -268
rect 100 -271 101 -270
rect 373 -271 374 -270
rect 401 -271 402 -270
rect 471 -271 472 -270
rect 485 -271 486 -270
rect 506 -271 507 -270
rect 516 -271 517 -270
rect 716 -271 717 -270
rect 726 -271 727 -270
rect 1143 -271 1144 -270
rect 124 -273 125 -272
rect 1052 -273 1053 -272
rect 1059 -273 1060 -272
rect 1227 -273 1228 -272
rect 128 -275 129 -274
rect 131 -275 132 -274
rect 142 -275 143 -274
rect 191 -275 192 -274
rect 219 -275 220 -274
rect 604 -275 605 -274
rect 663 -275 664 -274
rect 1066 -275 1067 -274
rect 1073 -275 1074 -274
rect 1241 -275 1242 -274
rect 128 -277 129 -276
rect 205 -277 206 -276
rect 240 -277 241 -276
rect 261 -277 262 -276
rect 289 -277 290 -276
rect 345 -277 346 -276
rect 359 -277 360 -276
rect 401 -277 402 -276
rect 457 -277 458 -276
rect 506 -277 507 -276
rect 530 -277 531 -276
rect 842 -277 843 -276
rect 849 -277 850 -276
rect 898 -277 899 -276
rect 954 -277 955 -276
rect 1129 -277 1130 -276
rect 149 -279 150 -278
rect 233 -279 234 -278
rect 254 -279 255 -278
rect 583 -279 584 -278
rect 604 -279 605 -278
rect 1045 -279 1046 -278
rect 1080 -279 1081 -278
rect 1269 -279 1270 -278
rect 156 -281 157 -280
rect 338 -281 339 -280
rect 488 -281 489 -280
rect 1038 -281 1039 -280
rect 1087 -281 1088 -280
rect 1290 -281 1291 -280
rect 163 -283 164 -282
rect 436 -283 437 -282
rect 467 -283 468 -282
rect 1087 -283 1088 -282
rect 1094 -283 1095 -282
rect 1283 -283 1284 -282
rect 82 -285 83 -284
rect 436 -285 437 -284
rect 492 -285 493 -284
rect 737 -285 738 -284
rect 744 -285 745 -284
rect 856 -285 857 -284
rect 877 -285 878 -284
rect 1066 -285 1067 -284
rect 163 -287 164 -286
rect 415 -287 416 -286
rect 541 -287 542 -286
rect 730 -287 731 -286
rect 765 -287 766 -286
rect 1276 -287 1277 -286
rect 184 -289 185 -288
rect 191 -289 192 -288
rect 198 -289 199 -288
rect 205 -289 206 -288
rect 212 -289 213 -288
rect 457 -289 458 -288
rect 513 -289 514 -288
rect 541 -289 542 -288
rect 544 -289 545 -288
rect 1150 -289 1151 -288
rect 58 -291 59 -290
rect 212 -291 213 -290
rect 254 -291 255 -290
rect 387 -291 388 -290
rect 408 -291 409 -290
rect 730 -291 731 -290
rect 768 -291 769 -290
rect 905 -291 906 -290
rect 933 -291 934 -290
rect 1080 -291 1081 -290
rect 107 -293 108 -292
rect 184 -293 185 -292
rect 268 -293 269 -292
rect 289 -293 290 -292
rect 296 -293 297 -292
rect 317 -293 318 -292
rect 320 -293 321 -292
rect 639 -293 640 -292
rect 646 -293 647 -292
rect 765 -293 766 -292
rect 779 -293 780 -292
rect 877 -293 878 -292
rect 884 -293 885 -292
rect 1094 -293 1095 -292
rect 107 -295 108 -294
rect 275 -295 276 -294
rect 303 -295 304 -294
rect 373 -295 374 -294
rect 387 -295 388 -294
rect 534 -295 535 -294
rect 548 -295 549 -294
rect 593 -295 594 -294
rect 597 -295 598 -294
rect 744 -295 745 -294
rect 751 -295 752 -294
rect 884 -295 885 -294
rect 891 -295 892 -294
rect 1045 -295 1046 -294
rect 114 -297 115 -296
rect 548 -297 549 -296
rect 562 -297 563 -296
rect 597 -297 598 -296
rect 625 -297 626 -296
rect 646 -297 647 -296
rect 702 -297 703 -296
rect 828 -297 829 -296
rect 831 -297 832 -296
rect 996 -297 997 -296
rect 1003 -297 1004 -296
rect 1171 -297 1172 -296
rect 135 -299 136 -298
rect 198 -299 199 -298
rect 247 -299 248 -298
rect 268 -299 269 -298
rect 275 -299 276 -298
rect 422 -299 423 -298
rect 471 -299 472 -298
rect 779 -299 780 -298
rect 786 -299 787 -298
rect 1059 -299 1060 -298
rect 131 -301 132 -300
rect 135 -301 136 -300
rect 177 -301 178 -300
rect 408 -301 409 -300
rect 415 -301 416 -300
rect 562 -301 563 -300
rect 569 -301 570 -300
rect 625 -301 626 -300
rect 632 -301 633 -300
rect 737 -301 738 -300
rect 772 -301 773 -300
rect 891 -301 892 -300
rect 940 -301 941 -300
rect 996 -301 997 -300
rect 1010 -301 1011 -300
rect 1199 -301 1200 -300
rect 177 -303 178 -302
rect 495 -303 496 -302
rect 499 -303 500 -302
rect 534 -303 535 -302
rect 569 -303 570 -302
rect 800 -303 801 -302
rect 807 -303 808 -302
rect 1073 -303 1074 -302
rect 236 -305 237 -304
rect 940 -305 941 -304
rect 968 -305 969 -304
rect 1157 -305 1158 -304
rect 303 -307 304 -306
rect 478 -307 479 -306
rect 513 -307 514 -306
rect 1010 -307 1011 -306
rect 1017 -307 1018 -306
rect 1234 -307 1235 -306
rect 114 -309 115 -308
rect 478 -309 479 -308
rect 520 -309 521 -308
rect 751 -309 752 -308
rect 793 -309 794 -308
rect 912 -309 913 -308
rect 968 -309 969 -308
rect 1122 -309 1123 -308
rect 317 -311 318 -310
rect 352 -311 353 -310
rect 366 -311 367 -310
rect 422 -311 423 -310
rect 464 -311 465 -310
rect 499 -311 500 -310
rect 520 -311 521 -310
rect 527 -311 528 -310
rect 576 -311 577 -310
rect 793 -311 794 -310
rect 814 -311 815 -310
rect 905 -311 906 -310
rect 961 -311 962 -310
rect 1122 -311 1123 -310
rect 310 -313 311 -312
rect 352 -313 353 -312
rect 404 -313 405 -312
rect 961 -313 962 -312
rect 975 -313 976 -312
rect 1164 -313 1165 -312
rect 310 -315 311 -314
rect 324 -315 325 -314
rect 485 -315 486 -314
rect 814 -315 815 -314
rect 821 -315 822 -314
rect 849 -315 850 -314
rect 863 -315 864 -314
rect 933 -315 934 -314
rect 982 -315 983 -314
rect 1192 -315 1193 -314
rect 324 -317 325 -316
rect 331 -317 332 -316
rect 527 -317 528 -316
rect 1220 -317 1221 -316
rect 583 -319 584 -318
rect 1101 -319 1102 -318
rect 632 -321 633 -320
rect 1108 -321 1109 -320
rect 586 -323 587 -322
rect 1108 -323 1109 -322
rect 586 -325 587 -324
rect 975 -325 976 -324
rect 989 -325 990 -324
rect 1255 -325 1256 -324
rect 639 -327 640 -326
rect 667 -327 668 -326
rect 674 -327 675 -326
rect 821 -327 822 -326
rect 835 -327 836 -326
rect 1129 -327 1130 -326
rect 607 -329 608 -328
rect 835 -329 836 -328
rect 842 -329 843 -328
rect 1115 -329 1116 -328
rect 611 -331 612 -330
rect 674 -331 675 -330
rect 684 -331 685 -330
rect 807 -331 808 -330
rect 870 -331 871 -330
rect 1003 -331 1004 -330
rect 1024 -331 1025 -330
rect 1248 -331 1249 -330
rect 72 -333 73 -332
rect 611 -333 612 -332
rect 618 -333 619 -332
rect 667 -333 668 -332
rect 688 -333 689 -332
rect 870 -333 871 -332
rect 919 -333 920 -332
rect 1115 -333 1116 -332
rect 450 -335 451 -334
rect 618 -335 619 -334
rect 653 -335 654 -334
rect 688 -335 689 -334
rect 695 -335 696 -334
rect 863 -335 864 -334
rect 926 -335 927 -334
rect 1101 -335 1102 -334
rect 226 -337 227 -336
rect 695 -337 696 -336
rect 709 -337 710 -336
rect 1017 -337 1018 -336
rect 226 -339 227 -338
rect 341 -339 342 -338
rect 446 -339 447 -338
rect 450 -339 451 -338
rect 488 -339 489 -338
rect 919 -339 920 -338
rect 555 -341 556 -340
rect 653 -341 654 -340
rect 660 -341 661 -340
rect 702 -341 703 -340
rect 719 -341 720 -340
rect 982 -341 983 -340
rect 394 -343 395 -342
rect 555 -343 556 -342
rect 590 -343 591 -342
rect 709 -343 710 -342
rect 723 -343 724 -342
rect 800 -343 801 -342
rect 845 -343 846 -342
rect 1024 -343 1025 -342
rect 173 -345 174 -344
rect 394 -345 395 -344
rect 590 -345 591 -344
rect 1213 -345 1214 -344
rect 758 -347 759 -346
rect 989 -347 990 -346
rect 380 -349 381 -348
rect 758 -349 759 -348
rect 786 -349 787 -348
rect 926 -349 927 -348
rect 170 -351 171 -350
rect 380 -351 381 -350
rect 51 -353 52 -352
rect 170 -353 171 -352
rect 58 -364 59 -363
rect 1059 -364 1060 -363
rect 1227 -364 1228 -363
rect 1311 -364 1312 -363
rect 1332 -364 1333 -363
rect 1374 -364 1375 -363
rect 65 -366 66 -365
rect 338 -366 339 -365
rect 366 -366 367 -365
rect 541 -366 542 -365
rect 558 -366 559 -365
rect 891 -366 892 -365
rect 919 -366 920 -365
rect 1318 -366 1319 -365
rect 79 -368 80 -367
rect 82 -368 83 -367
rect 96 -368 97 -367
rect 975 -368 976 -367
rect 1038 -368 1039 -367
rect 1297 -368 1298 -367
rect 1300 -368 1301 -367
rect 1304 -368 1305 -367
rect 114 -370 115 -369
rect 474 -370 475 -369
rect 485 -370 486 -369
rect 758 -370 759 -369
rect 786 -370 787 -369
rect 1171 -370 1172 -369
rect 1234 -370 1235 -369
rect 1325 -370 1326 -369
rect 124 -372 125 -371
rect 128 -372 129 -371
rect 149 -372 150 -371
rect 159 -372 160 -371
rect 163 -372 164 -371
rect 261 -372 262 -371
rect 296 -372 297 -371
rect 516 -372 517 -371
rect 530 -372 531 -371
rect 863 -372 864 -371
rect 891 -372 892 -371
rect 954 -372 955 -371
rect 996 -372 997 -371
rect 1171 -372 1172 -371
rect 1248 -372 1249 -371
rect 1339 -372 1340 -371
rect 128 -374 129 -373
rect 303 -374 304 -373
rect 310 -374 311 -373
rect 537 -374 538 -373
rect 565 -374 566 -373
rect 1143 -374 1144 -373
rect 1157 -374 1158 -373
rect 1248 -374 1249 -373
rect 1255 -374 1256 -373
rect 1346 -374 1347 -373
rect 152 -376 153 -375
rect 173 -376 174 -375
rect 184 -376 185 -375
rect 359 -376 360 -375
rect 380 -376 381 -375
rect 464 -376 465 -375
rect 488 -376 489 -375
rect 1087 -376 1088 -375
rect 1136 -376 1137 -375
rect 1234 -376 1235 -375
rect 1262 -376 1263 -375
rect 1353 -376 1354 -375
rect 163 -378 164 -377
rect 625 -378 626 -377
rect 677 -378 678 -377
rect 1073 -378 1074 -377
rect 1087 -378 1088 -377
rect 1213 -378 1214 -377
rect 1276 -378 1277 -377
rect 1360 -378 1361 -377
rect 170 -380 171 -379
rect 1241 -380 1242 -379
rect 1290 -380 1291 -379
rect 1367 -380 1368 -379
rect 170 -382 171 -381
rect 191 -382 192 -381
rect 198 -382 199 -381
rect 485 -382 486 -381
rect 513 -382 514 -381
rect 793 -382 794 -381
rect 800 -382 801 -381
rect 803 -382 804 -381
rect 831 -382 832 -381
rect 1003 -382 1004 -381
rect 1024 -382 1025 -381
rect 1073 -382 1074 -381
rect 1115 -382 1116 -381
rect 1213 -382 1214 -381
rect 184 -384 185 -383
rect 226 -384 227 -383
rect 247 -384 248 -383
rect 502 -384 503 -383
rect 516 -384 517 -383
rect 1227 -384 1228 -383
rect 191 -386 192 -385
rect 562 -386 563 -385
rect 579 -386 580 -385
rect 1283 -386 1284 -385
rect 198 -388 199 -387
rect 205 -388 206 -387
rect 219 -388 220 -387
rect 492 -388 493 -387
rect 534 -388 535 -387
rect 541 -388 542 -387
rect 562 -388 563 -387
rect 597 -388 598 -387
rect 604 -388 605 -387
rect 723 -388 724 -387
rect 726 -388 727 -387
rect 1122 -388 1123 -387
rect 1150 -388 1151 -387
rect 1241 -388 1242 -387
rect 124 -390 125 -389
rect 604 -390 605 -389
rect 607 -390 608 -389
rect 1059 -390 1060 -389
rect 1066 -390 1067 -389
rect 1136 -390 1137 -389
rect 1164 -390 1165 -389
rect 1262 -390 1263 -389
rect 135 -392 136 -391
rect 205 -392 206 -391
rect 219 -392 220 -391
rect 635 -392 636 -391
rect 684 -392 685 -391
rect 1080 -392 1081 -391
rect 1122 -392 1123 -391
rect 1178 -392 1179 -391
rect 1185 -392 1186 -391
rect 1276 -392 1277 -391
rect 135 -394 136 -393
rect 730 -394 731 -393
rect 754 -394 755 -393
rect 1220 -394 1221 -393
rect 226 -396 227 -395
rect 408 -396 409 -395
rect 457 -396 458 -395
rect 614 -396 615 -395
rect 632 -396 633 -395
rect 793 -396 794 -395
rect 800 -396 801 -395
rect 842 -396 843 -395
rect 849 -396 850 -395
rect 1066 -396 1067 -395
rect 1094 -396 1095 -395
rect 1185 -396 1186 -395
rect 1192 -396 1193 -395
rect 1283 -396 1284 -395
rect 296 -398 297 -397
rect 513 -398 514 -397
rect 576 -398 577 -397
rect 1164 -398 1165 -397
rect 1206 -398 1207 -397
rect 1290 -398 1291 -397
rect 303 -400 304 -399
rect 345 -400 346 -399
rect 373 -400 374 -399
rect 408 -400 409 -399
rect 481 -400 482 -399
rect 1080 -400 1081 -399
rect 1101 -400 1102 -399
rect 1192 -400 1193 -399
rect 310 -402 311 -401
rect 663 -402 664 -401
rect 716 -402 717 -401
rect 863 -402 864 -401
rect 898 -402 899 -401
rect 1255 -402 1256 -401
rect 324 -404 325 -403
rect 478 -404 479 -403
rect 576 -404 577 -403
rect 814 -404 815 -403
rect 828 -404 829 -403
rect 898 -404 899 -403
rect 905 -404 906 -403
rect 1150 -404 1151 -403
rect 107 -406 108 -405
rect 478 -406 479 -405
rect 579 -406 580 -405
rect 1206 -406 1207 -405
rect 107 -408 108 -407
rect 233 -408 234 -407
rect 289 -408 290 -407
rect 324 -408 325 -407
rect 331 -408 332 -407
rect 527 -408 528 -407
rect 583 -408 584 -407
rect 775 -408 776 -407
rect 803 -408 804 -407
rect 842 -408 843 -407
rect 849 -408 850 -407
rect 989 -408 990 -407
rect 1031 -408 1032 -407
rect 1038 -408 1039 -407
rect 1052 -408 1053 -407
rect 1094 -408 1095 -407
rect 1101 -408 1102 -407
rect 1199 -408 1200 -407
rect 177 -410 178 -409
rect 527 -410 528 -409
rect 583 -410 584 -409
rect 716 -410 717 -409
rect 719 -410 720 -409
rect 954 -410 955 -409
rect 968 -410 969 -409
rect 1003 -410 1004 -409
rect 1010 -410 1011 -409
rect 1052 -410 1053 -409
rect 1108 -410 1109 -409
rect 1199 -410 1200 -409
rect 156 -412 157 -411
rect 1108 -412 1109 -411
rect 131 -414 132 -413
rect 156 -414 157 -413
rect 177 -414 178 -413
rect 467 -414 468 -413
rect 586 -414 587 -413
rect 884 -414 885 -413
rect 912 -414 913 -413
rect 1143 -414 1144 -413
rect 233 -416 234 -415
rect 709 -416 710 -415
rect 723 -416 724 -415
rect 884 -416 885 -415
rect 926 -416 927 -415
rect 989 -416 990 -415
rect 338 -418 339 -417
rect 457 -418 458 -417
rect 520 -418 521 -417
rect 912 -418 913 -417
rect 940 -418 941 -417
rect 996 -418 997 -417
rect 345 -420 346 -419
rect 443 -420 444 -419
rect 506 -420 507 -419
rect 520 -420 521 -419
rect 597 -420 598 -419
rect 1045 -420 1046 -419
rect 149 -422 150 -421
rect 1045 -422 1046 -421
rect 373 -424 374 -423
rect 681 -424 682 -423
rect 702 -424 703 -423
rect 814 -424 815 -423
rect 835 -424 836 -423
rect 905 -424 906 -423
rect 982 -424 983 -423
rect 1024 -424 1025 -423
rect 380 -426 381 -425
rect 436 -426 437 -425
rect 611 -426 612 -425
rect 625 -426 626 -425
rect 632 -426 633 -425
rect 1017 -426 1018 -425
rect 387 -428 388 -427
rect 506 -428 507 -427
rect 635 -428 636 -427
rect 1269 -428 1270 -427
rect 352 -430 353 -429
rect 387 -430 388 -429
rect 394 -430 395 -429
rect 572 -430 573 -429
rect 642 -430 643 -429
rect 1010 -430 1011 -429
rect 72 -432 73 -431
rect 394 -432 395 -431
rect 401 -432 402 -431
rect 975 -432 976 -431
rect 72 -434 73 -433
rect 86 -434 87 -433
rect 100 -434 101 -433
rect 352 -434 353 -433
rect 401 -434 402 -433
rect 499 -434 500 -433
rect 660 -434 661 -433
rect 1178 -434 1179 -433
rect 86 -436 87 -435
rect 212 -436 213 -435
rect 422 -436 423 -435
rect 436 -436 437 -435
rect 499 -436 500 -435
rect 555 -436 556 -435
rect 660 -436 661 -435
rect 674 -436 675 -435
rect 684 -436 685 -435
rect 1269 -436 1270 -435
rect 100 -438 101 -437
rect 275 -438 276 -437
rect 415 -438 416 -437
rect 422 -438 423 -437
rect 429 -438 430 -437
rect 443 -438 444 -437
rect 555 -438 556 -437
rect 1115 -438 1116 -437
rect 212 -440 213 -439
rect 961 -440 962 -439
rect 254 -442 255 -441
rect 429 -442 430 -441
rect 667 -442 668 -441
rect 709 -442 710 -441
rect 730 -442 731 -441
rect 765 -442 766 -441
rect 772 -442 773 -441
rect 940 -442 941 -441
rect 947 -442 948 -441
rect 961 -442 962 -441
rect 254 -444 255 -443
rect 471 -444 472 -443
rect 534 -444 535 -443
rect 947 -444 948 -443
rect 317 -446 318 -445
rect 415 -446 416 -445
rect 667 -446 668 -445
rect 821 -446 822 -445
rect 870 -446 871 -445
rect 926 -446 927 -445
rect 933 -446 934 -445
rect 982 -446 983 -445
rect 268 -448 269 -447
rect 317 -448 318 -447
rect 355 -448 356 -447
rect 471 -448 472 -447
rect 590 -448 591 -447
rect 870 -448 871 -447
rect 877 -448 878 -447
rect 933 -448 934 -447
rect 93 -450 94 -449
rect 268 -450 269 -449
rect 590 -450 591 -449
rect 653 -450 654 -449
rect 688 -450 689 -449
rect 877 -450 878 -449
rect 887 -450 888 -449
rect 1017 -450 1018 -449
rect 51 -452 52 -451
rect 688 -452 689 -451
rect 702 -452 703 -451
rect 737 -452 738 -451
rect 744 -452 745 -451
rect 765 -452 766 -451
rect 789 -452 790 -451
rect 835 -452 836 -451
rect 569 -454 570 -453
rect 653 -454 654 -453
rect 674 -454 675 -453
rect 737 -454 738 -453
rect 751 -454 752 -453
rect 1031 -454 1032 -453
rect 142 -456 143 -455
rect 569 -456 570 -455
rect 695 -456 696 -455
rect 744 -456 745 -455
rect 758 -456 759 -455
rect 968 -456 969 -455
rect 142 -458 143 -457
rect 215 -458 216 -457
rect 695 -458 696 -457
rect 1157 -458 1158 -457
rect 789 -460 790 -459
rect 919 -460 920 -459
rect 807 -462 808 -461
rect 1220 -462 1221 -461
rect 779 -464 780 -463
rect 807 -464 808 -463
rect 821 -464 822 -463
rect 856 -464 857 -463
rect 639 -466 640 -465
rect 779 -466 780 -465
rect 639 -468 640 -467
rect 1129 -468 1130 -467
rect 611 -470 612 -469
rect 1129 -470 1130 -469
rect 646 -472 647 -471
rect 856 -472 857 -471
rect 618 -474 619 -473
rect 646 -474 647 -473
rect 450 -476 451 -475
rect 618 -476 619 -475
rect 450 -478 451 -477
rect 460 -478 461 -477
rect 58 -489 59 -488
rect 590 -489 591 -488
rect 611 -489 612 -488
rect 1297 -489 1298 -488
rect 1377 -489 1378 -488
rect 1381 -489 1382 -488
rect 65 -491 66 -490
rect 275 -491 276 -490
rect 310 -491 311 -490
rect 355 -491 356 -490
rect 373 -491 374 -490
rect 600 -491 601 -490
rect 625 -491 626 -490
rect 695 -491 696 -490
rect 698 -491 699 -490
rect 1318 -491 1319 -490
rect 51 -493 52 -492
rect 65 -493 66 -492
rect 68 -493 69 -492
rect 205 -493 206 -492
rect 212 -493 213 -492
rect 219 -493 220 -492
rect 233 -493 234 -492
rect 761 -493 762 -492
rect 768 -493 769 -492
rect 1325 -493 1326 -492
rect 72 -495 73 -494
rect 96 -495 97 -494
rect 114 -495 115 -494
rect 128 -495 129 -494
rect 131 -495 132 -494
rect 282 -495 283 -494
rect 338 -495 339 -494
rect 789 -495 790 -494
rect 831 -495 832 -494
rect 1283 -495 1284 -494
rect 1325 -495 1326 -494
rect 1353 -495 1354 -494
rect 72 -497 73 -496
rect 79 -497 80 -496
rect 124 -497 125 -496
rect 506 -497 507 -496
rect 513 -497 514 -496
rect 975 -497 976 -496
rect 978 -497 979 -496
rect 1283 -497 1284 -496
rect 128 -499 129 -498
rect 247 -499 248 -498
rect 254 -499 255 -498
rect 544 -499 545 -498
rect 569 -499 570 -498
rect 810 -499 811 -498
rect 884 -499 885 -498
rect 1367 -499 1368 -498
rect 152 -501 153 -500
rect 170 -501 171 -500
rect 177 -501 178 -500
rect 338 -501 339 -500
rect 373 -501 374 -500
rect 775 -501 776 -500
rect 782 -501 783 -500
rect 1143 -501 1144 -500
rect 152 -503 153 -502
rect 184 -503 185 -502
rect 198 -503 199 -502
rect 205 -503 206 -502
rect 215 -503 216 -502
rect 912 -503 913 -502
rect 954 -503 955 -502
rect 1143 -503 1144 -502
rect 156 -505 157 -504
rect 579 -505 580 -504
rect 586 -505 587 -504
rect 877 -505 878 -504
rect 887 -505 888 -504
rect 1388 -505 1389 -504
rect 163 -507 164 -506
rect 625 -507 626 -506
rect 646 -507 647 -506
rect 670 -507 671 -506
rect 688 -507 689 -506
rect 884 -507 885 -506
rect 891 -507 892 -506
rect 1374 -507 1375 -506
rect 163 -509 164 -508
rect 408 -509 409 -508
rect 460 -509 461 -508
rect 856 -509 857 -508
rect 870 -509 871 -508
rect 1367 -509 1368 -508
rect 156 -511 157 -510
rect 870 -511 871 -510
rect 912 -511 913 -510
rect 926 -511 927 -510
rect 968 -511 969 -510
rect 1318 -511 1319 -510
rect 177 -513 178 -512
rect 639 -513 640 -512
rect 688 -513 689 -512
rect 779 -513 780 -512
rect 786 -513 787 -512
rect 1213 -513 1214 -512
rect 184 -515 185 -514
rect 653 -515 654 -514
rect 705 -515 706 -514
rect 1031 -515 1032 -514
rect 1045 -515 1046 -514
rect 1472 -515 1473 -514
rect 219 -517 220 -516
rect 478 -517 479 -516
rect 499 -517 500 -516
rect 989 -517 990 -516
rect 1045 -517 1046 -516
rect 1353 -517 1354 -516
rect 222 -519 223 -518
rect 968 -519 969 -518
rect 989 -519 990 -518
rect 1003 -519 1004 -518
rect 1087 -519 1088 -518
rect 1297 -519 1298 -518
rect 240 -521 241 -520
rect 289 -521 290 -520
rect 296 -521 297 -520
rect 646 -521 647 -520
rect 653 -521 654 -520
rect 737 -521 738 -520
rect 754 -521 755 -520
rect 1059 -521 1060 -520
rect 1178 -521 1179 -520
rect 1213 -521 1214 -520
rect 243 -523 244 -522
rect 611 -523 612 -522
rect 614 -523 615 -522
rect 1059 -523 1060 -522
rect 1178 -523 1179 -522
rect 1234 -523 1235 -522
rect 268 -525 269 -524
rect 310 -525 311 -524
rect 380 -525 381 -524
rect 506 -525 507 -524
rect 513 -525 514 -524
rect 667 -525 668 -524
rect 716 -525 717 -524
rect 1255 -525 1256 -524
rect 268 -527 269 -526
rect 331 -527 332 -526
rect 359 -527 360 -526
rect 716 -527 717 -526
rect 719 -527 720 -526
rect 1150 -527 1151 -526
rect 1248 -527 1249 -526
rect 1255 -527 1256 -526
rect 107 -529 108 -528
rect 359 -529 360 -528
rect 397 -529 398 -528
rect 681 -529 682 -528
rect 737 -529 738 -528
rect 744 -529 745 -528
rect 751 -529 752 -528
rect 1234 -529 1235 -528
rect 1241 -529 1242 -528
rect 1248 -529 1249 -528
rect 107 -531 108 -530
rect 828 -531 829 -530
rect 835 -531 836 -530
rect 877 -531 878 -530
rect 901 -531 902 -530
rect 1031 -531 1032 -530
rect 1150 -531 1151 -530
rect 1164 -531 1165 -530
rect 159 -533 160 -532
rect 1241 -533 1242 -532
rect 296 -535 297 -534
rect 401 -535 402 -534
rect 408 -535 409 -534
rect 415 -535 416 -534
rect 499 -535 500 -534
rect 891 -535 892 -534
rect 926 -535 927 -534
rect 1080 -535 1081 -534
rect 1164 -535 1165 -534
rect 1171 -535 1172 -534
rect 317 -537 318 -536
rect 380 -537 381 -536
rect 401 -537 402 -536
rect 632 -537 633 -536
rect 733 -537 734 -536
rect 751 -537 752 -536
rect 772 -537 773 -536
rect 1017 -537 1018 -536
rect 1073 -537 1074 -536
rect 1080 -537 1081 -536
rect 1171 -537 1172 -536
rect 1185 -537 1186 -536
rect 303 -539 304 -538
rect 317 -539 318 -538
rect 324 -539 325 -538
rect 331 -539 332 -538
rect 366 -539 367 -538
rect 744 -539 745 -538
rect 786 -539 787 -538
rect 800 -539 801 -538
rect 814 -539 815 -538
rect 828 -539 829 -538
rect 835 -539 836 -538
rect 842 -539 843 -538
rect 856 -539 857 -538
rect 1052 -539 1053 -538
rect 1073 -539 1074 -538
rect 1108 -539 1109 -538
rect 1185 -539 1186 -538
rect 1199 -539 1200 -538
rect 261 -541 262 -540
rect 303 -541 304 -540
rect 324 -541 325 -540
rect 387 -541 388 -540
rect 415 -541 416 -540
rect 443 -541 444 -540
rect 502 -541 503 -540
rect 793 -541 794 -540
rect 821 -541 822 -540
rect 842 -541 843 -540
rect 919 -541 920 -540
rect 1017 -541 1018 -540
rect 1108 -541 1109 -540
rect 1192 -541 1193 -540
rect 387 -543 388 -542
rect 457 -543 458 -542
rect 502 -543 503 -542
rect 1276 -543 1277 -542
rect 443 -545 444 -544
rect 618 -545 619 -544
rect 674 -545 675 -544
rect 1052 -545 1053 -544
rect 1101 -545 1102 -544
rect 1192 -545 1193 -544
rect 1276 -545 1277 -544
rect 1304 -545 1305 -544
rect 450 -547 451 -546
rect 457 -547 458 -546
rect 492 -547 493 -546
rect 618 -547 619 -546
rect 660 -547 661 -546
rect 674 -547 675 -546
rect 730 -547 731 -546
rect 800 -547 801 -546
rect 807 -547 808 -546
rect 821 -547 822 -546
rect 919 -547 920 -546
rect 996 -547 997 -546
rect 1003 -547 1004 -546
rect 1024 -547 1025 -546
rect 1094 -547 1095 -546
rect 1101 -547 1102 -546
rect 1115 -547 1116 -546
rect 1199 -547 1200 -546
rect 1304 -547 1305 -546
rect 1311 -547 1312 -546
rect 121 -549 122 -548
rect 1115 -549 1116 -548
rect 1311 -549 1312 -548
rect 1339 -549 1340 -548
rect 121 -551 122 -550
rect 530 -551 531 -550
rect 534 -551 535 -550
rect 562 -551 563 -550
rect 590 -551 591 -550
rect 597 -551 598 -550
rect 604 -551 605 -550
rect 954 -551 955 -550
rect 975 -551 976 -550
rect 1087 -551 1088 -550
rect 1094 -551 1095 -550
rect 1129 -551 1130 -550
rect 1332 -551 1333 -550
rect 1339 -551 1340 -550
rect 93 -553 94 -552
rect 1332 -553 1333 -552
rect 142 -555 143 -554
rect 597 -555 598 -554
rect 635 -555 636 -554
rect 1129 -555 1130 -554
rect 135 -557 136 -556
rect 142 -557 143 -556
rect 394 -557 395 -556
rect 534 -557 535 -556
rect 537 -557 538 -556
rect 898 -557 899 -556
rect 940 -557 941 -556
rect 996 -557 997 -556
rect 135 -559 136 -558
rect 1262 -559 1263 -558
rect 149 -561 150 -560
rect 940 -561 941 -560
rect 149 -563 150 -562
rect 695 -563 696 -562
rect 779 -563 780 -562
rect 1262 -563 1263 -562
rect 191 -565 192 -564
rect 394 -565 395 -564
rect 429 -565 430 -564
rect 604 -565 605 -564
rect 639 -565 640 -564
rect 730 -565 731 -564
rect 793 -565 794 -564
rect 1269 -565 1270 -564
rect 191 -567 192 -566
rect 485 -567 486 -566
rect 492 -567 493 -566
rect 583 -567 584 -566
rect 660 -567 661 -566
rect 684 -567 685 -566
rect 1269 -567 1270 -566
rect 1290 -567 1291 -566
rect 345 -569 346 -568
rect 429 -569 430 -568
rect 436 -569 437 -568
rect 450 -569 451 -568
rect 471 -569 472 -568
rect 562 -569 563 -568
rect 583 -569 584 -568
rect 632 -569 633 -568
rect 1290 -569 1291 -568
rect 1360 -569 1361 -568
rect 198 -571 199 -570
rect 1360 -571 1361 -570
rect 250 -573 251 -572
rect 345 -573 346 -572
rect 352 -573 353 -572
rect 684 -573 685 -572
rect 422 -575 423 -574
rect 436 -575 437 -574
rect 464 -575 465 -574
rect 471 -575 472 -574
rect 485 -575 486 -574
rect 702 -575 703 -574
rect 100 -577 101 -576
rect 464 -577 465 -576
rect 478 -577 479 -576
rect 702 -577 703 -576
rect 86 -579 87 -578
rect 100 -579 101 -578
rect 422 -579 423 -578
rect 520 -579 521 -578
rect 527 -579 528 -578
rect 576 -579 577 -578
rect 79 -581 80 -580
rect 86 -581 87 -580
rect 520 -581 521 -580
rect 723 -581 724 -580
rect 527 -583 528 -582
rect 814 -583 815 -582
rect 548 -585 549 -584
rect 569 -585 570 -584
rect 723 -585 724 -584
rect 905 -585 906 -584
rect 226 -587 227 -586
rect 548 -587 549 -586
rect 555 -587 556 -586
rect 898 -587 899 -586
rect 905 -587 906 -586
rect 947 -587 948 -586
rect 40 -589 41 -588
rect 226 -589 227 -588
rect 541 -589 542 -588
rect 555 -589 556 -588
rect 947 -589 948 -588
rect 1010 -589 1011 -588
rect 40 -591 41 -590
rect 261 -591 262 -590
rect 541 -591 542 -590
rect 1220 -591 1221 -590
rect 1010 -593 1011 -592
rect 1122 -593 1123 -592
rect 1220 -593 1221 -592
rect 1227 -593 1228 -592
rect 807 -595 808 -594
rect 1227 -595 1228 -594
rect 961 -597 962 -596
rect 1122 -597 1123 -596
rect 961 -599 962 -598
rect 1066 -599 1067 -598
rect 1066 -601 1067 -600
rect 1136 -601 1137 -600
rect 1136 -603 1137 -602
rect 1157 -603 1158 -602
rect 1038 -605 1039 -604
rect 1157 -605 1158 -604
rect 758 -607 759 -606
rect 1038 -607 1039 -606
rect 758 -609 759 -608
rect 765 -609 766 -608
rect 765 -611 766 -610
rect 1024 -611 1025 -610
rect 44 -622 45 -621
rect 292 -622 293 -621
rect 387 -622 388 -621
rect 583 -622 584 -621
rect 649 -622 650 -621
rect 1115 -622 1116 -621
rect 1185 -622 1186 -621
rect 1395 -622 1396 -621
rect 1472 -622 1473 -621
rect 1633 -622 1634 -621
rect 51 -624 52 -623
rect 516 -624 517 -623
rect 527 -624 528 -623
rect 912 -624 913 -623
rect 975 -624 976 -623
rect 1045 -624 1046 -623
rect 1059 -624 1060 -623
rect 1185 -624 1186 -623
rect 1234 -624 1235 -623
rect 1500 -624 1501 -623
rect 51 -626 52 -625
rect 310 -626 311 -625
rect 397 -626 398 -625
rect 670 -626 671 -625
rect 684 -626 685 -625
rect 1255 -626 1256 -625
rect 1311 -626 1312 -625
rect 1409 -626 1410 -625
rect 72 -628 73 -627
rect 82 -628 83 -627
rect 107 -628 108 -627
rect 558 -628 559 -627
rect 698 -628 699 -627
rect 842 -628 843 -627
rect 887 -628 888 -627
rect 1101 -628 1102 -627
rect 1136 -628 1137 -627
rect 1234 -628 1235 -627
rect 1353 -628 1354 -627
rect 1381 -628 1382 -627
rect 1388 -628 1389 -627
rect 1570 -628 1571 -627
rect 65 -630 66 -629
rect 1101 -630 1102 -629
rect 1157 -630 1158 -629
rect 1311 -630 1312 -629
rect 1332 -630 1333 -629
rect 1381 -630 1382 -629
rect 65 -632 66 -631
rect 226 -632 227 -631
rect 233 -632 234 -631
rect 488 -632 489 -631
rect 537 -632 538 -631
rect 723 -632 724 -631
rect 730 -632 731 -631
rect 1213 -632 1214 -631
rect 1227 -632 1228 -631
rect 1255 -632 1256 -631
rect 1276 -632 1277 -631
rect 1353 -632 1354 -631
rect 1356 -632 1357 -631
rect 1367 -632 1368 -631
rect 72 -634 73 -633
rect 373 -634 374 -633
rect 429 -634 430 -633
rect 502 -634 503 -633
rect 541 -634 542 -633
rect 625 -634 626 -633
rect 702 -634 703 -633
rect 1374 -634 1375 -633
rect 82 -636 83 -635
rect 100 -636 101 -635
rect 114 -636 115 -635
rect 117 -636 118 -635
rect 128 -636 129 -635
rect 226 -636 227 -635
rect 243 -636 244 -635
rect 387 -636 388 -635
rect 432 -636 433 -635
rect 751 -636 752 -635
rect 772 -636 773 -635
rect 1339 -636 1340 -635
rect 1360 -636 1361 -635
rect 1521 -636 1522 -635
rect 86 -638 87 -637
rect 100 -638 101 -637
rect 128 -638 129 -637
rect 555 -638 556 -637
rect 702 -638 703 -637
rect 758 -638 759 -637
rect 768 -638 769 -637
rect 1360 -638 1361 -637
rect 86 -640 87 -639
rect 674 -640 675 -639
rect 705 -640 706 -639
rect 842 -640 843 -639
rect 898 -640 899 -639
rect 1010 -640 1011 -639
rect 1017 -640 1018 -639
rect 1115 -640 1116 -639
rect 1129 -640 1130 -639
rect 1227 -640 1228 -639
rect 1269 -640 1270 -639
rect 1339 -640 1340 -639
rect 138 -642 139 -641
rect 219 -642 220 -641
rect 247 -642 248 -641
rect 856 -642 857 -641
rect 863 -642 864 -641
rect 898 -642 899 -641
rect 940 -642 941 -641
rect 1010 -642 1011 -641
rect 1080 -642 1081 -641
rect 1136 -642 1137 -641
rect 1157 -642 1158 -641
rect 1164 -642 1165 -641
rect 1171 -642 1172 -641
rect 1276 -642 1277 -641
rect 1290 -642 1291 -641
rect 1388 -642 1389 -641
rect 107 -644 108 -643
rect 247 -644 248 -643
rect 250 -644 251 -643
rect 527 -644 528 -643
rect 555 -644 556 -643
rect 765 -644 766 -643
rect 772 -644 773 -643
rect 908 -644 909 -643
rect 954 -644 955 -643
rect 1045 -644 1046 -643
rect 1052 -644 1053 -643
rect 1164 -644 1165 -643
rect 1192 -644 1193 -643
rect 1332 -644 1333 -643
rect 142 -646 143 -645
rect 156 -646 157 -645
rect 159 -646 160 -645
rect 1402 -646 1403 -645
rect 149 -648 150 -647
rect 240 -648 241 -647
rect 250 -648 251 -647
rect 478 -648 479 -647
rect 485 -648 486 -647
rect 593 -648 594 -647
rect 674 -648 675 -647
rect 821 -648 822 -647
rect 831 -648 832 -647
rect 1178 -648 1179 -647
rect 1206 -648 1207 -647
rect 1269 -648 1270 -647
rect 1290 -648 1291 -647
rect 1304 -648 1305 -647
rect 1325 -648 1326 -647
rect 1374 -648 1375 -647
rect 152 -650 153 -649
rect 1199 -650 1200 -649
rect 1241 -650 1242 -649
rect 1304 -650 1305 -649
rect 156 -652 157 -651
rect 796 -652 797 -651
rect 807 -652 808 -651
rect 1346 -652 1347 -651
rect 163 -654 164 -653
rect 429 -654 430 -653
rect 443 -654 444 -653
rect 583 -654 584 -653
rect 586 -654 587 -653
rect 1199 -654 1200 -653
rect 1248 -654 1249 -653
rect 1346 -654 1347 -653
rect 163 -656 164 -655
rect 656 -656 657 -655
rect 695 -656 696 -655
rect 1129 -656 1130 -655
rect 1248 -656 1249 -655
rect 1426 -656 1427 -655
rect 58 -658 59 -657
rect 695 -658 696 -657
rect 709 -658 710 -657
rect 758 -658 759 -657
rect 775 -658 776 -657
rect 978 -658 979 -657
rect 982 -658 983 -657
rect 1052 -658 1053 -657
rect 1122 -658 1123 -657
rect 1206 -658 1207 -657
rect 58 -660 59 -659
rect 93 -660 94 -659
rect 170 -660 171 -659
rect 380 -660 381 -659
rect 415 -660 416 -659
rect 443 -660 444 -659
rect 471 -660 472 -659
rect 478 -660 479 -659
rect 565 -660 566 -659
rect 1192 -660 1193 -659
rect 187 -662 188 -661
rect 205 -662 206 -661
rect 219 -662 220 -661
rect 324 -662 325 -661
rect 345 -662 346 -661
rect 625 -662 626 -661
rect 716 -662 717 -661
rect 1325 -662 1326 -661
rect 124 -664 125 -663
rect 345 -664 346 -663
rect 373 -664 374 -663
rect 464 -664 465 -663
rect 471 -664 472 -663
rect 590 -664 591 -663
rect 607 -664 608 -663
rect 1241 -664 1242 -663
rect 149 -666 150 -665
rect 590 -666 591 -665
rect 716 -666 717 -665
rect 828 -666 829 -665
rect 856 -666 857 -665
rect 1367 -666 1368 -665
rect 201 -668 202 -667
rect 212 -668 213 -667
rect 268 -668 269 -667
rect 366 -668 367 -667
rect 380 -668 381 -667
rect 492 -668 493 -667
rect 719 -668 720 -667
rect 1094 -668 1095 -667
rect 205 -670 206 -669
rect 632 -670 633 -669
rect 723 -670 724 -669
rect 1297 -670 1298 -669
rect 212 -672 213 -671
rect 352 -672 353 -671
rect 401 -672 402 -671
rect 415 -672 416 -671
rect 464 -672 465 -671
rect 712 -672 713 -671
rect 726 -672 727 -671
rect 1017 -672 1018 -671
rect 1024 -672 1025 -671
rect 1122 -672 1123 -671
rect 268 -674 269 -673
rect 530 -674 531 -673
rect 733 -674 734 -673
rect 954 -674 955 -673
rect 961 -674 962 -673
rect 1178 -674 1179 -673
rect 275 -676 276 -675
rect 751 -676 752 -675
rect 779 -676 780 -675
rect 996 -676 997 -675
rect 1003 -676 1004 -675
rect 1213 -676 1214 -675
rect 254 -678 255 -677
rect 275 -678 276 -677
rect 282 -678 283 -677
rect 439 -678 440 -677
rect 611 -678 612 -677
rect 996 -678 997 -677
rect 1006 -678 1007 -677
rect 1143 -678 1144 -677
rect 282 -680 283 -679
rect 579 -680 580 -679
rect 737 -680 738 -679
rect 765 -680 766 -679
rect 786 -680 787 -679
rect 863 -680 864 -679
rect 877 -680 878 -679
rect 961 -680 962 -679
rect 968 -680 969 -679
rect 1080 -680 1081 -679
rect 121 -682 122 -681
rect 737 -682 738 -681
rect 744 -682 745 -681
rect 779 -682 780 -681
rect 793 -682 794 -681
rect 1416 -682 1417 -681
rect 121 -684 122 -683
rect 1073 -684 1074 -683
rect 296 -686 297 -685
rect 541 -686 542 -685
rect 646 -686 647 -685
rect 786 -686 787 -685
rect 793 -686 794 -685
rect 1318 -686 1319 -685
rect 289 -688 290 -687
rect 296 -688 297 -687
rect 310 -688 311 -687
rect 891 -688 892 -687
rect 905 -688 906 -687
rect 1024 -688 1025 -687
rect 1031 -688 1032 -687
rect 1143 -688 1144 -687
rect 1262 -688 1263 -687
rect 1318 -688 1319 -687
rect 317 -690 318 -689
rect 324 -690 325 -689
rect 352 -690 353 -689
rect 604 -690 605 -689
rect 618 -690 619 -689
rect 646 -690 647 -689
rect 733 -690 734 -689
rect 1073 -690 1074 -689
rect 1108 -690 1109 -689
rect 1262 -690 1263 -689
rect 317 -692 318 -691
rect 422 -692 423 -691
rect 513 -692 514 -691
rect 744 -692 745 -691
rect 800 -692 801 -691
rect 877 -692 878 -691
rect 884 -692 885 -691
rect 968 -692 969 -691
rect 989 -692 990 -691
rect 1094 -692 1095 -691
rect 401 -694 402 -693
rect 604 -694 605 -693
rect 660 -694 661 -693
rect 800 -694 801 -693
rect 807 -694 808 -693
rect 912 -694 913 -693
rect 933 -694 934 -693
rect 982 -694 983 -693
rect 992 -694 993 -693
rect 1150 -694 1151 -693
rect 408 -696 409 -695
rect 492 -696 493 -695
rect 513 -696 514 -695
rect 534 -696 535 -695
rect 576 -696 577 -695
rect 618 -696 619 -695
rect 660 -696 661 -695
rect 688 -696 689 -695
rect 814 -696 815 -695
rect 891 -696 892 -695
rect 905 -696 906 -695
rect 1283 -696 1284 -695
rect 68 -698 69 -697
rect 688 -698 689 -697
rect 821 -698 822 -697
rect 835 -698 836 -697
rect 884 -698 885 -697
rect 926 -698 927 -697
rect 1031 -698 1032 -697
rect 1059 -698 1060 -697
rect 1062 -698 1063 -697
rect 1297 -698 1298 -697
rect 96 -700 97 -699
rect 814 -700 815 -699
rect 828 -700 829 -699
rect 940 -700 941 -699
rect 1038 -700 1039 -699
rect 1171 -700 1172 -699
rect 1220 -700 1221 -699
rect 1283 -700 1284 -699
rect 135 -702 136 -701
rect 1038 -702 1039 -701
rect 1066 -702 1067 -701
rect 1108 -702 1109 -701
rect 135 -704 136 -703
rect 261 -704 262 -703
rect 359 -704 360 -703
rect 408 -704 409 -703
rect 422 -704 423 -703
rect 436 -704 437 -703
rect 520 -704 521 -703
rect 611 -704 612 -703
rect 667 -704 668 -703
rect 933 -704 934 -703
rect 1087 -704 1088 -703
rect 1220 -704 1221 -703
rect 184 -706 185 -705
rect 261 -706 262 -705
rect 359 -706 360 -705
rect 653 -706 654 -705
rect 667 -706 668 -705
rect 859 -706 860 -705
rect 870 -706 871 -705
rect 926 -706 927 -705
rect 947 -706 948 -705
rect 1087 -706 1088 -705
rect 436 -708 437 -707
rect 1150 -708 1151 -707
rect 520 -710 521 -709
rect 597 -710 598 -709
rect 653 -710 654 -709
rect 681 -710 682 -709
rect 835 -710 836 -709
rect 901 -710 902 -709
rect 919 -710 920 -709
rect 1066 -710 1067 -709
rect 534 -712 535 -711
rect 569 -712 570 -711
rect 849 -712 850 -711
rect 947 -712 948 -711
rect 548 -714 549 -713
rect 569 -714 570 -713
rect 709 -714 710 -713
rect 849 -714 850 -713
rect 919 -714 920 -713
rect 1430 -714 1431 -713
rect 548 -716 549 -715
rect 639 -716 640 -715
rect 394 -718 395 -717
rect 639 -718 640 -717
rect 177 -720 178 -719
rect 394 -720 395 -719
rect 562 -720 563 -719
rect 597 -720 598 -719
rect 177 -722 178 -721
rect 506 -722 507 -721
rect 191 -724 192 -723
rect 506 -724 507 -723
rect 191 -726 192 -725
rect 338 -726 339 -725
rect 303 -728 304 -727
rect 562 -728 563 -727
rect 303 -730 304 -729
rect 576 -730 577 -729
rect 331 -732 332 -731
rect 338 -732 339 -731
rect 184 -734 185 -733
rect 331 -734 332 -733
rect 37 -745 38 -744
rect 58 -745 59 -744
rect 79 -745 80 -744
rect 919 -745 920 -744
rect 922 -745 923 -744
rect 1402 -745 1403 -744
rect 1416 -745 1417 -744
rect 1608 -745 1609 -744
rect 1633 -745 1634 -744
rect 1696 -745 1697 -744
rect 44 -747 45 -746
rect 1556 -747 1557 -746
rect 1570 -747 1571 -746
rect 1626 -747 1627 -746
rect 44 -749 45 -748
rect 450 -749 451 -748
rect 467 -749 468 -748
rect 1437 -749 1438 -748
rect 1500 -749 1501 -748
rect 1619 -749 1620 -748
rect 58 -751 59 -750
rect 149 -751 150 -750
rect 166 -751 167 -750
rect 1458 -751 1459 -750
rect 1521 -751 1522 -750
rect 1591 -751 1592 -750
rect 1605 -751 1606 -750
rect 1612 -751 1613 -750
rect 82 -753 83 -752
rect 604 -753 605 -752
rect 607 -753 608 -752
rect 877 -753 878 -752
rect 884 -753 885 -752
rect 1521 -753 1522 -752
rect 93 -755 94 -754
rect 800 -755 801 -754
rect 821 -755 822 -754
rect 884 -755 885 -754
rect 905 -755 906 -754
rect 1346 -755 1347 -754
rect 1353 -755 1354 -754
rect 1549 -755 1550 -754
rect 93 -757 94 -756
rect 527 -757 528 -756
rect 537 -757 538 -756
rect 723 -757 724 -756
rect 730 -757 731 -756
rect 779 -757 780 -756
rect 782 -757 783 -756
rect 1220 -757 1221 -756
rect 1241 -757 1242 -756
rect 1416 -757 1417 -756
rect 1430 -757 1431 -756
rect 1633 -757 1634 -756
rect 33 -759 34 -758
rect 527 -759 528 -758
rect 558 -759 559 -758
rect 1507 -759 1508 -758
rect 103 -761 104 -760
rect 366 -761 367 -760
rect 485 -761 486 -760
rect 562 -761 563 -760
rect 565 -761 566 -760
rect 1094 -761 1095 -760
rect 1122 -761 1123 -760
rect 1542 -761 1543 -760
rect 124 -763 125 -762
rect 1570 -763 1571 -762
rect 128 -765 129 -764
rect 131 -765 132 -764
rect 138 -765 139 -764
rect 1360 -765 1361 -764
rect 1367 -765 1368 -764
rect 1577 -765 1578 -764
rect 128 -767 129 -766
rect 618 -767 619 -766
rect 632 -767 633 -766
rect 639 -767 640 -766
rect 649 -767 650 -766
rect 1367 -767 1368 -766
rect 1374 -767 1375 -766
rect 1584 -767 1585 -766
rect 142 -769 143 -768
rect 726 -769 727 -768
rect 730 -769 731 -768
rect 758 -769 759 -768
rect 765 -769 766 -768
rect 821 -769 822 -768
rect 828 -769 829 -768
rect 961 -769 962 -768
rect 1003 -769 1004 -768
rect 1426 -769 1427 -768
rect 149 -771 150 -770
rect 625 -771 626 -770
rect 628 -771 629 -770
rect 1374 -771 1375 -770
rect 1388 -771 1389 -770
rect 1514 -771 1515 -770
rect 184 -773 185 -772
rect 1493 -773 1494 -772
rect 184 -775 185 -774
rect 198 -775 199 -774
rect 205 -775 206 -774
rect 450 -775 451 -774
rect 488 -775 489 -774
rect 555 -775 556 -774
rect 576 -775 577 -774
rect 716 -775 717 -774
rect 733 -775 734 -774
rect 1423 -775 1424 -774
rect 187 -777 188 -776
rect 1213 -777 1214 -776
rect 1227 -777 1228 -776
rect 1388 -777 1389 -776
rect 191 -779 192 -778
rect 236 -779 237 -778
rect 240 -779 241 -778
rect 366 -779 367 -778
rect 471 -779 472 -778
rect 555 -779 556 -778
rect 576 -779 577 -778
rect 863 -779 864 -778
rect 870 -779 871 -778
rect 1444 -779 1445 -778
rect 191 -781 192 -780
rect 429 -781 430 -780
rect 471 -781 472 -780
rect 478 -781 479 -780
rect 499 -781 500 -780
rect 597 -781 598 -780
rect 625 -781 626 -780
rect 702 -781 703 -780
rect 709 -781 710 -780
rect 1276 -781 1277 -780
rect 1283 -781 1284 -780
rect 1472 -781 1473 -780
rect 198 -783 199 -782
rect 562 -783 563 -782
rect 579 -783 580 -782
rect 996 -783 997 -782
rect 1038 -783 1039 -782
rect 1094 -783 1095 -782
rect 1136 -783 1137 -782
rect 1227 -783 1228 -782
rect 1269 -783 1270 -782
rect 1465 -783 1466 -782
rect 205 -785 206 -784
rect 240 -785 241 -784
rect 247 -785 248 -784
rect 1199 -785 1200 -784
rect 1206 -785 1207 -784
rect 1346 -785 1347 -784
rect 1381 -785 1382 -784
rect 1423 -785 1424 -784
rect 233 -787 234 -786
rect 996 -787 997 -786
rect 1080 -787 1081 -786
rect 1122 -787 1123 -786
rect 1157 -787 1158 -786
rect 1353 -787 1354 -786
rect 23 -789 24 -788
rect 233 -789 234 -788
rect 250 -789 251 -788
rect 1486 -789 1487 -788
rect 79 -791 80 -790
rect 250 -791 251 -790
rect 275 -791 276 -790
rect 380 -791 381 -790
rect 429 -791 430 -790
rect 492 -791 493 -790
rect 534 -791 535 -790
rect 1080 -791 1081 -790
rect 1171 -791 1172 -790
rect 1402 -791 1403 -790
rect 135 -793 136 -792
rect 534 -793 535 -792
rect 583 -793 584 -792
rect 597 -793 598 -792
rect 642 -793 643 -792
rect 1206 -793 1207 -792
rect 1248 -793 1249 -792
rect 1269 -793 1270 -792
rect 1290 -793 1291 -792
rect 1479 -793 1480 -792
rect 65 -795 66 -794
rect 583 -795 584 -794
rect 590 -795 591 -794
rect 1563 -795 1564 -794
rect 65 -797 66 -796
rect 828 -797 829 -796
rect 842 -797 843 -796
rect 863 -797 864 -796
rect 877 -797 878 -796
rect 1199 -797 1200 -796
rect 1262 -797 1263 -796
rect 1381 -797 1382 -796
rect 170 -799 171 -798
rect 380 -799 381 -798
rect 408 -799 409 -798
rect 492 -799 493 -798
rect 569 -799 570 -798
rect 590 -799 591 -798
rect 593 -799 594 -798
rect 1136 -799 1137 -798
rect 1185 -799 1186 -798
rect 1262 -799 1263 -798
rect 1304 -799 1305 -798
rect 1500 -799 1501 -798
rect 275 -801 276 -800
rect 796 -801 797 -800
rect 814 -801 815 -800
rect 1220 -801 1221 -800
rect 1318 -801 1319 -800
rect 1430 -801 1431 -800
rect 289 -803 290 -802
rect 352 -803 353 -802
rect 359 -803 360 -802
rect 873 -803 874 -802
rect 908 -803 909 -802
rect 1283 -803 1284 -802
rect 1325 -803 1326 -802
rect 1451 -803 1452 -802
rect 163 -805 164 -804
rect 289 -805 290 -804
rect 310 -805 311 -804
rect 758 -805 759 -804
rect 765 -805 766 -804
rect 835 -805 836 -804
rect 842 -805 843 -804
rect 849 -805 850 -804
rect 856 -805 857 -804
rect 1276 -805 1277 -804
rect 1332 -805 1333 -804
rect 1528 -805 1529 -804
rect 261 -807 262 -806
rect 1325 -807 1326 -806
rect 1339 -807 1340 -806
rect 1535 -807 1536 -806
rect 261 -809 262 -808
rect 282 -809 283 -808
rect 310 -809 311 -808
rect 387 -809 388 -808
rect 408 -809 409 -808
rect 457 -809 458 -808
rect 541 -809 542 -808
rect 569 -809 570 -808
rect 586 -809 587 -808
rect 1318 -809 1319 -808
rect 268 -811 269 -810
rect 359 -811 360 -810
rect 387 -811 388 -810
rect 422 -811 423 -810
rect 432 -811 433 -810
rect 856 -811 857 -810
rect 859 -811 860 -810
rect 1409 -811 1410 -810
rect 177 -813 178 -812
rect 422 -813 423 -812
rect 457 -813 458 -812
rect 639 -813 640 -812
rect 646 -813 647 -812
rect 702 -813 703 -812
rect 716 -813 717 -812
rect 793 -813 794 -812
rect 912 -813 913 -812
rect 1395 -813 1396 -812
rect 177 -815 178 -814
rect 212 -815 213 -814
rect 254 -815 255 -814
rect 268 -815 269 -814
rect 282 -815 283 -814
rect 436 -815 437 -814
rect 513 -815 514 -814
rect 541 -815 542 -814
rect 565 -815 566 -814
rect 1185 -815 1186 -814
rect 1192 -815 1193 -814
rect 1290 -815 1291 -814
rect 1297 -815 1298 -814
rect 1409 -815 1410 -814
rect 110 -817 111 -816
rect 1297 -817 1298 -816
rect 156 -819 157 -818
rect 254 -819 255 -818
rect 317 -819 318 -818
rect 439 -819 440 -818
rect 653 -819 654 -818
rect 1241 -819 1242 -818
rect 1255 -819 1256 -818
rect 1395 -819 1396 -818
rect 156 -821 157 -820
rect 292 -821 293 -820
rect 345 -821 346 -820
rect 618 -821 619 -820
rect 656 -821 657 -820
rect 1178 -821 1179 -820
rect 1234 -821 1235 -820
rect 1339 -821 1340 -820
rect 135 -823 136 -822
rect 1234 -823 1235 -822
rect 212 -825 213 -824
rect 219 -825 220 -824
rect 226 -825 227 -824
rect 436 -825 437 -824
rect 660 -825 661 -824
rect 789 -825 790 -824
rect 887 -825 888 -824
rect 1178 -825 1179 -824
rect 121 -827 122 -826
rect 219 -827 220 -826
rect 345 -827 346 -826
rect 548 -827 549 -826
rect 667 -827 668 -826
rect 800 -827 801 -826
rect 912 -827 913 -826
rect 1164 -827 1165 -826
rect 114 -829 115 -828
rect 121 -829 122 -828
rect 131 -829 132 -828
rect 548 -829 549 -828
rect 667 -829 668 -828
rect 691 -829 692 -828
rect 695 -829 696 -828
rect 712 -829 713 -828
rect 740 -829 741 -828
rect 1360 -829 1361 -828
rect 51 -831 52 -830
rect 695 -831 696 -830
rect 751 -831 752 -830
rect 814 -831 815 -830
rect 919 -831 920 -830
rect 1150 -831 1151 -830
rect 100 -833 101 -832
rect 114 -833 115 -832
rect 170 -833 171 -832
rect 660 -833 661 -832
rect 681 -833 682 -832
rect 723 -833 724 -832
rect 772 -833 773 -832
rect 835 -833 836 -832
rect 929 -833 930 -832
rect 1311 -833 1312 -832
rect 51 -835 52 -834
rect 1311 -835 1312 -834
rect 100 -837 101 -836
rect 1248 -837 1249 -836
rect 352 -839 353 -838
rect 464 -839 465 -838
rect 681 -839 682 -838
rect 737 -839 738 -838
rect 744 -839 745 -838
rect 772 -839 773 -838
rect 786 -839 787 -838
rect 849 -839 850 -838
rect 954 -839 955 -838
rect 1003 -839 1004 -838
rect 1006 -839 1007 -838
rect 1304 -839 1305 -838
rect 72 -841 73 -840
rect 744 -841 745 -840
rect 786 -841 787 -840
rect 1213 -841 1214 -840
rect 72 -843 73 -842
rect 331 -843 332 -842
rect 415 -843 416 -842
rect 513 -843 514 -842
rect 688 -843 689 -842
rect 751 -843 752 -842
rect 933 -843 934 -842
rect 954 -843 955 -842
rect 982 -843 983 -842
rect 1038 -843 1039 -842
rect 1052 -843 1053 -842
rect 1150 -843 1151 -842
rect 296 -845 297 -844
rect 331 -845 332 -844
rect 401 -845 402 -844
rect 415 -845 416 -844
rect 688 -845 689 -844
rect 709 -845 710 -844
rect 831 -845 832 -844
rect 1052 -845 1053 -844
rect 1066 -845 1067 -844
rect 1157 -845 1158 -844
rect 324 -847 325 -846
rect 464 -847 465 -846
rect 831 -847 832 -846
rect 1255 -847 1256 -846
rect 324 -849 325 -848
rect 520 -849 521 -848
rect 891 -849 892 -848
rect 933 -849 934 -848
rect 1017 -849 1018 -848
rect 1066 -849 1067 -848
rect 1101 -849 1102 -848
rect 1192 -849 1193 -848
rect 401 -851 402 -850
rect 443 -851 444 -850
rect 506 -851 507 -850
rect 520 -851 521 -850
rect 611 -851 612 -850
rect 891 -851 892 -850
rect 926 -851 927 -850
rect 982 -851 983 -850
rect 989 -851 990 -850
rect 1101 -851 1102 -850
rect 1108 -851 1109 -850
rect 1332 -851 1333 -850
rect 86 -853 87 -852
rect 443 -853 444 -852
rect 611 -853 612 -852
rect 1143 -853 1144 -852
rect 107 -855 108 -854
rect 1143 -855 1144 -854
rect 107 -857 108 -856
rect 870 -857 871 -856
rect 989 -857 990 -856
rect 992 -857 993 -856
rect 1017 -857 1018 -856
rect 1059 -857 1060 -856
rect 1115 -857 1116 -856
rect 1164 -857 1165 -856
rect 373 -859 374 -858
rect 506 -859 507 -858
rect 1045 -859 1046 -858
rect 1108 -859 1109 -858
rect 1129 -859 1130 -858
rect 1171 -859 1172 -858
rect 373 -861 374 -860
rect 394 -861 395 -860
rect 1010 -861 1011 -860
rect 1045 -861 1046 -860
rect 1073 -861 1074 -860
rect 1115 -861 1116 -860
rect 229 -863 230 -862
rect 394 -863 395 -862
rect 968 -863 969 -862
rect 1010 -863 1011 -862
rect 1024 -863 1025 -862
rect 1073 -863 1074 -862
rect 1087 -863 1088 -862
rect 1129 -863 1130 -862
rect 478 -865 479 -864
rect 1024 -865 1025 -864
rect 1031 -865 1032 -864
rect 1087 -865 1088 -864
rect 940 -867 941 -866
rect 968 -867 969 -866
rect 975 -867 976 -866
rect 1031 -867 1032 -866
rect 674 -869 675 -868
rect 940 -869 941 -868
rect 674 -871 675 -870
rect 737 -871 738 -870
rect 898 -871 899 -870
rect 975 -871 976 -870
rect 898 -873 899 -872
rect 905 -873 906 -872
rect 30 -884 31 -883
rect 72 -884 73 -883
rect 89 -884 90 -883
rect 114 -884 115 -883
rect 135 -884 136 -883
rect 282 -884 283 -883
rect 292 -884 293 -883
rect 338 -884 339 -883
rect 450 -884 451 -883
rect 600 -884 601 -883
rect 618 -884 619 -883
rect 737 -884 738 -883
rect 740 -884 741 -883
rect 1500 -884 1501 -883
rect 1521 -884 1522 -883
rect 1675 -884 1676 -883
rect 1696 -884 1697 -883
rect 1724 -884 1725 -883
rect 65 -886 66 -885
rect 653 -886 654 -885
rect 663 -886 664 -885
rect 1577 -886 1578 -885
rect 1591 -886 1592 -885
rect 1608 -886 1609 -885
rect 1619 -886 1620 -885
rect 1717 -886 1718 -885
rect 65 -888 66 -887
rect 401 -888 402 -887
rect 422 -888 423 -887
rect 450 -888 451 -887
rect 457 -888 458 -887
rect 929 -888 930 -887
rect 957 -888 958 -887
rect 1535 -888 1536 -887
rect 1598 -888 1599 -887
rect 1626 -888 1627 -887
rect 1633 -888 1634 -887
rect 1710 -888 1711 -887
rect 72 -890 73 -889
rect 590 -890 591 -889
rect 597 -890 598 -889
rect 611 -890 612 -889
rect 635 -890 636 -889
rect 1549 -890 1550 -889
rect 86 -892 87 -891
rect 1591 -892 1592 -891
rect 103 -894 104 -893
rect 142 -894 143 -893
rect 149 -894 150 -893
rect 737 -894 738 -893
rect 761 -894 762 -893
rect 891 -894 892 -893
rect 905 -894 906 -893
rect 1528 -894 1529 -893
rect 107 -896 108 -895
rect 121 -896 122 -895
rect 135 -896 136 -895
rect 387 -896 388 -895
rect 422 -896 423 -895
rect 758 -896 759 -895
rect 761 -896 762 -895
rect 891 -896 892 -895
rect 898 -896 899 -895
rect 905 -896 906 -895
rect 908 -896 909 -895
rect 1332 -896 1333 -895
rect 1374 -896 1375 -895
rect 1521 -896 1522 -895
rect 110 -898 111 -897
rect 338 -898 339 -897
rect 387 -898 388 -897
rect 814 -898 815 -897
rect 873 -898 874 -897
rect 1654 -898 1655 -897
rect 114 -900 115 -899
rect 415 -900 416 -899
rect 457 -900 458 -899
rect 667 -900 668 -899
rect 691 -900 692 -899
rect 1157 -900 1158 -899
rect 1206 -900 1207 -899
rect 1500 -900 1501 -899
rect 1514 -900 1515 -899
rect 1696 -900 1697 -899
rect 142 -902 143 -901
rect 478 -902 479 -901
rect 499 -902 500 -901
rect 688 -902 689 -901
rect 705 -902 706 -901
rect 1192 -902 1193 -901
rect 1220 -902 1221 -901
rect 1549 -902 1550 -901
rect 149 -904 150 -903
rect 177 -904 178 -903
rect 184 -904 185 -903
rect 208 -904 209 -903
rect 226 -904 227 -903
rect 268 -904 269 -903
rect 296 -904 297 -903
rect 845 -904 846 -903
rect 877 -904 878 -903
rect 1150 -904 1151 -903
rect 1234 -904 1235 -903
rect 1626 -904 1627 -903
rect 128 -906 129 -905
rect 177 -906 178 -905
rect 184 -906 185 -905
rect 250 -906 251 -905
rect 261 -906 262 -905
rect 282 -906 283 -905
rect 303 -906 304 -905
rect 607 -906 608 -905
rect 611 -906 612 -905
rect 961 -906 962 -905
rect 964 -906 965 -905
rect 1647 -906 1648 -905
rect 128 -908 129 -907
rect 793 -908 794 -907
rect 796 -908 797 -907
rect 1346 -908 1347 -907
rect 1395 -908 1396 -907
rect 1528 -908 1529 -907
rect 138 -910 139 -909
rect 268 -910 269 -909
rect 303 -910 304 -909
rect 583 -910 584 -909
rect 586 -910 587 -909
rect 1542 -910 1543 -909
rect 163 -912 164 -911
rect 996 -912 997 -911
rect 1038 -912 1039 -911
rect 1157 -912 1158 -911
rect 1248 -912 1249 -911
rect 1374 -912 1375 -911
rect 1430 -912 1431 -911
rect 1535 -912 1536 -911
rect 163 -914 164 -913
rect 324 -914 325 -913
rect 331 -914 332 -913
rect 401 -914 402 -913
rect 415 -914 416 -913
rect 716 -914 717 -913
rect 768 -914 769 -913
rect 1633 -914 1634 -913
rect 93 -916 94 -915
rect 324 -916 325 -915
rect 373 -916 374 -915
rect 499 -916 500 -915
rect 548 -916 549 -915
rect 667 -916 668 -915
rect 786 -916 787 -915
rect 1584 -916 1585 -915
rect 86 -918 87 -917
rect 93 -918 94 -917
rect 166 -918 167 -917
rect 513 -918 514 -917
rect 548 -918 549 -917
rect 1682 -918 1683 -917
rect 170 -920 171 -919
rect 481 -920 482 -919
rect 513 -920 514 -919
rect 901 -920 902 -919
rect 912 -920 913 -919
rect 926 -920 927 -919
rect 933 -920 934 -919
rect 996 -920 997 -919
rect 1059 -920 1060 -919
rect 1465 -920 1466 -919
rect 1486 -920 1487 -919
rect 1605 -920 1606 -919
rect 170 -922 171 -921
rect 240 -922 241 -921
rect 247 -922 248 -921
rect 289 -922 290 -921
rect 310 -922 311 -921
rect 593 -922 594 -921
rect 646 -922 647 -921
rect 649 -922 650 -921
rect 733 -922 734 -921
rect 1486 -922 1487 -921
rect 1493 -922 1494 -921
rect 1668 -922 1669 -921
rect 191 -924 192 -923
rect 660 -924 661 -923
rect 765 -924 766 -923
rect 786 -924 787 -923
rect 810 -924 811 -923
rect 1703 -924 1704 -923
rect 79 -926 80 -925
rect 191 -926 192 -925
rect 198 -926 199 -925
rect 660 -926 661 -925
rect 765 -926 766 -925
rect 1325 -926 1326 -925
rect 1339 -926 1340 -925
rect 1465 -926 1466 -925
rect 79 -928 80 -927
rect 562 -928 563 -927
rect 576 -928 577 -927
rect 702 -928 703 -927
rect 856 -928 857 -927
rect 912 -928 913 -927
rect 919 -928 920 -927
rect 961 -928 962 -927
rect 968 -928 969 -927
rect 971 -928 972 -927
rect 975 -928 976 -927
rect 1038 -928 1039 -927
rect 1062 -928 1063 -927
rect 1388 -928 1389 -927
rect 1437 -928 1438 -927
rect 1584 -928 1585 -927
rect 124 -930 125 -929
rect 198 -930 199 -929
rect 205 -930 206 -929
rect 621 -930 622 -929
rect 646 -930 647 -929
rect 1094 -930 1095 -929
rect 1101 -930 1102 -929
rect 1234 -930 1235 -929
rect 1262 -930 1263 -929
rect 1395 -930 1396 -929
rect 1444 -930 1445 -929
rect 1661 -930 1662 -929
rect 226 -932 227 -931
rect 579 -932 580 -931
rect 583 -932 584 -931
rect 695 -932 696 -931
rect 772 -932 773 -931
rect 1388 -932 1389 -931
rect 1458 -932 1459 -931
rect 1619 -932 1620 -931
rect 229 -934 230 -933
rect 1143 -934 1144 -933
rect 1150 -934 1151 -933
rect 1381 -934 1382 -933
rect 1458 -934 1459 -933
rect 1507 -934 1508 -933
rect 121 -936 122 -935
rect 1507 -936 1508 -935
rect 233 -938 234 -937
rect 1570 -938 1571 -937
rect 89 -940 90 -939
rect 233 -940 234 -939
rect 236 -940 237 -939
rect 1640 -940 1641 -939
rect 240 -942 241 -941
rect 352 -942 353 -941
rect 373 -942 374 -941
rect 408 -942 409 -941
rect 436 -942 437 -941
rect 1220 -942 1221 -941
rect 1255 -942 1256 -941
rect 1570 -942 1571 -941
rect 261 -944 262 -943
rect 429 -944 430 -943
rect 436 -944 437 -943
rect 723 -944 724 -943
rect 730 -944 731 -943
rect 772 -944 773 -943
rect 856 -944 857 -943
rect 1514 -944 1515 -943
rect 289 -946 290 -945
rect 1248 -946 1249 -945
rect 1255 -946 1256 -945
rect 1269 -946 1270 -945
rect 1297 -946 1298 -945
rect 1689 -946 1690 -945
rect 37 -948 38 -947
rect 1297 -948 1298 -947
rect 1304 -948 1305 -947
rect 1444 -948 1445 -947
rect 313 -950 314 -949
rect 331 -950 332 -949
rect 345 -950 346 -949
rect 562 -950 563 -949
rect 576 -950 577 -949
rect 632 -950 633 -949
rect 709 -950 710 -949
rect 730 -950 731 -949
rect 863 -950 864 -949
rect 926 -950 927 -949
rect 940 -950 941 -949
rect 1143 -950 1144 -949
rect 1178 -950 1179 -949
rect 1304 -950 1305 -949
rect 1346 -950 1347 -949
rect 1367 -950 1368 -949
rect 1381 -950 1382 -949
rect 1612 -950 1613 -949
rect 317 -952 318 -951
rect 467 -952 468 -951
rect 474 -952 475 -951
rect 674 -952 675 -951
rect 800 -952 801 -951
rect 940 -952 941 -951
rect 968 -952 969 -951
rect 1017 -952 1018 -951
rect 1031 -952 1032 -951
rect 1339 -952 1340 -951
rect 1353 -952 1354 -951
rect 1493 -952 1494 -951
rect 345 -954 346 -953
rect 366 -954 367 -953
rect 394 -954 395 -953
rect 408 -954 409 -953
rect 429 -954 430 -953
rect 625 -954 626 -953
rect 632 -954 633 -953
rect 814 -954 815 -953
rect 849 -954 850 -953
rect 863 -954 864 -953
rect 870 -954 871 -953
rect 1437 -954 1438 -953
rect 107 -956 108 -955
rect 849 -956 850 -955
rect 870 -956 871 -955
rect 1178 -956 1179 -955
rect 1199 -956 1200 -955
rect 1325 -956 1326 -955
rect 1353 -956 1354 -955
rect 1409 -956 1410 -955
rect 352 -958 353 -957
rect 380 -958 381 -957
rect 394 -958 395 -957
rect 723 -958 724 -957
rect 800 -958 801 -957
rect 821 -958 822 -957
rect 877 -958 878 -957
rect 1416 -958 1417 -957
rect 366 -960 367 -959
rect 471 -960 472 -959
rect 478 -960 479 -959
rect 555 -960 556 -959
rect 604 -960 605 -959
rect 709 -960 710 -959
rect 751 -960 752 -959
rect 821 -960 822 -959
rect 884 -960 885 -959
rect 887 -960 888 -959
rect 898 -960 899 -959
rect 1241 -960 1242 -959
rect 1283 -960 1284 -959
rect 1409 -960 1410 -959
rect 37 -962 38 -961
rect 471 -962 472 -961
rect 520 -962 521 -961
rect 555 -962 556 -961
rect 604 -962 605 -961
rect 1577 -962 1578 -961
rect 380 -964 381 -963
rect 485 -964 486 -963
rect 492 -964 493 -963
rect 520 -964 521 -963
rect 527 -964 528 -963
rect 751 -964 752 -963
rect 884 -964 885 -963
rect 982 -964 983 -963
rect 1003 -964 1004 -963
rect 1094 -964 1095 -963
rect 1115 -964 1116 -963
rect 1262 -964 1263 -963
rect 1290 -964 1291 -963
rect 1416 -964 1417 -963
rect 44 -966 45 -965
rect 485 -966 486 -965
rect 534 -966 535 -965
rect 919 -966 920 -965
rect 947 -966 948 -965
rect 1031 -966 1032 -965
rect 1052 -966 1053 -965
rect 1199 -966 1200 -965
rect 1213 -966 1214 -965
rect 1612 -966 1613 -965
rect 44 -968 45 -967
rect 54 -968 55 -967
rect 58 -968 59 -967
rect 492 -968 493 -967
rect 537 -968 538 -967
rect 933 -968 934 -967
rect 975 -968 976 -967
rect 1430 -968 1431 -967
rect 54 -970 55 -969
rect 1556 -970 1557 -969
rect 58 -972 59 -971
rect 1136 -972 1137 -971
rect 1164 -972 1165 -971
rect 1290 -972 1291 -971
rect 100 -974 101 -973
rect 1556 -974 1557 -973
rect 23 -976 24 -975
rect 100 -976 101 -975
rect 219 -976 220 -975
rect 947 -976 948 -975
rect 978 -976 979 -975
rect 1601 -976 1602 -975
rect 359 -978 360 -977
rect 527 -978 528 -977
rect 551 -978 552 -977
rect 744 -978 745 -977
rect 880 -978 881 -977
rect 1115 -978 1116 -977
rect 1129 -978 1130 -977
rect 1269 -978 1270 -977
rect 212 -980 213 -979
rect 359 -980 360 -979
rect 443 -980 444 -979
rect 716 -980 717 -979
rect 744 -980 745 -979
rect 992 -980 993 -979
rect 1003 -980 1004 -979
rect 1108 -980 1109 -979
rect 1122 -980 1123 -979
rect 1129 -980 1130 -979
rect 1164 -980 1165 -979
rect 1171 -980 1172 -979
rect 156 -982 157 -981
rect 443 -982 444 -981
rect 467 -982 468 -981
rect 1241 -982 1242 -981
rect 156 -984 157 -983
rect 793 -984 794 -983
rect 835 -984 836 -983
rect 1122 -984 1123 -983
rect 212 -986 213 -985
rect 541 -986 542 -985
rect 614 -986 615 -985
rect 674 -986 675 -985
rect 835 -986 836 -985
rect 842 -986 843 -985
rect 971 -986 972 -985
rect 1017 -986 1018 -985
rect 1024 -986 1025 -985
rect 1136 -986 1137 -985
rect 541 -988 542 -987
rect 597 -988 598 -987
rect 618 -988 619 -987
rect 695 -988 696 -987
rect 796 -988 797 -987
rect 1024 -988 1025 -987
rect 1045 -988 1046 -987
rect 1171 -988 1172 -987
rect 625 -990 626 -989
rect 681 -990 682 -989
rect 842 -990 843 -989
rect 1332 -990 1333 -989
rect 639 -992 640 -991
rect 1367 -992 1368 -991
rect 639 -994 640 -993
rect 880 -994 881 -993
rect 954 -994 955 -993
rect 1045 -994 1046 -993
rect 1062 -994 1063 -993
rect 1472 -994 1473 -993
rect 681 -996 682 -995
rect 1283 -996 1284 -995
rect 789 -998 790 -997
rect 1472 -998 1473 -997
rect 954 -1000 955 -999
rect 1563 -1000 1564 -999
rect 989 -1002 990 -1001
rect 1052 -1002 1053 -1001
rect 1066 -1002 1067 -1001
rect 1192 -1002 1193 -1001
rect 1451 -1002 1452 -1001
rect 1563 -1002 1564 -1001
rect 989 -1004 990 -1003
rect 1542 -1004 1543 -1003
rect 1010 -1006 1011 -1005
rect 1101 -1006 1102 -1005
rect 1311 -1006 1312 -1005
rect 1451 -1006 1452 -1005
rect 534 -1008 535 -1007
rect 1311 -1008 1312 -1007
rect 1066 -1010 1067 -1009
rect 1402 -1010 1403 -1009
rect 1073 -1012 1074 -1011
rect 1206 -1012 1207 -1011
rect 1402 -1012 1403 -1011
rect 1423 -1012 1424 -1011
rect 628 -1014 629 -1013
rect 1073 -1014 1074 -1013
rect 1080 -1014 1081 -1013
rect 1213 -1014 1214 -1013
rect 779 -1016 780 -1015
rect 1080 -1016 1081 -1015
rect 779 -1018 780 -1017
rect 807 -1018 808 -1017
rect 828 -1018 829 -1017
rect 1423 -1018 1424 -1017
rect 807 -1020 808 -1019
rect 1010 -1020 1011 -1019
rect 828 -1022 829 -1021
rect 1360 -1022 1361 -1021
rect 1360 -1024 1361 -1023
rect 1479 -1024 1480 -1023
rect 1318 -1026 1319 -1025
rect 1479 -1026 1480 -1025
rect 1185 -1028 1186 -1027
rect 1318 -1028 1319 -1027
rect 1185 -1030 1186 -1029
rect 1227 -1030 1228 -1029
rect 1087 -1032 1088 -1031
rect 1227 -1032 1228 -1031
rect 201 -1034 202 -1033
rect 1087 -1034 1088 -1033
rect 44 -1045 45 -1044
rect 240 -1045 241 -1044
rect 261 -1045 262 -1044
rect 632 -1045 633 -1044
rect 681 -1045 682 -1044
rect 1143 -1045 1144 -1044
rect 1710 -1045 1711 -1044
rect 1731 -1045 1732 -1044
rect 65 -1047 66 -1046
rect 488 -1047 489 -1046
rect 499 -1047 500 -1046
rect 632 -1047 633 -1046
rect 681 -1047 682 -1046
rect 695 -1047 696 -1046
rect 719 -1047 720 -1046
rect 1521 -1047 1522 -1046
rect 65 -1049 66 -1048
rect 544 -1049 545 -1048
rect 579 -1049 580 -1048
rect 1367 -1049 1368 -1048
rect 86 -1051 87 -1050
rect 940 -1051 941 -1050
rect 957 -1051 958 -1050
rect 1626 -1051 1627 -1050
rect 89 -1053 90 -1052
rect 1514 -1053 1515 -1052
rect 1626 -1053 1627 -1052
rect 1668 -1053 1669 -1052
rect 93 -1055 94 -1054
rect 187 -1055 188 -1054
rect 198 -1055 199 -1054
rect 401 -1055 402 -1054
rect 408 -1055 409 -1054
rect 534 -1055 535 -1054
rect 590 -1055 591 -1054
rect 1500 -1055 1501 -1054
rect 51 -1057 52 -1056
rect 590 -1057 591 -1056
rect 597 -1057 598 -1056
rect 716 -1057 717 -1056
rect 723 -1057 724 -1056
rect 1549 -1057 1550 -1056
rect 51 -1059 52 -1058
rect 555 -1059 556 -1058
rect 600 -1059 601 -1058
rect 1010 -1059 1011 -1058
rect 1062 -1059 1063 -1058
rect 1521 -1059 1522 -1058
rect 93 -1061 94 -1060
rect 443 -1061 444 -1060
rect 450 -1061 451 -1060
rect 499 -1061 500 -1060
rect 513 -1061 514 -1060
rect 555 -1061 556 -1060
rect 569 -1061 570 -1060
rect 600 -1061 601 -1060
rect 614 -1061 615 -1060
rect 919 -1061 920 -1060
rect 940 -1061 941 -1060
rect 1038 -1061 1039 -1060
rect 1069 -1061 1070 -1060
rect 1696 -1061 1697 -1060
rect 54 -1063 55 -1062
rect 443 -1063 444 -1062
rect 450 -1063 451 -1062
rect 520 -1063 521 -1062
rect 527 -1063 528 -1062
rect 716 -1063 717 -1062
rect 726 -1063 727 -1062
rect 730 -1063 731 -1062
rect 751 -1063 752 -1062
rect 807 -1063 808 -1062
rect 810 -1063 811 -1062
rect 1045 -1063 1046 -1062
rect 1143 -1063 1144 -1062
rect 1234 -1063 1235 -1062
rect 1360 -1063 1361 -1062
rect 1549 -1063 1550 -1062
rect 100 -1065 101 -1064
rect 289 -1065 290 -1064
rect 292 -1065 293 -1064
rect 604 -1065 605 -1064
rect 702 -1065 703 -1064
rect 730 -1065 731 -1064
rect 751 -1065 752 -1064
rect 1381 -1065 1382 -1064
rect 1500 -1065 1501 -1064
rect 1612 -1065 1613 -1064
rect 103 -1067 104 -1066
rect 1388 -1067 1389 -1066
rect 1612 -1067 1613 -1066
rect 1654 -1067 1655 -1066
rect 107 -1069 108 -1068
rect 415 -1069 416 -1068
rect 464 -1069 465 -1068
rect 947 -1069 948 -1068
rect 971 -1069 972 -1068
rect 1048 -1069 1049 -1068
rect 1234 -1069 1235 -1068
rect 1650 -1069 1651 -1068
rect 107 -1071 108 -1070
rect 747 -1071 748 -1070
rect 758 -1071 759 -1070
rect 1227 -1071 1228 -1070
rect 1276 -1071 1277 -1070
rect 1360 -1071 1361 -1070
rect 1367 -1071 1368 -1070
rect 1465 -1071 1466 -1070
rect 89 -1073 90 -1072
rect 1465 -1073 1466 -1072
rect 110 -1075 111 -1074
rect 1479 -1075 1480 -1074
rect 121 -1077 122 -1076
rect 1220 -1077 1221 -1076
rect 1227 -1077 1228 -1076
rect 1290 -1077 1291 -1076
rect 1381 -1077 1382 -1076
rect 1535 -1077 1536 -1076
rect 121 -1079 122 -1078
rect 436 -1079 437 -1078
rect 478 -1079 479 -1078
rect 534 -1079 535 -1078
rect 621 -1079 622 -1078
rect 1276 -1079 1277 -1078
rect 1290 -1079 1291 -1078
rect 1409 -1079 1410 -1078
rect 1479 -1079 1480 -1078
rect 1640 -1079 1641 -1078
rect 128 -1081 129 -1080
rect 436 -1081 437 -1080
rect 506 -1081 507 -1080
rect 527 -1081 528 -1080
rect 621 -1081 622 -1080
rect 1122 -1081 1123 -1080
rect 1388 -1081 1389 -1080
rect 1430 -1081 1431 -1080
rect 1640 -1081 1641 -1080
rect 1675 -1081 1676 -1080
rect 128 -1083 129 -1082
rect 744 -1083 745 -1082
rect 768 -1083 769 -1082
rect 1339 -1083 1340 -1082
rect 1402 -1083 1403 -1082
rect 1654 -1083 1655 -1082
rect 135 -1085 136 -1084
rect 467 -1085 468 -1084
rect 506 -1085 507 -1084
rect 1241 -1085 1242 -1084
rect 1255 -1085 1256 -1084
rect 1430 -1085 1431 -1084
rect 1619 -1085 1620 -1084
rect 1675 -1085 1676 -1084
rect 135 -1087 136 -1086
rect 205 -1087 206 -1086
rect 208 -1087 209 -1086
rect 1311 -1087 1312 -1086
rect 1339 -1087 1340 -1086
rect 1374 -1087 1375 -1086
rect 1409 -1087 1410 -1086
rect 1451 -1087 1452 -1086
rect 142 -1089 143 -1088
rect 569 -1089 570 -1088
rect 628 -1089 629 -1088
rect 1451 -1089 1452 -1088
rect 142 -1091 143 -1090
rect 149 -1091 150 -1090
rect 166 -1091 167 -1090
rect 198 -1091 199 -1090
rect 219 -1091 220 -1090
rect 247 -1091 248 -1090
rect 261 -1091 262 -1090
rect 828 -1091 829 -1090
rect 845 -1091 846 -1090
rect 1150 -1091 1151 -1090
rect 1241 -1091 1242 -1090
rect 1297 -1091 1298 -1090
rect 1311 -1091 1312 -1090
rect 1437 -1091 1438 -1090
rect 149 -1093 150 -1092
rect 303 -1093 304 -1092
rect 310 -1093 311 -1092
rect 331 -1093 332 -1092
rect 359 -1093 360 -1092
rect 415 -1093 416 -1092
rect 513 -1093 514 -1092
rect 576 -1093 577 -1092
rect 702 -1093 703 -1092
rect 1423 -1093 1424 -1092
rect 1437 -1093 1438 -1092
rect 1458 -1093 1459 -1092
rect 170 -1095 171 -1094
rect 408 -1095 409 -1094
rect 516 -1095 517 -1094
rect 758 -1095 759 -1094
rect 786 -1095 787 -1094
rect 842 -1095 843 -1094
rect 859 -1095 860 -1094
rect 1514 -1095 1515 -1094
rect 170 -1097 171 -1096
rect 191 -1097 192 -1096
rect 212 -1097 213 -1096
rect 303 -1097 304 -1096
rect 331 -1097 332 -1096
rect 345 -1097 346 -1096
rect 359 -1097 360 -1096
rect 485 -1097 486 -1096
rect 520 -1097 521 -1096
rect 541 -1097 542 -1096
rect 733 -1097 734 -1096
rect 1220 -1097 1221 -1096
rect 1297 -1097 1298 -1096
rect 1416 -1097 1417 -1096
rect 1458 -1097 1459 -1096
rect 1472 -1097 1473 -1096
rect 47 -1099 48 -1098
rect 541 -1099 542 -1098
rect 744 -1099 745 -1098
rect 996 -1099 997 -1098
rect 1010 -1099 1011 -1098
rect 1094 -1099 1095 -1098
rect 1122 -1099 1123 -1098
rect 1178 -1099 1179 -1098
rect 1346 -1099 1347 -1098
rect 1423 -1099 1424 -1098
rect 1472 -1099 1473 -1098
rect 1528 -1099 1529 -1098
rect 79 -1101 80 -1100
rect 191 -1101 192 -1100
rect 212 -1101 213 -1100
rect 254 -1101 255 -1100
rect 282 -1101 283 -1100
rect 345 -1101 346 -1100
rect 366 -1101 367 -1100
rect 474 -1101 475 -1100
rect 485 -1101 486 -1100
rect 1535 -1101 1536 -1100
rect 79 -1103 80 -1102
rect 1556 -1103 1557 -1102
rect 163 -1105 164 -1104
rect 254 -1105 255 -1104
rect 275 -1105 276 -1104
rect 282 -1105 283 -1104
rect 289 -1105 290 -1104
rect 317 -1105 318 -1104
rect 366 -1105 367 -1104
rect 551 -1105 552 -1104
rect 793 -1105 794 -1104
rect 1584 -1105 1585 -1104
rect 114 -1107 115 -1106
rect 317 -1107 318 -1106
rect 380 -1107 381 -1106
rect 695 -1107 696 -1106
rect 807 -1107 808 -1106
rect 1073 -1107 1074 -1106
rect 1115 -1107 1116 -1106
rect 1584 -1107 1585 -1106
rect 114 -1109 115 -1108
rect 779 -1109 780 -1108
rect 842 -1109 843 -1108
rect 1045 -1109 1046 -1108
rect 1073 -1109 1074 -1108
rect 1087 -1109 1088 -1108
rect 1115 -1109 1116 -1108
rect 1171 -1109 1172 -1108
rect 1178 -1109 1179 -1108
rect 1213 -1109 1214 -1108
rect 1332 -1109 1333 -1108
rect 1346 -1109 1347 -1108
rect 1374 -1109 1375 -1108
rect 1605 -1109 1606 -1108
rect 156 -1111 157 -1110
rect 275 -1111 276 -1110
rect 380 -1111 381 -1110
rect 467 -1111 468 -1110
rect 723 -1111 724 -1110
rect 1213 -1111 1214 -1110
rect 1528 -1111 1529 -1110
rect 1542 -1111 1543 -1110
rect 1556 -1111 1557 -1110
rect 1577 -1111 1578 -1110
rect 156 -1113 157 -1112
rect 646 -1113 647 -1112
rect 772 -1113 773 -1112
rect 779 -1113 780 -1112
rect 849 -1113 850 -1112
rect 1332 -1113 1333 -1112
rect 1542 -1113 1543 -1112
rect 1661 -1113 1662 -1112
rect 75 -1115 76 -1114
rect 849 -1115 850 -1114
rect 856 -1115 857 -1114
rect 1094 -1115 1095 -1114
rect 1150 -1115 1151 -1114
rect 1248 -1115 1249 -1114
rect 177 -1117 178 -1116
rect 625 -1117 626 -1116
rect 646 -1117 647 -1116
rect 667 -1117 668 -1116
rect 674 -1117 675 -1116
rect 772 -1117 773 -1116
rect 835 -1117 836 -1116
rect 856 -1117 857 -1116
rect 870 -1117 871 -1116
rect 1059 -1117 1060 -1116
rect 1164 -1117 1165 -1116
rect 1171 -1117 1172 -1116
rect 1248 -1117 1249 -1116
rect 1325 -1117 1326 -1116
rect 177 -1119 178 -1118
rect 1664 -1119 1665 -1118
rect 201 -1121 202 -1120
rect 1087 -1121 1088 -1120
rect 1164 -1121 1165 -1120
rect 1262 -1121 1263 -1120
rect 201 -1123 202 -1122
rect 457 -1123 458 -1122
rect 537 -1123 538 -1122
rect 674 -1123 675 -1122
rect 821 -1123 822 -1122
rect 870 -1123 871 -1122
rect 873 -1123 874 -1122
rect 1493 -1123 1494 -1122
rect 205 -1125 206 -1124
rect 1605 -1125 1606 -1124
rect 236 -1127 237 -1126
rect 1255 -1127 1256 -1126
rect 1353 -1127 1354 -1126
rect 1493 -1127 1494 -1126
rect 240 -1129 241 -1128
rect 639 -1129 640 -1128
rect 667 -1129 668 -1128
rect 688 -1129 689 -1128
rect 821 -1129 822 -1128
rect 1101 -1129 1102 -1128
rect 1185 -1129 1186 -1128
rect 1262 -1129 1263 -1128
rect 1353 -1129 1354 -1128
rect 1395 -1129 1396 -1128
rect 58 -1131 59 -1130
rect 688 -1131 689 -1130
rect 835 -1131 836 -1130
rect 968 -1131 969 -1130
rect 975 -1131 976 -1130
rect 1031 -1131 1032 -1130
rect 1038 -1131 1039 -1130
rect 1206 -1131 1207 -1130
rect 1395 -1131 1396 -1130
rect 1444 -1131 1445 -1130
rect 58 -1133 59 -1132
rect 663 -1133 664 -1132
rect 877 -1133 878 -1132
rect 1619 -1133 1620 -1132
rect 247 -1135 248 -1134
rect 268 -1135 269 -1134
rect 387 -1135 388 -1134
rect 604 -1135 605 -1134
rect 625 -1135 626 -1134
rect 954 -1135 955 -1134
rect 978 -1135 979 -1134
rect 1577 -1135 1578 -1134
rect 163 -1137 164 -1136
rect 268 -1137 269 -1136
rect 394 -1137 395 -1136
rect 880 -1137 881 -1136
rect 894 -1137 895 -1136
rect 1416 -1137 1417 -1136
rect 1444 -1137 1445 -1136
rect 1507 -1137 1508 -1136
rect 226 -1139 227 -1138
rect 387 -1139 388 -1138
rect 394 -1139 395 -1138
rect 754 -1139 755 -1138
rect 877 -1139 878 -1138
rect 884 -1139 885 -1138
rect 898 -1139 899 -1138
rect 1633 -1139 1634 -1138
rect 30 -1141 31 -1140
rect 226 -1141 227 -1140
rect 401 -1141 402 -1140
rect 593 -1141 594 -1140
rect 639 -1141 640 -1140
rect 737 -1141 738 -1140
rect 898 -1141 899 -1140
rect 1507 -1141 1508 -1140
rect 1598 -1141 1599 -1140
rect 1633 -1141 1634 -1140
rect 30 -1143 31 -1142
rect 583 -1143 584 -1142
rect 709 -1143 710 -1142
rect 737 -1143 738 -1142
rect 912 -1143 913 -1142
rect 968 -1143 969 -1142
rect 989 -1143 990 -1142
rect 1689 -1143 1690 -1142
rect 233 -1145 234 -1144
rect 583 -1145 584 -1144
rect 709 -1145 710 -1144
rect 1066 -1145 1067 -1144
rect 1101 -1145 1102 -1144
rect 1157 -1145 1158 -1144
rect 1563 -1145 1564 -1144
rect 1598 -1145 1599 -1144
rect 422 -1147 423 -1146
rect 786 -1147 787 -1146
rect 912 -1147 913 -1146
rect 926 -1147 927 -1146
rect 933 -1147 934 -1146
rect 1325 -1147 1326 -1146
rect 1563 -1147 1564 -1146
rect 1591 -1147 1592 -1146
rect 422 -1149 423 -1148
rect 548 -1149 549 -1148
rect 726 -1149 727 -1148
rect 926 -1149 927 -1148
rect 947 -1149 948 -1148
rect 982 -1149 983 -1148
rect 989 -1149 990 -1148
rect 1402 -1149 1403 -1148
rect 1591 -1149 1592 -1148
rect 1647 -1149 1648 -1148
rect 324 -1151 325 -1150
rect 548 -1151 549 -1150
rect 765 -1151 766 -1150
rect 933 -1151 934 -1150
rect 954 -1151 955 -1150
rect 1570 -1151 1571 -1150
rect 1647 -1151 1648 -1150
rect 1717 -1151 1718 -1150
rect 100 -1153 101 -1152
rect 324 -1153 325 -1152
rect 429 -1153 430 -1152
rect 793 -1153 794 -1152
rect 814 -1153 815 -1152
rect 982 -1153 983 -1152
rect 992 -1153 993 -1152
rect 1206 -1153 1207 -1152
rect 1570 -1153 1571 -1152
rect 1682 -1153 1683 -1152
rect 373 -1155 374 -1154
rect 429 -1155 430 -1154
rect 457 -1155 458 -1154
rect 611 -1155 612 -1154
rect 814 -1155 815 -1154
rect 863 -1155 864 -1154
rect 919 -1155 920 -1154
rect 961 -1155 962 -1154
rect 992 -1155 993 -1154
rect 1486 -1155 1487 -1154
rect 373 -1157 374 -1156
rect 660 -1157 661 -1156
rect 800 -1157 801 -1156
rect 863 -1157 864 -1156
rect 996 -1157 997 -1156
rect 1024 -1157 1025 -1156
rect 1031 -1157 1032 -1156
rect 1108 -1157 1109 -1156
rect 1157 -1157 1158 -1156
rect 1283 -1157 1284 -1156
rect 1486 -1157 1487 -1156
rect 1703 -1157 1704 -1156
rect 338 -1159 339 -1158
rect 800 -1159 801 -1158
rect 831 -1159 832 -1158
rect 961 -1159 962 -1158
rect 1003 -1159 1004 -1158
rect 1185 -1159 1186 -1158
rect 1283 -1159 1284 -1158
rect 1318 -1159 1319 -1158
rect 184 -1161 185 -1160
rect 338 -1161 339 -1160
rect 471 -1161 472 -1160
rect 884 -1161 885 -1160
rect 957 -1161 958 -1160
rect 1318 -1161 1319 -1160
rect 37 -1163 38 -1162
rect 471 -1163 472 -1162
rect 562 -1163 563 -1162
rect 765 -1163 766 -1162
rect 1003 -1163 1004 -1162
rect 1052 -1163 1053 -1162
rect 37 -1165 38 -1164
rect 72 -1165 73 -1164
rect 124 -1165 125 -1164
rect 1052 -1165 1053 -1164
rect 184 -1167 185 -1166
rect 478 -1167 479 -1166
rect 492 -1167 493 -1166
rect 562 -1167 563 -1166
rect 611 -1167 612 -1166
rect 891 -1167 892 -1166
rect 1017 -1167 1018 -1166
rect 1066 -1167 1067 -1166
rect 492 -1169 493 -1168
rect 761 -1169 762 -1168
rect 1017 -1169 1018 -1168
rect 1080 -1169 1081 -1168
rect 635 -1171 636 -1170
rect 1108 -1171 1109 -1170
rect 660 -1173 661 -1172
rect 1199 -1173 1200 -1172
rect 901 -1175 902 -1174
rect 1199 -1175 1200 -1174
rect 1024 -1177 1025 -1176
rect 1136 -1177 1137 -1176
rect 1080 -1179 1081 -1178
rect 1269 -1179 1270 -1178
rect 1136 -1181 1137 -1180
rect 1192 -1181 1193 -1180
rect 1269 -1181 1270 -1180
rect 1304 -1181 1305 -1180
rect 597 -1183 598 -1182
rect 1192 -1183 1193 -1182
rect 607 -1185 608 -1184
rect 1304 -1185 1305 -1184
rect 23 -1196 24 -1195
rect 65 -1196 66 -1195
rect 79 -1196 80 -1195
rect 100 -1196 101 -1195
rect 124 -1196 125 -1195
rect 1115 -1196 1116 -1195
rect 1486 -1196 1487 -1195
rect 1689 -1196 1690 -1195
rect 1717 -1196 1718 -1195
rect 1724 -1196 1725 -1195
rect 1731 -1196 1732 -1195
rect 1738 -1196 1739 -1195
rect 30 -1198 31 -1197
rect 89 -1198 90 -1197
rect 93 -1198 94 -1197
rect 145 -1198 146 -1197
rect 149 -1198 150 -1197
rect 205 -1198 206 -1197
rect 208 -1198 209 -1197
rect 793 -1198 794 -1197
rect 810 -1198 811 -1197
rect 835 -1198 836 -1197
rect 873 -1198 874 -1197
rect 1598 -1198 1599 -1197
rect 1605 -1198 1606 -1197
rect 1682 -1198 1683 -1197
rect 30 -1200 31 -1199
rect 488 -1200 489 -1199
rect 506 -1200 507 -1199
rect 695 -1200 696 -1199
rect 723 -1200 724 -1199
rect 1185 -1200 1186 -1199
rect 1451 -1200 1452 -1199
rect 1486 -1200 1487 -1199
rect 1500 -1200 1501 -1199
rect 1598 -1200 1599 -1199
rect 1619 -1200 1620 -1199
rect 1668 -1200 1669 -1199
rect 1675 -1200 1676 -1199
rect 1731 -1200 1732 -1199
rect 58 -1202 59 -1201
rect 121 -1202 122 -1201
rect 135 -1202 136 -1201
rect 513 -1202 514 -1201
rect 541 -1202 542 -1201
rect 709 -1202 710 -1201
rect 744 -1202 745 -1201
rect 1136 -1202 1137 -1201
rect 1185 -1202 1186 -1201
rect 1325 -1202 1326 -1201
rect 1465 -1202 1466 -1201
rect 1619 -1202 1620 -1201
rect 1654 -1202 1655 -1201
rect 1675 -1202 1676 -1201
rect 58 -1204 59 -1203
rect 247 -1204 248 -1203
rect 250 -1204 251 -1203
rect 352 -1204 353 -1203
rect 380 -1204 381 -1203
rect 723 -1204 724 -1203
rect 744 -1204 745 -1203
rect 779 -1204 780 -1203
rect 814 -1204 815 -1203
rect 898 -1204 899 -1203
rect 901 -1204 902 -1203
rect 1444 -1204 1445 -1203
rect 1591 -1204 1592 -1203
rect 1605 -1204 1606 -1203
rect 1661 -1204 1662 -1203
rect 1724 -1204 1725 -1203
rect 65 -1206 66 -1205
rect 201 -1206 202 -1205
rect 205 -1206 206 -1205
rect 576 -1206 577 -1205
rect 593 -1206 594 -1205
rect 1402 -1206 1403 -1205
rect 1416 -1206 1417 -1205
rect 1465 -1206 1466 -1205
rect 1542 -1206 1543 -1205
rect 1661 -1206 1662 -1205
rect 96 -1208 97 -1207
rect 1514 -1208 1515 -1207
rect 1528 -1208 1529 -1207
rect 1542 -1208 1543 -1207
rect 121 -1210 122 -1209
rect 1521 -1210 1522 -1209
rect 135 -1212 136 -1211
rect 359 -1212 360 -1211
rect 380 -1212 381 -1211
rect 387 -1212 388 -1211
rect 422 -1212 423 -1211
rect 516 -1212 517 -1211
rect 530 -1212 531 -1211
rect 1136 -1212 1137 -1211
rect 1206 -1212 1207 -1211
rect 1444 -1212 1445 -1211
rect 1521 -1212 1522 -1211
rect 1570 -1212 1571 -1211
rect 142 -1214 143 -1213
rect 149 -1214 150 -1213
rect 163 -1214 164 -1213
rect 1297 -1214 1298 -1213
rect 1325 -1214 1326 -1213
rect 1395 -1214 1396 -1213
rect 1416 -1214 1417 -1213
rect 1479 -1214 1480 -1213
rect 142 -1216 143 -1215
rect 1122 -1216 1123 -1215
rect 1129 -1216 1130 -1215
rect 1206 -1216 1207 -1215
rect 1241 -1216 1242 -1215
rect 1297 -1216 1298 -1215
rect 1339 -1216 1340 -1215
rect 1402 -1216 1403 -1215
rect 1409 -1216 1410 -1215
rect 1479 -1216 1480 -1215
rect 124 -1218 125 -1217
rect 1409 -1218 1410 -1217
rect 1437 -1218 1438 -1217
rect 1654 -1218 1655 -1217
rect 163 -1220 164 -1219
rect 1192 -1220 1193 -1219
rect 1213 -1220 1214 -1219
rect 1241 -1220 1242 -1219
rect 1290 -1220 1291 -1219
rect 1437 -1220 1438 -1219
rect 166 -1222 167 -1221
rect 485 -1222 486 -1221
rect 492 -1222 493 -1221
rect 779 -1222 780 -1221
rect 814 -1222 815 -1221
rect 1640 -1222 1641 -1221
rect 166 -1224 167 -1223
rect 464 -1224 465 -1223
rect 492 -1224 493 -1223
rect 639 -1224 640 -1223
rect 674 -1224 675 -1223
rect 716 -1224 717 -1223
rect 768 -1224 769 -1223
rect 1696 -1224 1697 -1223
rect 184 -1226 185 -1225
rect 688 -1226 689 -1225
rect 695 -1226 696 -1225
rect 978 -1226 979 -1225
rect 982 -1226 983 -1225
rect 999 -1226 1000 -1225
rect 1013 -1226 1014 -1225
rect 1367 -1226 1368 -1225
rect 1374 -1226 1375 -1225
rect 1640 -1226 1641 -1225
rect 82 -1228 83 -1227
rect 184 -1228 185 -1227
rect 198 -1228 199 -1227
rect 467 -1228 468 -1227
rect 513 -1228 514 -1227
rect 1500 -1228 1501 -1227
rect 198 -1230 199 -1229
rect 625 -1230 626 -1229
rect 639 -1230 640 -1229
rect 653 -1230 654 -1229
rect 709 -1230 710 -1229
rect 719 -1230 720 -1229
rect 772 -1230 773 -1229
rect 835 -1230 836 -1229
rect 894 -1230 895 -1229
rect 912 -1230 913 -1229
rect 936 -1230 937 -1229
rect 1626 -1230 1627 -1229
rect 156 -1232 157 -1231
rect 625 -1232 626 -1231
rect 646 -1232 647 -1231
rect 674 -1232 675 -1231
rect 828 -1232 829 -1231
rect 1514 -1232 1515 -1231
rect 1535 -1232 1536 -1231
rect 1626 -1232 1627 -1231
rect 156 -1234 157 -1233
rect 618 -1234 619 -1233
rect 646 -1234 647 -1233
rect 663 -1234 664 -1233
rect 831 -1234 832 -1233
rect 940 -1234 941 -1233
rect 957 -1234 958 -1233
rect 1577 -1234 1578 -1233
rect 233 -1236 234 -1235
rect 331 -1236 332 -1235
rect 352 -1236 353 -1235
rect 450 -1236 451 -1235
rect 478 -1236 479 -1235
rect 772 -1236 773 -1235
rect 884 -1236 885 -1235
rect 940 -1236 941 -1235
rect 971 -1236 972 -1235
rect 1584 -1236 1585 -1235
rect 212 -1238 213 -1237
rect 331 -1238 332 -1237
rect 387 -1238 388 -1237
rect 499 -1238 500 -1237
rect 576 -1238 577 -1237
rect 1528 -1238 1529 -1237
rect 191 -1240 192 -1239
rect 212 -1240 213 -1239
rect 233 -1240 234 -1239
rect 499 -1240 500 -1239
rect 597 -1240 598 -1239
rect 1577 -1240 1578 -1239
rect 177 -1242 178 -1241
rect 191 -1242 192 -1241
rect 236 -1242 237 -1241
rect 1451 -1242 1452 -1241
rect 1472 -1242 1473 -1241
rect 1535 -1242 1536 -1241
rect 177 -1244 178 -1243
rect 219 -1244 220 -1243
rect 240 -1244 241 -1243
rect 618 -1244 619 -1243
rect 653 -1244 654 -1243
rect 950 -1244 951 -1243
rect 975 -1244 976 -1243
rect 1192 -1244 1193 -1243
rect 1276 -1244 1277 -1243
rect 1290 -1244 1291 -1243
rect 1356 -1244 1357 -1243
rect 1584 -1244 1585 -1243
rect 219 -1246 220 -1245
rect 817 -1246 818 -1245
rect 821 -1246 822 -1245
rect 884 -1246 885 -1245
rect 898 -1246 899 -1245
rect 905 -1246 906 -1245
rect 975 -1246 976 -1245
rect 992 -1246 993 -1245
rect 1045 -1246 1046 -1245
rect 1556 -1246 1557 -1245
rect 152 -1248 153 -1247
rect 905 -1248 906 -1247
rect 982 -1248 983 -1247
rect 1262 -1248 1263 -1247
rect 1381 -1248 1382 -1247
rect 1570 -1248 1571 -1247
rect 240 -1250 241 -1249
rect 621 -1250 622 -1249
rect 821 -1250 822 -1249
rect 1010 -1250 1011 -1249
rect 1031 -1250 1032 -1249
rect 1262 -1250 1263 -1249
rect 1395 -1250 1396 -1249
rect 1734 -1250 1735 -1249
rect 254 -1252 255 -1251
rect 345 -1252 346 -1251
rect 394 -1252 395 -1251
rect 464 -1252 465 -1251
rect 478 -1252 479 -1251
rect 527 -1252 528 -1251
rect 544 -1252 545 -1251
rect 1381 -1252 1382 -1251
rect 1423 -1252 1424 -1251
rect 1472 -1252 1473 -1251
rect 1556 -1252 1557 -1251
rect 1647 -1252 1648 -1251
rect 37 -1254 38 -1253
rect 527 -1254 528 -1253
rect 562 -1254 563 -1253
rect 597 -1254 598 -1253
rect 611 -1254 612 -1253
rect 691 -1254 692 -1253
rect 989 -1254 990 -1253
rect 1059 -1254 1060 -1253
rect 1080 -1254 1081 -1253
rect 1367 -1254 1368 -1253
rect 1388 -1254 1389 -1253
rect 1423 -1254 1424 -1253
rect 1612 -1254 1613 -1253
rect 1647 -1254 1648 -1253
rect 37 -1256 38 -1255
rect 548 -1256 549 -1255
rect 614 -1256 615 -1255
rect 1591 -1256 1592 -1255
rect 278 -1258 279 -1257
rect 807 -1258 808 -1257
rect 989 -1258 990 -1257
rect 1087 -1258 1088 -1257
rect 1108 -1258 1109 -1257
rect 1339 -1258 1340 -1257
rect 1549 -1258 1550 -1257
rect 1612 -1258 1613 -1257
rect 310 -1260 311 -1259
rect 509 -1260 510 -1259
rect 548 -1260 549 -1259
rect 555 -1260 556 -1259
rect 751 -1260 752 -1259
rect 1388 -1260 1389 -1259
rect 1493 -1260 1494 -1259
rect 1549 -1260 1550 -1259
rect 310 -1262 311 -1261
rect 460 -1262 461 -1261
rect 471 -1262 472 -1261
rect 562 -1262 563 -1261
rect 751 -1262 752 -1261
rect 758 -1262 759 -1261
rect 807 -1262 808 -1261
rect 1115 -1262 1116 -1261
rect 1129 -1262 1130 -1261
rect 1227 -1262 1228 -1261
rect 1255 -1262 1256 -1261
rect 1493 -1262 1494 -1261
rect 317 -1264 318 -1263
rect 726 -1264 727 -1263
rect 1003 -1264 1004 -1263
rect 1059 -1264 1060 -1263
rect 1108 -1264 1109 -1263
rect 1353 -1264 1354 -1263
rect 282 -1266 283 -1265
rect 317 -1266 318 -1265
rect 324 -1266 325 -1265
rect 359 -1266 360 -1265
rect 394 -1266 395 -1265
rect 870 -1266 871 -1265
rect 1003 -1266 1004 -1265
rect 1234 -1266 1235 -1265
rect 1353 -1266 1354 -1265
rect 1374 -1266 1375 -1265
rect 170 -1268 171 -1267
rect 324 -1268 325 -1267
rect 345 -1268 346 -1267
rect 408 -1268 409 -1267
rect 429 -1268 430 -1267
rect 516 -1268 517 -1267
rect 555 -1268 556 -1267
rect 831 -1268 832 -1267
rect 870 -1268 871 -1267
rect 1017 -1268 1018 -1267
rect 1024 -1268 1025 -1267
rect 1087 -1268 1088 -1267
rect 1143 -1268 1144 -1267
rect 1213 -1268 1214 -1267
rect 1220 -1268 1221 -1267
rect 1276 -1268 1277 -1267
rect 170 -1270 171 -1269
rect 604 -1270 605 -1269
rect 877 -1270 878 -1269
rect 1220 -1270 1221 -1269
rect 282 -1272 283 -1271
rect 985 -1272 986 -1271
rect 996 -1272 997 -1271
rect 1024 -1272 1025 -1271
rect 1045 -1272 1046 -1271
rect 1164 -1272 1165 -1271
rect 1171 -1272 1172 -1271
rect 1255 -1272 1256 -1271
rect 338 -1274 339 -1273
rect 429 -1274 430 -1273
rect 443 -1274 444 -1273
rect 446 -1274 447 -1273
rect 450 -1274 451 -1273
rect 583 -1274 584 -1273
rect 590 -1274 591 -1273
rect 877 -1274 878 -1273
rect 933 -1274 934 -1273
rect 996 -1274 997 -1273
rect 1010 -1274 1011 -1273
rect 1080 -1274 1081 -1273
rect 1094 -1274 1095 -1273
rect 1171 -1274 1172 -1273
rect 1199 -1274 1200 -1273
rect 1227 -1274 1228 -1273
rect 86 -1276 87 -1275
rect 583 -1276 584 -1275
rect 933 -1276 934 -1275
rect 1066 -1276 1067 -1275
rect 1094 -1276 1095 -1275
rect 1157 -1276 1158 -1275
rect 1164 -1276 1165 -1275
rect 1178 -1276 1179 -1275
rect 261 -1278 262 -1277
rect 338 -1278 339 -1277
rect 408 -1278 409 -1277
rect 415 -1278 416 -1277
rect 443 -1278 444 -1277
rect 520 -1278 521 -1277
rect 534 -1278 535 -1277
rect 604 -1278 605 -1277
rect 947 -1278 948 -1277
rect 1017 -1278 1018 -1277
rect 1048 -1278 1049 -1277
rect 1430 -1278 1431 -1277
rect 44 -1280 45 -1279
rect 534 -1280 535 -1279
rect 569 -1280 570 -1279
rect 758 -1280 759 -1279
rect 947 -1280 948 -1279
rect 1713 -1280 1714 -1279
rect 44 -1282 45 -1281
rect 75 -1282 76 -1281
rect 226 -1282 227 -1281
rect 569 -1282 570 -1281
rect 954 -1282 955 -1281
rect 1234 -1282 1235 -1281
rect 1360 -1282 1361 -1281
rect 1430 -1282 1431 -1281
rect 75 -1284 76 -1283
rect 86 -1284 87 -1283
rect 226 -1284 227 -1283
rect 457 -1284 458 -1283
rect 471 -1284 472 -1283
rect 747 -1284 748 -1283
rect 863 -1284 864 -1283
rect 954 -1284 955 -1283
rect 961 -1284 962 -1283
rect 1066 -1284 1067 -1283
rect 1101 -1284 1102 -1283
rect 1143 -1284 1144 -1283
rect 1150 -1284 1151 -1283
rect 1199 -1284 1200 -1283
rect 1304 -1284 1305 -1283
rect 1360 -1284 1361 -1283
rect 261 -1286 262 -1285
rect 422 -1286 423 -1285
rect 425 -1286 426 -1285
rect 1304 -1286 1305 -1285
rect 415 -1288 416 -1287
rect 681 -1288 682 -1287
rect 702 -1288 703 -1287
rect 961 -1288 962 -1287
rect 968 -1288 969 -1287
rect 1178 -1288 1179 -1287
rect 366 -1290 367 -1289
rect 681 -1290 682 -1289
rect 800 -1290 801 -1289
rect 863 -1290 864 -1289
rect 919 -1290 920 -1289
rect 968 -1290 969 -1289
rect 999 -1290 1000 -1289
rect 1031 -1290 1032 -1289
rect 1038 -1290 1039 -1289
rect 1150 -1290 1151 -1289
rect 1157 -1290 1158 -1289
rect 1283 -1290 1284 -1289
rect 128 -1292 129 -1291
rect 800 -1292 801 -1291
rect 842 -1292 843 -1291
rect 1101 -1292 1102 -1291
rect 107 -1294 108 -1293
rect 128 -1294 129 -1293
rect 303 -1294 304 -1293
rect 366 -1294 367 -1293
rect 509 -1294 510 -1293
rect 667 -1294 668 -1293
rect 842 -1294 843 -1293
rect 856 -1294 857 -1293
rect 1052 -1294 1053 -1293
rect 1122 -1294 1123 -1293
rect 107 -1296 108 -1295
rect 268 -1296 269 -1295
rect 303 -1296 304 -1295
rect 401 -1296 402 -1295
rect 628 -1296 629 -1295
rect 667 -1296 668 -1295
rect 828 -1296 829 -1295
rect 856 -1296 857 -1295
rect 1052 -1296 1053 -1295
rect 1563 -1296 1564 -1295
rect 114 -1298 115 -1297
rect 401 -1298 402 -1297
rect 632 -1298 633 -1297
rect 702 -1298 703 -1297
rect 849 -1298 850 -1297
rect 919 -1298 920 -1297
rect 1055 -1298 1056 -1297
rect 1311 -1298 1312 -1297
rect 1507 -1298 1508 -1297
rect 1563 -1298 1564 -1297
rect 114 -1300 115 -1299
rect 688 -1300 689 -1299
rect 765 -1300 766 -1299
rect 849 -1300 850 -1299
rect 1073 -1300 1074 -1299
rect 1283 -1300 1284 -1299
rect 1311 -1300 1312 -1299
rect 1346 -1300 1347 -1299
rect 1458 -1300 1459 -1299
rect 1507 -1300 1508 -1299
rect 268 -1302 269 -1301
rect 289 -1302 290 -1301
rect 373 -1302 374 -1301
rect 632 -1302 633 -1301
rect 660 -1302 661 -1301
rect 1038 -1302 1039 -1301
rect 1458 -1302 1459 -1301
rect 1664 -1302 1665 -1301
rect 51 -1304 52 -1303
rect 289 -1304 290 -1303
rect 373 -1304 374 -1303
rect 436 -1304 437 -1303
rect 660 -1304 661 -1303
rect 737 -1304 738 -1303
rect 765 -1304 766 -1303
rect 912 -1304 913 -1303
rect 51 -1306 52 -1305
rect 614 -1306 615 -1305
rect 730 -1306 731 -1305
rect 737 -1306 738 -1305
rect 786 -1306 787 -1305
rect 1073 -1306 1074 -1305
rect 257 -1308 258 -1307
rect 436 -1308 437 -1307
rect 481 -1308 482 -1307
rect 730 -1308 731 -1307
rect 786 -1308 787 -1307
rect 1248 -1308 1249 -1307
rect 891 -1310 892 -1309
rect 1346 -1310 1347 -1309
rect 891 -1312 892 -1311
rect 926 -1312 927 -1311
rect 1248 -1312 1249 -1311
rect 1332 -1312 1333 -1311
rect 82 -1314 83 -1313
rect 926 -1314 927 -1313
rect 1269 -1314 1270 -1313
rect 1332 -1314 1333 -1313
rect 93 -1316 94 -1315
rect 1269 -1316 1270 -1315
rect 16 -1327 17 -1326
rect 51 -1327 52 -1326
rect 58 -1327 59 -1326
rect 422 -1327 423 -1326
rect 478 -1327 479 -1326
rect 1374 -1327 1375 -1326
rect 1493 -1327 1494 -1326
rect 1731 -1327 1732 -1326
rect 1738 -1327 1739 -1326
rect 1745 -1327 1746 -1326
rect 37 -1329 38 -1328
rect 422 -1329 423 -1328
rect 478 -1329 479 -1328
rect 520 -1329 521 -1328
rect 579 -1329 580 -1328
rect 1276 -1329 1277 -1328
rect 1346 -1329 1347 -1328
rect 1706 -1329 1707 -1328
rect 1717 -1329 1718 -1328
rect 1734 -1329 1735 -1328
rect 37 -1331 38 -1330
rect 229 -1331 230 -1330
rect 233 -1331 234 -1330
rect 282 -1331 283 -1330
rect 289 -1331 290 -1330
rect 527 -1331 528 -1330
rect 597 -1331 598 -1330
rect 765 -1331 766 -1330
rect 768 -1331 769 -1330
rect 1171 -1331 1172 -1330
rect 1276 -1331 1277 -1330
rect 1360 -1331 1361 -1330
rect 1493 -1331 1494 -1330
rect 1521 -1331 1522 -1330
rect 1626 -1331 1627 -1330
rect 1720 -1331 1721 -1330
rect 44 -1333 45 -1332
rect 72 -1333 73 -1332
rect 82 -1333 83 -1332
rect 1297 -1333 1298 -1332
rect 1521 -1333 1522 -1332
rect 1591 -1333 1592 -1332
rect 1675 -1333 1676 -1332
rect 1703 -1333 1704 -1332
rect 44 -1335 45 -1334
rect 198 -1335 199 -1334
rect 240 -1335 241 -1334
rect 831 -1335 832 -1334
rect 873 -1335 874 -1334
rect 1423 -1335 1424 -1334
rect 1584 -1335 1585 -1334
rect 1626 -1335 1627 -1334
rect 1682 -1335 1683 -1334
rect 1717 -1335 1718 -1334
rect 51 -1337 52 -1336
rect 625 -1337 626 -1336
rect 628 -1337 629 -1336
rect 779 -1337 780 -1336
rect 786 -1337 787 -1336
rect 842 -1337 843 -1336
rect 901 -1337 902 -1336
rect 1094 -1337 1095 -1336
rect 1125 -1337 1126 -1336
rect 1591 -1337 1592 -1336
rect 1696 -1337 1697 -1336
rect 1710 -1337 1711 -1336
rect 75 -1339 76 -1338
rect 240 -1339 241 -1338
rect 250 -1339 251 -1338
rect 1304 -1339 1305 -1338
rect 1699 -1339 1700 -1338
rect 1724 -1339 1725 -1338
rect 82 -1341 83 -1340
rect 1339 -1341 1340 -1340
rect 86 -1343 87 -1342
rect 96 -1343 97 -1342
rect 124 -1343 125 -1342
rect 149 -1343 150 -1342
rect 170 -1343 171 -1342
rect 733 -1343 734 -1342
rect 765 -1343 766 -1342
rect 1374 -1343 1375 -1342
rect 93 -1345 94 -1344
rect 1262 -1345 1263 -1344
rect 1283 -1345 1284 -1344
rect 1675 -1345 1676 -1344
rect 96 -1347 97 -1346
rect 324 -1347 325 -1346
rect 366 -1347 367 -1346
rect 576 -1347 577 -1346
rect 590 -1347 591 -1346
rect 625 -1347 626 -1346
rect 632 -1347 633 -1346
rect 786 -1347 787 -1346
rect 796 -1347 797 -1346
rect 1360 -1347 1361 -1346
rect 107 -1349 108 -1348
rect 170 -1349 171 -1348
rect 177 -1349 178 -1348
rect 236 -1349 237 -1348
rect 264 -1349 265 -1348
rect 317 -1349 318 -1348
rect 324 -1349 325 -1348
rect 541 -1349 542 -1348
rect 548 -1349 549 -1348
rect 576 -1349 577 -1348
rect 597 -1349 598 -1348
rect 1101 -1349 1102 -1348
rect 1136 -1349 1137 -1348
rect 1724 -1349 1725 -1348
rect 107 -1351 108 -1350
rect 1507 -1351 1508 -1350
rect 135 -1353 136 -1352
rect 457 -1353 458 -1352
rect 460 -1353 461 -1352
rect 1346 -1353 1347 -1352
rect 135 -1355 136 -1354
rect 502 -1355 503 -1354
rect 506 -1355 507 -1354
rect 632 -1355 633 -1354
rect 653 -1355 654 -1354
rect 817 -1355 818 -1354
rect 821 -1355 822 -1354
rect 1192 -1355 1193 -1354
rect 1262 -1355 1263 -1354
rect 1318 -1355 1319 -1354
rect 1339 -1355 1340 -1354
rect 1549 -1355 1550 -1354
rect 142 -1357 143 -1356
rect 807 -1357 808 -1356
rect 828 -1357 829 -1356
rect 1640 -1357 1641 -1356
rect 30 -1359 31 -1358
rect 142 -1359 143 -1358
rect 149 -1359 150 -1358
rect 562 -1359 563 -1358
rect 593 -1359 594 -1358
rect 1640 -1359 1641 -1358
rect 26 -1361 27 -1360
rect 30 -1361 31 -1360
rect 177 -1361 178 -1360
rect 184 -1361 185 -1360
rect 191 -1361 192 -1360
rect 198 -1361 199 -1360
rect 219 -1361 220 -1360
rect 506 -1361 507 -1360
rect 520 -1361 521 -1360
rect 891 -1361 892 -1360
rect 947 -1361 948 -1360
rect 1542 -1361 1543 -1360
rect 117 -1363 118 -1362
rect 1542 -1363 1543 -1362
rect 163 -1365 164 -1364
rect 184 -1365 185 -1364
rect 219 -1365 220 -1364
rect 254 -1365 255 -1364
rect 275 -1365 276 -1364
rect 450 -1365 451 -1364
rect 457 -1365 458 -1364
rect 730 -1365 731 -1364
rect 779 -1365 780 -1364
rect 835 -1365 836 -1364
rect 891 -1365 892 -1364
rect 989 -1365 990 -1364
rect 1010 -1365 1011 -1364
rect 1213 -1365 1214 -1364
rect 1297 -1365 1298 -1364
rect 1311 -1365 1312 -1364
rect 114 -1367 115 -1366
rect 254 -1367 255 -1366
rect 275 -1367 276 -1366
rect 331 -1367 332 -1366
rect 366 -1367 367 -1366
rect 691 -1367 692 -1366
rect 695 -1367 696 -1366
rect 894 -1367 895 -1366
rect 947 -1367 948 -1366
rect 968 -1367 969 -1366
rect 978 -1367 979 -1366
rect 1612 -1367 1613 -1366
rect 156 -1369 157 -1368
rect 163 -1369 164 -1368
rect 247 -1369 248 -1368
rect 1318 -1369 1319 -1368
rect 1612 -1369 1613 -1368
rect 1633 -1369 1634 -1368
rect 156 -1371 157 -1370
rect 191 -1371 192 -1370
rect 247 -1371 248 -1370
rect 278 -1371 279 -1370
rect 282 -1371 283 -1370
rect 345 -1371 346 -1370
rect 373 -1371 374 -1370
rect 1507 -1371 1508 -1370
rect 1605 -1371 1606 -1370
rect 1633 -1371 1634 -1370
rect 289 -1373 290 -1372
rect 418 -1373 419 -1372
rect 436 -1373 437 -1372
rect 541 -1373 542 -1372
rect 548 -1373 549 -1372
rect 555 -1373 556 -1372
rect 562 -1373 563 -1372
rect 604 -1373 605 -1372
rect 614 -1373 615 -1372
rect 821 -1373 822 -1372
rect 828 -1373 829 -1372
rect 863 -1373 864 -1372
rect 968 -1373 969 -1372
rect 1024 -1373 1025 -1372
rect 1027 -1373 1028 -1372
rect 1584 -1373 1585 -1372
rect 296 -1375 297 -1374
rect 611 -1375 612 -1374
rect 618 -1375 619 -1374
rect 663 -1375 664 -1374
rect 667 -1375 668 -1374
rect 989 -1375 990 -1374
rect 1045 -1375 1046 -1374
rect 1048 -1375 1049 -1374
rect 1055 -1375 1056 -1374
rect 1332 -1375 1333 -1374
rect 1416 -1375 1417 -1374
rect 1605 -1375 1606 -1374
rect 303 -1377 304 -1376
rect 345 -1377 346 -1376
rect 352 -1377 353 -1376
rect 614 -1377 615 -1376
rect 639 -1377 640 -1376
rect 667 -1377 668 -1376
rect 688 -1377 689 -1376
rect 1479 -1377 1480 -1376
rect 317 -1379 318 -1378
rect 789 -1379 790 -1378
rect 835 -1379 836 -1378
rect 936 -1379 937 -1378
rect 982 -1379 983 -1378
rect 1416 -1379 1417 -1378
rect 1479 -1379 1480 -1378
rect 1514 -1379 1515 -1378
rect 331 -1381 332 -1380
rect 499 -1381 500 -1380
rect 590 -1381 591 -1380
rect 1514 -1381 1515 -1380
rect 352 -1383 353 -1382
rect 408 -1383 409 -1382
rect 415 -1383 416 -1382
rect 436 -1383 437 -1382
rect 450 -1383 451 -1382
rect 772 -1383 773 -1382
rect 863 -1383 864 -1382
rect 1108 -1383 1109 -1382
rect 1129 -1383 1130 -1382
rect 1192 -1383 1193 -1382
rect 1213 -1383 1214 -1382
rect 1255 -1383 1256 -1382
rect 1304 -1383 1305 -1382
rect 1409 -1383 1410 -1382
rect 338 -1385 339 -1384
rect 408 -1385 409 -1384
rect 415 -1385 416 -1384
rect 534 -1385 535 -1384
rect 604 -1385 605 -1384
rect 635 -1385 636 -1384
rect 639 -1385 640 -1384
rect 1073 -1385 1074 -1384
rect 1094 -1385 1095 -1384
rect 1206 -1385 1207 -1384
rect 1255 -1385 1256 -1384
rect 1402 -1385 1403 -1384
rect 261 -1387 262 -1386
rect 338 -1387 339 -1386
rect 373 -1387 374 -1386
rect 583 -1387 584 -1386
rect 611 -1387 612 -1386
rect 1423 -1387 1424 -1386
rect 261 -1389 262 -1388
rect 1101 -1389 1102 -1388
rect 1146 -1389 1147 -1388
rect 1654 -1389 1655 -1388
rect 387 -1391 388 -1390
rect 527 -1391 528 -1390
rect 534 -1391 535 -1390
rect 856 -1391 857 -1390
rect 877 -1391 878 -1390
rect 936 -1391 937 -1390
rect 940 -1391 941 -1390
rect 982 -1391 983 -1390
rect 985 -1391 986 -1390
rect 1689 -1391 1690 -1390
rect 303 -1393 304 -1392
rect 387 -1393 388 -1392
rect 394 -1393 395 -1392
rect 1010 -1393 1011 -1392
rect 1017 -1393 1018 -1392
rect 1108 -1393 1109 -1392
rect 1171 -1393 1172 -1392
rect 1241 -1393 1242 -1392
rect 1311 -1393 1312 -1392
rect 1444 -1393 1445 -1392
rect 1654 -1393 1655 -1392
rect 1661 -1393 1662 -1392
rect 205 -1395 206 -1394
rect 394 -1395 395 -1394
rect 401 -1395 402 -1394
rect 842 -1395 843 -1394
rect 877 -1395 878 -1394
rect 898 -1395 899 -1394
rect 905 -1395 906 -1394
rect 1073 -1395 1074 -1394
rect 1139 -1395 1140 -1394
rect 1241 -1395 1242 -1394
rect 1325 -1395 1326 -1394
rect 1409 -1395 1410 -1394
rect 79 -1397 80 -1396
rect 898 -1397 899 -1396
rect 940 -1397 941 -1396
rect 961 -1397 962 -1396
rect 1017 -1397 1018 -1396
rect 1066 -1397 1067 -1396
rect 1069 -1397 1070 -1396
rect 1647 -1397 1648 -1396
rect 110 -1399 111 -1398
rect 205 -1399 206 -1398
rect 401 -1399 402 -1398
rect 443 -1399 444 -1398
rect 464 -1399 465 -1398
rect 618 -1399 619 -1398
rect 653 -1399 654 -1398
rect 709 -1399 710 -1398
rect 719 -1399 720 -1398
rect 954 -1399 955 -1398
rect 1045 -1399 1046 -1398
rect 1087 -1399 1088 -1398
rect 1185 -1399 1186 -1398
rect 1283 -1399 1284 -1398
rect 1332 -1399 1333 -1398
rect 1388 -1399 1389 -1398
rect 1402 -1399 1403 -1398
rect 1458 -1399 1459 -1398
rect 1619 -1399 1620 -1398
rect 1647 -1399 1648 -1398
rect 121 -1401 122 -1400
rect 1388 -1401 1389 -1400
rect 1458 -1401 1459 -1400
rect 1486 -1401 1487 -1400
rect 121 -1403 122 -1402
rect 380 -1403 381 -1402
rect 464 -1403 465 -1402
rect 646 -1403 647 -1402
rect 660 -1403 661 -1402
rect 1220 -1403 1221 -1402
rect 1353 -1403 1354 -1402
rect 1661 -1403 1662 -1402
rect 128 -1405 129 -1404
rect 646 -1405 647 -1404
rect 660 -1405 661 -1404
rect 975 -1405 976 -1404
rect 1087 -1405 1088 -1404
rect 1150 -1405 1151 -1404
rect 1185 -1405 1186 -1404
rect 1381 -1405 1382 -1404
rect 1486 -1405 1487 -1404
rect 1528 -1405 1529 -1404
rect 128 -1407 129 -1406
rect 359 -1407 360 -1406
rect 380 -1407 381 -1406
rect 429 -1407 430 -1406
rect 485 -1407 486 -1406
rect 726 -1407 727 -1406
rect 730 -1407 731 -1406
rect 1549 -1407 1550 -1406
rect 23 -1409 24 -1408
rect 485 -1409 486 -1408
rect 499 -1409 500 -1408
rect 1619 -1409 1620 -1408
rect 65 -1411 66 -1410
rect 429 -1411 430 -1410
rect 513 -1411 514 -1410
rect 1066 -1411 1067 -1410
rect 1206 -1411 1207 -1410
rect 1290 -1411 1291 -1410
rect 1353 -1411 1354 -1410
rect 1437 -1411 1438 -1410
rect 1528 -1411 1529 -1410
rect 1570 -1411 1571 -1410
rect 65 -1413 66 -1412
rect 222 -1413 223 -1412
rect 226 -1413 227 -1412
rect 443 -1413 444 -1412
rect 555 -1413 556 -1412
rect 1689 -1413 1690 -1412
rect 310 -1415 311 -1414
rect 359 -1415 360 -1414
rect 583 -1415 584 -1414
rect 1013 -1415 1014 -1414
rect 1048 -1415 1049 -1414
rect 1150 -1415 1151 -1414
rect 1157 -1415 1158 -1414
rect 1290 -1415 1291 -1414
rect 310 -1417 311 -1416
rect 471 -1417 472 -1416
rect 677 -1417 678 -1416
rect 1220 -1417 1221 -1416
rect 1248 -1417 1249 -1416
rect 1381 -1417 1382 -1416
rect 58 -1419 59 -1418
rect 471 -1419 472 -1418
rect 688 -1419 689 -1418
rect 702 -1419 703 -1418
rect 709 -1419 710 -1418
rect 716 -1419 717 -1418
rect 723 -1419 724 -1418
rect 793 -1419 794 -1418
rect 800 -1419 801 -1418
rect 1129 -1419 1130 -1418
rect 1248 -1419 1249 -1418
rect 1395 -1419 1396 -1418
rect 695 -1421 696 -1420
rect 758 -1421 759 -1420
rect 800 -1421 801 -1420
rect 849 -1421 850 -1420
rect 866 -1421 867 -1420
rect 1570 -1421 1571 -1420
rect 702 -1423 703 -1422
rect 1031 -1423 1032 -1422
rect 1395 -1423 1396 -1422
rect 1451 -1423 1452 -1422
rect 61 -1425 62 -1424
rect 1031 -1425 1032 -1424
rect 1430 -1425 1431 -1424
rect 1451 -1425 1452 -1424
rect 716 -1427 717 -1426
rect 1157 -1427 1158 -1426
rect 1430 -1427 1431 -1426
rect 1465 -1427 1466 -1426
rect 226 -1429 227 -1428
rect 1465 -1429 1466 -1428
rect 723 -1431 724 -1430
rect 1367 -1431 1368 -1430
rect 744 -1433 745 -1432
rect 793 -1433 794 -1432
rect 814 -1433 815 -1432
rect 905 -1433 906 -1432
rect 919 -1433 920 -1432
rect 961 -1433 962 -1432
rect 975 -1433 976 -1432
rect 996 -1433 997 -1432
rect 1367 -1433 1368 -1432
rect 1472 -1433 1473 -1432
rect 737 -1435 738 -1434
rect 744 -1435 745 -1434
rect 751 -1435 752 -1434
rect 772 -1435 773 -1434
rect 814 -1435 815 -1434
rect 884 -1435 885 -1434
rect 919 -1435 920 -1434
rect 1059 -1435 1060 -1434
rect 1472 -1435 1473 -1434
rect 1500 -1435 1501 -1434
rect 145 -1437 146 -1436
rect 751 -1437 752 -1436
rect 758 -1437 759 -1436
rect 870 -1437 871 -1436
rect 933 -1437 934 -1436
rect 1437 -1437 1438 -1436
rect 1500 -1437 1501 -1436
rect 1535 -1437 1536 -1436
rect 569 -1439 570 -1438
rect 737 -1439 738 -1438
rect 824 -1439 825 -1438
rect 1444 -1439 1445 -1438
rect 1535 -1439 1536 -1438
rect 1577 -1439 1578 -1438
rect 509 -1441 510 -1440
rect 569 -1441 570 -1440
rect 681 -1441 682 -1440
rect 884 -1441 885 -1440
rect 933 -1441 934 -1440
rect 1682 -1441 1683 -1440
rect 674 -1443 675 -1442
rect 681 -1443 682 -1442
rect 849 -1443 850 -1442
rect 926 -1443 927 -1442
rect 954 -1443 955 -1442
rect 1143 -1443 1144 -1442
rect 1577 -1443 1578 -1442
rect 1598 -1443 1599 -1442
rect 492 -1445 493 -1444
rect 674 -1445 675 -1444
rect 856 -1445 857 -1444
rect 870 -1445 871 -1444
rect 926 -1445 927 -1444
rect 1003 -1445 1004 -1444
rect 1059 -1445 1060 -1444
rect 1122 -1445 1123 -1444
rect 1143 -1445 1144 -1444
rect 1325 -1445 1326 -1444
rect 1563 -1445 1564 -1444
rect 1598 -1445 1599 -1444
rect 86 -1447 87 -1446
rect 1122 -1447 1123 -1446
rect 1227 -1447 1228 -1446
rect 1563 -1447 1564 -1446
rect 93 -1449 94 -1448
rect 492 -1449 493 -1448
rect 530 -1449 531 -1448
rect 1227 -1449 1228 -1448
rect 996 -1451 997 -1450
rect 1038 -1451 1039 -1450
rect 1003 -1453 1004 -1452
rect 1199 -1453 1200 -1452
rect 600 -1455 601 -1454
rect 1199 -1455 1200 -1454
rect 1038 -1457 1039 -1456
rect 1115 -1457 1116 -1456
rect 1115 -1459 1116 -1458
rect 1164 -1459 1165 -1458
rect 1164 -1461 1165 -1460
rect 1234 -1461 1235 -1460
rect 1080 -1463 1081 -1462
rect 1234 -1463 1235 -1462
rect 1080 -1465 1081 -1464
rect 1178 -1465 1179 -1464
rect 1052 -1467 1053 -1466
rect 1178 -1467 1179 -1466
rect 912 -1469 913 -1468
rect 1052 -1469 1053 -1468
rect 642 -1471 643 -1470
rect 912 -1471 913 -1470
rect 16 -1482 17 -1481
rect 765 -1482 766 -1481
rect 786 -1482 787 -1481
rect 863 -1482 864 -1481
rect 870 -1482 871 -1481
rect 919 -1482 920 -1481
rect 1024 -1482 1025 -1481
rect 1094 -1482 1095 -1481
rect 1104 -1482 1105 -1481
rect 1339 -1482 1340 -1481
rect 1745 -1482 1746 -1481
rect 1752 -1482 1753 -1481
rect 23 -1484 24 -1483
rect 75 -1484 76 -1483
rect 96 -1484 97 -1483
rect 1640 -1484 1641 -1483
rect 30 -1486 31 -1485
rect 82 -1486 83 -1485
rect 107 -1486 108 -1485
rect 415 -1486 416 -1485
rect 418 -1486 419 -1485
rect 765 -1486 766 -1485
rect 786 -1486 787 -1485
rect 905 -1486 906 -1485
rect 1024 -1486 1025 -1485
rect 1087 -1486 1088 -1485
rect 1118 -1486 1119 -1485
rect 1710 -1486 1711 -1485
rect 58 -1488 59 -1487
rect 1689 -1488 1690 -1487
rect 61 -1490 62 -1489
rect 117 -1490 118 -1489
rect 142 -1490 143 -1489
rect 208 -1490 209 -1489
rect 226 -1490 227 -1489
rect 359 -1490 360 -1489
rect 373 -1490 374 -1489
rect 761 -1490 762 -1489
rect 863 -1490 864 -1489
rect 940 -1490 941 -1489
rect 1073 -1490 1074 -1489
rect 1713 -1490 1714 -1489
rect 68 -1492 69 -1491
rect 548 -1492 549 -1491
rect 555 -1492 556 -1491
rect 611 -1492 612 -1491
rect 621 -1492 622 -1491
rect 709 -1492 710 -1491
rect 719 -1492 720 -1491
rect 1563 -1492 1564 -1491
rect 1640 -1492 1641 -1491
rect 1668 -1492 1669 -1491
rect 72 -1494 73 -1493
rect 366 -1494 367 -1493
rect 390 -1494 391 -1493
rect 429 -1494 430 -1493
rect 443 -1494 444 -1493
rect 544 -1494 545 -1493
rect 562 -1494 563 -1493
rect 709 -1494 710 -1493
rect 733 -1494 734 -1493
rect 919 -1494 920 -1493
rect 1073 -1494 1074 -1493
rect 1143 -1494 1144 -1493
rect 1153 -1494 1154 -1493
rect 1332 -1494 1333 -1493
rect 1339 -1494 1340 -1493
rect 1416 -1494 1417 -1493
rect 1493 -1494 1494 -1493
rect 1689 -1494 1690 -1493
rect 44 -1496 45 -1495
rect 72 -1496 73 -1495
rect 107 -1496 108 -1495
rect 366 -1496 367 -1495
rect 394 -1496 395 -1495
rect 768 -1496 769 -1495
rect 866 -1496 867 -1495
rect 1094 -1496 1095 -1495
rect 1122 -1496 1123 -1495
rect 1262 -1496 1263 -1495
rect 1311 -1496 1312 -1495
rect 1332 -1496 1333 -1495
rect 1416 -1496 1417 -1495
rect 1486 -1496 1487 -1495
rect 1493 -1496 1494 -1495
rect 1535 -1496 1536 -1495
rect 1563 -1496 1564 -1495
rect 1591 -1496 1592 -1495
rect 1612 -1496 1613 -1495
rect 1668 -1496 1669 -1495
rect 44 -1498 45 -1497
rect 369 -1498 370 -1497
rect 394 -1498 395 -1497
rect 471 -1498 472 -1497
rect 474 -1498 475 -1497
rect 961 -1498 962 -1497
rect 989 -1498 990 -1497
rect 1122 -1498 1123 -1497
rect 1125 -1498 1126 -1497
rect 1703 -1498 1704 -1497
rect 30 -1500 31 -1499
rect 471 -1500 472 -1499
rect 492 -1500 493 -1499
rect 901 -1500 902 -1499
rect 905 -1500 906 -1499
rect 926 -1500 927 -1499
rect 961 -1500 962 -1499
rect 968 -1500 969 -1499
rect 975 -1500 976 -1499
rect 989 -1500 990 -1499
rect 1087 -1500 1088 -1499
rect 1171 -1500 1172 -1499
rect 1311 -1500 1312 -1499
rect 1325 -1500 1326 -1499
rect 1486 -1500 1487 -1499
rect 1605 -1500 1606 -1499
rect 114 -1502 115 -1501
rect 436 -1502 437 -1501
rect 443 -1502 444 -1501
rect 1703 -1502 1704 -1501
rect 114 -1504 115 -1503
rect 670 -1504 671 -1503
rect 677 -1504 678 -1503
rect 1549 -1504 1550 -1503
rect 1556 -1504 1557 -1503
rect 1605 -1504 1606 -1503
rect 142 -1506 143 -1505
rect 401 -1506 402 -1505
rect 422 -1506 423 -1505
rect 593 -1506 594 -1505
rect 607 -1506 608 -1505
rect 667 -1506 668 -1505
rect 730 -1506 731 -1505
rect 1262 -1506 1263 -1505
rect 1325 -1506 1326 -1505
rect 1402 -1506 1403 -1505
rect 1500 -1506 1501 -1505
rect 1612 -1506 1613 -1505
rect 51 -1508 52 -1507
rect 401 -1508 402 -1507
rect 436 -1508 437 -1507
rect 929 -1508 930 -1507
rect 975 -1508 976 -1507
rect 1346 -1508 1347 -1507
rect 1402 -1508 1403 -1507
rect 1472 -1508 1473 -1507
rect 1535 -1508 1536 -1507
rect 1577 -1508 1578 -1507
rect 1584 -1508 1585 -1507
rect 1591 -1508 1592 -1507
rect 156 -1510 157 -1509
rect 1556 -1510 1557 -1509
rect 1570 -1510 1571 -1509
rect 1577 -1510 1578 -1509
rect 1584 -1510 1585 -1509
rect 1598 -1510 1599 -1509
rect 156 -1512 157 -1511
rect 212 -1512 213 -1511
rect 226 -1512 227 -1511
rect 257 -1512 258 -1511
rect 261 -1512 262 -1511
rect 282 -1512 283 -1511
rect 296 -1512 297 -1511
rect 618 -1512 619 -1511
rect 632 -1512 633 -1511
rect 1045 -1512 1046 -1511
rect 1048 -1512 1049 -1511
rect 1570 -1512 1571 -1511
rect 1598 -1512 1599 -1511
rect 1619 -1512 1620 -1511
rect 159 -1514 160 -1513
rect 583 -1514 584 -1513
rect 635 -1514 636 -1513
rect 1507 -1514 1508 -1513
rect 1549 -1514 1550 -1513
rect 1720 -1514 1721 -1513
rect 149 -1516 150 -1515
rect 583 -1516 584 -1515
rect 639 -1516 640 -1515
rect 1706 -1516 1707 -1515
rect 149 -1518 150 -1517
rect 558 -1518 559 -1517
rect 562 -1518 563 -1517
rect 681 -1518 682 -1517
rect 712 -1518 713 -1517
rect 1500 -1518 1501 -1517
rect 1619 -1518 1620 -1517
rect 1633 -1518 1634 -1517
rect 191 -1520 192 -1519
rect 219 -1520 220 -1519
rect 229 -1520 230 -1519
rect 982 -1520 983 -1519
rect 1045 -1520 1046 -1519
rect 1129 -1520 1130 -1519
rect 1139 -1520 1140 -1519
rect 1451 -1520 1452 -1519
rect 1472 -1520 1473 -1519
rect 1654 -1520 1655 -1519
rect 194 -1522 195 -1521
rect 534 -1522 535 -1521
rect 541 -1522 542 -1521
rect 555 -1522 556 -1521
rect 576 -1522 577 -1521
rect 597 -1522 598 -1521
rect 604 -1522 605 -1521
rect 681 -1522 682 -1521
rect 730 -1522 731 -1521
rect 779 -1522 780 -1521
rect 796 -1522 797 -1521
rect 1633 -1522 1634 -1521
rect 79 -1524 80 -1523
rect 576 -1524 577 -1523
rect 604 -1524 605 -1523
rect 1682 -1524 1683 -1523
rect 79 -1526 80 -1525
rect 163 -1526 164 -1525
rect 212 -1526 213 -1525
rect 240 -1526 241 -1525
rect 268 -1526 269 -1525
rect 282 -1526 283 -1525
rect 310 -1526 311 -1525
rect 415 -1526 416 -1525
rect 450 -1526 451 -1525
rect 492 -1526 493 -1525
rect 499 -1526 500 -1525
rect 618 -1526 619 -1525
rect 639 -1526 640 -1525
rect 660 -1526 661 -1525
rect 747 -1526 748 -1525
rect 814 -1526 815 -1525
rect 870 -1526 871 -1525
rect 1017 -1526 1018 -1525
rect 1020 -1526 1021 -1525
rect 1654 -1526 1655 -1525
rect 121 -1528 122 -1527
rect 240 -1528 241 -1527
rect 299 -1528 300 -1527
rect 310 -1528 311 -1527
rect 331 -1528 332 -1527
rect 422 -1528 423 -1527
rect 450 -1528 451 -1527
rect 674 -1528 675 -1527
rect 779 -1528 780 -1527
rect 800 -1528 801 -1527
rect 891 -1528 892 -1527
rect 1136 -1528 1137 -1527
rect 1143 -1528 1144 -1527
rect 1206 -1528 1207 -1527
rect 1283 -1528 1284 -1527
rect 1682 -1528 1683 -1527
rect 93 -1530 94 -1529
rect 121 -1530 122 -1529
rect 163 -1530 164 -1529
rect 590 -1530 591 -1529
rect 660 -1530 661 -1529
rect 695 -1530 696 -1529
rect 719 -1530 720 -1529
rect 1283 -1530 1284 -1529
rect 1346 -1530 1347 -1529
rect 1423 -1530 1424 -1529
rect 1451 -1530 1452 -1529
rect 1542 -1530 1543 -1529
rect 93 -1532 94 -1531
rect 625 -1532 626 -1531
rect 674 -1532 675 -1531
rect 737 -1532 738 -1531
rect 793 -1532 794 -1531
rect 814 -1532 815 -1531
rect 891 -1532 892 -1531
rect 996 -1532 997 -1531
rect 1017 -1532 1018 -1531
rect 1675 -1532 1676 -1531
rect 51 -1534 52 -1533
rect 793 -1534 794 -1533
rect 800 -1534 801 -1533
rect 842 -1534 843 -1533
rect 898 -1534 899 -1533
rect 947 -1534 948 -1533
rect 982 -1534 983 -1533
rect 1157 -1534 1158 -1533
rect 1171 -1534 1172 -1533
rect 1234 -1534 1235 -1533
rect 1258 -1534 1259 -1533
rect 1423 -1534 1424 -1533
rect 1521 -1534 1522 -1533
rect 1542 -1534 1543 -1533
rect 1626 -1534 1627 -1533
rect 1675 -1534 1676 -1533
rect 205 -1536 206 -1535
rect 331 -1536 332 -1535
rect 338 -1536 339 -1535
rect 373 -1536 374 -1535
rect 464 -1536 465 -1535
rect 632 -1536 633 -1535
rect 737 -1536 738 -1535
rect 968 -1536 969 -1535
rect 996 -1536 997 -1535
rect 1059 -1536 1060 -1535
rect 1062 -1536 1063 -1535
rect 1157 -1536 1158 -1535
rect 1199 -1536 1200 -1535
rect 1507 -1536 1508 -1535
rect 1521 -1536 1522 -1535
rect 1661 -1536 1662 -1535
rect 191 -1538 192 -1537
rect 1199 -1538 1200 -1537
rect 1206 -1538 1207 -1537
rect 1360 -1538 1361 -1537
rect 1661 -1538 1662 -1537
rect 1710 -1538 1711 -1537
rect 205 -1540 206 -1539
rect 912 -1540 913 -1539
rect 926 -1540 927 -1539
rect 1290 -1540 1291 -1539
rect 219 -1542 220 -1541
rect 247 -1542 248 -1541
rect 303 -1542 304 -1541
rect 464 -1542 465 -1541
rect 502 -1542 503 -1541
rect 688 -1542 689 -1541
rect 758 -1542 759 -1541
rect 912 -1542 913 -1541
rect 933 -1542 934 -1541
rect 1626 -1542 1627 -1541
rect 184 -1544 185 -1543
rect 247 -1544 248 -1543
rect 324 -1544 325 -1543
rect 695 -1544 696 -1543
rect 758 -1544 759 -1543
rect 1185 -1544 1186 -1543
rect 1227 -1544 1228 -1543
rect 1360 -1544 1361 -1543
rect 135 -1546 136 -1545
rect 184 -1546 185 -1545
rect 233 -1546 234 -1545
rect 303 -1546 304 -1545
rect 338 -1546 339 -1545
rect 383 -1546 384 -1545
rect 506 -1546 507 -1545
rect 716 -1546 717 -1545
rect 842 -1546 843 -1545
rect 1066 -1546 1067 -1545
rect 1129 -1546 1130 -1545
rect 1213 -1546 1214 -1545
rect 1227 -1546 1228 -1545
rect 1724 -1546 1725 -1545
rect 37 -1548 38 -1547
rect 135 -1548 136 -1547
rect 233 -1548 234 -1547
rect 387 -1548 388 -1547
rect 457 -1548 458 -1547
rect 506 -1548 507 -1547
rect 520 -1548 521 -1547
rect 1146 -1548 1147 -1547
rect 1185 -1548 1186 -1547
rect 1241 -1548 1242 -1547
rect 1290 -1548 1291 -1547
rect 1297 -1548 1298 -1547
rect 86 -1550 87 -1549
rect 387 -1550 388 -1549
rect 457 -1550 458 -1549
rect 485 -1550 486 -1549
rect 527 -1550 528 -1549
rect 534 -1550 535 -1549
rect 569 -1550 570 -1549
rect 597 -1550 598 -1549
rect 625 -1550 626 -1549
rect 740 -1550 741 -1549
rect 933 -1550 934 -1549
rect 936 -1550 937 -1549
rect 947 -1550 948 -1549
rect 1031 -1550 1032 -1549
rect 1213 -1550 1214 -1549
rect 1353 -1550 1354 -1549
rect 65 -1552 66 -1551
rect 569 -1552 570 -1551
rect 590 -1552 591 -1551
rect 807 -1552 808 -1551
rect 1031 -1552 1032 -1551
rect 1115 -1552 1116 -1551
rect 1234 -1552 1235 -1551
rect 1255 -1552 1256 -1551
rect 1297 -1552 1298 -1551
rect 1395 -1552 1396 -1551
rect 65 -1554 66 -1553
rect 940 -1554 941 -1553
rect 1241 -1554 1242 -1553
rect 1318 -1554 1319 -1553
rect 1353 -1554 1354 -1553
rect 1437 -1554 1438 -1553
rect 86 -1556 87 -1555
rect 835 -1556 836 -1555
rect 873 -1556 874 -1555
rect 1255 -1556 1256 -1555
rect 1318 -1556 1319 -1555
rect 1374 -1556 1375 -1555
rect 1437 -1556 1438 -1555
rect 1528 -1556 1529 -1555
rect 128 -1558 129 -1557
rect 520 -1558 521 -1557
rect 527 -1558 528 -1557
rect 1717 -1558 1718 -1557
rect 128 -1560 129 -1559
rect 275 -1560 276 -1559
rect 345 -1560 346 -1559
rect 429 -1560 430 -1559
rect 485 -1560 486 -1559
rect 751 -1560 752 -1559
rect 807 -1560 808 -1559
rect 1696 -1560 1697 -1559
rect 170 -1562 171 -1561
rect 835 -1562 836 -1561
rect 1115 -1562 1116 -1561
rect 1528 -1562 1529 -1561
rect 170 -1564 171 -1563
rect 352 -1564 353 -1563
rect 359 -1564 360 -1563
rect 478 -1564 479 -1563
rect 667 -1564 668 -1563
rect 1066 -1564 1067 -1563
rect 1367 -1564 1368 -1563
rect 1374 -1564 1375 -1563
rect 254 -1566 255 -1565
rect 324 -1566 325 -1565
rect 352 -1566 353 -1565
rect 380 -1566 381 -1565
rect 478 -1566 479 -1565
rect 828 -1566 829 -1565
rect 1367 -1566 1368 -1565
rect 1444 -1566 1445 -1565
rect 275 -1568 276 -1567
rect 317 -1568 318 -1567
rect 380 -1568 381 -1567
rect 726 -1568 727 -1567
rect 751 -1568 752 -1567
rect 772 -1568 773 -1567
rect 821 -1568 822 -1567
rect 1395 -1568 1396 -1567
rect 1430 -1568 1431 -1567
rect 1444 -1568 1445 -1567
rect 289 -1570 290 -1569
rect 345 -1570 346 -1569
rect 688 -1570 689 -1569
rect 1010 -1570 1011 -1569
rect 1430 -1570 1431 -1569
rect 1465 -1570 1466 -1569
rect 177 -1572 178 -1571
rect 289 -1572 290 -1571
rect 614 -1572 615 -1571
rect 1465 -1572 1466 -1571
rect 177 -1574 178 -1573
rect 411 -1574 412 -1573
rect 716 -1574 717 -1573
rect 1108 -1574 1109 -1573
rect 723 -1576 724 -1575
rect 1717 -1576 1718 -1575
rect 723 -1578 724 -1577
rect 744 -1578 745 -1577
rect 772 -1578 773 -1577
rect 856 -1578 857 -1577
rect 1010 -1578 1011 -1577
rect 1052 -1578 1053 -1577
rect 1108 -1578 1109 -1577
rect 1192 -1578 1193 -1577
rect 548 -1580 549 -1579
rect 744 -1580 745 -1579
rect 821 -1580 822 -1579
rect 1164 -1580 1165 -1579
rect 1192 -1580 1193 -1579
rect 1269 -1580 1270 -1579
rect 614 -1582 615 -1581
rect 1269 -1582 1270 -1581
rect 726 -1584 727 -1583
rect 954 -1584 955 -1583
rect 1052 -1584 1053 -1583
rect 1080 -1584 1081 -1583
rect 1164 -1584 1165 -1583
rect 1220 -1584 1221 -1583
rect 828 -1586 829 -1585
rect 877 -1586 878 -1585
rect 954 -1586 955 -1585
rect 1101 -1586 1102 -1585
rect 1220 -1586 1221 -1585
rect 1248 -1586 1249 -1585
rect 849 -1588 850 -1587
rect 856 -1588 857 -1587
rect 877 -1588 878 -1587
rect 884 -1588 885 -1587
rect 1080 -1588 1081 -1587
rect 1150 -1588 1151 -1587
rect 1248 -1588 1249 -1587
rect 1304 -1588 1305 -1587
rect 702 -1590 703 -1589
rect 884 -1590 885 -1589
rect 1101 -1590 1102 -1589
rect 1381 -1590 1382 -1589
rect 292 -1592 293 -1591
rect 702 -1592 703 -1591
rect 849 -1592 850 -1591
rect 1003 -1592 1004 -1591
rect 1304 -1592 1305 -1591
rect 1409 -1592 1410 -1591
rect 541 -1594 542 -1593
rect 1409 -1594 1410 -1593
rect 1003 -1596 1004 -1595
rect 1038 -1596 1039 -1595
rect 1381 -1596 1382 -1595
rect 1458 -1596 1459 -1595
rect 1038 -1598 1039 -1597
rect 1178 -1598 1179 -1597
rect 1458 -1598 1459 -1597
rect 1479 -1598 1480 -1597
rect 1178 -1600 1179 -1599
rect 1276 -1600 1277 -1599
rect 1479 -1600 1480 -1599
rect 1647 -1600 1648 -1599
rect 264 -1602 265 -1601
rect 1647 -1602 1648 -1601
rect 1276 -1604 1277 -1603
rect 1388 -1604 1389 -1603
rect 1388 -1606 1389 -1605
rect 1514 -1606 1515 -1605
rect 642 -1608 643 -1607
rect 1514 -1608 1515 -1607
rect 16 -1619 17 -1618
rect 30 -1619 31 -1618
rect 37 -1619 38 -1618
rect 289 -1619 290 -1618
rect 296 -1619 297 -1618
rect 383 -1619 384 -1618
rect 411 -1619 412 -1618
rect 744 -1619 745 -1618
rect 758 -1619 759 -1618
rect 1104 -1619 1105 -1618
rect 1115 -1619 1116 -1618
rect 1318 -1619 1319 -1618
rect 1381 -1619 1382 -1618
rect 1384 -1619 1385 -1618
rect 1479 -1619 1480 -1618
rect 1724 -1619 1725 -1618
rect 1752 -1619 1753 -1618
rect 1766 -1619 1767 -1618
rect 44 -1621 45 -1620
rect 254 -1621 255 -1620
rect 268 -1621 269 -1620
rect 310 -1621 311 -1620
rect 317 -1621 318 -1620
rect 915 -1621 916 -1620
rect 929 -1621 930 -1620
rect 1682 -1621 1683 -1620
rect 1717 -1621 1718 -1620
rect 1780 -1621 1781 -1620
rect 44 -1623 45 -1622
rect 345 -1623 346 -1622
rect 348 -1623 349 -1622
rect 919 -1623 920 -1622
rect 996 -1623 997 -1622
rect 1773 -1623 1774 -1622
rect 58 -1625 59 -1624
rect 1542 -1625 1543 -1624
rect 1626 -1625 1627 -1624
rect 1731 -1625 1732 -1624
rect 65 -1627 66 -1626
rect 495 -1627 496 -1626
rect 513 -1627 514 -1626
rect 726 -1627 727 -1626
rect 730 -1627 731 -1626
rect 758 -1627 759 -1626
rect 761 -1627 762 -1626
rect 1661 -1627 1662 -1626
rect 1668 -1627 1669 -1626
rect 1703 -1627 1704 -1626
rect 79 -1629 80 -1628
rect 264 -1629 265 -1628
rect 268 -1629 269 -1628
rect 320 -1629 321 -1628
rect 324 -1629 325 -1628
rect 366 -1629 367 -1628
rect 369 -1629 370 -1628
rect 415 -1629 416 -1628
rect 432 -1629 433 -1628
rect 457 -1629 458 -1628
rect 478 -1629 479 -1628
rect 614 -1629 615 -1628
rect 667 -1629 668 -1628
rect 814 -1629 815 -1628
rect 828 -1629 829 -1628
rect 894 -1629 895 -1628
rect 919 -1629 920 -1628
rect 922 -1629 923 -1628
rect 975 -1629 976 -1628
rect 1661 -1629 1662 -1628
rect 23 -1631 24 -1630
rect 366 -1631 367 -1630
rect 387 -1631 388 -1630
rect 457 -1631 458 -1630
rect 513 -1631 514 -1630
rect 607 -1631 608 -1630
rect 667 -1631 668 -1630
rect 695 -1631 696 -1630
rect 712 -1631 713 -1630
rect 1024 -1631 1025 -1630
rect 1048 -1631 1049 -1630
rect 1612 -1631 1613 -1630
rect 1640 -1631 1641 -1630
rect 1738 -1631 1739 -1630
rect 61 -1633 62 -1632
rect 387 -1633 388 -1632
rect 450 -1633 451 -1632
rect 789 -1633 790 -1632
rect 793 -1633 794 -1632
rect 1395 -1633 1396 -1632
rect 1486 -1633 1487 -1632
rect 1668 -1633 1669 -1632
rect 79 -1635 80 -1634
rect 548 -1635 549 -1634
rect 562 -1635 563 -1634
rect 1318 -1635 1319 -1634
rect 1381 -1635 1382 -1634
rect 1402 -1635 1403 -1634
rect 1500 -1635 1501 -1634
rect 1626 -1635 1627 -1634
rect 1640 -1635 1641 -1634
rect 1675 -1635 1676 -1634
rect 121 -1637 122 -1636
rect 544 -1637 545 -1636
rect 548 -1637 549 -1636
rect 555 -1637 556 -1636
rect 576 -1637 577 -1636
rect 926 -1637 927 -1636
rect 975 -1637 976 -1636
rect 1458 -1637 1459 -1636
rect 1514 -1637 1515 -1636
rect 1682 -1637 1683 -1636
rect 121 -1639 122 -1638
rect 716 -1639 717 -1638
rect 726 -1639 727 -1638
rect 898 -1639 899 -1638
rect 996 -1639 997 -1638
rect 1038 -1639 1039 -1638
rect 1059 -1639 1060 -1638
rect 1444 -1639 1445 -1638
rect 1521 -1639 1522 -1638
rect 1717 -1639 1718 -1638
rect 135 -1641 136 -1640
rect 618 -1641 619 -1640
rect 674 -1641 675 -1640
rect 740 -1641 741 -1640
rect 803 -1641 804 -1640
rect 814 -1641 815 -1640
rect 863 -1641 864 -1640
rect 1059 -1641 1060 -1640
rect 1115 -1641 1116 -1640
rect 1458 -1641 1459 -1640
rect 1591 -1641 1592 -1640
rect 1675 -1641 1676 -1640
rect 135 -1643 136 -1642
rect 681 -1643 682 -1642
rect 702 -1643 703 -1642
rect 793 -1643 794 -1642
rect 807 -1643 808 -1642
rect 1024 -1643 1025 -1642
rect 1118 -1643 1119 -1642
rect 1234 -1643 1235 -1642
rect 1241 -1643 1242 -1642
rect 1486 -1643 1487 -1642
rect 1598 -1643 1599 -1642
rect 1703 -1643 1704 -1642
rect 156 -1645 157 -1644
rect 415 -1645 416 -1644
rect 450 -1645 451 -1644
rect 747 -1645 748 -1644
rect 807 -1645 808 -1644
rect 898 -1645 899 -1644
rect 992 -1645 993 -1644
rect 1591 -1645 1592 -1644
rect 1647 -1645 1648 -1644
rect 1752 -1645 1753 -1644
rect 156 -1647 157 -1646
rect 982 -1647 983 -1646
rect 1052 -1647 1053 -1646
rect 1241 -1647 1242 -1646
rect 1251 -1647 1252 -1646
rect 1689 -1647 1690 -1646
rect 170 -1649 171 -1648
rect 324 -1649 325 -1648
rect 338 -1649 339 -1648
rect 716 -1649 717 -1648
rect 733 -1649 734 -1648
rect 968 -1649 969 -1648
rect 982 -1649 983 -1648
rect 1017 -1649 1018 -1648
rect 1101 -1649 1102 -1648
rect 1647 -1649 1648 -1648
rect 1654 -1649 1655 -1648
rect 1759 -1649 1760 -1648
rect 170 -1651 171 -1650
rect 331 -1651 332 -1650
rect 338 -1651 339 -1650
rect 646 -1651 647 -1650
rect 709 -1651 710 -1650
rect 1038 -1651 1039 -1650
rect 1101 -1651 1102 -1650
rect 1171 -1651 1172 -1650
rect 1213 -1651 1214 -1650
rect 1500 -1651 1501 -1650
rect 1689 -1651 1690 -1650
rect 1710 -1651 1711 -1650
rect 191 -1653 192 -1652
rect 271 -1653 272 -1652
rect 289 -1653 290 -1652
rect 849 -1653 850 -1652
rect 863 -1653 864 -1652
rect 884 -1653 885 -1652
rect 887 -1653 888 -1652
rect 1430 -1653 1431 -1652
rect 1437 -1653 1438 -1652
rect 1521 -1653 1522 -1652
rect 1619 -1653 1620 -1652
rect 1710 -1653 1711 -1652
rect 191 -1655 192 -1654
rect 870 -1655 871 -1654
rect 968 -1655 969 -1654
rect 989 -1655 990 -1654
rect 1010 -1655 1011 -1654
rect 1052 -1655 1053 -1654
rect 1153 -1655 1154 -1654
rect 1332 -1655 1333 -1654
rect 1367 -1655 1368 -1654
rect 1430 -1655 1431 -1654
rect 1465 -1655 1466 -1654
rect 1598 -1655 1599 -1654
rect 194 -1657 195 -1656
rect 1556 -1657 1557 -1656
rect 205 -1659 206 -1658
rect 1234 -1659 1235 -1658
rect 1255 -1659 1256 -1658
rect 1472 -1659 1473 -1658
rect 1493 -1659 1494 -1658
rect 1556 -1659 1557 -1658
rect 51 -1661 52 -1660
rect 205 -1661 206 -1660
rect 208 -1661 209 -1660
rect 1696 -1661 1697 -1660
rect 51 -1663 52 -1662
rect 408 -1663 409 -1662
rect 422 -1663 423 -1662
rect 709 -1663 710 -1662
rect 737 -1663 738 -1662
rect 1605 -1663 1606 -1662
rect 177 -1665 178 -1664
rect 1255 -1665 1256 -1664
rect 1262 -1665 1263 -1664
rect 1444 -1665 1445 -1664
rect 1507 -1665 1508 -1664
rect 1619 -1665 1620 -1664
rect 212 -1667 213 -1666
rect 310 -1667 311 -1666
rect 331 -1667 332 -1666
rect 978 -1667 979 -1666
rect 1066 -1667 1067 -1666
rect 1472 -1667 1473 -1666
rect 1563 -1667 1564 -1666
rect 1696 -1667 1697 -1666
rect 86 -1669 87 -1668
rect 212 -1669 213 -1668
rect 226 -1669 227 -1668
rect 576 -1669 577 -1668
rect 597 -1669 598 -1668
rect 600 -1669 601 -1668
rect 604 -1669 605 -1668
rect 1122 -1669 1123 -1668
rect 1206 -1669 1207 -1668
rect 1332 -1669 1333 -1668
rect 1367 -1669 1368 -1668
rect 1549 -1669 1550 -1668
rect 1563 -1669 1564 -1668
rect 1706 -1669 1707 -1668
rect 86 -1671 87 -1670
rect 142 -1671 143 -1670
rect 184 -1671 185 -1670
rect 226 -1671 227 -1670
rect 233 -1671 234 -1670
rect 1017 -1671 1018 -1670
rect 1066 -1671 1067 -1670
rect 1437 -1671 1438 -1670
rect 1535 -1671 1536 -1670
rect 1549 -1671 1550 -1670
rect 1584 -1671 1585 -1670
rect 1605 -1671 1606 -1670
rect 142 -1673 143 -1672
rect 163 -1673 164 -1672
rect 184 -1673 185 -1672
rect 198 -1673 199 -1672
rect 233 -1673 234 -1672
rect 261 -1673 262 -1672
rect 278 -1673 279 -1672
rect 1010 -1673 1011 -1672
rect 1073 -1673 1074 -1672
rect 1122 -1673 1123 -1672
rect 1157 -1673 1158 -1672
rect 1206 -1673 1207 -1672
rect 1269 -1673 1270 -1672
rect 1542 -1673 1543 -1672
rect 107 -1675 108 -1674
rect 163 -1675 164 -1674
rect 240 -1675 241 -1674
rect 422 -1675 423 -1674
rect 436 -1675 437 -1674
rect 989 -1675 990 -1674
rect 1073 -1675 1074 -1674
rect 1227 -1675 1228 -1674
rect 1276 -1675 1277 -1674
rect 1479 -1675 1480 -1674
rect 100 -1677 101 -1676
rect 107 -1677 108 -1676
rect 149 -1677 150 -1676
rect 198 -1677 199 -1676
rect 240 -1677 241 -1676
rect 282 -1677 283 -1676
rect 296 -1677 297 -1676
rect 429 -1677 430 -1676
rect 436 -1677 437 -1676
rect 660 -1677 661 -1676
rect 772 -1677 773 -1676
rect 849 -1677 850 -1676
rect 870 -1677 871 -1676
rect 877 -1677 878 -1676
rect 905 -1677 906 -1676
rect 1262 -1677 1263 -1676
rect 1304 -1677 1305 -1676
rect 1395 -1677 1396 -1676
rect 1416 -1677 1417 -1676
rect 1493 -1677 1494 -1676
rect 100 -1679 101 -1678
rect 429 -1679 430 -1678
rect 478 -1679 479 -1678
rect 681 -1679 682 -1678
rect 751 -1679 752 -1678
rect 772 -1679 773 -1678
rect 782 -1679 783 -1678
rect 1584 -1679 1585 -1678
rect 149 -1681 150 -1680
rect 677 -1681 678 -1680
rect 751 -1681 752 -1680
rect 842 -1681 843 -1680
rect 877 -1681 878 -1680
rect 891 -1681 892 -1680
rect 905 -1681 906 -1680
rect 954 -1681 955 -1680
rect 1020 -1681 1021 -1680
rect 1276 -1681 1277 -1680
rect 1339 -1681 1340 -1680
rect 1416 -1681 1417 -1680
rect 1423 -1681 1424 -1680
rect 1514 -1681 1515 -1680
rect 282 -1683 283 -1682
rect 464 -1683 465 -1682
rect 492 -1683 493 -1682
rect 1654 -1683 1655 -1682
rect 359 -1685 360 -1684
rect 464 -1685 465 -1684
rect 471 -1685 472 -1684
rect 492 -1685 493 -1684
rect 499 -1685 500 -1684
rect 695 -1685 696 -1684
rect 796 -1685 797 -1684
rect 1213 -1685 1214 -1684
rect 1339 -1685 1340 -1684
rect 1346 -1685 1347 -1684
rect 1353 -1685 1354 -1684
rect 1423 -1685 1424 -1684
rect 352 -1687 353 -1686
rect 471 -1687 472 -1686
rect 499 -1687 500 -1686
rect 520 -1687 521 -1686
rect 527 -1687 528 -1686
rect 1633 -1687 1634 -1686
rect 219 -1689 220 -1688
rect 352 -1689 353 -1688
rect 359 -1689 360 -1688
rect 1045 -1689 1046 -1688
rect 1118 -1689 1119 -1688
rect 1507 -1689 1508 -1688
rect 1570 -1689 1571 -1688
rect 1633 -1689 1634 -1688
rect 219 -1691 220 -1690
rect 275 -1691 276 -1690
rect 380 -1691 381 -1690
rect 527 -1691 528 -1690
rect 534 -1691 535 -1690
rect 555 -1691 556 -1690
rect 562 -1691 563 -1690
rect 740 -1691 741 -1690
rect 884 -1691 885 -1690
rect 954 -1691 955 -1690
rect 1150 -1691 1151 -1690
rect 1353 -1691 1354 -1690
rect 1374 -1691 1375 -1690
rect 1465 -1691 1466 -1690
rect 1528 -1691 1529 -1690
rect 1570 -1691 1571 -1690
rect 173 -1693 174 -1692
rect 275 -1693 276 -1692
rect 380 -1693 381 -1692
rect 481 -1693 482 -1692
rect 520 -1693 521 -1692
rect 723 -1693 724 -1692
rect 912 -1693 913 -1692
rect 1157 -1693 1158 -1692
rect 1164 -1693 1165 -1692
rect 1227 -1693 1228 -1692
rect 1283 -1693 1284 -1692
rect 1346 -1693 1347 -1692
rect 1374 -1693 1375 -1692
rect 1409 -1693 1410 -1692
rect 177 -1695 178 -1694
rect 1528 -1695 1529 -1694
rect 443 -1697 444 -1696
rect 842 -1697 843 -1696
rect 873 -1697 874 -1696
rect 1409 -1697 1410 -1696
rect 443 -1699 444 -1698
rect 530 -1699 531 -1698
rect 534 -1699 535 -1698
rect 565 -1699 566 -1698
rect 569 -1699 570 -1698
rect 660 -1699 661 -1698
rect 723 -1699 724 -1698
rect 856 -1699 857 -1698
rect 940 -1699 941 -1698
rect 1045 -1699 1046 -1698
rect 1087 -1699 1088 -1698
rect 1150 -1699 1151 -1698
rect 1178 -1699 1179 -1698
rect 1304 -1699 1305 -1698
rect 1388 -1699 1389 -1698
rect 1535 -1699 1536 -1698
rect 530 -1701 531 -1700
rect 835 -1701 836 -1700
rect 929 -1701 930 -1700
rect 1087 -1701 1088 -1700
rect 1108 -1701 1109 -1700
rect 1164 -1701 1165 -1700
rect 1185 -1701 1186 -1700
rect 1269 -1701 1270 -1700
rect 1297 -1701 1298 -1700
rect 1388 -1701 1389 -1700
rect 128 -1703 129 -1702
rect 835 -1703 836 -1702
rect 940 -1703 941 -1702
rect 947 -1703 948 -1702
rect 1094 -1703 1095 -1702
rect 1185 -1703 1186 -1702
rect 1199 -1703 1200 -1702
rect 1283 -1703 1284 -1702
rect 1290 -1703 1291 -1702
rect 1297 -1703 1298 -1702
rect 93 -1705 94 -1704
rect 128 -1705 129 -1704
rect 541 -1705 542 -1704
rect 1577 -1705 1578 -1704
rect 93 -1707 94 -1706
rect 730 -1707 731 -1706
rect 765 -1707 766 -1706
rect 856 -1707 857 -1706
rect 1108 -1707 1109 -1706
rect 1143 -1707 1144 -1706
rect 1192 -1707 1193 -1706
rect 1290 -1707 1291 -1706
rect 1451 -1707 1452 -1706
rect 1577 -1707 1578 -1706
rect 96 -1709 97 -1708
rect 947 -1709 948 -1708
rect 1129 -1709 1130 -1708
rect 1143 -1709 1144 -1708
rect 1360 -1709 1361 -1708
rect 1451 -1709 1452 -1708
rect 159 -1711 160 -1710
rect 1129 -1711 1130 -1710
rect 1136 -1711 1137 -1710
rect 1199 -1711 1200 -1710
rect 1325 -1711 1326 -1710
rect 1360 -1711 1361 -1710
rect 247 -1713 248 -1712
rect 1136 -1713 1137 -1712
rect 1311 -1713 1312 -1712
rect 1325 -1713 1326 -1712
rect 247 -1715 248 -1714
rect 257 -1715 258 -1714
rect 506 -1715 507 -1714
rect 765 -1715 766 -1714
rect 821 -1715 822 -1714
rect 1192 -1715 1193 -1714
rect 1248 -1715 1249 -1714
rect 1311 -1715 1312 -1714
rect 394 -1717 395 -1716
rect 506 -1717 507 -1716
rect 544 -1717 545 -1716
rect 618 -1717 619 -1716
rect 621 -1717 622 -1716
rect 1171 -1717 1172 -1716
rect 394 -1719 395 -1718
rect 401 -1719 402 -1718
rect 569 -1719 570 -1718
rect 719 -1719 720 -1718
rect 800 -1719 801 -1718
rect 821 -1719 822 -1718
rect 828 -1719 829 -1718
rect 1094 -1719 1095 -1718
rect 401 -1721 402 -1720
rect 541 -1721 542 -1720
rect 583 -1721 584 -1720
rect 604 -1721 605 -1720
rect 611 -1721 612 -1720
rect 1612 -1721 1613 -1720
rect 114 -1723 115 -1722
rect 611 -1723 612 -1722
rect 646 -1723 647 -1722
rect 653 -1723 654 -1722
rect 670 -1723 671 -1722
rect 1178 -1723 1179 -1722
rect 114 -1725 115 -1724
rect 590 -1725 591 -1724
rect 597 -1725 598 -1724
rect 625 -1725 626 -1724
rect 653 -1725 654 -1724
rect 786 -1725 787 -1724
rect 800 -1725 801 -1724
rect 1080 -1725 1081 -1724
rect 303 -1727 304 -1726
rect 583 -1727 584 -1726
rect 590 -1727 591 -1726
rect 688 -1727 689 -1726
rect 1031 -1727 1032 -1726
rect 1080 -1727 1081 -1726
rect 1384 -1727 1385 -1726
rect 1402 -1727 1403 -1726
rect 303 -1729 304 -1728
rect 1748 -1729 1749 -1728
rect 688 -1731 689 -1730
rect 779 -1731 780 -1730
rect 926 -1731 927 -1730
rect 1031 -1731 1032 -1730
rect 485 -1733 486 -1732
rect 779 -1733 780 -1732
rect 345 -1735 346 -1734
rect 485 -1735 486 -1734
rect 30 -1746 31 -1745
rect 128 -1746 129 -1745
rect 159 -1746 160 -1745
rect 530 -1746 531 -1745
rect 541 -1746 542 -1745
rect 765 -1746 766 -1745
rect 810 -1746 811 -1745
rect 877 -1746 878 -1745
rect 884 -1746 885 -1745
rect 940 -1746 941 -1745
rect 978 -1746 979 -1745
rect 1598 -1746 1599 -1745
rect 1682 -1746 1683 -1745
rect 1794 -1746 1795 -1745
rect 58 -1748 59 -1747
rect 499 -1748 500 -1747
rect 502 -1748 503 -1747
rect 842 -1748 843 -1747
rect 866 -1748 867 -1747
rect 1808 -1748 1809 -1747
rect 61 -1750 62 -1749
rect 352 -1750 353 -1749
rect 401 -1750 402 -1749
rect 940 -1750 941 -1749
rect 989 -1750 990 -1749
rect 1647 -1750 1648 -1749
rect 1748 -1750 1749 -1749
rect 1766 -1750 1767 -1749
rect 1780 -1750 1781 -1749
rect 1815 -1750 1816 -1749
rect 65 -1752 66 -1751
rect 254 -1752 255 -1751
rect 275 -1752 276 -1751
rect 415 -1752 416 -1751
rect 450 -1752 451 -1751
rect 1248 -1752 1249 -1751
rect 1367 -1752 1368 -1751
rect 1682 -1752 1683 -1751
rect 1752 -1752 1753 -1751
rect 1766 -1752 1767 -1751
rect 65 -1754 66 -1753
rect 170 -1754 171 -1753
rect 177 -1754 178 -1753
rect 1626 -1754 1627 -1753
rect 1738 -1754 1739 -1753
rect 1752 -1754 1753 -1753
rect 107 -1756 108 -1755
rect 128 -1756 129 -1755
rect 159 -1756 160 -1755
rect 296 -1756 297 -1755
rect 324 -1756 325 -1755
rect 481 -1756 482 -1755
rect 618 -1756 619 -1755
rect 730 -1756 731 -1755
rect 740 -1756 741 -1755
rect 1059 -1756 1060 -1755
rect 1069 -1756 1070 -1755
rect 1535 -1756 1536 -1755
rect 1612 -1756 1613 -1755
rect 1647 -1756 1648 -1755
rect 1710 -1756 1711 -1755
rect 1738 -1756 1739 -1755
rect 107 -1758 108 -1757
rect 1192 -1758 1193 -1757
rect 1199 -1758 1200 -1757
rect 1248 -1758 1249 -1757
rect 1332 -1758 1333 -1757
rect 1367 -1758 1368 -1757
rect 1374 -1758 1375 -1757
rect 1535 -1758 1536 -1757
rect 1605 -1758 1606 -1757
rect 1612 -1758 1613 -1757
rect 1626 -1758 1627 -1757
rect 1640 -1758 1641 -1757
rect 1696 -1758 1697 -1757
rect 1710 -1758 1711 -1757
rect 110 -1760 111 -1759
rect 254 -1760 255 -1759
rect 275 -1760 276 -1759
rect 800 -1760 801 -1759
rect 814 -1760 815 -1759
rect 842 -1760 843 -1759
rect 870 -1760 871 -1759
rect 1059 -1760 1060 -1759
rect 1080 -1760 1081 -1759
rect 1115 -1760 1116 -1759
rect 1160 -1760 1161 -1759
rect 1213 -1760 1214 -1759
rect 1374 -1760 1375 -1759
rect 1493 -1760 1494 -1759
rect 1528 -1760 1529 -1759
rect 1640 -1760 1641 -1759
rect 114 -1762 115 -1761
rect 618 -1762 619 -1761
rect 667 -1762 668 -1761
rect 765 -1762 766 -1761
rect 793 -1762 794 -1761
rect 877 -1762 878 -1761
rect 887 -1762 888 -1761
rect 1318 -1762 1319 -1761
rect 1444 -1762 1445 -1761
rect 1493 -1762 1494 -1761
rect 1528 -1762 1529 -1761
rect 1619 -1762 1620 -1761
rect 1633 -1762 1634 -1761
rect 1696 -1762 1697 -1761
rect 114 -1764 115 -1763
rect 366 -1764 367 -1763
rect 408 -1764 409 -1763
rect 485 -1764 486 -1763
rect 625 -1764 626 -1763
rect 667 -1764 668 -1763
rect 677 -1764 678 -1763
rect 772 -1764 773 -1763
rect 800 -1764 801 -1763
rect 1045 -1764 1046 -1763
rect 1073 -1764 1074 -1763
rect 1080 -1764 1081 -1763
rect 1108 -1764 1109 -1763
rect 1199 -1764 1200 -1763
rect 1276 -1764 1277 -1763
rect 1318 -1764 1319 -1763
rect 1430 -1764 1431 -1763
rect 1444 -1764 1445 -1763
rect 1563 -1764 1564 -1763
rect 1605 -1764 1606 -1763
rect 149 -1766 150 -1765
rect 1073 -1766 1074 -1765
rect 1111 -1766 1112 -1765
rect 1668 -1766 1669 -1765
rect 149 -1768 150 -1767
rect 184 -1768 185 -1767
rect 191 -1768 192 -1767
rect 436 -1768 437 -1767
rect 478 -1768 479 -1767
rect 1780 -1768 1781 -1767
rect 170 -1770 171 -1769
rect 810 -1770 811 -1769
rect 821 -1770 822 -1769
rect 870 -1770 871 -1769
rect 891 -1770 892 -1769
rect 1479 -1770 1480 -1769
rect 1549 -1770 1550 -1769
rect 1668 -1770 1669 -1769
rect 180 -1772 181 -1771
rect 422 -1772 423 -1771
rect 436 -1772 437 -1771
rect 443 -1772 444 -1771
rect 625 -1772 626 -1771
rect 726 -1772 727 -1771
rect 733 -1772 734 -1771
rect 1479 -1772 1480 -1771
rect 1584 -1772 1585 -1771
rect 1619 -1772 1620 -1771
rect 180 -1774 181 -1773
rect 1661 -1774 1662 -1773
rect 184 -1776 185 -1775
rect 548 -1776 549 -1775
rect 688 -1776 689 -1775
rect 982 -1776 983 -1775
rect 989 -1776 990 -1775
rect 1031 -1776 1032 -1775
rect 1041 -1776 1042 -1775
rect 1269 -1776 1270 -1775
rect 1279 -1776 1280 -1775
rect 1549 -1776 1550 -1775
rect 1570 -1776 1571 -1775
rect 1661 -1776 1662 -1775
rect 191 -1778 192 -1777
rect 1654 -1778 1655 -1777
rect 208 -1780 209 -1779
rect 541 -1780 542 -1779
rect 548 -1780 549 -1779
rect 1010 -1780 1011 -1779
rect 1017 -1780 1018 -1779
rect 1213 -1780 1214 -1779
rect 1234 -1780 1235 -1779
rect 1430 -1780 1431 -1779
rect 1521 -1780 1522 -1779
rect 1584 -1780 1585 -1779
rect 1591 -1780 1592 -1779
rect 1654 -1780 1655 -1779
rect 233 -1782 234 -1781
rect 341 -1782 342 -1781
rect 348 -1782 349 -1781
rect 835 -1782 836 -1781
rect 849 -1782 850 -1781
rect 891 -1782 892 -1781
rect 915 -1782 916 -1781
rect 1388 -1782 1389 -1781
rect 1507 -1782 1508 -1781
rect 1591 -1782 1592 -1781
rect 233 -1784 234 -1783
rect 432 -1784 433 -1783
rect 576 -1784 577 -1783
rect 688 -1784 689 -1783
rect 695 -1784 696 -1783
rect 786 -1784 787 -1783
rect 821 -1784 822 -1783
rect 1283 -1784 1284 -1783
rect 1381 -1784 1382 -1783
rect 1521 -1784 1522 -1783
rect 1556 -1784 1557 -1783
rect 1570 -1784 1571 -1783
rect 268 -1786 269 -1785
rect 366 -1786 367 -1785
rect 411 -1786 412 -1785
rect 803 -1786 804 -1785
rect 824 -1786 825 -1785
rect 1633 -1786 1634 -1785
rect 268 -1788 269 -1787
rect 569 -1788 570 -1787
rect 576 -1788 577 -1787
rect 894 -1788 895 -1787
rect 919 -1788 920 -1787
rect 1724 -1788 1725 -1787
rect 282 -1790 283 -1789
rect 296 -1790 297 -1789
rect 317 -1790 318 -1789
rect 478 -1790 479 -1789
rect 632 -1790 633 -1789
rect 695 -1790 696 -1789
rect 702 -1790 703 -1789
rect 1171 -1790 1172 -1789
rect 1220 -1790 1221 -1789
rect 1234 -1790 1235 -1789
rect 1269 -1790 1270 -1789
rect 1311 -1790 1312 -1789
rect 1465 -1790 1466 -1789
rect 1507 -1790 1508 -1789
rect 1703 -1790 1704 -1789
rect 1724 -1790 1725 -1789
rect 156 -1792 157 -1791
rect 1465 -1792 1466 -1791
rect 1675 -1792 1676 -1791
rect 1703 -1792 1704 -1791
rect 156 -1794 157 -1793
rect 632 -1794 633 -1793
rect 639 -1794 640 -1793
rect 702 -1794 703 -1793
rect 709 -1794 710 -1793
rect 793 -1794 794 -1793
rect 828 -1794 829 -1793
rect 1157 -1794 1158 -1793
rect 1171 -1794 1172 -1793
rect 1804 -1794 1805 -1793
rect 198 -1796 199 -1795
rect 317 -1796 318 -1795
rect 324 -1796 325 -1795
rect 394 -1796 395 -1795
rect 415 -1796 416 -1795
rect 922 -1796 923 -1795
rect 926 -1796 927 -1795
rect 1136 -1796 1137 -1795
rect 1157 -1796 1158 -1795
rect 1416 -1796 1417 -1795
rect 1675 -1796 1676 -1795
rect 1689 -1796 1690 -1795
rect 198 -1798 199 -1797
rect 513 -1798 514 -1797
rect 639 -1798 640 -1797
rect 646 -1798 647 -1797
rect 709 -1798 710 -1797
rect 1066 -1798 1067 -1797
rect 1115 -1798 1116 -1797
rect 1164 -1798 1165 -1797
rect 1178 -1798 1179 -1797
rect 1220 -1798 1221 -1797
rect 1276 -1798 1277 -1797
rect 1689 -1798 1690 -1797
rect 247 -1800 248 -1799
rect 282 -1800 283 -1799
rect 289 -1800 290 -1799
rect 1136 -1800 1137 -1799
rect 1283 -1800 1284 -1799
rect 1290 -1800 1291 -1799
rect 1416 -1800 1417 -1799
rect 1745 -1800 1746 -1799
rect 121 -1802 122 -1801
rect 289 -1802 290 -1801
rect 310 -1802 311 -1801
rect 394 -1802 395 -1801
rect 422 -1802 423 -1801
rect 674 -1802 675 -1801
rect 716 -1802 717 -1801
rect 1010 -1802 1011 -1801
rect 1017 -1802 1018 -1801
rect 1486 -1802 1487 -1801
rect 1731 -1802 1732 -1801
rect 1745 -1802 1746 -1801
rect 93 -1804 94 -1803
rect 716 -1804 717 -1803
rect 737 -1804 738 -1803
rect 1381 -1804 1382 -1803
rect 1717 -1804 1718 -1803
rect 1731 -1804 1732 -1803
rect 93 -1806 94 -1805
rect 257 -1806 258 -1805
rect 303 -1806 304 -1805
rect 737 -1806 738 -1805
rect 744 -1806 745 -1805
rect 912 -1806 913 -1805
rect 919 -1806 920 -1805
rect 1776 -1806 1777 -1805
rect 79 -1808 80 -1807
rect 303 -1808 304 -1807
rect 331 -1808 332 -1807
rect 352 -1808 353 -1807
rect 359 -1808 360 -1807
rect 485 -1808 486 -1807
rect 674 -1808 675 -1807
rect 1108 -1808 1109 -1807
rect 1153 -1808 1154 -1807
rect 1486 -1808 1487 -1807
rect 79 -1810 80 -1809
rect 380 -1810 381 -1809
rect 446 -1810 447 -1809
rect 1556 -1810 1557 -1809
rect 121 -1812 122 -1811
rect 506 -1812 507 -1811
rect 744 -1812 745 -1811
rect 751 -1812 752 -1811
rect 758 -1812 759 -1811
rect 814 -1812 815 -1811
rect 828 -1812 829 -1811
rect 1787 -1812 1788 -1811
rect 135 -1814 136 -1813
rect 758 -1814 759 -1813
rect 772 -1814 773 -1813
rect 1801 -1814 1802 -1813
rect 100 -1816 101 -1815
rect 135 -1816 136 -1815
rect 205 -1816 206 -1815
rect 310 -1816 311 -1815
rect 331 -1816 332 -1815
rect 443 -1816 444 -1815
rect 464 -1816 465 -1815
rect 513 -1816 514 -1815
rect 611 -1816 612 -1815
rect 751 -1816 752 -1815
rect 789 -1816 790 -1815
rect 1717 -1816 1718 -1815
rect 100 -1818 101 -1817
rect 226 -1818 227 -1817
rect 338 -1818 339 -1817
rect 474 -1818 475 -1817
rect 506 -1818 507 -1817
rect 555 -1818 556 -1817
rect 597 -1818 598 -1817
rect 611 -1818 612 -1817
rect 849 -1818 850 -1817
rect 1087 -1818 1088 -1817
rect 1101 -1818 1102 -1817
rect 1178 -1818 1179 -1817
rect 1290 -1818 1291 -1817
rect 1773 -1818 1774 -1817
rect 86 -1820 87 -1819
rect 555 -1820 556 -1819
rect 597 -1820 598 -1819
rect 779 -1820 780 -1819
rect 863 -1820 864 -1819
rect 1101 -1820 1102 -1819
rect 1542 -1820 1543 -1819
rect 1773 -1820 1774 -1819
rect 72 -1822 73 -1821
rect 86 -1822 87 -1821
rect 205 -1822 206 -1821
rect 1255 -1822 1256 -1821
rect 1458 -1822 1459 -1821
rect 1542 -1822 1543 -1821
rect 44 -1824 45 -1823
rect 72 -1824 73 -1823
rect 212 -1824 213 -1823
rect 779 -1824 780 -1823
rect 863 -1824 864 -1823
rect 1262 -1824 1263 -1823
rect 1423 -1824 1424 -1823
rect 1458 -1824 1459 -1823
rect 44 -1826 45 -1825
rect 163 -1826 164 -1825
rect 212 -1826 213 -1825
rect 492 -1826 493 -1825
rect 912 -1826 913 -1825
rect 954 -1826 955 -1825
rect 982 -1826 983 -1825
rect 1241 -1826 1242 -1825
rect 1339 -1826 1340 -1825
rect 1423 -1826 1424 -1825
rect 163 -1828 164 -1827
rect 831 -1828 832 -1827
rect 926 -1828 927 -1827
rect 1577 -1828 1578 -1827
rect 219 -1830 220 -1829
rect 226 -1830 227 -1829
rect 338 -1830 339 -1829
rect 467 -1830 468 -1829
rect 471 -1830 472 -1829
rect 569 -1830 570 -1829
rect 831 -1830 832 -1829
rect 1332 -1830 1333 -1829
rect 1402 -1830 1403 -1829
rect 1577 -1830 1578 -1829
rect 219 -1832 220 -1831
rect 691 -1832 692 -1831
rect 929 -1832 930 -1831
rect 1500 -1832 1501 -1831
rect 359 -1834 360 -1833
rect 373 -1834 374 -1833
rect 380 -1834 381 -1833
rect 457 -1834 458 -1833
rect 492 -1834 493 -1833
rect 527 -1834 528 -1833
rect 936 -1834 937 -1833
rect 1150 -1834 1151 -1833
rect 1206 -1834 1207 -1833
rect 1255 -1834 1256 -1833
rect 1395 -1834 1396 -1833
rect 1402 -1834 1403 -1833
rect 37 -1836 38 -1835
rect 527 -1836 528 -1835
rect 947 -1836 948 -1835
rect 1388 -1836 1389 -1835
rect 37 -1838 38 -1837
rect 51 -1838 52 -1837
rect 247 -1838 248 -1837
rect 457 -1838 458 -1837
rect 898 -1838 899 -1837
rect 947 -1838 948 -1837
rect 975 -1838 976 -1837
rect 1150 -1838 1151 -1837
rect 1206 -1838 1207 -1837
rect 1304 -1838 1305 -1837
rect 1346 -1838 1347 -1837
rect 1395 -1838 1396 -1837
rect 51 -1840 52 -1839
rect 142 -1840 143 -1839
rect 373 -1840 374 -1839
rect 562 -1840 563 -1839
rect 898 -1840 899 -1839
rect 929 -1840 930 -1839
rect 933 -1840 934 -1839
rect 1346 -1840 1347 -1839
rect 142 -1842 143 -1841
rect 177 -1842 178 -1841
rect 401 -1842 402 -1841
rect 471 -1842 472 -1841
rect 562 -1842 563 -1841
rect 649 -1842 650 -1841
rect 856 -1842 857 -1841
rect 933 -1842 934 -1841
rect 996 -1842 997 -1841
rect 1192 -1842 1193 -1841
rect 1227 -1842 1228 -1841
rect 1262 -1842 1263 -1841
rect 1297 -1842 1298 -1841
rect 1304 -1842 1305 -1841
rect 429 -1844 430 -1843
rect 464 -1844 465 -1843
rect 656 -1844 657 -1843
rect 1227 -1844 1228 -1843
rect 1251 -1844 1252 -1843
rect 1339 -1844 1340 -1843
rect 681 -1846 682 -1845
rect 856 -1846 857 -1845
rect 961 -1846 962 -1845
rect 996 -1846 997 -1845
rect 1003 -1846 1004 -1845
rect 1031 -1846 1032 -1845
rect 1038 -1846 1039 -1845
rect 1087 -1846 1088 -1845
rect 1143 -1846 1144 -1845
rect 1241 -1846 1242 -1845
rect 1297 -1846 1298 -1845
rect 1514 -1846 1515 -1845
rect 345 -1848 346 -1847
rect 1038 -1848 1039 -1847
rect 1045 -1848 1046 -1847
rect 1563 -1848 1564 -1847
rect 583 -1850 584 -1849
rect 681 -1850 682 -1849
rect 835 -1850 836 -1849
rect 1003 -1850 1004 -1849
rect 1024 -1850 1025 -1849
rect 1164 -1850 1165 -1849
rect 1353 -1850 1354 -1849
rect 1514 -1850 1515 -1849
rect 583 -1852 584 -1851
rect 590 -1852 591 -1851
rect 653 -1852 654 -1851
rect 961 -1852 962 -1851
rect 968 -1852 969 -1851
rect 1024 -1852 1025 -1851
rect 1027 -1852 1028 -1851
rect 1598 -1852 1599 -1851
rect 450 -1854 451 -1853
rect 653 -1854 654 -1853
rect 968 -1854 969 -1853
rect 985 -1854 986 -1853
rect 1048 -1854 1049 -1853
rect 1500 -1854 1501 -1853
rect 590 -1856 591 -1855
rect 660 -1856 661 -1855
rect 1066 -1856 1067 -1855
rect 1129 -1856 1130 -1855
rect 1353 -1856 1354 -1855
rect 1472 -1856 1473 -1855
rect 660 -1858 661 -1857
rect 782 -1858 783 -1857
rect 905 -1858 906 -1857
rect 1129 -1858 1130 -1857
rect 1451 -1858 1452 -1857
rect 1472 -1858 1473 -1857
rect 807 -1860 808 -1859
rect 1451 -1860 1452 -1859
rect 905 -1862 906 -1861
rect 1437 -1862 1438 -1861
rect 1094 -1864 1095 -1863
rect 1143 -1864 1144 -1863
rect 1409 -1864 1410 -1863
rect 1437 -1864 1438 -1863
rect 194 -1866 195 -1865
rect 1409 -1866 1410 -1865
rect 1094 -1868 1095 -1867
rect 1122 -1868 1123 -1867
rect 1122 -1870 1123 -1869
rect 1185 -1870 1186 -1869
rect 1185 -1872 1186 -1871
rect 1360 -1872 1361 -1871
rect 1325 -1874 1326 -1873
rect 1360 -1874 1361 -1873
rect 723 -1876 724 -1875
rect 1325 -1876 1326 -1875
rect 387 -1878 388 -1877
rect 723 -1878 724 -1877
rect 387 -1880 388 -1879
rect 520 -1880 521 -1879
rect 250 -1882 251 -1881
rect 520 -1882 521 -1881
rect 51 -1893 52 -1892
rect 215 -1893 216 -1892
rect 233 -1893 234 -1892
rect 887 -1893 888 -1892
rect 905 -1893 906 -1892
rect 1199 -1893 1200 -1892
rect 1216 -1893 1217 -1892
rect 1227 -1893 1228 -1892
rect 1276 -1893 1277 -1892
rect 1577 -1893 1578 -1892
rect 1654 -1893 1655 -1892
rect 1804 -1893 1805 -1892
rect 51 -1895 52 -1894
rect 268 -1895 269 -1894
rect 303 -1895 304 -1894
rect 474 -1895 475 -1894
rect 478 -1895 479 -1894
rect 905 -1895 906 -1894
rect 919 -1895 920 -1894
rect 982 -1895 983 -1894
rect 1017 -1895 1018 -1894
rect 1164 -1895 1165 -1894
rect 1276 -1895 1277 -1894
rect 1416 -1895 1417 -1894
rect 1773 -1895 1774 -1894
rect 1794 -1895 1795 -1894
rect 68 -1897 69 -1896
rect 548 -1897 549 -1896
rect 572 -1897 573 -1896
rect 1346 -1897 1347 -1896
rect 1381 -1897 1382 -1896
rect 1384 -1897 1385 -1896
rect 1409 -1897 1410 -1896
rect 1776 -1897 1777 -1896
rect 1794 -1897 1795 -1896
rect 1808 -1897 1809 -1896
rect 72 -1899 73 -1898
rect 107 -1899 108 -1898
rect 135 -1899 136 -1898
rect 261 -1899 262 -1898
rect 303 -1899 304 -1898
rect 562 -1899 563 -1898
rect 593 -1899 594 -1898
rect 1451 -1899 1452 -1898
rect 1493 -1899 1494 -1898
rect 1808 -1899 1809 -1898
rect 72 -1901 73 -1900
rect 149 -1901 150 -1900
rect 156 -1901 157 -1900
rect 233 -1901 234 -1900
rect 250 -1901 251 -1900
rect 548 -1901 549 -1900
rect 562 -1901 563 -1900
rect 947 -1901 948 -1900
rect 954 -1901 955 -1900
rect 968 -1901 969 -1900
rect 1024 -1901 1025 -1900
rect 1759 -1901 1760 -1900
rect 79 -1903 80 -1902
rect 338 -1903 339 -1902
rect 345 -1903 346 -1902
rect 828 -1903 829 -1902
rect 831 -1903 832 -1902
rect 1101 -1903 1102 -1902
rect 1111 -1903 1112 -1902
rect 1724 -1903 1725 -1902
rect 79 -1905 80 -1904
rect 611 -1905 612 -1904
rect 646 -1905 647 -1904
rect 779 -1905 780 -1904
rect 796 -1905 797 -1904
rect 842 -1905 843 -1904
rect 849 -1905 850 -1904
rect 1199 -1905 1200 -1904
rect 1279 -1905 1280 -1904
rect 1724 -1905 1725 -1904
rect 86 -1907 87 -1906
rect 107 -1907 108 -1906
rect 135 -1907 136 -1906
rect 401 -1907 402 -1906
rect 436 -1907 437 -1906
rect 999 -1907 1000 -1906
rect 1024 -1907 1025 -1906
rect 1143 -1907 1144 -1906
rect 1153 -1907 1154 -1906
rect 1731 -1907 1732 -1906
rect 86 -1909 87 -1908
rect 310 -1909 311 -1908
rect 324 -1909 325 -1908
rect 467 -1909 468 -1908
rect 499 -1909 500 -1908
rect 866 -1909 867 -1908
rect 922 -1909 923 -1908
rect 985 -1909 986 -1908
rect 1031 -1909 1032 -1908
rect 1101 -1909 1102 -1908
rect 1115 -1909 1116 -1908
rect 1227 -1909 1228 -1908
rect 1314 -1909 1315 -1908
rect 1633 -1909 1634 -1908
rect 1731 -1909 1732 -1908
rect 1752 -1909 1753 -1908
rect 89 -1911 90 -1910
rect 1164 -1911 1165 -1910
rect 1353 -1911 1354 -1910
rect 1493 -1911 1494 -1910
rect 1633 -1911 1634 -1910
rect 1647 -1911 1648 -1910
rect 1752 -1911 1753 -1910
rect 1780 -1911 1781 -1910
rect 100 -1913 101 -1912
rect 446 -1913 447 -1912
rect 464 -1913 465 -1912
rect 877 -1913 878 -1912
rect 926 -1913 927 -1912
rect 996 -1913 997 -1912
rect 1003 -1913 1004 -1912
rect 1115 -1913 1116 -1912
rect 1139 -1913 1140 -1912
rect 1773 -1913 1774 -1912
rect 1780 -1913 1781 -1912
rect 1801 -1913 1802 -1912
rect 100 -1915 101 -1914
rect 1577 -1915 1578 -1914
rect 1801 -1915 1802 -1914
rect 1815 -1915 1816 -1914
rect 110 -1917 111 -1916
rect 436 -1917 437 -1916
rect 509 -1917 510 -1916
rect 1346 -1917 1347 -1916
rect 1381 -1917 1382 -1916
rect 1507 -1917 1508 -1916
rect 142 -1919 143 -1918
rect 1654 -1919 1655 -1918
rect 142 -1921 143 -1920
rect 1556 -1921 1557 -1920
rect 145 -1923 146 -1922
rect 310 -1923 311 -1922
rect 324 -1923 325 -1922
rect 394 -1923 395 -1922
rect 527 -1923 528 -1922
rect 1689 -1923 1690 -1922
rect 149 -1925 150 -1924
rect 208 -1925 209 -1924
rect 212 -1925 213 -1924
rect 443 -1925 444 -1924
rect 527 -1925 528 -1924
rect 674 -1925 675 -1924
rect 723 -1925 724 -1924
rect 947 -1925 948 -1924
rect 957 -1925 958 -1924
rect 1318 -1925 1319 -1924
rect 1409 -1925 1410 -1924
rect 1521 -1925 1522 -1924
rect 1626 -1925 1627 -1924
rect 1689 -1925 1690 -1924
rect 156 -1927 157 -1926
rect 184 -1927 185 -1926
rect 191 -1927 192 -1926
rect 268 -1927 269 -1926
rect 334 -1927 335 -1926
rect 443 -1927 444 -1926
rect 541 -1927 542 -1926
rect 611 -1927 612 -1926
rect 618 -1927 619 -1926
rect 926 -1927 927 -1926
rect 929 -1927 930 -1926
rect 1003 -1927 1004 -1926
rect 1027 -1927 1028 -1926
rect 1647 -1927 1648 -1926
rect 128 -1929 129 -1928
rect 184 -1929 185 -1928
rect 191 -1929 192 -1928
rect 415 -1929 416 -1928
rect 506 -1929 507 -1928
rect 541 -1929 542 -1928
rect 597 -1929 598 -1928
rect 779 -1929 780 -1928
rect 800 -1929 801 -1928
rect 975 -1929 976 -1928
rect 1031 -1929 1032 -1928
rect 1080 -1929 1081 -1928
rect 1143 -1929 1144 -1928
rect 1248 -1929 1249 -1928
rect 1318 -1929 1319 -1928
rect 1360 -1929 1361 -1928
rect 1374 -1929 1375 -1928
rect 1521 -1929 1522 -1928
rect 1626 -1929 1627 -1928
rect 1675 -1929 1676 -1928
rect 152 -1931 153 -1930
rect 415 -1931 416 -1930
rect 457 -1931 458 -1930
rect 597 -1931 598 -1930
rect 618 -1931 619 -1930
rect 639 -1931 640 -1930
rect 653 -1931 654 -1930
rect 1213 -1931 1214 -1930
rect 1248 -1931 1249 -1930
rect 1262 -1931 1263 -1930
rect 1360 -1931 1361 -1930
rect 1444 -1931 1445 -1930
rect 1675 -1931 1676 -1930
rect 1710 -1931 1711 -1930
rect 37 -1933 38 -1932
rect 457 -1933 458 -1932
rect 506 -1933 507 -1932
rect 1759 -1933 1760 -1932
rect 159 -1935 160 -1934
rect 863 -1935 864 -1934
rect 901 -1935 902 -1934
rect 1556 -1935 1557 -1934
rect 1710 -1935 1711 -1934
rect 1745 -1935 1746 -1934
rect 163 -1937 164 -1936
rect 247 -1937 248 -1936
rect 254 -1937 255 -1936
rect 1048 -1937 1049 -1936
rect 1059 -1937 1060 -1936
rect 1353 -1937 1354 -1936
rect 1374 -1937 1375 -1936
rect 1395 -1937 1396 -1936
rect 1423 -1937 1424 -1936
rect 1444 -1937 1445 -1936
rect 163 -1939 164 -1938
rect 341 -1939 342 -1938
rect 345 -1939 346 -1938
rect 429 -1939 430 -1938
rect 632 -1939 633 -1938
rect 646 -1939 647 -1938
rect 653 -1939 654 -1938
rect 1041 -1939 1042 -1938
rect 1045 -1939 1046 -1938
rect 1297 -1939 1298 -1938
rect 1395 -1939 1396 -1938
rect 1500 -1939 1501 -1938
rect 93 -1941 94 -1940
rect 1500 -1941 1501 -1940
rect 93 -1943 94 -1942
rect 177 -1943 178 -1942
rect 198 -1943 199 -1942
rect 429 -1943 430 -1942
rect 632 -1943 633 -1942
rect 702 -1943 703 -1942
rect 793 -1943 794 -1942
rect 800 -1943 801 -1942
rect 807 -1943 808 -1942
rect 961 -1943 962 -1942
rect 968 -1943 969 -1942
rect 1332 -1943 1333 -1942
rect 1423 -1943 1424 -1942
rect 1514 -1943 1515 -1942
rect 103 -1945 104 -1944
rect 1332 -1945 1333 -1944
rect 1437 -1945 1438 -1944
rect 1451 -1945 1452 -1944
rect 1514 -1945 1515 -1944
rect 1535 -1945 1536 -1944
rect 170 -1947 171 -1946
rect 401 -1947 402 -1946
rect 460 -1947 461 -1946
rect 702 -1947 703 -1946
rect 807 -1947 808 -1946
rect 891 -1947 892 -1946
rect 933 -1947 934 -1946
rect 940 -1947 941 -1946
rect 975 -1947 976 -1946
rect 1339 -1947 1340 -1946
rect 1402 -1947 1403 -1946
rect 1437 -1947 1438 -1946
rect 1535 -1947 1536 -1946
rect 1563 -1947 1564 -1946
rect 110 -1949 111 -1948
rect 1402 -1949 1403 -1948
rect 1563 -1949 1564 -1948
rect 1570 -1949 1571 -1948
rect 170 -1951 171 -1950
rect 226 -1951 227 -1950
rect 247 -1951 248 -1950
rect 275 -1951 276 -1950
rect 373 -1951 374 -1950
rect 376 -1951 377 -1950
rect 380 -1951 381 -1950
rect 478 -1951 479 -1950
rect 639 -1951 640 -1950
rect 821 -1951 822 -1950
rect 824 -1951 825 -1950
rect 884 -1951 885 -1950
rect 891 -1951 892 -1950
rect 1458 -1951 1459 -1950
rect 114 -1953 115 -1952
rect 821 -1953 822 -1952
rect 835 -1953 836 -1952
rect 908 -1953 909 -1952
rect 1010 -1953 1011 -1952
rect 1045 -1953 1046 -1952
rect 1080 -1953 1081 -1952
rect 1108 -1953 1109 -1952
rect 1157 -1953 1158 -1952
rect 1185 -1953 1186 -1952
rect 1206 -1953 1207 -1952
rect 1339 -1953 1340 -1952
rect 1430 -1953 1431 -1952
rect 1458 -1953 1459 -1952
rect 114 -1955 115 -1954
rect 282 -1955 283 -1954
rect 373 -1955 374 -1954
rect 492 -1955 493 -1954
rect 667 -1955 668 -1954
rect 674 -1955 675 -1954
rect 719 -1955 720 -1954
rect 1108 -1955 1109 -1954
rect 1122 -1955 1123 -1954
rect 1430 -1955 1431 -1954
rect 131 -1957 132 -1956
rect 226 -1957 227 -1956
rect 254 -1957 255 -1956
rect 534 -1957 535 -1956
rect 667 -1957 668 -1956
rect 758 -1957 759 -1956
rect 786 -1957 787 -1956
rect 940 -1957 941 -1956
rect 989 -1957 990 -1956
rect 1010 -1957 1011 -1956
rect 1020 -1957 1021 -1956
rect 1059 -1957 1060 -1956
rect 1087 -1957 1088 -1956
rect 1122 -1957 1123 -1956
rect 1129 -1957 1130 -1956
rect 1157 -1957 1158 -1956
rect 1206 -1957 1207 -1956
rect 1241 -1957 1242 -1956
rect 1262 -1957 1263 -1956
rect 1486 -1957 1487 -1956
rect 177 -1959 178 -1958
rect 894 -1959 895 -1958
rect 989 -1959 990 -1958
rect 1584 -1959 1585 -1958
rect 180 -1961 181 -1960
rect 793 -1961 794 -1960
rect 814 -1961 815 -1960
rect 842 -1961 843 -1960
rect 877 -1961 878 -1960
rect 884 -1961 885 -1960
rect 1052 -1961 1053 -1960
rect 1185 -1961 1186 -1960
rect 1241 -1961 1242 -1960
rect 1255 -1961 1256 -1960
rect 1297 -1961 1298 -1960
rect 1325 -1961 1326 -1960
rect 1486 -1961 1487 -1960
rect 1619 -1961 1620 -1960
rect 180 -1963 181 -1962
rect 422 -1963 423 -1962
rect 485 -1963 486 -1962
rect 492 -1963 493 -1962
rect 534 -1963 535 -1962
rect 555 -1963 556 -1962
rect 590 -1963 591 -1962
rect 786 -1963 787 -1962
rect 810 -1963 811 -1962
rect 1325 -1963 1326 -1962
rect 1528 -1963 1529 -1962
rect 1584 -1963 1585 -1962
rect 1619 -1963 1620 -1962
rect 1640 -1963 1641 -1962
rect 58 -1965 59 -1964
rect 555 -1965 556 -1964
rect 758 -1965 759 -1964
rect 1066 -1965 1067 -1964
rect 1073 -1965 1074 -1964
rect 1129 -1965 1130 -1964
rect 1220 -1965 1221 -1964
rect 1255 -1965 1256 -1964
rect 1311 -1965 1312 -1964
rect 1570 -1965 1571 -1964
rect 1640 -1965 1641 -1964
rect 1682 -1965 1683 -1964
rect 58 -1967 59 -1966
rect 709 -1967 710 -1966
rect 814 -1967 815 -1966
rect 856 -1967 857 -1966
rect 1052 -1967 1053 -1966
rect 1136 -1967 1137 -1966
rect 1192 -1967 1193 -1966
rect 1220 -1967 1221 -1966
rect 1269 -1967 1270 -1966
rect 1311 -1967 1312 -1966
rect 1384 -1967 1385 -1966
rect 1507 -1967 1508 -1966
rect 1528 -1967 1529 -1966
rect 1549 -1967 1550 -1966
rect 1682 -1967 1683 -1966
rect 1717 -1967 1718 -1966
rect 198 -1969 199 -1968
rect 761 -1969 762 -1968
rect 838 -1969 839 -1968
rect 1388 -1969 1389 -1968
rect 1542 -1969 1543 -1968
rect 1549 -1969 1550 -1968
rect 205 -1971 206 -1970
rect 289 -1971 290 -1970
rect 387 -1971 388 -1970
rect 464 -1971 465 -1970
rect 649 -1971 650 -1970
rect 1717 -1971 1718 -1970
rect 212 -1973 213 -1972
rect 1598 -1973 1599 -1972
rect 219 -1975 220 -1974
rect 1087 -1975 1088 -1974
rect 1178 -1975 1179 -1974
rect 1269 -1975 1270 -1974
rect 1388 -1975 1389 -1974
rect 1472 -1975 1473 -1974
rect 1598 -1975 1599 -1974
rect 1612 -1975 1613 -1974
rect 219 -1977 220 -1976
rect 380 -1977 381 -1976
rect 394 -1977 395 -1976
rect 716 -1977 717 -1976
rect 856 -1977 857 -1976
rect 870 -1977 871 -1976
rect 1017 -1977 1018 -1976
rect 1136 -1977 1137 -1976
rect 1178 -1977 1179 -1976
rect 1367 -1977 1368 -1976
rect 1465 -1977 1466 -1976
rect 1472 -1977 1473 -1976
rect 1612 -1977 1613 -1976
rect 1661 -1977 1662 -1976
rect 264 -1979 265 -1978
rect 289 -1979 290 -1978
rect 422 -1979 423 -1978
rect 730 -1979 731 -1978
rect 870 -1979 871 -1978
rect 936 -1979 937 -1978
rect 1038 -1979 1039 -1978
rect 1542 -1979 1543 -1978
rect 1661 -1979 1662 -1978
rect 1703 -1979 1704 -1978
rect 275 -1981 276 -1980
rect 359 -1981 360 -1980
rect 709 -1981 710 -1980
rect 898 -1981 899 -1980
rect 1038 -1981 1039 -1980
rect 1696 -1981 1697 -1980
rect 1703 -1981 1704 -1980
rect 1738 -1981 1739 -1980
rect 282 -1983 283 -1982
rect 471 -1983 472 -1982
rect 716 -1983 717 -1982
rect 849 -1983 850 -1982
rect 1066 -1983 1067 -1982
rect 1290 -1983 1291 -1982
rect 1293 -1983 1294 -1982
rect 1696 -1983 1697 -1982
rect 1738 -1983 1739 -1982
rect 1766 -1983 1767 -1982
rect 359 -1985 360 -1984
rect 688 -1985 689 -1984
rect 723 -1985 724 -1984
rect 898 -1985 899 -1984
rect 1073 -1985 1074 -1984
rect 1094 -1985 1095 -1984
rect 1192 -1985 1193 -1984
rect 1416 -1985 1417 -1984
rect 1465 -1985 1466 -1984
rect 1605 -1985 1606 -1984
rect 1766 -1985 1767 -1984
rect 1787 -1985 1788 -1984
rect 366 -1987 367 -1986
rect 471 -1987 472 -1986
rect 583 -1987 584 -1986
rect 1094 -1987 1095 -1986
rect 1304 -1987 1305 -1986
rect 1367 -1987 1368 -1986
rect 1591 -1987 1592 -1986
rect 1605 -1987 1606 -1986
rect 317 -1989 318 -1988
rect 366 -1989 367 -1988
rect 583 -1989 584 -1988
rect 625 -1989 626 -1988
rect 628 -1989 629 -1988
rect 1304 -1989 1305 -1988
rect 317 -1991 318 -1990
rect 408 -1991 409 -1990
rect 625 -1991 626 -1990
rect 695 -1991 696 -1990
rect 730 -1991 731 -1990
rect 1150 -1991 1151 -1990
rect 1160 -1991 1161 -1990
rect 1591 -1991 1592 -1990
rect 352 -1993 353 -1992
rect 408 -1993 409 -1992
rect 576 -1993 577 -1992
rect 695 -1993 696 -1992
rect 919 -1993 920 -1992
rect 1787 -1993 1788 -1992
rect 30 -1995 31 -1994
rect 576 -1995 577 -1994
rect 681 -1995 682 -1994
rect 688 -1995 689 -1994
rect 961 -1995 962 -1994
rect 1150 -1995 1151 -1994
rect 30 -1997 31 -1996
rect 331 -1997 332 -1996
rect 681 -1997 682 -1996
rect 765 -1997 766 -1996
rect 44 -1999 45 -1998
rect 331 -1999 332 -1998
rect 744 -1999 745 -1998
rect 765 -1999 766 -1998
rect 44 -2001 45 -2000
rect 530 -2001 531 -2000
rect 660 -2001 661 -2000
rect 744 -2001 745 -2000
rect 124 -2003 125 -2002
rect 352 -2003 353 -2002
rect 520 -2003 521 -2002
rect 660 -2003 661 -2002
rect 513 -2005 514 -2004
rect 520 -2005 521 -2004
rect 450 -2007 451 -2006
rect 513 -2007 514 -2006
rect 450 -2009 451 -2008
rect 569 -2009 570 -2008
rect 121 -2011 122 -2010
rect 569 -2011 570 -2010
rect 121 -2013 122 -2012
rect 1479 -2013 1480 -2012
rect 656 -2015 657 -2014
rect 1479 -2015 1480 -2014
rect 37 -2026 38 -2025
rect 625 -2026 626 -2025
rect 667 -2026 668 -2025
rect 670 -2026 671 -2025
rect 702 -2026 703 -2025
rect 957 -2026 958 -2025
rect 964 -2026 965 -2025
rect 1052 -2026 1053 -2025
rect 1062 -2026 1063 -2025
rect 1080 -2026 1081 -2025
rect 1139 -2026 1140 -2025
rect 1437 -2026 1438 -2025
rect 1479 -2026 1480 -2025
rect 1748 -2026 1749 -2025
rect 44 -2028 45 -2027
rect 712 -2028 713 -2027
rect 719 -2028 720 -2027
rect 926 -2028 927 -2027
rect 929 -2028 930 -2027
rect 1430 -2028 1431 -2027
rect 1591 -2028 1592 -2027
rect 1594 -2028 1595 -2027
rect 1713 -2028 1714 -2027
rect 1794 -2028 1795 -2027
rect 44 -2030 45 -2029
rect 180 -2030 181 -2029
rect 222 -2030 223 -2029
rect 247 -2030 248 -2029
rect 278 -2030 279 -2029
rect 1164 -2030 1165 -2029
rect 1195 -2030 1196 -2029
rect 1444 -2030 1445 -2029
rect 1591 -2030 1592 -2029
rect 1605 -2030 1606 -2029
rect 1745 -2030 1746 -2029
rect 1780 -2030 1781 -2029
rect 51 -2032 52 -2031
rect 177 -2032 178 -2031
rect 229 -2032 230 -2031
rect 1199 -2032 1200 -2031
rect 1213 -2032 1214 -2031
rect 1682 -2032 1683 -2031
rect 51 -2034 52 -2033
rect 275 -2034 276 -2033
rect 331 -2034 332 -2033
rect 471 -2034 472 -2033
rect 516 -2034 517 -2033
rect 940 -2034 941 -2033
rect 954 -2034 955 -2033
rect 1339 -2034 1340 -2033
rect 1423 -2034 1424 -2033
rect 1437 -2034 1438 -2033
rect 1444 -2034 1445 -2033
rect 1521 -2034 1522 -2033
rect 1682 -2034 1683 -2033
rect 1710 -2034 1711 -2033
rect 61 -2036 62 -2035
rect 1094 -2036 1095 -2035
rect 1157 -2036 1158 -2035
rect 1479 -2036 1480 -2035
rect 72 -2038 73 -2037
rect 201 -2038 202 -2037
rect 240 -2038 241 -2037
rect 250 -2038 251 -2037
rect 331 -2038 332 -2037
rect 460 -2038 461 -2037
rect 464 -2038 465 -2037
rect 506 -2038 507 -2037
rect 520 -2038 521 -2037
rect 523 -2038 524 -2037
rect 555 -2038 556 -2037
rect 586 -2038 587 -2037
rect 590 -2038 591 -2037
rect 597 -2038 598 -2037
rect 614 -2038 615 -2037
rect 975 -2038 976 -2037
rect 996 -2038 997 -2037
rect 1339 -2038 1340 -2037
rect 1395 -2038 1396 -2037
rect 1423 -2038 1424 -2037
rect 1430 -2038 1431 -2037
rect 1514 -2038 1515 -2037
rect 72 -2040 73 -2039
rect 261 -2040 262 -2039
rect 338 -2040 339 -2039
rect 593 -2040 594 -2039
rect 667 -2040 668 -2039
rect 730 -2040 731 -2039
rect 751 -2040 752 -2039
rect 894 -2040 895 -2039
rect 898 -2040 899 -2039
rect 1297 -2040 1298 -2039
rect 1314 -2040 1315 -2039
rect 1703 -2040 1704 -2039
rect 100 -2042 101 -2041
rect 422 -2042 423 -2041
rect 520 -2042 521 -2041
rect 534 -2042 535 -2041
rect 558 -2042 559 -2041
rect 1521 -2042 1522 -2041
rect 1703 -2042 1704 -2041
rect 1724 -2042 1725 -2041
rect 103 -2044 104 -2043
rect 863 -2044 864 -2043
rect 877 -2044 878 -2043
rect 961 -2044 962 -2043
rect 996 -2044 997 -2043
rect 1178 -2044 1179 -2043
rect 1195 -2044 1196 -2043
rect 1668 -2044 1669 -2043
rect 1724 -2044 1725 -2043
rect 1787 -2044 1788 -2043
rect 103 -2046 104 -2045
rect 191 -2046 192 -2045
rect 205 -2046 206 -2045
rect 464 -2046 465 -2045
rect 702 -2046 703 -2045
rect 1451 -2046 1452 -2045
rect 1514 -2046 1515 -2045
rect 1570 -2046 1571 -2045
rect 1594 -2046 1595 -2045
rect 1605 -2046 1606 -2045
rect 1626 -2046 1627 -2045
rect 1668 -2046 1669 -2045
rect 110 -2048 111 -2047
rect 149 -2048 150 -2047
rect 177 -2048 178 -2047
rect 583 -2048 584 -2047
rect 751 -2048 752 -2047
rect 772 -2048 773 -2047
rect 786 -2048 787 -2047
rect 992 -2048 993 -2047
rect 999 -2048 1000 -2047
rect 1738 -2048 1739 -2047
rect 114 -2050 115 -2049
rect 597 -2050 598 -2049
rect 761 -2050 762 -2049
rect 835 -2050 836 -2049
rect 856 -2050 857 -2049
rect 863 -2050 864 -2049
rect 887 -2050 888 -2049
rect 1619 -2050 1620 -2049
rect 1626 -2050 1627 -2049
rect 1661 -2050 1662 -2049
rect 1738 -2050 1739 -2049
rect 1808 -2050 1809 -2049
rect 114 -2052 115 -2051
rect 653 -2052 654 -2051
rect 786 -2052 787 -2051
rect 884 -2052 885 -2051
rect 905 -2052 906 -2051
rect 954 -2052 955 -2051
rect 999 -2052 1000 -2051
rect 1115 -2052 1116 -2051
rect 1157 -2052 1158 -2051
rect 1171 -2052 1172 -2051
rect 1199 -2052 1200 -2051
rect 1332 -2052 1333 -2051
rect 1395 -2052 1396 -2051
rect 1409 -2052 1410 -2051
rect 1451 -2052 1452 -2051
rect 1458 -2052 1459 -2051
rect 1570 -2052 1571 -2051
rect 1577 -2052 1578 -2051
rect 1619 -2052 1620 -2051
rect 1640 -2052 1641 -2051
rect 1661 -2052 1662 -2051
rect 1759 -2052 1760 -2051
rect 121 -2054 122 -2053
rect 1500 -2054 1501 -2053
rect 1507 -2054 1508 -2053
rect 1640 -2054 1641 -2053
rect 121 -2056 122 -2055
rect 457 -2056 458 -2055
rect 572 -2056 573 -2055
rect 653 -2056 654 -2055
rect 695 -2056 696 -2055
rect 884 -2056 885 -2055
rect 912 -2056 913 -2055
rect 940 -2056 941 -2055
rect 1017 -2056 1018 -2055
rect 1038 -2056 1039 -2055
rect 1052 -2056 1053 -2055
rect 1101 -2056 1102 -2055
rect 1164 -2056 1165 -2055
rect 1248 -2056 1249 -2055
rect 1293 -2056 1294 -2055
rect 1367 -2056 1368 -2055
rect 1409 -2056 1410 -2055
rect 1416 -2056 1417 -2055
rect 1458 -2056 1459 -2055
rect 1528 -2056 1529 -2055
rect 1577 -2056 1578 -2055
rect 1598 -2056 1599 -2055
rect 124 -2058 125 -2057
rect 205 -2058 206 -2057
rect 219 -2058 220 -2057
rect 1297 -2058 1298 -2057
rect 1332 -2058 1333 -2057
rect 1388 -2058 1389 -2057
rect 1500 -2058 1501 -2057
rect 1696 -2058 1697 -2057
rect 124 -2060 125 -2059
rect 310 -2060 311 -2059
rect 338 -2060 339 -2059
rect 1108 -2060 1109 -2059
rect 1171 -2060 1172 -2059
rect 1241 -2060 1242 -2059
rect 1283 -2060 1284 -2059
rect 1367 -2060 1368 -2059
rect 1507 -2060 1508 -2059
rect 1563 -2060 1564 -2059
rect 1584 -2060 1585 -2059
rect 1598 -2060 1599 -2059
rect 1689 -2060 1690 -2059
rect 1696 -2060 1697 -2059
rect 131 -2062 132 -2061
rect 562 -2062 563 -2061
rect 569 -2062 570 -2061
rect 1248 -2062 1249 -2061
rect 1283 -2062 1284 -2061
rect 1318 -2062 1319 -2061
rect 1563 -2062 1564 -2061
rect 1612 -2062 1613 -2061
rect 1689 -2062 1690 -2061
rect 1717 -2062 1718 -2061
rect 131 -2064 132 -2063
rect 1654 -2064 1655 -2063
rect 135 -2066 136 -2065
rect 275 -2066 276 -2065
rect 359 -2066 360 -2065
rect 387 -2066 388 -2065
rect 394 -2066 395 -2065
rect 803 -2066 804 -2065
rect 817 -2066 818 -2065
rect 870 -2066 871 -2065
rect 873 -2066 874 -2065
rect 1528 -2066 1529 -2065
rect 1612 -2066 1613 -2065
rect 1647 -2066 1648 -2065
rect 1654 -2066 1655 -2065
rect 1752 -2066 1753 -2065
rect 30 -2068 31 -2067
rect 135 -2068 136 -2067
rect 142 -2068 143 -2067
rect 905 -2068 906 -2067
rect 912 -2068 913 -2067
rect 947 -2068 948 -2067
rect 968 -2068 969 -2067
rect 1108 -2068 1109 -2067
rect 1241 -2068 1242 -2067
rect 1276 -2068 1277 -2067
rect 1318 -2068 1319 -2067
rect 1381 -2068 1382 -2067
rect 1647 -2068 1648 -2067
rect 1731 -2068 1732 -2067
rect 30 -2070 31 -2069
rect 96 -2070 97 -2069
rect 142 -2070 143 -2069
rect 723 -2070 724 -2069
rect 793 -2070 794 -2069
rect 828 -2070 829 -2069
rect 831 -2070 832 -2069
rect 1255 -2070 1256 -2069
rect 1381 -2070 1382 -2069
rect 1542 -2070 1543 -2069
rect 1731 -2070 1732 -2069
rect 1801 -2070 1802 -2069
rect 145 -2072 146 -2071
rect 1003 -2072 1004 -2071
rect 1024 -2072 1025 -2071
rect 1115 -2072 1116 -2071
rect 1255 -2072 1256 -2071
rect 1311 -2072 1312 -2071
rect 184 -2074 185 -2073
rect 310 -2074 311 -2073
rect 317 -2074 318 -2073
rect 359 -2074 360 -2073
rect 366 -2074 367 -2073
rect 509 -2074 510 -2073
rect 548 -2074 549 -2073
rect 1584 -2074 1585 -2073
rect 184 -2076 185 -2075
rect 212 -2076 213 -2075
rect 233 -2076 234 -2075
rect 877 -2076 878 -2075
rect 922 -2076 923 -2075
rect 1185 -2076 1186 -2075
rect 1290 -2076 1291 -2075
rect 1542 -2076 1543 -2075
rect 65 -2078 66 -2077
rect 212 -2078 213 -2077
rect 240 -2078 241 -2077
rect 292 -2078 293 -2077
rect 317 -2078 318 -2077
rect 324 -2078 325 -2077
rect 366 -2078 367 -2077
rect 485 -2078 486 -2077
rect 541 -2078 542 -2077
rect 548 -2078 549 -2077
rect 628 -2078 629 -2077
rect 723 -2078 724 -2077
rect 796 -2078 797 -2077
rect 1213 -2078 1214 -2077
rect 65 -2080 66 -2079
rect 705 -2080 706 -2079
rect 709 -2080 710 -2079
rect 1017 -2080 1018 -2079
rect 1024 -2080 1025 -2079
rect 1143 -2080 1144 -2079
rect 1185 -2080 1186 -2079
rect 1269 -2080 1270 -2079
rect 86 -2082 87 -2081
rect 233 -2082 234 -2081
rect 247 -2082 248 -2081
rect 471 -2082 472 -2081
rect 541 -2082 542 -2081
rect 821 -2082 822 -2081
rect 835 -2082 836 -2081
rect 1027 -2082 1028 -2081
rect 1073 -2082 1074 -2081
rect 1136 -2082 1137 -2081
rect 1143 -2082 1144 -2081
rect 1304 -2082 1305 -2081
rect 86 -2084 87 -2083
rect 625 -2084 626 -2083
rect 695 -2084 696 -2083
rect 737 -2084 738 -2083
rect 821 -2084 822 -2083
rect 1472 -2084 1473 -2083
rect 191 -2086 192 -2085
rect 450 -2086 451 -2085
rect 457 -2086 458 -2085
rect 604 -2086 605 -2085
rect 681 -2086 682 -2085
rect 737 -2086 738 -2085
rect 856 -2086 857 -2085
rect 891 -2086 892 -2085
rect 919 -2086 920 -2085
rect 1290 -2086 1291 -2085
rect 1304 -2086 1305 -2085
rect 1360 -2086 1361 -2085
rect 1472 -2086 1473 -2085
rect 1493 -2086 1494 -2085
rect 93 -2088 94 -2087
rect 919 -2088 920 -2087
rect 933 -2088 934 -2087
rect 968 -2088 969 -2087
rect 989 -2088 990 -2087
rect 1276 -2088 1277 -2087
rect 1493 -2088 1494 -2087
rect 1556 -2088 1557 -2087
rect 93 -2090 94 -2089
rect 1633 -2090 1634 -2089
rect 163 -2092 164 -2091
rect 604 -2092 605 -2091
rect 660 -2092 661 -2091
rect 681 -2092 682 -2091
rect 807 -2092 808 -2091
rect 933 -2092 934 -2091
rect 947 -2092 948 -2091
rect 982 -2092 983 -2091
rect 1031 -2092 1032 -2091
rect 1073 -2092 1074 -2091
rect 1080 -2092 1081 -2091
rect 1129 -2092 1130 -2091
rect 1262 -2092 1263 -2091
rect 1360 -2092 1361 -2091
rect 1486 -2092 1487 -2091
rect 1556 -2092 1557 -2091
rect 1633 -2092 1634 -2091
rect 1675 -2092 1676 -2091
rect 163 -2094 164 -2093
rect 975 -2094 976 -2093
rect 978 -2094 979 -2093
rect 1262 -2094 1263 -2093
rect 1269 -2094 1270 -2093
rect 1325 -2094 1326 -2093
rect 1675 -2094 1676 -2093
rect 1766 -2094 1767 -2093
rect 198 -2096 199 -2095
rect 387 -2096 388 -2095
rect 394 -2096 395 -2095
rect 513 -2096 514 -2095
rect 555 -2096 556 -2095
rect 989 -2096 990 -2095
rect 1010 -2096 1011 -2095
rect 1031 -2096 1032 -2095
rect 1087 -2096 1088 -2095
rect 1416 -2096 1417 -2095
rect 198 -2098 199 -2097
rect 219 -2098 220 -2097
rect 254 -2098 255 -2097
rect 562 -2098 563 -2097
rect 583 -2098 584 -2097
rect 1486 -2098 1487 -2097
rect 254 -2100 255 -2099
rect 576 -2100 577 -2099
rect 807 -2100 808 -2099
rect 849 -2100 850 -2099
rect 891 -2100 892 -2099
rect 1132 -2100 1133 -2099
rect 1325 -2100 1326 -2099
rect 1353 -2100 1354 -2099
rect 156 -2102 157 -2101
rect 576 -2102 577 -2101
rect 716 -2102 717 -2101
rect 1353 -2102 1354 -2101
rect 58 -2104 59 -2103
rect 156 -2104 157 -2103
rect 268 -2104 269 -2103
rect 422 -2104 423 -2103
rect 429 -2104 430 -2103
rect 569 -2104 570 -2103
rect 716 -2104 717 -2103
rect 1192 -2104 1193 -2103
rect 226 -2106 227 -2105
rect 268 -2106 269 -2105
rect 282 -2106 283 -2105
rect 485 -2106 486 -2105
rect 814 -2106 815 -2105
rect 849 -2106 850 -2105
rect 982 -2106 983 -2105
rect 1059 -2106 1060 -2105
rect 1087 -2106 1088 -2105
rect 1227 -2106 1228 -2105
rect 226 -2108 227 -2107
rect 1178 -2108 1179 -2107
rect 1227 -2108 1228 -2107
rect 1710 -2108 1711 -2107
rect 282 -2110 283 -2109
rect 527 -2110 528 -2109
rect 1010 -2110 1011 -2109
rect 1374 -2110 1375 -2109
rect 289 -2112 290 -2111
rect 660 -2112 661 -2111
rect 1059 -2112 1060 -2111
rect 1388 -2112 1389 -2111
rect 170 -2114 171 -2113
rect 289 -2114 290 -2113
rect 324 -2114 325 -2113
rect 373 -2114 374 -2113
rect 380 -2114 381 -2113
rect 814 -2114 815 -2113
rect 1094 -2114 1095 -2113
rect 1122 -2114 1123 -2113
rect 1129 -2114 1130 -2113
rect 1773 -2114 1774 -2113
rect 170 -2116 171 -2115
rect 478 -2116 479 -2115
rect 527 -2116 528 -2115
rect 779 -2116 780 -2115
rect 1101 -2116 1102 -2115
rect 1150 -2116 1151 -2115
rect 1374 -2116 1375 -2115
rect 1465 -2116 1466 -2115
rect 107 -2118 108 -2117
rect 1465 -2118 1466 -2117
rect 107 -2120 108 -2119
rect 688 -2120 689 -2119
rect 758 -2120 759 -2119
rect 1150 -2120 1151 -2119
rect 345 -2122 346 -2121
rect 478 -2122 479 -2121
rect 499 -2122 500 -2121
rect 688 -2122 689 -2121
rect 765 -2122 766 -2121
rect 779 -2122 780 -2121
rect 345 -2124 346 -2123
rect 443 -2124 444 -2123
rect 499 -2124 500 -2123
rect 611 -2124 612 -2123
rect 765 -2124 766 -2123
rect 800 -2124 801 -2123
rect 303 -2126 304 -2125
rect 443 -2126 444 -2125
rect 492 -2126 493 -2125
rect 611 -2126 612 -2125
rect 303 -2128 304 -2127
rect 901 -2128 902 -2127
rect 352 -2130 353 -2129
rect 758 -2130 759 -2129
rect 352 -2132 353 -2131
rect 513 -2132 514 -2131
rect 373 -2134 374 -2133
rect 1346 -2134 1347 -2133
rect 128 -2136 129 -2135
rect 1346 -2136 1347 -2135
rect 128 -2138 129 -2137
rect 261 -2138 262 -2137
rect 380 -2138 381 -2137
rect 646 -2138 647 -2137
rect 401 -2140 402 -2139
rect 492 -2140 493 -2139
rect 646 -2140 647 -2139
rect 674 -2140 675 -2139
rect 79 -2142 80 -2141
rect 401 -2142 402 -2141
rect 408 -2142 409 -2141
rect 450 -2142 451 -2141
rect 674 -2142 675 -2141
rect 1125 -2142 1126 -2141
rect 79 -2144 80 -2143
rect 415 -2144 416 -2143
rect 418 -2144 419 -2143
rect 1003 -2144 1004 -2143
rect 408 -2146 409 -2145
rect 628 -2146 629 -2145
rect 429 -2148 430 -2147
rect 1311 -2148 1312 -2147
rect 436 -2150 437 -2149
rect 772 -2150 773 -2149
rect 436 -2152 437 -2151
rect 639 -2152 640 -2151
rect 618 -2154 619 -2153
rect 639 -2154 640 -2153
rect 618 -2156 619 -2155
rect 1045 -2156 1046 -2155
rect 1045 -2158 1046 -2157
rect 1220 -2158 1221 -2157
rect 1206 -2160 1207 -2159
rect 1220 -2160 1221 -2159
rect 1206 -2162 1207 -2161
rect 1234 -2162 1235 -2161
rect 1234 -2164 1235 -2163
rect 1402 -2164 1403 -2163
rect 1402 -2166 1403 -2165
rect 1535 -2166 1536 -2165
rect 1535 -2168 1536 -2167
rect 1549 -2168 1550 -2167
rect 152 -2170 153 -2169
rect 1549 -2170 1550 -2169
rect 51 -2181 52 -2180
rect 415 -2181 416 -2180
rect 418 -2181 419 -2180
rect 800 -2181 801 -2180
rect 803 -2181 804 -2180
rect 1689 -2181 1690 -2180
rect 1696 -2181 1697 -2180
rect 1710 -2181 1711 -2180
rect 58 -2183 59 -2182
rect 135 -2183 136 -2182
rect 145 -2183 146 -2182
rect 905 -2183 906 -2182
rect 940 -2183 941 -2182
rect 1059 -2183 1060 -2182
rect 1125 -2183 1126 -2182
rect 1423 -2183 1424 -2182
rect 1640 -2183 1641 -2182
rect 1717 -2183 1718 -2182
rect 72 -2185 73 -2184
rect 628 -2185 629 -2184
rect 660 -2185 661 -2184
rect 828 -2185 829 -2184
rect 866 -2185 867 -2184
rect 1339 -2185 1340 -2184
rect 1409 -2185 1410 -2184
rect 1412 -2185 1413 -2184
rect 1650 -2185 1651 -2184
rect 1668 -2185 1669 -2184
rect 1671 -2185 1672 -2184
rect 1738 -2185 1739 -2184
rect 93 -2187 94 -2186
rect 310 -2187 311 -2186
rect 317 -2187 318 -2186
rect 376 -2187 377 -2186
rect 380 -2187 381 -2186
rect 926 -2187 927 -2186
rect 943 -2187 944 -2186
rect 1087 -2187 1088 -2186
rect 1132 -2187 1133 -2186
rect 1682 -2187 1683 -2186
rect 1689 -2187 1690 -2186
rect 1724 -2187 1725 -2186
rect 93 -2189 94 -2188
rect 1202 -2189 1203 -2188
rect 1262 -2189 1263 -2188
rect 1682 -2189 1683 -2188
rect 1696 -2189 1697 -2188
rect 1731 -2189 1732 -2188
rect 100 -2191 101 -2190
rect 1041 -2191 1042 -2190
rect 1059 -2191 1060 -2190
rect 1066 -2191 1067 -2190
rect 1087 -2191 1088 -2190
rect 1122 -2191 1123 -2190
rect 1150 -2191 1151 -2190
rect 1339 -2191 1340 -2190
rect 1388 -2191 1389 -2190
rect 1668 -2191 1669 -2190
rect 61 -2193 62 -2192
rect 100 -2193 101 -2192
rect 107 -2193 108 -2192
rect 408 -2193 409 -2192
rect 492 -2193 493 -2192
rect 583 -2193 584 -2192
rect 586 -2193 587 -2192
rect 933 -2193 934 -2192
rect 975 -2193 976 -2192
rect 1367 -2193 1368 -2192
rect 1388 -2193 1389 -2192
rect 1444 -2193 1445 -2192
rect 110 -2195 111 -2194
rect 198 -2195 199 -2194
rect 201 -2195 202 -2194
rect 422 -2195 423 -2194
rect 499 -2195 500 -2194
rect 824 -2195 825 -2194
rect 873 -2195 874 -2194
rect 1297 -2195 1298 -2194
rect 1311 -2195 1312 -2194
rect 1507 -2195 1508 -2194
rect 72 -2197 73 -2196
rect 873 -2197 874 -2196
rect 877 -2197 878 -2196
rect 926 -2197 927 -2196
rect 933 -2197 934 -2196
rect 982 -2197 983 -2196
rect 999 -2197 1000 -2196
rect 1080 -2197 1081 -2196
rect 1150 -2197 1151 -2196
rect 1720 -2197 1721 -2196
rect 114 -2199 115 -2198
rect 422 -2199 423 -2198
rect 499 -2199 500 -2198
rect 506 -2199 507 -2198
rect 513 -2199 514 -2198
rect 1122 -2199 1123 -2198
rect 1174 -2199 1175 -2198
rect 1248 -2199 1249 -2198
rect 1262 -2199 1263 -2198
rect 1353 -2199 1354 -2198
rect 1409 -2199 1410 -2198
rect 1486 -2199 1487 -2198
rect 1507 -2199 1508 -2198
rect 1542 -2199 1543 -2198
rect 114 -2201 115 -2200
rect 614 -2201 615 -2200
rect 618 -2201 619 -2200
rect 670 -2201 671 -2200
rect 688 -2201 689 -2200
rect 870 -2201 871 -2200
rect 877 -2201 878 -2200
rect 1227 -2201 1228 -2200
rect 1248 -2201 1249 -2200
rect 1269 -2201 1270 -2200
rect 1311 -2201 1312 -2200
rect 1332 -2201 1333 -2200
rect 1353 -2201 1354 -2200
rect 1465 -2201 1466 -2200
rect 1542 -2201 1543 -2200
rect 1598 -2201 1599 -2200
rect 121 -2203 122 -2202
rect 457 -2203 458 -2202
rect 506 -2203 507 -2202
rect 576 -2203 577 -2202
rect 583 -2203 584 -2202
rect 590 -2203 591 -2202
rect 604 -2203 605 -2202
rect 838 -2203 839 -2202
rect 905 -2203 906 -2202
rect 961 -2203 962 -2202
rect 975 -2203 976 -2202
rect 1038 -2203 1039 -2202
rect 1066 -2203 1067 -2202
rect 1108 -2203 1109 -2202
rect 1227 -2203 1228 -2202
rect 1416 -2203 1417 -2202
rect 1444 -2203 1445 -2202
rect 1451 -2203 1452 -2202
rect 1598 -2203 1599 -2202
rect 1633 -2203 1634 -2202
rect 44 -2205 45 -2204
rect 457 -2205 458 -2204
rect 495 -2205 496 -2204
rect 590 -2205 591 -2204
rect 611 -2205 612 -2204
rect 632 -2205 633 -2204
rect 660 -2205 661 -2204
rect 912 -2205 913 -2204
rect 961 -2205 962 -2204
rect 1003 -2205 1004 -2204
rect 1020 -2205 1021 -2204
rect 1297 -2205 1298 -2204
rect 1318 -2205 1319 -2204
rect 1367 -2205 1368 -2204
rect 1374 -2205 1375 -2204
rect 1465 -2205 1466 -2204
rect 44 -2207 45 -2206
rect 96 -2207 97 -2206
rect 128 -2207 129 -2206
rect 135 -2207 136 -2206
rect 156 -2207 157 -2206
rect 408 -2207 409 -2206
rect 513 -2207 514 -2206
rect 520 -2207 521 -2206
rect 534 -2207 535 -2206
rect 558 -2207 559 -2206
rect 618 -2207 619 -2206
rect 646 -2207 647 -2206
rect 688 -2207 689 -2206
rect 807 -2207 808 -2206
rect 817 -2207 818 -2206
rect 1640 -2207 1641 -2206
rect 128 -2209 129 -2208
rect 653 -2209 654 -2208
rect 691 -2209 692 -2208
rect 723 -2209 724 -2208
rect 761 -2209 762 -2208
rect 1017 -2209 1018 -2208
rect 1027 -2209 1028 -2208
rect 1220 -2209 1221 -2208
rect 1314 -2209 1315 -2208
rect 1374 -2209 1375 -2208
rect 1381 -2209 1382 -2208
rect 1416 -2209 1417 -2208
rect 131 -2211 132 -2210
rect 149 -2211 150 -2210
rect 156 -2211 157 -2210
rect 464 -2211 465 -2210
rect 520 -2211 521 -2210
rect 569 -2211 570 -2210
rect 597 -2211 598 -2210
rect 646 -2211 647 -2210
rect 698 -2211 699 -2210
rect 786 -2211 787 -2210
rect 807 -2211 808 -2210
rect 863 -2211 864 -2210
rect 978 -2211 979 -2210
rect 1703 -2211 1704 -2210
rect 65 -2213 66 -2212
rect 863 -2213 864 -2212
rect 982 -2213 983 -2212
rect 1052 -2213 1053 -2212
rect 1062 -2213 1063 -2212
rect 1318 -2213 1319 -2212
rect 1332 -2213 1333 -2212
rect 1430 -2213 1431 -2212
rect 65 -2215 66 -2214
rect 282 -2215 283 -2214
rect 285 -2215 286 -2214
rect 1528 -2215 1529 -2214
rect 124 -2217 125 -2216
rect 1430 -2217 1431 -2216
rect 1528 -2217 1529 -2216
rect 1626 -2217 1627 -2216
rect 138 -2219 139 -2218
rect 653 -2219 654 -2218
rect 709 -2219 710 -2218
rect 1451 -2219 1452 -2218
rect 1626 -2219 1627 -2218
rect 1675 -2219 1676 -2218
rect 163 -2221 164 -2220
rect 247 -2221 248 -2220
rect 254 -2221 255 -2220
rect 338 -2221 339 -2220
rect 359 -2221 360 -2220
rect 380 -2221 381 -2220
rect 394 -2221 395 -2220
rect 579 -2221 580 -2220
rect 600 -2221 601 -2220
rect 1052 -2221 1053 -2220
rect 1080 -2221 1081 -2220
rect 1136 -2221 1137 -2220
rect 1381 -2221 1382 -2220
rect 1395 -2221 1396 -2220
rect 163 -2223 164 -2222
rect 737 -2223 738 -2222
rect 786 -2223 787 -2222
rect 849 -2223 850 -2222
rect 1003 -2223 1004 -2222
rect 1073 -2223 1074 -2222
rect 1108 -2223 1109 -2222
rect 1195 -2223 1196 -2222
rect 1395 -2223 1396 -2222
rect 1437 -2223 1438 -2222
rect 170 -2225 171 -2224
rect 415 -2225 416 -2224
rect 464 -2225 465 -2224
rect 667 -2225 668 -2224
rect 674 -2225 675 -2224
rect 849 -2225 850 -2224
rect 1017 -2225 1018 -2224
rect 1472 -2225 1473 -2224
rect 30 -2227 31 -2226
rect 170 -2227 171 -2226
rect 177 -2227 178 -2226
rect 642 -2227 643 -2226
rect 667 -2227 668 -2226
rect 919 -2227 920 -2226
rect 1024 -2227 1025 -2226
rect 1220 -2227 1221 -2226
rect 1437 -2227 1438 -2226
rect 1556 -2227 1557 -2226
rect 30 -2229 31 -2228
rect 208 -2229 209 -2228
rect 212 -2229 213 -2228
rect 289 -2229 290 -2228
rect 296 -2229 297 -2228
rect 299 -2229 300 -2228
rect 303 -2229 304 -2228
rect 702 -2229 703 -2228
rect 709 -2229 710 -2228
rect 898 -2229 899 -2228
rect 1027 -2229 1028 -2228
rect 1164 -2229 1165 -2228
rect 1556 -2229 1557 -2228
rect 1577 -2229 1578 -2228
rect 177 -2231 178 -2230
rect 695 -2231 696 -2230
rect 716 -2231 717 -2230
rect 919 -2231 920 -2230
rect 1073 -2231 1074 -2230
rect 1178 -2231 1179 -2230
rect 1577 -2231 1578 -2230
rect 1661 -2231 1662 -2230
rect 215 -2233 216 -2232
rect 1010 -2233 1011 -2232
rect 1115 -2233 1116 -2232
rect 1633 -2233 1634 -2232
rect 226 -2235 227 -2234
rect 541 -2235 542 -2234
rect 555 -2235 556 -2234
rect 639 -2235 640 -2234
rect 681 -2235 682 -2234
rect 702 -2235 703 -2234
rect 737 -2235 738 -2234
rect 1024 -2235 1025 -2234
rect 1115 -2235 1116 -2234
rect 1157 -2235 1158 -2234
rect 1178 -2235 1179 -2234
rect 1290 -2235 1291 -2234
rect 1535 -2235 1536 -2234
rect 1661 -2235 1662 -2234
rect 226 -2237 227 -2236
rect 240 -2237 241 -2236
rect 261 -2237 262 -2236
rect 373 -2237 374 -2236
rect 394 -2237 395 -2236
rect 450 -2237 451 -2236
rect 509 -2237 510 -2236
rect 716 -2237 717 -2236
rect 821 -2237 822 -2236
rect 1423 -2237 1424 -2236
rect 229 -2239 230 -2238
rect 1472 -2239 1473 -2238
rect 233 -2241 234 -2240
rect 1136 -2241 1137 -2240
rect 1143 -2241 1144 -2240
rect 1164 -2241 1165 -2240
rect 1199 -2241 1200 -2240
rect 1290 -2241 1291 -2240
rect 233 -2243 234 -2242
rect 912 -2243 913 -2242
rect 989 -2243 990 -2242
rect 1157 -2243 1158 -2242
rect 1206 -2243 1207 -2242
rect 1535 -2243 1536 -2242
rect 240 -2245 241 -2244
rect 597 -2245 598 -2244
rect 625 -2245 626 -2244
rect 1479 -2245 1480 -2244
rect 261 -2247 262 -2246
rect 1192 -2247 1193 -2246
rect 1206 -2247 1207 -2246
rect 1241 -2247 1242 -2246
rect 1479 -2247 1480 -2246
rect 1493 -2247 1494 -2246
rect 268 -2249 269 -2248
rect 275 -2249 276 -2248
rect 282 -2249 283 -2248
rect 954 -2249 955 -2248
rect 989 -2249 990 -2248
rect 1094 -2249 1095 -2248
rect 1143 -2249 1144 -2248
rect 1185 -2249 1186 -2248
rect 1241 -2249 1242 -2248
rect 1276 -2249 1277 -2248
rect 1493 -2249 1494 -2248
rect 1570 -2249 1571 -2248
rect 268 -2251 269 -2250
rect 345 -2251 346 -2250
rect 359 -2251 360 -2250
rect 831 -2251 832 -2250
rect 898 -2251 899 -2250
rect 968 -2251 969 -2250
rect 996 -2251 997 -2250
rect 1185 -2251 1186 -2250
rect 1276 -2251 1277 -2250
rect 1458 -2251 1459 -2250
rect 1570 -2251 1571 -2250
rect 1591 -2251 1592 -2250
rect 79 -2253 80 -2252
rect 345 -2253 346 -2252
rect 401 -2253 402 -2252
rect 569 -2253 570 -2252
rect 628 -2253 629 -2252
rect 1269 -2253 1270 -2252
rect 1591 -2253 1592 -2252
rect 1612 -2253 1613 -2252
rect 79 -2255 80 -2254
rect 1521 -2255 1522 -2254
rect 1605 -2255 1606 -2254
rect 1612 -2255 1613 -2254
rect 103 -2257 104 -2256
rect 1458 -2257 1459 -2256
rect 1521 -2257 1522 -2256
rect 1584 -2257 1585 -2256
rect 1605 -2257 1606 -2256
rect 1647 -2257 1648 -2256
rect 250 -2259 251 -2258
rect 401 -2259 402 -2258
rect 471 -2259 472 -2258
rect 968 -2259 969 -2258
rect 996 -2259 997 -2258
rect 1101 -2259 1102 -2258
rect 1584 -2259 1585 -2258
rect 1619 -2259 1620 -2258
rect 1647 -2259 1648 -2258
rect 1675 -2259 1676 -2258
rect 296 -2261 297 -2260
rect 429 -2261 430 -2260
rect 471 -2261 472 -2260
rect 772 -2261 773 -2260
rect 821 -2261 822 -2260
rect 856 -2261 857 -2260
rect 929 -2261 930 -2260
rect 1192 -2261 1193 -2260
rect 1619 -2261 1620 -2260
rect 1654 -2261 1655 -2260
rect 257 -2263 258 -2262
rect 772 -2263 773 -2262
rect 856 -2263 857 -2262
rect 947 -2263 948 -2262
rect 954 -2263 955 -2262
rect 1213 -2263 1214 -2262
rect 1412 -2263 1413 -2262
rect 1486 -2263 1487 -2262
rect 303 -2265 304 -2264
rect 443 -2265 444 -2264
rect 534 -2265 535 -2264
rect 730 -2265 731 -2264
rect 814 -2265 815 -2264
rect 947 -2265 948 -2264
rect 1010 -2265 1011 -2264
rect 1713 -2265 1714 -2264
rect 191 -2267 192 -2266
rect 443 -2267 444 -2266
rect 541 -2267 542 -2266
rect 842 -2267 843 -2266
rect 1094 -2267 1095 -2266
rect 1171 -2267 1172 -2266
rect 1213 -2267 1214 -2266
rect 1255 -2267 1256 -2266
rect 149 -2269 150 -2268
rect 191 -2269 192 -2268
rect 310 -2269 311 -2268
rect 331 -2269 332 -2268
rect 338 -2269 339 -2268
rect 352 -2269 353 -2268
rect 548 -2269 549 -2268
rect 555 -2269 556 -2268
rect 632 -2269 633 -2268
rect 891 -2269 892 -2268
rect 1255 -2269 1256 -2268
rect 1346 -2269 1347 -2268
rect 86 -2271 87 -2270
rect 352 -2271 353 -2270
rect 681 -2271 682 -2270
rect 751 -2271 752 -2270
rect 758 -2271 759 -2270
rect 842 -2271 843 -2270
rect 1234 -2271 1235 -2270
rect 1346 -2271 1347 -2270
rect 86 -2273 87 -2272
rect 677 -2273 678 -2272
rect 705 -2273 706 -2272
rect 1101 -2273 1102 -2272
rect 1234 -2273 1235 -2272
rect 1325 -2273 1326 -2272
rect 152 -2275 153 -2274
rect 548 -2275 549 -2274
rect 730 -2275 731 -2274
rect 779 -2275 780 -2274
rect 793 -2275 794 -2274
rect 891 -2275 892 -2274
rect 1283 -2275 1284 -2274
rect 1325 -2275 1326 -2274
rect 205 -2277 206 -2276
rect 751 -2277 752 -2276
rect 814 -2277 815 -2276
rect 884 -2277 885 -2276
rect 1283 -2277 1284 -2276
rect 1304 -2277 1305 -2276
rect 317 -2279 318 -2278
rect 366 -2279 367 -2278
rect 527 -2279 528 -2278
rect 758 -2279 759 -2278
rect 884 -2279 885 -2278
rect 1045 -2279 1046 -2278
rect 1304 -2279 1305 -2278
rect 1360 -2279 1361 -2278
rect 142 -2281 143 -2280
rect 527 -2281 528 -2280
rect 604 -2281 605 -2280
rect 779 -2281 780 -2280
rect 1031 -2281 1032 -2280
rect 1045 -2281 1046 -2280
rect 1360 -2281 1361 -2280
rect 1402 -2281 1403 -2280
rect 142 -2283 143 -2282
rect 723 -2283 724 -2282
rect 744 -2283 745 -2282
rect 793 -2283 794 -2282
rect 1031 -2283 1032 -2282
rect 1129 -2283 1130 -2282
rect 1402 -2283 1403 -2282
rect 1500 -2283 1501 -2282
rect 205 -2285 206 -2284
rect 1129 -2285 1130 -2284
rect 1500 -2285 1501 -2284
rect 1514 -2285 1515 -2284
rect 324 -2287 325 -2286
rect 516 -2287 517 -2286
rect 744 -2287 745 -2286
rect 765 -2287 766 -2286
rect 324 -2289 325 -2288
rect 485 -2289 486 -2288
rect 765 -2289 766 -2288
rect 835 -2289 836 -2288
rect 331 -2291 332 -2290
rect 436 -2291 437 -2290
rect 485 -2291 486 -2290
rect 1038 -2291 1039 -2290
rect 366 -2293 367 -2292
rect 387 -2293 388 -2292
rect 436 -2293 437 -2292
rect 562 -2293 563 -2292
rect 835 -2293 836 -2292
rect 1514 -2293 1515 -2292
rect 37 -2295 38 -2294
rect 562 -2295 563 -2294
rect 387 -2297 388 -2296
rect 478 -2297 479 -2296
rect 450 -2299 451 -2298
rect 478 -2299 479 -2298
rect 30 -2310 31 -2309
rect 149 -2310 150 -2309
rect 205 -2310 206 -2309
rect 219 -2310 220 -2309
rect 254 -2310 255 -2309
rect 523 -2310 524 -2309
rect 548 -2310 549 -2309
rect 943 -2310 944 -2309
rect 971 -2310 972 -2309
rect 1094 -2310 1095 -2309
rect 1174 -2310 1175 -2309
rect 1493 -2310 1494 -2309
rect 1622 -2310 1623 -2309
rect 1696 -2310 1697 -2309
rect 51 -2312 52 -2311
rect 359 -2312 360 -2311
rect 387 -2312 388 -2311
rect 548 -2312 549 -2311
rect 576 -2312 577 -2311
rect 828 -2312 829 -2311
rect 835 -2312 836 -2311
rect 1451 -2312 1452 -2311
rect 1493 -2312 1494 -2311
rect 1542 -2312 1543 -2311
rect 1647 -2312 1648 -2311
rect 1689 -2312 1690 -2311
rect 65 -2314 66 -2313
rect 68 -2314 69 -2313
rect 79 -2314 80 -2313
rect 562 -2314 563 -2313
rect 597 -2314 598 -2313
rect 761 -2314 762 -2313
rect 779 -2314 780 -2313
rect 1346 -2314 1347 -2313
rect 1451 -2314 1452 -2313
rect 1654 -2314 1655 -2313
rect 65 -2316 66 -2315
rect 261 -2316 262 -2315
rect 285 -2316 286 -2315
rect 310 -2316 311 -2315
rect 317 -2316 318 -2315
rect 586 -2316 587 -2315
rect 625 -2316 626 -2315
rect 751 -2316 752 -2315
rect 821 -2316 822 -2315
rect 828 -2316 829 -2315
rect 859 -2316 860 -2315
rect 1430 -2316 1431 -2315
rect 1542 -2316 1543 -2315
rect 1584 -2316 1585 -2315
rect 79 -2318 80 -2317
rect 401 -2318 402 -2317
rect 415 -2318 416 -2317
rect 600 -2318 601 -2317
rect 635 -2318 636 -2317
rect 674 -2318 675 -2317
rect 677 -2318 678 -2317
rect 730 -2318 731 -2317
rect 740 -2318 741 -2317
rect 1633 -2318 1634 -2317
rect 128 -2320 129 -2319
rect 702 -2320 703 -2319
rect 705 -2320 706 -2319
rect 807 -2320 808 -2319
rect 866 -2320 867 -2319
rect 1248 -2320 1249 -2319
rect 1251 -2320 1252 -2319
rect 1325 -2320 1326 -2319
rect 1346 -2320 1347 -2319
rect 1374 -2320 1375 -2319
rect 1430 -2320 1431 -2319
rect 1458 -2320 1459 -2319
rect 1612 -2320 1613 -2319
rect 1633 -2320 1634 -2319
rect 114 -2322 115 -2321
rect 807 -2322 808 -2321
rect 873 -2322 874 -2321
rect 1304 -2322 1305 -2321
rect 1374 -2322 1375 -2321
rect 1395 -2322 1396 -2321
rect 1444 -2322 1445 -2321
rect 1458 -2322 1459 -2321
rect 1612 -2322 1613 -2321
rect 1640 -2322 1641 -2321
rect 114 -2324 115 -2323
rect 408 -2324 409 -2323
rect 450 -2324 451 -2323
rect 1136 -2324 1137 -2323
rect 1171 -2324 1172 -2323
rect 1654 -2324 1655 -2323
rect 135 -2326 136 -2325
rect 541 -2326 542 -2325
rect 562 -2326 563 -2325
rect 891 -2326 892 -2325
rect 912 -2326 913 -2325
rect 1290 -2326 1291 -2325
rect 1444 -2326 1445 -2325
rect 1472 -2326 1473 -2325
rect 149 -2328 150 -2327
rect 1066 -2328 1067 -2327
rect 1073 -2328 1074 -2327
rect 1136 -2328 1137 -2327
rect 1164 -2328 1165 -2327
rect 1171 -2328 1172 -2327
rect 1199 -2328 1200 -2327
rect 1535 -2328 1536 -2327
rect 208 -2330 209 -2329
rect 464 -2330 465 -2329
rect 492 -2330 493 -2329
rect 1041 -2330 1042 -2329
rect 1052 -2330 1053 -2329
rect 1094 -2330 1095 -2329
rect 1129 -2330 1130 -2329
rect 1584 -2330 1585 -2329
rect 215 -2332 216 -2331
rect 324 -2332 325 -2331
rect 359 -2332 360 -2331
rect 534 -2332 535 -2331
rect 541 -2332 542 -2331
rect 569 -2332 570 -2331
rect 579 -2332 580 -2331
rect 1052 -2332 1053 -2331
rect 1073 -2332 1074 -2331
rect 1080 -2332 1081 -2331
rect 1122 -2332 1123 -2331
rect 1129 -2332 1130 -2331
rect 1157 -2332 1158 -2331
rect 1164 -2332 1165 -2331
rect 1202 -2332 1203 -2331
rect 1381 -2332 1382 -2331
rect 1472 -2332 1473 -2331
rect 1507 -2332 1508 -2331
rect 1535 -2332 1536 -2331
rect 1591 -2332 1592 -2331
rect 86 -2334 87 -2333
rect 569 -2334 570 -2333
rect 590 -2334 591 -2333
rect 625 -2334 626 -2333
rect 639 -2334 640 -2333
rect 842 -2334 843 -2333
rect 891 -2334 892 -2333
rect 898 -2334 899 -2333
rect 912 -2334 913 -2333
rect 1293 -2334 1294 -2333
rect 1591 -2334 1592 -2333
rect 1605 -2334 1606 -2333
rect 72 -2336 73 -2335
rect 590 -2336 591 -2335
rect 639 -2336 640 -2335
rect 681 -2336 682 -2335
rect 684 -2336 685 -2335
rect 821 -2336 822 -2335
rect 842 -2336 843 -2335
rect 905 -2336 906 -2335
rect 915 -2336 916 -2335
rect 1416 -2336 1417 -2335
rect 1605 -2336 1606 -2335
rect 1671 -2336 1672 -2335
rect 72 -2338 73 -2337
rect 632 -2338 633 -2337
rect 667 -2338 668 -2337
rect 856 -2338 857 -2337
rect 989 -2338 990 -2337
rect 992 -2338 993 -2337
rect 1017 -2338 1018 -2337
rect 1108 -2338 1109 -2337
rect 1122 -2338 1123 -2337
rect 1577 -2338 1578 -2337
rect 86 -2340 87 -2339
rect 229 -2340 230 -2339
rect 233 -2340 234 -2339
rect 254 -2340 255 -2339
rect 261 -2340 262 -2339
rect 275 -2340 276 -2339
rect 289 -2340 290 -2339
rect 408 -2340 409 -2339
rect 436 -2340 437 -2339
rect 492 -2340 493 -2339
rect 495 -2340 496 -2339
rect 646 -2340 647 -2339
rect 681 -2340 682 -2339
rect 1157 -2340 1158 -2339
rect 1185 -2340 1186 -2339
rect 1507 -2340 1508 -2339
rect 117 -2342 118 -2341
rect 289 -2342 290 -2341
rect 296 -2342 297 -2341
rect 576 -2342 577 -2341
rect 632 -2342 633 -2341
rect 954 -2342 955 -2341
rect 975 -2342 976 -2341
rect 1108 -2342 1109 -2341
rect 1185 -2342 1186 -2341
rect 1367 -2342 1368 -2341
rect 142 -2344 143 -2343
rect 233 -2344 234 -2343
rect 247 -2344 248 -2343
rect 324 -2344 325 -2343
rect 373 -2344 374 -2343
rect 464 -2344 465 -2343
rect 478 -2344 479 -2343
rect 905 -2344 906 -2343
rect 975 -2344 976 -2343
rect 982 -2344 983 -2343
rect 989 -2344 990 -2343
rect 1003 -2344 1004 -2343
rect 1020 -2344 1021 -2343
rect 1059 -2344 1060 -2343
rect 1206 -2344 1207 -2343
rect 1244 -2344 1245 -2343
rect 1248 -2344 1249 -2343
rect 1626 -2344 1627 -2343
rect 142 -2346 143 -2345
rect 240 -2346 241 -2345
rect 247 -2346 248 -2345
rect 331 -2346 332 -2345
rect 373 -2346 374 -2345
rect 604 -2346 605 -2345
rect 688 -2346 689 -2345
rect 786 -2346 787 -2345
rect 849 -2346 850 -2345
rect 982 -2346 983 -2345
rect 1003 -2346 1004 -2345
rect 1031 -2346 1032 -2345
rect 1038 -2346 1039 -2345
rect 1388 -2346 1389 -2345
rect 1570 -2346 1571 -2345
rect 1626 -2346 1627 -2345
rect 170 -2348 171 -2347
rect 275 -2348 276 -2347
rect 282 -2348 283 -2347
rect 954 -2348 955 -2347
rect 996 -2348 997 -2347
rect 1031 -2348 1032 -2347
rect 1045 -2348 1046 -2347
rect 1080 -2348 1081 -2347
rect 1206 -2348 1207 -2347
rect 1363 -2348 1364 -2347
rect 1367 -2348 1368 -2347
rect 1500 -2348 1501 -2347
rect 170 -2350 171 -2349
rect 191 -2350 192 -2349
rect 219 -2350 220 -2349
rect 226 -2350 227 -2349
rect 240 -2350 241 -2349
rect 366 -2350 367 -2349
rect 380 -2350 381 -2349
rect 401 -2350 402 -2349
rect 422 -2350 423 -2349
rect 646 -2350 647 -2349
rect 691 -2350 692 -2349
rect 779 -2350 780 -2349
rect 786 -2350 787 -2349
rect 1668 -2350 1669 -2349
rect 184 -2352 185 -2351
rect 191 -2352 192 -2351
rect 226 -2352 227 -2351
rect 968 -2352 969 -2351
rect 1059 -2352 1060 -2351
rect 1227 -2352 1228 -2351
rect 1237 -2352 1238 -2351
rect 1486 -2352 1487 -2351
rect 184 -2354 185 -2353
rect 485 -2354 486 -2353
rect 506 -2354 507 -2353
rect 702 -2354 703 -2353
rect 709 -2354 710 -2353
rect 1045 -2354 1046 -2353
rect 1150 -2354 1151 -2353
rect 1227 -2354 1228 -2353
rect 1241 -2354 1242 -2353
rect 1479 -2354 1480 -2353
rect 1486 -2354 1487 -2353
rect 1650 -2354 1651 -2353
rect 268 -2356 269 -2355
rect 415 -2356 416 -2355
rect 422 -2356 423 -2355
rect 457 -2356 458 -2355
rect 506 -2356 507 -2355
rect 555 -2356 556 -2355
rect 604 -2356 605 -2355
rect 611 -2356 612 -2355
rect 621 -2356 622 -2355
rect 1500 -2356 1501 -2355
rect 1650 -2356 1651 -2355
rect 1661 -2356 1662 -2355
rect 268 -2358 269 -2357
rect 835 -2358 836 -2357
rect 838 -2358 839 -2357
rect 1570 -2358 1571 -2357
rect 1661 -2358 1662 -2357
rect 1682 -2358 1683 -2357
rect 282 -2360 283 -2359
rect 1479 -2360 1480 -2359
rect 296 -2362 297 -2361
rect 338 -2362 339 -2361
rect 345 -2362 346 -2361
rect 688 -2362 689 -2361
rect 695 -2362 696 -2361
rect 877 -2362 878 -2361
rect 947 -2362 948 -2361
rect 1038 -2362 1039 -2361
rect 1150 -2362 1151 -2361
rect 1381 -2362 1382 -2361
rect 1388 -2362 1389 -2361
rect 1409 -2362 1410 -2361
rect 100 -2364 101 -2363
rect 695 -2364 696 -2363
rect 709 -2364 710 -2363
rect 793 -2364 794 -2363
rect 800 -2364 801 -2363
rect 877 -2364 878 -2363
rect 947 -2364 948 -2363
rect 961 -2364 962 -2363
rect 992 -2364 993 -2363
rect 996 -2364 997 -2363
rect 1241 -2364 1242 -2363
rect 1297 -2364 1298 -2363
rect 1318 -2364 1319 -2363
rect 1416 -2364 1417 -2363
rect 100 -2366 101 -2365
rect 814 -2366 815 -2365
rect 870 -2366 871 -2365
rect 1297 -2366 1298 -2365
rect 1318 -2366 1319 -2365
rect 1332 -2366 1333 -2365
rect 1339 -2366 1340 -2365
rect 1409 -2366 1410 -2365
rect 310 -2368 311 -2367
rect 471 -2368 472 -2367
rect 509 -2368 510 -2367
rect 513 -2368 514 -2367
rect 534 -2368 535 -2367
rect 929 -2368 930 -2367
rect 1269 -2368 1270 -2367
rect 1325 -2368 1326 -2367
rect 1332 -2368 1333 -2367
rect 1353 -2368 1354 -2367
rect 58 -2370 59 -2369
rect 513 -2370 514 -2369
rect 611 -2370 612 -2369
rect 793 -2370 794 -2369
rect 870 -2370 871 -2369
rect 1024 -2370 1025 -2369
rect 1255 -2370 1256 -2369
rect 1269 -2370 1270 -2369
rect 1283 -2370 1284 -2369
rect 1304 -2370 1305 -2369
rect 1339 -2370 1340 -2369
rect 1360 -2370 1361 -2369
rect 44 -2372 45 -2371
rect 58 -2372 59 -2371
rect 317 -2372 318 -2371
rect 670 -2372 671 -2371
rect 716 -2372 717 -2371
rect 800 -2372 801 -2371
rect 926 -2372 927 -2371
rect 961 -2372 962 -2371
rect 1234 -2372 1235 -2371
rect 1255 -2372 1256 -2371
rect 1262 -2372 1263 -2371
rect 1283 -2372 1284 -2371
rect 1290 -2372 1291 -2371
rect 1528 -2372 1529 -2371
rect 44 -2374 45 -2373
rect 782 -2374 783 -2373
rect 898 -2374 899 -2373
rect 926 -2374 927 -2373
rect 1017 -2374 1018 -2373
rect 1234 -2374 1235 -2373
rect 1353 -2374 1354 -2373
rect 1423 -2374 1424 -2373
rect 1528 -2374 1529 -2373
rect 1549 -2374 1550 -2373
rect 331 -2376 332 -2375
rect 649 -2376 650 -2375
rect 653 -2376 654 -2375
rect 1024 -2376 1025 -2375
rect 1192 -2376 1193 -2375
rect 1423 -2376 1424 -2375
rect 1549 -2376 1550 -2375
rect 1556 -2376 1557 -2375
rect 107 -2378 108 -2377
rect 653 -2378 654 -2377
rect 660 -2378 661 -2377
rect 814 -2378 815 -2377
rect 1178 -2378 1179 -2377
rect 1192 -2378 1193 -2377
rect 1213 -2378 1214 -2377
rect 1262 -2378 1263 -2377
rect 1402 -2378 1403 -2377
rect 1556 -2378 1557 -2377
rect 138 -2380 139 -2379
rect 1178 -2380 1179 -2379
rect 1213 -2380 1214 -2379
rect 1521 -2380 1522 -2379
rect 163 -2382 164 -2381
rect 660 -2382 661 -2381
rect 723 -2382 724 -2381
rect 1066 -2382 1067 -2381
rect 1276 -2382 1277 -2381
rect 1402 -2382 1403 -2381
rect 1521 -2382 1522 -2381
rect 1563 -2382 1564 -2381
rect 163 -2384 164 -2383
rect 429 -2384 430 -2383
rect 436 -2384 437 -2383
rect 520 -2384 521 -2383
rect 583 -2384 584 -2383
rect 716 -2384 717 -2383
rect 723 -2384 724 -2383
rect 1675 -2384 1676 -2383
rect 338 -2386 339 -2385
rect 352 -2386 353 -2385
rect 366 -2386 367 -2385
rect 527 -2386 528 -2385
rect 730 -2386 731 -2385
rect 884 -2386 885 -2385
rect 1202 -2386 1203 -2385
rect 1276 -2386 1277 -2385
rect 1563 -2386 1564 -2385
rect 1598 -2386 1599 -2385
rect 156 -2388 157 -2387
rect 352 -2388 353 -2387
rect 380 -2388 381 -2387
rect 1104 -2388 1105 -2387
rect 1598 -2388 1599 -2387
rect 1619 -2388 1620 -2387
rect 156 -2390 157 -2389
rect 733 -2390 734 -2389
rect 747 -2390 748 -2389
rect 1395 -2390 1396 -2389
rect 345 -2392 346 -2391
rect 583 -2392 584 -2391
rect 751 -2392 752 -2391
rect 863 -2392 864 -2391
rect 387 -2394 388 -2393
rect 394 -2394 395 -2393
rect 404 -2394 405 -2393
rect 429 -2394 430 -2393
rect 443 -2394 444 -2393
rect 478 -2394 479 -2393
rect 520 -2394 521 -2393
rect 555 -2394 556 -2393
rect 744 -2394 745 -2393
rect 863 -2394 864 -2393
rect 128 -2396 129 -2395
rect 744 -2396 745 -2395
rect 758 -2396 759 -2395
rect 884 -2396 885 -2395
rect 443 -2398 444 -2397
rect 940 -2398 941 -2397
rect 450 -2400 451 -2399
rect 1619 -2400 1620 -2399
rect 453 -2402 454 -2401
rect 737 -2402 738 -2401
rect 758 -2402 759 -2401
rect 765 -2402 766 -2401
rect 775 -2402 776 -2401
rect 1577 -2402 1578 -2401
rect 394 -2404 395 -2403
rect 737 -2404 738 -2403
rect 765 -2404 766 -2403
rect 772 -2404 773 -2403
rect 933 -2404 934 -2403
rect 940 -2404 941 -2403
rect 457 -2406 458 -2405
rect 1010 -2406 1011 -2405
rect 471 -2408 472 -2407
rect 618 -2408 619 -2407
rect 642 -2408 643 -2407
rect 933 -2408 934 -2407
rect 1010 -2408 1011 -2407
rect 1101 -2408 1102 -2407
rect 121 -2410 122 -2409
rect 618 -2410 619 -2409
rect 121 -2412 122 -2411
rect 212 -2412 213 -2411
rect 527 -2412 528 -2411
rect 772 -2412 773 -2411
rect 198 -2414 199 -2413
rect 212 -2414 213 -2413
rect 93 -2416 94 -2415
rect 198 -2416 199 -2415
rect 93 -2418 94 -2417
rect 177 -2418 178 -2417
rect 152 -2420 153 -2419
rect 177 -2420 178 -2419
rect 44 -2431 45 -2430
rect 530 -2431 531 -2430
rect 562 -2431 563 -2430
rect 1395 -2431 1396 -2430
rect 1615 -2431 1616 -2430
rect 1633 -2431 1634 -2430
rect 93 -2433 94 -2432
rect 117 -2433 118 -2432
rect 121 -2433 122 -2432
rect 775 -2433 776 -2432
rect 831 -2433 832 -2432
rect 1213 -2433 1214 -2432
rect 1234 -2433 1235 -2432
rect 1587 -2433 1588 -2432
rect 1622 -2433 1623 -2432
rect 1661 -2433 1662 -2432
rect 93 -2435 94 -2434
rect 443 -2435 444 -2434
rect 471 -2435 472 -2434
rect 614 -2435 615 -2434
rect 674 -2435 675 -2434
rect 740 -2435 741 -2434
rect 747 -2435 748 -2434
rect 1577 -2435 1578 -2434
rect 1626 -2435 1627 -2434
rect 1643 -2435 1644 -2434
rect 107 -2437 108 -2436
rect 1514 -2437 1515 -2436
rect 1577 -2437 1578 -2436
rect 1584 -2437 1585 -2436
rect 107 -2439 108 -2438
rect 110 -2439 111 -2438
rect 121 -2439 122 -2438
rect 723 -2439 724 -2438
rect 737 -2439 738 -2438
rect 1227 -2439 1228 -2438
rect 1248 -2439 1249 -2438
rect 1605 -2439 1606 -2438
rect 135 -2441 136 -2440
rect 646 -2441 647 -2440
rect 674 -2441 675 -2440
rect 1027 -2441 1028 -2440
rect 1066 -2441 1067 -2440
rect 1122 -2441 1123 -2440
rect 1185 -2441 1186 -2440
rect 1213 -2441 1214 -2440
rect 1251 -2441 1252 -2440
rect 1409 -2441 1410 -2440
rect 1549 -2441 1550 -2440
rect 1605 -2441 1606 -2440
rect 135 -2443 136 -2442
rect 457 -2443 458 -2442
rect 520 -2443 521 -2442
rect 660 -2443 661 -2442
rect 681 -2443 682 -2442
rect 863 -2443 864 -2442
rect 901 -2443 902 -2442
rect 975 -2443 976 -2442
rect 989 -2443 990 -2442
rect 1066 -2443 1067 -2442
rect 1104 -2443 1105 -2442
rect 1262 -2443 1263 -2442
rect 1290 -2443 1291 -2442
rect 1416 -2443 1417 -2442
rect 1549 -2443 1550 -2442
rect 1570 -2443 1571 -2442
rect 142 -2445 143 -2444
rect 481 -2445 482 -2444
rect 572 -2445 573 -2444
rect 716 -2445 717 -2444
rect 723 -2445 724 -2444
rect 1188 -2445 1189 -2444
rect 1199 -2445 1200 -2444
rect 1437 -2445 1438 -2444
rect 142 -2447 143 -2446
rect 387 -2447 388 -2446
rect 394 -2447 395 -2446
rect 471 -2447 472 -2446
rect 569 -2447 570 -2446
rect 716 -2447 717 -2446
rect 733 -2447 734 -2446
rect 1570 -2447 1571 -2446
rect 163 -2449 164 -2448
rect 810 -2449 811 -2448
rect 821 -2449 822 -2448
rect 989 -2449 990 -2448
rect 1013 -2449 1014 -2448
rect 1528 -2449 1529 -2448
rect 163 -2451 164 -2450
rect 390 -2451 391 -2450
rect 394 -2451 395 -2450
rect 632 -2451 633 -2450
rect 639 -2451 640 -2450
rect 646 -2451 647 -2450
rect 681 -2451 682 -2450
rect 684 -2451 685 -2450
rect 688 -2451 689 -2450
rect 803 -2451 804 -2450
rect 821 -2451 822 -2450
rect 1405 -2451 1406 -2450
rect 1493 -2451 1494 -2450
rect 1528 -2451 1529 -2450
rect 170 -2453 171 -2452
rect 257 -2453 258 -2452
rect 282 -2453 283 -2452
rect 772 -2453 773 -2452
rect 835 -2453 836 -2452
rect 1045 -2453 1046 -2452
rect 1164 -2453 1165 -2452
rect 1199 -2453 1200 -2452
rect 1220 -2453 1221 -2452
rect 1290 -2453 1291 -2452
rect 1332 -2453 1333 -2452
rect 1395 -2453 1396 -2452
rect 1486 -2453 1487 -2452
rect 1493 -2453 1494 -2452
rect 51 -2455 52 -2454
rect 170 -2455 171 -2454
rect 219 -2455 220 -2454
rect 226 -2455 227 -2454
rect 229 -2455 230 -2454
rect 1650 -2455 1651 -2454
rect 51 -2457 52 -2456
rect 401 -2457 402 -2456
rect 404 -2457 405 -2456
rect 429 -2457 430 -2456
rect 583 -2457 584 -2456
rect 1486 -2457 1487 -2456
rect 114 -2459 115 -2458
rect 219 -2459 220 -2458
rect 240 -2459 241 -2458
rect 429 -2459 430 -2458
rect 583 -2459 584 -2458
rect 709 -2459 710 -2458
rect 740 -2459 741 -2458
rect 842 -2459 843 -2458
rect 849 -2459 850 -2458
rect 1297 -2459 1298 -2458
rect 1339 -2459 1340 -2458
rect 1409 -2459 1410 -2458
rect 58 -2461 59 -2460
rect 114 -2461 115 -2460
rect 128 -2461 129 -2460
rect 835 -2461 836 -2460
rect 849 -2461 850 -2460
rect 877 -2461 878 -2460
rect 919 -2461 920 -2460
rect 1325 -2461 1326 -2460
rect 1346 -2461 1347 -2460
rect 1416 -2461 1417 -2460
rect 58 -2463 59 -2462
rect 285 -2463 286 -2462
rect 303 -2463 304 -2462
rect 730 -2463 731 -2462
rect 758 -2463 759 -2462
rect 772 -2463 773 -2462
rect 828 -2463 829 -2462
rect 842 -2463 843 -2462
rect 852 -2463 853 -2462
rect 1108 -2463 1109 -2462
rect 1192 -2463 1193 -2462
rect 1297 -2463 1298 -2462
rect 1318 -2463 1319 -2462
rect 1325 -2463 1326 -2462
rect 1353 -2463 1354 -2462
rect 1437 -2463 1438 -2462
rect 79 -2465 80 -2464
rect 758 -2465 759 -2464
rect 856 -2465 857 -2464
rect 1514 -2465 1515 -2464
rect 79 -2467 80 -2466
rect 247 -2467 248 -2466
rect 254 -2467 255 -2466
rect 282 -2467 283 -2466
rect 303 -2467 304 -2466
rect 1125 -2467 1126 -2466
rect 1143 -2467 1144 -2466
rect 1192 -2467 1193 -2466
rect 1206 -2467 1207 -2466
rect 1339 -2467 1340 -2466
rect 1360 -2467 1361 -2466
rect 1563 -2467 1564 -2466
rect 247 -2469 248 -2468
rect 478 -2469 479 -2468
rect 576 -2469 577 -2468
rect 730 -2469 731 -2468
rect 793 -2469 794 -2468
rect 856 -2469 857 -2468
rect 929 -2469 930 -2468
rect 1402 -2469 1403 -2468
rect 1563 -2469 1564 -2468
rect 1612 -2469 1613 -2468
rect 254 -2471 255 -2470
rect 859 -2471 860 -2470
rect 933 -2471 934 -2470
rect 1108 -2471 1109 -2470
rect 1171 -2471 1172 -2470
rect 1360 -2471 1361 -2470
rect 1374 -2471 1375 -2470
rect 1381 -2471 1382 -2470
rect 1384 -2471 1385 -2470
rect 1591 -2471 1592 -2470
rect 338 -2473 339 -2472
rect 457 -2473 458 -2472
rect 523 -2473 524 -2472
rect 576 -2473 577 -2472
rect 586 -2473 587 -2472
rect 1227 -2473 1228 -2472
rect 1241 -2473 1242 -2472
rect 1346 -2473 1347 -2472
rect 324 -2475 325 -2474
rect 338 -2475 339 -2474
rect 359 -2475 360 -2474
rect 478 -2475 479 -2474
rect 600 -2475 601 -2474
rect 961 -2475 962 -2474
rect 1024 -2475 1025 -2474
rect 1101 -2475 1102 -2474
rect 1150 -2475 1151 -2474
rect 1171 -2475 1172 -2474
rect 1202 -2475 1203 -2474
rect 1241 -2475 1242 -2474
rect 1251 -2475 1252 -2474
rect 1262 -2475 1263 -2474
rect 1269 -2475 1270 -2474
rect 1318 -2475 1319 -2474
rect 233 -2477 234 -2476
rect 324 -2477 325 -2476
rect 359 -2477 360 -2476
rect 464 -2477 465 -2476
rect 604 -2477 605 -2476
rect 660 -2477 661 -2476
rect 667 -2477 668 -2476
rect 877 -2477 878 -2476
rect 905 -2477 906 -2476
rect 961 -2477 962 -2476
rect 1024 -2477 1025 -2476
rect 1507 -2477 1508 -2476
rect 233 -2479 234 -2478
rect 373 -2479 374 -2478
rect 380 -2479 381 -2478
rect 863 -2479 864 -2478
rect 898 -2479 899 -2478
rect 905 -2479 906 -2478
rect 947 -2479 948 -2478
rect 975 -2479 976 -2478
rect 1038 -2479 1039 -2478
rect 1185 -2479 1186 -2478
rect 1206 -2479 1207 -2478
rect 1640 -2479 1641 -2478
rect 296 -2481 297 -2480
rect 373 -2481 374 -2480
rect 380 -2481 381 -2480
rect 702 -2481 703 -2480
rect 709 -2481 710 -2480
rect 765 -2481 766 -2480
rect 793 -2481 794 -2480
rect 800 -2481 801 -2480
rect 828 -2481 829 -2480
rect 1381 -2481 1382 -2480
rect 1507 -2481 1508 -2480
rect 1535 -2481 1536 -2480
rect 1640 -2481 1641 -2480
rect 1654 -2481 1655 -2480
rect 173 -2483 174 -2482
rect 296 -2483 297 -2482
rect 366 -2483 367 -2482
rect 562 -2483 563 -2482
rect 618 -2483 619 -2482
rect 919 -2483 920 -2482
rect 947 -2483 948 -2482
rect 1094 -2483 1095 -2482
rect 1178 -2483 1179 -2482
rect 1269 -2483 1270 -2482
rect 1276 -2483 1277 -2482
rect 1591 -2483 1592 -2482
rect 366 -2485 367 -2484
rect 499 -2485 500 -2484
rect 618 -2485 619 -2484
rect 625 -2485 626 -2484
rect 639 -2485 640 -2484
rect 838 -2485 839 -2484
rect 891 -2485 892 -2484
rect 1276 -2485 1277 -2484
rect 1283 -2485 1284 -2484
rect 1332 -2485 1333 -2484
rect 1535 -2485 1536 -2484
rect 1556 -2485 1557 -2484
rect 401 -2487 402 -2486
rect 436 -2487 437 -2486
rect 464 -2487 465 -2486
rect 653 -2487 654 -2486
rect 695 -2487 696 -2486
rect 933 -2487 934 -2486
rect 996 -2487 997 -2486
rect 1038 -2487 1039 -2486
rect 1045 -2487 1046 -2486
rect 1087 -2487 1088 -2486
rect 1129 -2487 1130 -2486
rect 1178 -2487 1179 -2486
rect 1220 -2487 1221 -2486
rect 1237 -2487 1238 -2486
rect 1304 -2487 1305 -2486
rect 1353 -2487 1354 -2486
rect 1556 -2487 1557 -2486
rect 1598 -2487 1599 -2486
rect 128 -2489 129 -2488
rect 996 -2489 997 -2488
rect 1052 -2489 1053 -2488
rect 1150 -2489 1151 -2488
rect 1304 -2489 1305 -2488
rect 1311 -2489 1312 -2488
rect 1458 -2489 1459 -2488
rect 1598 -2489 1599 -2488
rect 408 -2491 409 -2490
rect 443 -2491 444 -2490
rect 485 -2491 486 -2490
rect 604 -2491 605 -2490
rect 621 -2491 622 -2490
rect 688 -2491 689 -2490
rect 702 -2491 703 -2490
rect 807 -2491 808 -2490
rect 870 -2491 871 -2490
rect 891 -2491 892 -2490
rect 926 -2491 927 -2490
rect 1094 -2491 1095 -2490
rect 1146 -2491 1147 -2490
rect 1458 -2491 1459 -2490
rect 65 -2493 66 -2492
rect 485 -2493 486 -2492
rect 499 -2493 500 -2492
rect 541 -2493 542 -2492
rect 569 -2493 570 -2492
rect 1129 -2493 1130 -2492
rect 1255 -2493 1256 -2492
rect 1311 -2493 1312 -2492
rect 65 -2495 66 -2494
rect 1619 -2495 1620 -2494
rect 310 -2497 311 -2496
rect 408 -2497 409 -2496
rect 436 -2497 437 -2496
rect 450 -2497 451 -2496
rect 513 -2497 514 -2496
rect 695 -2497 696 -2496
rect 737 -2497 738 -2496
rect 1612 -2497 1613 -2496
rect 198 -2499 199 -2498
rect 310 -2499 311 -2498
rect 352 -2499 353 -2498
rect 541 -2499 542 -2498
rect 611 -2499 612 -2498
rect 1255 -2499 1256 -2498
rect 89 -2501 90 -2500
rect 352 -2501 353 -2500
rect 450 -2501 451 -2500
rect 565 -2501 566 -2500
rect 625 -2501 626 -2500
rect 912 -2501 913 -2500
rect 1052 -2501 1053 -2500
rect 1080 -2501 1081 -2500
rect 198 -2503 199 -2502
rect 205 -2503 206 -2502
rect 492 -2503 493 -2502
rect 513 -2503 514 -2502
rect 527 -2503 528 -2502
rect 1283 -2503 1284 -2502
rect 205 -2505 206 -2504
rect 212 -2505 213 -2504
rect 345 -2505 346 -2504
rect 527 -2505 528 -2504
rect 548 -2505 549 -2504
rect 611 -2505 612 -2504
rect 649 -2505 650 -2504
rect 1374 -2505 1375 -2504
rect 212 -2507 213 -2506
rect 275 -2507 276 -2506
rect 289 -2507 290 -2506
rect 345 -2507 346 -2506
rect 492 -2507 493 -2506
rect 786 -2507 787 -2506
rect 800 -2507 801 -2506
rect 1451 -2507 1452 -2506
rect 240 -2509 241 -2508
rect 289 -2509 290 -2508
rect 548 -2509 549 -2508
rect 597 -2509 598 -2508
rect 653 -2509 654 -2508
rect 779 -2509 780 -2508
rect 807 -2509 808 -2508
rect 1542 -2509 1543 -2508
rect 275 -2511 276 -2510
rect 422 -2511 423 -2510
rect 506 -2511 507 -2510
rect 597 -2511 598 -2510
rect 744 -2511 745 -2510
rect 1087 -2511 1088 -2510
rect 1367 -2511 1368 -2510
rect 1451 -2511 1452 -2510
rect 1521 -2511 1522 -2510
rect 1542 -2511 1543 -2510
rect 86 -2513 87 -2512
rect 506 -2513 507 -2512
rect 565 -2513 566 -2512
rect 632 -2513 633 -2512
rect 765 -2513 766 -2512
rect 1647 -2513 1648 -2512
rect 86 -2515 87 -2514
rect 520 -2515 521 -2514
rect 779 -2515 780 -2514
rect 1363 -2515 1364 -2514
rect 1479 -2515 1480 -2514
rect 1521 -2515 1522 -2514
rect 156 -2517 157 -2516
rect 422 -2517 423 -2516
rect 814 -2517 815 -2516
rect 870 -2517 871 -2516
rect 884 -2517 885 -2516
rect 926 -2517 927 -2516
rect 1010 -2517 1011 -2516
rect 1080 -2517 1081 -2516
rect 1157 -2517 1158 -2516
rect 1367 -2517 1368 -2516
rect 1472 -2517 1473 -2516
rect 1479 -2517 1480 -2516
rect 100 -2519 101 -2518
rect 156 -2519 157 -2518
rect 268 -2519 269 -2518
rect 814 -2519 815 -2518
rect 884 -2519 885 -2518
rect 1003 -2519 1004 -2518
rect 1073 -2519 1074 -2518
rect 1164 -2519 1165 -2518
rect 1465 -2519 1466 -2518
rect 1472 -2519 1473 -2518
rect 100 -2521 101 -2520
rect 331 -2521 332 -2520
rect 534 -2521 535 -2520
rect 1010 -2521 1011 -2520
rect 1073 -2521 1074 -2520
rect 1136 -2521 1137 -2520
rect 1430 -2521 1431 -2520
rect 1465 -2521 1466 -2520
rect 72 -2523 73 -2522
rect 534 -2523 535 -2522
rect 786 -2523 787 -2522
rect 1157 -2523 1158 -2522
rect 1423 -2523 1424 -2522
rect 1430 -2523 1431 -2522
rect 72 -2525 73 -2524
rect 261 -2525 262 -2524
rect 331 -2525 332 -2524
rect 415 -2525 416 -2524
rect 912 -2525 913 -2524
rect 954 -2525 955 -2524
rect 968 -2525 969 -2524
rect 1003 -2525 1004 -2524
rect 1388 -2525 1389 -2524
rect 1423 -2525 1424 -2524
rect 149 -2527 150 -2526
rect 1136 -2527 1137 -2526
rect 149 -2529 150 -2528
rect 191 -2529 192 -2528
rect 261 -2529 262 -2528
rect 317 -2529 318 -2528
rect 555 -2529 556 -2528
rect 1388 -2529 1389 -2528
rect 184 -2531 185 -2530
rect 268 -2531 269 -2530
rect 278 -2531 279 -2530
rect 555 -2531 556 -2530
rect 751 -2531 752 -2530
rect 954 -2531 955 -2530
rect 968 -2531 969 -2530
rect 982 -2531 983 -2530
rect 177 -2533 178 -2532
rect 184 -2533 185 -2532
rect 191 -2533 192 -2532
rect 744 -2533 745 -2532
rect 982 -2533 983 -2532
rect 1017 -2533 1018 -2532
rect 177 -2535 178 -2534
rect 215 -2535 216 -2534
rect 317 -2535 318 -2534
rect 387 -2535 388 -2534
rect 1017 -2535 1018 -2534
rect 1059 -2535 1060 -2534
rect 1031 -2537 1032 -2536
rect 1059 -2537 1060 -2536
rect 971 -2539 972 -2538
rect 1031 -2539 1032 -2538
rect 44 -2550 45 -2549
rect 303 -2550 304 -2549
rect 387 -2550 388 -2549
rect 639 -2550 640 -2549
rect 656 -2550 657 -2549
rect 1549 -2550 1550 -2549
rect 1556 -2550 1557 -2549
rect 1559 -2550 1560 -2549
rect 1584 -2550 1585 -2549
rect 1605 -2550 1606 -2549
rect 1629 -2550 1630 -2549
rect 1640 -2550 1641 -2549
rect 72 -2552 73 -2551
rect 292 -2552 293 -2551
rect 303 -2552 304 -2551
rect 425 -2552 426 -2551
rect 457 -2552 458 -2551
rect 478 -2552 479 -2551
rect 527 -2552 528 -2551
rect 681 -2552 682 -2551
rect 730 -2552 731 -2551
rect 1465 -2552 1466 -2551
rect 1472 -2552 1473 -2551
rect 1549 -2552 1550 -2551
rect 1556 -2552 1557 -2551
rect 1612 -2552 1613 -2551
rect 72 -2554 73 -2553
rect 618 -2554 619 -2553
rect 625 -2554 626 -2553
rect 807 -2554 808 -2553
rect 849 -2554 850 -2553
rect 898 -2554 899 -2553
rect 950 -2554 951 -2553
rect 1479 -2554 1480 -2553
rect 1514 -2554 1515 -2553
rect 1584 -2554 1585 -2553
rect 1591 -2554 1592 -2553
rect 1619 -2554 1620 -2553
rect 86 -2556 87 -2555
rect 180 -2556 181 -2555
rect 212 -2556 213 -2555
rect 296 -2556 297 -2555
rect 352 -2556 353 -2555
rect 681 -2556 682 -2555
rect 737 -2556 738 -2555
rect 1486 -2556 1487 -2555
rect 1559 -2556 1560 -2555
rect 1612 -2556 1613 -2555
rect 86 -2558 87 -2557
rect 646 -2558 647 -2557
rect 737 -2558 738 -2557
rect 901 -2558 902 -2557
rect 971 -2558 972 -2557
rect 1122 -2558 1123 -2557
rect 1143 -2558 1144 -2557
rect 1325 -2558 1326 -2557
rect 1405 -2558 1406 -2557
rect 1542 -2558 1543 -2557
rect 1598 -2558 1599 -2557
rect 1626 -2558 1627 -2557
rect 93 -2560 94 -2559
rect 212 -2560 213 -2559
rect 233 -2560 234 -2559
rect 667 -2560 668 -2559
rect 744 -2560 745 -2559
rect 1101 -2560 1102 -2559
rect 1136 -2560 1137 -2559
rect 1143 -2560 1144 -2559
rect 1188 -2560 1189 -2559
rect 1430 -2560 1431 -2559
rect 1444 -2560 1445 -2559
rect 1479 -2560 1480 -2559
rect 1507 -2560 1508 -2559
rect 1542 -2560 1543 -2559
rect 1577 -2560 1578 -2559
rect 1598 -2560 1599 -2559
rect 93 -2562 94 -2561
rect 530 -2562 531 -2561
rect 534 -2562 535 -2561
rect 747 -2562 748 -2561
rect 789 -2562 790 -2561
rect 1276 -2562 1277 -2561
rect 1304 -2562 1305 -2561
rect 1402 -2562 1403 -2561
rect 1409 -2562 1410 -2561
rect 1486 -2562 1487 -2561
rect 121 -2564 122 -2563
rect 831 -2564 832 -2563
rect 835 -2564 836 -2563
rect 849 -2564 850 -2563
rect 887 -2564 888 -2563
rect 1297 -2564 1298 -2563
rect 1304 -2564 1305 -2563
rect 1437 -2564 1438 -2563
rect 1458 -2564 1459 -2563
rect 1514 -2564 1515 -2563
rect 65 -2566 66 -2565
rect 121 -2566 122 -2565
rect 135 -2566 136 -2565
rect 828 -2566 829 -2565
rect 901 -2566 902 -2565
rect 1066 -2566 1067 -2565
rect 1073 -2566 1074 -2565
rect 1465 -2566 1466 -2565
rect 65 -2568 66 -2567
rect 100 -2568 101 -2567
rect 135 -2568 136 -2567
rect 177 -2568 178 -2567
rect 201 -2568 202 -2567
rect 1444 -2568 1445 -2567
rect 100 -2570 101 -2569
rect 107 -2570 108 -2569
rect 142 -2570 143 -2569
rect 415 -2570 416 -2569
rect 422 -2570 423 -2569
rect 646 -2570 647 -2569
rect 667 -2570 668 -2569
rect 716 -2570 717 -2569
rect 730 -2570 731 -2569
rect 744 -2570 745 -2569
rect 758 -2570 759 -2569
rect 835 -2570 836 -2569
rect 954 -2570 955 -2569
rect 1325 -2570 1326 -2569
rect 1388 -2570 1389 -2569
rect 1437 -2570 1438 -2569
rect 107 -2572 108 -2571
rect 131 -2572 132 -2571
rect 142 -2572 143 -2571
rect 205 -2572 206 -2571
rect 215 -2572 216 -2571
rect 422 -2572 423 -2571
rect 450 -2572 451 -2571
rect 1122 -2572 1123 -2571
rect 1129 -2572 1130 -2571
rect 1136 -2572 1137 -2571
rect 1234 -2572 1235 -2571
rect 1591 -2572 1592 -2571
rect 152 -2574 153 -2573
rect 1507 -2574 1508 -2573
rect 163 -2576 164 -2575
rect 236 -2576 237 -2575
rect 254 -2576 255 -2575
rect 961 -2576 962 -2575
rect 978 -2576 979 -2575
rect 1283 -2576 1284 -2575
rect 1346 -2576 1347 -2575
rect 1388 -2576 1389 -2575
rect 1409 -2576 1410 -2575
rect 1570 -2576 1571 -2575
rect 226 -2578 227 -2577
rect 254 -2578 255 -2577
rect 275 -2578 276 -2577
rect 758 -2578 759 -2577
rect 803 -2578 804 -2577
rect 1360 -2578 1361 -2577
rect 1423 -2578 1424 -2577
rect 1458 -2578 1459 -2577
rect 198 -2580 199 -2579
rect 226 -2580 227 -2579
rect 268 -2580 269 -2579
rect 275 -2580 276 -2579
rect 278 -2580 279 -2579
rect 688 -2580 689 -2579
rect 828 -2580 829 -2579
rect 877 -2580 878 -2579
rect 926 -2580 927 -2579
rect 954 -2580 955 -2579
rect 961 -2580 962 -2579
rect 1059 -2580 1060 -2579
rect 1066 -2580 1067 -2579
rect 1087 -2580 1088 -2579
rect 1090 -2580 1091 -2579
rect 1535 -2580 1536 -2579
rect 268 -2582 269 -2581
rect 376 -2582 377 -2581
rect 380 -2582 381 -2581
rect 534 -2582 535 -2581
rect 562 -2582 563 -2581
rect 590 -2582 591 -2581
rect 597 -2582 598 -2581
rect 1577 -2582 1578 -2581
rect 247 -2584 248 -2583
rect 590 -2584 591 -2583
rect 600 -2584 601 -2583
rect 1472 -2584 1473 -2583
rect 247 -2586 248 -2585
rect 310 -2586 311 -2585
rect 317 -2586 318 -2585
rect 352 -2586 353 -2585
rect 390 -2586 391 -2585
rect 408 -2586 409 -2585
rect 450 -2586 451 -2585
rect 957 -2586 958 -2585
rect 996 -2586 997 -2585
rect 1563 -2586 1564 -2585
rect 89 -2588 90 -2587
rect 1563 -2588 1564 -2587
rect 191 -2590 192 -2589
rect 310 -2590 311 -2589
rect 345 -2590 346 -2589
rect 380 -2590 381 -2589
rect 394 -2590 395 -2589
rect 415 -2590 416 -2589
rect 457 -2590 458 -2589
rect 485 -2590 486 -2589
rect 492 -2590 493 -2589
rect 618 -2590 619 -2589
rect 625 -2590 626 -2589
rect 709 -2590 710 -2589
rect 880 -2590 881 -2589
rect 996 -2590 997 -2589
rect 1017 -2590 1018 -2589
rect 1297 -2590 1298 -2589
rect 1318 -2590 1319 -2589
rect 1360 -2590 1361 -2589
rect 1374 -2590 1375 -2589
rect 1423 -2590 1424 -2589
rect 58 -2592 59 -2591
rect 191 -2592 192 -2591
rect 282 -2592 283 -2591
rect 443 -2592 444 -2591
rect 464 -2592 465 -2591
rect 562 -2592 563 -2591
rect 565 -2592 566 -2591
rect 1535 -2592 1536 -2591
rect 58 -2594 59 -2593
rect 324 -2594 325 -2593
rect 345 -2594 346 -2593
rect 373 -2594 374 -2593
rect 401 -2594 402 -2593
rect 408 -2594 409 -2593
rect 464 -2594 465 -2593
rect 821 -2594 822 -2593
rect 905 -2594 906 -2593
rect 1059 -2594 1060 -2593
rect 1073 -2594 1074 -2593
rect 1227 -2594 1228 -2593
rect 1251 -2594 1252 -2593
rect 1528 -2594 1529 -2593
rect 233 -2596 234 -2595
rect 324 -2596 325 -2595
rect 401 -2596 402 -2595
rect 541 -2596 542 -2595
rect 555 -2596 556 -2595
rect 709 -2596 710 -2595
rect 786 -2596 787 -2595
rect 1017 -2596 1018 -2595
rect 1024 -2596 1025 -2595
rect 1521 -2596 1522 -2595
rect 257 -2598 258 -2597
rect 443 -2598 444 -2597
rect 481 -2598 482 -2597
rect 492 -2598 493 -2597
rect 502 -2598 503 -2597
rect 597 -2598 598 -2597
rect 611 -2598 612 -2597
rect 639 -2598 640 -2597
rect 688 -2598 689 -2597
rect 814 -2598 815 -2597
rect 821 -2598 822 -2597
rect 891 -2598 892 -2597
rect 905 -2598 906 -2597
rect 975 -2598 976 -2597
rect 1027 -2598 1028 -2597
rect 1339 -2598 1340 -2597
rect 1493 -2598 1494 -2597
rect 1521 -2598 1522 -2597
rect 156 -2600 157 -2599
rect 611 -2600 612 -2599
rect 614 -2600 615 -2599
rect 1283 -2600 1284 -2599
rect 1339 -2600 1340 -2599
rect 1615 -2600 1616 -2599
rect 156 -2602 157 -2601
rect 205 -2602 206 -2601
rect 261 -2602 262 -2601
rect 282 -2602 283 -2601
rect 289 -2602 290 -2601
rect 317 -2602 318 -2601
rect 485 -2602 486 -2601
rect 674 -2602 675 -2601
rect 786 -2602 787 -2601
rect 793 -2602 794 -2601
rect 814 -2602 815 -2601
rect 842 -2602 843 -2601
rect 877 -2602 878 -2601
rect 891 -2602 892 -2601
rect 912 -2602 913 -2601
rect 926 -2602 927 -2601
rect 1038 -2602 1039 -2601
rect 1101 -2602 1102 -2601
rect 1129 -2602 1130 -2601
rect 1262 -2602 1263 -2601
rect 1269 -2602 1270 -2601
rect 1318 -2602 1319 -2601
rect 1416 -2602 1417 -2601
rect 1493 -2602 1494 -2601
rect 1500 -2602 1501 -2601
rect 1528 -2602 1529 -2601
rect 163 -2604 164 -2603
rect 975 -2604 976 -2603
rect 1038 -2604 1039 -2603
rect 1115 -2604 1116 -2603
rect 1178 -2604 1179 -2603
rect 1374 -2604 1375 -2603
rect 1451 -2604 1452 -2603
rect 1500 -2604 1501 -2603
rect 240 -2606 241 -2605
rect 842 -2606 843 -2605
rect 912 -2606 913 -2605
rect 933 -2606 934 -2605
rect 1045 -2606 1046 -2605
rect 1430 -2606 1431 -2605
rect 219 -2608 220 -2607
rect 240 -2608 241 -2607
rect 261 -2608 262 -2607
rect 604 -2608 605 -2607
rect 733 -2608 734 -2607
rect 1178 -2608 1179 -2607
rect 1220 -2608 1221 -2607
rect 1262 -2608 1263 -2607
rect 1269 -2608 1270 -2607
rect 1636 -2608 1637 -2607
rect 219 -2610 220 -2609
rect 264 -2610 265 -2609
rect 289 -2610 290 -2609
rect 338 -2610 339 -2609
rect 520 -2610 521 -2609
rect 674 -2610 675 -2609
rect 733 -2610 734 -2609
rect 1241 -2610 1242 -2609
rect 1255 -2610 1256 -2609
rect 1346 -2610 1347 -2609
rect 1367 -2610 1368 -2609
rect 1416 -2610 1417 -2609
rect 338 -2612 339 -2611
rect 499 -2612 500 -2611
rect 520 -2612 521 -2611
rect 544 -2612 545 -2611
rect 555 -2612 556 -2611
rect 569 -2612 570 -2611
rect 572 -2612 573 -2611
rect 660 -2612 661 -2611
rect 793 -2612 794 -2611
rect 1010 -2612 1011 -2611
rect 1052 -2612 1053 -2611
rect 1146 -2612 1147 -2611
rect 1171 -2612 1172 -2611
rect 1220 -2612 1221 -2611
rect 1227 -2612 1228 -2611
rect 1248 -2612 1249 -2611
rect 1276 -2612 1277 -2611
rect 1587 -2612 1588 -2611
rect 499 -2614 500 -2613
rect 541 -2614 542 -2613
rect 569 -2614 570 -2613
rect 723 -2614 724 -2613
rect 800 -2614 801 -2613
rect 1045 -2614 1046 -2613
rect 1087 -2614 1088 -2613
rect 1234 -2614 1235 -2613
rect 1241 -2614 1242 -2613
rect 1381 -2614 1382 -2613
rect 1395 -2614 1396 -2613
rect 1451 -2614 1452 -2613
rect 471 -2616 472 -2615
rect 723 -2616 724 -2615
rect 863 -2616 864 -2615
rect 1248 -2616 1249 -2615
rect 1332 -2616 1333 -2615
rect 1367 -2616 1368 -2615
rect 359 -2618 360 -2617
rect 471 -2618 472 -2617
rect 583 -2618 584 -2617
rect 754 -2618 755 -2617
rect 863 -2618 864 -2617
rect 870 -2618 871 -2617
rect 884 -2618 885 -2617
rect 933 -2618 934 -2617
rect 940 -2618 941 -2617
rect 1010 -2618 1011 -2617
rect 1031 -2618 1032 -2617
rect 1052 -2618 1053 -2617
rect 1108 -2618 1109 -2617
rect 1171 -2618 1172 -2617
rect 1213 -2618 1214 -2617
rect 1255 -2618 1256 -2617
rect 1290 -2618 1291 -2617
rect 1332 -2618 1333 -2617
rect 1353 -2618 1354 -2617
rect 1395 -2618 1396 -2617
rect 208 -2620 209 -2619
rect 1108 -2620 1109 -2619
rect 1115 -2620 1116 -2619
rect 1199 -2620 1200 -2619
rect 1311 -2620 1312 -2619
rect 1353 -2620 1354 -2619
rect 359 -2622 360 -2621
rect 418 -2622 419 -2621
rect 583 -2622 584 -2621
rect 653 -2622 654 -2621
rect 660 -2622 661 -2621
rect 947 -2622 948 -2621
rect 1031 -2622 1032 -2621
rect 1206 -2622 1207 -2621
rect 331 -2624 332 -2623
rect 653 -2624 654 -2623
rect 670 -2624 671 -2623
rect 1381 -2624 1382 -2623
rect 79 -2626 80 -2625
rect 331 -2626 332 -2625
rect 604 -2626 605 -2625
rect 702 -2626 703 -2625
rect 740 -2626 741 -2625
rect 1206 -2626 1207 -2625
rect 79 -2628 80 -2627
rect 128 -2628 129 -2627
rect 702 -2628 703 -2627
rect 989 -2628 990 -2627
rect 1080 -2628 1081 -2627
rect 1213 -2628 1214 -2627
rect 803 -2630 804 -2629
rect 1290 -2630 1291 -2629
rect 810 -2632 811 -2631
rect 947 -2632 948 -2631
rect 989 -2632 990 -2631
rect 1003 -2632 1004 -2631
rect 1164 -2632 1165 -2631
rect 1199 -2632 1200 -2631
rect 856 -2634 857 -2633
rect 870 -2634 871 -2633
rect 884 -2634 885 -2633
rect 1094 -2634 1095 -2633
rect 1157 -2634 1158 -2633
rect 1164 -2634 1165 -2633
rect 1192 -2634 1193 -2633
rect 1311 -2634 1312 -2633
rect 170 -2636 171 -2635
rect 1094 -2636 1095 -2635
rect 1150 -2636 1151 -2635
rect 1157 -2636 1158 -2635
rect 170 -2638 171 -2637
rect 184 -2638 185 -2637
rect 751 -2638 752 -2637
rect 1192 -2638 1193 -2637
rect 184 -2640 185 -2639
rect 719 -2640 720 -2639
rect 859 -2640 860 -2639
rect 1080 -2640 1081 -2639
rect 1150 -2640 1151 -2639
rect 1605 -2640 1606 -2639
rect 506 -2642 507 -2641
rect 751 -2642 752 -2641
rect 919 -2642 920 -2641
rect 940 -2642 941 -2641
rect 982 -2642 983 -2641
rect 1003 -2642 1004 -2641
rect 506 -2644 507 -2643
rect 548 -2644 549 -2643
rect 919 -2644 920 -2643
rect 1153 -2644 1154 -2643
rect 436 -2646 437 -2645
rect 548 -2646 549 -2645
rect 968 -2646 969 -2645
rect 982 -2646 983 -2645
rect 436 -2648 437 -2647
rect 513 -2648 514 -2647
rect 968 -2648 969 -2647
rect 1185 -2648 1186 -2647
rect 513 -2650 514 -2649
rect 576 -2650 577 -2649
rect 1185 -2650 1186 -2649
rect 1570 -2650 1571 -2649
rect 576 -2652 577 -2651
rect 765 -2652 766 -2651
rect 765 -2654 766 -2653
rect 772 -2654 773 -2653
rect 695 -2656 696 -2655
rect 772 -2656 773 -2655
rect 695 -2658 696 -2657
rect 779 -2658 780 -2657
rect 51 -2660 52 -2659
rect 779 -2660 780 -2659
rect 51 -2662 52 -2661
rect 149 -2662 150 -2661
rect 114 -2664 115 -2663
rect 149 -2664 150 -2663
rect 114 -2666 115 -2665
rect 366 -2666 367 -2665
rect 366 -2668 367 -2667
rect 898 -2668 899 -2667
rect 44 -2679 45 -2678
rect 747 -2679 748 -2678
rect 782 -2679 783 -2678
rect 1584 -2679 1585 -2678
rect 44 -2681 45 -2680
rect 394 -2681 395 -2680
rect 397 -2681 398 -2680
rect 429 -2681 430 -2680
rect 436 -2681 437 -2680
rect 499 -2681 500 -2680
rect 534 -2681 535 -2680
rect 646 -2681 647 -2680
rect 649 -2681 650 -2680
rect 772 -2681 773 -2680
rect 786 -2681 787 -2680
rect 884 -2681 885 -2680
rect 908 -2681 909 -2680
rect 1297 -2681 1298 -2680
rect 1524 -2681 1525 -2680
rect 1598 -2681 1599 -2680
rect 51 -2683 52 -2682
rect 201 -2683 202 -2682
rect 205 -2683 206 -2682
rect 345 -2683 346 -2682
rect 394 -2683 395 -2682
rect 1188 -2683 1189 -2682
rect 1262 -2683 1263 -2682
rect 1300 -2683 1301 -2682
rect 58 -2685 59 -2684
rect 236 -2685 237 -2684
rect 264 -2685 265 -2684
rect 1283 -2685 1284 -2684
rect 58 -2687 59 -2686
rect 128 -2687 129 -2686
rect 135 -2687 136 -2686
rect 177 -2687 178 -2686
rect 198 -2687 199 -2686
rect 310 -2687 311 -2686
rect 331 -2687 332 -2686
rect 429 -2687 430 -2686
rect 446 -2687 447 -2686
rect 1507 -2687 1508 -2686
rect 72 -2689 73 -2688
rect 677 -2689 678 -2688
rect 681 -2689 682 -2688
rect 772 -2689 773 -2688
rect 786 -2689 787 -2688
rect 1465 -2689 1466 -2688
rect 1507 -2689 1508 -2688
rect 1605 -2689 1606 -2688
rect 72 -2691 73 -2690
rect 170 -2691 171 -2690
rect 177 -2691 178 -2690
rect 443 -2691 444 -2690
rect 499 -2691 500 -2690
rect 793 -2691 794 -2690
rect 800 -2691 801 -2690
rect 1171 -2691 1172 -2690
rect 1185 -2691 1186 -2690
rect 1549 -2691 1550 -2690
rect 79 -2693 80 -2692
rect 373 -2693 374 -2692
rect 408 -2693 409 -2692
rect 422 -2693 423 -2692
rect 534 -2693 535 -2692
rect 807 -2693 808 -2692
rect 817 -2693 818 -2692
rect 1486 -2693 1487 -2692
rect 79 -2695 80 -2694
rect 765 -2695 766 -2694
rect 793 -2695 794 -2694
rect 814 -2695 815 -2694
rect 877 -2695 878 -2694
rect 1010 -2695 1011 -2694
rect 1024 -2695 1025 -2694
rect 1465 -2695 1466 -2694
rect 1486 -2695 1487 -2694
rect 1577 -2695 1578 -2694
rect 86 -2697 87 -2696
rect 565 -2697 566 -2696
rect 576 -2697 577 -2696
rect 716 -2697 717 -2696
rect 730 -2697 731 -2696
rect 1153 -2697 1154 -2696
rect 1185 -2697 1186 -2696
rect 1339 -2697 1340 -2696
rect 86 -2699 87 -2698
rect 100 -2699 101 -2698
rect 114 -2699 115 -2698
rect 331 -2699 332 -2698
rect 345 -2699 346 -2698
rect 352 -2699 353 -2698
rect 373 -2699 374 -2698
rect 415 -2699 416 -2698
rect 422 -2699 423 -2698
rect 541 -2699 542 -2698
rect 576 -2699 577 -2698
rect 695 -2699 696 -2698
rect 709 -2699 710 -2698
rect 733 -2699 734 -2698
rect 737 -2699 738 -2698
rect 898 -2699 899 -2698
rect 940 -2699 941 -2698
rect 950 -2699 951 -2698
rect 957 -2699 958 -2698
rect 1311 -2699 1312 -2698
rect 65 -2701 66 -2700
rect 114 -2701 115 -2700
rect 124 -2701 125 -2700
rect 198 -2701 199 -2700
rect 205 -2701 206 -2700
rect 240 -2701 241 -2700
rect 264 -2701 265 -2700
rect 296 -2701 297 -2700
rect 310 -2701 311 -2700
rect 611 -2701 612 -2700
rect 653 -2701 654 -2700
rect 800 -2701 801 -2700
rect 845 -2701 846 -2700
rect 898 -2701 899 -2700
rect 933 -2701 934 -2700
rect 940 -2701 941 -2700
rect 968 -2701 969 -2700
rect 996 -2701 997 -2700
rect 1010 -2701 1011 -2700
rect 1626 -2701 1627 -2700
rect 65 -2703 66 -2702
rect 152 -2703 153 -2702
rect 156 -2703 157 -2702
rect 618 -2703 619 -2702
rect 653 -2703 654 -2702
rect 1143 -2703 1144 -2702
rect 1150 -2703 1151 -2702
rect 1612 -2703 1613 -2702
rect 93 -2705 94 -2704
rect 159 -2705 160 -2704
rect 170 -2705 171 -2704
rect 450 -2705 451 -2704
rect 464 -2705 465 -2704
rect 541 -2705 542 -2704
rect 569 -2705 570 -2704
rect 618 -2705 619 -2704
rect 656 -2705 657 -2704
rect 1052 -2705 1053 -2704
rect 1073 -2705 1074 -2704
rect 1171 -2705 1172 -2704
rect 1241 -2705 1242 -2704
rect 1339 -2705 1340 -2704
rect 93 -2707 94 -2706
rect 247 -2707 248 -2706
rect 296 -2707 297 -2706
rect 471 -2707 472 -2706
rect 520 -2707 521 -2706
rect 877 -2707 878 -2706
rect 880 -2707 881 -2706
rect 1374 -2707 1375 -2706
rect 100 -2709 101 -2708
rect 208 -2709 209 -2708
rect 212 -2709 213 -2708
rect 247 -2709 248 -2708
rect 352 -2709 353 -2708
rect 401 -2709 402 -2708
rect 415 -2709 416 -2708
rect 555 -2709 556 -2708
rect 569 -2709 570 -2708
rect 590 -2709 591 -2708
rect 604 -2709 605 -2708
rect 737 -2709 738 -2708
rect 744 -2709 745 -2708
rect 761 -2709 762 -2708
rect 765 -2709 766 -2708
rect 821 -2709 822 -2708
rect 880 -2709 881 -2708
rect 1101 -2709 1102 -2708
rect 1150 -2709 1151 -2708
rect 1381 -2709 1382 -2708
rect 128 -2711 129 -2710
rect 436 -2711 437 -2710
rect 450 -2711 451 -2710
rect 506 -2711 507 -2710
rect 555 -2711 556 -2710
rect 723 -2711 724 -2710
rect 744 -2711 745 -2710
rect 1430 -2711 1431 -2710
rect 135 -2713 136 -2712
rect 639 -2713 640 -2712
rect 660 -2713 661 -2712
rect 1090 -2713 1091 -2712
rect 1101 -2713 1102 -2712
rect 1206 -2713 1207 -2712
rect 1241 -2713 1242 -2712
rect 1353 -2713 1354 -2712
rect 1381 -2713 1382 -2712
rect 1542 -2713 1543 -2712
rect 142 -2715 143 -2714
rect 261 -2715 262 -2714
rect 401 -2715 402 -2714
rect 492 -2715 493 -2714
rect 506 -2715 507 -2714
rect 667 -2715 668 -2714
rect 674 -2715 675 -2714
rect 814 -2715 815 -2714
rect 821 -2715 822 -2714
rect 849 -2715 850 -2714
rect 884 -2715 885 -2714
rect 947 -2715 948 -2714
rect 954 -2715 955 -2714
rect 1143 -2715 1144 -2714
rect 1188 -2715 1189 -2714
rect 1374 -2715 1375 -2714
rect 1430 -2715 1431 -2714
rect 1514 -2715 1515 -2714
rect 142 -2717 143 -2716
rect 289 -2717 290 -2716
rect 425 -2717 426 -2716
rect 604 -2717 605 -2716
rect 611 -2717 612 -2716
rect 919 -2717 920 -2716
rect 926 -2717 927 -2716
rect 1052 -2717 1053 -2716
rect 1087 -2717 1088 -2716
rect 1178 -2717 1179 -2716
rect 1262 -2717 1263 -2716
rect 1367 -2717 1368 -2716
rect 1514 -2717 1515 -2716
rect 1619 -2717 1620 -2716
rect 149 -2719 150 -2718
rect 856 -2719 857 -2718
rect 870 -2719 871 -2718
rect 919 -2719 920 -2718
rect 933 -2719 934 -2718
rect 982 -2719 983 -2718
rect 996 -2719 997 -2718
rect 1003 -2719 1004 -2718
rect 1024 -2719 1025 -2718
rect 1108 -2719 1109 -2718
rect 1129 -2719 1130 -2718
rect 1206 -2719 1207 -2718
rect 1283 -2719 1284 -2718
rect 1451 -2719 1452 -2718
rect 149 -2721 150 -2720
rect 268 -2721 269 -2720
rect 464 -2721 465 -2720
rect 597 -2721 598 -2720
rect 625 -2721 626 -2720
rect 723 -2721 724 -2720
rect 779 -2721 780 -2720
rect 1073 -2721 1074 -2720
rect 1108 -2721 1109 -2720
rect 1192 -2721 1193 -2720
rect 1311 -2721 1312 -2720
rect 1395 -2721 1396 -2720
rect 1451 -2721 1452 -2720
rect 1528 -2721 1529 -2720
rect 156 -2723 157 -2722
rect 1269 -2723 1270 -2722
rect 1353 -2723 1354 -2722
rect 1444 -2723 1445 -2722
rect 163 -2725 164 -2724
rect 268 -2725 269 -2724
rect 387 -2725 388 -2724
rect 597 -2725 598 -2724
rect 660 -2725 661 -2724
rect 1591 -2725 1592 -2724
rect 163 -2727 164 -2726
rect 219 -2727 220 -2726
rect 226 -2727 227 -2726
rect 240 -2727 241 -2726
rect 387 -2727 388 -2726
rect 548 -2727 549 -2726
rect 562 -2727 563 -2726
rect 639 -2727 640 -2726
rect 663 -2727 664 -2726
rect 870 -2727 871 -2726
rect 901 -2727 902 -2726
rect 1269 -2727 1270 -2726
rect 1367 -2727 1368 -2726
rect 1458 -2727 1459 -2726
rect 138 -2729 139 -2728
rect 1458 -2729 1459 -2728
rect 215 -2731 216 -2730
rect 254 -2731 255 -2730
rect 408 -2731 409 -2730
rect 562 -2731 563 -2730
rect 681 -2731 682 -2730
rect 751 -2731 752 -2730
rect 849 -2731 850 -2730
rect 989 -2731 990 -2730
rect 1115 -2731 1116 -2730
rect 1129 -2731 1130 -2730
rect 1192 -2731 1193 -2730
rect 1423 -2731 1424 -2730
rect 1444 -2731 1445 -2730
rect 1629 -2731 1630 -2730
rect 219 -2733 220 -2732
rect 303 -2733 304 -2732
rect 366 -2733 367 -2732
rect 751 -2733 752 -2732
rect 856 -2733 857 -2732
rect 863 -2733 864 -2732
rect 905 -2733 906 -2732
rect 1178 -2733 1179 -2732
rect 1395 -2733 1396 -2732
rect 1472 -2733 1473 -2732
rect 226 -2735 227 -2734
rect 233 -2735 234 -2734
rect 254 -2735 255 -2734
rect 282 -2735 283 -2734
rect 303 -2735 304 -2734
rect 338 -2735 339 -2734
rect 471 -2735 472 -2734
rect 485 -2735 486 -2734
rect 492 -2735 493 -2734
rect 614 -2735 615 -2734
rect 691 -2735 692 -2734
rect 1080 -2735 1081 -2734
rect 1115 -2735 1116 -2734
rect 1227 -2735 1228 -2734
rect 1472 -2735 1473 -2734
rect 1556 -2735 1557 -2734
rect 212 -2737 213 -2736
rect 485 -2737 486 -2736
rect 527 -2737 528 -2736
rect 625 -2737 626 -2736
rect 695 -2737 696 -2736
rect 1094 -2737 1095 -2736
rect 1227 -2737 1228 -2736
rect 1325 -2737 1326 -2736
rect 324 -2739 325 -2738
rect 366 -2739 367 -2738
rect 478 -2739 479 -2738
rect 520 -2739 521 -2738
rect 527 -2739 528 -2738
rect 632 -2739 633 -2738
rect 702 -2739 703 -2738
rect 926 -2739 927 -2738
rect 954 -2739 955 -2738
rect 1136 -2739 1137 -2738
rect 1255 -2739 1256 -2738
rect 1325 -2739 1326 -2738
rect 292 -2741 293 -2740
rect 478 -2741 479 -2740
rect 548 -2741 549 -2740
rect 842 -2741 843 -2740
rect 859 -2741 860 -2740
rect 1423 -2741 1424 -2740
rect 324 -2743 325 -2742
rect 513 -2743 514 -2742
rect 583 -2743 584 -2742
rect 632 -2743 633 -2742
rect 702 -2743 703 -2742
rect 758 -2743 759 -2742
rect 842 -2743 843 -2742
rect 1059 -2743 1060 -2742
rect 1080 -2743 1081 -2742
rect 1157 -2743 1158 -2742
rect 1255 -2743 1256 -2742
rect 1360 -2743 1361 -2742
rect 338 -2745 339 -2744
rect 359 -2745 360 -2744
rect 457 -2745 458 -2744
rect 513 -2745 514 -2744
rect 583 -2745 584 -2744
rect 688 -2745 689 -2744
rect 709 -2745 710 -2744
rect 835 -2745 836 -2744
rect 863 -2745 864 -2744
rect 1157 -2745 1158 -2744
rect 1160 -2745 1161 -2744
rect 1360 -2745 1361 -2744
rect 184 -2747 185 -2746
rect 359 -2747 360 -2746
rect 380 -2747 381 -2746
rect 457 -2747 458 -2746
rect 758 -2747 759 -2746
rect 1346 -2747 1347 -2746
rect 184 -2749 185 -2748
rect 803 -2749 804 -2748
rect 828 -2749 829 -2748
rect 835 -2749 836 -2748
rect 891 -2749 892 -2748
rect 905 -2749 906 -2748
rect 961 -2749 962 -2748
rect 982 -2749 983 -2748
rect 989 -2749 990 -2748
rect 1017 -2749 1018 -2748
rect 1059 -2749 1060 -2748
rect 1220 -2749 1221 -2748
rect 1346 -2749 1347 -2748
rect 1437 -2749 1438 -2748
rect 121 -2751 122 -2750
rect 891 -2751 892 -2750
rect 971 -2751 972 -2750
rect 1038 -2751 1039 -2750
rect 1094 -2751 1095 -2750
rect 1164 -2751 1165 -2750
rect 1220 -2751 1221 -2750
rect 1636 -2751 1637 -2750
rect 121 -2753 122 -2752
rect 131 -2753 132 -2752
rect 317 -2753 318 -2752
rect 380 -2753 381 -2752
rect 779 -2753 780 -2752
rect 961 -2753 962 -2752
rect 975 -2753 976 -2752
rect 1045 -2753 1046 -2752
rect 1136 -2753 1137 -2752
rect 1234 -2753 1235 -2752
rect 1437 -2753 1438 -2752
rect 1521 -2753 1522 -2752
rect 107 -2755 108 -2754
rect 131 -2755 132 -2754
rect 191 -2755 192 -2754
rect 317 -2755 318 -2754
rect 828 -2755 829 -2754
rect 912 -2755 913 -2754
rect 947 -2755 948 -2754
rect 1521 -2755 1522 -2754
rect 107 -2757 108 -2756
rect 191 -2757 192 -2756
rect 289 -2757 290 -2756
rect 975 -2757 976 -2756
rect 978 -2757 979 -2756
rect 1493 -2757 1494 -2756
rect 667 -2759 668 -2758
rect 912 -2759 913 -2758
rect 1017 -2759 1018 -2758
rect 1031 -2759 1032 -2758
rect 1038 -2759 1039 -2758
rect 1122 -2759 1123 -2758
rect 1164 -2759 1165 -2758
rect 1248 -2759 1249 -2758
rect 1493 -2759 1494 -2758
rect 1570 -2759 1571 -2758
rect 1031 -2761 1032 -2760
rect 1066 -2761 1067 -2760
rect 1122 -2761 1123 -2760
rect 1276 -2761 1277 -2760
rect 1045 -2763 1046 -2762
rect 1213 -2763 1214 -2762
rect 1234 -2763 1235 -2762
rect 1332 -2763 1333 -2762
rect 1066 -2765 1067 -2764
rect 1199 -2765 1200 -2764
rect 1213 -2765 1214 -2764
rect 1318 -2765 1319 -2764
rect 1332 -2765 1333 -2764
rect 1409 -2765 1410 -2764
rect 1199 -2767 1200 -2766
rect 1290 -2767 1291 -2766
rect 1318 -2767 1319 -2766
rect 1416 -2767 1417 -2766
rect 887 -2769 888 -2768
rect 1416 -2769 1417 -2768
rect 1248 -2771 1249 -2770
rect 1633 -2771 1634 -2770
rect 1276 -2773 1277 -2772
rect 1388 -2773 1389 -2772
rect 1409 -2773 1410 -2772
rect 1500 -2773 1501 -2772
rect 1290 -2775 1291 -2774
rect 1535 -2775 1536 -2774
rect 1304 -2777 1305 -2776
rect 1388 -2777 1389 -2776
rect 1402 -2777 1403 -2776
rect 1500 -2777 1501 -2776
rect 674 -2779 675 -2778
rect 1304 -2779 1305 -2778
rect 1402 -2779 1403 -2778
rect 1479 -2779 1480 -2778
rect 1479 -2781 1480 -2780
rect 1563 -2781 1564 -2780
rect 58 -2792 59 -2791
rect 236 -2792 237 -2791
rect 247 -2792 248 -2791
rect 292 -2792 293 -2791
rect 303 -2792 304 -2791
rect 558 -2792 559 -2791
rect 593 -2792 594 -2791
rect 730 -2792 731 -2791
rect 747 -2792 748 -2791
rect 1143 -2792 1144 -2791
rect 1160 -2792 1161 -2791
rect 1500 -2792 1501 -2791
rect 65 -2794 66 -2793
rect 138 -2794 139 -2793
rect 149 -2794 150 -2793
rect 282 -2794 283 -2793
rect 285 -2794 286 -2793
rect 366 -2794 367 -2793
rect 380 -2794 381 -2793
rect 446 -2794 447 -2793
rect 499 -2794 500 -2793
rect 789 -2794 790 -2793
rect 810 -2794 811 -2793
rect 1479 -2794 1480 -2793
rect 86 -2796 87 -2795
rect 107 -2796 108 -2795
rect 110 -2796 111 -2795
rect 828 -2796 829 -2795
rect 845 -2796 846 -2795
rect 996 -2796 997 -2795
rect 1006 -2796 1007 -2795
rect 1325 -2796 1326 -2795
rect 86 -2798 87 -2797
rect 317 -2798 318 -2797
rect 324 -2798 325 -2797
rect 705 -2798 706 -2797
rect 730 -2798 731 -2797
rect 737 -2798 738 -2797
rect 772 -2798 773 -2797
rect 922 -2798 923 -2797
rect 996 -2798 997 -2797
rect 1136 -2798 1137 -2797
rect 1297 -2798 1298 -2797
rect 1381 -2798 1382 -2797
rect 93 -2800 94 -2799
rect 838 -2800 839 -2799
rect 866 -2800 867 -2799
rect 1486 -2800 1487 -2799
rect 93 -2802 94 -2801
rect 184 -2802 185 -2801
rect 198 -2802 199 -2801
rect 292 -2802 293 -2801
rect 310 -2802 311 -2801
rect 324 -2802 325 -2801
rect 331 -2802 332 -2801
rect 495 -2802 496 -2801
rect 499 -2802 500 -2801
rect 670 -2802 671 -2801
rect 688 -2802 689 -2801
rect 723 -2802 724 -2801
rect 737 -2802 738 -2801
rect 751 -2802 752 -2801
rect 772 -2802 773 -2801
rect 884 -2802 885 -2801
rect 898 -2802 899 -2801
rect 1185 -2802 1186 -2801
rect 1297 -2802 1298 -2801
rect 1395 -2802 1396 -2801
rect 107 -2804 108 -2803
rect 352 -2804 353 -2803
rect 366 -2804 367 -2803
rect 422 -2804 423 -2803
rect 429 -2804 430 -2803
rect 660 -2804 661 -2803
rect 688 -2804 689 -2803
rect 1150 -2804 1151 -2803
rect 1185 -2804 1186 -2803
rect 1255 -2804 1256 -2803
rect 1325 -2804 1326 -2803
rect 1437 -2804 1438 -2803
rect 100 -2806 101 -2805
rect 429 -2806 430 -2805
rect 443 -2806 444 -2805
rect 908 -2806 909 -2805
rect 912 -2806 913 -2805
rect 1157 -2806 1158 -2805
rect 1255 -2806 1256 -2805
rect 1311 -2806 1312 -2805
rect 1363 -2806 1364 -2805
rect 1395 -2806 1396 -2805
rect 114 -2808 115 -2807
rect 117 -2808 118 -2807
rect 121 -2808 122 -2807
rect 653 -2808 654 -2807
rect 723 -2808 724 -2807
rect 1010 -2808 1011 -2807
rect 1020 -2808 1021 -2807
rect 1507 -2808 1508 -2807
rect 114 -2810 115 -2809
rect 275 -2810 276 -2809
rect 310 -2810 311 -2809
rect 408 -2810 409 -2809
rect 443 -2810 444 -2809
rect 492 -2810 493 -2809
rect 506 -2810 507 -2809
rect 779 -2810 780 -2809
rect 828 -2810 829 -2809
rect 849 -2810 850 -2809
rect 898 -2810 899 -2809
rect 954 -2810 955 -2809
rect 1010 -2810 1011 -2809
rect 1164 -2810 1165 -2809
rect 1311 -2810 1312 -2809
rect 1430 -2810 1431 -2809
rect 117 -2812 118 -2811
rect 275 -2812 276 -2811
rect 338 -2812 339 -2811
rect 422 -2812 423 -2811
rect 506 -2812 507 -2811
rect 625 -2812 626 -2811
rect 653 -2812 654 -2811
rect 1003 -2812 1004 -2811
rect 1097 -2812 1098 -2811
rect 1283 -2812 1284 -2811
rect 1381 -2812 1382 -2811
rect 1521 -2812 1522 -2811
rect 124 -2814 125 -2813
rect 331 -2814 332 -2813
rect 345 -2814 346 -2813
rect 590 -2814 591 -2813
rect 597 -2814 598 -2813
rect 807 -2814 808 -2813
rect 842 -2814 843 -2813
rect 884 -2814 885 -2813
rect 1003 -2814 1004 -2813
rect 1101 -2814 1102 -2813
rect 1129 -2814 1130 -2813
rect 1143 -2814 1144 -2813
rect 1150 -2814 1151 -2813
rect 1269 -2814 1270 -2813
rect 1283 -2814 1284 -2813
rect 1374 -2814 1375 -2813
rect 1430 -2814 1431 -2813
rect 1493 -2814 1494 -2813
rect 44 -2816 45 -2815
rect 124 -2816 125 -2815
rect 128 -2816 129 -2815
rect 513 -2816 514 -2815
rect 520 -2816 521 -2815
rect 562 -2816 563 -2815
rect 565 -2816 566 -2815
rect 1269 -2816 1270 -2815
rect 1374 -2816 1375 -2815
rect 1465 -2816 1466 -2815
rect 103 -2818 104 -2817
rect 128 -2818 129 -2817
rect 135 -2818 136 -2817
rect 660 -2818 661 -2817
rect 744 -2818 745 -2817
rect 1157 -2818 1158 -2817
rect 1164 -2818 1165 -2817
rect 1276 -2818 1277 -2817
rect 135 -2820 136 -2819
rect 569 -2820 570 -2819
rect 590 -2820 591 -2819
rect 604 -2820 605 -2819
rect 625 -2820 626 -2819
rect 947 -2820 948 -2819
rect 1101 -2820 1102 -2819
rect 1262 -2820 1263 -2819
rect 1276 -2820 1277 -2819
rect 1367 -2820 1368 -2819
rect 142 -2822 143 -2821
rect 338 -2822 339 -2821
rect 345 -2822 346 -2821
rect 401 -2822 402 -2821
rect 408 -2822 409 -2821
rect 485 -2822 486 -2821
rect 513 -2822 514 -2821
rect 709 -2822 710 -2821
rect 744 -2822 745 -2821
rect 1094 -2822 1095 -2821
rect 1129 -2822 1130 -2821
rect 1213 -2822 1214 -2821
rect 1262 -2822 1263 -2821
rect 1360 -2822 1361 -2821
rect 1367 -2822 1368 -2821
rect 1458 -2822 1459 -2821
rect 142 -2824 143 -2823
rect 149 -2824 150 -2823
rect 156 -2824 157 -2823
rect 555 -2824 556 -2823
rect 597 -2824 598 -2823
rect 681 -2824 682 -2823
rect 709 -2824 710 -2823
rect 880 -2824 881 -2823
rect 1136 -2824 1137 -2823
rect 1300 -2824 1301 -2823
rect 159 -2826 160 -2825
rect 856 -2826 857 -2825
rect 1213 -2826 1214 -2825
rect 1339 -2826 1340 -2825
rect 170 -2828 171 -2827
rect 303 -2828 304 -2827
rect 317 -2828 318 -2827
rect 1094 -2828 1095 -2827
rect 170 -2830 171 -2829
rect 250 -2830 251 -2829
rect 261 -2830 262 -2829
rect 541 -2830 542 -2829
rect 548 -2830 549 -2829
rect 667 -2830 668 -2829
rect 681 -2830 682 -2829
rect 947 -2830 948 -2829
rect 177 -2832 178 -2831
rect 478 -2832 479 -2831
rect 520 -2832 521 -2831
rect 765 -2832 766 -2831
rect 779 -2832 780 -2831
rect 891 -2832 892 -2831
rect 177 -2834 178 -2833
rect 450 -2834 451 -2833
rect 471 -2834 472 -2833
rect 485 -2834 486 -2833
rect 527 -2834 528 -2833
rect 562 -2834 563 -2833
rect 632 -2834 633 -2833
rect 667 -2834 668 -2833
rect 765 -2834 766 -2833
rect 863 -2834 864 -2833
rect 891 -2834 892 -2833
rect 989 -2834 990 -2833
rect 184 -2836 185 -2835
rect 205 -2836 206 -2835
rect 212 -2836 213 -2835
rect 1290 -2836 1291 -2835
rect 72 -2838 73 -2837
rect 205 -2838 206 -2837
rect 212 -2838 213 -2837
rect 282 -2838 283 -2837
rect 352 -2838 353 -2837
rect 457 -2838 458 -2837
rect 527 -2838 528 -2837
rect 957 -2838 958 -2837
rect 989 -2838 990 -2837
rect 1087 -2838 1088 -2837
rect 72 -2840 73 -2839
rect 163 -2840 164 -2839
rect 191 -2840 192 -2839
rect 198 -2840 199 -2839
rect 215 -2840 216 -2839
rect 677 -2840 678 -2839
rect 800 -2840 801 -2839
rect 807 -2840 808 -2839
rect 842 -2840 843 -2839
rect 982 -2840 983 -2839
rect 163 -2842 164 -2841
rect 268 -2842 269 -2841
rect 380 -2842 381 -2841
rect 642 -2842 643 -2841
rect 663 -2842 664 -2841
rect 1339 -2842 1340 -2841
rect 191 -2844 192 -2843
rect 208 -2844 209 -2843
rect 233 -2844 234 -2843
rect 751 -2844 752 -2843
rect 800 -2844 801 -2843
rect 940 -2844 941 -2843
rect 954 -2844 955 -2843
rect 1087 -2844 1088 -2843
rect 226 -2846 227 -2845
rect 233 -2846 234 -2845
rect 247 -2846 248 -2845
rect 695 -2846 696 -2845
rect 845 -2846 846 -2845
rect 940 -2846 941 -2845
rect 982 -2846 983 -2845
rect 1066 -2846 1067 -2845
rect 226 -2848 227 -2847
rect 618 -2848 619 -2847
rect 632 -2848 633 -2847
rect 1024 -2848 1025 -2847
rect 1066 -2848 1067 -2847
rect 1220 -2848 1221 -2847
rect 254 -2850 255 -2849
rect 268 -2850 269 -2849
rect 387 -2850 388 -2849
rect 814 -2850 815 -2849
rect 849 -2850 850 -2849
rect 1073 -2850 1074 -2849
rect 219 -2852 220 -2851
rect 387 -2852 388 -2851
rect 401 -2852 402 -2851
rect 464 -2852 465 -2851
rect 534 -2852 535 -2851
rect 824 -2852 825 -2851
rect 856 -2852 857 -2851
rect 961 -2852 962 -2851
rect 1073 -2852 1074 -2851
rect 1241 -2852 1242 -2851
rect 219 -2854 220 -2853
rect 817 -2854 818 -2853
rect 912 -2854 913 -2853
rect 1290 -2854 1291 -2853
rect 229 -2856 230 -2855
rect 464 -2856 465 -2855
rect 534 -2856 535 -2855
rect 702 -2856 703 -2855
rect 761 -2856 762 -2855
rect 1220 -2856 1221 -2855
rect 1241 -2856 1242 -2855
rect 1353 -2856 1354 -2855
rect 240 -2858 241 -2857
rect 254 -2858 255 -2857
rect 264 -2858 265 -2857
rect 359 -2858 360 -2857
rect 436 -2858 437 -2857
rect 471 -2858 472 -2857
rect 541 -2858 542 -2857
rect 646 -2858 647 -2857
rect 674 -2858 675 -2857
rect 702 -2858 703 -2857
rect 761 -2858 762 -2857
rect 1052 -2858 1053 -2857
rect 1353 -2858 1354 -2857
rect 1472 -2858 1473 -2857
rect 79 -2860 80 -2859
rect 436 -2860 437 -2859
rect 450 -2860 451 -2859
rect 576 -2860 577 -2859
rect 618 -2860 619 -2859
rect 639 -2860 640 -2859
rect 695 -2860 696 -2859
rect 793 -2860 794 -2859
rect 814 -2860 815 -2859
rect 919 -2860 920 -2859
rect 961 -2860 962 -2859
rect 1045 -2860 1046 -2859
rect 1052 -2860 1053 -2859
rect 1227 -2860 1228 -2859
rect 79 -2862 80 -2861
rect 278 -2862 279 -2861
rect 359 -2862 360 -2861
rect 415 -2862 416 -2861
rect 457 -2862 458 -2861
rect 915 -2862 916 -2861
rect 919 -2862 920 -2861
rect 1122 -2862 1123 -2861
rect 121 -2864 122 -2863
rect 646 -2864 647 -2863
rect 793 -2864 794 -2863
rect 835 -2864 836 -2863
rect 877 -2864 878 -2863
rect 1227 -2864 1228 -2863
rect 240 -2866 241 -2865
rect 870 -2866 871 -2865
rect 1045 -2866 1046 -2865
rect 1199 -2866 1200 -2865
rect 394 -2868 395 -2867
rect 415 -2868 416 -2867
rect 548 -2868 549 -2867
rect 716 -2868 717 -2867
rect 786 -2868 787 -2867
rect 877 -2868 878 -2867
rect 1122 -2868 1123 -2867
rect 1318 -2868 1319 -2867
rect 145 -2870 146 -2869
rect 394 -2870 395 -2869
rect 555 -2870 556 -2869
rect 604 -2870 605 -2869
rect 611 -2870 612 -2869
rect 639 -2870 640 -2869
rect 716 -2870 717 -2869
rect 758 -2870 759 -2869
rect 786 -2870 787 -2869
rect 821 -2870 822 -2869
rect 870 -2870 871 -2869
rect 926 -2870 927 -2869
rect 1192 -2870 1193 -2869
rect 1199 -2870 1200 -2869
rect 1318 -2870 1319 -2869
rect 1388 -2870 1389 -2869
rect 569 -2872 570 -2871
rect 835 -2872 836 -2871
rect 926 -2872 927 -2871
rect 933 -2872 934 -2871
rect 1017 -2872 1018 -2871
rect 1192 -2872 1193 -2871
rect 1332 -2872 1333 -2871
rect 1388 -2872 1389 -2871
rect 576 -2874 577 -2873
rect 1038 -2874 1039 -2873
rect 1332 -2874 1333 -2873
rect 1444 -2874 1445 -2873
rect 583 -2876 584 -2875
rect 611 -2876 612 -2875
rect 821 -2876 822 -2875
rect 1108 -2876 1109 -2875
rect 933 -2878 934 -2877
rect 975 -2878 976 -2877
rect 1017 -2878 1018 -2877
rect 1024 -2878 1025 -2877
rect 1038 -2878 1039 -2877
rect 1206 -2878 1207 -2877
rect 975 -2880 976 -2879
rect 1059 -2880 1060 -2879
rect 1108 -2880 1109 -2879
rect 1234 -2880 1235 -2879
rect 1059 -2882 1060 -2881
rect 1080 -2882 1081 -2881
rect 1206 -2882 1207 -2881
rect 1402 -2882 1403 -2881
rect 1080 -2884 1081 -2883
rect 1171 -2884 1172 -2883
rect 1234 -2884 1235 -2883
rect 1346 -2884 1347 -2883
rect 1402 -2884 1403 -2883
rect 1514 -2884 1515 -2883
rect 1171 -2886 1172 -2885
rect 1248 -2886 1249 -2885
rect 1346 -2886 1347 -2885
rect 1451 -2886 1452 -2885
rect 1248 -2888 1249 -2887
rect 1409 -2888 1410 -2887
rect 905 -2890 906 -2889
rect 1409 -2890 1410 -2889
rect 905 -2892 906 -2891
rect 968 -2892 969 -2891
rect 968 -2894 969 -2893
rect 1115 -2894 1116 -2893
rect 1115 -2896 1116 -2895
rect 1178 -2896 1179 -2895
rect 1178 -2898 1179 -2897
rect 1304 -2898 1305 -2897
rect 1304 -2900 1305 -2899
rect 1423 -2900 1424 -2899
rect 1416 -2902 1417 -2901
rect 1423 -2902 1424 -2901
rect 1031 -2904 1032 -2903
rect 1416 -2904 1417 -2903
rect 663 -2906 664 -2905
rect 1031 -2906 1032 -2905
rect 72 -2917 73 -2916
rect 247 -2917 248 -2916
rect 250 -2917 251 -2916
rect 569 -2917 570 -2916
rect 583 -2917 584 -2916
rect 954 -2917 955 -2916
rect 957 -2917 958 -2916
rect 1185 -2917 1186 -2916
rect 1227 -2917 1228 -2916
rect 1230 -2917 1231 -2916
rect 1360 -2917 1361 -2916
rect 1430 -2917 1431 -2916
rect 93 -2919 94 -2918
rect 124 -2919 125 -2918
rect 166 -2919 167 -2918
rect 576 -2919 577 -2918
rect 586 -2919 587 -2918
rect 618 -2919 619 -2918
rect 754 -2919 755 -2918
rect 793 -2919 794 -2918
rect 800 -2919 801 -2918
rect 1094 -2919 1095 -2918
rect 1097 -2919 1098 -2918
rect 1248 -2919 1249 -2918
rect 1360 -2919 1361 -2918
rect 1409 -2919 1410 -2918
rect 93 -2921 94 -2920
rect 205 -2921 206 -2920
rect 208 -2921 209 -2920
rect 310 -2921 311 -2920
rect 436 -2921 437 -2920
rect 702 -2921 703 -2920
rect 765 -2921 766 -2920
rect 793 -2921 794 -2920
rect 838 -2921 839 -2920
rect 1192 -2921 1193 -2920
rect 1227 -2921 1228 -2920
rect 1255 -2921 1256 -2920
rect 1409 -2921 1410 -2920
rect 1423 -2921 1424 -2920
rect 100 -2923 101 -2922
rect 149 -2923 150 -2922
rect 184 -2923 185 -2922
rect 285 -2923 286 -2922
rect 289 -2923 290 -2922
rect 296 -2923 297 -2922
rect 310 -2923 311 -2922
rect 324 -2923 325 -2922
rect 457 -2923 458 -2922
rect 824 -2923 825 -2922
rect 838 -2923 839 -2922
rect 884 -2923 885 -2922
rect 891 -2923 892 -2922
rect 894 -2923 895 -2922
rect 912 -2923 913 -2922
rect 1171 -2923 1172 -2922
rect 1185 -2923 1186 -2922
rect 1213 -2923 1214 -2922
rect 1248 -2923 1249 -2922
rect 1297 -2923 1298 -2922
rect 103 -2925 104 -2924
rect 744 -2925 745 -2924
rect 768 -2925 769 -2924
rect 1115 -2925 1116 -2924
rect 1192 -2925 1193 -2924
rect 1234 -2925 1235 -2924
rect 1276 -2925 1277 -2924
rect 1297 -2925 1298 -2924
rect 121 -2927 122 -2926
rect 849 -2927 850 -2926
rect 884 -2927 885 -2926
rect 926 -2927 927 -2926
rect 947 -2927 948 -2926
rect 982 -2927 983 -2926
rect 1017 -2927 1018 -2926
rect 1059 -2927 1060 -2926
rect 1076 -2927 1077 -2926
rect 1220 -2927 1221 -2926
rect 1234 -2927 1235 -2926
rect 1290 -2927 1291 -2926
rect 121 -2929 122 -2928
rect 212 -2929 213 -2928
rect 219 -2929 220 -2928
rect 576 -2929 577 -2928
rect 604 -2929 605 -2928
rect 618 -2929 619 -2928
rect 667 -2929 668 -2928
rect 702 -2929 703 -2928
rect 744 -2929 745 -2928
rect 751 -2929 752 -2928
rect 789 -2929 790 -2928
rect 1080 -2929 1081 -2928
rect 1087 -2929 1088 -2928
rect 1115 -2929 1116 -2928
rect 1213 -2929 1214 -2928
rect 1241 -2929 1242 -2928
rect 1269 -2929 1270 -2928
rect 1276 -2929 1277 -2928
rect 142 -2931 143 -2930
rect 436 -2931 437 -2930
rect 457 -2931 458 -2930
rect 590 -2931 591 -2930
rect 604 -2931 605 -2930
rect 737 -2931 738 -2930
rect 821 -2931 822 -2930
rect 982 -2931 983 -2930
rect 1024 -2931 1025 -2930
rect 1059 -2931 1060 -2930
rect 1080 -2931 1081 -2930
rect 1129 -2931 1130 -2930
rect 1220 -2931 1221 -2930
rect 1262 -2931 1263 -2930
rect 1269 -2931 1270 -2930
rect 1325 -2931 1326 -2930
rect 107 -2933 108 -2932
rect 590 -2933 591 -2932
rect 611 -2933 612 -2932
rect 642 -2933 643 -2932
rect 646 -2933 647 -2932
rect 667 -2933 668 -2932
rect 681 -2933 682 -2932
rect 849 -2933 850 -2932
rect 891 -2933 892 -2932
rect 905 -2933 906 -2932
rect 912 -2933 913 -2932
rect 989 -2933 990 -2932
rect 1094 -2933 1095 -2932
rect 1157 -2933 1158 -2932
rect 1206 -2933 1207 -2932
rect 1325 -2933 1326 -2932
rect 107 -2935 108 -2934
rect 548 -2935 549 -2934
rect 597 -2935 598 -2934
rect 611 -2935 612 -2934
rect 691 -2935 692 -2934
rect 1087 -2935 1088 -2934
rect 1101 -2935 1102 -2934
rect 1171 -2935 1172 -2934
rect 1230 -2935 1231 -2934
rect 1255 -2935 1256 -2934
rect 1262 -2935 1263 -2934
rect 1311 -2935 1312 -2934
rect 142 -2937 143 -2936
rect 646 -2937 647 -2936
rect 709 -2937 710 -2936
rect 737 -2937 738 -2936
rect 807 -2937 808 -2936
rect 1024 -2937 1025 -2936
rect 1052 -2937 1053 -2936
rect 1157 -2937 1158 -2936
rect 1241 -2937 1242 -2936
rect 1332 -2937 1333 -2936
rect 184 -2939 185 -2938
rect 639 -2939 640 -2938
rect 772 -2939 773 -2938
rect 807 -2939 808 -2938
rect 821 -2939 822 -2938
rect 870 -2939 871 -2938
rect 898 -2939 899 -2938
rect 947 -2939 948 -2938
rect 954 -2939 955 -2938
rect 961 -2939 962 -2938
rect 989 -2939 990 -2938
rect 1045 -2939 1046 -2938
rect 1066 -2939 1067 -2938
rect 1101 -2939 1102 -2938
rect 1129 -2939 1130 -2938
rect 1164 -2939 1165 -2938
rect 1304 -2939 1305 -2938
rect 1332 -2939 1333 -2938
rect 208 -2941 209 -2940
rect 233 -2941 234 -2940
rect 240 -2941 241 -2940
rect 800 -2941 801 -2940
rect 835 -2941 836 -2940
rect 1052 -2941 1053 -2940
rect 1108 -2941 1109 -2940
rect 1164 -2941 1165 -2940
rect 1311 -2941 1312 -2940
rect 1388 -2941 1389 -2940
rect 212 -2943 213 -2942
rect 366 -2943 367 -2942
rect 411 -2943 412 -2942
rect 1290 -2943 1291 -2942
rect 1388 -2943 1389 -2942
rect 1416 -2943 1417 -2942
rect 222 -2945 223 -2944
rect 450 -2945 451 -2944
rect 495 -2945 496 -2944
rect 926 -2945 927 -2944
rect 950 -2945 951 -2944
rect 1045 -2945 1046 -2944
rect 1143 -2945 1144 -2944
rect 1206 -2945 1207 -2944
rect 226 -2947 227 -2946
rect 268 -2947 269 -2946
rect 275 -2947 276 -2946
rect 583 -2947 584 -2946
rect 597 -2947 598 -2946
rect 625 -2947 626 -2946
rect 639 -2947 640 -2946
rect 660 -2947 661 -2946
rect 688 -2947 689 -2946
rect 835 -2947 836 -2946
rect 842 -2947 843 -2946
rect 1395 -2947 1396 -2946
rect 163 -2949 164 -2948
rect 268 -2949 269 -2948
rect 275 -2949 276 -2948
rect 422 -2949 423 -2948
rect 443 -2949 444 -2948
rect 681 -2949 682 -2948
rect 751 -2949 752 -2948
rect 1066 -2949 1067 -2948
rect 1143 -2949 1144 -2948
rect 1150 -2949 1151 -2948
rect 163 -2951 164 -2950
rect 380 -2951 381 -2950
rect 443 -2951 444 -2950
rect 471 -2951 472 -2950
rect 513 -2951 514 -2950
rect 625 -2951 626 -2950
rect 660 -2951 661 -2950
rect 1395 -2951 1396 -2950
rect 135 -2953 136 -2952
rect 471 -2953 472 -2952
rect 520 -2953 521 -2952
rect 649 -2953 650 -2952
rect 772 -2953 773 -2952
rect 786 -2953 787 -2952
rect 842 -2953 843 -2952
rect 856 -2953 857 -2952
rect 870 -2953 871 -2952
rect 1122 -2953 1123 -2952
rect 135 -2955 136 -2954
rect 653 -2955 654 -2954
rect 898 -2955 899 -2954
rect 933 -2955 934 -2954
rect 961 -2955 962 -2954
rect 975 -2955 976 -2954
rect 1017 -2955 1018 -2954
rect 1122 -2955 1123 -2954
rect 149 -2957 150 -2956
rect 856 -2957 857 -2956
rect 915 -2957 916 -2956
rect 1038 -2957 1039 -2956
rect 191 -2959 192 -2958
rect 422 -2959 423 -2958
rect 464 -2959 465 -2958
rect 933 -2959 934 -2958
rect 1031 -2959 1032 -2958
rect 1304 -2959 1305 -2958
rect 191 -2961 192 -2960
rect 198 -2961 199 -2960
rect 229 -2961 230 -2960
rect 632 -2961 633 -2960
rect 786 -2961 787 -2960
rect 975 -2961 976 -2960
rect 1038 -2961 1039 -2960
rect 1073 -2961 1074 -2960
rect 86 -2963 87 -2962
rect 198 -2963 199 -2962
rect 233 -2963 234 -2962
rect 292 -2963 293 -2962
rect 296 -2963 297 -2962
rect 688 -2963 689 -2962
rect 919 -2963 920 -2962
rect 1003 -2963 1004 -2962
rect 1073 -2963 1074 -2962
rect 1318 -2963 1319 -2962
rect 79 -2965 80 -2964
rect 86 -2965 87 -2964
rect 219 -2965 220 -2964
rect 919 -2965 920 -2964
rect 940 -2965 941 -2964
rect 1031 -2965 1032 -2964
rect 1283 -2965 1284 -2964
rect 1318 -2965 1319 -2964
rect 240 -2967 241 -2966
rect 373 -2967 374 -2966
rect 387 -2967 388 -2966
rect 653 -2967 654 -2966
rect 674 -2967 675 -2966
rect 940 -2967 941 -2966
rect 1003 -2967 1004 -2966
rect 1010 -2967 1011 -2966
rect 1283 -2967 1284 -2966
rect 1339 -2967 1340 -2966
rect 170 -2969 171 -2968
rect 387 -2969 388 -2968
rect 401 -2969 402 -2968
rect 513 -2969 514 -2968
rect 520 -2969 521 -2968
rect 866 -2969 867 -2968
rect 1339 -2969 1340 -2968
rect 1346 -2969 1347 -2968
rect 170 -2971 171 -2970
rect 873 -2971 874 -2970
rect 1346 -2971 1347 -2970
rect 1381 -2971 1382 -2970
rect 247 -2973 248 -2972
rect 761 -2973 762 -2972
rect 282 -2975 283 -2974
rect 747 -2975 748 -2974
rect 254 -2977 255 -2976
rect 282 -2977 283 -2976
rect 289 -2977 290 -2976
rect 663 -2977 664 -2976
rect 674 -2977 675 -2976
rect 915 -2977 916 -2976
rect 254 -2979 255 -2978
rect 278 -2979 279 -2978
rect 303 -2979 304 -2978
rect 366 -2979 367 -2978
rect 373 -2979 374 -2978
rect 394 -2979 395 -2978
rect 464 -2979 465 -2978
rect 485 -2979 486 -2978
rect 534 -2979 535 -2978
rect 569 -2979 570 -2978
rect 632 -2979 633 -2978
rect 1108 -2979 1109 -2978
rect 261 -2981 262 -2980
rect 534 -2981 535 -2980
rect 548 -2981 549 -2980
rect 877 -2981 878 -2980
rect 261 -2983 262 -2982
rect 380 -2983 381 -2982
rect 394 -2983 395 -2982
rect 408 -2983 409 -2982
rect 485 -2983 486 -2982
rect 716 -2983 717 -2982
rect 303 -2985 304 -2984
rect 317 -2985 318 -2984
rect 324 -2985 325 -2984
rect 506 -2985 507 -2984
rect 555 -2985 556 -2984
rect 866 -2985 867 -2984
rect 317 -2987 318 -2986
rect 338 -2987 339 -2986
rect 345 -2987 346 -2986
rect 450 -2987 451 -2986
rect 562 -2987 563 -2986
rect 709 -2987 710 -2986
rect 716 -2987 717 -2986
rect 863 -2987 864 -2986
rect 145 -2989 146 -2988
rect 338 -2989 339 -2988
rect 345 -2989 346 -2988
rect 499 -2989 500 -2988
rect 695 -2989 696 -2988
rect 863 -2989 864 -2988
rect 264 -2991 265 -2990
rect 562 -2991 563 -2990
rect 698 -2991 699 -2990
rect 1010 -2991 1011 -2990
rect 359 -2993 360 -2992
rect 401 -2993 402 -2992
rect 408 -2993 409 -2992
rect 877 -2993 878 -2992
rect 359 -2995 360 -2994
rect 478 -2995 479 -2994
rect 499 -2995 500 -2994
rect 635 -2995 636 -2994
rect 705 -2995 706 -2994
rect 1381 -2995 1382 -2994
rect 429 -2997 430 -2996
rect 695 -2997 696 -2996
rect 177 -2999 178 -2998
rect 429 -2999 430 -2998
rect 478 -2999 479 -2998
rect 541 -2999 542 -2998
rect 156 -3001 157 -3000
rect 177 -3001 178 -3000
rect 541 -3001 542 -3000
rect 723 -3001 724 -3000
rect 156 -3003 157 -3002
rect 352 -3003 353 -3002
rect 723 -3003 724 -3002
rect 730 -3003 731 -3002
rect 352 -3005 353 -3004
rect 415 -3005 416 -3004
rect 730 -3005 731 -3004
rect 814 -3005 815 -3004
rect 331 -3007 332 -3006
rect 415 -3007 416 -3006
rect 779 -3007 780 -3006
rect 814 -3007 815 -3006
rect 114 -3009 115 -3008
rect 331 -3009 332 -3008
rect 779 -3009 780 -3008
rect 922 -3009 923 -3008
rect 114 -3011 115 -3010
rect 1020 -3011 1021 -3010
rect 922 -3013 923 -3012
rect 1353 -3013 1354 -3012
rect 1353 -3015 1354 -3014
rect 1367 -3015 1368 -3014
rect 1367 -3017 1368 -3016
rect 1374 -3017 1375 -3016
rect 1374 -3019 1375 -3018
rect 1402 -3019 1403 -3018
rect 758 -3021 759 -3020
rect 1402 -3021 1403 -3020
rect 527 -3023 528 -3022
rect 758 -3023 759 -3022
rect 527 -3025 528 -3024
rect 663 -3025 664 -3024
rect 86 -3036 87 -3035
rect 149 -3036 150 -3035
rect 156 -3036 157 -3035
rect 408 -3036 409 -3035
rect 411 -3036 412 -3035
rect 653 -3036 654 -3035
rect 660 -3036 661 -3035
rect 982 -3036 983 -3035
rect 1017 -3036 1018 -3035
rect 1045 -3036 1046 -3035
rect 1073 -3036 1074 -3035
rect 1402 -3036 1403 -3035
rect 93 -3038 94 -3037
rect 810 -3038 811 -3037
rect 835 -3038 836 -3037
rect 1171 -3038 1172 -3037
rect 100 -3040 101 -3039
rect 152 -3040 153 -3039
rect 198 -3040 199 -3039
rect 208 -3040 209 -3039
rect 275 -3040 276 -3039
rect 278 -3040 279 -3039
rect 289 -3040 290 -3039
rect 506 -3040 507 -3039
rect 516 -3040 517 -3039
rect 541 -3040 542 -3039
rect 555 -3040 556 -3039
rect 653 -3040 654 -3039
rect 660 -3040 661 -3039
rect 877 -3040 878 -3039
rect 919 -3040 920 -3039
rect 1332 -3040 1333 -3039
rect 100 -3042 101 -3041
rect 128 -3042 129 -3041
rect 135 -3042 136 -3041
rect 205 -3042 206 -3041
rect 275 -3042 276 -3041
rect 366 -3042 367 -3041
rect 422 -3042 423 -3041
rect 915 -3042 916 -3041
rect 926 -3042 927 -3041
rect 1335 -3042 1336 -3041
rect 107 -3044 108 -3043
rect 222 -3044 223 -3043
rect 310 -3044 311 -3043
rect 411 -3044 412 -3043
rect 471 -3044 472 -3043
rect 541 -3044 542 -3043
rect 576 -3044 577 -3043
rect 632 -3044 633 -3043
rect 681 -3044 682 -3043
rect 695 -3044 696 -3043
rect 698 -3044 699 -3043
rect 989 -3044 990 -3043
rect 1020 -3044 1021 -3043
rect 1276 -3044 1277 -3043
rect 107 -3046 108 -3045
rect 261 -3046 262 -3045
rect 310 -3046 311 -3045
rect 866 -3046 867 -3045
rect 873 -3046 874 -3045
rect 1395 -3046 1396 -3045
rect 128 -3048 129 -3047
rect 233 -3048 234 -3047
rect 324 -3048 325 -3047
rect 838 -3048 839 -3047
rect 863 -3048 864 -3047
rect 1325 -3048 1326 -3047
rect 135 -3050 136 -3049
rect 1209 -3050 1210 -3049
rect 1241 -3050 1242 -3049
rect 1276 -3050 1277 -3049
rect 1325 -3050 1326 -3049
rect 1381 -3050 1382 -3049
rect 149 -3052 150 -3051
rect 922 -3052 923 -3051
rect 926 -3052 927 -3051
rect 996 -3052 997 -3051
rect 1038 -3052 1039 -3051
rect 1073 -3052 1074 -3051
rect 1136 -3052 1137 -3051
rect 1171 -3052 1172 -3051
rect 1241 -3052 1242 -3051
rect 1269 -3052 1270 -3051
rect 170 -3054 171 -3053
rect 198 -3054 199 -3053
rect 229 -3054 230 -3053
rect 261 -3054 262 -3053
rect 327 -3054 328 -3053
rect 646 -3054 647 -3053
rect 691 -3054 692 -3053
rect 1255 -3054 1256 -3053
rect 170 -3056 171 -3055
rect 247 -3056 248 -3055
rect 338 -3056 339 -3055
rect 471 -3056 472 -3055
rect 513 -3056 514 -3055
rect 555 -3056 556 -3055
rect 583 -3056 584 -3055
rect 989 -3056 990 -3055
rect 1038 -3056 1039 -3055
rect 1066 -3056 1067 -3055
rect 1115 -3056 1116 -3055
rect 1136 -3056 1137 -3055
rect 1150 -3056 1151 -3055
rect 1297 -3056 1298 -3055
rect 184 -3058 185 -3057
rect 289 -3058 290 -3057
rect 338 -3058 339 -3057
rect 527 -3058 528 -3057
rect 534 -3058 535 -3057
rect 607 -3058 608 -3057
rect 618 -3058 619 -3057
rect 649 -3058 650 -3057
rect 698 -3058 699 -3057
rect 1178 -3058 1179 -3057
rect 1234 -3058 1235 -3057
rect 1255 -3058 1256 -3057
rect 1297 -3058 1298 -3057
rect 1332 -3058 1333 -3057
rect 184 -3060 185 -3059
rect 226 -3060 227 -3059
rect 233 -3060 234 -3059
rect 254 -3060 255 -3059
rect 345 -3060 346 -3059
rect 509 -3060 510 -3059
rect 527 -3060 528 -3059
rect 590 -3060 591 -3059
rect 618 -3060 619 -3059
rect 765 -3060 766 -3059
rect 789 -3060 790 -3059
rect 870 -3060 871 -3059
rect 877 -3060 878 -3059
rect 1220 -3060 1221 -3059
rect 121 -3062 122 -3061
rect 226 -3062 227 -3061
rect 345 -3062 346 -3061
rect 436 -3062 437 -3061
rect 443 -3062 444 -3061
rect 576 -3062 577 -3061
rect 590 -3062 591 -3061
rect 1087 -3062 1088 -3061
rect 1150 -3062 1151 -3061
rect 1206 -3062 1207 -3061
rect 1220 -3062 1221 -3061
rect 1227 -3062 1228 -3061
rect 121 -3064 122 -3063
rect 219 -3064 220 -3063
rect 331 -3064 332 -3063
rect 436 -3064 437 -3063
rect 464 -3064 465 -3063
rect 513 -3064 514 -3063
rect 534 -3064 535 -3063
rect 597 -3064 598 -3063
rect 635 -3064 636 -3063
rect 681 -3064 682 -3063
rect 730 -3064 731 -3063
rect 733 -3064 734 -3063
rect 740 -3064 741 -3063
rect 947 -3064 948 -3063
rect 982 -3064 983 -3063
rect 1202 -3064 1203 -3063
rect 1213 -3064 1214 -3063
rect 1227 -3064 1228 -3063
rect 166 -3066 167 -3065
rect 331 -3066 332 -3065
rect 352 -3066 353 -3065
rect 366 -3066 367 -3065
rect 380 -3066 381 -3065
rect 464 -3066 465 -3065
rect 478 -3066 479 -3065
rect 583 -3066 584 -3065
rect 597 -3066 598 -3065
rect 667 -3066 668 -3065
rect 730 -3066 731 -3065
rect 793 -3066 794 -3065
rect 796 -3066 797 -3065
rect 1234 -3066 1235 -3065
rect 177 -3068 178 -3067
rect 254 -3068 255 -3067
rect 257 -3068 258 -3067
rect 478 -3068 479 -3067
rect 520 -3068 521 -3067
rect 667 -3068 668 -3067
rect 744 -3068 745 -3067
rect 765 -3068 766 -3067
rect 835 -3068 836 -3067
rect 842 -3068 843 -3067
rect 863 -3068 864 -3067
rect 891 -3068 892 -3067
rect 898 -3068 899 -3067
rect 919 -3068 920 -3067
rect 1045 -3068 1046 -3067
rect 1101 -3068 1102 -3067
rect 1178 -3068 1179 -3067
rect 1367 -3068 1368 -3067
rect 177 -3070 178 -3069
rect 499 -3070 500 -3069
rect 520 -3070 521 -3069
rect 639 -3070 640 -3069
rect 649 -3070 650 -3069
rect 1087 -3070 1088 -3069
rect 1101 -3070 1102 -3069
rect 1122 -3070 1123 -3069
rect 1213 -3070 1214 -3069
rect 1304 -3070 1305 -3069
rect 1367 -3070 1368 -3069
rect 1388 -3070 1389 -3069
rect 282 -3072 283 -3071
rect 352 -3072 353 -3071
rect 380 -3072 381 -3071
rect 457 -3072 458 -3071
rect 499 -3072 500 -3071
rect 604 -3072 605 -3071
rect 611 -3072 612 -3071
rect 639 -3072 640 -3071
rect 744 -3072 745 -3071
rect 1157 -3072 1158 -3071
rect 1304 -3072 1305 -3071
rect 1353 -3072 1354 -3071
rect 394 -3074 395 -3073
rect 422 -3074 423 -3073
rect 429 -3074 430 -3073
rect 457 -3074 458 -3073
rect 548 -3074 549 -3073
rect 611 -3074 612 -3073
rect 733 -3074 734 -3073
rect 793 -3074 794 -3073
rect 842 -3074 843 -3073
rect 905 -3074 906 -3073
rect 933 -3074 934 -3073
rect 1157 -3074 1158 -3073
rect 1353 -3074 1354 -3073
rect 1360 -3074 1361 -3073
rect 303 -3076 304 -3075
rect 548 -3076 549 -3075
rect 747 -3076 748 -3075
rect 1269 -3076 1270 -3075
rect 1360 -3076 1361 -3075
rect 1374 -3076 1375 -3075
rect 303 -3078 304 -3077
rect 387 -3078 388 -3077
rect 394 -3078 395 -3077
rect 761 -3078 762 -3077
rect 887 -3078 888 -3077
rect 947 -3078 948 -3077
rect 1059 -3078 1060 -3077
rect 1066 -3078 1067 -3077
rect 1122 -3078 1123 -3077
rect 1129 -3078 1130 -3077
rect 1374 -3078 1375 -3077
rect 1409 -3078 1410 -3077
rect 401 -3080 402 -3079
rect 429 -3080 430 -3079
rect 751 -3080 752 -3079
rect 779 -3080 780 -3079
rect 891 -3080 892 -3079
rect 954 -3080 955 -3079
rect 1059 -3080 1060 -3079
rect 1080 -3080 1081 -3079
rect 1108 -3080 1109 -3079
rect 1129 -3080 1130 -3079
rect 296 -3082 297 -3081
rect 401 -3082 402 -3081
rect 415 -3082 416 -3081
rect 443 -3082 444 -3081
rect 772 -3082 773 -3081
rect 779 -3082 780 -3081
rect 898 -3082 899 -3081
rect 1199 -3082 1200 -3081
rect 296 -3084 297 -3083
rect 373 -3084 374 -3083
rect 415 -3084 416 -3083
rect 754 -3084 755 -3083
rect 758 -3084 759 -3083
rect 772 -3084 773 -3083
rect 901 -3084 902 -3083
rect 1115 -3084 1116 -3083
rect 373 -3086 374 -3085
rect 688 -3086 689 -3085
rect 905 -3086 906 -3085
rect 1024 -3086 1025 -3085
rect 1080 -3086 1081 -3085
rect 1143 -3086 1144 -3085
rect 688 -3088 689 -3087
rect 723 -3088 724 -3087
rect 933 -3088 934 -3087
rect 961 -3088 962 -3087
rect 1024 -3088 1025 -3087
rect 1052 -3088 1053 -3087
rect 1108 -3088 1109 -3087
rect 1192 -3088 1193 -3087
rect 674 -3090 675 -3089
rect 1052 -3090 1053 -3089
rect 1143 -3090 1144 -3089
rect 1185 -3090 1186 -3089
rect 1192 -3090 1193 -3089
rect 1290 -3090 1291 -3089
rect 674 -3092 675 -3091
rect 702 -3092 703 -3091
rect 716 -3092 717 -3091
rect 723 -3092 724 -3091
rect 940 -3092 941 -3091
rect 961 -3092 962 -3091
rect 1003 -3092 1004 -3091
rect 1185 -3092 1186 -3091
rect 1290 -3092 1291 -3091
rect 1339 -3092 1340 -3091
rect 485 -3094 486 -3093
rect 716 -3094 717 -3093
rect 940 -3094 941 -3093
rect 968 -3094 969 -3093
rect 1003 -3094 1004 -3093
rect 1031 -3094 1032 -3093
rect 1339 -3094 1340 -3093
rect 1346 -3094 1347 -3093
rect 317 -3096 318 -3095
rect 485 -3096 486 -3095
rect 702 -3096 703 -3095
rect 709 -3096 710 -3095
rect 912 -3096 913 -3095
rect 968 -3096 969 -3095
rect 1031 -3096 1032 -3095
rect 1094 -3096 1095 -3095
rect 163 -3098 164 -3097
rect 1094 -3098 1095 -3097
rect 163 -3100 164 -3099
rect 268 -3100 269 -3099
rect 317 -3100 318 -3099
rect 359 -3100 360 -3099
rect 562 -3100 563 -3099
rect 709 -3100 710 -3099
rect 912 -3100 913 -3099
rect 1164 -3100 1165 -3099
rect 212 -3102 213 -3101
rect 268 -3102 269 -3101
rect 324 -3102 325 -3101
rect 562 -3102 563 -3101
rect 954 -3102 955 -3101
rect 975 -3102 976 -3101
rect 1164 -3102 1165 -3101
rect 1262 -3102 1263 -3101
rect 191 -3104 192 -3103
rect 212 -3104 213 -3103
rect 240 -3104 241 -3103
rect 359 -3104 360 -3103
rect 975 -3104 976 -3103
rect 1010 -3104 1011 -3103
rect 1248 -3104 1249 -3103
rect 1262 -3104 1263 -3103
rect 156 -3106 157 -3105
rect 191 -3106 192 -3105
rect 240 -3106 241 -3105
rect 1153 -3106 1154 -3105
rect 695 -3108 696 -3107
rect 1248 -3108 1249 -3107
rect 1010 -3110 1011 -3109
rect 1318 -3110 1319 -3109
rect 1311 -3112 1312 -3111
rect 1318 -3112 1319 -3111
rect 884 -3114 885 -3113
rect 1311 -3114 1312 -3113
rect 856 -3116 857 -3115
rect 884 -3116 885 -3115
rect 849 -3118 850 -3117
rect 856 -3118 857 -3117
rect 828 -3120 829 -3119
rect 849 -3120 850 -3119
rect 814 -3122 815 -3121
rect 828 -3122 829 -3121
rect 814 -3124 815 -3123
rect 821 -3124 822 -3123
rect 737 -3126 738 -3125
rect 821 -3126 822 -3125
rect 492 -3128 493 -3127
rect 737 -3128 738 -3127
rect 492 -3130 493 -3129
rect 786 -3130 787 -3129
rect 786 -3132 787 -3131
rect 800 -3132 801 -3131
rect 800 -3134 801 -3133
rect 807 -3134 808 -3133
rect 807 -3136 808 -3135
rect 996 -3136 997 -3135
rect 100 -3147 101 -3146
rect 159 -3147 160 -3146
rect 184 -3147 185 -3146
rect 324 -3147 325 -3146
rect 331 -3147 332 -3146
rect 390 -3147 391 -3146
rect 394 -3147 395 -3146
rect 754 -3147 755 -3146
rect 758 -3147 759 -3146
rect 814 -3147 815 -3146
rect 898 -3147 899 -3146
rect 1171 -3147 1172 -3146
rect 1199 -3147 1200 -3146
rect 1220 -3147 1221 -3146
rect 1293 -3147 1294 -3146
rect 1339 -3147 1340 -3146
rect 1346 -3147 1347 -3146
rect 1360 -3147 1361 -3146
rect 107 -3149 108 -3148
rect 285 -3149 286 -3148
rect 296 -3149 297 -3148
rect 695 -3149 696 -3148
rect 698 -3149 699 -3148
rect 968 -3149 969 -3148
rect 1171 -3149 1172 -3148
rect 1213 -3149 1214 -3148
rect 1335 -3149 1336 -3148
rect 1367 -3149 1368 -3148
rect 114 -3151 115 -3150
rect 187 -3151 188 -3150
rect 191 -3151 192 -3150
rect 250 -3151 251 -3150
rect 254 -3151 255 -3150
rect 373 -3151 374 -3150
rect 387 -3151 388 -3150
rect 485 -3151 486 -3150
rect 492 -3151 493 -3150
rect 810 -3151 811 -3150
rect 870 -3151 871 -3150
rect 898 -3151 899 -3150
rect 912 -3151 913 -3150
rect 1199 -3151 1200 -3150
rect 1206 -3151 1207 -3150
rect 1241 -3151 1242 -3150
rect 1360 -3151 1361 -3150
rect 1374 -3151 1375 -3150
rect 121 -3153 122 -3152
rect 222 -3153 223 -3152
rect 247 -3153 248 -3152
rect 352 -3153 353 -3152
rect 373 -3153 374 -3152
rect 429 -3153 430 -3152
rect 460 -3153 461 -3152
rect 527 -3153 528 -3152
rect 593 -3153 594 -3152
rect 1286 -3153 1287 -3152
rect 177 -3155 178 -3154
rect 387 -3155 388 -3154
rect 394 -3155 395 -3154
rect 457 -3155 458 -3154
rect 464 -3155 465 -3154
rect 544 -3155 545 -3154
rect 607 -3155 608 -3154
rect 1157 -3155 1158 -3154
rect 1206 -3155 1207 -3154
rect 1276 -3155 1277 -3154
rect 177 -3157 178 -3156
rect 768 -3157 769 -3156
rect 807 -3157 808 -3156
rect 894 -3157 895 -3156
rect 915 -3157 916 -3156
rect 1230 -3157 1231 -3156
rect 1241 -3157 1242 -3156
rect 1318 -3157 1319 -3156
rect 191 -3159 192 -3158
rect 747 -3159 748 -3158
rect 758 -3159 759 -3158
rect 849 -3159 850 -3158
rect 870 -3159 871 -3158
rect 884 -3159 885 -3158
rect 943 -3159 944 -3158
rect 1136 -3159 1137 -3158
rect 1209 -3159 1210 -3158
rect 1220 -3159 1221 -3158
rect 1276 -3159 1277 -3158
rect 1325 -3159 1326 -3158
rect 198 -3161 199 -3160
rect 226 -3161 227 -3160
rect 233 -3161 234 -3160
rect 247 -3161 248 -3160
rect 275 -3161 276 -3160
rect 296 -3161 297 -3160
rect 327 -3161 328 -3160
rect 485 -3161 486 -3160
rect 492 -3161 493 -3160
rect 611 -3161 612 -3160
rect 618 -3161 619 -3160
rect 1010 -3161 1011 -3160
rect 1059 -3161 1060 -3160
rect 1136 -3161 1137 -3160
rect 1213 -3161 1214 -3160
rect 1304 -3161 1305 -3160
rect 128 -3163 129 -3162
rect 198 -3163 199 -3162
rect 219 -3163 220 -3162
rect 289 -3163 290 -3162
rect 331 -3163 332 -3162
rect 380 -3163 381 -3162
rect 401 -3163 402 -3162
rect 618 -3163 619 -3162
rect 635 -3163 636 -3162
rect 828 -3163 829 -3162
rect 849 -3163 850 -3162
rect 975 -3163 976 -3162
rect 1234 -3163 1235 -3162
rect 1304 -3163 1305 -3162
rect 135 -3165 136 -3164
rect 275 -3165 276 -3164
rect 338 -3165 339 -3164
rect 590 -3165 591 -3164
rect 611 -3165 612 -3164
rect 681 -3165 682 -3164
rect 695 -3165 696 -3164
rect 772 -3165 773 -3164
rect 810 -3165 811 -3164
rect 1185 -3165 1186 -3164
rect 1234 -3165 1235 -3164
rect 1290 -3165 1291 -3164
rect 184 -3167 185 -3166
rect 289 -3167 290 -3166
rect 338 -3167 339 -3166
rect 366 -3167 367 -3166
rect 401 -3167 402 -3166
rect 436 -3167 437 -3166
rect 464 -3167 465 -3166
rect 1332 -3167 1333 -3166
rect 233 -3169 234 -3168
rect 282 -3169 283 -3168
rect 345 -3169 346 -3168
rect 747 -3169 748 -3168
rect 772 -3169 773 -3168
rect 786 -3169 787 -3168
rect 877 -3169 878 -3168
rect 1059 -3169 1060 -3168
rect 1108 -3169 1109 -3168
rect 1185 -3169 1186 -3168
rect 282 -3171 283 -3170
rect 324 -3171 325 -3170
rect 345 -3171 346 -3170
rect 450 -3171 451 -3170
rect 506 -3171 507 -3170
rect 744 -3171 745 -3170
rect 761 -3171 762 -3170
rect 786 -3171 787 -3170
rect 877 -3171 878 -3170
rect 954 -3171 955 -3170
rect 968 -3171 969 -3170
rect 982 -3171 983 -3170
rect 1108 -3171 1109 -3170
rect 1227 -3171 1228 -3170
rect 205 -3173 206 -3172
rect 450 -3173 451 -3172
rect 471 -3173 472 -3172
rect 506 -3173 507 -3172
rect 520 -3173 521 -3172
rect 737 -3173 738 -3172
rect 740 -3173 741 -3172
rect 1157 -3173 1158 -3172
rect 205 -3175 206 -3174
rect 261 -3175 262 -3174
rect 352 -3175 353 -3174
rect 534 -3175 535 -3174
rect 590 -3175 591 -3174
rect 744 -3175 745 -3174
rect 884 -3175 885 -3174
rect 891 -3175 892 -3174
rect 905 -3175 906 -3174
rect 954 -3175 955 -3174
rect 975 -3175 976 -3174
rect 1024 -3175 1025 -3174
rect 142 -3177 143 -3176
rect 261 -3177 262 -3176
rect 317 -3177 318 -3176
rect 891 -3177 892 -3176
rect 905 -3177 906 -3176
rect 933 -3177 934 -3176
rect 982 -3177 983 -3176
rect 1017 -3177 1018 -3176
rect 1024 -3177 1025 -3176
rect 1101 -3177 1102 -3176
rect 240 -3179 241 -3178
rect 317 -3179 318 -3178
rect 359 -3179 360 -3178
rect 380 -3179 381 -3178
rect 415 -3179 416 -3178
rect 429 -3179 430 -3178
rect 471 -3179 472 -3178
rect 555 -3179 556 -3178
rect 625 -3179 626 -3178
rect 737 -3179 738 -3178
rect 919 -3179 920 -3178
rect 1010 -3179 1011 -3178
rect 1101 -3179 1102 -3178
rect 1143 -3179 1144 -3178
rect 240 -3181 241 -3180
rect 604 -3181 605 -3180
rect 646 -3181 647 -3180
rect 765 -3181 766 -3180
rect 919 -3181 920 -3180
rect 1202 -3181 1203 -3180
rect 359 -3183 360 -3182
rect 411 -3183 412 -3182
rect 422 -3183 423 -3182
rect 436 -3183 437 -3182
rect 443 -3183 444 -3182
rect 604 -3183 605 -3182
rect 646 -3183 647 -3182
rect 709 -3183 710 -3182
rect 716 -3183 717 -3182
rect 901 -3183 902 -3182
rect 926 -3183 927 -3182
rect 933 -3183 934 -3182
rect 996 -3183 997 -3182
rect 1017 -3183 1018 -3182
rect 1143 -3183 1144 -3182
rect 1262 -3183 1263 -3182
rect 366 -3185 367 -3184
rect 639 -3185 640 -3184
rect 667 -3185 668 -3184
rect 828 -3185 829 -3184
rect 926 -3185 927 -3184
rect 1003 -3185 1004 -3184
rect 1150 -3185 1151 -3184
rect 1202 -3185 1203 -3184
rect 408 -3187 409 -3186
rect 415 -3187 416 -3186
rect 422 -3187 423 -3186
rect 499 -3187 500 -3186
rect 513 -3187 514 -3186
rect 625 -3187 626 -3186
rect 667 -3187 668 -3186
rect 793 -3187 794 -3186
rect 961 -3187 962 -3186
rect 1262 -3187 1263 -3186
rect 163 -3189 164 -3188
rect 408 -3189 409 -3188
rect 443 -3189 444 -3188
rect 457 -3189 458 -3188
rect 513 -3189 514 -3188
rect 653 -3189 654 -3188
rect 681 -3189 682 -3188
rect 751 -3189 752 -3188
rect 765 -3189 766 -3188
rect 1311 -3189 1312 -3188
rect 156 -3191 157 -3190
rect 163 -3191 164 -3190
rect 303 -3191 304 -3190
rect 499 -3191 500 -3190
rect 520 -3191 521 -3190
rect 548 -3191 549 -3190
rect 555 -3191 556 -3190
rect 569 -3191 570 -3190
rect 597 -3191 598 -3190
rect 639 -3191 640 -3190
rect 709 -3191 710 -3190
rect 1178 -3191 1179 -3190
rect 303 -3193 304 -3192
rect 310 -3193 311 -3192
rect 527 -3193 528 -3192
rect 541 -3193 542 -3192
rect 548 -3193 549 -3192
rect 576 -3193 577 -3192
rect 597 -3193 598 -3192
rect 807 -3193 808 -3192
rect 996 -3193 997 -3192
rect 1094 -3193 1095 -3192
rect 1150 -3193 1151 -3192
rect 1269 -3193 1270 -3192
rect 149 -3195 150 -3194
rect 310 -3195 311 -3194
rect 534 -3195 535 -3194
rect 821 -3195 822 -3194
rect 947 -3195 948 -3194
rect 1094 -3195 1095 -3194
rect 562 -3197 563 -3196
rect 653 -3197 654 -3196
rect 716 -3197 717 -3196
rect 730 -3197 731 -3196
rect 751 -3197 752 -3196
rect 1178 -3197 1179 -3196
rect 562 -3199 563 -3198
rect 583 -3199 584 -3198
rect 730 -3199 731 -3198
rect 779 -3199 780 -3198
rect 793 -3199 794 -3198
rect 800 -3199 801 -3198
rect 821 -3199 822 -3198
rect 835 -3199 836 -3198
rect 940 -3199 941 -3198
rect 947 -3199 948 -3198
rect 1003 -3199 1004 -3198
rect 1073 -3199 1074 -3198
rect 170 -3201 171 -3200
rect 800 -3201 801 -3200
rect 835 -3201 836 -3200
rect 856 -3201 857 -3200
rect 940 -3201 941 -3200
rect 1066 -3201 1067 -3200
rect 170 -3203 171 -3202
rect 723 -3203 724 -3202
rect 856 -3203 857 -3202
rect 989 -3203 990 -3202
rect 1031 -3203 1032 -3202
rect 1073 -3203 1074 -3202
rect 478 -3205 479 -3204
rect 779 -3205 780 -3204
rect 989 -3205 990 -3204
rect 1038 -3205 1039 -3204
rect 1066 -3205 1067 -3204
rect 1255 -3205 1256 -3204
rect 478 -3207 479 -3206
rect 1129 -3207 1130 -3206
rect 516 -3209 517 -3208
rect 583 -3209 584 -3208
rect 723 -3209 724 -3208
rect 1087 -3209 1088 -3208
rect 1129 -3209 1130 -3208
rect 1248 -3209 1249 -3208
rect 569 -3211 570 -3210
rect 632 -3211 633 -3210
rect 814 -3211 815 -3210
rect 1255 -3211 1256 -3210
rect 229 -3213 230 -3212
rect 632 -3213 633 -3212
rect 1031 -3213 1032 -3212
rect 1115 -3213 1116 -3212
rect 1248 -3213 1249 -3212
rect 1283 -3213 1284 -3212
rect 576 -3215 577 -3214
rect 702 -3215 703 -3214
rect 961 -3215 962 -3214
rect 1115 -3215 1116 -3214
rect 1269 -3215 1270 -3214
rect 1283 -3215 1284 -3214
rect 688 -3217 689 -3216
rect 702 -3217 703 -3216
rect 1038 -3217 1039 -3216
rect 1052 -3217 1053 -3216
rect 1087 -3217 1088 -3216
rect 1290 -3217 1291 -3216
rect 660 -3219 661 -3218
rect 688 -3219 689 -3218
rect 1052 -3219 1053 -3218
rect 1080 -3219 1081 -3218
rect 660 -3221 661 -3220
rect 674 -3221 675 -3220
rect 1080 -3221 1081 -3220
rect 1122 -3221 1123 -3220
rect 674 -3223 675 -3222
rect 1167 -3223 1168 -3222
rect 1122 -3225 1123 -3224
rect 1164 -3225 1165 -3224
rect 1164 -3227 1165 -3226
rect 1192 -3227 1193 -3226
rect 796 -3229 797 -3228
rect 1192 -3229 1193 -3228
rect 156 -3240 157 -3239
rect 212 -3240 213 -3239
rect 219 -3240 220 -3239
rect 460 -3240 461 -3239
rect 499 -3240 500 -3239
rect 709 -3240 710 -3239
rect 712 -3240 713 -3239
rect 1255 -3240 1256 -3239
rect 1290 -3240 1291 -3239
rect 1304 -3240 1305 -3239
rect 1339 -3240 1340 -3239
rect 1360 -3240 1361 -3239
rect 163 -3242 164 -3241
rect 201 -3242 202 -3241
rect 212 -3242 213 -3241
rect 240 -3242 241 -3241
rect 243 -3242 244 -3241
rect 324 -3242 325 -3241
rect 352 -3242 353 -3241
rect 663 -3242 664 -3241
rect 733 -3242 734 -3241
rect 814 -3242 815 -3241
rect 838 -3242 839 -3241
rect 1192 -3242 1193 -3241
rect 1199 -3242 1200 -3241
rect 1206 -3242 1207 -3241
rect 1227 -3242 1228 -3241
rect 1283 -3242 1284 -3241
rect 1293 -3242 1294 -3241
rect 1297 -3242 1298 -3241
rect 1346 -3242 1347 -3241
rect 1349 -3242 1350 -3241
rect 163 -3244 164 -3243
rect 366 -3244 367 -3243
rect 394 -3244 395 -3243
rect 544 -3244 545 -3243
rect 548 -3244 549 -3243
rect 576 -3244 577 -3243
rect 632 -3244 633 -3243
rect 681 -3244 682 -3243
rect 744 -3244 745 -3243
rect 1066 -3244 1067 -3243
rect 1136 -3244 1137 -3243
rect 1255 -3244 1256 -3243
rect 1346 -3244 1347 -3243
rect 1353 -3244 1354 -3243
rect 170 -3246 171 -3245
rect 481 -3246 482 -3245
rect 499 -3246 500 -3245
rect 747 -3246 748 -3245
rect 751 -3246 752 -3245
rect 772 -3246 773 -3245
rect 807 -3246 808 -3245
rect 1227 -3246 1228 -3245
rect 1349 -3246 1350 -3245
rect 1353 -3246 1354 -3245
rect 170 -3248 171 -3247
rect 656 -3248 657 -3247
rect 667 -3248 668 -3247
rect 751 -3248 752 -3247
rect 758 -3248 759 -3247
rect 772 -3248 773 -3247
rect 807 -3248 808 -3247
rect 894 -3248 895 -3247
rect 933 -3248 934 -3247
rect 1066 -3248 1067 -3247
rect 1164 -3248 1165 -3247
rect 1234 -3248 1235 -3247
rect 177 -3250 178 -3249
rect 394 -3250 395 -3249
rect 408 -3250 409 -3249
rect 478 -3250 479 -3249
rect 541 -3250 542 -3249
rect 737 -3250 738 -3249
rect 758 -3250 759 -3249
rect 793 -3250 794 -3249
rect 810 -3250 811 -3249
rect 1038 -3250 1039 -3249
rect 1045 -3250 1046 -3249
rect 1258 -3250 1259 -3249
rect 177 -3252 178 -3251
rect 282 -3252 283 -3251
rect 289 -3252 290 -3251
rect 814 -3252 815 -3251
rect 863 -3252 864 -3251
rect 933 -3252 934 -3251
rect 947 -3252 948 -3251
rect 1038 -3252 1039 -3251
rect 1143 -3252 1144 -3251
rect 1164 -3252 1165 -3251
rect 1178 -3252 1179 -3251
rect 1206 -3252 1207 -3251
rect 1220 -3252 1221 -3251
rect 1234 -3252 1235 -3251
rect 187 -3254 188 -3253
rect 254 -3254 255 -3253
rect 282 -3254 283 -3253
rect 296 -3254 297 -3253
rect 317 -3254 318 -3253
rect 366 -3254 367 -3253
rect 408 -3254 409 -3253
rect 436 -3254 437 -3253
rect 450 -3254 451 -3253
rect 579 -3254 580 -3253
rect 618 -3254 619 -3253
rect 744 -3254 745 -3253
rect 765 -3254 766 -3253
rect 786 -3254 787 -3253
rect 793 -3254 794 -3253
rect 828 -3254 829 -3253
rect 863 -3254 864 -3253
rect 884 -3254 885 -3253
rect 891 -3254 892 -3253
rect 1003 -3254 1004 -3253
rect 1024 -3254 1025 -3253
rect 1192 -3254 1193 -3253
rect 1213 -3254 1214 -3253
rect 1220 -3254 1221 -3253
rect 198 -3256 199 -3255
rect 219 -3256 220 -3255
rect 247 -3256 248 -3255
rect 254 -3256 255 -3255
rect 296 -3256 297 -3255
rect 443 -3256 444 -3255
rect 450 -3256 451 -3255
rect 520 -3256 521 -3255
rect 541 -3256 542 -3255
rect 569 -3256 570 -3255
rect 618 -3256 619 -3255
rect 912 -3256 913 -3255
rect 947 -3256 948 -3255
rect 1087 -3256 1088 -3255
rect 1108 -3256 1109 -3255
rect 1143 -3256 1144 -3255
rect 1213 -3256 1214 -3255
rect 1248 -3256 1249 -3255
rect 205 -3258 206 -3257
rect 289 -3258 290 -3257
rect 303 -3258 304 -3257
rect 317 -3258 318 -3257
rect 324 -3258 325 -3257
rect 345 -3258 346 -3257
rect 352 -3258 353 -3257
rect 513 -3258 514 -3257
rect 548 -3258 549 -3257
rect 562 -3258 563 -3257
rect 709 -3258 710 -3257
rect 1024 -3258 1025 -3257
rect 1059 -3258 1060 -3257
rect 1108 -3258 1109 -3257
rect 205 -3260 206 -3259
rect 226 -3260 227 -3259
rect 247 -3260 248 -3259
rect 646 -3260 647 -3259
rect 737 -3260 738 -3259
rect 1272 -3260 1273 -3259
rect 198 -3262 199 -3261
rect 226 -3262 227 -3261
rect 303 -3262 304 -3261
rect 380 -3262 381 -3261
rect 387 -3262 388 -3261
rect 520 -3262 521 -3261
rect 562 -3262 563 -3261
rect 754 -3262 755 -3261
rect 768 -3262 769 -3261
rect 898 -3262 899 -3261
rect 912 -3262 913 -3261
rect 926 -3262 927 -3261
rect 954 -3262 955 -3261
rect 1178 -3262 1179 -3261
rect 191 -3264 192 -3263
rect 380 -3264 381 -3263
rect 387 -3264 388 -3263
rect 779 -3264 780 -3263
rect 786 -3264 787 -3263
rect 919 -3264 920 -3263
rect 954 -3264 955 -3263
rect 1136 -3264 1137 -3263
rect 191 -3266 192 -3265
rect 275 -3266 276 -3265
rect 331 -3266 332 -3265
rect 345 -3266 346 -3265
rect 415 -3266 416 -3265
rect 670 -3266 671 -3265
rect 779 -3266 780 -3265
rect 842 -3266 843 -3265
rect 870 -3266 871 -3265
rect 961 -3266 962 -3265
rect 964 -3266 965 -3265
rect 1185 -3266 1186 -3265
rect 275 -3268 276 -3267
rect 359 -3268 360 -3267
rect 415 -3268 416 -3267
rect 660 -3268 661 -3267
rect 800 -3268 801 -3267
rect 926 -3268 927 -3267
rect 996 -3268 997 -3267
rect 1045 -3268 1046 -3267
rect 1059 -3268 1060 -3267
rect 1073 -3268 1074 -3267
rect 1171 -3268 1172 -3267
rect 1185 -3268 1186 -3267
rect 331 -3270 332 -3269
rect 464 -3270 465 -3269
rect 478 -3270 479 -3269
rect 639 -3270 640 -3269
rect 646 -3270 647 -3269
rect 695 -3270 696 -3269
rect 828 -3270 829 -3269
rect 849 -3270 850 -3269
rect 856 -3270 857 -3269
rect 961 -3270 962 -3269
rect 996 -3270 997 -3269
rect 1031 -3270 1032 -3269
rect 1052 -3270 1053 -3269
rect 1073 -3270 1074 -3269
rect 1157 -3270 1158 -3269
rect 1171 -3270 1172 -3269
rect 184 -3272 185 -3271
rect 695 -3272 696 -3271
rect 842 -3272 843 -3271
rect 968 -3272 969 -3271
rect 982 -3272 983 -3271
rect 1031 -3272 1032 -3271
rect 1052 -3272 1053 -3271
rect 1150 -3272 1151 -3271
rect 184 -3274 185 -3273
rect 233 -3274 234 -3273
rect 310 -3274 311 -3273
rect 464 -3274 465 -3273
rect 485 -3274 486 -3273
rect 569 -3274 570 -3273
rect 614 -3274 615 -3273
rect 898 -3274 899 -3273
rect 919 -3274 920 -3273
rect 975 -3274 976 -3273
rect 982 -3274 983 -3273
rect 989 -3274 990 -3273
rect 1010 -3274 1011 -3273
rect 1248 -3274 1249 -3273
rect 233 -3276 234 -3275
rect 940 -3276 941 -3275
rect 968 -3276 969 -3275
rect 1122 -3276 1123 -3275
rect 1129 -3276 1130 -3275
rect 1150 -3276 1151 -3275
rect 310 -3278 311 -3277
rect 597 -3278 598 -3277
rect 625 -3278 626 -3277
rect 639 -3278 640 -3277
rect 660 -3278 661 -3277
rect 1129 -3278 1130 -3277
rect 359 -3280 360 -3279
rect 590 -3280 591 -3279
rect 625 -3280 626 -3279
rect 691 -3280 692 -3279
rect 821 -3280 822 -3279
rect 975 -3280 976 -3279
rect 989 -3280 990 -3279
rect 1202 -3280 1203 -3279
rect 422 -3282 423 -3281
rect 488 -3282 489 -3281
rect 513 -3282 514 -3281
rect 653 -3282 654 -3281
rect 667 -3282 668 -3281
rect 800 -3282 801 -3281
rect 884 -3282 885 -3281
rect 905 -3282 906 -3281
rect 940 -3282 941 -3281
rect 1003 -3282 1004 -3281
rect 1017 -3282 1018 -3281
rect 1087 -3282 1088 -3281
rect 1115 -3282 1116 -3281
rect 1122 -3282 1123 -3281
rect 422 -3284 423 -3283
rect 555 -3284 556 -3283
rect 583 -3284 584 -3283
rect 597 -3284 598 -3283
rect 653 -3284 654 -3283
rect 859 -3284 860 -3283
rect 877 -3284 878 -3283
rect 905 -3284 906 -3283
rect 1017 -3284 1018 -3283
rect 1080 -3284 1081 -3283
rect 1094 -3284 1095 -3283
rect 1115 -3284 1116 -3283
rect 429 -3286 430 -3285
rect 555 -3286 556 -3285
rect 583 -3286 584 -3285
rect 611 -3286 612 -3285
rect 681 -3286 682 -3285
rect 821 -3286 822 -3285
rect 877 -3286 878 -3285
rect 1262 -3286 1263 -3285
rect 429 -3288 430 -3287
rect 824 -3288 825 -3287
rect 1006 -3288 1007 -3287
rect 1080 -3288 1081 -3287
rect 1262 -3288 1263 -3287
rect 1276 -3288 1277 -3287
rect 436 -3290 437 -3289
rect 492 -3290 493 -3289
rect 534 -3290 535 -3289
rect 590 -3290 591 -3289
rect 611 -3290 612 -3289
rect 891 -3290 892 -3289
rect 1027 -3290 1028 -3289
rect 1157 -3290 1158 -3289
rect 1269 -3290 1270 -3289
rect 1276 -3290 1277 -3289
rect 261 -3292 262 -3291
rect 492 -3292 493 -3291
rect 688 -3292 689 -3291
rect 849 -3292 850 -3291
rect 261 -3294 262 -3293
rect 401 -3294 402 -3293
rect 443 -3294 444 -3293
rect 506 -3294 507 -3293
rect 688 -3294 689 -3293
rect 1010 -3294 1011 -3293
rect 338 -3296 339 -3295
rect 401 -3296 402 -3295
rect 457 -3296 458 -3295
rect 1094 -3296 1095 -3295
rect 338 -3298 339 -3297
rect 471 -3298 472 -3297
rect 485 -3298 486 -3297
rect 723 -3298 724 -3297
rect 457 -3300 458 -3299
rect 604 -3300 605 -3299
rect 716 -3300 717 -3299
rect 723 -3300 724 -3299
rect 471 -3302 472 -3301
rect 537 -3302 538 -3301
rect 604 -3302 605 -3301
rect 835 -3302 836 -3301
rect 506 -3304 507 -3303
rect 674 -3304 675 -3303
rect 716 -3304 717 -3303
rect 730 -3304 731 -3303
rect 674 -3306 675 -3305
rect 873 -3306 874 -3305
rect 156 -3317 157 -3316
rect 271 -3317 272 -3316
rect 303 -3317 304 -3316
rect 485 -3317 486 -3316
rect 520 -3317 521 -3316
rect 558 -3317 559 -3316
rect 576 -3317 577 -3316
rect 614 -3317 615 -3316
rect 653 -3317 654 -3316
rect 849 -3317 850 -3316
rect 856 -3317 857 -3316
rect 1143 -3317 1144 -3316
rect 1181 -3317 1182 -3316
rect 1262 -3317 1263 -3316
rect 1269 -3317 1270 -3316
rect 1290 -3317 1291 -3316
rect 163 -3319 164 -3318
rect 425 -3319 426 -3318
rect 436 -3319 437 -3318
rect 485 -3319 486 -3318
rect 544 -3319 545 -3318
rect 751 -3319 752 -3318
rect 761 -3319 762 -3318
rect 905 -3319 906 -3318
rect 1003 -3319 1004 -3318
rect 1073 -3319 1074 -3318
rect 1136 -3319 1137 -3318
rect 1241 -3319 1242 -3318
rect 1272 -3319 1273 -3318
rect 1276 -3319 1277 -3318
rect 177 -3321 178 -3320
rect 579 -3321 580 -3320
rect 611 -3321 612 -3320
rect 639 -3321 640 -3320
rect 660 -3321 661 -3320
rect 779 -3321 780 -3320
rect 786 -3321 787 -3320
rect 821 -3321 822 -3320
rect 824 -3321 825 -3320
rect 1066 -3321 1067 -3320
rect 1073 -3321 1074 -3320
rect 1150 -3321 1151 -3320
rect 184 -3323 185 -3322
rect 243 -3323 244 -3322
rect 261 -3323 262 -3322
rect 394 -3323 395 -3322
rect 411 -3323 412 -3322
rect 873 -3323 874 -3322
rect 891 -3323 892 -3322
rect 1031 -3323 1032 -3322
rect 1038 -3323 1039 -3322
rect 1041 -3323 1042 -3322
rect 1055 -3323 1056 -3322
rect 1087 -3323 1088 -3322
rect 1139 -3323 1140 -3322
rect 1157 -3323 1158 -3322
rect 198 -3325 199 -3324
rect 219 -3325 220 -3324
rect 226 -3325 227 -3324
rect 240 -3325 241 -3324
rect 282 -3325 283 -3324
rect 303 -3325 304 -3324
rect 359 -3325 360 -3324
rect 667 -3325 668 -3324
rect 670 -3325 671 -3324
rect 1178 -3325 1179 -3324
rect 226 -3327 227 -3326
rect 310 -3327 311 -3326
rect 387 -3327 388 -3326
rect 859 -3327 860 -3326
rect 870 -3327 871 -3326
rect 1192 -3327 1193 -3326
rect 275 -3329 276 -3328
rect 359 -3329 360 -3328
rect 387 -3329 388 -3328
rect 478 -3329 479 -3328
rect 513 -3329 514 -3328
rect 639 -3329 640 -3328
rect 660 -3329 661 -3328
rect 737 -3329 738 -3328
rect 751 -3329 752 -3328
rect 772 -3329 773 -3328
rect 779 -3329 780 -3328
rect 814 -3329 815 -3328
rect 835 -3329 836 -3328
rect 1248 -3329 1249 -3328
rect 275 -3331 276 -3330
rect 345 -3331 346 -3330
rect 394 -3331 395 -3330
rect 506 -3331 507 -3330
rect 513 -3331 514 -3330
rect 653 -3331 654 -3330
rect 667 -3331 668 -3330
rect 723 -3331 724 -3330
rect 737 -3331 738 -3330
rect 765 -3331 766 -3330
rect 807 -3331 808 -3330
rect 814 -3331 815 -3330
rect 835 -3331 836 -3330
rect 926 -3331 927 -3330
rect 947 -3331 948 -3330
rect 1087 -3331 1088 -3330
rect 1192 -3331 1193 -3330
rect 1213 -3331 1214 -3330
rect 282 -3333 283 -3332
rect 296 -3333 297 -3332
rect 310 -3333 311 -3332
rect 317 -3333 318 -3332
rect 345 -3333 346 -3332
rect 373 -3333 374 -3332
rect 422 -3333 423 -3332
rect 537 -3333 538 -3332
rect 569 -3333 570 -3332
rect 772 -3333 773 -3332
rect 838 -3333 839 -3332
rect 1115 -3333 1116 -3332
rect 219 -3335 220 -3334
rect 569 -3335 570 -3334
rect 572 -3335 573 -3334
rect 723 -3335 724 -3334
rect 761 -3335 762 -3334
rect 1045 -3335 1046 -3334
rect 296 -3337 297 -3336
rect 324 -3337 325 -3336
rect 373 -3337 374 -3336
rect 401 -3337 402 -3336
rect 436 -3337 437 -3336
rect 464 -3337 465 -3336
rect 478 -3337 479 -3336
rect 541 -3337 542 -3336
rect 632 -3337 633 -3336
rect 807 -3337 808 -3336
rect 849 -3337 850 -3336
rect 961 -3337 962 -3336
rect 1003 -3337 1004 -3336
rect 1052 -3337 1053 -3336
rect 317 -3339 318 -3338
rect 408 -3339 409 -3338
rect 506 -3339 507 -3338
rect 541 -3339 542 -3338
rect 632 -3339 633 -3338
rect 730 -3339 731 -3338
rect 765 -3339 766 -3338
rect 793 -3339 794 -3338
rect 856 -3339 857 -3338
rect 940 -3339 941 -3338
rect 947 -3339 948 -3338
rect 968 -3339 969 -3338
rect 1024 -3339 1025 -3338
rect 1234 -3339 1235 -3338
rect 324 -3341 325 -3340
rect 471 -3341 472 -3340
rect 534 -3341 535 -3340
rect 786 -3341 787 -3340
rect 870 -3341 871 -3340
rect 1094 -3341 1095 -3340
rect 170 -3343 171 -3342
rect 471 -3343 472 -3342
rect 534 -3343 535 -3342
rect 548 -3343 549 -3342
rect 681 -3343 682 -3342
rect 968 -3343 969 -3342
rect 1027 -3343 1028 -3342
rect 1185 -3343 1186 -3342
rect 331 -3345 332 -3344
rect 793 -3345 794 -3344
rect 884 -3345 885 -3344
rect 1031 -3345 1032 -3344
rect 1045 -3345 1046 -3344
rect 1108 -3345 1109 -3344
rect 1185 -3345 1186 -3344
rect 1199 -3345 1200 -3344
rect 331 -3347 332 -3346
rect 443 -3347 444 -3346
rect 548 -3347 549 -3346
rect 625 -3347 626 -3346
rect 688 -3347 689 -3346
rect 702 -3347 703 -3346
rect 730 -3347 731 -3346
rect 744 -3347 745 -3346
rect 884 -3347 885 -3346
rect 1010 -3347 1011 -3346
rect 1052 -3347 1053 -3346
rect 1255 -3347 1256 -3346
rect 380 -3349 381 -3348
rect 401 -3349 402 -3348
rect 408 -3349 409 -3348
rect 464 -3349 465 -3348
rect 492 -3349 493 -3348
rect 625 -3349 626 -3348
rect 702 -3349 703 -3348
rect 716 -3349 717 -3348
rect 744 -3349 745 -3348
rect 877 -3349 878 -3348
rect 891 -3349 892 -3348
rect 912 -3349 913 -3348
rect 926 -3349 927 -3348
rect 1227 -3349 1228 -3348
rect 380 -3351 381 -3350
rect 499 -3351 500 -3350
rect 597 -3351 598 -3350
rect 681 -3351 682 -3350
rect 691 -3351 692 -3350
rect 716 -3351 717 -3350
rect 877 -3351 878 -3350
rect 982 -3351 983 -3350
rect 1094 -3351 1095 -3350
rect 1122 -3351 1123 -3350
rect 443 -3353 444 -3352
rect 527 -3353 528 -3352
rect 618 -3353 619 -3352
rect 688 -3353 689 -3352
rect 894 -3353 895 -3352
rect 933 -3353 934 -3352
rect 940 -3353 941 -3352
rect 1080 -3353 1081 -3352
rect 1122 -3353 1123 -3352
rect 1220 -3353 1221 -3352
rect 450 -3355 451 -3354
rect 499 -3355 500 -3354
rect 527 -3355 528 -3354
rect 663 -3355 664 -3354
rect 898 -3355 899 -3354
rect 1069 -3355 1070 -3354
rect 1080 -3355 1081 -3354
rect 1101 -3355 1102 -3354
rect 233 -3357 234 -3356
rect 450 -3357 451 -3356
rect 457 -3357 458 -3356
rect 597 -3357 598 -3356
rect 898 -3357 899 -3356
rect 954 -3357 955 -3356
rect 961 -3357 962 -3356
rect 1206 -3357 1207 -3356
rect 233 -3359 234 -3358
rect 338 -3359 339 -3358
rect 422 -3359 423 -3358
rect 457 -3359 458 -3358
rect 492 -3359 493 -3358
rect 604 -3359 605 -3358
rect 758 -3359 759 -3358
rect 954 -3359 955 -3358
rect 975 -3359 976 -3358
rect 1010 -3359 1011 -3358
rect 1017 -3359 1018 -3358
rect 1101 -3359 1102 -3358
rect 338 -3361 339 -3360
rect 562 -3361 563 -3360
rect 576 -3361 577 -3360
rect 604 -3361 605 -3360
rect 674 -3361 675 -3360
rect 975 -3361 976 -3360
rect 982 -3361 983 -3360
rect 1171 -3361 1172 -3360
rect 247 -3363 248 -3362
rect 674 -3363 675 -3362
rect 905 -3363 906 -3362
rect 919 -3363 920 -3362
rect 933 -3363 934 -3362
rect 989 -3363 990 -3362
rect 1013 -3363 1014 -3362
rect 1017 -3363 1018 -3362
rect 191 -3365 192 -3364
rect 247 -3365 248 -3364
rect 352 -3365 353 -3364
rect 562 -3365 563 -3364
rect 583 -3365 584 -3364
rect 618 -3365 619 -3364
rect 912 -3365 913 -3364
rect 996 -3365 997 -3364
rect 352 -3367 353 -3366
rect 555 -3367 556 -3366
rect 583 -3367 584 -3366
rect 709 -3367 710 -3366
rect 800 -3367 801 -3366
rect 996 -3367 997 -3366
rect 415 -3369 416 -3368
rect 555 -3369 556 -3368
rect 590 -3369 591 -3368
rect 709 -3369 710 -3368
rect 800 -3369 801 -3368
rect 863 -3369 864 -3368
rect 919 -3369 920 -3368
rect 1066 -3369 1067 -3368
rect 404 -3371 405 -3370
rect 590 -3371 591 -3370
rect 695 -3371 696 -3370
rect 863 -3371 864 -3370
rect 989 -3371 990 -3370
rect 1059 -3371 1060 -3370
rect 415 -3373 416 -3372
rect 429 -3373 430 -3372
rect 656 -3373 657 -3372
rect 695 -3373 696 -3372
rect 1059 -3373 1060 -3372
rect 1129 -3373 1130 -3372
rect 366 -3375 367 -3374
rect 429 -3375 430 -3374
rect 520 -3375 521 -3374
rect 656 -3375 657 -3374
rect 1129 -3375 1130 -3374
rect 1164 -3375 1165 -3374
rect 289 -3377 290 -3376
rect 366 -3377 367 -3376
rect 268 -3379 269 -3378
rect 289 -3379 290 -3378
rect 198 -3390 199 -3389
rect 292 -3390 293 -3389
rect 296 -3390 297 -3389
rect 446 -3390 447 -3389
rect 457 -3390 458 -3389
rect 460 -3390 461 -3389
rect 492 -3390 493 -3389
rect 656 -3390 657 -3389
rect 723 -3390 724 -3389
rect 758 -3390 759 -3389
rect 793 -3390 794 -3389
rect 870 -3390 871 -3389
rect 1013 -3390 1014 -3389
rect 1087 -3390 1088 -3389
rect 1101 -3390 1102 -3389
rect 1136 -3390 1137 -3389
rect 1178 -3390 1179 -3389
rect 1185 -3390 1186 -3389
rect 1346 -3390 1347 -3389
rect 1349 -3390 1350 -3389
rect 205 -3392 206 -3391
rect 278 -3392 279 -3391
rect 317 -3392 318 -3391
rect 408 -3392 409 -3391
rect 422 -3392 423 -3391
rect 723 -3392 724 -3391
rect 737 -3392 738 -3391
rect 793 -3392 794 -3391
rect 807 -3392 808 -3391
rect 810 -3392 811 -3391
rect 824 -3392 825 -3391
rect 898 -3392 899 -3391
rect 1027 -3392 1028 -3391
rect 1122 -3392 1123 -3391
rect 1181 -3392 1182 -3391
rect 1192 -3392 1193 -3391
rect 1346 -3392 1347 -3391
rect 1353 -3392 1354 -3391
rect 212 -3394 213 -3393
rect 268 -3394 269 -3393
rect 271 -3394 272 -3393
rect 691 -3394 692 -3393
rect 737 -3394 738 -3393
rect 975 -3394 976 -3393
rect 1066 -3394 1067 -3393
rect 1080 -3394 1081 -3393
rect 1087 -3394 1088 -3393
rect 1094 -3394 1095 -3393
rect 1115 -3394 1116 -3393
rect 1129 -3394 1130 -3393
rect 219 -3396 220 -3395
rect 502 -3396 503 -3395
rect 530 -3396 531 -3395
rect 576 -3396 577 -3395
rect 579 -3396 580 -3395
rect 646 -3396 647 -3395
rect 649 -3396 650 -3395
rect 961 -3396 962 -3395
rect 1010 -3396 1011 -3395
rect 1094 -3396 1095 -3395
rect 247 -3398 248 -3397
rect 474 -3398 475 -3397
rect 555 -3398 556 -3397
rect 590 -3398 591 -3397
rect 597 -3398 598 -3397
rect 646 -3398 647 -3397
rect 653 -3398 654 -3397
rect 996 -3398 997 -3397
rect 1010 -3398 1011 -3397
rect 1045 -3398 1046 -3397
rect 240 -3400 241 -3399
rect 247 -3400 248 -3399
rect 261 -3400 262 -3399
rect 289 -3400 290 -3399
rect 324 -3400 325 -3399
rect 348 -3400 349 -3399
rect 366 -3400 367 -3399
rect 404 -3400 405 -3399
rect 408 -3400 409 -3399
rect 429 -3400 430 -3399
rect 450 -3400 451 -3399
rect 492 -3400 493 -3399
rect 558 -3400 559 -3399
rect 590 -3400 591 -3399
rect 667 -3400 668 -3399
rect 758 -3400 759 -3399
rect 807 -3400 808 -3399
rect 877 -3400 878 -3399
rect 933 -3400 934 -3399
rect 975 -3400 976 -3399
rect 1031 -3400 1032 -3399
rect 1045 -3400 1046 -3399
rect 226 -3402 227 -3401
rect 366 -3402 367 -3401
rect 387 -3402 388 -3401
rect 429 -3402 430 -3401
rect 450 -3402 451 -3401
rect 611 -3402 612 -3401
rect 667 -3402 668 -3401
rect 786 -3402 787 -3401
rect 859 -3402 860 -3401
rect 873 -3402 874 -3401
rect 877 -3402 878 -3401
rect 891 -3402 892 -3401
rect 961 -3402 962 -3401
rect 1024 -3402 1025 -3401
rect 1031 -3402 1032 -3401
rect 1059 -3402 1060 -3401
rect 254 -3404 255 -3403
rect 261 -3404 262 -3403
rect 282 -3404 283 -3403
rect 317 -3404 318 -3403
rect 359 -3404 360 -3403
rect 387 -3404 388 -3403
rect 401 -3404 402 -3403
rect 478 -3404 479 -3403
rect 485 -3404 486 -3403
rect 597 -3404 598 -3403
rect 716 -3404 717 -3403
rect 933 -3404 934 -3403
rect 968 -3404 969 -3403
rect 1024 -3404 1025 -3403
rect 303 -3406 304 -3405
rect 324 -3406 325 -3405
rect 345 -3406 346 -3405
rect 359 -3406 360 -3405
rect 415 -3406 416 -3405
rect 422 -3406 423 -3405
rect 457 -3406 458 -3405
rect 527 -3406 528 -3405
rect 548 -3406 549 -3405
rect 611 -3406 612 -3405
rect 716 -3406 717 -3405
rect 772 -3406 773 -3405
rect 786 -3406 787 -3405
rect 800 -3406 801 -3405
rect 863 -3406 864 -3405
rect 887 -3406 888 -3405
rect 968 -3406 969 -3405
rect 989 -3406 990 -3405
rect 233 -3408 234 -3407
rect 345 -3408 346 -3407
rect 373 -3408 374 -3407
rect 415 -3408 416 -3407
rect 478 -3408 479 -3407
rect 506 -3408 507 -3407
rect 541 -3408 542 -3407
rect 548 -3408 549 -3407
rect 569 -3408 570 -3407
rect 618 -3408 619 -3407
rect 660 -3408 661 -3407
rect 772 -3408 773 -3407
rect 800 -3408 801 -3407
rect 814 -3408 815 -3407
rect 863 -3408 864 -3407
rect 919 -3408 920 -3407
rect 1349 -3408 1350 -3407
rect 1353 -3408 1354 -3407
rect 373 -3410 374 -3409
rect 796 -3410 797 -3409
rect 919 -3410 920 -3409
rect 947 -3410 948 -3409
rect 394 -3412 395 -3411
rect 569 -3412 570 -3411
rect 572 -3412 573 -3411
rect 957 -3412 958 -3411
rect 338 -3414 339 -3413
rect 394 -3414 395 -3413
rect 485 -3414 486 -3413
rect 499 -3414 500 -3413
rect 506 -3414 507 -3413
rect 604 -3414 605 -3413
rect 618 -3414 619 -3413
rect 695 -3414 696 -3413
rect 940 -3414 941 -3413
rect 947 -3414 948 -3413
rect 310 -3416 311 -3415
rect 338 -3416 339 -3415
rect 436 -3416 437 -3415
rect 604 -3416 605 -3415
rect 632 -3416 633 -3415
rect 695 -3416 696 -3415
rect 905 -3416 906 -3415
rect 940 -3416 941 -3415
rect 310 -3418 311 -3417
rect 331 -3418 332 -3417
rect 380 -3418 381 -3417
rect 436 -3418 437 -3417
rect 499 -3418 500 -3417
rect 779 -3418 780 -3417
rect 856 -3418 857 -3417
rect 905 -3418 906 -3417
rect 331 -3420 332 -3419
rect 513 -3420 514 -3419
rect 541 -3420 542 -3419
rect 639 -3420 640 -3419
rect 674 -3420 675 -3419
rect 814 -3420 815 -3419
rect 380 -3422 381 -3421
rect 464 -3422 465 -3421
rect 513 -3422 514 -3421
rect 520 -3422 521 -3421
rect 562 -3422 563 -3421
rect 660 -3422 661 -3421
rect 674 -3422 675 -3421
rect 751 -3422 752 -3421
rect 352 -3424 353 -3423
rect 562 -3424 563 -3423
rect 576 -3424 577 -3423
rect 625 -3424 626 -3423
rect 632 -3424 633 -3423
rect 835 -3424 836 -3423
rect 352 -3426 353 -3425
rect 411 -3426 412 -3425
rect 443 -3426 444 -3425
rect 520 -3426 521 -3425
rect 625 -3426 626 -3425
rect 709 -3426 710 -3425
rect 835 -3426 836 -3425
rect 842 -3426 843 -3425
rect 464 -3428 465 -3427
rect 471 -3428 472 -3427
rect 639 -3428 640 -3427
rect 765 -3428 766 -3427
rect 842 -3428 843 -3427
rect 926 -3428 927 -3427
rect 471 -3430 472 -3429
rect 534 -3430 535 -3429
rect 688 -3430 689 -3429
rect 779 -3430 780 -3429
rect 912 -3430 913 -3429
rect 926 -3430 927 -3429
rect 534 -3432 535 -3431
rect 583 -3432 584 -3431
rect 702 -3432 703 -3431
rect 751 -3432 752 -3431
rect 765 -3432 766 -3431
rect 828 -3432 829 -3431
rect 912 -3432 913 -3431
rect 982 -3432 983 -3431
rect 583 -3434 584 -3433
rect 744 -3434 745 -3433
rect 828 -3434 829 -3433
rect 884 -3434 885 -3433
rect 982 -3434 983 -3433
rect 1038 -3434 1039 -3433
rect 702 -3436 703 -3435
rect 730 -3436 731 -3435
rect 744 -3436 745 -3435
rect 1017 -3436 1018 -3435
rect 1038 -3436 1039 -3435
rect 1073 -3436 1074 -3435
rect 709 -3438 710 -3437
rect 821 -3438 822 -3437
rect 884 -3438 885 -3437
rect 954 -3438 955 -3437
rect 730 -3440 731 -3439
rect 849 -3440 850 -3439
rect 740 -3442 741 -3441
rect 849 -3442 850 -3441
rect 275 -3453 276 -3452
rect 289 -3453 290 -3452
rect 292 -3453 293 -3452
rect 310 -3453 311 -3452
rect 331 -3453 332 -3452
rect 366 -3453 367 -3452
rect 380 -3453 381 -3452
rect 383 -3453 384 -3452
rect 464 -3453 465 -3452
rect 467 -3453 468 -3452
rect 513 -3453 514 -3452
rect 579 -3453 580 -3452
rect 611 -3453 612 -3452
rect 649 -3453 650 -3452
rect 677 -3453 678 -3452
rect 957 -3453 958 -3452
rect 989 -3453 990 -3452
rect 1010 -3453 1011 -3452
rect 1045 -3453 1046 -3452
rect 1052 -3453 1053 -3452
rect 1080 -3453 1081 -3452
rect 1087 -3453 1088 -3452
rect 1094 -3453 1095 -3452
rect 1122 -3453 1123 -3452
rect 1136 -3453 1137 -3452
rect 1150 -3453 1151 -3452
rect 1339 -3453 1340 -3452
rect 1342 -3453 1343 -3452
rect 317 -3455 318 -3454
rect 331 -3455 332 -3454
rect 338 -3455 339 -3454
rect 345 -3455 346 -3454
rect 359 -3455 360 -3454
rect 362 -3455 363 -3454
rect 380 -3455 381 -3454
rect 436 -3455 437 -3454
rect 513 -3455 514 -3454
rect 534 -3455 535 -3454
rect 611 -3455 612 -3454
rect 667 -3455 668 -3454
rect 688 -3455 689 -3454
rect 702 -3455 703 -3454
rect 726 -3455 727 -3454
rect 807 -3455 808 -3454
rect 817 -3455 818 -3454
rect 863 -3455 864 -3454
rect 870 -3455 871 -3454
rect 884 -3455 885 -3454
rect 898 -3455 899 -3454
rect 982 -3455 983 -3454
rect 996 -3455 997 -3454
rect 1038 -3455 1039 -3454
rect 1087 -3455 1088 -3454
rect 1171 -3455 1172 -3454
rect 1339 -3455 1340 -3454
rect 1346 -3455 1347 -3454
rect 324 -3457 325 -3456
rect 338 -3457 339 -3456
rect 359 -3457 360 -3456
rect 387 -3457 388 -3456
rect 408 -3457 409 -3456
rect 464 -3457 465 -3456
rect 478 -3457 479 -3456
rect 534 -3457 535 -3456
rect 604 -3457 605 -3456
rect 667 -3457 668 -3456
rect 681 -3457 682 -3456
rect 688 -3457 689 -3456
rect 691 -3457 692 -3456
rect 842 -3457 843 -3456
rect 849 -3457 850 -3456
rect 901 -3457 902 -3456
rect 905 -3457 906 -3456
rect 999 -3457 1000 -3456
rect 1010 -3457 1011 -3456
rect 1031 -3457 1032 -3456
rect 1108 -3457 1109 -3456
rect 1115 -3457 1116 -3456
rect 1346 -3457 1347 -3456
rect 1353 -3457 1354 -3456
rect 408 -3459 409 -3458
rect 450 -3459 451 -3458
rect 478 -3459 479 -3458
rect 548 -3459 549 -3458
rect 597 -3459 598 -3458
rect 604 -3459 605 -3458
rect 628 -3459 629 -3458
rect 1027 -3459 1028 -3458
rect 422 -3461 423 -3460
rect 450 -3461 451 -3460
rect 499 -3461 500 -3460
rect 548 -3461 549 -3460
rect 562 -3461 563 -3460
rect 597 -3461 598 -3460
rect 646 -3461 647 -3460
rect 737 -3461 738 -3460
rect 751 -3461 752 -3460
rect 754 -3461 755 -3460
rect 779 -3461 780 -3460
rect 863 -3461 864 -3460
rect 877 -3461 878 -3460
rect 887 -3461 888 -3460
rect 905 -3461 906 -3460
rect 912 -3461 913 -3460
rect 926 -3461 927 -3460
rect 929 -3461 930 -3460
rect 933 -3461 934 -3460
rect 936 -3461 937 -3460
rect 940 -3461 941 -3460
rect 943 -3461 944 -3460
rect 954 -3461 955 -3460
rect 982 -3461 983 -3460
rect 436 -3463 437 -3462
rect 471 -3463 472 -3462
rect 520 -3463 521 -3462
rect 583 -3463 584 -3462
rect 653 -3463 654 -3462
rect 702 -3463 703 -3462
rect 751 -3463 752 -3462
rect 758 -3463 759 -3462
rect 779 -3463 780 -3462
rect 824 -3463 825 -3462
rect 835 -3463 836 -3462
rect 856 -3463 857 -3462
rect 891 -3463 892 -3462
rect 912 -3463 913 -3462
rect 926 -3463 927 -3462
rect 968 -3463 969 -3462
rect 401 -3465 402 -3464
rect 471 -3465 472 -3464
rect 527 -3465 528 -3464
rect 576 -3465 577 -3464
rect 590 -3465 591 -3464
rect 653 -3465 654 -3464
rect 660 -3465 661 -3464
rect 681 -3465 682 -3464
rect 695 -3465 696 -3464
rect 740 -3465 741 -3464
rect 772 -3465 773 -3464
rect 835 -3465 836 -3464
rect 933 -3465 934 -3464
rect 961 -3465 962 -3464
rect 425 -3467 426 -3466
rect 520 -3467 521 -3466
rect 530 -3467 531 -3466
rect 660 -3467 661 -3466
rect 674 -3467 675 -3466
rect 737 -3467 738 -3466
rect 772 -3467 773 -3466
rect 859 -3467 860 -3466
rect 940 -3467 941 -3466
rect 947 -3467 948 -3466
rect 954 -3467 955 -3466
rect 975 -3467 976 -3466
rect 443 -3469 444 -3468
rect 590 -3469 591 -3468
rect 786 -3469 787 -3468
rect 870 -3469 871 -3468
rect 1342 -3469 1343 -3468
rect 1353 -3469 1354 -3468
rect 443 -3471 444 -3470
rect 457 -3471 458 -3470
rect 506 -3471 507 -3470
rect 527 -3471 528 -3470
rect 562 -3471 563 -3470
rect 618 -3471 619 -3470
rect 793 -3471 794 -3470
rect 821 -3471 822 -3470
rect 828 -3471 829 -3470
rect 856 -3471 857 -3470
rect 422 -3473 423 -3472
rect 506 -3473 507 -3472
rect 618 -3473 619 -3472
rect 625 -3473 626 -3472
rect 723 -3473 724 -3472
rect 821 -3473 822 -3472
rect 446 -3475 447 -3474
rect 499 -3475 500 -3474
rect 583 -3475 584 -3474
rect 625 -3475 626 -3474
rect 800 -3475 801 -3474
rect 842 -3475 843 -3474
rect 457 -3477 458 -3476
rect 485 -3477 486 -3476
rect 709 -3477 710 -3476
rect 800 -3477 801 -3476
rect 807 -3477 808 -3476
rect 1174 -3477 1175 -3476
rect 485 -3479 486 -3478
rect 541 -3479 542 -3478
rect 709 -3479 710 -3478
rect 730 -3479 731 -3478
rect 814 -3479 815 -3478
rect 877 -3479 878 -3478
rect 541 -3481 542 -3480
rect 569 -3481 570 -3480
rect 695 -3481 696 -3480
rect 814 -3481 815 -3480
rect 569 -3483 570 -3482
rect 632 -3483 633 -3482
rect 716 -3483 717 -3482
rect 730 -3483 731 -3482
rect 555 -3485 556 -3484
rect 632 -3485 633 -3484
rect 639 -3485 640 -3484
rect 716 -3485 717 -3484
rect 492 -3487 493 -3486
rect 555 -3487 556 -3486
rect 639 -3487 640 -3486
rect 849 -3487 850 -3486
rect 429 -3489 430 -3488
rect 492 -3489 493 -3488
rect 394 -3491 395 -3490
rect 429 -3491 430 -3490
rect 352 -3493 353 -3492
rect 394 -3493 395 -3492
rect 352 -3495 353 -3494
rect 373 -3495 374 -3494
rect 373 -3497 374 -3496
rect 415 -3497 416 -3496
rect 415 -3499 416 -3498
rect 537 -3499 538 -3498
rect 254 -3510 255 -3509
rect 296 -3510 297 -3509
rect 352 -3510 353 -3509
rect 534 -3510 535 -3509
rect 555 -3510 556 -3509
rect 625 -3510 626 -3509
rect 639 -3510 640 -3509
rect 688 -3510 689 -3509
rect 691 -3510 692 -3509
rect 772 -3510 773 -3509
rect 821 -3510 822 -3509
rect 922 -3510 923 -3509
rect 947 -3510 948 -3509
rect 954 -3510 955 -3509
rect 968 -3510 969 -3509
rect 975 -3510 976 -3509
rect 982 -3510 983 -3509
rect 1006 -3510 1007 -3509
rect 1059 -3510 1060 -3509
rect 1087 -3510 1088 -3509
rect 1122 -3510 1123 -3509
rect 1160 -3510 1161 -3509
rect 1171 -3510 1172 -3509
rect 1178 -3510 1179 -3509
rect 1339 -3510 1340 -3509
rect 1349 -3510 1350 -3509
rect 268 -3512 269 -3511
rect 275 -3512 276 -3511
rect 401 -3512 402 -3511
rect 425 -3512 426 -3511
rect 429 -3512 430 -3511
rect 562 -3512 563 -3511
rect 576 -3512 577 -3511
rect 604 -3512 605 -3511
rect 618 -3512 619 -3511
rect 625 -3512 626 -3511
rect 653 -3512 654 -3511
rect 688 -3512 689 -3511
rect 730 -3512 731 -3511
rect 733 -3512 734 -3511
rect 849 -3512 850 -3511
rect 898 -3512 899 -3511
rect 933 -3512 934 -3511
rect 947 -3512 948 -3511
rect 961 -3512 962 -3511
rect 968 -3512 969 -3511
rect 996 -3512 997 -3511
rect 1010 -3512 1011 -3511
rect 1346 -3512 1347 -3511
rect 1353 -3512 1354 -3511
rect 387 -3514 388 -3513
rect 401 -3514 402 -3513
rect 422 -3514 423 -3513
rect 478 -3514 479 -3513
rect 495 -3514 496 -3513
rect 642 -3514 643 -3513
rect 660 -3514 661 -3513
rect 723 -3514 724 -3513
rect 730 -3514 731 -3513
rect 744 -3514 745 -3513
rect 842 -3514 843 -3513
rect 849 -3514 850 -3513
rect 870 -3514 871 -3513
rect 884 -3514 885 -3513
rect 912 -3514 913 -3513
rect 933 -3514 934 -3513
rect 1003 -3514 1004 -3513
rect 1010 -3514 1011 -3513
rect 373 -3516 374 -3515
rect 422 -3516 423 -3515
rect 429 -3516 430 -3515
rect 604 -3516 605 -3515
rect 667 -3516 668 -3515
rect 726 -3516 727 -3515
rect 737 -3516 738 -3515
rect 744 -3516 745 -3515
rect 856 -3516 857 -3515
rect 870 -3516 871 -3515
rect 877 -3516 878 -3515
rect 891 -3516 892 -3515
rect 912 -3516 913 -3515
rect 926 -3516 927 -3515
rect 450 -3518 451 -3517
rect 492 -3518 493 -3517
rect 499 -3518 500 -3517
rect 534 -3518 535 -3517
rect 548 -3518 549 -3517
rect 576 -3518 577 -3517
rect 590 -3518 591 -3517
rect 639 -3518 640 -3517
rect 667 -3518 668 -3517
rect 807 -3518 808 -3517
rect 863 -3518 864 -3517
rect 877 -3518 878 -3517
rect 919 -3518 920 -3517
rect 926 -3518 927 -3517
rect 394 -3520 395 -3519
rect 450 -3520 451 -3519
rect 453 -3520 454 -3519
rect 478 -3520 479 -3519
rect 485 -3520 486 -3519
rect 492 -3520 493 -3519
rect 499 -3520 500 -3519
rect 565 -3520 566 -3519
rect 597 -3520 598 -3519
rect 628 -3520 629 -3519
rect 674 -3520 675 -3519
rect 681 -3520 682 -3519
rect 733 -3520 734 -3519
rect 737 -3520 738 -3519
rect 835 -3520 836 -3519
rect 863 -3520 864 -3519
rect 359 -3522 360 -3521
rect 394 -3522 395 -3521
rect 457 -3522 458 -3521
rect 548 -3522 549 -3521
rect 555 -3522 556 -3521
rect 569 -3522 570 -3521
rect 600 -3522 601 -3521
rect 646 -3522 647 -3521
rect 677 -3522 678 -3521
rect 943 -3522 944 -3521
rect 338 -3524 339 -3523
rect 359 -3524 360 -3523
rect 408 -3524 409 -3523
rect 457 -3524 458 -3523
rect 513 -3524 514 -3523
rect 562 -3524 563 -3523
rect 569 -3524 570 -3523
rect 583 -3524 584 -3523
rect 632 -3524 633 -3523
rect 681 -3524 682 -3523
rect 800 -3524 801 -3523
rect 835 -3524 836 -3523
rect 408 -3526 409 -3525
rect 464 -3526 465 -3525
rect 467 -3526 468 -3525
rect 583 -3526 584 -3525
rect 443 -3528 444 -3527
rect 513 -3528 514 -3527
rect 520 -3528 521 -3527
rect 579 -3528 580 -3527
rect 366 -3530 367 -3529
rect 443 -3530 444 -3529
rect 464 -3530 465 -3529
rect 544 -3530 545 -3529
rect 436 -3532 437 -3531
rect 520 -3532 521 -3531
rect 527 -3532 528 -3531
rect 590 -3532 591 -3531
rect 415 -3534 416 -3533
rect 436 -3534 437 -3533
rect 527 -3534 528 -3533
rect 541 -3534 542 -3533
rect 380 -3536 381 -3535
rect 415 -3536 416 -3535
rect 541 -3536 542 -3535
rect 695 -3536 696 -3535
rect 345 -3538 346 -3537
rect 380 -3538 381 -3537
rect 695 -3538 696 -3537
rect 716 -3538 717 -3537
rect 331 -3540 332 -3539
rect 345 -3540 346 -3539
rect 716 -3540 717 -3539
rect 779 -3540 780 -3539
rect 247 -3551 248 -3550
rect 257 -3551 258 -3550
rect 296 -3551 297 -3550
rect 310 -3551 311 -3550
rect 327 -3551 328 -3550
rect 366 -3551 367 -3550
rect 394 -3551 395 -3550
rect 432 -3551 433 -3550
rect 457 -3551 458 -3550
rect 600 -3551 601 -3550
rect 604 -3551 605 -3550
rect 646 -3551 647 -3550
rect 677 -3551 678 -3550
rect 940 -3551 941 -3550
rect 1006 -3551 1007 -3550
rect 1010 -3551 1011 -3550
rect 1038 -3551 1039 -3550
rect 1059 -3551 1060 -3550
rect 1080 -3551 1081 -3550
rect 1087 -3551 1088 -3550
rect 1150 -3551 1151 -3550
rect 1157 -3551 1158 -3550
rect 345 -3553 346 -3552
rect 352 -3553 353 -3552
rect 380 -3553 381 -3552
rect 394 -3553 395 -3552
rect 443 -3553 444 -3552
rect 457 -3553 458 -3552
rect 485 -3553 486 -3552
rect 506 -3553 507 -3552
rect 544 -3553 545 -3552
rect 576 -3553 577 -3552
rect 583 -3553 584 -3552
rect 597 -3553 598 -3552
rect 618 -3553 619 -3552
rect 667 -3553 668 -3552
rect 681 -3553 682 -3552
rect 688 -3553 689 -3552
rect 695 -3553 696 -3552
rect 698 -3553 699 -3552
rect 723 -3553 724 -3552
rect 726 -3553 727 -3552
rect 849 -3553 850 -3552
rect 856 -3553 857 -3552
rect 870 -3553 871 -3552
rect 901 -3553 902 -3552
rect 912 -3553 913 -3552
rect 919 -3553 920 -3552
rect 933 -3553 934 -3552
rect 947 -3553 948 -3552
rect 488 -3555 489 -3554
rect 534 -3555 535 -3554
rect 562 -3555 563 -3554
rect 628 -3555 629 -3554
rect 639 -3555 640 -3554
rect 660 -3555 661 -3554
rect 695 -3555 696 -3554
rect 702 -3555 703 -3554
rect 723 -3555 724 -3554
rect 730 -3555 731 -3554
rect 835 -3555 836 -3554
rect 849 -3555 850 -3554
rect 863 -3555 864 -3554
rect 919 -3555 920 -3554
rect 450 -3557 451 -3556
rect 562 -3557 563 -3556
rect 702 -3557 703 -3556
rect 716 -3557 717 -3556
rect 730 -3557 731 -3556
rect 737 -3557 738 -3556
rect 884 -3557 885 -3556
rect 922 -3557 923 -3556
rect 450 -3559 451 -3558
rect 453 -3559 454 -3558
rect 464 -3559 465 -3558
rect 488 -3559 489 -3558
rect 492 -3559 493 -3558
rect 534 -3559 535 -3558
rect 709 -3559 710 -3558
rect 716 -3559 717 -3558
rect 737 -3559 738 -3558
rect 751 -3559 752 -3558
rect 891 -3559 892 -3558
rect 912 -3559 913 -3558
rect 436 -3561 437 -3560
rect 464 -3561 465 -3560
rect 478 -3561 479 -3560
rect 492 -3561 493 -3560
rect 499 -3561 500 -3560
rect 506 -3561 507 -3560
rect 751 -3561 752 -3560
rect 758 -3561 759 -3560
rect 877 -3561 878 -3560
rect 891 -3561 892 -3560
rect 898 -3561 899 -3560
rect 982 -3561 983 -3560
rect 415 -3563 416 -3562
rect 436 -3563 437 -3562
rect 471 -3563 472 -3562
rect 499 -3563 500 -3562
rect 744 -3563 745 -3562
rect 758 -3563 759 -3562
rect 408 -3565 409 -3564
rect 415 -3565 416 -3564
rect 422 -3565 423 -3564
rect 471 -3565 472 -3564
rect 478 -3565 479 -3564
rect 541 -3565 542 -3564
rect 726 -3565 727 -3564
rect 744 -3565 745 -3564
rect 376 -3567 377 -3566
rect 408 -3567 409 -3566
rect 541 -3567 542 -3566
rect 555 -3567 556 -3566
rect 555 -3569 556 -3568
rect 569 -3569 570 -3568
rect 548 -3571 549 -3570
rect 569 -3571 570 -3570
rect 527 -3573 528 -3572
rect 548 -3573 549 -3572
rect 513 -3575 514 -3574
rect 527 -3575 528 -3574
rect 513 -3577 514 -3576
rect 590 -3577 591 -3576
rect 264 -3588 265 -3587
rect 268 -3588 269 -3587
rect 310 -3588 311 -3587
rect 327 -3588 328 -3587
rect 359 -3588 360 -3587
rect 376 -3588 377 -3587
rect 394 -3588 395 -3587
rect 401 -3588 402 -3587
rect 408 -3588 409 -3587
rect 446 -3588 447 -3587
rect 450 -3588 451 -3587
rect 457 -3588 458 -3587
rect 492 -3588 493 -3587
rect 516 -3588 517 -3587
rect 520 -3588 521 -3587
rect 544 -3588 545 -3587
rect 562 -3588 563 -3587
rect 677 -3588 678 -3587
rect 751 -3588 752 -3587
rect 754 -3588 755 -3587
rect 758 -3588 759 -3587
rect 772 -3588 773 -3587
rect 849 -3588 850 -3587
rect 863 -3588 864 -3587
rect 905 -3588 906 -3587
rect 908 -3588 909 -3587
rect 912 -3588 913 -3587
rect 919 -3588 920 -3587
rect 940 -3588 941 -3587
rect 1045 -3588 1046 -3587
rect 1083 -3588 1084 -3587
rect 1087 -3588 1088 -3587
rect 324 -3590 325 -3589
rect 327 -3590 328 -3589
rect 366 -3590 367 -3589
rect 404 -3590 405 -3589
rect 408 -3590 409 -3589
rect 415 -3590 416 -3589
rect 436 -3590 437 -3589
rect 457 -3590 458 -3589
rect 471 -3590 472 -3589
rect 492 -3590 493 -3589
rect 506 -3590 507 -3589
rect 520 -3590 521 -3589
rect 534 -3590 535 -3589
rect 562 -3590 563 -3589
rect 569 -3590 570 -3589
rect 576 -3590 577 -3589
rect 597 -3590 598 -3589
rect 604 -3590 605 -3589
rect 611 -3590 612 -3589
rect 614 -3590 615 -3589
rect 646 -3590 647 -3589
rect 681 -3590 682 -3589
rect 744 -3590 745 -3589
rect 758 -3590 759 -3589
rect 891 -3590 892 -3589
rect 905 -3590 906 -3589
rect 968 -3590 969 -3589
rect 982 -3590 983 -3589
rect 985 -3590 986 -3589
rect 989 -3590 990 -3589
rect 1031 -3590 1032 -3589
rect 1038 -3590 1039 -3589
rect 443 -3592 444 -3591
rect 478 -3592 479 -3591
rect 499 -3592 500 -3591
rect 506 -3592 507 -3591
rect 516 -3592 517 -3591
rect 541 -3592 542 -3591
rect 548 -3592 549 -3591
rect 569 -3592 570 -3591
rect 597 -3592 598 -3591
rect 618 -3592 619 -3591
rect 660 -3592 661 -3591
rect 674 -3592 675 -3591
rect 737 -3592 738 -3591
rect 744 -3592 745 -3591
rect 751 -3592 752 -3591
rect 765 -3592 766 -3591
rect 975 -3592 976 -3591
rect 982 -3592 983 -3591
rect 464 -3594 465 -3593
rect 471 -3594 472 -3593
rect 548 -3594 549 -3593
rect 555 -3594 556 -3593
rect 730 -3594 731 -3593
rect 737 -3594 738 -3593
rect 754 -3594 755 -3593
rect 765 -3594 766 -3593
rect 901 -3594 902 -3593
rect 975 -3594 976 -3593
rect 527 -3596 528 -3595
rect 555 -3596 556 -3595
rect 723 -3596 724 -3595
rect 730 -3596 731 -3595
rect 709 -3598 710 -3597
rect 723 -3598 724 -3597
rect 688 -3600 689 -3599
rect 709 -3600 710 -3599
rect 401 -3611 402 -3610
rect 404 -3611 405 -3610
rect 457 -3611 458 -3610
rect 464 -3611 465 -3610
rect 492 -3611 493 -3610
rect 513 -3611 514 -3610
rect 520 -3611 521 -3610
rect 527 -3611 528 -3610
rect 541 -3611 542 -3610
rect 548 -3611 549 -3610
rect 555 -3611 556 -3610
rect 583 -3611 584 -3610
rect 590 -3611 591 -3610
rect 597 -3611 598 -3610
rect 604 -3611 605 -3610
rect 611 -3611 612 -3610
rect 684 -3611 685 -3610
rect 800 -3611 801 -3610
rect 926 -3611 927 -3610
rect 933 -3611 934 -3610
rect 975 -3611 976 -3610
rect 1003 -3611 1004 -3610
rect 1045 -3611 1046 -3610
rect 1080 -3611 1081 -3610
rect 401 -3613 402 -3612
rect 408 -3613 409 -3612
rect 506 -3613 507 -3612
rect 516 -3613 517 -3612
rect 709 -3613 710 -3612
rect 712 -3613 713 -3612
rect 730 -3613 731 -3612
rect 775 -3613 776 -3612
rect 919 -3613 920 -3612
rect 926 -3613 927 -3612
rect 1052 -3613 1053 -3612
rect 1059 -3613 1060 -3612
rect 709 -3615 710 -3614
rect 716 -3615 717 -3614
rect 751 -3615 752 -3614
rect 761 -3615 762 -3614
rect 712 -3617 713 -3616
rect 716 -3617 717 -3616
rect 737 -3617 738 -3616
rect 751 -3617 752 -3616
rect 758 -3617 759 -3616
rect 765 -3617 766 -3616
rect 744 -3619 745 -3618
rect 758 -3619 759 -3618
rect 765 -3619 766 -3618
rect 772 -3619 773 -3618
rect 723 -3621 724 -3620
rect 744 -3621 745 -3620
rect 702 -3623 703 -3622
rect 723 -3623 724 -3622
rect 695 -3625 696 -3624
rect 702 -3625 703 -3624
rect 471 -3636 472 -3635
rect 474 -3636 475 -3635
rect 562 -3636 563 -3635
rect 572 -3636 573 -3635
rect 583 -3636 584 -3635
rect 597 -3636 598 -3635
rect 719 -3636 720 -3635
rect 723 -3636 724 -3635
rect 744 -3636 745 -3635
rect 772 -3636 773 -3635
rect 856 -3636 857 -3635
rect 859 -3636 860 -3635
rect 926 -3636 927 -3635
rect 929 -3636 930 -3635
rect 982 -3636 983 -3635
rect 989 -3636 990 -3635
rect 1031 -3636 1032 -3635
rect 1034 -3636 1035 -3635
rect 1055 -3636 1056 -3635
rect 1059 -3636 1060 -3635
rect 1080 -3636 1081 -3635
rect 1094 -3636 1095 -3635
rect 1108 -3636 1109 -3635
rect 1111 -3636 1112 -3635
rect 576 -3638 577 -3637
rect 583 -3638 584 -3637
rect 709 -3638 710 -3637
rect 723 -3638 724 -3637
rect 800 -3638 801 -3637
rect 926 -3638 927 -3637
rect 985 -3638 986 -3637
rect 1052 -3638 1053 -3637
rect 569 -3640 570 -3639
rect 576 -3640 577 -3639
rect 702 -3640 703 -3639
rect 709 -3640 710 -3639
rect 1003 -3640 1004 -3639
rect 1031 -3640 1032 -3639
rect 464 -3651 465 -3650
rect 474 -3651 475 -3650
rect 527 -3651 528 -3650
rect 534 -3651 535 -3650
rect 569 -3651 570 -3650
rect 576 -3651 577 -3650
rect 583 -3651 584 -3650
rect 590 -3651 591 -3650
rect 709 -3651 710 -3650
rect 719 -3651 720 -3650
rect 765 -3651 766 -3650
rect 772 -3651 773 -3650
rect 856 -3651 857 -3650
rect 863 -3651 864 -3650
rect 929 -3651 930 -3650
rect 933 -3651 934 -3650
rect 985 -3651 986 -3650
rect 989 -3651 990 -3650
rect 1094 -3651 1095 -3650
rect 1108 -3651 1109 -3650
rect 586 -3653 587 -3652
rect 597 -3653 598 -3652
rect 716 -3653 717 -3652
rect 723 -3653 724 -3652
rect 758 -3653 759 -3652
rect 765 -3653 766 -3652
rect 751 -3655 752 -3654
rect 758 -3655 759 -3654
rect 404 -3666 405 -3665
rect 408 -3666 409 -3665
rect 527 -3666 528 -3665
rect 534 -3666 535 -3665
rect 758 -3666 759 -3665
rect 765 -3666 766 -3665
rect 768 -3666 769 -3665
rect 772 -3666 773 -3665
<< metal2 >>
rect 226 -7 227 1
rect 331 -7 332 1
rect 366 -7 367 1
rect 404 -7 405 1
rect 415 -7 416 1
rect 562 -7 563 1
rect 590 -7 591 1
rect 642 -7 643 1
rect 667 -7 668 1
rect 674 -7 675 1
rect 705 -7 706 1
rect 828 -7 829 1
rect 254 -7 255 -1
rect 380 -7 381 -1
rect 401 -7 402 -1
rect 450 -7 451 -1
rect 457 -7 458 -1
rect 471 -7 472 -1
rect 492 -7 493 -1
rect 537 -7 538 -1
rect 765 -7 766 -1
rect 800 -7 801 -1
rect 803 -7 804 -1
rect 842 -7 843 -1
rect 275 -7 276 -3
rect 460 -7 461 -3
rect 506 -7 507 -3
rect 513 -7 514 -3
rect 516 -7 517 -3
rect 527 -7 528 -3
rect 534 -7 535 -3
rect 569 -7 570 -3
rect 317 -7 318 -5
rect 373 -7 374 -5
rect 429 -7 430 -5
rect 436 -7 437 -5
rect 135 -36 136 -16
rect 222 -36 223 -16
rect 303 -36 304 -16
rect 317 -17 318 -15
rect 327 -36 328 -16
rect 380 -36 381 -16
rect 383 -17 384 -15
rect 534 -36 535 -16
rect 541 -17 542 -15
rect 548 -36 549 -16
rect 565 -17 566 -15
rect 709 -36 710 -16
rect 765 -17 766 -15
rect 765 -36 766 -16
rect 765 -17 766 -15
rect 765 -36 766 -16
rect 775 -36 776 -16
rect 800 -36 801 -16
rect 821 -36 822 -16
rect 919 -36 920 -16
rect 191 -36 192 -18
rect 226 -19 227 -15
rect 310 -36 311 -18
rect 338 -36 339 -18
rect 345 -36 346 -18
rect 366 -19 367 -15
rect 373 -36 374 -18
rect 443 -19 444 -15
rect 450 -19 451 -15
rect 520 -36 521 -18
rect 527 -19 528 -15
rect 541 -36 542 -18
rect 569 -19 570 -15
rect 583 -36 584 -18
rect 632 -36 633 -18
rect 667 -36 668 -18
rect 674 -19 675 -15
rect 695 -36 696 -18
rect 782 -36 783 -18
rect 793 -36 794 -18
rect 828 -19 829 -15
rect 877 -36 878 -18
rect 205 -36 206 -20
rect 254 -21 255 -15
rect 331 -21 332 -15
rect 478 -36 479 -20
rect 488 -36 489 -20
rect 555 -36 556 -20
rect 569 -36 570 -20
rect 705 -21 706 -15
rect 842 -21 843 -15
rect 856 -36 857 -20
rect 212 -36 213 -22
rect 275 -23 276 -15
rect 331 -36 332 -22
rect 404 -36 405 -22
rect 408 -36 409 -22
rect 464 -36 465 -22
rect 471 -23 472 -15
rect 471 -36 472 -22
rect 471 -23 472 -15
rect 471 -36 472 -22
rect 492 -23 493 -15
rect 492 -36 493 -22
rect 492 -23 493 -15
rect 492 -36 493 -22
rect 506 -23 507 -15
rect 513 -36 514 -22
rect 576 -36 577 -22
rect 590 -23 591 -15
rect 635 -36 636 -22
rect 653 -36 654 -22
rect 660 -36 661 -22
rect 761 -36 762 -22
rect 226 -36 227 -24
rect 296 -36 297 -24
rect 352 -36 353 -24
rect 415 -25 416 -15
rect 436 -25 437 -15
rect 446 -25 447 -15
rect 450 -36 451 -24
rect 527 -36 528 -24
rect 639 -25 640 -15
rect 702 -36 703 -24
rect 254 -36 255 -26
rect 366 -36 367 -26
rect 376 -27 377 -15
rect 422 -36 423 -26
rect 443 -36 444 -26
rect 684 -36 685 -26
rect 299 -36 300 -28
rect 415 -36 416 -28
rect 457 -29 458 -15
rect 646 -36 647 -28
rect 317 -36 318 -30
rect 446 -36 447 -30
rect 618 -31 619 -15
rect 639 -36 640 -30
rect 387 -36 388 -32
rect 394 -33 395 -15
rect 401 -36 402 -32
rect 457 -36 458 -32
rect 618 -36 619 -32
rect 786 -36 787 -32
rect 359 -36 360 -34
rect 394 -36 395 -34
rect 79 -85 80 -45
rect 236 -46 237 -44
rect 268 -85 269 -45
rect 331 -46 332 -44
rect 345 -46 346 -44
rect 345 -85 346 -45
rect 345 -46 346 -44
rect 345 -85 346 -45
rect 380 -46 381 -44
rect 446 -85 447 -45
rect 450 -46 451 -44
rect 604 -85 605 -45
rect 618 -46 619 -44
rect 807 -85 808 -45
rect 856 -46 857 -44
rect 863 -85 864 -45
rect 877 -46 878 -44
rect 905 -85 906 -45
rect 919 -46 920 -44
rect 968 -85 969 -45
rect 100 -85 101 -47
rect 135 -48 136 -44
rect 142 -85 143 -47
rect 327 -48 328 -44
rect 380 -85 381 -47
rect 572 -85 573 -47
rect 576 -48 577 -44
rect 597 -85 598 -47
rect 632 -85 633 -47
rect 653 -48 654 -44
rect 667 -48 668 -44
rect 723 -85 724 -47
rect 758 -85 759 -47
rect 870 -85 871 -47
rect 128 -85 129 -49
rect 236 -85 237 -49
rect 278 -85 279 -49
rect 303 -50 304 -44
rect 310 -50 311 -44
rect 310 -85 311 -49
rect 310 -50 311 -44
rect 310 -85 311 -49
rect 324 -85 325 -49
rect 474 -85 475 -49
rect 478 -50 479 -44
rect 611 -85 612 -49
rect 639 -50 640 -44
rect 688 -85 689 -49
rect 695 -50 696 -44
rect 751 -85 752 -49
rect 761 -50 762 -44
rect 891 -85 892 -49
rect 149 -85 150 -51
rect 317 -52 318 -44
rect 397 -52 398 -44
rect 401 -85 402 -51
rect 408 -52 409 -44
rect 506 -85 507 -51
rect 541 -52 542 -44
rect 562 -85 563 -51
rect 576 -85 577 -51
rect 583 -52 584 -44
rect 590 -52 591 -44
rect 653 -85 654 -51
rect 660 -52 661 -44
rect 667 -85 668 -51
rect 702 -52 703 -44
rect 744 -85 745 -51
rect 765 -52 766 -44
rect 772 -85 773 -51
rect 786 -52 787 -44
rect 856 -85 857 -51
rect 156 -85 157 -53
rect 254 -54 255 -44
rect 289 -85 290 -53
rect 366 -54 367 -44
rect 422 -54 423 -44
rect 467 -54 468 -44
rect 485 -85 486 -53
rect 642 -85 643 -53
rect 702 -85 703 -53
rect 824 -54 825 -44
rect 163 -85 164 -55
rect 180 -56 181 -44
rect 184 -85 185 -55
rect 191 -56 192 -44
rect 219 -85 220 -55
rect 453 -56 454 -44
rect 464 -56 465 -44
rect 695 -85 696 -55
rect 709 -56 710 -44
rect 786 -85 787 -55
rect 793 -56 794 -44
rect 814 -85 815 -55
rect 170 -85 171 -57
rect 296 -58 297 -44
rect 303 -85 304 -57
rect 359 -58 360 -44
rect 366 -85 367 -57
rect 478 -85 479 -57
rect 499 -85 500 -57
rect 569 -58 570 -44
rect 625 -85 626 -57
rect 765 -85 766 -57
rect 800 -58 801 -44
rect 821 -85 822 -57
rect 177 -60 178 -44
rect 198 -85 199 -59
rect 222 -60 223 -44
rect 359 -85 360 -59
rect 415 -60 416 -44
rect 422 -85 423 -59
rect 436 -85 437 -59
rect 471 -60 472 -44
rect 520 -60 521 -44
rect 709 -85 710 -59
rect 177 -85 178 -61
rect 464 -85 465 -61
rect 527 -62 528 -44
rect 541 -85 542 -61
rect 555 -62 556 -44
rect 716 -85 717 -61
rect 180 -85 181 -63
rect 205 -64 206 -44
rect 226 -64 227 -44
rect 254 -85 255 -63
rect 261 -85 262 -63
rect 296 -85 297 -63
rect 317 -85 318 -63
rect 352 -64 353 -44
rect 369 -64 370 -44
rect 520 -85 521 -63
rect 527 -85 528 -63
rect 740 -85 741 -63
rect 191 -85 192 -65
rect 212 -66 213 -44
rect 226 -85 227 -65
rect 583 -85 584 -65
rect 646 -66 647 -44
rect 800 -85 801 -65
rect 205 -85 206 -67
rect 373 -68 374 -44
rect 415 -85 416 -67
rect 457 -68 458 -44
rect 534 -68 535 -44
rect 660 -85 661 -67
rect 681 -68 682 -44
rect 793 -85 794 -67
rect 229 -85 230 -69
rect 429 -85 430 -69
rect 450 -85 451 -69
rect 488 -70 489 -44
rect 513 -70 514 -44
rect 534 -85 535 -69
rect 548 -70 549 -44
rect 555 -85 556 -69
rect 569 -85 570 -69
rect 618 -85 619 -69
rect 646 -85 647 -69
rect 782 -85 783 -69
rect 243 -85 244 -71
rect 352 -85 353 -71
rect 369 -85 370 -71
rect 779 -85 780 -71
rect 331 -85 332 -73
rect 681 -85 682 -73
rect 338 -76 339 -44
rect 408 -85 409 -75
rect 457 -85 458 -75
rect 628 -85 629 -75
rect 338 -85 339 -77
rect 621 -78 622 -44
rect 373 -85 374 -79
rect 387 -80 388 -44
rect 492 -80 493 -44
rect 513 -85 514 -79
rect 548 -85 549 -79
rect 593 -80 594 -44
rect 492 -85 493 -81
rect 733 -85 734 -81
rect 593 -85 594 -83
rect 674 -85 675 -83
rect 79 -95 80 -93
rect 390 -156 391 -94
rect 418 -156 419 -94
rect 758 -156 759 -94
rect 814 -95 815 -93
rect 849 -156 850 -94
rect 856 -95 857 -93
rect 919 -156 920 -94
rect 940 -156 941 -94
rect 975 -156 976 -94
rect 114 -97 115 -93
rect 338 -97 339 -93
rect 352 -97 353 -93
rect 394 -156 395 -96
rect 432 -156 433 -96
rect 709 -97 710 -93
rect 730 -97 731 -93
rect 772 -97 773 -93
rect 842 -156 843 -96
rect 947 -156 948 -96
rect 968 -97 969 -93
rect 1003 -156 1004 -96
rect 100 -99 101 -93
rect 114 -156 115 -98
rect 128 -99 129 -93
rect 226 -99 227 -93
rect 250 -156 251 -98
rect 730 -156 731 -98
rect 744 -99 745 -93
rect 835 -156 836 -98
rect 870 -99 871 -93
rect 954 -156 955 -98
rect 100 -156 101 -100
rect 117 -101 118 -93
rect 149 -101 150 -93
rect 334 -101 335 -93
rect 352 -156 353 -100
rect 415 -101 416 -93
rect 443 -101 444 -93
rect 709 -156 710 -100
rect 744 -156 745 -100
rect 786 -101 787 -93
rect 863 -101 864 -93
rect 870 -156 871 -100
rect 891 -101 892 -93
rect 961 -156 962 -100
rect 156 -103 157 -93
rect 236 -103 237 -93
rect 240 -103 241 -93
rect 443 -156 444 -102
rect 446 -103 447 -93
rect 548 -103 549 -93
rect 558 -156 559 -102
rect 968 -156 969 -102
rect 163 -105 164 -93
rect 163 -156 164 -104
rect 163 -105 164 -93
rect 163 -156 164 -104
rect 205 -105 206 -93
rect 338 -156 339 -104
rect 453 -105 454 -93
rect 716 -105 717 -93
rect 723 -105 724 -93
rect 863 -156 864 -104
rect 905 -105 906 -93
rect 926 -156 927 -104
rect 205 -156 206 -106
rect 275 -107 276 -93
rect 282 -107 283 -93
rect 310 -107 311 -93
rect 324 -107 325 -93
rect 327 -125 328 -106
rect 506 -107 507 -93
rect 779 -156 780 -106
rect 793 -107 794 -93
rect 905 -156 906 -106
rect 149 -156 150 -108
rect 275 -156 276 -108
rect 292 -156 293 -108
rect 408 -109 409 -93
rect 499 -109 500 -93
rect 506 -156 507 -108
rect 513 -109 514 -93
rect 625 -156 626 -108
rect 642 -109 643 -93
rect 828 -156 829 -108
rect 145 -111 146 -93
rect 408 -156 409 -110
rect 513 -156 514 -110
rect 684 -156 685 -110
rect 688 -111 689 -93
rect 814 -156 815 -110
rect 821 -111 822 -93
rect 891 -156 892 -110
rect 170 -113 171 -93
rect 282 -156 283 -112
rect 296 -113 297 -93
rect 415 -156 416 -112
rect 562 -113 563 -93
rect 639 -156 640 -112
rect 646 -113 647 -93
rect 649 -113 650 -93
rect 660 -113 661 -93
rect 982 -156 983 -112
rect 170 -156 171 -114
rect 467 -156 468 -114
rect 485 -115 486 -93
rect 562 -156 563 -114
rect 569 -115 570 -93
rect 933 -156 934 -114
rect 215 -117 216 -93
rect 226 -156 227 -116
rect 268 -117 269 -93
rect 299 -117 300 -93
rect 303 -117 304 -93
rect 366 -117 367 -93
rect 569 -156 570 -116
rect 632 -117 633 -93
rect 646 -156 647 -116
rect 653 -117 654 -93
rect 660 -156 661 -116
rect 740 -117 741 -93
rect 751 -117 752 -93
rect 898 -156 899 -116
rect 177 -119 178 -93
rect 299 -156 300 -118
rect 310 -156 311 -118
rect 317 -119 318 -93
rect 324 -156 325 -118
rect 471 -119 472 -93
rect 632 -156 633 -118
rect 653 -156 654 -118
rect 807 -119 808 -93
rect 177 -156 178 -120
rect 261 -121 262 -93
rect 268 -156 269 -120
rect 303 -156 304 -120
rect 359 -121 360 -93
rect 499 -156 500 -120
rect 548 -156 549 -120
rect 751 -156 752 -120
rect 754 -156 755 -120
rect 821 -156 822 -120
rect 191 -123 192 -93
rect 261 -156 262 -122
rect 278 -123 279 -93
rect 296 -156 297 -122
rect 345 -123 346 -93
rect 359 -156 360 -122
rect 471 -156 472 -122
rect 611 -123 612 -93
rect 618 -123 619 -93
rect 884 -156 885 -122
rect 142 -125 143 -93
rect 345 -156 346 -124
rect 450 -125 451 -93
rect 618 -156 619 -124
rect 649 -156 650 -124
rect 807 -156 808 -124
rect 184 -127 185 -93
rect 191 -156 192 -126
rect 212 -127 213 -93
rect 366 -156 367 -126
rect 436 -127 437 -93
rect 450 -156 451 -126
rect 534 -127 535 -93
rect 611 -156 612 -126
rect 667 -127 668 -93
rect 989 -156 990 -126
rect 184 -156 185 -128
rect 474 -156 475 -128
rect 555 -129 556 -93
rect 667 -156 668 -128
rect 674 -129 675 -93
rect 772 -156 773 -128
rect 198 -131 199 -93
rect 212 -156 213 -130
rect 254 -131 255 -93
rect 317 -156 318 -130
rect 457 -131 458 -93
rect 534 -156 535 -130
rect 583 -131 584 -93
rect 877 -156 878 -130
rect 198 -156 199 -132
rect 219 -133 220 -93
rect 240 -156 241 -132
rect 254 -156 255 -132
rect 285 -133 286 -93
rect 436 -156 437 -132
rect 457 -156 458 -132
rect 509 -156 510 -132
rect 583 -156 584 -132
rect 604 -133 605 -93
rect 674 -156 675 -132
rect 761 -133 762 -93
rect 765 -133 766 -93
rect 786 -156 787 -132
rect 219 -156 220 -134
rect 271 -156 272 -134
rect 285 -156 286 -134
rect 331 -156 332 -134
rect 492 -135 493 -93
rect 604 -156 605 -134
rect 688 -156 689 -134
rect 702 -135 703 -93
rect 716 -156 717 -134
rect 800 -135 801 -93
rect 422 -137 423 -93
rect 492 -156 493 -136
rect 520 -137 521 -93
rect 800 -156 801 -136
rect 401 -139 402 -93
rect 422 -156 423 -138
rect 520 -156 521 -138
rect 527 -139 528 -93
rect 590 -139 591 -93
rect 681 -139 682 -93
rect 695 -139 696 -93
rect 912 -156 913 -138
rect 373 -141 374 -93
rect 401 -156 402 -140
rect 429 -141 430 -93
rect 527 -156 528 -140
rect 597 -141 598 -93
rect 723 -156 724 -140
rect 289 -143 290 -93
rect 373 -156 374 -142
rect 429 -156 430 -142
rect 793 -156 794 -142
rect 233 -156 234 -144
rect 289 -156 290 -144
rect 478 -145 479 -93
rect 590 -156 591 -144
rect 681 -156 682 -144
rect 765 -156 766 -144
rect 478 -156 479 -146
rect 576 -147 577 -93
rect 702 -156 703 -146
rect 737 -156 738 -146
rect 464 -149 465 -93
rect 576 -156 577 -148
rect 464 -156 465 -150
rect 856 -156 857 -150
rect 541 -153 542 -93
rect 597 -156 598 -152
rect 488 -156 489 -154
rect 541 -156 542 -154
rect 72 -251 73 -165
rect 432 -166 433 -164
rect 450 -166 451 -164
rect 481 -251 482 -165
rect 495 -251 496 -165
rect 590 -166 591 -164
rect 618 -166 619 -164
rect 863 -166 864 -164
rect 870 -166 871 -164
rect 940 -251 941 -165
rect 954 -166 955 -164
rect 1087 -251 1088 -165
rect 100 -168 101 -164
rect 128 -251 129 -167
rect 135 -251 136 -167
rect 352 -168 353 -164
rect 390 -168 391 -164
rect 436 -168 437 -164
rect 453 -251 454 -167
rect 527 -168 528 -164
rect 541 -168 542 -164
rect 555 -251 556 -167
rect 618 -251 619 -167
rect 716 -168 717 -164
rect 730 -168 731 -164
rect 1122 -251 1123 -167
rect 100 -251 101 -169
rect 114 -170 115 -164
rect 124 -251 125 -169
rect 1052 -251 1053 -169
rect 107 -251 108 -171
rect 870 -251 871 -171
rect 877 -172 878 -164
rect 1031 -251 1032 -171
rect 110 -251 111 -173
rect 418 -174 419 -164
rect 457 -174 458 -164
rect 590 -251 591 -173
rect 621 -174 622 -164
rect 1129 -251 1130 -173
rect 114 -251 115 -175
rect 492 -176 493 -164
rect 509 -176 510 -164
rect 1080 -251 1081 -175
rect 149 -178 150 -164
rect 247 -178 248 -164
rect 254 -251 255 -177
rect 429 -178 430 -164
rect 467 -178 468 -164
rect 674 -178 675 -164
rect 695 -178 696 -164
rect 712 -178 713 -164
rect 730 -251 731 -177
rect 982 -178 983 -164
rect 1003 -178 1004 -164
rect 1059 -251 1060 -177
rect 156 -180 157 -164
rect 492 -251 493 -179
rect 506 -180 507 -164
rect 674 -251 675 -179
rect 695 -251 696 -179
rect 989 -180 990 -164
rect 996 -180 997 -164
rect 1003 -251 1004 -179
rect 170 -182 171 -164
rect 289 -182 290 -164
rect 310 -182 311 -164
rect 341 -251 342 -181
rect 352 -251 353 -181
rect 488 -182 489 -164
rect 506 -251 507 -181
rect 520 -182 521 -164
rect 625 -182 626 -164
rect 625 -251 626 -181
rect 625 -182 626 -164
rect 625 -251 626 -181
rect 632 -182 633 -164
rect 716 -251 717 -181
rect 786 -182 787 -164
rect 863 -251 864 -181
rect 884 -182 885 -164
rect 1073 -251 1074 -181
rect 166 -251 167 -183
rect 520 -251 521 -183
rect 562 -184 563 -164
rect 632 -251 633 -183
rect 667 -184 668 -164
rect 670 -200 671 -183
rect 828 -184 829 -164
rect 1045 -251 1046 -183
rect 173 -251 174 -185
rect 292 -186 293 -164
rect 310 -251 311 -185
rect 474 -186 475 -164
rect 488 -251 489 -185
rect 698 -186 699 -164
rect 835 -186 836 -164
rect 884 -251 885 -185
rect 891 -186 892 -164
rect 1017 -251 1018 -185
rect 184 -188 185 -164
rect 450 -251 451 -187
rect 471 -251 472 -187
rect 541 -251 542 -187
rect 562 -251 563 -187
rect 702 -188 703 -164
rect 814 -188 815 -164
rect 891 -251 892 -187
rect 898 -188 899 -164
rect 1066 -251 1067 -187
rect 163 -190 164 -164
rect 184 -251 185 -189
rect 198 -190 199 -164
rect 198 -251 199 -189
rect 198 -190 199 -164
rect 198 -251 199 -189
rect 208 -251 209 -189
rect 212 -190 213 -164
rect 219 -190 220 -164
rect 247 -251 248 -189
rect 261 -190 262 -164
rect 436 -251 437 -189
rect 639 -190 640 -164
rect 702 -251 703 -189
rect 814 -251 815 -189
rect 828 -251 829 -189
rect 856 -190 857 -164
rect 982 -251 983 -189
rect 163 -251 164 -191
rect 835 -251 836 -191
rect 905 -192 906 -164
rect 989 -251 990 -191
rect 177 -194 178 -164
rect 639 -251 640 -193
rect 667 -251 668 -193
rect 744 -194 745 -164
rect 758 -194 759 -164
rect 856 -251 857 -193
rect 912 -194 913 -164
rect 1108 -251 1109 -193
rect 177 -251 178 -195
rect 303 -196 304 -164
rect 324 -196 325 -164
rect 457 -251 458 -195
rect 653 -196 654 -164
rect 758 -251 759 -195
rect 779 -196 780 -164
rect 912 -251 913 -195
rect 919 -196 920 -164
rect 1024 -251 1025 -195
rect 121 -251 122 -197
rect 324 -251 325 -197
rect 380 -198 381 -164
rect 527 -251 528 -197
rect 597 -198 598 -164
rect 653 -251 654 -197
rect 744 -251 745 -197
rect 793 -198 794 -164
rect 905 -251 906 -197
rect 926 -198 927 -164
rect 1010 -251 1011 -197
rect 212 -251 213 -199
rect 366 -200 367 -164
rect 380 -251 381 -199
rect 422 -200 423 -164
rect 432 -251 433 -199
rect 597 -251 598 -199
rect 712 -251 713 -199
rect 793 -251 794 -199
rect 821 -200 822 -164
rect 898 -251 899 -199
rect 933 -200 934 -164
rect 1094 -251 1095 -199
rect 219 -251 220 -201
rect 268 -251 269 -201
rect 282 -202 283 -164
rect 373 -202 374 -164
rect 394 -202 395 -164
rect 464 -202 465 -164
rect 737 -202 738 -164
rect 779 -251 780 -201
rect 842 -202 843 -164
rect 926 -251 927 -201
rect 943 -202 944 -164
rect 954 -251 955 -201
rect 961 -202 962 -164
rect 1038 -251 1039 -201
rect 222 -251 223 -203
rect 303 -251 304 -203
rect 331 -204 332 -164
rect 422 -251 423 -203
rect 464 -251 465 -203
rect 478 -204 479 -164
rect 611 -204 612 -164
rect 737 -251 738 -203
rect 754 -204 755 -164
rect 933 -251 934 -203
rect 947 -204 948 -164
rect 996 -251 997 -203
rect 226 -206 227 -164
rect 275 -206 276 -164
rect 285 -251 286 -205
rect 558 -206 559 -164
rect 681 -206 682 -164
rect 961 -251 962 -205
rect 968 -206 969 -164
rect 1115 -251 1116 -205
rect 226 -251 227 -207
rect 548 -208 549 -164
rect 681 -251 682 -207
rect 947 -251 948 -207
rect 975 -208 976 -164
rect 999 -208 1000 -164
rect 240 -210 241 -164
rect 275 -251 276 -209
rect 289 -251 290 -209
rect 611 -251 612 -209
rect 705 -210 706 -164
rect 968 -251 969 -209
rect 250 -212 251 -164
rect 282 -251 283 -211
rect 317 -212 318 -164
rect 975 -251 976 -211
rect 261 -251 262 -213
rect 429 -251 430 -213
rect 478 -251 479 -213
rect 877 -251 878 -213
rect 271 -216 272 -164
rect 331 -251 332 -215
rect 359 -216 360 -164
rect 373 -251 374 -215
rect 394 -251 395 -215
rect 408 -216 409 -164
rect 415 -251 416 -215
rect 513 -216 514 -164
rect 548 -251 549 -215
rect 583 -216 584 -164
rect 772 -216 773 -164
rect 821 -251 822 -215
rect 849 -216 850 -164
rect 919 -251 920 -215
rect 205 -218 206 -164
rect 359 -251 360 -217
rect 366 -251 367 -217
rect 684 -251 685 -217
rect 723 -218 724 -164
rect 772 -251 773 -217
rect 205 -251 206 -219
rect 485 -220 486 -164
rect 513 -251 514 -219
rect 660 -220 661 -164
rect 765 -220 766 -164
rect 849 -251 850 -219
rect 257 -222 258 -164
rect 408 -251 409 -221
rect 604 -222 605 -164
rect 660 -251 661 -221
rect 765 -251 766 -221
rect 786 -251 787 -221
rect 345 -224 346 -164
rect 583 -251 584 -223
rect 646 -224 647 -164
rect 723 -251 724 -223
rect 278 -226 279 -164
rect 345 -251 346 -225
rect 401 -226 402 -164
rect 404 -251 405 -225
rect 569 -226 570 -164
rect 604 -251 605 -225
rect 401 -251 402 -227
rect 751 -251 752 -227
rect 534 -230 535 -164
rect 569 -251 570 -229
rect 576 -230 577 -164
rect 646 -251 647 -229
rect 233 -232 234 -164
rect 576 -251 577 -231
rect 191 -234 192 -164
rect 233 -251 234 -233
rect 534 -251 535 -233
rect 807 -234 808 -164
rect 191 -251 192 -235
rect 446 -251 447 -235
rect 800 -236 801 -164
rect 807 -251 808 -235
rect 709 -238 710 -164
rect 800 -251 801 -237
rect 387 -240 388 -164
rect 709 -251 710 -239
rect 387 -251 388 -241
rect 499 -242 500 -164
rect 443 -244 444 -164
rect 499 -251 500 -243
rect 296 -246 297 -164
rect 443 -251 444 -245
rect 296 -251 297 -247
rect 338 -248 339 -164
rect 338 -251 339 -249
rect 1101 -251 1102 -249
rect 54 -261 55 -259
rect 282 -261 283 -259
rect 296 -261 297 -259
rect 443 -354 444 -260
rect 481 -261 482 -259
rect 576 -261 577 -259
rect 614 -261 615 -259
rect 1031 -261 1032 -259
rect 1038 -261 1039 -259
rect 1206 -354 1207 -260
rect 72 -263 73 -259
rect 121 -354 122 -262
rect 124 -263 125 -259
rect 208 -263 209 -259
rect 219 -263 220 -259
rect 912 -263 913 -259
rect 947 -263 948 -259
rect 1031 -354 1032 -262
rect 1052 -263 1053 -259
rect 1262 -354 1263 -262
rect 79 -354 80 -264
rect 1185 -354 1186 -264
rect 86 -354 87 -266
rect 100 -267 101 -259
rect 110 -267 111 -259
rect 338 -267 339 -259
rect 345 -267 346 -259
rect 429 -354 430 -266
rect 481 -354 482 -266
rect 856 -267 857 -259
rect 898 -267 899 -259
rect 947 -354 948 -266
rect 954 -267 955 -259
rect 1136 -354 1137 -266
rect 93 -354 94 -268
rect 579 -354 580 -268
rect 635 -354 636 -268
rect 1178 -354 1179 -268
rect 100 -354 101 -270
rect 373 -271 374 -259
rect 401 -271 402 -259
rect 471 -271 472 -259
rect 485 -271 486 -259
rect 506 -271 507 -259
rect 516 -271 517 -259
rect 716 -271 717 -259
rect 726 -354 727 -270
rect 1143 -354 1144 -270
rect 124 -354 125 -272
rect 1052 -354 1053 -272
rect 1059 -273 1060 -259
rect 1227 -354 1228 -272
rect 128 -275 129 -259
rect 131 -301 132 -274
rect 142 -354 143 -274
rect 191 -275 192 -259
rect 219 -354 220 -274
rect 604 -275 605 -259
rect 663 -354 664 -274
rect 1066 -275 1067 -259
rect 1073 -275 1074 -259
rect 1241 -354 1242 -274
rect 128 -354 129 -276
rect 205 -277 206 -259
rect 240 -354 241 -276
rect 261 -277 262 -259
rect 289 -277 290 -259
rect 345 -354 346 -276
rect 359 -277 360 -259
rect 401 -354 402 -276
rect 457 -277 458 -259
rect 506 -354 507 -276
rect 530 -354 531 -276
rect 842 -277 843 -259
rect 849 -277 850 -259
rect 898 -354 899 -276
rect 954 -354 955 -276
rect 1129 -277 1130 -259
rect 149 -354 150 -278
rect 233 -279 234 -259
rect 254 -279 255 -259
rect 583 -279 584 -259
rect 604 -354 605 -278
rect 1045 -279 1046 -259
rect 1080 -279 1081 -259
rect 1269 -354 1270 -278
rect 156 -354 157 -280
rect 338 -354 339 -280
rect 488 -281 489 -259
rect 1038 -354 1039 -280
rect 1087 -281 1088 -259
rect 1290 -354 1291 -280
rect 163 -283 164 -259
rect 436 -283 437 -259
rect 467 -354 468 -282
rect 1087 -354 1088 -282
rect 1094 -283 1095 -259
rect 1283 -354 1284 -282
rect 82 -354 83 -284
rect 436 -354 437 -284
rect 492 -285 493 -259
rect 737 -285 738 -259
rect 744 -285 745 -259
rect 856 -354 857 -284
rect 877 -285 878 -259
rect 1066 -354 1067 -284
rect 163 -354 164 -286
rect 415 -287 416 -259
rect 541 -287 542 -259
rect 730 -287 731 -259
rect 765 -287 766 -259
rect 1276 -354 1277 -286
rect 184 -289 185 -259
rect 191 -354 192 -288
rect 198 -289 199 -259
rect 205 -354 206 -288
rect 212 -289 213 -259
rect 457 -354 458 -288
rect 513 -289 514 -259
rect 541 -354 542 -288
rect 544 -289 545 -259
rect 1150 -354 1151 -288
rect 58 -354 59 -290
rect 212 -354 213 -290
rect 254 -354 255 -290
rect 387 -291 388 -259
rect 408 -291 409 -259
rect 730 -354 731 -290
rect 768 -291 769 -259
rect 905 -291 906 -259
rect 933 -291 934 -259
rect 1080 -354 1081 -290
rect 107 -293 108 -259
rect 184 -354 185 -292
rect 268 -293 269 -259
rect 289 -354 290 -292
rect 296 -354 297 -292
rect 317 -293 318 -259
rect 320 -293 321 -259
rect 639 -293 640 -259
rect 646 -293 647 -259
rect 765 -354 766 -292
rect 779 -293 780 -259
rect 877 -354 878 -292
rect 884 -293 885 -259
rect 1094 -354 1095 -292
rect 107 -354 108 -294
rect 275 -295 276 -259
rect 303 -295 304 -259
rect 373 -354 374 -294
rect 387 -354 388 -294
rect 534 -295 535 -259
rect 548 -295 549 -259
rect 593 -354 594 -294
rect 597 -295 598 -259
rect 744 -354 745 -294
rect 751 -295 752 -259
rect 884 -354 885 -294
rect 891 -295 892 -259
rect 1045 -354 1046 -294
rect 114 -297 115 -259
rect 548 -354 549 -296
rect 562 -297 563 -259
rect 597 -354 598 -296
rect 625 -297 626 -259
rect 646 -354 647 -296
rect 702 -297 703 -259
rect 828 -354 829 -296
rect 831 -297 832 -259
rect 996 -297 997 -259
rect 1003 -297 1004 -259
rect 1171 -354 1172 -296
rect 135 -299 136 -259
rect 198 -354 199 -298
rect 247 -299 248 -259
rect 268 -354 269 -298
rect 275 -354 276 -298
rect 422 -299 423 -259
rect 471 -354 472 -298
rect 779 -354 780 -298
rect 786 -299 787 -259
rect 1059 -354 1060 -298
rect 135 -354 136 -300
rect 177 -301 178 -259
rect 408 -354 409 -300
rect 415 -354 416 -300
rect 562 -354 563 -300
rect 569 -301 570 -259
rect 625 -354 626 -300
rect 632 -301 633 -259
rect 737 -354 738 -300
rect 772 -301 773 -259
rect 891 -354 892 -300
rect 940 -301 941 -259
rect 996 -354 997 -300
rect 1010 -301 1011 -259
rect 1199 -354 1200 -300
rect 177 -354 178 -302
rect 495 -303 496 -259
rect 499 -303 500 -259
rect 534 -354 535 -302
rect 569 -354 570 -302
rect 800 -303 801 -259
rect 807 -303 808 -259
rect 1073 -354 1074 -302
rect 236 -354 237 -304
rect 940 -354 941 -304
rect 968 -305 969 -259
rect 1157 -354 1158 -304
rect 303 -354 304 -306
rect 478 -307 479 -259
rect 513 -354 514 -306
rect 1010 -354 1011 -306
rect 1017 -307 1018 -259
rect 1234 -354 1235 -306
rect 114 -354 115 -308
rect 478 -354 479 -308
rect 520 -309 521 -259
rect 751 -354 752 -308
rect 793 -309 794 -259
rect 912 -354 913 -308
rect 968 -354 969 -308
rect 1122 -309 1123 -259
rect 317 -354 318 -310
rect 352 -311 353 -259
rect 366 -311 367 -259
rect 422 -354 423 -310
rect 464 -311 465 -259
rect 499 -354 500 -310
rect 520 -354 521 -310
rect 527 -311 528 -259
rect 576 -354 577 -310
rect 793 -354 794 -310
rect 814 -311 815 -259
rect 905 -354 906 -310
rect 961 -311 962 -259
rect 1122 -354 1123 -310
rect 310 -313 311 -259
rect 352 -354 353 -312
rect 404 -313 405 -259
rect 961 -354 962 -312
rect 975 -313 976 -259
rect 1164 -354 1165 -312
rect 310 -354 311 -314
rect 324 -315 325 -259
rect 485 -354 486 -314
rect 814 -354 815 -314
rect 821 -315 822 -259
rect 849 -354 850 -314
rect 863 -315 864 -259
rect 933 -354 934 -314
rect 982 -315 983 -259
rect 1192 -354 1193 -314
rect 324 -354 325 -316
rect 331 -317 332 -259
rect 527 -354 528 -316
rect 1220 -354 1221 -316
rect 583 -354 584 -318
rect 1101 -319 1102 -259
rect 632 -354 633 -320
rect 1108 -321 1109 -259
rect 586 -323 587 -259
rect 1108 -354 1109 -322
rect 586 -354 587 -324
rect 975 -354 976 -324
rect 989 -325 990 -259
rect 1255 -354 1256 -324
rect 639 -354 640 -326
rect 667 -327 668 -259
rect 674 -327 675 -259
rect 821 -354 822 -326
rect 835 -327 836 -259
rect 1129 -354 1130 -326
rect 607 -354 608 -328
rect 835 -354 836 -328
rect 842 -354 843 -328
rect 1115 -329 1116 -259
rect 611 -331 612 -259
rect 674 -354 675 -330
rect 684 -354 685 -330
rect 807 -354 808 -330
rect 870 -331 871 -259
rect 1003 -354 1004 -330
rect 1024 -331 1025 -259
rect 1248 -354 1249 -330
rect 72 -354 73 -332
rect 611 -354 612 -332
rect 618 -333 619 -259
rect 667 -354 668 -332
rect 688 -333 689 -259
rect 870 -354 871 -332
rect 919 -333 920 -259
rect 1115 -354 1116 -332
rect 450 -335 451 -259
rect 618 -354 619 -334
rect 653 -335 654 -259
rect 688 -354 689 -334
rect 695 -335 696 -259
rect 863 -354 864 -334
rect 926 -335 927 -259
rect 1101 -354 1102 -334
rect 226 -337 227 -259
rect 695 -354 696 -336
rect 709 -337 710 -259
rect 1017 -354 1018 -336
rect 226 -354 227 -338
rect 341 -339 342 -259
rect 446 -339 447 -259
rect 450 -354 451 -338
rect 488 -354 489 -338
rect 919 -354 920 -338
rect 555 -341 556 -259
rect 653 -354 654 -340
rect 660 -341 661 -259
rect 702 -354 703 -340
rect 719 -354 720 -340
rect 982 -354 983 -340
rect 394 -343 395 -259
rect 555 -354 556 -342
rect 590 -343 591 -259
rect 709 -354 710 -342
rect 723 -343 724 -259
rect 800 -354 801 -342
rect 845 -343 846 -259
rect 1024 -354 1025 -342
rect 173 -345 174 -259
rect 394 -354 395 -344
rect 590 -354 591 -344
rect 1213 -354 1214 -344
rect 758 -347 759 -259
rect 989 -354 990 -346
rect 380 -349 381 -259
rect 758 -354 759 -348
rect 786 -354 787 -348
rect 926 -354 927 -348
rect 170 -351 171 -259
rect 380 -354 381 -350
rect 51 -354 52 -352
rect 170 -354 171 -352
rect 58 -364 59 -362
rect 1059 -364 1060 -362
rect 1227 -364 1228 -362
rect 1311 -479 1312 -363
rect 1332 -479 1333 -363
rect 1374 -479 1375 -363
rect 65 -479 66 -365
rect 338 -366 339 -362
rect 366 -479 367 -365
rect 541 -366 542 -362
rect 548 -366 549 -362
rect 548 -479 549 -365
rect 548 -366 549 -362
rect 548 -479 549 -365
rect 558 -479 559 -365
rect 891 -366 892 -362
rect 919 -366 920 -362
rect 1318 -479 1319 -365
rect 79 -479 80 -367
rect 82 -368 83 -362
rect 96 -479 97 -367
rect 975 -368 976 -362
rect 1038 -368 1039 -362
rect 1297 -479 1298 -367
rect 1300 -368 1301 -362
rect 1304 -479 1305 -367
rect 114 -370 115 -362
rect 474 -370 475 -362
rect 485 -370 486 -362
rect 758 -370 759 -362
rect 786 -479 787 -369
rect 1171 -370 1172 -362
rect 1234 -370 1235 -362
rect 1325 -479 1326 -369
rect 124 -372 125 -362
rect 128 -372 129 -362
rect 149 -372 150 -362
rect 159 -372 160 -362
rect 163 -372 164 -362
rect 261 -479 262 -371
rect 296 -372 297 -362
rect 516 -372 517 -362
rect 530 -372 531 -362
rect 863 -372 864 -362
rect 891 -479 892 -371
rect 954 -372 955 -362
rect 996 -372 997 -362
rect 1171 -479 1172 -371
rect 1248 -372 1249 -362
rect 1339 -479 1340 -371
rect 128 -479 129 -373
rect 303 -374 304 -362
rect 310 -374 311 -362
rect 537 -479 538 -373
rect 565 -374 566 -362
rect 1143 -374 1144 -362
rect 1157 -374 1158 -362
rect 1248 -479 1249 -373
rect 1255 -374 1256 -362
rect 1346 -479 1347 -373
rect 152 -479 153 -375
rect 173 -376 174 -362
rect 184 -376 185 -362
rect 359 -479 360 -375
rect 380 -376 381 -362
rect 464 -479 465 -375
rect 488 -376 489 -362
rect 1087 -376 1088 -362
rect 1136 -376 1137 -362
rect 1234 -479 1235 -375
rect 1262 -376 1263 -362
rect 1353 -479 1354 -375
rect 163 -479 164 -377
rect 625 -378 626 -362
rect 677 -479 678 -377
rect 1073 -378 1074 -362
rect 1087 -479 1088 -377
rect 1213 -378 1214 -362
rect 1276 -378 1277 -362
rect 1360 -479 1361 -377
rect 170 -380 171 -362
rect 1241 -380 1242 -362
rect 1290 -380 1291 -362
rect 1367 -479 1368 -379
rect 170 -479 171 -381
rect 191 -382 192 -362
rect 198 -382 199 -362
rect 485 -479 486 -381
rect 513 -382 514 -362
rect 793 -382 794 -362
rect 800 -382 801 -362
rect 803 -408 804 -381
rect 831 -479 832 -381
rect 1003 -382 1004 -362
rect 1024 -382 1025 -362
rect 1073 -479 1074 -381
rect 1115 -382 1116 -362
rect 1213 -479 1214 -381
rect 184 -479 185 -383
rect 226 -384 227 -362
rect 240 -384 241 -362
rect 240 -479 241 -383
rect 240 -384 241 -362
rect 240 -479 241 -383
rect 247 -479 248 -383
rect 502 -479 503 -383
rect 516 -479 517 -383
rect 1227 -479 1228 -383
rect 191 -479 192 -385
rect 562 -386 563 -362
rect 579 -386 580 -362
rect 1283 -386 1284 -362
rect 198 -479 199 -387
rect 205 -388 206 -362
rect 219 -388 220 -362
rect 492 -479 493 -387
rect 534 -388 535 -362
rect 541 -479 542 -387
rect 562 -479 563 -387
rect 597 -388 598 -362
rect 604 -388 605 -362
rect 723 -388 724 -362
rect 726 -388 727 -362
rect 1122 -388 1123 -362
rect 1150 -388 1151 -362
rect 1241 -479 1242 -387
rect 124 -479 125 -389
rect 604 -479 605 -389
rect 607 -390 608 -362
rect 1059 -479 1060 -389
rect 1066 -390 1067 -362
rect 1136 -479 1137 -389
rect 1164 -390 1165 -362
rect 1262 -479 1263 -389
rect 135 -392 136 -362
rect 205 -479 206 -391
rect 219 -479 220 -391
rect 635 -392 636 -362
rect 684 -392 685 -362
rect 1080 -392 1081 -362
rect 1122 -479 1123 -391
rect 1178 -392 1179 -362
rect 1185 -392 1186 -362
rect 1276 -479 1277 -391
rect 135 -479 136 -393
rect 730 -394 731 -362
rect 754 -479 755 -393
rect 1220 -394 1221 -362
rect 226 -479 227 -395
rect 408 -396 409 -362
rect 457 -396 458 -362
rect 614 -479 615 -395
rect 632 -396 633 -362
rect 793 -479 794 -395
rect 800 -479 801 -395
rect 842 -396 843 -362
rect 849 -396 850 -362
rect 1066 -479 1067 -395
rect 1094 -396 1095 -362
rect 1185 -479 1186 -395
rect 1192 -396 1193 -362
rect 1283 -479 1284 -395
rect 296 -479 297 -397
rect 513 -479 514 -397
rect 576 -398 577 -362
rect 1164 -479 1165 -397
rect 1206 -398 1207 -362
rect 1290 -479 1291 -397
rect 303 -479 304 -399
rect 345 -400 346 -362
rect 373 -400 374 -362
rect 408 -479 409 -399
rect 481 -400 482 -362
rect 1080 -479 1081 -399
rect 1101 -400 1102 -362
rect 1192 -479 1193 -399
rect 310 -479 311 -401
rect 663 -402 664 -362
rect 716 -402 717 -362
rect 863 -479 864 -401
rect 898 -402 899 -362
rect 1255 -479 1256 -401
rect 324 -404 325 -362
rect 478 -404 479 -362
rect 576 -479 577 -403
rect 814 -404 815 -362
rect 828 -404 829 -362
rect 898 -479 899 -403
rect 905 -404 906 -362
rect 1150 -479 1151 -403
rect 107 -406 108 -362
rect 478 -479 479 -405
rect 579 -479 580 -405
rect 1206 -479 1207 -405
rect 107 -479 108 -407
rect 233 -408 234 -362
rect 289 -408 290 -362
rect 324 -479 325 -407
rect 331 -479 332 -407
rect 527 -408 528 -362
rect 583 -408 584 -362
rect 775 -408 776 -362
rect 842 -479 843 -407
rect 849 -479 850 -407
rect 989 -408 990 -362
rect 1031 -408 1032 -362
rect 1038 -479 1039 -407
rect 1052 -408 1053 -362
rect 1094 -479 1095 -407
rect 1101 -479 1102 -407
rect 1199 -408 1200 -362
rect 177 -410 178 -362
rect 527 -479 528 -409
rect 583 -479 584 -409
rect 716 -479 717 -409
rect 719 -479 720 -409
rect 954 -479 955 -409
rect 968 -410 969 -362
rect 1003 -479 1004 -409
rect 1010 -410 1011 -362
rect 1052 -479 1053 -409
rect 1108 -410 1109 -362
rect 1199 -479 1200 -409
rect 156 -412 157 -362
rect 1108 -479 1109 -411
rect 131 -479 132 -413
rect 156 -479 157 -413
rect 177 -479 178 -413
rect 467 -414 468 -362
rect 586 -414 587 -362
rect 884 -414 885 -362
rect 912 -414 913 -362
rect 1143 -479 1144 -413
rect 233 -479 234 -415
rect 709 -416 710 -362
rect 723 -479 724 -415
rect 884 -479 885 -415
rect 926 -416 927 -362
rect 989 -479 990 -415
rect 338 -479 339 -417
rect 457 -479 458 -417
rect 520 -418 521 -362
rect 912 -479 913 -417
rect 940 -418 941 -362
rect 996 -479 997 -417
rect 345 -479 346 -419
rect 443 -420 444 -362
rect 506 -420 507 -362
rect 520 -479 521 -419
rect 597 -479 598 -419
rect 1045 -420 1046 -362
rect 149 -479 150 -421
rect 1045 -479 1046 -421
rect 373 -479 374 -423
rect 681 -424 682 -362
rect 702 -424 703 -362
rect 814 -479 815 -423
rect 835 -424 836 -362
rect 905 -479 906 -423
rect 982 -424 983 -362
rect 1024 -479 1025 -423
rect 380 -479 381 -425
rect 436 -426 437 -362
rect 611 -426 612 -362
rect 625 -479 626 -425
rect 632 -479 633 -425
rect 1017 -426 1018 -362
rect 387 -428 388 -362
rect 506 -479 507 -427
rect 635 -479 636 -427
rect 1269 -428 1270 -362
rect 352 -430 353 -362
rect 387 -479 388 -429
rect 394 -430 395 -362
rect 572 -430 573 -362
rect 642 -479 643 -429
rect 1010 -479 1011 -429
rect 72 -432 73 -362
rect 394 -479 395 -431
rect 401 -432 402 -362
rect 975 -479 976 -431
rect 72 -479 73 -433
rect 86 -434 87 -362
rect 100 -434 101 -362
rect 352 -479 353 -433
rect 401 -479 402 -433
rect 499 -434 500 -362
rect 660 -434 661 -362
rect 1178 -479 1179 -433
rect 86 -479 87 -435
rect 212 -436 213 -362
rect 422 -436 423 -362
rect 436 -479 437 -435
rect 499 -479 500 -435
rect 555 -436 556 -362
rect 660 -479 661 -435
rect 674 -436 675 -362
rect 684 -479 685 -435
rect 1269 -479 1270 -435
rect 100 -479 101 -437
rect 275 -438 276 -362
rect 415 -438 416 -362
rect 422 -479 423 -437
rect 429 -438 430 -362
rect 443 -479 444 -437
rect 555 -479 556 -437
rect 1115 -479 1116 -437
rect 212 -479 213 -439
rect 961 -440 962 -362
rect 254 -442 255 -362
rect 429 -479 430 -441
rect 667 -442 668 -362
rect 709 -479 710 -441
rect 730 -479 731 -441
rect 765 -442 766 -362
rect 772 -442 773 -362
rect 940 -479 941 -441
rect 947 -442 948 -362
rect 961 -479 962 -441
rect 254 -479 255 -443
rect 471 -444 472 -362
rect 534 -479 535 -443
rect 947 -479 948 -443
rect 317 -446 318 -362
rect 415 -479 416 -445
rect 667 -479 668 -445
rect 821 -446 822 -362
rect 870 -446 871 -362
rect 926 -479 927 -445
rect 933 -446 934 -362
rect 982 -479 983 -445
rect 268 -448 269 -362
rect 317 -479 318 -447
rect 355 -479 356 -447
rect 471 -479 472 -447
rect 590 -448 591 -362
rect 870 -479 871 -447
rect 877 -448 878 -362
rect 933 -479 934 -447
rect 93 -450 94 -362
rect 268 -479 269 -449
rect 590 -479 591 -449
rect 653 -450 654 -362
rect 688 -450 689 -362
rect 877 -479 878 -449
rect 887 -479 888 -449
rect 1017 -479 1018 -449
rect 51 -452 52 -362
rect 688 -479 689 -451
rect 702 -479 703 -451
rect 737 -452 738 -362
rect 744 -452 745 -362
rect 765 -479 766 -451
rect 789 -452 790 -362
rect 835 -479 836 -451
rect 569 -454 570 -362
rect 653 -479 654 -453
rect 674 -479 675 -453
rect 737 -479 738 -453
rect 751 -454 752 -362
rect 1031 -479 1032 -453
rect 142 -456 143 -362
rect 569 -479 570 -455
rect 695 -456 696 -362
rect 744 -479 745 -455
rect 758 -479 759 -455
rect 968 -479 969 -455
rect 142 -479 143 -457
rect 215 -479 216 -457
rect 695 -479 696 -457
rect 1157 -479 1158 -457
rect 789 -479 790 -459
rect 919 -479 920 -459
rect 807 -462 808 -362
rect 1220 -479 1221 -461
rect 779 -464 780 -362
rect 807 -479 808 -463
rect 821 -479 822 -463
rect 856 -464 857 -362
rect 639 -466 640 -362
rect 779 -479 780 -465
rect 639 -479 640 -467
rect 1129 -468 1130 -362
rect 611 -479 612 -469
rect 1129 -479 1130 -469
rect 646 -472 647 -362
rect 856 -479 857 -471
rect 618 -474 619 -362
rect 646 -479 647 -473
rect 450 -476 451 -362
rect 618 -479 619 -475
rect 450 -479 451 -477
rect 460 -479 461 -477
rect 58 -612 59 -488
rect 590 -489 591 -487
rect 611 -489 612 -487
rect 1297 -489 1298 -487
rect 1346 -489 1347 -487
rect 1346 -612 1347 -488
rect 1346 -489 1347 -487
rect 1346 -612 1347 -488
rect 1377 -489 1378 -487
rect 1381 -612 1382 -488
rect 65 -491 66 -487
rect 275 -612 276 -490
rect 310 -491 311 -487
rect 355 -491 356 -487
rect 373 -491 374 -487
rect 600 -491 601 -487
rect 625 -491 626 -487
rect 695 -491 696 -487
rect 698 -612 699 -490
rect 1318 -491 1319 -487
rect 51 -612 52 -492
rect 65 -612 66 -492
rect 68 -612 69 -492
rect 205 -493 206 -487
rect 212 -612 213 -492
rect 219 -493 220 -487
rect 233 -493 234 -487
rect 761 -493 762 -487
rect 768 -612 769 -492
rect 1325 -493 1326 -487
rect 72 -495 73 -487
rect 96 -495 97 -487
rect 114 -612 115 -494
rect 128 -495 129 -487
rect 131 -495 132 -487
rect 282 -612 283 -494
rect 338 -495 339 -487
rect 789 -495 790 -487
rect 831 -495 832 -487
rect 1283 -495 1284 -487
rect 1325 -612 1326 -494
rect 1353 -495 1354 -487
rect 72 -612 73 -496
rect 79 -497 80 -487
rect 124 -497 125 -487
rect 506 -497 507 -487
rect 513 -497 514 -487
rect 975 -497 976 -487
rect 978 -612 979 -496
rect 1283 -612 1284 -496
rect 128 -612 129 -498
rect 247 -499 248 -487
rect 254 -499 255 -487
rect 544 -612 545 -498
rect 569 -499 570 -487
rect 810 -612 811 -498
rect 849 -499 850 -487
rect 849 -612 850 -498
rect 849 -499 850 -487
rect 849 -612 850 -498
rect 863 -499 864 -487
rect 863 -612 864 -498
rect 863 -499 864 -487
rect 863 -612 864 -498
rect 884 -499 885 -487
rect 1367 -499 1368 -487
rect 152 -501 153 -487
rect 170 -501 171 -487
rect 177 -501 178 -487
rect 338 -612 339 -500
rect 373 -612 374 -500
rect 775 -612 776 -500
rect 782 -612 783 -500
rect 1143 -501 1144 -487
rect 1206 -501 1207 -487
rect 1206 -612 1207 -500
rect 1206 -501 1207 -487
rect 1206 -612 1207 -500
rect 152 -612 153 -502
rect 184 -503 185 -487
rect 198 -503 199 -487
rect 205 -612 206 -502
rect 215 -503 216 -487
rect 912 -503 913 -487
rect 933 -503 934 -487
rect 933 -612 934 -502
rect 933 -503 934 -487
rect 933 -612 934 -502
rect 954 -503 955 -487
rect 1143 -612 1144 -502
rect 156 -505 157 -487
rect 579 -505 580 -487
rect 586 -612 587 -504
rect 877 -505 878 -487
rect 887 -505 888 -487
rect 1388 -612 1389 -504
rect 163 -507 164 -487
rect 625 -612 626 -506
rect 646 -507 647 -487
rect 670 -612 671 -506
rect 688 -507 689 -487
rect 884 -612 885 -506
rect 891 -507 892 -487
rect 1374 -612 1375 -506
rect 163 -612 164 -508
rect 408 -509 409 -487
rect 460 -509 461 -487
rect 856 -509 857 -487
rect 870 -509 871 -487
rect 1367 -612 1368 -508
rect 156 -612 157 -510
rect 870 -612 871 -510
rect 912 -612 913 -510
rect 926 -511 927 -487
rect 968 -511 969 -487
rect 1318 -612 1319 -510
rect 177 -612 178 -512
rect 639 -513 640 -487
rect 688 -612 689 -512
rect 779 -513 780 -487
rect 786 -513 787 -487
rect 1213 -513 1214 -487
rect 184 -612 185 -514
rect 653 -515 654 -487
rect 705 -612 706 -514
rect 1031 -515 1032 -487
rect 1045 -515 1046 -487
rect 1472 -612 1473 -514
rect 219 -612 220 -516
rect 478 -517 479 -487
rect 499 -517 500 -487
rect 989 -517 990 -487
rect 1045 -612 1046 -516
rect 1353 -612 1354 -516
rect 222 -612 223 -518
rect 968 -612 969 -518
rect 982 -519 983 -487
rect 982 -612 983 -518
rect 982 -519 983 -487
rect 982 -612 983 -518
rect 989 -612 990 -518
rect 1003 -519 1004 -487
rect 1087 -519 1088 -487
rect 1297 -612 1298 -518
rect 240 -521 241 -487
rect 289 -612 290 -520
rect 296 -521 297 -487
rect 646 -612 647 -520
rect 653 -612 654 -520
rect 737 -521 738 -487
rect 754 -521 755 -487
rect 1059 -521 1060 -487
rect 1178 -521 1179 -487
rect 1213 -612 1214 -520
rect 243 -612 244 -522
rect 611 -612 612 -522
rect 614 -523 615 -487
rect 1059 -612 1060 -522
rect 1178 -612 1179 -522
rect 1234 -523 1235 -487
rect 268 -525 269 -487
rect 310 -612 311 -524
rect 380 -525 381 -487
rect 506 -612 507 -524
rect 513 -612 514 -524
rect 667 -525 668 -487
rect 709 -525 710 -487
rect 709 -612 710 -524
rect 709 -525 710 -487
rect 709 -612 710 -524
rect 716 -525 717 -487
rect 1255 -525 1256 -487
rect 268 -612 269 -526
rect 331 -527 332 -487
rect 359 -527 360 -487
rect 716 -612 717 -526
rect 719 -527 720 -487
rect 1150 -527 1151 -487
rect 1248 -527 1249 -487
rect 1255 -612 1256 -526
rect 107 -529 108 -487
rect 359 -612 360 -528
rect 397 -612 398 -528
rect 681 -612 682 -528
rect 737 -612 738 -528
rect 744 -529 745 -487
rect 751 -529 752 -487
rect 1234 -612 1235 -528
rect 1241 -529 1242 -487
rect 1248 -612 1249 -528
rect 107 -612 108 -530
rect 828 -531 829 -487
rect 835 -531 836 -487
rect 877 -612 878 -530
rect 901 -612 902 -530
rect 1031 -612 1032 -530
rect 1150 -612 1151 -530
rect 1164 -531 1165 -487
rect 159 -612 160 -532
rect 1241 -612 1242 -532
rect 296 -612 297 -534
rect 401 -535 402 -487
rect 408 -612 409 -534
rect 415 -535 416 -487
rect 499 -612 500 -534
rect 891 -612 892 -534
rect 926 -612 927 -534
rect 1080 -535 1081 -487
rect 1164 -612 1165 -534
rect 1171 -535 1172 -487
rect 317 -537 318 -487
rect 380 -612 381 -536
rect 401 -612 402 -536
rect 632 -537 633 -487
rect 733 -612 734 -536
rect 751 -612 752 -536
rect 772 -537 773 -487
rect 1017 -537 1018 -487
rect 1073 -537 1074 -487
rect 1080 -612 1081 -536
rect 1171 -612 1172 -536
rect 1185 -537 1186 -487
rect 303 -539 304 -487
rect 317 -612 318 -538
rect 324 -539 325 -487
rect 331 -612 332 -538
rect 366 -539 367 -487
rect 744 -612 745 -538
rect 786 -612 787 -538
rect 800 -539 801 -487
rect 814 -539 815 -487
rect 828 -612 829 -538
rect 835 -612 836 -538
rect 842 -539 843 -487
rect 856 -612 857 -538
rect 1052 -539 1053 -487
rect 1073 -612 1074 -538
rect 1108 -539 1109 -487
rect 1185 -612 1186 -538
rect 1199 -539 1200 -487
rect 261 -541 262 -487
rect 303 -612 304 -540
rect 324 -612 325 -540
rect 387 -541 388 -487
rect 415 -612 416 -540
rect 443 -541 444 -487
rect 502 -541 503 -487
rect 793 -541 794 -487
rect 821 -541 822 -487
rect 842 -612 843 -540
rect 919 -541 920 -487
rect 1017 -612 1018 -540
rect 1108 -612 1109 -540
rect 1192 -541 1193 -487
rect 387 -612 388 -542
rect 457 -543 458 -487
rect 502 -612 503 -542
rect 1276 -543 1277 -487
rect 443 -612 444 -544
rect 618 -545 619 -487
rect 674 -545 675 -487
rect 1052 -612 1053 -544
rect 1101 -545 1102 -487
rect 1192 -612 1193 -544
rect 1276 -612 1277 -544
rect 1304 -545 1305 -487
rect 450 -547 451 -487
rect 457 -612 458 -546
rect 492 -547 493 -487
rect 618 -612 619 -546
rect 660 -547 661 -487
rect 674 -612 675 -546
rect 730 -547 731 -487
rect 800 -612 801 -546
rect 807 -547 808 -487
rect 821 -612 822 -546
rect 919 -612 920 -546
rect 996 -547 997 -487
rect 1003 -612 1004 -546
rect 1024 -547 1025 -487
rect 1094 -547 1095 -487
rect 1101 -612 1102 -546
rect 1115 -547 1116 -487
rect 1199 -612 1200 -546
rect 1304 -612 1305 -546
rect 1311 -547 1312 -487
rect 121 -549 122 -487
rect 1115 -612 1116 -548
rect 1311 -612 1312 -548
rect 1339 -549 1340 -487
rect 121 -612 122 -550
rect 530 -612 531 -550
rect 534 -551 535 -487
rect 562 -551 563 -487
rect 590 -612 591 -550
rect 597 -551 598 -487
rect 604 -551 605 -487
rect 954 -612 955 -550
rect 975 -612 976 -550
rect 1087 -612 1088 -550
rect 1094 -612 1095 -550
rect 1129 -551 1130 -487
rect 1332 -551 1333 -487
rect 1339 -612 1340 -550
rect 93 -553 94 -487
rect 1332 -612 1333 -552
rect 142 -555 143 -487
rect 597 -612 598 -554
rect 635 -555 636 -487
rect 1129 -612 1130 -554
rect 135 -557 136 -487
rect 142 -612 143 -556
rect 394 -557 395 -487
rect 534 -612 535 -556
rect 537 -557 538 -487
rect 898 -557 899 -487
rect 940 -557 941 -487
rect 996 -612 997 -556
rect 135 -612 136 -558
rect 1262 -559 1263 -487
rect 149 -561 150 -487
rect 940 -612 941 -560
rect 149 -612 150 -562
rect 695 -612 696 -562
rect 779 -612 780 -562
rect 1262 -612 1263 -562
rect 191 -565 192 -487
rect 394 -612 395 -564
rect 429 -565 430 -487
rect 604 -612 605 -564
rect 639 -612 640 -564
rect 730 -612 731 -564
rect 793 -612 794 -564
rect 1269 -565 1270 -487
rect 191 -612 192 -566
rect 485 -567 486 -487
rect 492 -612 493 -566
rect 583 -567 584 -487
rect 660 -612 661 -566
rect 684 -567 685 -487
rect 1269 -612 1270 -566
rect 1290 -567 1291 -487
rect 345 -569 346 -487
rect 429 -612 430 -568
rect 436 -569 437 -487
rect 450 -612 451 -568
rect 471 -569 472 -487
rect 562 -612 563 -568
rect 583 -612 584 -568
rect 632 -612 633 -568
rect 1290 -612 1291 -568
rect 1360 -569 1361 -487
rect 198 -612 199 -570
rect 1360 -612 1361 -570
rect 250 -612 251 -572
rect 345 -612 346 -572
rect 352 -612 353 -572
rect 684 -612 685 -572
rect 422 -575 423 -487
rect 436 -612 437 -574
rect 464 -575 465 -487
rect 471 -612 472 -574
rect 485 -612 486 -574
rect 702 -575 703 -487
rect 100 -577 101 -487
rect 464 -612 465 -576
rect 478 -612 479 -576
rect 702 -612 703 -576
rect 86 -579 87 -487
rect 100 -612 101 -578
rect 422 -612 423 -578
rect 520 -579 521 -487
rect 527 -579 528 -487
rect 576 -612 577 -578
rect 79 -612 80 -580
rect 86 -612 87 -580
rect 520 -612 521 -580
rect 723 -581 724 -487
rect 527 -612 528 -582
rect 814 -612 815 -582
rect 548 -585 549 -487
rect 569 -612 570 -584
rect 723 -612 724 -584
rect 905 -585 906 -487
rect 226 -587 227 -487
rect 548 -612 549 -586
rect 555 -587 556 -487
rect 898 -612 899 -586
rect 905 -612 906 -586
rect 947 -587 948 -487
rect 40 -589 41 -487
rect 226 -612 227 -588
rect 541 -589 542 -487
rect 555 -612 556 -588
rect 947 -612 948 -588
rect 1010 -589 1011 -487
rect 40 -612 41 -590
rect 261 -612 262 -590
rect 541 -612 542 -590
rect 1220 -591 1221 -487
rect 1010 -612 1011 -592
rect 1122 -593 1123 -487
rect 1220 -612 1221 -592
rect 1227 -593 1228 -487
rect 807 -612 808 -594
rect 1227 -612 1228 -594
rect 961 -597 962 -487
rect 1122 -612 1123 -596
rect 961 -612 962 -598
rect 1066 -599 1067 -487
rect 1066 -612 1067 -600
rect 1136 -601 1137 -487
rect 1136 -612 1137 -602
rect 1157 -603 1158 -487
rect 1038 -605 1039 -487
rect 1157 -612 1158 -604
rect 758 -607 759 -487
rect 1038 -612 1039 -606
rect 758 -612 759 -608
rect 765 -609 766 -487
rect 765 -612 766 -610
rect 1024 -612 1025 -610
rect 44 -735 45 -621
rect 292 -735 293 -621
rect 387 -622 388 -620
rect 583 -622 584 -620
rect 649 -735 650 -621
rect 1115 -622 1116 -620
rect 1185 -622 1186 -620
rect 1395 -735 1396 -621
rect 1472 -622 1473 -620
rect 1633 -735 1634 -621
rect 51 -624 52 -620
rect 516 -624 517 -620
rect 527 -624 528 -620
rect 912 -624 913 -620
rect 975 -735 976 -623
rect 1045 -624 1046 -620
rect 1059 -624 1060 -620
rect 1185 -735 1186 -623
rect 1234 -624 1235 -620
rect 1500 -735 1501 -623
rect 51 -735 52 -625
rect 310 -626 311 -620
rect 397 -626 398 -620
rect 670 -626 671 -620
rect 684 -626 685 -620
rect 1255 -626 1256 -620
rect 1311 -626 1312 -620
rect 1409 -735 1410 -625
rect 72 -628 73 -620
rect 82 -628 83 -620
rect 107 -628 108 -620
rect 558 -735 559 -627
rect 698 -628 699 -620
rect 842 -628 843 -620
rect 887 -735 888 -627
rect 1101 -628 1102 -620
rect 1136 -628 1137 -620
rect 1234 -735 1235 -627
rect 1353 -628 1354 -620
rect 1381 -628 1382 -620
rect 1388 -628 1389 -620
rect 1570 -735 1571 -627
rect 65 -630 66 -620
rect 1101 -735 1102 -629
rect 1157 -630 1158 -620
rect 1311 -735 1312 -629
rect 1332 -630 1333 -620
rect 1381 -735 1382 -629
rect 65 -735 66 -631
rect 226 -632 227 -620
rect 233 -735 234 -631
rect 488 -735 489 -631
rect 537 -735 538 -631
rect 723 -632 724 -620
rect 730 -735 731 -631
rect 1213 -632 1214 -620
rect 1227 -632 1228 -620
rect 1255 -735 1256 -631
rect 1276 -632 1277 -620
rect 1353 -735 1354 -631
rect 1356 -632 1357 -620
rect 1367 -632 1368 -620
rect 72 -735 73 -633
rect 373 -634 374 -620
rect 429 -634 430 -620
rect 502 -634 503 -620
rect 541 -634 542 -620
rect 625 -634 626 -620
rect 702 -634 703 -620
rect 1374 -634 1375 -620
rect 82 -735 83 -635
rect 100 -636 101 -620
rect 114 -735 115 -635
rect 117 -636 118 -620
rect 128 -636 129 -620
rect 226 -735 227 -635
rect 243 -636 244 -620
rect 387 -735 388 -635
rect 432 -735 433 -635
rect 751 -636 752 -620
rect 772 -636 773 -620
rect 1339 -636 1340 -620
rect 1360 -636 1361 -620
rect 1521 -735 1522 -635
rect 86 -638 87 -620
rect 100 -735 101 -637
rect 128 -735 129 -637
rect 555 -638 556 -620
rect 702 -735 703 -637
rect 758 -638 759 -620
rect 768 -638 769 -620
rect 1360 -735 1361 -637
rect 86 -735 87 -639
rect 674 -640 675 -620
rect 705 -640 706 -620
rect 842 -735 843 -639
rect 898 -640 899 -620
rect 1010 -640 1011 -620
rect 1017 -640 1018 -620
rect 1115 -735 1116 -639
rect 1129 -640 1130 -620
rect 1227 -735 1228 -639
rect 1269 -640 1270 -620
rect 1339 -735 1340 -639
rect 138 -642 139 -620
rect 219 -642 220 -620
rect 247 -642 248 -620
rect 856 -642 857 -620
rect 863 -642 864 -620
rect 898 -735 899 -641
rect 940 -642 941 -620
rect 1010 -735 1011 -641
rect 1080 -642 1081 -620
rect 1136 -735 1137 -641
rect 1157 -735 1158 -641
rect 1164 -642 1165 -620
rect 1171 -642 1172 -620
rect 1276 -735 1277 -641
rect 1290 -642 1291 -620
rect 1388 -735 1389 -641
rect 107 -735 108 -643
rect 247 -735 248 -643
rect 250 -644 251 -620
rect 527 -735 528 -643
rect 555 -735 556 -643
rect 765 -644 766 -620
rect 772 -735 773 -643
rect 908 -735 909 -643
rect 954 -644 955 -620
rect 1045 -735 1046 -643
rect 1052 -644 1053 -620
rect 1164 -735 1165 -643
rect 1192 -644 1193 -620
rect 1332 -735 1333 -643
rect 142 -646 143 -620
rect 156 -646 157 -620
rect 159 -646 160 -620
rect 1402 -735 1403 -645
rect 149 -648 150 -620
rect 240 -735 241 -647
rect 250 -735 251 -647
rect 478 -648 479 -620
rect 485 -648 486 -620
rect 593 -735 594 -647
rect 674 -735 675 -647
rect 821 -648 822 -620
rect 831 -735 832 -647
rect 1178 -648 1179 -620
rect 1206 -648 1207 -620
rect 1269 -735 1270 -647
rect 1290 -735 1291 -647
rect 1304 -648 1305 -620
rect 1325 -648 1326 -620
rect 1374 -735 1375 -647
rect 152 -650 153 -620
rect 1199 -650 1200 -620
rect 1241 -650 1242 -620
rect 1304 -735 1305 -649
rect 156 -735 157 -651
rect 796 -652 797 -620
rect 807 -652 808 -620
rect 1346 -652 1347 -620
rect 163 -654 164 -620
rect 429 -735 430 -653
rect 443 -654 444 -620
rect 583 -735 584 -653
rect 586 -654 587 -620
rect 1199 -735 1200 -653
rect 1248 -654 1249 -620
rect 1346 -735 1347 -653
rect 163 -735 164 -655
rect 656 -735 657 -655
rect 695 -656 696 -620
rect 1129 -735 1130 -655
rect 1248 -735 1249 -655
rect 1426 -735 1427 -655
rect 58 -658 59 -620
rect 695 -735 696 -657
rect 709 -658 710 -620
rect 758 -735 759 -657
rect 775 -658 776 -620
rect 978 -658 979 -620
rect 982 -658 983 -620
rect 1052 -735 1053 -657
rect 1122 -658 1123 -620
rect 1206 -735 1207 -657
rect 58 -735 59 -659
rect 93 -735 94 -659
rect 170 -735 171 -659
rect 380 -660 381 -620
rect 415 -660 416 -620
rect 443 -735 444 -659
rect 450 -660 451 -620
rect 450 -735 451 -659
rect 450 -660 451 -620
rect 450 -735 451 -659
rect 457 -660 458 -620
rect 457 -735 458 -659
rect 457 -660 458 -620
rect 457 -735 458 -659
rect 471 -660 472 -620
rect 478 -735 479 -659
rect 565 -735 566 -659
rect 1192 -735 1193 -659
rect 187 -735 188 -661
rect 205 -662 206 -620
rect 219 -735 220 -661
rect 324 -662 325 -620
rect 345 -662 346 -620
rect 625 -735 626 -661
rect 716 -662 717 -620
rect 1325 -735 1326 -661
rect 124 -735 125 -663
rect 345 -735 346 -663
rect 373 -735 374 -663
rect 464 -664 465 -620
rect 471 -735 472 -663
rect 590 -664 591 -620
rect 607 -735 608 -663
rect 1241 -735 1242 -663
rect 149 -735 150 -665
rect 590 -735 591 -665
rect 716 -735 717 -665
rect 828 -666 829 -620
rect 856 -735 857 -665
rect 1367 -735 1368 -665
rect 198 -668 199 -620
rect 198 -735 199 -667
rect 198 -668 199 -620
rect 198 -735 199 -667
rect 201 -668 202 -620
rect 212 -668 213 -620
rect 268 -668 269 -620
rect 366 -735 367 -667
rect 380 -735 381 -667
rect 492 -668 493 -620
rect 719 -668 720 -620
rect 1094 -668 1095 -620
rect 205 -735 206 -669
rect 632 -670 633 -620
rect 723 -735 724 -669
rect 1297 -670 1298 -620
rect 212 -735 213 -671
rect 352 -672 353 -620
rect 401 -672 402 -620
rect 415 -735 416 -671
rect 464 -735 465 -671
rect 712 -735 713 -671
rect 726 -735 727 -671
rect 1017 -735 1018 -671
rect 1024 -672 1025 -620
rect 1122 -735 1123 -671
rect 268 -735 269 -673
rect 530 -674 531 -620
rect 733 -674 734 -620
rect 954 -735 955 -673
rect 961 -674 962 -620
rect 1178 -735 1179 -673
rect 275 -676 276 -620
rect 751 -735 752 -675
rect 779 -676 780 -620
rect 996 -676 997 -620
rect 1003 -676 1004 -620
rect 1213 -735 1214 -675
rect 254 -735 255 -677
rect 275 -735 276 -677
rect 282 -678 283 -620
rect 439 -735 440 -677
rect 611 -678 612 -620
rect 996 -735 997 -677
rect 1006 -735 1007 -677
rect 1143 -678 1144 -620
rect 282 -735 283 -679
rect 579 -735 580 -679
rect 737 -680 738 -620
rect 765 -735 766 -679
rect 786 -680 787 -620
rect 863 -735 864 -679
rect 877 -680 878 -620
rect 961 -735 962 -679
rect 968 -680 969 -620
rect 1080 -735 1081 -679
rect 121 -682 122 -620
rect 737 -735 738 -681
rect 744 -682 745 -620
rect 779 -735 780 -681
rect 793 -682 794 -620
rect 1416 -735 1417 -681
rect 121 -735 122 -683
rect 1073 -684 1074 -620
rect 296 -686 297 -620
rect 541 -735 542 -685
rect 646 -686 647 -620
rect 786 -735 787 -685
rect 793 -735 794 -685
rect 1318 -686 1319 -620
rect 289 -688 290 -620
rect 296 -735 297 -687
rect 310 -735 311 -687
rect 891 -688 892 -620
rect 905 -688 906 -620
rect 1024 -735 1025 -687
rect 1031 -688 1032 -620
rect 1143 -735 1144 -687
rect 1262 -688 1263 -620
rect 1318 -735 1319 -687
rect 317 -690 318 -620
rect 324 -735 325 -689
rect 352 -735 353 -689
rect 604 -690 605 -620
rect 618 -690 619 -620
rect 646 -735 647 -689
rect 733 -735 734 -689
rect 1073 -735 1074 -689
rect 1108 -690 1109 -620
rect 1262 -735 1263 -689
rect 317 -735 318 -691
rect 422 -692 423 -620
rect 513 -692 514 -620
rect 744 -735 745 -691
rect 800 -692 801 -620
rect 877 -735 878 -691
rect 884 -692 885 -620
rect 968 -735 969 -691
rect 989 -692 990 -620
rect 1094 -735 1095 -691
rect 401 -735 402 -693
rect 604 -735 605 -693
rect 660 -694 661 -620
rect 800 -735 801 -693
rect 807 -735 808 -693
rect 912 -735 913 -693
rect 933 -694 934 -620
rect 982 -735 983 -693
rect 992 -735 993 -693
rect 1150 -694 1151 -620
rect 408 -696 409 -620
rect 492 -735 493 -695
rect 513 -735 514 -695
rect 534 -696 535 -620
rect 576 -696 577 -620
rect 618 -735 619 -695
rect 660 -735 661 -695
rect 688 -696 689 -620
rect 814 -696 815 -620
rect 891 -735 892 -695
rect 905 -735 906 -695
rect 1283 -696 1284 -620
rect 68 -698 69 -620
rect 688 -735 689 -697
rect 821 -735 822 -697
rect 835 -698 836 -620
rect 884 -735 885 -697
rect 926 -698 927 -620
rect 1031 -735 1032 -697
rect 1059 -735 1060 -697
rect 1062 -735 1063 -697
rect 1297 -735 1298 -697
rect 96 -735 97 -699
rect 814 -735 815 -699
rect 828 -735 829 -699
rect 940 -735 941 -699
rect 1038 -700 1039 -620
rect 1171 -735 1172 -699
rect 1220 -700 1221 -620
rect 1283 -735 1284 -699
rect 135 -702 136 -620
rect 1038 -735 1039 -701
rect 1066 -702 1067 -620
rect 1108 -735 1109 -701
rect 135 -735 136 -703
rect 261 -704 262 -620
rect 359 -704 360 -620
rect 408 -735 409 -703
rect 422 -735 423 -703
rect 436 -704 437 -620
rect 520 -704 521 -620
rect 611 -735 612 -703
rect 667 -704 668 -620
rect 933 -735 934 -703
rect 1087 -704 1088 -620
rect 1220 -735 1221 -703
rect 184 -706 185 -620
rect 261 -735 262 -705
rect 359 -735 360 -705
rect 653 -706 654 -620
rect 667 -735 668 -705
rect 859 -735 860 -705
rect 870 -706 871 -620
rect 926 -735 927 -705
rect 947 -706 948 -620
rect 1087 -735 1088 -705
rect 436 -735 437 -707
rect 1150 -735 1151 -707
rect 520 -735 521 -709
rect 597 -710 598 -620
rect 653 -735 654 -709
rect 681 -735 682 -709
rect 835 -735 836 -709
rect 901 -710 902 -620
rect 919 -710 920 -620
rect 1066 -735 1067 -709
rect 534 -735 535 -711
rect 569 -712 570 -620
rect 849 -712 850 -620
rect 947 -735 948 -711
rect 548 -714 549 -620
rect 569 -735 570 -713
rect 709 -735 710 -713
rect 849 -735 850 -713
rect 919 -735 920 -713
rect 1430 -735 1431 -713
rect 548 -735 549 -715
rect 639 -716 640 -620
rect 394 -718 395 -620
rect 639 -735 640 -717
rect 177 -720 178 -620
rect 394 -735 395 -719
rect 562 -720 563 -620
rect 597 -735 598 -719
rect 177 -735 178 -721
rect 506 -722 507 -620
rect 191 -724 192 -620
rect 506 -735 507 -723
rect 191 -735 192 -725
rect 338 -726 339 -620
rect 303 -728 304 -620
rect 562 -735 563 -727
rect 303 -735 304 -729
rect 576 -735 577 -729
rect 331 -732 332 -620
rect 338 -735 339 -731
rect 184 -735 185 -733
rect 331 -735 332 -733
rect 37 -874 38 -744
rect 58 -745 59 -743
rect 79 -745 80 -743
rect 919 -745 920 -743
rect 922 -745 923 -743
rect 1402 -745 1403 -743
rect 1416 -745 1417 -743
rect 1608 -874 1609 -744
rect 1633 -745 1634 -743
rect 1696 -874 1697 -744
rect 44 -747 45 -743
rect 1556 -874 1557 -746
rect 1570 -747 1571 -743
rect 1626 -874 1627 -746
rect 44 -874 45 -748
rect 450 -749 451 -743
rect 467 -874 468 -748
rect 1437 -874 1438 -748
rect 1500 -749 1501 -743
rect 1619 -874 1620 -748
rect 58 -874 59 -750
rect 149 -751 150 -743
rect 166 -874 167 -750
rect 1458 -874 1459 -750
rect 1521 -751 1522 -743
rect 1591 -874 1592 -750
rect 1605 -874 1606 -750
rect 1612 -874 1613 -750
rect 82 -753 83 -743
rect 604 -874 605 -752
rect 607 -753 608 -743
rect 877 -753 878 -743
rect 884 -753 885 -743
rect 1521 -874 1522 -752
rect 93 -755 94 -743
rect 800 -755 801 -743
rect 807 -755 808 -743
rect 807 -874 808 -754
rect 807 -755 808 -743
rect 807 -874 808 -754
rect 821 -755 822 -743
rect 884 -874 885 -754
rect 905 -755 906 -743
rect 1346 -755 1347 -743
rect 1353 -755 1354 -743
rect 1549 -874 1550 -754
rect 93 -874 94 -756
rect 527 -757 528 -743
rect 537 -757 538 -743
rect 723 -757 724 -743
rect 730 -757 731 -743
rect 779 -757 780 -743
rect 782 -874 783 -756
rect 1220 -757 1221 -743
rect 1241 -757 1242 -743
rect 1416 -874 1417 -756
rect 1430 -757 1431 -743
rect 1633 -874 1634 -756
rect 33 -874 34 -758
rect 527 -874 528 -758
rect 558 -759 559 -743
rect 1507 -874 1508 -758
rect 103 -874 104 -760
rect 366 -761 367 -743
rect 485 -874 486 -760
rect 562 -761 563 -743
rect 565 -761 566 -743
rect 1094 -761 1095 -743
rect 1122 -761 1123 -743
rect 1542 -874 1543 -760
rect 124 -763 125 -743
rect 1570 -874 1571 -762
rect 128 -765 129 -743
rect 131 -829 132 -764
rect 138 -874 139 -764
rect 1360 -765 1361 -743
rect 1367 -765 1368 -743
rect 1577 -874 1578 -764
rect 128 -874 129 -766
rect 618 -767 619 -743
rect 632 -874 633 -766
rect 639 -767 640 -743
rect 649 -767 650 -743
rect 1367 -874 1368 -766
rect 1374 -767 1375 -743
rect 1584 -874 1585 -766
rect 142 -874 143 -768
rect 726 -769 727 -743
rect 730 -874 731 -768
rect 758 -769 759 -743
rect 765 -769 766 -743
rect 821 -874 822 -768
rect 828 -769 829 -743
rect 961 -769 962 -743
rect 1003 -769 1004 -743
rect 1426 -769 1427 -743
rect 149 -874 150 -770
rect 625 -771 626 -743
rect 628 -874 629 -770
rect 1374 -874 1375 -770
rect 1388 -771 1389 -743
rect 1514 -874 1515 -770
rect 184 -773 185 -743
rect 1493 -874 1494 -772
rect 184 -874 185 -774
rect 198 -775 199 -743
rect 205 -775 206 -743
rect 450 -874 451 -774
rect 488 -775 489 -743
rect 555 -775 556 -743
rect 576 -775 577 -743
rect 716 -775 717 -743
rect 733 -775 734 -743
rect 1423 -775 1424 -743
rect 187 -777 188 -743
rect 1213 -777 1214 -743
rect 1227 -777 1228 -743
rect 1388 -874 1389 -776
rect 191 -779 192 -743
rect 236 -874 237 -778
rect 240 -779 241 -743
rect 366 -874 367 -778
rect 471 -779 472 -743
rect 555 -874 556 -778
rect 576 -874 577 -778
rect 863 -779 864 -743
rect 870 -779 871 -743
rect 1444 -874 1445 -778
rect 191 -874 192 -780
rect 429 -781 430 -743
rect 471 -874 472 -780
rect 478 -781 479 -743
rect 499 -874 500 -780
rect 597 -781 598 -743
rect 625 -874 626 -780
rect 702 -781 703 -743
rect 709 -781 710 -743
rect 1276 -781 1277 -743
rect 1283 -781 1284 -743
rect 1472 -874 1473 -780
rect 198 -874 199 -782
rect 562 -874 563 -782
rect 579 -783 580 -743
rect 996 -783 997 -743
rect 1038 -783 1039 -743
rect 1094 -874 1095 -782
rect 1136 -783 1137 -743
rect 1227 -874 1228 -782
rect 1269 -783 1270 -743
rect 1465 -874 1466 -782
rect 205 -874 206 -784
rect 240 -874 241 -784
rect 247 -874 248 -784
rect 1199 -785 1200 -743
rect 1206 -785 1207 -743
rect 1346 -874 1347 -784
rect 1381 -785 1382 -743
rect 1423 -874 1424 -784
rect 233 -787 234 -743
rect 996 -874 997 -786
rect 1080 -787 1081 -743
rect 1122 -874 1123 -786
rect 1157 -787 1158 -743
rect 1353 -874 1354 -786
rect 23 -874 24 -788
rect 233 -874 234 -788
rect 250 -789 251 -743
rect 1486 -874 1487 -788
rect 79 -874 80 -790
rect 250 -874 251 -790
rect 275 -791 276 -743
rect 380 -791 381 -743
rect 429 -874 430 -790
rect 492 -791 493 -743
rect 534 -791 535 -743
rect 1080 -874 1081 -790
rect 1171 -791 1172 -743
rect 1402 -874 1403 -790
rect 135 -793 136 -743
rect 534 -874 535 -792
rect 583 -793 584 -743
rect 597 -874 598 -792
rect 642 -874 643 -792
rect 1206 -874 1207 -792
rect 1248 -793 1249 -743
rect 1269 -874 1270 -792
rect 1290 -793 1291 -743
rect 1479 -874 1480 -792
rect 65 -795 66 -743
rect 583 -874 584 -794
rect 590 -795 591 -743
rect 1563 -874 1564 -794
rect 65 -874 66 -796
rect 828 -874 829 -796
rect 842 -797 843 -743
rect 863 -874 864 -796
rect 877 -874 878 -796
rect 1199 -874 1200 -796
rect 1262 -797 1263 -743
rect 1381 -874 1382 -796
rect 170 -799 171 -743
rect 380 -874 381 -798
rect 408 -799 409 -743
rect 492 -874 493 -798
rect 569 -799 570 -743
rect 590 -874 591 -798
rect 593 -799 594 -743
rect 1136 -874 1137 -798
rect 1185 -799 1186 -743
rect 1262 -874 1263 -798
rect 1304 -799 1305 -743
rect 1500 -874 1501 -798
rect 275 -874 276 -800
rect 796 -801 797 -743
rect 814 -801 815 -743
rect 1220 -874 1221 -800
rect 1318 -801 1319 -743
rect 1430 -874 1431 -800
rect 289 -803 290 -743
rect 352 -803 353 -743
rect 359 -803 360 -743
rect 873 -803 874 -743
rect 908 -874 909 -802
rect 1283 -874 1284 -802
rect 1325 -803 1326 -743
rect 1451 -874 1452 -802
rect 163 -805 164 -743
rect 289 -874 290 -804
rect 303 -805 304 -743
rect 303 -874 304 -804
rect 303 -805 304 -743
rect 303 -874 304 -804
rect 310 -805 311 -743
rect 758 -874 759 -804
rect 765 -874 766 -804
rect 835 -805 836 -743
rect 842 -874 843 -804
rect 849 -805 850 -743
rect 856 -805 857 -743
rect 1276 -874 1277 -804
rect 1332 -805 1333 -743
rect 1528 -874 1529 -804
rect 261 -807 262 -743
rect 1325 -874 1326 -806
rect 1339 -807 1340 -743
rect 1535 -874 1536 -806
rect 261 -874 262 -808
rect 282 -809 283 -743
rect 310 -874 311 -808
rect 387 -809 388 -743
rect 408 -874 409 -808
rect 457 -809 458 -743
rect 541 -809 542 -743
rect 569 -874 570 -808
rect 586 -874 587 -808
rect 1318 -874 1319 -808
rect 268 -811 269 -743
rect 359 -874 360 -810
rect 387 -874 388 -810
rect 422 -811 423 -743
rect 432 -811 433 -743
rect 856 -874 857 -810
rect 859 -811 860 -743
rect 1409 -811 1410 -743
rect 177 -813 178 -743
rect 422 -874 423 -812
rect 457 -874 458 -812
rect 639 -874 640 -812
rect 646 -874 647 -812
rect 702 -874 703 -812
rect 716 -874 717 -812
rect 793 -874 794 -812
rect 912 -813 913 -743
rect 1395 -813 1396 -743
rect 177 -874 178 -814
rect 212 -815 213 -743
rect 254 -815 255 -743
rect 268 -874 269 -814
rect 282 -874 283 -814
rect 436 -815 437 -743
rect 513 -815 514 -743
rect 541 -874 542 -814
rect 565 -874 566 -814
rect 1185 -874 1186 -814
rect 1192 -815 1193 -743
rect 1290 -874 1291 -814
rect 1297 -815 1298 -743
rect 1409 -874 1410 -814
rect 110 -874 111 -816
rect 1297 -874 1298 -816
rect 156 -819 157 -743
rect 254 -874 255 -818
rect 317 -819 318 -743
rect 439 -819 440 -743
rect 653 -819 654 -743
rect 1241 -874 1242 -818
rect 1255 -819 1256 -743
rect 1395 -874 1396 -818
rect 156 -874 157 -820
rect 292 -821 293 -743
rect 338 -821 339 -743
rect 338 -874 339 -820
rect 338 -821 339 -743
rect 338 -874 339 -820
rect 345 -821 346 -743
rect 618 -874 619 -820
rect 656 -821 657 -743
rect 1178 -821 1179 -743
rect 1234 -821 1235 -743
rect 1339 -874 1340 -820
rect 135 -874 136 -822
rect 1234 -874 1235 -822
rect 212 -874 213 -824
rect 219 -825 220 -743
rect 226 -825 227 -743
rect 436 -874 437 -824
rect 660 -825 661 -743
rect 789 -874 790 -824
rect 887 -825 888 -743
rect 1178 -874 1179 -824
rect 121 -827 122 -743
rect 219 -874 220 -826
rect 345 -874 346 -826
rect 548 -827 549 -743
rect 667 -827 668 -743
rect 800 -874 801 -826
rect 912 -874 913 -826
rect 1164 -827 1165 -743
rect 114 -829 115 -743
rect 121 -874 122 -828
rect 548 -874 549 -828
rect 667 -874 668 -828
rect 691 -874 692 -828
rect 695 -829 696 -743
rect 712 -829 713 -743
rect 740 -874 741 -828
rect 1360 -874 1361 -828
rect 51 -831 52 -743
rect 695 -874 696 -830
rect 751 -831 752 -743
rect 814 -874 815 -830
rect 919 -874 920 -830
rect 1150 -831 1151 -743
rect 100 -833 101 -743
rect 114 -874 115 -832
rect 170 -874 171 -832
rect 660 -874 661 -832
rect 681 -833 682 -743
rect 723 -874 724 -832
rect 772 -833 773 -743
rect 835 -874 836 -832
rect 929 -874 930 -832
rect 1311 -833 1312 -743
rect 51 -874 52 -834
rect 1311 -874 1312 -834
rect 100 -874 101 -836
rect 1248 -874 1249 -836
rect 352 -874 353 -838
rect 464 -839 465 -743
rect 681 -874 682 -838
rect 737 -839 738 -743
rect 744 -839 745 -743
rect 772 -874 773 -838
rect 786 -839 787 -743
rect 849 -874 850 -838
rect 947 -839 948 -743
rect 947 -874 948 -838
rect 947 -839 948 -743
rect 947 -874 948 -838
rect 954 -839 955 -743
rect 1003 -874 1004 -838
rect 1006 -839 1007 -743
rect 1304 -874 1305 -838
rect 72 -841 73 -743
rect 744 -874 745 -840
rect 786 -874 787 -840
rect 1213 -874 1214 -840
rect 72 -874 73 -842
rect 331 -843 332 -743
rect 415 -843 416 -743
rect 513 -874 514 -842
rect 688 -843 689 -743
rect 751 -874 752 -842
rect 933 -843 934 -743
rect 954 -874 955 -842
rect 982 -843 983 -743
rect 1038 -874 1039 -842
rect 1052 -843 1053 -743
rect 1150 -874 1151 -842
rect 296 -845 297 -743
rect 331 -874 332 -844
rect 401 -845 402 -743
rect 415 -874 416 -844
rect 688 -874 689 -844
rect 709 -874 710 -844
rect 831 -845 832 -743
rect 1052 -874 1053 -844
rect 1066 -845 1067 -743
rect 1157 -874 1158 -844
rect 324 -847 325 -743
rect 464 -874 465 -846
rect 831 -874 832 -846
rect 1255 -874 1256 -846
rect 324 -874 325 -848
rect 520 -849 521 -743
rect 891 -849 892 -743
rect 933 -874 934 -848
rect 1017 -849 1018 -743
rect 1066 -874 1067 -848
rect 1101 -849 1102 -743
rect 1192 -874 1193 -848
rect 401 -874 402 -850
rect 443 -851 444 -743
rect 506 -851 507 -743
rect 520 -874 521 -850
rect 611 -851 612 -743
rect 891 -874 892 -850
rect 926 -851 927 -743
rect 982 -874 983 -850
rect 989 -851 990 -743
rect 1101 -874 1102 -850
rect 1108 -851 1109 -743
rect 1332 -874 1333 -850
rect 86 -853 87 -743
rect 443 -874 444 -852
rect 611 -874 612 -852
rect 1143 -853 1144 -743
rect 107 -855 108 -743
rect 1143 -874 1144 -854
rect 107 -874 108 -856
rect 870 -874 871 -856
rect 989 -874 990 -856
rect 992 -857 993 -743
rect 1017 -874 1018 -856
rect 1059 -874 1060 -856
rect 1115 -857 1116 -743
rect 1164 -874 1165 -856
rect 373 -859 374 -743
rect 506 -874 507 -858
rect 1045 -859 1046 -743
rect 1108 -874 1109 -858
rect 1129 -859 1130 -743
rect 1171 -874 1172 -858
rect 373 -874 374 -860
rect 394 -861 395 -743
rect 1010 -861 1011 -743
rect 1045 -874 1046 -860
rect 1073 -861 1074 -743
rect 1115 -874 1116 -860
rect 229 -874 230 -862
rect 394 -874 395 -862
rect 968 -863 969 -743
rect 1010 -874 1011 -862
rect 1024 -863 1025 -743
rect 1073 -874 1074 -862
rect 1087 -863 1088 -743
rect 1129 -874 1130 -862
rect 478 -874 479 -864
rect 1024 -874 1025 -864
rect 1031 -865 1032 -743
rect 1087 -874 1088 -864
rect 940 -867 941 -743
rect 968 -874 969 -866
rect 975 -867 976 -743
rect 1031 -874 1032 -866
rect 674 -869 675 -743
rect 940 -874 941 -868
rect 674 -874 675 -870
rect 737 -874 738 -870
rect 898 -871 899 -743
rect 975 -874 976 -870
rect 898 -874 899 -872
rect 905 -874 906 -872
rect 30 -1035 31 -883
rect 72 -884 73 -882
rect 89 -884 90 -882
rect 114 -884 115 -882
rect 135 -884 136 -882
rect 282 -884 283 -882
rect 292 -1035 293 -883
rect 338 -884 339 -882
rect 450 -884 451 -882
rect 600 -1035 601 -883
rect 618 -884 619 -882
rect 737 -884 738 -882
rect 740 -884 741 -882
rect 1500 -884 1501 -882
rect 1521 -884 1522 -882
rect 1675 -1035 1676 -883
rect 1696 -884 1697 -882
rect 1724 -1035 1725 -883
rect 65 -886 66 -882
rect 653 -1035 654 -885
rect 663 -886 664 -882
rect 1577 -886 1578 -882
rect 1591 -886 1592 -882
rect 1608 -886 1609 -882
rect 1619 -886 1620 -882
rect 1717 -1035 1718 -885
rect 65 -1035 66 -887
rect 401 -888 402 -882
rect 422 -888 423 -882
rect 450 -1035 451 -887
rect 457 -888 458 -882
rect 929 -888 930 -882
rect 957 -1035 958 -887
rect 1535 -888 1536 -882
rect 1598 -1035 1599 -887
rect 1626 -888 1627 -882
rect 1633 -888 1634 -882
rect 1710 -1035 1711 -887
rect 72 -1035 73 -889
rect 590 -890 591 -882
rect 597 -890 598 -882
rect 611 -890 612 -882
rect 635 -1035 636 -889
rect 1549 -890 1550 -882
rect 86 -892 87 -882
rect 1591 -1035 1592 -891
rect 103 -894 104 -882
rect 142 -894 143 -882
rect 149 -894 150 -882
rect 737 -1035 738 -893
rect 761 -894 762 -882
rect 891 -894 892 -882
rect 905 -894 906 -882
rect 1528 -894 1529 -882
rect 107 -896 108 -882
rect 121 -896 122 -882
rect 135 -1035 136 -895
rect 387 -896 388 -882
rect 422 -1035 423 -895
rect 758 -896 759 -882
rect 761 -1035 762 -895
rect 891 -1035 892 -895
rect 898 -896 899 -882
rect 905 -1035 906 -895
rect 908 -896 909 -882
rect 1332 -896 1333 -882
rect 1374 -896 1375 -882
rect 1521 -1035 1522 -895
rect 110 -1035 111 -897
rect 338 -1035 339 -897
rect 387 -1035 388 -897
rect 814 -898 815 -882
rect 873 -1035 874 -897
rect 1654 -1035 1655 -897
rect 114 -1035 115 -899
rect 415 -900 416 -882
rect 457 -1035 458 -899
rect 667 -900 668 -882
rect 691 -900 692 -882
rect 1157 -900 1158 -882
rect 1206 -900 1207 -882
rect 1500 -1035 1501 -899
rect 1514 -900 1515 -882
rect 1696 -1035 1697 -899
rect 142 -1035 143 -901
rect 478 -902 479 -882
rect 499 -902 500 -882
rect 688 -1035 689 -901
rect 705 -902 706 -882
rect 1192 -902 1193 -882
rect 1220 -902 1221 -882
rect 1549 -1035 1550 -901
rect 149 -1035 150 -903
rect 177 -904 178 -882
rect 184 -904 185 -882
rect 208 -904 209 -882
rect 226 -904 227 -882
rect 268 -904 269 -882
rect 275 -904 276 -882
rect 275 -1035 276 -903
rect 275 -904 276 -882
rect 275 -1035 276 -903
rect 296 -1035 297 -903
rect 845 -1035 846 -903
rect 877 -904 878 -882
rect 1150 -904 1151 -882
rect 1234 -904 1235 -882
rect 1626 -1035 1627 -903
rect 128 -906 129 -882
rect 177 -1035 178 -905
rect 184 -1035 185 -905
rect 250 -906 251 -882
rect 254 -906 255 -882
rect 254 -1035 255 -905
rect 254 -906 255 -882
rect 254 -1035 255 -905
rect 261 -906 262 -882
rect 282 -1035 283 -905
rect 303 -906 304 -882
rect 607 -1035 608 -905
rect 611 -1035 612 -905
rect 961 -906 962 -882
rect 964 -906 965 -882
rect 1647 -1035 1648 -905
rect 128 -1035 129 -907
rect 793 -908 794 -882
rect 796 -908 797 -882
rect 1346 -908 1347 -882
rect 1395 -908 1396 -882
rect 1528 -1035 1529 -907
rect 138 -910 139 -882
rect 268 -1035 269 -909
rect 303 -1035 304 -909
rect 583 -910 584 -882
rect 586 -910 587 -882
rect 1542 -910 1543 -882
rect 163 -912 164 -882
rect 996 -912 997 -882
rect 1038 -912 1039 -882
rect 1157 -1035 1158 -911
rect 1248 -912 1249 -882
rect 1374 -1035 1375 -911
rect 1430 -912 1431 -882
rect 1535 -1035 1536 -911
rect 163 -1035 164 -913
rect 324 -914 325 -882
rect 331 -914 332 -882
rect 401 -1035 402 -913
rect 415 -1035 416 -913
rect 716 -914 717 -882
rect 768 -1035 769 -913
rect 1633 -1035 1634 -913
rect 93 -916 94 -882
rect 324 -1035 325 -915
rect 373 -916 374 -882
rect 499 -1035 500 -915
rect 506 -916 507 -882
rect 506 -1035 507 -915
rect 506 -916 507 -882
rect 506 -1035 507 -915
rect 548 -916 549 -882
rect 667 -1035 668 -915
rect 786 -916 787 -882
rect 1584 -916 1585 -882
rect 86 -1035 87 -917
rect 93 -1035 94 -917
rect 166 -918 167 -882
rect 513 -918 514 -882
rect 548 -1035 549 -917
rect 1682 -1035 1683 -917
rect 170 -920 171 -882
rect 481 -920 482 -882
rect 513 -1035 514 -919
rect 901 -1035 902 -919
rect 912 -920 913 -882
rect 926 -920 927 -882
rect 933 -920 934 -882
rect 996 -1035 997 -919
rect 1059 -920 1060 -882
rect 1465 -920 1466 -882
rect 1486 -920 1487 -882
rect 1605 -1035 1606 -919
rect 170 -1035 171 -921
rect 240 -922 241 -882
rect 247 -1035 248 -921
rect 289 -922 290 -882
rect 310 -922 311 -882
rect 593 -1035 594 -921
rect 646 -922 647 -882
rect 649 -986 650 -921
rect 733 -1035 734 -921
rect 1486 -1035 1487 -921
rect 1493 -922 1494 -882
rect 1668 -1035 1669 -921
rect 191 -924 192 -882
rect 660 -924 661 -882
rect 765 -924 766 -882
rect 786 -1035 787 -923
rect 810 -1035 811 -923
rect 1703 -1035 1704 -923
rect 79 -926 80 -882
rect 191 -1035 192 -925
rect 198 -926 199 -882
rect 660 -1035 661 -925
rect 765 -1035 766 -925
rect 1325 -926 1326 -882
rect 1339 -926 1340 -882
rect 1465 -1035 1466 -925
rect 79 -1035 80 -927
rect 562 -928 563 -882
rect 569 -928 570 -882
rect 569 -1035 570 -927
rect 569 -928 570 -882
rect 569 -1035 570 -927
rect 576 -928 577 -882
rect 702 -1035 703 -927
rect 856 -928 857 -882
rect 912 -1035 913 -927
rect 919 -928 920 -882
rect 961 -1035 962 -927
rect 968 -928 969 -882
rect 971 -986 972 -927
rect 975 -928 976 -882
rect 1038 -1035 1039 -927
rect 1062 -928 1063 -882
rect 1388 -928 1389 -882
rect 1437 -928 1438 -882
rect 1584 -1035 1585 -927
rect 124 -1035 125 -929
rect 198 -1035 199 -929
rect 205 -1035 206 -929
rect 621 -1035 622 -929
rect 646 -1035 647 -929
rect 1094 -930 1095 -882
rect 1101 -930 1102 -882
rect 1234 -1035 1235 -929
rect 1262 -930 1263 -882
rect 1395 -1035 1396 -929
rect 1444 -930 1445 -882
rect 1661 -1035 1662 -929
rect 226 -1035 227 -931
rect 579 -932 580 -882
rect 583 -1035 584 -931
rect 695 -932 696 -882
rect 772 -932 773 -882
rect 1388 -1035 1389 -931
rect 1458 -932 1459 -882
rect 1619 -1035 1620 -931
rect 229 -934 230 -882
rect 1143 -934 1144 -882
rect 1150 -1035 1151 -933
rect 1381 -934 1382 -882
rect 1458 -1035 1459 -933
rect 1507 -934 1508 -882
rect 121 -1035 122 -935
rect 1507 -1035 1508 -935
rect 233 -938 234 -882
rect 1570 -938 1571 -882
rect 89 -1035 90 -939
rect 233 -1035 234 -939
rect 236 -940 237 -882
rect 1640 -1035 1641 -939
rect 240 -1035 241 -941
rect 352 -942 353 -882
rect 373 -1035 374 -941
rect 408 -942 409 -882
rect 436 -942 437 -882
rect 1220 -1035 1221 -941
rect 1255 -942 1256 -882
rect 1570 -1035 1571 -941
rect 261 -1035 262 -943
rect 429 -944 430 -882
rect 436 -1035 437 -943
rect 723 -944 724 -882
rect 730 -944 731 -882
rect 772 -1035 773 -943
rect 856 -1035 857 -943
rect 1514 -1035 1515 -943
rect 289 -1035 290 -945
rect 1248 -1035 1249 -945
rect 1255 -1035 1256 -945
rect 1269 -946 1270 -882
rect 1276 -946 1277 -882
rect 1276 -1035 1277 -945
rect 1276 -946 1277 -882
rect 1276 -1035 1277 -945
rect 1297 -946 1298 -882
rect 1689 -1035 1690 -945
rect 37 -948 38 -882
rect 1297 -1035 1298 -947
rect 1304 -948 1305 -882
rect 1444 -1035 1445 -947
rect 313 -1035 314 -949
rect 331 -1035 332 -949
rect 345 -950 346 -882
rect 562 -1035 563 -949
rect 576 -1035 577 -949
rect 632 -950 633 -882
rect 709 -950 710 -882
rect 730 -1035 731 -949
rect 863 -950 864 -882
rect 926 -1035 927 -949
rect 940 -950 941 -882
rect 1143 -1035 1144 -949
rect 1178 -950 1179 -882
rect 1304 -1035 1305 -949
rect 1346 -1035 1347 -949
rect 1367 -950 1368 -882
rect 1381 -1035 1382 -949
rect 1612 -950 1613 -882
rect 317 -1035 318 -951
rect 467 -952 468 -882
rect 474 -1035 475 -951
rect 674 -952 675 -882
rect 800 -952 801 -882
rect 940 -1035 941 -951
rect 968 -1035 969 -951
rect 1017 -952 1018 -882
rect 1031 -952 1032 -882
rect 1339 -1035 1340 -951
rect 1353 -952 1354 -882
rect 1493 -1035 1494 -951
rect 345 -1035 346 -953
rect 366 -954 367 -882
rect 394 -954 395 -882
rect 408 -1035 409 -953
rect 429 -1035 430 -953
rect 625 -954 626 -882
rect 632 -1035 633 -953
rect 814 -1035 815 -953
rect 849 -954 850 -882
rect 863 -1035 864 -953
rect 870 -954 871 -882
rect 1437 -1035 1438 -953
rect 107 -1035 108 -955
rect 849 -1035 850 -955
rect 870 -1035 871 -955
rect 1178 -1035 1179 -955
rect 1199 -956 1200 -882
rect 1325 -1035 1326 -955
rect 1353 -1035 1354 -955
rect 1409 -956 1410 -882
rect 352 -1035 353 -957
rect 380 -958 381 -882
rect 394 -1035 395 -957
rect 723 -1035 724 -957
rect 800 -1035 801 -957
rect 821 -958 822 -882
rect 877 -1035 878 -957
rect 1416 -958 1417 -882
rect 366 -1035 367 -959
rect 471 -960 472 -882
rect 478 -1035 479 -959
rect 555 -960 556 -882
rect 604 -960 605 -882
rect 709 -1035 710 -959
rect 751 -960 752 -882
rect 821 -1035 822 -959
rect 884 -960 885 -882
rect 887 -986 888 -959
rect 898 -1035 899 -959
rect 1241 -960 1242 -882
rect 1283 -960 1284 -882
rect 1409 -1035 1410 -959
rect 37 -1035 38 -961
rect 471 -1035 472 -961
rect 520 -962 521 -882
rect 555 -1035 556 -961
rect 604 -1035 605 -961
rect 1577 -1035 1578 -961
rect 380 -1035 381 -963
rect 485 -964 486 -882
rect 492 -964 493 -882
rect 520 -1035 521 -963
rect 527 -964 528 -882
rect 751 -1035 752 -963
rect 884 -1035 885 -963
rect 982 -964 983 -882
rect 1003 -964 1004 -882
rect 1094 -1035 1095 -963
rect 1115 -964 1116 -882
rect 1262 -1035 1263 -963
rect 1290 -964 1291 -882
rect 1416 -1035 1417 -963
rect 44 -966 45 -882
rect 485 -1035 486 -965
rect 534 -966 535 -882
rect 919 -1035 920 -965
rect 947 -966 948 -882
rect 1031 -1035 1032 -965
rect 1052 -966 1053 -882
rect 1199 -1035 1200 -965
rect 1213 -966 1214 -882
rect 1612 -1035 1613 -965
rect 44 -1035 45 -967
rect 54 -968 55 -882
rect 58 -968 59 -882
rect 492 -1035 493 -967
rect 537 -1035 538 -967
rect 933 -1035 934 -967
rect 975 -1035 976 -967
rect 1430 -1035 1431 -967
rect 54 -1035 55 -969
rect 1556 -970 1557 -882
rect 58 -1035 59 -971
rect 1136 -972 1137 -882
rect 1164 -972 1165 -882
rect 1290 -1035 1291 -971
rect 100 -974 101 -882
rect 1556 -1035 1557 -973
rect 23 -976 24 -882
rect 100 -1035 101 -975
rect 219 -976 220 -882
rect 947 -1035 948 -975
rect 978 -1035 979 -975
rect 1601 -976 1602 -882
rect 359 -978 360 -882
rect 527 -1035 528 -977
rect 551 -1035 552 -977
rect 744 -978 745 -882
rect 880 -978 881 -882
rect 1115 -1035 1116 -977
rect 1129 -978 1130 -882
rect 1269 -1035 1270 -977
rect 212 -980 213 -882
rect 359 -1035 360 -979
rect 443 -980 444 -882
rect 716 -1035 717 -979
rect 744 -1035 745 -979
rect 992 -1035 993 -979
rect 1003 -1035 1004 -979
rect 1108 -980 1109 -882
rect 1122 -980 1123 -882
rect 1129 -1035 1130 -979
rect 1164 -1035 1165 -979
rect 1171 -980 1172 -882
rect 156 -982 157 -882
rect 443 -1035 444 -981
rect 467 -1035 468 -981
rect 1241 -1035 1242 -981
rect 156 -1035 157 -983
rect 793 -1035 794 -983
rect 835 -984 836 -882
rect 1122 -1035 1123 -983
rect 212 -1035 213 -985
rect 541 -986 542 -882
rect 614 -986 615 -882
rect 674 -1035 675 -985
rect 835 -1035 836 -985
rect 842 -986 843 -882
rect 1017 -1035 1018 -985
rect 1024 -986 1025 -882
rect 1136 -1035 1137 -985
rect 541 -1035 542 -987
rect 597 -1035 598 -987
rect 618 -1035 619 -987
rect 695 -1035 696 -987
rect 796 -1035 797 -987
rect 1024 -1035 1025 -987
rect 1045 -988 1046 -882
rect 1171 -1035 1172 -987
rect 625 -1035 626 -989
rect 681 -990 682 -882
rect 842 -1035 843 -989
rect 1332 -1035 1333 -989
rect 639 -992 640 -882
rect 1367 -1035 1368 -991
rect 639 -1035 640 -993
rect 880 -1035 881 -993
rect 954 -994 955 -882
rect 1045 -1035 1046 -993
rect 1062 -1035 1063 -993
rect 1472 -994 1473 -882
rect 681 -1035 682 -995
rect 1283 -1035 1284 -995
rect 789 -998 790 -882
rect 1472 -1035 1473 -997
rect 954 -1035 955 -999
rect 1563 -1000 1564 -882
rect 989 -1002 990 -882
rect 1052 -1035 1053 -1001
rect 1066 -1002 1067 -882
rect 1192 -1035 1193 -1001
rect 1451 -1002 1452 -882
rect 1563 -1035 1564 -1001
rect 989 -1035 990 -1003
rect 1542 -1035 1543 -1003
rect 1010 -1006 1011 -882
rect 1101 -1035 1102 -1005
rect 1311 -1006 1312 -882
rect 1451 -1035 1452 -1005
rect 534 -1035 535 -1007
rect 1311 -1035 1312 -1007
rect 1066 -1035 1067 -1009
rect 1402 -1010 1403 -882
rect 1073 -1012 1074 -882
rect 1206 -1035 1207 -1011
rect 1402 -1035 1403 -1011
rect 1423 -1012 1424 -882
rect 628 -1014 629 -882
rect 1073 -1035 1074 -1013
rect 1080 -1014 1081 -882
rect 1213 -1035 1214 -1013
rect 779 -1016 780 -882
rect 1080 -1035 1081 -1015
rect 779 -1035 780 -1017
rect 807 -1018 808 -882
rect 828 -1018 829 -882
rect 1423 -1035 1424 -1017
rect 807 -1035 808 -1019
rect 1010 -1035 1011 -1019
rect 828 -1035 829 -1021
rect 1360 -1022 1361 -882
rect 1360 -1035 1361 -1023
rect 1479 -1024 1480 -882
rect 1318 -1026 1319 -882
rect 1479 -1035 1480 -1025
rect 1185 -1028 1186 -882
rect 1318 -1035 1319 -1027
rect 1185 -1035 1186 -1029
rect 1227 -1030 1228 -882
rect 1087 -1032 1088 -882
rect 1227 -1035 1228 -1031
rect 201 -1035 202 -1033
rect 1087 -1035 1088 -1033
rect 44 -1186 45 -1044
rect 240 -1045 241 -1043
rect 261 -1045 262 -1043
rect 632 -1045 633 -1043
rect 653 -1045 654 -1043
rect 653 -1186 654 -1044
rect 653 -1045 654 -1043
rect 653 -1186 654 -1044
rect 681 -1045 682 -1043
rect 1143 -1045 1144 -1043
rect 1710 -1045 1711 -1043
rect 1731 -1186 1732 -1044
rect 65 -1047 66 -1043
rect 488 -1186 489 -1046
rect 499 -1047 500 -1043
rect 632 -1186 633 -1046
rect 681 -1186 682 -1046
rect 695 -1047 696 -1043
rect 719 -1186 720 -1046
rect 1521 -1047 1522 -1043
rect 1724 -1047 1725 -1043
rect 1724 -1186 1725 -1046
rect 1724 -1047 1725 -1043
rect 1724 -1186 1725 -1046
rect 65 -1186 66 -1048
rect 544 -1186 545 -1048
rect 579 -1186 580 -1048
rect 1367 -1049 1368 -1043
rect 86 -1051 87 -1043
rect 940 -1051 941 -1043
rect 957 -1051 958 -1043
rect 1626 -1051 1627 -1043
rect 89 -1053 90 -1043
rect 1514 -1053 1515 -1043
rect 1626 -1186 1627 -1052
rect 1668 -1053 1669 -1043
rect 93 -1055 94 -1043
rect 187 -1186 188 -1054
rect 198 -1055 199 -1043
rect 401 -1055 402 -1043
rect 408 -1055 409 -1043
rect 534 -1055 535 -1043
rect 590 -1055 591 -1043
rect 1500 -1055 1501 -1043
rect 51 -1057 52 -1043
rect 590 -1186 591 -1056
rect 597 -1057 598 -1043
rect 716 -1057 717 -1043
rect 723 -1057 724 -1043
rect 1549 -1057 1550 -1043
rect 51 -1186 52 -1058
rect 555 -1059 556 -1043
rect 600 -1059 601 -1043
rect 1010 -1059 1011 -1043
rect 1062 -1059 1063 -1043
rect 1521 -1186 1522 -1058
rect 93 -1186 94 -1060
rect 443 -1061 444 -1043
rect 450 -1061 451 -1043
rect 499 -1186 500 -1060
rect 513 -1061 514 -1043
rect 555 -1186 556 -1060
rect 569 -1061 570 -1043
rect 600 -1186 601 -1060
rect 614 -1186 615 -1060
rect 919 -1061 920 -1043
rect 940 -1186 941 -1060
rect 1038 -1061 1039 -1043
rect 1069 -1061 1070 -1043
rect 1696 -1061 1697 -1043
rect 54 -1063 55 -1043
rect 443 -1186 444 -1062
rect 450 -1186 451 -1062
rect 520 -1063 521 -1043
rect 527 -1063 528 -1043
rect 716 -1186 717 -1062
rect 726 -1063 727 -1043
rect 730 -1063 731 -1043
rect 751 -1063 752 -1043
rect 807 -1063 808 -1043
rect 810 -1063 811 -1043
rect 1045 -1063 1046 -1043
rect 1129 -1063 1130 -1043
rect 1129 -1186 1130 -1062
rect 1129 -1063 1130 -1043
rect 1129 -1186 1130 -1062
rect 1143 -1186 1144 -1062
rect 1234 -1063 1235 -1043
rect 1360 -1063 1361 -1043
rect 1549 -1186 1550 -1062
rect 100 -1065 101 -1043
rect 289 -1065 290 -1043
rect 292 -1065 293 -1043
rect 604 -1065 605 -1043
rect 702 -1065 703 -1043
rect 730 -1186 731 -1064
rect 751 -1186 752 -1064
rect 1381 -1065 1382 -1043
rect 1500 -1186 1501 -1064
rect 1612 -1065 1613 -1043
rect 103 -1186 104 -1066
rect 1388 -1067 1389 -1043
rect 1612 -1186 1613 -1066
rect 1654 -1067 1655 -1043
rect 107 -1069 108 -1043
rect 415 -1069 416 -1043
rect 464 -1186 465 -1068
rect 947 -1069 948 -1043
rect 971 -1186 972 -1068
rect 1048 -1186 1049 -1068
rect 1234 -1186 1235 -1068
rect 1650 -1186 1651 -1068
rect 107 -1186 108 -1070
rect 747 -1186 748 -1070
rect 758 -1071 759 -1043
rect 1227 -1071 1228 -1043
rect 1276 -1071 1277 -1043
rect 1360 -1186 1361 -1070
rect 1367 -1186 1368 -1070
rect 1465 -1071 1466 -1043
rect 89 -1186 90 -1072
rect 1465 -1186 1466 -1072
rect 110 -1075 111 -1043
rect 1479 -1075 1480 -1043
rect 121 -1077 122 -1043
rect 1220 -1077 1221 -1043
rect 1227 -1186 1228 -1076
rect 1290 -1077 1291 -1043
rect 1381 -1186 1382 -1076
rect 1535 -1077 1536 -1043
rect 121 -1186 122 -1078
rect 436 -1079 437 -1043
rect 478 -1079 479 -1043
rect 534 -1186 535 -1078
rect 621 -1079 622 -1043
rect 1276 -1186 1277 -1078
rect 1290 -1186 1291 -1078
rect 1409 -1079 1410 -1043
rect 1479 -1186 1480 -1078
rect 1640 -1079 1641 -1043
rect 128 -1081 129 -1043
rect 436 -1186 437 -1080
rect 506 -1081 507 -1043
rect 527 -1186 528 -1080
rect 621 -1186 622 -1080
rect 1122 -1081 1123 -1043
rect 1388 -1186 1389 -1080
rect 1430 -1081 1431 -1043
rect 1640 -1186 1641 -1080
rect 1675 -1081 1676 -1043
rect 128 -1186 129 -1082
rect 744 -1083 745 -1043
rect 768 -1083 769 -1043
rect 1339 -1083 1340 -1043
rect 1402 -1083 1403 -1043
rect 1654 -1186 1655 -1082
rect 135 -1085 136 -1043
rect 467 -1085 468 -1043
rect 506 -1186 507 -1084
rect 1241 -1085 1242 -1043
rect 1255 -1085 1256 -1043
rect 1430 -1186 1431 -1084
rect 1619 -1085 1620 -1043
rect 1675 -1186 1676 -1084
rect 135 -1186 136 -1086
rect 205 -1087 206 -1043
rect 208 -1186 209 -1086
rect 1311 -1087 1312 -1043
rect 1339 -1186 1340 -1086
rect 1374 -1087 1375 -1043
rect 1409 -1186 1410 -1086
rect 1451 -1087 1452 -1043
rect 142 -1089 143 -1043
rect 569 -1186 570 -1088
rect 628 -1089 629 -1043
rect 1451 -1186 1452 -1088
rect 142 -1186 143 -1090
rect 149 -1091 150 -1043
rect 166 -1186 167 -1090
rect 198 -1186 199 -1090
rect 219 -1186 220 -1090
rect 247 -1091 248 -1043
rect 261 -1186 262 -1090
rect 828 -1186 829 -1090
rect 845 -1091 846 -1043
rect 1150 -1091 1151 -1043
rect 1241 -1186 1242 -1090
rect 1297 -1091 1298 -1043
rect 1311 -1186 1312 -1090
rect 1437 -1091 1438 -1043
rect 149 -1186 150 -1092
rect 303 -1093 304 -1043
rect 310 -1186 311 -1092
rect 331 -1093 332 -1043
rect 352 -1093 353 -1043
rect 352 -1186 353 -1092
rect 352 -1093 353 -1043
rect 352 -1186 353 -1092
rect 359 -1093 360 -1043
rect 415 -1186 416 -1092
rect 513 -1186 514 -1092
rect 576 -1093 577 -1043
rect 702 -1186 703 -1092
rect 1423 -1093 1424 -1043
rect 1437 -1186 1438 -1092
rect 1458 -1093 1459 -1043
rect 170 -1095 171 -1043
rect 408 -1186 409 -1094
rect 516 -1186 517 -1094
rect 758 -1186 759 -1094
rect 786 -1095 787 -1043
rect 842 -1095 843 -1043
rect 859 -1095 860 -1043
rect 1514 -1186 1515 -1094
rect 170 -1186 171 -1096
rect 191 -1097 192 -1043
rect 212 -1097 213 -1043
rect 303 -1186 304 -1096
rect 331 -1186 332 -1096
rect 345 -1097 346 -1043
rect 359 -1186 360 -1096
rect 485 -1097 486 -1043
rect 520 -1186 521 -1096
rect 541 -1097 542 -1043
rect 733 -1097 734 -1043
rect 1220 -1186 1221 -1096
rect 1297 -1186 1298 -1096
rect 1416 -1097 1417 -1043
rect 1458 -1186 1459 -1096
rect 1472 -1097 1473 -1043
rect 47 -1099 48 -1043
rect 541 -1186 542 -1098
rect 744 -1186 745 -1098
rect 996 -1099 997 -1043
rect 1010 -1186 1011 -1098
rect 1094 -1099 1095 -1043
rect 1122 -1186 1123 -1098
rect 1178 -1099 1179 -1043
rect 1346 -1099 1347 -1043
rect 1423 -1186 1424 -1098
rect 1472 -1186 1473 -1098
rect 1528 -1099 1529 -1043
rect 79 -1101 80 -1043
rect 191 -1186 192 -1100
rect 212 -1186 213 -1100
rect 254 -1101 255 -1043
rect 282 -1101 283 -1043
rect 345 -1186 346 -1100
rect 366 -1101 367 -1043
rect 474 -1101 475 -1043
rect 485 -1186 486 -1100
rect 1535 -1186 1536 -1100
rect 79 -1186 80 -1102
rect 1556 -1103 1557 -1043
rect 163 -1105 164 -1043
rect 254 -1186 255 -1104
rect 275 -1105 276 -1043
rect 282 -1186 283 -1104
rect 289 -1186 290 -1104
rect 317 -1105 318 -1043
rect 366 -1186 367 -1104
rect 551 -1105 552 -1043
rect 793 -1105 794 -1043
rect 1584 -1105 1585 -1043
rect 114 -1107 115 -1043
rect 317 -1186 318 -1106
rect 380 -1107 381 -1043
rect 695 -1186 696 -1106
rect 807 -1186 808 -1106
rect 1073 -1107 1074 -1043
rect 1115 -1107 1116 -1043
rect 1584 -1186 1585 -1106
rect 114 -1186 115 -1108
rect 779 -1109 780 -1043
rect 842 -1186 843 -1108
rect 1045 -1186 1046 -1108
rect 1073 -1186 1074 -1108
rect 1087 -1109 1088 -1043
rect 1115 -1186 1116 -1108
rect 1171 -1109 1172 -1043
rect 1178 -1186 1179 -1108
rect 1213 -1109 1214 -1043
rect 1332 -1109 1333 -1043
rect 1346 -1186 1347 -1108
rect 1374 -1186 1375 -1108
rect 1605 -1109 1606 -1043
rect 156 -1111 157 -1043
rect 275 -1186 276 -1110
rect 296 -1111 297 -1043
rect 296 -1186 297 -1110
rect 296 -1111 297 -1043
rect 296 -1186 297 -1110
rect 380 -1186 381 -1110
rect 467 -1186 468 -1110
rect 723 -1186 724 -1110
rect 1213 -1186 1214 -1110
rect 1528 -1186 1529 -1110
rect 1542 -1111 1543 -1043
rect 1556 -1186 1557 -1110
rect 1577 -1111 1578 -1043
rect 156 -1186 157 -1112
rect 646 -1113 647 -1043
rect 772 -1113 773 -1043
rect 779 -1186 780 -1112
rect 849 -1113 850 -1043
rect 1332 -1186 1333 -1112
rect 1542 -1186 1543 -1112
rect 1661 -1113 1662 -1043
rect 75 -1186 76 -1114
rect 849 -1186 850 -1114
rect 856 -1115 857 -1043
rect 1094 -1186 1095 -1114
rect 1150 -1186 1151 -1114
rect 1248 -1115 1249 -1043
rect 177 -1117 178 -1043
rect 625 -1117 626 -1043
rect 646 -1186 647 -1116
rect 667 -1117 668 -1043
rect 674 -1117 675 -1043
rect 772 -1186 773 -1116
rect 835 -1117 836 -1043
rect 856 -1186 857 -1116
rect 870 -1117 871 -1043
rect 1059 -1186 1060 -1116
rect 1164 -1117 1165 -1043
rect 1171 -1186 1172 -1116
rect 1248 -1186 1249 -1116
rect 1325 -1117 1326 -1043
rect 177 -1186 178 -1118
rect 1664 -1186 1665 -1118
rect 201 -1121 202 -1043
rect 1087 -1186 1088 -1120
rect 1164 -1186 1165 -1120
rect 1262 -1121 1263 -1043
rect 201 -1186 202 -1122
rect 457 -1123 458 -1043
rect 537 -1123 538 -1043
rect 674 -1186 675 -1122
rect 821 -1123 822 -1043
rect 870 -1186 871 -1122
rect 873 -1123 874 -1043
rect 1493 -1123 1494 -1043
rect 205 -1186 206 -1124
rect 1605 -1186 1606 -1124
rect 236 -1186 237 -1126
rect 1255 -1186 1256 -1126
rect 1353 -1127 1354 -1043
rect 1493 -1186 1494 -1126
rect 240 -1186 241 -1128
rect 639 -1129 640 -1043
rect 667 -1186 668 -1128
rect 688 -1129 689 -1043
rect 821 -1186 822 -1128
rect 1101 -1129 1102 -1043
rect 1185 -1129 1186 -1043
rect 1262 -1186 1263 -1128
rect 1353 -1186 1354 -1128
rect 1395 -1129 1396 -1043
rect 58 -1131 59 -1043
rect 688 -1186 689 -1130
rect 835 -1186 836 -1130
rect 968 -1131 969 -1043
rect 975 -1186 976 -1130
rect 1031 -1131 1032 -1043
rect 1038 -1186 1039 -1130
rect 1206 -1131 1207 -1043
rect 1395 -1186 1396 -1130
rect 1444 -1131 1445 -1043
rect 58 -1186 59 -1132
rect 663 -1186 664 -1132
rect 877 -1133 878 -1043
rect 1619 -1186 1620 -1132
rect 247 -1186 248 -1134
rect 268 -1135 269 -1043
rect 387 -1135 388 -1043
rect 604 -1186 605 -1134
rect 625 -1186 626 -1134
rect 954 -1135 955 -1043
rect 978 -1135 979 -1043
rect 1577 -1186 1578 -1134
rect 163 -1186 164 -1136
rect 268 -1186 269 -1136
rect 394 -1137 395 -1043
rect 880 -1137 881 -1043
rect 894 -1186 895 -1136
rect 1416 -1186 1417 -1136
rect 1444 -1186 1445 -1136
rect 1507 -1137 1508 -1043
rect 226 -1139 227 -1043
rect 387 -1186 388 -1138
rect 394 -1186 395 -1138
rect 754 -1186 755 -1138
rect 877 -1186 878 -1138
rect 884 -1139 885 -1043
rect 898 -1139 899 -1043
rect 1633 -1139 1634 -1043
rect 30 -1141 31 -1043
rect 226 -1186 227 -1140
rect 401 -1186 402 -1140
rect 593 -1141 594 -1043
rect 639 -1186 640 -1140
rect 737 -1141 738 -1043
rect 898 -1186 899 -1140
rect 1507 -1186 1508 -1140
rect 1598 -1141 1599 -1043
rect 1633 -1186 1634 -1140
rect 30 -1186 31 -1142
rect 583 -1143 584 -1043
rect 709 -1143 710 -1043
rect 737 -1186 738 -1142
rect 905 -1143 906 -1043
rect 905 -1186 906 -1142
rect 905 -1143 906 -1043
rect 905 -1186 906 -1142
rect 912 -1143 913 -1043
rect 968 -1186 969 -1142
rect 989 -1143 990 -1043
rect 1689 -1143 1690 -1043
rect 233 -1145 234 -1043
rect 583 -1186 584 -1144
rect 709 -1186 710 -1144
rect 1066 -1145 1067 -1043
rect 1101 -1186 1102 -1144
rect 1157 -1145 1158 -1043
rect 1563 -1145 1564 -1043
rect 1598 -1186 1599 -1144
rect 422 -1147 423 -1043
rect 786 -1186 787 -1146
rect 912 -1186 913 -1146
rect 926 -1147 927 -1043
rect 933 -1147 934 -1043
rect 1325 -1186 1326 -1146
rect 1563 -1186 1564 -1146
rect 1591 -1147 1592 -1043
rect 422 -1186 423 -1148
rect 548 -1149 549 -1043
rect 726 -1186 727 -1148
rect 926 -1186 927 -1148
rect 947 -1186 948 -1148
rect 982 -1149 983 -1043
rect 989 -1186 990 -1148
rect 1402 -1186 1403 -1148
rect 1591 -1186 1592 -1148
rect 1647 -1149 1648 -1043
rect 324 -1151 325 -1043
rect 548 -1186 549 -1150
rect 765 -1151 766 -1043
rect 933 -1186 934 -1150
rect 954 -1186 955 -1150
rect 1570 -1151 1571 -1043
rect 1647 -1186 1648 -1150
rect 1717 -1151 1718 -1043
rect 100 -1186 101 -1152
rect 324 -1186 325 -1152
rect 429 -1153 430 -1043
rect 793 -1186 794 -1152
rect 814 -1153 815 -1043
rect 982 -1186 983 -1152
rect 992 -1153 993 -1043
rect 1206 -1186 1207 -1152
rect 1570 -1186 1571 -1152
rect 1682 -1153 1683 -1043
rect 373 -1155 374 -1043
rect 429 -1186 430 -1154
rect 457 -1186 458 -1154
rect 611 -1155 612 -1043
rect 814 -1186 815 -1154
rect 863 -1155 864 -1043
rect 919 -1186 920 -1154
rect 961 -1155 962 -1043
rect 992 -1186 993 -1154
rect 1486 -1155 1487 -1043
rect 373 -1186 374 -1156
rect 660 -1157 661 -1043
rect 800 -1157 801 -1043
rect 863 -1186 864 -1156
rect 996 -1186 997 -1156
rect 1024 -1157 1025 -1043
rect 1031 -1186 1032 -1156
rect 1108 -1157 1109 -1043
rect 1157 -1186 1158 -1156
rect 1283 -1157 1284 -1043
rect 1486 -1186 1487 -1156
rect 1703 -1157 1704 -1043
rect 338 -1159 339 -1043
rect 800 -1186 801 -1158
rect 831 -1159 832 -1043
rect 961 -1186 962 -1158
rect 1003 -1159 1004 -1043
rect 1185 -1186 1186 -1158
rect 1283 -1186 1284 -1158
rect 1318 -1159 1319 -1043
rect 184 -1161 185 -1043
rect 338 -1186 339 -1160
rect 471 -1161 472 -1043
rect 884 -1186 885 -1160
rect 957 -1186 958 -1160
rect 1318 -1186 1319 -1160
rect 37 -1163 38 -1043
rect 471 -1186 472 -1162
rect 562 -1163 563 -1043
rect 765 -1186 766 -1162
rect 1003 -1186 1004 -1162
rect 1052 -1163 1053 -1043
rect 37 -1186 38 -1164
rect 72 -1165 73 -1043
rect 124 -1186 125 -1164
rect 1052 -1186 1053 -1164
rect 184 -1186 185 -1166
rect 478 -1186 479 -1166
rect 492 -1167 493 -1043
rect 562 -1186 563 -1166
rect 611 -1186 612 -1166
rect 891 -1167 892 -1043
rect 1017 -1167 1018 -1043
rect 1066 -1186 1067 -1166
rect 492 -1186 493 -1168
rect 761 -1169 762 -1043
rect 1017 -1186 1018 -1168
rect 1080 -1169 1081 -1043
rect 635 -1171 636 -1043
rect 1108 -1186 1109 -1170
rect 660 -1186 661 -1172
rect 1199 -1173 1200 -1043
rect 901 -1186 902 -1174
rect 1199 -1186 1200 -1174
rect 1024 -1186 1025 -1176
rect 1136 -1177 1137 -1043
rect 1080 -1186 1081 -1178
rect 1269 -1179 1270 -1043
rect 1136 -1186 1137 -1180
rect 1192 -1181 1193 -1043
rect 1269 -1186 1270 -1180
rect 1304 -1181 1305 -1043
rect 597 -1186 598 -1182
rect 1192 -1186 1193 -1182
rect 607 -1185 608 -1043
rect 1304 -1186 1305 -1184
rect 23 -1317 24 -1195
rect 65 -1196 66 -1194
rect 79 -1317 80 -1195
rect 100 -1317 101 -1195
rect 124 -1196 125 -1194
rect 1115 -1196 1116 -1194
rect 1318 -1196 1319 -1194
rect 1318 -1317 1319 -1195
rect 1318 -1196 1319 -1194
rect 1318 -1317 1319 -1195
rect 1486 -1196 1487 -1194
rect 1689 -1317 1690 -1195
rect 1717 -1317 1718 -1195
rect 1724 -1196 1725 -1194
rect 1731 -1196 1732 -1194
rect 1738 -1317 1739 -1195
rect 30 -1198 31 -1194
rect 89 -1198 90 -1194
rect 93 -1198 94 -1194
rect 145 -1317 146 -1197
rect 149 -1198 150 -1194
rect 205 -1198 206 -1194
rect 208 -1198 209 -1194
rect 793 -1198 794 -1194
rect 810 -1317 811 -1197
rect 835 -1198 836 -1194
rect 873 -1198 874 -1194
rect 1598 -1198 1599 -1194
rect 1605 -1198 1606 -1194
rect 1682 -1317 1683 -1197
rect 30 -1317 31 -1199
rect 488 -1200 489 -1194
rect 506 -1317 507 -1199
rect 695 -1200 696 -1194
rect 723 -1200 724 -1194
rect 1185 -1200 1186 -1194
rect 1451 -1200 1452 -1194
rect 1486 -1317 1487 -1199
rect 1500 -1200 1501 -1194
rect 1598 -1317 1599 -1199
rect 1619 -1200 1620 -1194
rect 1668 -1317 1669 -1199
rect 1675 -1200 1676 -1194
rect 1731 -1317 1732 -1199
rect 58 -1202 59 -1194
rect 121 -1202 122 -1194
rect 135 -1202 136 -1194
rect 513 -1202 514 -1194
rect 541 -1317 542 -1201
rect 709 -1202 710 -1194
rect 744 -1202 745 -1194
rect 1136 -1202 1137 -1194
rect 1185 -1317 1186 -1201
rect 1325 -1202 1326 -1194
rect 1465 -1202 1466 -1194
rect 1619 -1317 1620 -1201
rect 1633 -1202 1634 -1194
rect 1633 -1317 1634 -1201
rect 1633 -1202 1634 -1194
rect 1633 -1317 1634 -1201
rect 1654 -1202 1655 -1194
rect 1675 -1317 1676 -1201
rect 58 -1317 59 -1203
rect 247 -1204 248 -1194
rect 250 -1317 251 -1203
rect 352 -1204 353 -1194
rect 380 -1204 381 -1194
rect 723 -1317 724 -1203
rect 744 -1317 745 -1203
rect 779 -1204 780 -1194
rect 814 -1204 815 -1194
rect 898 -1204 899 -1194
rect 901 -1204 902 -1194
rect 1444 -1204 1445 -1194
rect 1591 -1204 1592 -1194
rect 1605 -1317 1606 -1203
rect 1661 -1204 1662 -1194
rect 1724 -1317 1725 -1203
rect 65 -1317 66 -1205
rect 201 -1206 202 -1194
rect 205 -1317 206 -1205
rect 576 -1206 577 -1194
rect 593 -1317 594 -1205
rect 1402 -1206 1403 -1194
rect 1416 -1206 1417 -1194
rect 1465 -1317 1466 -1205
rect 1542 -1206 1543 -1194
rect 1661 -1317 1662 -1205
rect 96 -1317 97 -1207
rect 1514 -1208 1515 -1194
rect 1528 -1208 1529 -1194
rect 1542 -1317 1543 -1207
rect 121 -1317 122 -1209
rect 1521 -1210 1522 -1194
rect 135 -1317 136 -1211
rect 359 -1212 360 -1194
rect 380 -1317 381 -1211
rect 387 -1212 388 -1194
rect 422 -1212 423 -1194
rect 516 -1212 517 -1194
rect 530 -1317 531 -1211
rect 1136 -1317 1137 -1211
rect 1206 -1212 1207 -1194
rect 1444 -1317 1445 -1211
rect 1521 -1317 1522 -1211
rect 1570 -1212 1571 -1194
rect 142 -1214 143 -1194
rect 149 -1317 150 -1213
rect 163 -1214 164 -1194
rect 1297 -1214 1298 -1194
rect 1325 -1317 1326 -1213
rect 1395 -1214 1396 -1194
rect 1416 -1317 1417 -1213
rect 1479 -1214 1480 -1194
rect 142 -1317 143 -1215
rect 1122 -1216 1123 -1194
rect 1129 -1216 1130 -1194
rect 1206 -1317 1207 -1215
rect 1241 -1216 1242 -1194
rect 1297 -1317 1298 -1215
rect 1339 -1216 1340 -1194
rect 1402 -1317 1403 -1215
rect 1409 -1216 1410 -1194
rect 1479 -1317 1480 -1215
rect 124 -1317 125 -1217
rect 1409 -1317 1410 -1217
rect 1437 -1218 1438 -1194
rect 1654 -1317 1655 -1217
rect 163 -1317 164 -1219
rect 1192 -1220 1193 -1194
rect 1213 -1220 1214 -1194
rect 1241 -1317 1242 -1219
rect 1290 -1220 1291 -1194
rect 1437 -1317 1438 -1219
rect 166 -1222 167 -1194
rect 485 -1317 486 -1221
rect 492 -1222 493 -1194
rect 779 -1317 780 -1221
rect 814 -1317 815 -1221
rect 1640 -1222 1641 -1194
rect 166 -1317 167 -1223
rect 464 -1224 465 -1194
rect 492 -1317 493 -1223
rect 639 -1224 640 -1194
rect 674 -1224 675 -1194
rect 716 -1317 717 -1223
rect 768 -1317 769 -1223
rect 1696 -1317 1697 -1223
rect 184 -1226 185 -1194
rect 688 -1226 689 -1194
rect 695 -1317 696 -1225
rect 978 -1317 979 -1225
rect 982 -1226 983 -1194
rect 999 -1226 1000 -1194
rect 1013 -1317 1014 -1225
rect 1367 -1226 1368 -1194
rect 1374 -1226 1375 -1194
rect 1640 -1317 1641 -1225
rect 82 -1228 83 -1194
rect 184 -1317 185 -1227
rect 198 -1228 199 -1194
rect 467 -1228 468 -1194
rect 513 -1317 514 -1227
rect 1500 -1317 1501 -1227
rect 198 -1317 199 -1229
rect 625 -1230 626 -1194
rect 639 -1317 640 -1229
rect 653 -1230 654 -1194
rect 709 -1317 710 -1229
rect 719 -1230 720 -1194
rect 772 -1230 773 -1194
rect 835 -1317 836 -1229
rect 894 -1230 895 -1194
rect 912 -1230 913 -1194
rect 936 -1317 937 -1229
rect 1626 -1230 1627 -1194
rect 156 -1232 157 -1194
rect 625 -1317 626 -1231
rect 646 -1232 647 -1194
rect 674 -1317 675 -1231
rect 828 -1232 829 -1194
rect 1514 -1317 1515 -1231
rect 1535 -1232 1536 -1194
rect 1626 -1317 1627 -1231
rect 156 -1317 157 -1233
rect 618 -1234 619 -1194
rect 646 -1317 647 -1233
rect 663 -1234 664 -1194
rect 831 -1234 832 -1194
rect 940 -1234 941 -1194
rect 957 -1234 958 -1194
rect 1577 -1234 1578 -1194
rect 233 -1236 234 -1194
rect 331 -1236 332 -1194
rect 352 -1317 353 -1235
rect 450 -1236 451 -1194
rect 478 -1236 479 -1194
rect 772 -1317 773 -1235
rect 884 -1236 885 -1194
rect 940 -1317 941 -1235
rect 971 -1236 972 -1194
rect 1584 -1236 1585 -1194
rect 212 -1238 213 -1194
rect 331 -1317 332 -1237
rect 387 -1317 388 -1237
rect 499 -1238 500 -1194
rect 576 -1317 577 -1237
rect 1528 -1317 1529 -1237
rect 191 -1240 192 -1194
rect 212 -1317 213 -1239
rect 233 -1317 234 -1239
rect 499 -1317 500 -1239
rect 597 -1240 598 -1194
rect 1577 -1317 1578 -1239
rect 177 -1242 178 -1194
rect 191 -1317 192 -1241
rect 236 -1242 237 -1194
rect 1451 -1317 1452 -1241
rect 1472 -1242 1473 -1194
rect 1535 -1317 1536 -1241
rect 177 -1317 178 -1243
rect 219 -1244 220 -1194
rect 240 -1244 241 -1194
rect 618 -1317 619 -1243
rect 653 -1317 654 -1243
rect 950 -1317 951 -1243
rect 975 -1244 976 -1194
rect 1192 -1317 1193 -1243
rect 1276 -1244 1277 -1194
rect 1290 -1317 1291 -1243
rect 1356 -1317 1357 -1243
rect 1584 -1317 1585 -1243
rect 219 -1317 220 -1245
rect 817 -1317 818 -1245
rect 821 -1246 822 -1194
rect 884 -1317 885 -1245
rect 898 -1317 899 -1245
rect 905 -1246 906 -1194
rect 975 -1317 976 -1245
rect 992 -1246 993 -1194
rect 1045 -1246 1046 -1194
rect 1556 -1246 1557 -1194
rect 152 -1248 153 -1194
rect 905 -1317 906 -1247
rect 982 -1317 983 -1247
rect 1262 -1248 1263 -1194
rect 1381 -1248 1382 -1194
rect 1570 -1317 1571 -1247
rect 240 -1317 241 -1249
rect 621 -1250 622 -1194
rect 821 -1317 822 -1249
rect 1010 -1250 1011 -1194
rect 1031 -1250 1032 -1194
rect 1262 -1317 1263 -1249
rect 1395 -1317 1396 -1249
rect 1734 -1317 1735 -1249
rect 254 -1317 255 -1251
rect 345 -1252 346 -1194
rect 394 -1252 395 -1194
rect 464 -1317 465 -1251
rect 478 -1317 479 -1251
rect 527 -1252 528 -1194
rect 544 -1252 545 -1194
rect 1381 -1317 1382 -1251
rect 1423 -1252 1424 -1194
rect 1472 -1317 1473 -1251
rect 1556 -1317 1557 -1251
rect 1647 -1252 1648 -1194
rect 37 -1254 38 -1194
rect 527 -1317 528 -1253
rect 562 -1254 563 -1194
rect 597 -1317 598 -1253
rect 611 -1254 612 -1194
rect 691 -1317 692 -1253
rect 989 -1254 990 -1194
rect 1059 -1254 1060 -1194
rect 1080 -1254 1081 -1194
rect 1367 -1317 1368 -1253
rect 1388 -1254 1389 -1194
rect 1423 -1317 1424 -1253
rect 1612 -1254 1613 -1194
rect 1647 -1317 1648 -1253
rect 37 -1317 38 -1255
rect 548 -1256 549 -1194
rect 614 -1256 615 -1194
rect 1591 -1317 1592 -1255
rect 278 -1258 279 -1194
rect 807 -1258 808 -1194
rect 989 -1317 990 -1257
rect 1087 -1258 1088 -1194
rect 1108 -1258 1109 -1194
rect 1339 -1317 1340 -1257
rect 1549 -1258 1550 -1194
rect 1612 -1317 1613 -1257
rect 296 -1260 297 -1194
rect 296 -1317 297 -1259
rect 296 -1260 297 -1194
rect 296 -1317 297 -1259
rect 310 -1260 311 -1194
rect 509 -1260 510 -1194
rect 548 -1317 549 -1259
rect 555 -1260 556 -1194
rect 751 -1260 752 -1194
rect 1388 -1317 1389 -1259
rect 1493 -1260 1494 -1194
rect 1549 -1317 1550 -1259
rect 310 -1317 311 -1261
rect 460 -1317 461 -1261
rect 471 -1262 472 -1194
rect 562 -1317 563 -1261
rect 751 -1317 752 -1261
rect 758 -1262 759 -1194
rect 807 -1317 808 -1261
rect 1115 -1317 1116 -1261
rect 1129 -1317 1130 -1261
rect 1227 -1262 1228 -1194
rect 1255 -1262 1256 -1194
rect 1493 -1317 1494 -1261
rect 317 -1264 318 -1194
rect 726 -1264 727 -1194
rect 1003 -1264 1004 -1194
rect 1059 -1317 1060 -1263
rect 1108 -1317 1109 -1263
rect 1353 -1264 1354 -1194
rect 282 -1266 283 -1194
rect 317 -1317 318 -1265
rect 324 -1266 325 -1194
rect 359 -1317 360 -1265
rect 394 -1317 395 -1265
rect 870 -1266 871 -1194
rect 1003 -1317 1004 -1265
rect 1234 -1266 1235 -1194
rect 1353 -1317 1354 -1265
rect 1374 -1317 1375 -1265
rect 170 -1268 171 -1194
rect 324 -1317 325 -1267
rect 345 -1317 346 -1267
rect 408 -1268 409 -1194
rect 429 -1268 430 -1194
rect 516 -1317 517 -1267
rect 555 -1317 556 -1267
rect 831 -1317 832 -1267
rect 870 -1317 871 -1267
rect 1017 -1268 1018 -1194
rect 1024 -1268 1025 -1194
rect 1087 -1317 1088 -1267
rect 1143 -1268 1144 -1194
rect 1213 -1317 1214 -1267
rect 1220 -1268 1221 -1194
rect 1276 -1317 1277 -1267
rect 170 -1317 171 -1269
rect 604 -1270 605 -1194
rect 877 -1270 878 -1194
rect 1220 -1317 1221 -1269
rect 282 -1317 283 -1271
rect 985 -1317 986 -1271
rect 996 -1272 997 -1194
rect 1024 -1317 1025 -1271
rect 1045 -1317 1046 -1271
rect 1164 -1272 1165 -1194
rect 1171 -1272 1172 -1194
rect 1255 -1317 1256 -1271
rect 338 -1274 339 -1194
rect 429 -1317 430 -1273
rect 443 -1274 444 -1194
rect 446 -1290 447 -1273
rect 450 -1317 451 -1273
rect 583 -1274 584 -1194
rect 590 -1274 591 -1194
rect 877 -1317 878 -1273
rect 933 -1274 934 -1194
rect 996 -1317 997 -1273
rect 1010 -1317 1011 -1273
rect 1080 -1317 1081 -1273
rect 1094 -1274 1095 -1194
rect 1171 -1317 1172 -1273
rect 1199 -1274 1200 -1194
rect 1227 -1317 1228 -1273
rect 86 -1276 87 -1194
rect 583 -1317 584 -1275
rect 933 -1317 934 -1275
rect 1066 -1276 1067 -1194
rect 1094 -1317 1095 -1275
rect 1157 -1276 1158 -1194
rect 1164 -1317 1165 -1275
rect 1178 -1276 1179 -1194
rect 261 -1278 262 -1194
rect 338 -1317 339 -1277
rect 408 -1317 409 -1277
rect 415 -1278 416 -1194
rect 443 -1317 444 -1277
rect 534 -1278 535 -1194
rect 604 -1317 605 -1277
rect 947 -1278 948 -1194
rect 1017 -1317 1018 -1277
rect 1048 -1278 1049 -1194
rect 1430 -1278 1431 -1194
rect 44 -1280 45 -1194
rect 534 -1317 535 -1279
rect 569 -1280 570 -1194
rect 758 -1317 759 -1279
rect 947 -1317 948 -1279
rect 1713 -1317 1714 -1279
rect 44 -1317 45 -1281
rect 75 -1282 76 -1194
rect 226 -1282 227 -1194
rect 569 -1317 570 -1281
rect 954 -1282 955 -1194
rect 1234 -1317 1235 -1281
rect 1360 -1282 1361 -1194
rect 1430 -1317 1431 -1281
rect 75 -1317 76 -1283
rect 86 -1317 87 -1283
rect 226 -1317 227 -1283
rect 457 -1284 458 -1194
rect 471 -1317 472 -1283
rect 747 -1284 748 -1194
rect 863 -1284 864 -1194
rect 954 -1317 955 -1283
rect 961 -1284 962 -1194
rect 1066 -1317 1067 -1283
rect 1101 -1284 1102 -1194
rect 1143 -1317 1144 -1283
rect 1150 -1284 1151 -1194
rect 1199 -1317 1200 -1283
rect 1304 -1284 1305 -1194
rect 1360 -1317 1361 -1283
rect 261 -1317 262 -1285
rect 422 -1317 423 -1285
rect 425 -1317 426 -1285
rect 1304 -1317 1305 -1285
rect 415 -1317 416 -1287
rect 681 -1288 682 -1194
rect 702 -1288 703 -1194
rect 961 -1317 962 -1287
rect 968 -1288 969 -1194
rect 1178 -1317 1179 -1287
rect 366 -1290 367 -1194
rect 681 -1317 682 -1289
rect 800 -1290 801 -1194
rect 863 -1317 864 -1289
rect 919 -1290 920 -1194
rect 968 -1317 969 -1289
rect 999 -1317 1000 -1289
rect 1031 -1317 1032 -1289
rect 1038 -1290 1039 -1194
rect 1150 -1317 1151 -1289
rect 1157 -1317 1158 -1289
rect 1283 -1290 1284 -1194
rect 128 -1292 129 -1194
rect 800 -1317 801 -1291
rect 842 -1292 843 -1194
rect 1101 -1317 1102 -1291
rect 107 -1294 108 -1194
rect 128 -1317 129 -1293
rect 303 -1294 304 -1194
rect 366 -1317 367 -1293
rect 509 -1317 510 -1293
rect 667 -1294 668 -1194
rect 842 -1317 843 -1293
rect 856 -1294 857 -1194
rect 1052 -1294 1053 -1194
rect 1122 -1317 1123 -1293
rect 107 -1317 108 -1295
rect 268 -1296 269 -1194
rect 303 -1317 304 -1295
rect 401 -1296 402 -1194
rect 628 -1317 629 -1295
rect 667 -1317 668 -1295
rect 828 -1317 829 -1295
rect 856 -1317 857 -1295
rect 1052 -1317 1053 -1295
rect 1563 -1296 1564 -1194
rect 114 -1298 115 -1194
rect 401 -1317 402 -1297
rect 632 -1298 633 -1194
rect 702 -1317 703 -1297
rect 849 -1298 850 -1194
rect 919 -1317 920 -1297
rect 1055 -1317 1056 -1297
rect 1311 -1298 1312 -1194
rect 1507 -1298 1508 -1194
rect 1563 -1317 1564 -1297
rect 114 -1317 115 -1299
rect 688 -1317 689 -1299
rect 765 -1300 766 -1194
rect 849 -1317 850 -1299
rect 1073 -1300 1074 -1194
rect 1283 -1317 1284 -1299
rect 1311 -1317 1312 -1299
rect 1346 -1300 1347 -1194
rect 1458 -1300 1459 -1194
rect 1507 -1317 1508 -1299
rect 268 -1317 269 -1301
rect 289 -1302 290 -1194
rect 373 -1302 374 -1194
rect 632 -1317 633 -1301
rect 660 -1302 661 -1194
rect 1038 -1317 1039 -1301
rect 1458 -1317 1459 -1301
rect 1664 -1302 1665 -1194
rect 51 -1304 52 -1194
rect 289 -1317 290 -1303
rect 373 -1317 374 -1303
rect 436 -1304 437 -1194
rect 660 -1317 661 -1303
rect 737 -1304 738 -1194
rect 765 -1317 766 -1303
rect 912 -1317 913 -1303
rect 51 -1317 52 -1305
rect 614 -1317 615 -1305
rect 730 -1306 731 -1194
rect 737 -1317 738 -1305
rect 786 -1306 787 -1194
rect 1073 -1317 1074 -1305
rect 257 -1308 258 -1194
rect 436 -1317 437 -1307
rect 481 -1317 482 -1307
rect 730 -1317 731 -1307
rect 786 -1317 787 -1307
rect 1248 -1308 1249 -1194
rect 891 -1310 892 -1194
rect 1346 -1317 1347 -1309
rect 891 -1317 892 -1311
rect 926 -1312 927 -1194
rect 1248 -1317 1249 -1311
rect 1332 -1312 1333 -1194
rect 82 -1317 83 -1313
rect 926 -1317 927 -1313
rect 1269 -1314 1270 -1194
rect 1332 -1317 1333 -1313
rect 93 -1317 94 -1315
rect 1269 -1317 1270 -1315
rect 16 -1472 17 -1326
rect 51 -1327 52 -1325
rect 58 -1327 59 -1325
rect 422 -1327 423 -1325
rect 478 -1327 479 -1325
rect 1374 -1327 1375 -1325
rect 1493 -1327 1494 -1325
rect 1731 -1327 1732 -1325
rect 1738 -1327 1739 -1325
rect 1745 -1472 1746 -1326
rect 37 -1329 38 -1325
rect 422 -1472 423 -1328
rect 478 -1472 479 -1328
rect 520 -1329 521 -1325
rect 579 -1329 580 -1325
rect 1276 -1329 1277 -1325
rect 1346 -1329 1347 -1325
rect 1706 -1329 1707 -1325
rect 1717 -1329 1718 -1325
rect 1734 -1329 1735 -1325
rect 37 -1472 38 -1330
rect 229 -1472 230 -1330
rect 233 -1472 234 -1330
rect 282 -1331 283 -1325
rect 289 -1331 290 -1325
rect 527 -1331 528 -1325
rect 597 -1331 598 -1325
rect 765 -1331 766 -1325
rect 768 -1331 769 -1325
rect 1171 -1331 1172 -1325
rect 1269 -1331 1270 -1325
rect 1269 -1472 1270 -1330
rect 1269 -1331 1270 -1325
rect 1269 -1472 1270 -1330
rect 1276 -1472 1277 -1330
rect 1360 -1331 1361 -1325
rect 1493 -1472 1494 -1330
rect 1521 -1331 1522 -1325
rect 1556 -1331 1557 -1325
rect 1556 -1472 1557 -1330
rect 1556 -1331 1557 -1325
rect 1556 -1472 1557 -1330
rect 1626 -1331 1627 -1325
rect 1720 -1472 1721 -1330
rect 44 -1333 45 -1325
rect 72 -1333 73 -1325
rect 82 -1333 83 -1325
rect 1297 -1333 1298 -1325
rect 1521 -1472 1522 -1332
rect 1591 -1333 1592 -1325
rect 1668 -1333 1669 -1325
rect 1668 -1472 1669 -1332
rect 1668 -1333 1669 -1325
rect 1668 -1472 1669 -1332
rect 1675 -1333 1676 -1325
rect 1703 -1472 1704 -1332
rect 44 -1472 45 -1334
rect 198 -1335 199 -1325
rect 212 -1335 213 -1325
rect 212 -1472 213 -1334
rect 212 -1335 213 -1325
rect 212 -1472 213 -1334
rect 240 -1335 241 -1325
rect 831 -1335 832 -1325
rect 873 -1472 874 -1334
rect 1423 -1335 1424 -1325
rect 1584 -1335 1585 -1325
rect 1626 -1472 1627 -1334
rect 1682 -1335 1683 -1325
rect 1717 -1472 1718 -1334
rect 51 -1472 52 -1336
rect 625 -1337 626 -1325
rect 628 -1337 629 -1325
rect 779 -1337 780 -1325
rect 786 -1337 787 -1325
rect 842 -1337 843 -1325
rect 901 -1472 902 -1336
rect 1094 -1337 1095 -1325
rect 1125 -1472 1126 -1336
rect 1591 -1472 1592 -1336
rect 1696 -1337 1697 -1325
rect 1710 -1472 1711 -1336
rect 75 -1472 76 -1338
rect 240 -1472 241 -1338
rect 250 -1339 251 -1325
rect 1304 -1339 1305 -1325
rect 1699 -1472 1700 -1338
rect 1724 -1339 1725 -1325
rect 82 -1472 83 -1340
rect 1339 -1341 1340 -1325
rect 86 -1343 87 -1325
rect 96 -1343 97 -1325
rect 100 -1343 101 -1325
rect 100 -1472 101 -1342
rect 100 -1343 101 -1325
rect 100 -1472 101 -1342
rect 124 -1343 125 -1325
rect 149 -1343 150 -1325
rect 170 -1343 171 -1325
rect 733 -1472 734 -1342
rect 765 -1472 766 -1342
rect 1374 -1472 1375 -1342
rect 93 -1345 94 -1325
rect 1262 -1345 1263 -1325
rect 1283 -1345 1284 -1325
rect 1675 -1472 1676 -1344
rect 96 -1472 97 -1346
rect 324 -1347 325 -1325
rect 366 -1347 367 -1325
rect 576 -1347 577 -1325
rect 590 -1347 591 -1325
rect 625 -1472 626 -1346
rect 632 -1347 633 -1325
rect 786 -1472 787 -1346
rect 796 -1347 797 -1325
rect 1360 -1472 1361 -1346
rect 107 -1349 108 -1325
rect 170 -1472 171 -1348
rect 177 -1349 178 -1325
rect 236 -1349 237 -1325
rect 264 -1472 265 -1348
rect 317 -1349 318 -1325
rect 324 -1472 325 -1348
rect 541 -1349 542 -1325
rect 548 -1349 549 -1325
rect 576 -1472 577 -1348
rect 597 -1472 598 -1348
rect 1101 -1349 1102 -1325
rect 1136 -1349 1137 -1325
rect 1724 -1472 1725 -1348
rect 107 -1472 108 -1350
rect 1507 -1351 1508 -1325
rect 135 -1353 136 -1325
rect 457 -1353 458 -1325
rect 460 -1353 461 -1325
rect 1346 -1472 1347 -1352
rect 135 -1472 136 -1354
rect 502 -1472 503 -1354
rect 506 -1355 507 -1325
rect 632 -1472 633 -1354
rect 653 -1355 654 -1325
rect 817 -1355 818 -1325
rect 821 -1355 822 -1325
rect 1192 -1355 1193 -1325
rect 1262 -1472 1263 -1354
rect 1318 -1355 1319 -1325
rect 1339 -1472 1340 -1354
rect 1549 -1355 1550 -1325
rect 142 -1357 143 -1325
rect 807 -1472 808 -1356
rect 828 -1357 829 -1325
rect 1640 -1357 1641 -1325
rect 30 -1359 31 -1325
rect 142 -1472 143 -1358
rect 149 -1472 150 -1358
rect 562 -1359 563 -1325
rect 593 -1472 594 -1358
rect 1640 -1472 1641 -1358
rect 26 -1472 27 -1360
rect 30 -1472 31 -1360
rect 177 -1472 178 -1360
rect 184 -1361 185 -1325
rect 191 -1361 192 -1325
rect 198 -1472 199 -1360
rect 219 -1361 220 -1325
rect 506 -1472 507 -1360
rect 520 -1472 521 -1360
rect 891 -1361 892 -1325
rect 947 -1361 948 -1325
rect 1542 -1361 1543 -1325
rect 117 -1472 118 -1362
rect 1542 -1472 1543 -1362
rect 163 -1365 164 -1325
rect 184 -1472 185 -1364
rect 219 -1472 220 -1364
rect 254 -1365 255 -1325
rect 268 -1365 269 -1325
rect 268 -1472 269 -1364
rect 268 -1365 269 -1325
rect 268 -1472 269 -1364
rect 275 -1365 276 -1325
rect 450 -1365 451 -1325
rect 457 -1472 458 -1364
rect 730 -1365 731 -1325
rect 779 -1472 780 -1364
rect 835 -1365 836 -1325
rect 891 -1472 892 -1364
rect 989 -1365 990 -1325
rect 1010 -1365 1011 -1325
rect 1213 -1365 1214 -1325
rect 1297 -1472 1298 -1364
rect 1311 -1365 1312 -1325
rect 114 -1367 115 -1325
rect 254 -1472 255 -1366
rect 275 -1472 276 -1366
rect 331 -1367 332 -1325
rect 366 -1472 367 -1366
rect 691 -1367 692 -1325
rect 695 -1367 696 -1325
rect 894 -1472 895 -1366
rect 947 -1472 948 -1366
rect 968 -1367 969 -1325
rect 978 -1367 979 -1325
rect 1612 -1367 1613 -1325
rect 156 -1369 157 -1325
rect 163 -1472 164 -1368
rect 247 -1369 248 -1325
rect 1318 -1472 1319 -1368
rect 1612 -1472 1613 -1368
rect 1633 -1369 1634 -1325
rect 156 -1472 157 -1370
rect 191 -1472 192 -1370
rect 247 -1472 248 -1370
rect 278 -1371 279 -1325
rect 282 -1472 283 -1370
rect 345 -1371 346 -1325
rect 373 -1371 374 -1325
rect 1507 -1472 1508 -1370
rect 1605 -1371 1606 -1325
rect 1633 -1472 1634 -1370
rect 289 -1472 290 -1372
rect 418 -1472 419 -1372
rect 436 -1373 437 -1325
rect 541 -1472 542 -1372
rect 548 -1472 549 -1372
rect 555 -1373 556 -1325
rect 562 -1472 563 -1372
rect 604 -1373 605 -1325
rect 614 -1373 615 -1325
rect 821 -1472 822 -1372
rect 828 -1472 829 -1372
rect 863 -1373 864 -1325
rect 968 -1472 969 -1372
rect 1024 -1373 1025 -1325
rect 1027 -1472 1028 -1372
rect 1584 -1472 1585 -1372
rect 296 -1375 297 -1325
rect 611 -1375 612 -1325
rect 618 -1375 619 -1325
rect 663 -1375 664 -1325
rect 667 -1375 668 -1325
rect 989 -1472 990 -1374
rect 1045 -1375 1046 -1325
rect 1048 -1415 1049 -1374
rect 1055 -1375 1056 -1325
rect 1332 -1375 1333 -1325
rect 1416 -1375 1417 -1325
rect 1605 -1472 1606 -1374
rect 303 -1377 304 -1325
rect 345 -1472 346 -1376
rect 352 -1377 353 -1325
rect 614 -1472 615 -1376
rect 639 -1377 640 -1325
rect 667 -1472 668 -1376
rect 688 -1377 689 -1325
rect 1479 -1377 1480 -1325
rect 317 -1472 318 -1378
rect 789 -1379 790 -1325
rect 835 -1472 836 -1378
rect 936 -1379 937 -1325
rect 982 -1379 983 -1325
rect 1416 -1472 1417 -1378
rect 1479 -1472 1480 -1378
rect 1514 -1379 1515 -1325
rect 331 -1472 332 -1380
rect 499 -1381 500 -1325
rect 590 -1472 591 -1380
rect 1514 -1472 1515 -1380
rect 352 -1472 353 -1382
rect 408 -1383 409 -1325
rect 415 -1383 416 -1325
rect 436 -1472 437 -1382
rect 450 -1472 451 -1382
rect 772 -1383 773 -1325
rect 863 -1472 864 -1382
rect 1108 -1383 1109 -1325
rect 1129 -1383 1130 -1325
rect 1192 -1472 1193 -1382
rect 1213 -1472 1214 -1382
rect 1255 -1383 1256 -1325
rect 1304 -1472 1305 -1382
rect 1409 -1383 1410 -1325
rect 338 -1385 339 -1325
rect 408 -1472 409 -1384
rect 415 -1472 416 -1384
rect 534 -1385 535 -1325
rect 604 -1472 605 -1384
rect 635 -1472 636 -1384
rect 639 -1472 640 -1384
rect 1073 -1385 1074 -1325
rect 1094 -1472 1095 -1384
rect 1206 -1385 1207 -1325
rect 1255 -1472 1256 -1384
rect 1402 -1385 1403 -1325
rect 261 -1387 262 -1325
rect 338 -1472 339 -1386
rect 373 -1472 374 -1386
rect 583 -1387 584 -1325
rect 611 -1472 612 -1386
rect 1423 -1472 1424 -1386
rect 261 -1472 262 -1388
rect 1101 -1472 1102 -1388
rect 1146 -1472 1147 -1388
rect 1654 -1389 1655 -1325
rect 387 -1391 388 -1325
rect 527 -1472 528 -1390
rect 534 -1472 535 -1390
rect 856 -1391 857 -1325
rect 877 -1391 878 -1325
rect 936 -1472 937 -1390
rect 940 -1391 941 -1325
rect 982 -1472 983 -1390
rect 985 -1391 986 -1325
rect 1689 -1391 1690 -1325
rect 303 -1472 304 -1392
rect 387 -1472 388 -1392
rect 394 -1393 395 -1325
rect 1010 -1472 1011 -1392
rect 1017 -1393 1018 -1325
rect 1108 -1472 1109 -1392
rect 1171 -1472 1172 -1392
rect 1241 -1393 1242 -1325
rect 1311 -1472 1312 -1392
rect 1444 -1393 1445 -1325
rect 1654 -1472 1655 -1392
rect 1661 -1393 1662 -1325
rect 205 -1395 206 -1325
rect 394 -1472 395 -1394
rect 401 -1395 402 -1325
rect 842 -1472 843 -1394
rect 877 -1472 878 -1394
rect 898 -1395 899 -1325
rect 905 -1395 906 -1325
rect 1073 -1472 1074 -1394
rect 1139 -1472 1140 -1394
rect 1241 -1472 1242 -1394
rect 1325 -1395 1326 -1325
rect 1409 -1472 1410 -1394
rect 79 -1472 80 -1396
rect 898 -1472 899 -1396
rect 940 -1472 941 -1396
rect 961 -1397 962 -1325
rect 1017 -1472 1018 -1396
rect 1066 -1397 1067 -1325
rect 1069 -1472 1070 -1396
rect 1647 -1397 1648 -1325
rect 110 -1472 111 -1398
rect 205 -1472 206 -1398
rect 401 -1472 402 -1398
rect 443 -1399 444 -1325
rect 464 -1399 465 -1325
rect 618 -1472 619 -1398
rect 653 -1472 654 -1398
rect 709 -1399 710 -1325
rect 719 -1472 720 -1398
rect 954 -1399 955 -1325
rect 1045 -1472 1046 -1398
rect 1087 -1399 1088 -1325
rect 1185 -1399 1186 -1325
rect 1283 -1472 1284 -1398
rect 1332 -1472 1333 -1398
rect 1388 -1399 1389 -1325
rect 1402 -1472 1403 -1398
rect 1458 -1399 1459 -1325
rect 1619 -1399 1620 -1325
rect 1647 -1472 1648 -1398
rect 121 -1401 122 -1325
rect 1388 -1472 1389 -1400
rect 1458 -1472 1459 -1400
rect 1486 -1401 1487 -1325
rect 121 -1472 122 -1402
rect 380 -1403 381 -1325
rect 464 -1472 465 -1402
rect 646 -1403 647 -1325
rect 660 -1403 661 -1325
rect 1220 -1403 1221 -1325
rect 1353 -1403 1354 -1325
rect 1661 -1472 1662 -1402
rect 128 -1405 129 -1325
rect 646 -1472 647 -1404
rect 660 -1472 661 -1404
rect 975 -1405 976 -1325
rect 1087 -1472 1088 -1404
rect 1150 -1405 1151 -1325
rect 1185 -1472 1186 -1404
rect 1381 -1405 1382 -1325
rect 1486 -1472 1487 -1404
rect 1528 -1405 1529 -1325
rect 128 -1472 129 -1406
rect 359 -1407 360 -1325
rect 380 -1472 381 -1406
rect 429 -1407 430 -1325
rect 485 -1407 486 -1325
rect 726 -1472 727 -1406
rect 730 -1472 731 -1406
rect 1549 -1472 1550 -1406
rect 23 -1409 24 -1325
rect 485 -1472 486 -1408
rect 499 -1472 500 -1408
rect 1619 -1472 1620 -1408
rect 65 -1411 66 -1325
rect 429 -1472 430 -1410
rect 513 -1472 514 -1410
rect 1066 -1472 1067 -1410
rect 1206 -1472 1207 -1410
rect 1290 -1411 1291 -1325
rect 1353 -1472 1354 -1410
rect 1437 -1411 1438 -1325
rect 1528 -1472 1529 -1410
rect 1570 -1411 1571 -1325
rect 65 -1472 66 -1412
rect 222 -1472 223 -1412
rect 226 -1413 227 -1325
rect 443 -1472 444 -1412
rect 555 -1472 556 -1412
rect 1689 -1472 1690 -1412
rect 310 -1415 311 -1325
rect 359 -1472 360 -1414
rect 583 -1472 584 -1414
rect 1013 -1415 1014 -1325
rect 1150 -1472 1151 -1414
rect 1157 -1415 1158 -1325
rect 1290 -1472 1291 -1414
rect 310 -1472 311 -1416
rect 471 -1417 472 -1325
rect 677 -1472 678 -1416
rect 1220 -1472 1221 -1416
rect 1248 -1417 1249 -1325
rect 1381 -1472 1382 -1416
rect 58 -1472 59 -1418
rect 471 -1472 472 -1418
rect 688 -1472 689 -1418
rect 702 -1419 703 -1325
rect 709 -1472 710 -1418
rect 716 -1419 717 -1325
rect 723 -1419 724 -1325
rect 793 -1419 794 -1325
rect 800 -1419 801 -1325
rect 1129 -1472 1130 -1418
rect 1248 -1472 1249 -1418
rect 1395 -1419 1396 -1325
rect 695 -1472 696 -1420
rect 758 -1421 759 -1325
rect 800 -1472 801 -1420
rect 849 -1421 850 -1325
rect 866 -1472 867 -1420
rect 1570 -1472 1571 -1420
rect 702 -1472 703 -1422
rect 1031 -1423 1032 -1325
rect 1395 -1472 1396 -1422
rect 1451 -1423 1452 -1325
rect 61 -1472 62 -1424
rect 1031 -1472 1032 -1424
rect 1430 -1425 1431 -1325
rect 1451 -1472 1452 -1424
rect 716 -1472 717 -1426
rect 1157 -1472 1158 -1426
rect 1430 -1472 1431 -1426
rect 1465 -1427 1466 -1325
rect 226 -1472 227 -1428
rect 1465 -1472 1466 -1428
rect 723 -1472 724 -1430
rect 1367 -1431 1368 -1325
rect 744 -1433 745 -1325
rect 793 -1472 794 -1432
rect 814 -1433 815 -1325
rect 905 -1472 906 -1432
rect 919 -1433 920 -1325
rect 961 -1472 962 -1432
rect 975 -1472 976 -1432
rect 996 -1433 997 -1325
rect 1367 -1472 1368 -1432
rect 1472 -1433 1473 -1325
rect 737 -1435 738 -1325
rect 744 -1472 745 -1434
rect 751 -1435 752 -1325
rect 772 -1472 773 -1434
rect 814 -1472 815 -1434
rect 884 -1435 885 -1325
rect 919 -1472 920 -1434
rect 1059 -1435 1060 -1325
rect 1472 -1472 1473 -1434
rect 1500 -1435 1501 -1325
rect 145 -1437 146 -1325
rect 751 -1472 752 -1436
rect 758 -1472 759 -1436
rect 870 -1437 871 -1325
rect 933 -1437 934 -1325
rect 1437 -1472 1438 -1436
rect 1500 -1472 1501 -1436
rect 1535 -1437 1536 -1325
rect 569 -1439 570 -1325
rect 737 -1472 738 -1438
rect 824 -1439 825 -1325
rect 1444 -1472 1445 -1438
rect 1535 -1472 1536 -1438
rect 1577 -1439 1578 -1325
rect 509 -1441 510 -1325
rect 569 -1472 570 -1440
rect 681 -1441 682 -1325
rect 884 -1472 885 -1440
rect 933 -1472 934 -1440
rect 1682 -1472 1683 -1440
rect 674 -1443 675 -1325
rect 681 -1472 682 -1442
rect 849 -1472 850 -1442
rect 926 -1443 927 -1325
rect 954 -1472 955 -1442
rect 1143 -1443 1144 -1325
rect 1577 -1472 1578 -1442
rect 1598 -1443 1599 -1325
rect 492 -1445 493 -1325
rect 674 -1472 675 -1444
rect 856 -1472 857 -1444
rect 870 -1472 871 -1444
rect 926 -1472 927 -1444
rect 1003 -1445 1004 -1325
rect 1059 -1472 1060 -1444
rect 1122 -1445 1123 -1325
rect 1143 -1472 1144 -1444
rect 1325 -1472 1326 -1444
rect 1563 -1445 1564 -1325
rect 1598 -1472 1599 -1444
rect 86 -1472 87 -1446
rect 1122 -1472 1123 -1446
rect 1227 -1447 1228 -1325
rect 1563 -1472 1564 -1446
rect 93 -1472 94 -1448
rect 492 -1472 493 -1448
rect 530 -1449 531 -1325
rect 1227 -1472 1228 -1448
rect 996 -1472 997 -1450
rect 1038 -1451 1039 -1325
rect 1003 -1472 1004 -1452
rect 1199 -1453 1200 -1325
rect 600 -1472 601 -1454
rect 1199 -1472 1200 -1454
rect 1038 -1472 1039 -1456
rect 1115 -1457 1116 -1325
rect 1115 -1472 1116 -1458
rect 1164 -1459 1165 -1325
rect 1164 -1472 1165 -1460
rect 1234 -1461 1235 -1325
rect 1080 -1463 1081 -1325
rect 1234 -1472 1235 -1462
rect 1080 -1472 1081 -1464
rect 1178 -1465 1179 -1325
rect 1052 -1467 1053 -1325
rect 1178 -1472 1179 -1466
rect 912 -1469 913 -1325
rect 1052 -1472 1053 -1468
rect 642 -1472 643 -1470
rect 912 -1472 913 -1470
rect 16 -1482 17 -1480
rect 765 -1482 766 -1480
rect 786 -1482 787 -1480
rect 863 -1482 864 -1480
rect 870 -1482 871 -1480
rect 919 -1482 920 -1480
rect 1024 -1482 1025 -1480
rect 1094 -1482 1095 -1480
rect 1104 -1609 1105 -1481
rect 1339 -1482 1340 -1480
rect 1745 -1482 1746 -1480
rect 1752 -1609 1753 -1481
rect 23 -1609 24 -1483
rect 75 -1484 76 -1480
rect 96 -1609 97 -1483
rect 1640 -1484 1641 -1480
rect 30 -1486 31 -1480
rect 82 -1486 83 -1480
rect 100 -1486 101 -1480
rect 100 -1609 101 -1485
rect 100 -1486 101 -1480
rect 100 -1609 101 -1485
rect 107 -1486 108 -1480
rect 415 -1486 416 -1480
rect 418 -1486 419 -1480
rect 765 -1609 766 -1485
rect 786 -1609 787 -1485
rect 905 -1486 906 -1480
rect 1024 -1609 1025 -1485
rect 1087 -1486 1088 -1480
rect 1118 -1609 1119 -1485
rect 1710 -1486 1711 -1480
rect 58 -1609 59 -1487
rect 1689 -1488 1690 -1480
rect 61 -1609 62 -1489
rect 117 -1490 118 -1480
rect 142 -1490 143 -1480
rect 208 -1609 209 -1489
rect 226 -1490 227 -1480
rect 359 -1490 360 -1480
rect 373 -1490 374 -1480
rect 761 -1609 762 -1489
rect 863 -1609 864 -1489
rect 940 -1490 941 -1480
rect 1073 -1490 1074 -1480
rect 1713 -1609 1714 -1489
rect 68 -1609 69 -1491
rect 548 -1492 549 -1480
rect 555 -1492 556 -1480
rect 611 -1609 612 -1491
rect 621 -1609 622 -1491
rect 709 -1492 710 -1480
rect 719 -1492 720 -1480
rect 1563 -1492 1564 -1480
rect 1640 -1609 1641 -1491
rect 1668 -1492 1669 -1480
rect 72 -1494 73 -1480
rect 366 -1494 367 -1480
rect 390 -1494 391 -1480
rect 429 -1494 430 -1480
rect 443 -1494 444 -1480
rect 544 -1609 545 -1493
rect 562 -1494 563 -1480
rect 709 -1609 710 -1493
rect 733 -1494 734 -1480
rect 919 -1609 920 -1493
rect 1073 -1609 1074 -1493
rect 1143 -1494 1144 -1480
rect 1153 -1609 1154 -1493
rect 1332 -1494 1333 -1480
rect 1339 -1609 1340 -1493
rect 1416 -1494 1417 -1480
rect 1493 -1494 1494 -1480
rect 1689 -1609 1690 -1493
rect 44 -1496 45 -1480
rect 72 -1609 73 -1495
rect 107 -1609 108 -1495
rect 366 -1609 367 -1495
rect 394 -1496 395 -1480
rect 768 -1496 769 -1480
rect 866 -1496 867 -1480
rect 1094 -1609 1095 -1495
rect 1122 -1496 1123 -1480
rect 1262 -1496 1263 -1480
rect 1311 -1496 1312 -1480
rect 1332 -1609 1333 -1495
rect 1416 -1609 1417 -1495
rect 1486 -1496 1487 -1480
rect 1493 -1609 1494 -1495
rect 1535 -1496 1536 -1480
rect 1563 -1609 1564 -1495
rect 1591 -1496 1592 -1480
rect 1612 -1496 1613 -1480
rect 1668 -1609 1669 -1495
rect 44 -1609 45 -1497
rect 369 -1609 370 -1497
rect 394 -1609 395 -1497
rect 471 -1498 472 -1480
rect 474 -1609 475 -1497
rect 961 -1498 962 -1480
rect 989 -1498 990 -1480
rect 1122 -1609 1123 -1497
rect 1125 -1498 1126 -1480
rect 1703 -1498 1704 -1480
rect 30 -1609 31 -1499
rect 471 -1609 472 -1499
rect 492 -1500 493 -1480
rect 901 -1500 902 -1480
rect 905 -1609 906 -1499
rect 926 -1500 927 -1480
rect 961 -1609 962 -1499
rect 968 -1500 969 -1480
rect 975 -1500 976 -1480
rect 989 -1609 990 -1499
rect 1087 -1609 1088 -1499
rect 1171 -1500 1172 -1480
rect 1311 -1609 1312 -1499
rect 1325 -1500 1326 -1480
rect 1486 -1609 1487 -1499
rect 1605 -1500 1606 -1480
rect 114 -1502 115 -1480
rect 436 -1502 437 -1480
rect 443 -1609 444 -1501
rect 1703 -1609 1704 -1501
rect 114 -1609 115 -1503
rect 670 -1609 671 -1503
rect 677 -1504 678 -1480
rect 1549 -1504 1550 -1480
rect 1556 -1504 1557 -1480
rect 1605 -1609 1606 -1503
rect 142 -1609 143 -1505
rect 401 -1506 402 -1480
rect 408 -1506 409 -1480
rect 408 -1609 409 -1505
rect 408 -1506 409 -1480
rect 408 -1609 409 -1505
rect 422 -1506 423 -1480
rect 593 -1506 594 -1480
rect 607 -1609 608 -1505
rect 667 -1506 668 -1480
rect 730 -1506 731 -1480
rect 1262 -1609 1263 -1505
rect 1325 -1609 1326 -1505
rect 1402 -1506 1403 -1480
rect 1500 -1506 1501 -1480
rect 1612 -1609 1613 -1505
rect 51 -1508 52 -1480
rect 401 -1609 402 -1507
rect 436 -1609 437 -1507
rect 929 -1609 930 -1507
rect 975 -1609 976 -1507
rect 1346 -1508 1347 -1480
rect 1402 -1609 1403 -1507
rect 1472 -1508 1473 -1480
rect 1535 -1609 1536 -1507
rect 1577 -1508 1578 -1480
rect 1584 -1508 1585 -1480
rect 1591 -1609 1592 -1507
rect 156 -1510 157 -1480
rect 1556 -1609 1557 -1509
rect 1570 -1510 1571 -1480
rect 1577 -1609 1578 -1509
rect 1584 -1609 1585 -1509
rect 1598 -1510 1599 -1480
rect 156 -1609 157 -1511
rect 212 -1512 213 -1480
rect 226 -1609 227 -1511
rect 257 -1609 258 -1511
rect 261 -1609 262 -1511
rect 282 -1512 283 -1480
rect 296 -1609 297 -1511
rect 618 -1512 619 -1480
rect 632 -1512 633 -1480
rect 1045 -1512 1046 -1480
rect 1048 -1609 1049 -1511
rect 1570 -1609 1571 -1511
rect 1598 -1609 1599 -1511
rect 1619 -1512 1620 -1480
rect 159 -1514 160 -1480
rect 583 -1514 584 -1480
rect 635 -1514 636 -1480
rect 1507 -1514 1508 -1480
rect 1549 -1609 1550 -1513
rect 1720 -1514 1721 -1480
rect 149 -1516 150 -1480
rect 583 -1609 584 -1515
rect 639 -1516 640 -1480
rect 1706 -1609 1707 -1515
rect 149 -1609 150 -1517
rect 558 -1518 559 -1480
rect 562 -1609 563 -1517
rect 681 -1518 682 -1480
rect 712 -1609 713 -1517
rect 1500 -1609 1501 -1517
rect 1619 -1609 1620 -1517
rect 1633 -1518 1634 -1480
rect 191 -1520 192 -1480
rect 219 -1520 220 -1480
rect 229 -1520 230 -1480
rect 982 -1520 983 -1480
rect 1045 -1609 1046 -1519
rect 1129 -1520 1130 -1480
rect 1139 -1520 1140 -1480
rect 1451 -1520 1452 -1480
rect 1472 -1609 1473 -1519
rect 1654 -1520 1655 -1480
rect 194 -1609 195 -1521
rect 534 -1522 535 -1480
rect 541 -1522 542 -1480
rect 555 -1609 556 -1521
rect 576 -1522 577 -1480
rect 597 -1522 598 -1480
rect 604 -1522 605 -1480
rect 681 -1609 682 -1521
rect 730 -1609 731 -1521
rect 779 -1522 780 -1480
rect 796 -1609 797 -1521
rect 1633 -1609 1634 -1521
rect 79 -1524 80 -1480
rect 576 -1609 577 -1523
rect 604 -1609 605 -1523
rect 1682 -1524 1683 -1480
rect 79 -1609 80 -1525
rect 163 -1526 164 -1480
rect 198 -1526 199 -1480
rect 198 -1609 199 -1525
rect 198 -1526 199 -1480
rect 198 -1609 199 -1525
rect 212 -1609 213 -1525
rect 240 -1526 241 -1480
rect 268 -1526 269 -1480
rect 282 -1609 283 -1525
rect 310 -1526 311 -1480
rect 415 -1609 416 -1525
rect 450 -1526 451 -1480
rect 492 -1609 493 -1525
rect 499 -1609 500 -1525
rect 618 -1609 619 -1525
rect 639 -1609 640 -1525
rect 660 -1526 661 -1480
rect 747 -1609 748 -1525
rect 814 -1526 815 -1480
rect 870 -1609 871 -1525
rect 1017 -1526 1018 -1480
rect 1020 -1609 1021 -1525
rect 1654 -1609 1655 -1525
rect 121 -1528 122 -1480
rect 240 -1609 241 -1527
rect 299 -1528 300 -1480
rect 310 -1609 311 -1527
rect 331 -1528 332 -1480
rect 422 -1609 423 -1527
rect 450 -1609 451 -1527
rect 674 -1528 675 -1480
rect 779 -1609 780 -1527
rect 800 -1528 801 -1480
rect 891 -1528 892 -1480
rect 1136 -1609 1137 -1527
rect 1143 -1609 1144 -1527
rect 1206 -1528 1207 -1480
rect 1283 -1528 1284 -1480
rect 1682 -1609 1683 -1527
rect 93 -1530 94 -1480
rect 121 -1609 122 -1529
rect 163 -1609 164 -1529
rect 590 -1530 591 -1480
rect 646 -1530 647 -1480
rect 646 -1609 647 -1529
rect 646 -1530 647 -1480
rect 646 -1609 647 -1529
rect 653 -1530 654 -1480
rect 653 -1609 654 -1529
rect 653 -1530 654 -1480
rect 653 -1609 654 -1529
rect 660 -1609 661 -1529
rect 695 -1530 696 -1480
rect 719 -1609 720 -1529
rect 1283 -1609 1284 -1529
rect 1346 -1609 1347 -1529
rect 1423 -1530 1424 -1480
rect 1451 -1609 1452 -1529
rect 1542 -1530 1543 -1480
rect 93 -1609 94 -1531
rect 625 -1532 626 -1480
rect 674 -1609 675 -1531
rect 737 -1532 738 -1480
rect 793 -1532 794 -1480
rect 814 -1609 815 -1531
rect 891 -1609 892 -1531
rect 996 -1532 997 -1480
rect 1017 -1609 1018 -1531
rect 1675 -1532 1676 -1480
rect 51 -1609 52 -1533
rect 793 -1609 794 -1533
rect 800 -1609 801 -1533
rect 842 -1534 843 -1480
rect 898 -1609 899 -1533
rect 947 -1534 948 -1480
rect 982 -1609 983 -1533
rect 1157 -1534 1158 -1480
rect 1171 -1609 1172 -1533
rect 1234 -1534 1235 -1480
rect 1258 -1609 1259 -1533
rect 1423 -1609 1424 -1533
rect 1521 -1534 1522 -1480
rect 1542 -1609 1543 -1533
rect 1626 -1534 1627 -1480
rect 1675 -1609 1676 -1533
rect 205 -1536 206 -1480
rect 331 -1609 332 -1535
rect 338 -1536 339 -1480
rect 373 -1609 374 -1535
rect 464 -1536 465 -1480
rect 632 -1609 633 -1535
rect 737 -1609 738 -1535
rect 968 -1609 969 -1535
rect 996 -1609 997 -1535
rect 1059 -1536 1060 -1480
rect 1062 -1609 1063 -1535
rect 1157 -1609 1158 -1535
rect 1199 -1536 1200 -1480
rect 1507 -1609 1508 -1535
rect 1521 -1609 1522 -1535
rect 1661 -1536 1662 -1480
rect 191 -1609 192 -1537
rect 1199 -1609 1200 -1537
rect 1206 -1609 1207 -1537
rect 1360 -1538 1361 -1480
rect 1661 -1609 1662 -1537
rect 1710 -1609 1711 -1537
rect 205 -1609 206 -1539
rect 912 -1540 913 -1480
rect 926 -1609 927 -1539
rect 1290 -1540 1291 -1480
rect 219 -1609 220 -1541
rect 247 -1542 248 -1480
rect 303 -1542 304 -1480
rect 464 -1609 465 -1541
rect 502 -1542 503 -1480
rect 688 -1542 689 -1480
rect 758 -1542 759 -1480
rect 912 -1609 913 -1541
rect 933 -1542 934 -1480
rect 1626 -1609 1627 -1541
rect 184 -1544 185 -1480
rect 247 -1609 248 -1543
rect 324 -1544 325 -1480
rect 695 -1609 696 -1543
rect 758 -1609 759 -1543
rect 1185 -1544 1186 -1480
rect 1227 -1544 1228 -1480
rect 1360 -1609 1361 -1543
rect 135 -1546 136 -1480
rect 184 -1609 185 -1545
rect 233 -1546 234 -1480
rect 303 -1609 304 -1545
rect 338 -1609 339 -1545
rect 383 -1609 384 -1545
rect 506 -1546 507 -1480
rect 716 -1546 717 -1480
rect 842 -1609 843 -1545
rect 1066 -1546 1067 -1480
rect 1129 -1609 1130 -1545
rect 1213 -1546 1214 -1480
rect 1227 -1609 1228 -1545
rect 1724 -1546 1725 -1480
rect 37 -1548 38 -1480
rect 135 -1609 136 -1547
rect 233 -1609 234 -1547
rect 387 -1548 388 -1480
rect 457 -1548 458 -1480
rect 506 -1609 507 -1547
rect 513 -1548 514 -1480
rect 513 -1609 514 -1547
rect 513 -1548 514 -1480
rect 513 -1609 514 -1547
rect 520 -1548 521 -1480
rect 1146 -1548 1147 -1480
rect 1185 -1609 1186 -1547
rect 1241 -1548 1242 -1480
rect 1290 -1609 1291 -1547
rect 1297 -1548 1298 -1480
rect 86 -1550 87 -1480
rect 387 -1609 388 -1549
rect 457 -1609 458 -1549
rect 485 -1550 486 -1480
rect 527 -1550 528 -1480
rect 534 -1609 535 -1549
rect 569 -1550 570 -1480
rect 597 -1609 598 -1549
rect 625 -1609 626 -1549
rect 740 -1609 741 -1549
rect 933 -1609 934 -1549
rect 936 -1550 937 -1480
rect 947 -1609 948 -1549
rect 1031 -1550 1032 -1480
rect 1213 -1609 1214 -1549
rect 1353 -1550 1354 -1480
rect 65 -1552 66 -1480
rect 569 -1609 570 -1551
rect 590 -1609 591 -1551
rect 807 -1552 808 -1480
rect 1031 -1609 1032 -1551
rect 1115 -1552 1116 -1480
rect 1234 -1609 1235 -1551
rect 1255 -1552 1256 -1480
rect 1297 -1609 1298 -1551
rect 1395 -1552 1396 -1480
rect 65 -1609 66 -1553
rect 940 -1609 941 -1553
rect 1241 -1609 1242 -1553
rect 1318 -1554 1319 -1480
rect 1353 -1609 1354 -1553
rect 1437 -1554 1438 -1480
rect 86 -1609 87 -1555
rect 835 -1556 836 -1480
rect 873 -1556 874 -1480
rect 1255 -1609 1256 -1555
rect 1318 -1609 1319 -1555
rect 1374 -1556 1375 -1480
rect 1437 -1609 1438 -1555
rect 1528 -1556 1529 -1480
rect 128 -1558 129 -1480
rect 520 -1609 521 -1557
rect 527 -1609 528 -1557
rect 1717 -1558 1718 -1480
rect 128 -1609 129 -1559
rect 275 -1560 276 -1480
rect 345 -1560 346 -1480
rect 429 -1609 430 -1559
rect 485 -1609 486 -1559
rect 751 -1560 752 -1480
rect 807 -1609 808 -1559
rect 1696 -1609 1697 -1559
rect 170 -1562 171 -1480
rect 835 -1609 836 -1561
rect 1115 -1609 1116 -1561
rect 1528 -1609 1529 -1561
rect 170 -1609 171 -1563
rect 352 -1564 353 -1480
rect 359 -1609 360 -1563
rect 478 -1564 479 -1480
rect 667 -1609 668 -1563
rect 1066 -1609 1067 -1563
rect 1367 -1564 1368 -1480
rect 1374 -1609 1375 -1563
rect 254 -1566 255 -1480
rect 324 -1609 325 -1565
rect 352 -1609 353 -1565
rect 380 -1566 381 -1480
rect 478 -1609 479 -1565
rect 828 -1566 829 -1480
rect 1367 -1609 1368 -1565
rect 1444 -1566 1445 -1480
rect 275 -1609 276 -1567
rect 317 -1568 318 -1480
rect 380 -1609 381 -1567
rect 726 -1568 727 -1480
rect 751 -1609 752 -1567
rect 772 -1568 773 -1480
rect 821 -1568 822 -1480
rect 1395 -1609 1396 -1567
rect 1430 -1568 1431 -1480
rect 1444 -1609 1445 -1567
rect 289 -1570 290 -1480
rect 345 -1609 346 -1569
rect 688 -1609 689 -1569
rect 1010 -1570 1011 -1480
rect 1430 -1609 1431 -1569
rect 1465 -1570 1466 -1480
rect 177 -1572 178 -1480
rect 289 -1609 290 -1571
rect 614 -1572 615 -1480
rect 1465 -1609 1466 -1571
rect 177 -1609 178 -1573
rect 411 -1574 412 -1480
rect 716 -1609 717 -1573
rect 1108 -1574 1109 -1480
rect 723 -1576 724 -1480
rect 1717 -1609 1718 -1575
rect 723 -1609 724 -1577
rect 744 -1578 745 -1480
rect 772 -1609 773 -1577
rect 856 -1578 857 -1480
rect 1010 -1609 1011 -1577
rect 1052 -1578 1053 -1480
rect 1108 -1609 1109 -1577
rect 1192 -1578 1193 -1480
rect 548 -1609 549 -1579
rect 744 -1609 745 -1579
rect 821 -1609 822 -1579
rect 1164 -1580 1165 -1480
rect 1192 -1609 1193 -1579
rect 1269 -1580 1270 -1480
rect 614 -1609 615 -1581
rect 1269 -1609 1270 -1581
rect 726 -1609 727 -1583
rect 954 -1584 955 -1480
rect 1052 -1609 1053 -1583
rect 1080 -1584 1081 -1480
rect 1164 -1609 1165 -1583
rect 1220 -1584 1221 -1480
rect 828 -1609 829 -1585
rect 877 -1586 878 -1480
rect 954 -1609 955 -1585
rect 1101 -1586 1102 -1480
rect 1220 -1609 1221 -1585
rect 1248 -1586 1249 -1480
rect 849 -1588 850 -1480
rect 856 -1609 857 -1587
rect 877 -1609 878 -1587
rect 884 -1588 885 -1480
rect 1080 -1609 1081 -1587
rect 1150 -1588 1151 -1480
rect 1248 -1609 1249 -1587
rect 1304 -1588 1305 -1480
rect 702 -1590 703 -1480
rect 884 -1609 885 -1589
rect 1101 -1609 1102 -1589
rect 1381 -1590 1382 -1480
rect 292 -1609 293 -1591
rect 702 -1609 703 -1591
rect 849 -1609 850 -1591
rect 1003 -1592 1004 -1480
rect 1304 -1609 1305 -1591
rect 1409 -1592 1410 -1480
rect 541 -1609 542 -1593
rect 1409 -1609 1410 -1593
rect 1003 -1609 1004 -1595
rect 1038 -1596 1039 -1480
rect 1381 -1609 1382 -1595
rect 1458 -1596 1459 -1480
rect 1038 -1609 1039 -1597
rect 1178 -1598 1179 -1480
rect 1458 -1609 1459 -1597
rect 1479 -1598 1480 -1480
rect 1178 -1609 1179 -1599
rect 1276 -1600 1277 -1480
rect 1479 -1609 1480 -1599
rect 1647 -1600 1648 -1480
rect 264 -1602 265 -1480
rect 1647 -1609 1648 -1601
rect 1276 -1609 1277 -1603
rect 1388 -1604 1389 -1480
rect 1388 -1609 1389 -1605
rect 1514 -1606 1515 -1480
rect 642 -1608 643 -1480
rect 1514 -1609 1515 -1607
rect 16 -1736 17 -1618
rect 30 -1619 31 -1617
rect 37 -1736 38 -1618
rect 289 -1619 290 -1617
rect 296 -1619 297 -1617
rect 383 -1619 384 -1617
rect 411 -1736 412 -1618
rect 744 -1736 745 -1618
rect 758 -1619 759 -1617
rect 1104 -1619 1105 -1617
rect 1115 -1619 1116 -1617
rect 1318 -1619 1319 -1617
rect 1381 -1619 1382 -1617
rect 1384 -1619 1385 -1617
rect 1479 -1619 1480 -1617
rect 1724 -1736 1725 -1618
rect 1752 -1619 1753 -1617
rect 1766 -1736 1767 -1618
rect 44 -1621 45 -1617
rect 254 -1621 255 -1617
rect 268 -1621 269 -1617
rect 310 -1621 311 -1617
rect 317 -1736 318 -1620
rect 915 -1736 916 -1620
rect 929 -1621 930 -1617
rect 1682 -1621 1683 -1617
rect 1717 -1621 1718 -1617
rect 1780 -1736 1781 -1620
rect 44 -1736 45 -1622
rect 345 -1623 346 -1617
rect 348 -1736 349 -1622
rect 919 -1623 920 -1617
rect 933 -1623 934 -1617
rect 933 -1736 934 -1622
rect 933 -1623 934 -1617
rect 933 -1736 934 -1622
rect 961 -1623 962 -1617
rect 961 -1736 962 -1622
rect 961 -1623 962 -1617
rect 961 -1736 962 -1622
rect 996 -1623 997 -1617
rect 1773 -1736 1774 -1622
rect 58 -1736 59 -1624
rect 1542 -1625 1543 -1617
rect 1626 -1625 1627 -1617
rect 1731 -1736 1732 -1624
rect 65 -1736 66 -1626
rect 495 -1627 496 -1617
rect 513 -1627 514 -1617
rect 726 -1627 727 -1617
rect 730 -1627 731 -1617
rect 758 -1736 759 -1626
rect 761 -1627 762 -1617
rect 1661 -1627 1662 -1617
rect 1668 -1627 1669 -1617
rect 1703 -1627 1704 -1617
rect 72 -1629 73 -1617
rect 72 -1736 73 -1628
rect 72 -1629 73 -1617
rect 72 -1736 73 -1628
rect 79 -1629 80 -1617
rect 264 -1736 265 -1628
rect 268 -1736 269 -1628
rect 320 -1629 321 -1617
rect 324 -1629 325 -1617
rect 366 -1629 367 -1617
rect 369 -1629 370 -1617
rect 415 -1629 416 -1617
rect 432 -1736 433 -1628
rect 457 -1629 458 -1617
rect 478 -1629 479 -1617
rect 614 -1629 615 -1617
rect 632 -1629 633 -1617
rect 632 -1736 633 -1628
rect 632 -1629 633 -1617
rect 632 -1736 633 -1628
rect 639 -1629 640 -1617
rect 639 -1736 640 -1628
rect 639 -1629 640 -1617
rect 639 -1736 640 -1628
rect 667 -1629 668 -1617
rect 814 -1629 815 -1617
rect 828 -1629 829 -1617
rect 894 -1736 895 -1628
rect 919 -1736 920 -1628
rect 922 -1736 923 -1628
rect 975 -1629 976 -1617
rect 1661 -1736 1662 -1628
rect 23 -1631 24 -1617
rect 366 -1736 367 -1630
rect 373 -1631 374 -1617
rect 373 -1736 374 -1630
rect 373 -1631 374 -1617
rect 373 -1736 374 -1630
rect 387 -1631 388 -1617
rect 457 -1736 458 -1630
rect 513 -1736 514 -1630
rect 607 -1631 608 -1617
rect 667 -1736 668 -1630
rect 695 -1631 696 -1617
rect 712 -1631 713 -1617
rect 1024 -1631 1025 -1617
rect 1048 -1631 1049 -1617
rect 1612 -1631 1613 -1617
rect 1640 -1631 1641 -1617
rect 1738 -1736 1739 -1630
rect 61 -1736 62 -1632
rect 387 -1736 388 -1632
rect 450 -1633 451 -1617
rect 789 -1736 790 -1632
rect 793 -1633 794 -1617
rect 1395 -1633 1396 -1617
rect 1486 -1633 1487 -1617
rect 1668 -1736 1669 -1632
rect 79 -1736 80 -1634
rect 548 -1635 549 -1617
rect 562 -1635 563 -1617
rect 1318 -1736 1319 -1634
rect 1381 -1736 1382 -1634
rect 1402 -1635 1403 -1617
rect 1500 -1635 1501 -1617
rect 1626 -1736 1627 -1634
rect 1640 -1736 1641 -1634
rect 1675 -1635 1676 -1617
rect 121 -1637 122 -1617
rect 544 -1637 545 -1617
rect 548 -1736 549 -1636
rect 555 -1637 556 -1617
rect 576 -1637 577 -1617
rect 926 -1637 927 -1617
rect 975 -1736 976 -1636
rect 1458 -1637 1459 -1617
rect 1514 -1637 1515 -1617
rect 1682 -1736 1683 -1636
rect 121 -1736 122 -1638
rect 716 -1639 717 -1617
rect 726 -1736 727 -1638
rect 898 -1639 899 -1617
rect 996 -1736 997 -1638
rect 1038 -1639 1039 -1617
rect 1059 -1639 1060 -1617
rect 1444 -1639 1445 -1617
rect 1521 -1639 1522 -1617
rect 1717 -1736 1718 -1638
rect 135 -1641 136 -1617
rect 618 -1641 619 -1617
rect 674 -1641 675 -1617
rect 740 -1641 741 -1617
rect 803 -1736 804 -1640
rect 814 -1736 815 -1640
rect 863 -1641 864 -1617
rect 1059 -1736 1060 -1640
rect 1115 -1736 1116 -1640
rect 1458 -1736 1459 -1640
rect 1591 -1641 1592 -1617
rect 1675 -1736 1676 -1640
rect 135 -1736 136 -1642
rect 681 -1643 682 -1617
rect 702 -1643 703 -1617
rect 793 -1736 794 -1642
rect 807 -1643 808 -1617
rect 1024 -1736 1025 -1642
rect 1118 -1643 1119 -1617
rect 1234 -1643 1235 -1617
rect 1241 -1643 1242 -1617
rect 1486 -1736 1487 -1642
rect 1598 -1643 1599 -1617
rect 1703 -1736 1704 -1642
rect 156 -1645 157 -1617
rect 415 -1736 416 -1644
rect 450 -1736 451 -1644
rect 747 -1645 748 -1617
rect 807 -1736 808 -1644
rect 898 -1736 899 -1644
rect 992 -1736 993 -1644
rect 1591 -1736 1592 -1644
rect 1647 -1645 1648 -1617
rect 1752 -1736 1753 -1644
rect 156 -1736 157 -1646
rect 982 -1647 983 -1617
rect 1003 -1647 1004 -1617
rect 1003 -1736 1004 -1646
rect 1003 -1647 1004 -1617
rect 1003 -1736 1004 -1646
rect 1052 -1647 1053 -1617
rect 1241 -1736 1242 -1646
rect 1251 -1736 1252 -1646
rect 1689 -1647 1690 -1617
rect 170 -1649 171 -1617
rect 324 -1736 325 -1648
rect 338 -1649 339 -1617
rect 716 -1736 717 -1648
rect 733 -1736 734 -1648
rect 968 -1649 969 -1617
rect 982 -1736 983 -1648
rect 1017 -1649 1018 -1617
rect 1101 -1649 1102 -1617
rect 1647 -1736 1648 -1648
rect 1654 -1649 1655 -1617
rect 1759 -1736 1760 -1648
rect 170 -1736 171 -1650
rect 331 -1651 332 -1617
rect 338 -1736 339 -1650
rect 646 -1651 647 -1617
rect 709 -1651 710 -1617
rect 1038 -1736 1039 -1650
rect 1101 -1736 1102 -1650
rect 1171 -1651 1172 -1617
rect 1213 -1651 1214 -1617
rect 1500 -1736 1501 -1650
rect 1689 -1736 1690 -1650
rect 1710 -1651 1711 -1617
rect 191 -1653 192 -1617
rect 271 -1653 272 -1617
rect 289 -1736 290 -1652
rect 849 -1653 850 -1617
rect 863 -1736 864 -1652
rect 884 -1653 885 -1617
rect 887 -1736 888 -1652
rect 1430 -1653 1431 -1617
rect 1437 -1653 1438 -1617
rect 1521 -1736 1522 -1652
rect 1619 -1653 1620 -1617
rect 1710 -1736 1711 -1652
rect 191 -1736 192 -1654
rect 870 -1655 871 -1617
rect 968 -1736 969 -1654
rect 989 -1655 990 -1617
rect 1010 -1655 1011 -1617
rect 1052 -1736 1053 -1654
rect 1153 -1655 1154 -1617
rect 1332 -1655 1333 -1617
rect 1367 -1655 1368 -1617
rect 1430 -1736 1431 -1654
rect 1465 -1655 1466 -1617
rect 1598 -1736 1599 -1654
rect 194 -1657 195 -1617
rect 1556 -1657 1557 -1617
rect 205 -1659 206 -1617
rect 1234 -1736 1235 -1658
rect 1255 -1659 1256 -1617
rect 1472 -1659 1473 -1617
rect 1493 -1659 1494 -1617
rect 1556 -1736 1557 -1658
rect 51 -1661 52 -1617
rect 205 -1736 206 -1660
rect 208 -1661 209 -1617
rect 1696 -1661 1697 -1617
rect 51 -1736 52 -1662
rect 408 -1663 409 -1617
rect 422 -1663 423 -1617
rect 709 -1736 710 -1662
rect 737 -1663 738 -1617
rect 1605 -1663 1606 -1617
rect 177 -1665 178 -1617
rect 1255 -1736 1256 -1664
rect 1262 -1665 1263 -1617
rect 1444 -1736 1445 -1664
rect 1507 -1665 1508 -1617
rect 1619 -1736 1620 -1664
rect 212 -1667 213 -1617
rect 310 -1736 311 -1666
rect 331 -1736 332 -1666
rect 978 -1736 979 -1666
rect 1066 -1667 1067 -1617
rect 1472 -1736 1473 -1666
rect 1563 -1667 1564 -1617
rect 1696 -1736 1697 -1666
rect 86 -1669 87 -1617
rect 212 -1736 213 -1668
rect 226 -1669 227 -1617
rect 576 -1736 577 -1668
rect 597 -1669 598 -1617
rect 600 -1727 601 -1668
rect 604 -1669 605 -1617
rect 1122 -1669 1123 -1617
rect 1206 -1669 1207 -1617
rect 1332 -1736 1333 -1668
rect 1367 -1736 1368 -1668
rect 1549 -1669 1550 -1617
rect 1563 -1736 1564 -1668
rect 1706 -1669 1707 -1617
rect 86 -1736 87 -1670
rect 142 -1671 143 -1617
rect 184 -1671 185 -1617
rect 226 -1736 227 -1670
rect 233 -1671 234 -1617
rect 1017 -1736 1018 -1670
rect 1066 -1736 1067 -1670
rect 1437 -1736 1438 -1670
rect 1535 -1671 1536 -1617
rect 1549 -1736 1550 -1670
rect 1584 -1671 1585 -1617
rect 1605 -1736 1606 -1670
rect 142 -1736 143 -1672
rect 163 -1673 164 -1617
rect 184 -1736 185 -1672
rect 198 -1673 199 -1617
rect 233 -1736 234 -1672
rect 261 -1673 262 -1617
rect 278 -1736 279 -1672
rect 1010 -1736 1011 -1672
rect 1073 -1673 1074 -1617
rect 1122 -1736 1123 -1672
rect 1157 -1673 1158 -1617
rect 1206 -1736 1207 -1672
rect 1220 -1673 1221 -1617
rect 1220 -1736 1221 -1672
rect 1220 -1673 1221 -1617
rect 1220 -1736 1221 -1672
rect 1269 -1673 1270 -1617
rect 1542 -1736 1543 -1672
rect 107 -1675 108 -1617
rect 163 -1736 164 -1674
rect 240 -1675 241 -1617
rect 422 -1736 423 -1674
rect 436 -1675 437 -1617
rect 989 -1736 990 -1674
rect 1073 -1736 1074 -1674
rect 1227 -1675 1228 -1617
rect 1276 -1675 1277 -1617
rect 1479 -1736 1480 -1674
rect 100 -1677 101 -1617
rect 107 -1736 108 -1676
rect 149 -1677 150 -1617
rect 198 -1736 199 -1676
rect 240 -1736 241 -1676
rect 282 -1677 283 -1617
rect 296 -1736 297 -1676
rect 429 -1677 430 -1617
rect 436 -1736 437 -1676
rect 660 -1677 661 -1617
rect 772 -1677 773 -1617
rect 849 -1736 850 -1676
rect 870 -1736 871 -1676
rect 877 -1677 878 -1617
rect 905 -1677 906 -1617
rect 1262 -1736 1263 -1676
rect 1304 -1677 1305 -1617
rect 1395 -1736 1396 -1676
rect 1416 -1677 1417 -1617
rect 1493 -1736 1494 -1676
rect 100 -1736 101 -1678
rect 429 -1736 430 -1678
rect 478 -1736 479 -1678
rect 681 -1736 682 -1678
rect 751 -1679 752 -1617
rect 772 -1736 773 -1678
rect 782 -1736 783 -1678
rect 1584 -1736 1585 -1678
rect 149 -1736 150 -1680
rect 677 -1736 678 -1680
rect 751 -1736 752 -1680
rect 842 -1681 843 -1617
rect 877 -1736 878 -1680
rect 891 -1681 892 -1617
rect 905 -1736 906 -1680
rect 954 -1681 955 -1617
rect 1020 -1681 1021 -1617
rect 1276 -1736 1277 -1680
rect 1339 -1681 1340 -1617
rect 1416 -1736 1417 -1680
rect 1423 -1681 1424 -1617
rect 1514 -1736 1515 -1680
rect 282 -1736 283 -1682
rect 464 -1683 465 -1617
rect 492 -1683 493 -1617
rect 1654 -1736 1655 -1682
rect 359 -1685 360 -1617
rect 464 -1736 465 -1684
rect 471 -1685 472 -1617
rect 492 -1736 493 -1684
rect 499 -1685 500 -1617
rect 695 -1736 696 -1684
rect 796 -1685 797 -1617
rect 1213 -1736 1214 -1684
rect 1339 -1736 1340 -1684
rect 1346 -1685 1347 -1617
rect 1353 -1685 1354 -1617
rect 1423 -1736 1424 -1684
rect 352 -1687 353 -1617
rect 471 -1736 472 -1686
rect 499 -1736 500 -1686
rect 520 -1687 521 -1617
rect 527 -1687 528 -1617
rect 1633 -1687 1634 -1617
rect 219 -1689 220 -1617
rect 352 -1736 353 -1688
rect 359 -1736 360 -1688
rect 1045 -1689 1046 -1617
rect 1118 -1736 1119 -1688
rect 1507 -1736 1508 -1688
rect 1570 -1689 1571 -1617
rect 1633 -1736 1634 -1688
rect 219 -1736 220 -1690
rect 275 -1691 276 -1617
rect 380 -1691 381 -1617
rect 527 -1736 528 -1690
rect 534 -1691 535 -1617
rect 555 -1736 556 -1690
rect 562 -1736 563 -1690
rect 740 -1736 741 -1690
rect 884 -1736 885 -1690
rect 954 -1736 955 -1690
rect 1150 -1691 1151 -1617
rect 1353 -1736 1354 -1690
rect 1374 -1691 1375 -1617
rect 1465 -1736 1466 -1690
rect 1528 -1691 1529 -1617
rect 1570 -1736 1571 -1690
rect 173 -1736 174 -1692
rect 275 -1736 276 -1692
rect 380 -1736 381 -1692
rect 481 -1736 482 -1692
rect 520 -1736 521 -1692
rect 723 -1693 724 -1617
rect 912 -1693 913 -1617
rect 1157 -1736 1158 -1692
rect 1164 -1693 1165 -1617
rect 1227 -1736 1228 -1692
rect 1283 -1693 1284 -1617
rect 1346 -1736 1347 -1692
rect 1374 -1736 1375 -1692
rect 1409 -1693 1410 -1617
rect 177 -1736 178 -1694
rect 1528 -1736 1529 -1694
rect 443 -1697 444 -1617
rect 842 -1736 843 -1696
rect 873 -1736 874 -1696
rect 1409 -1736 1410 -1696
rect 443 -1736 444 -1698
rect 530 -1699 531 -1617
rect 534 -1736 535 -1698
rect 565 -1699 566 -1617
rect 569 -1699 570 -1617
rect 660 -1736 661 -1698
rect 723 -1736 724 -1698
rect 856 -1699 857 -1617
rect 940 -1699 941 -1617
rect 1045 -1736 1046 -1698
rect 1087 -1699 1088 -1617
rect 1150 -1736 1151 -1698
rect 1178 -1699 1179 -1617
rect 1304 -1736 1305 -1698
rect 1388 -1699 1389 -1617
rect 1535 -1736 1536 -1698
rect 530 -1736 531 -1700
rect 835 -1701 836 -1617
rect 929 -1736 930 -1700
rect 1087 -1736 1088 -1700
rect 1108 -1701 1109 -1617
rect 1164 -1736 1165 -1700
rect 1185 -1701 1186 -1617
rect 1269 -1736 1270 -1700
rect 1297 -1701 1298 -1617
rect 1388 -1736 1389 -1700
rect 128 -1703 129 -1617
rect 835 -1736 836 -1702
rect 940 -1736 941 -1702
rect 947 -1703 948 -1617
rect 1094 -1703 1095 -1617
rect 1185 -1736 1186 -1702
rect 1199 -1703 1200 -1617
rect 1283 -1736 1284 -1702
rect 1290 -1703 1291 -1617
rect 1297 -1736 1298 -1702
rect 93 -1705 94 -1617
rect 128 -1736 129 -1704
rect 541 -1705 542 -1617
rect 1577 -1705 1578 -1617
rect 93 -1736 94 -1706
rect 730 -1736 731 -1706
rect 765 -1707 766 -1617
rect 856 -1736 857 -1706
rect 1108 -1736 1109 -1706
rect 1143 -1707 1144 -1617
rect 1192 -1707 1193 -1617
rect 1290 -1736 1291 -1706
rect 1451 -1707 1452 -1617
rect 1577 -1736 1578 -1706
rect 96 -1709 97 -1617
rect 947 -1736 948 -1708
rect 1129 -1709 1130 -1617
rect 1143 -1736 1144 -1708
rect 1360 -1709 1361 -1617
rect 1451 -1736 1452 -1708
rect 159 -1736 160 -1710
rect 1129 -1736 1130 -1710
rect 1136 -1711 1137 -1617
rect 1199 -1736 1200 -1710
rect 1325 -1711 1326 -1617
rect 1360 -1736 1361 -1710
rect 247 -1713 248 -1617
rect 1136 -1736 1137 -1712
rect 1311 -1713 1312 -1617
rect 1325 -1736 1326 -1712
rect 247 -1736 248 -1714
rect 257 -1736 258 -1714
rect 506 -1715 507 -1617
rect 765 -1736 766 -1714
rect 821 -1715 822 -1617
rect 1192 -1736 1193 -1714
rect 1248 -1715 1249 -1617
rect 1311 -1736 1312 -1714
rect 394 -1717 395 -1617
rect 506 -1736 507 -1716
rect 544 -1736 545 -1716
rect 618 -1736 619 -1716
rect 621 -1717 622 -1617
rect 1171 -1736 1172 -1716
rect 394 -1736 395 -1718
rect 401 -1719 402 -1617
rect 569 -1736 570 -1718
rect 719 -1719 720 -1617
rect 800 -1719 801 -1617
rect 821 -1736 822 -1718
rect 828 -1736 829 -1718
rect 1094 -1736 1095 -1718
rect 401 -1736 402 -1720
rect 541 -1736 542 -1720
rect 583 -1721 584 -1617
rect 604 -1736 605 -1720
rect 611 -1721 612 -1617
rect 1612 -1736 1613 -1720
rect 114 -1723 115 -1617
rect 611 -1736 612 -1722
rect 646 -1736 647 -1722
rect 653 -1723 654 -1617
rect 670 -1723 671 -1617
rect 1178 -1736 1179 -1722
rect 114 -1736 115 -1724
rect 590 -1725 591 -1617
rect 597 -1736 598 -1724
rect 653 -1736 654 -1724
rect 786 -1725 787 -1617
rect 800 -1736 801 -1724
rect 1080 -1725 1081 -1617
rect 303 -1727 304 -1617
rect 583 -1736 584 -1726
rect 590 -1736 591 -1726
rect 688 -1727 689 -1617
rect 1031 -1727 1032 -1617
rect 1080 -1736 1081 -1726
rect 1384 -1736 1385 -1726
rect 1402 -1736 1403 -1726
rect 303 -1736 304 -1728
rect 1748 -1736 1749 -1728
rect 688 -1736 689 -1730
rect 779 -1731 780 -1617
rect 926 -1736 927 -1730
rect 1031 -1736 1032 -1730
rect 485 -1733 486 -1617
rect 779 -1736 780 -1732
rect 345 -1736 346 -1734
rect 485 -1736 486 -1734
rect 30 -1883 31 -1745
rect 128 -1746 129 -1744
rect 159 -1746 160 -1744
rect 530 -1746 531 -1744
rect 534 -1746 535 -1744
rect 534 -1883 535 -1745
rect 534 -1746 535 -1744
rect 534 -1883 535 -1745
rect 541 -1746 542 -1744
rect 765 -1746 766 -1744
rect 810 -1746 811 -1744
rect 877 -1746 878 -1744
rect 884 -1883 885 -1745
rect 940 -1746 941 -1744
rect 978 -1746 979 -1744
rect 1598 -1746 1599 -1744
rect 1682 -1746 1683 -1744
rect 1794 -1883 1795 -1745
rect 58 -1883 59 -1747
rect 499 -1748 500 -1744
rect 502 -1883 503 -1747
rect 842 -1748 843 -1744
rect 866 -1883 867 -1747
rect 1808 -1883 1809 -1747
rect 61 -1750 62 -1744
rect 352 -1750 353 -1744
rect 401 -1750 402 -1744
rect 940 -1883 941 -1749
rect 989 -1750 990 -1744
rect 1647 -1750 1648 -1744
rect 1748 -1750 1749 -1744
rect 1766 -1750 1767 -1744
rect 1780 -1750 1781 -1744
rect 1815 -1883 1816 -1749
rect 65 -1752 66 -1744
rect 254 -1752 255 -1744
rect 264 -1752 265 -1744
rect 264 -1883 265 -1751
rect 264 -1752 265 -1744
rect 264 -1883 265 -1751
rect 275 -1752 276 -1744
rect 415 -1752 416 -1744
rect 450 -1752 451 -1744
rect 1248 -1752 1249 -1744
rect 1367 -1752 1368 -1744
rect 1682 -1883 1683 -1751
rect 1752 -1752 1753 -1744
rect 1766 -1883 1767 -1751
rect 65 -1883 66 -1753
rect 170 -1754 171 -1744
rect 177 -1754 178 -1744
rect 1626 -1754 1627 -1744
rect 1738 -1754 1739 -1744
rect 1752 -1883 1753 -1753
rect 1759 -1754 1760 -1744
rect 1759 -1883 1760 -1753
rect 1759 -1754 1760 -1744
rect 1759 -1883 1760 -1753
rect 107 -1756 108 -1744
rect 128 -1883 129 -1755
rect 159 -1883 160 -1755
rect 296 -1756 297 -1744
rect 324 -1756 325 -1744
rect 481 -1756 482 -1744
rect 604 -1756 605 -1744
rect 604 -1883 605 -1755
rect 604 -1756 605 -1744
rect 604 -1883 605 -1755
rect 618 -1756 619 -1744
rect 730 -1883 731 -1755
rect 740 -1756 741 -1744
rect 1059 -1756 1060 -1744
rect 1069 -1756 1070 -1744
rect 1535 -1756 1536 -1744
rect 1612 -1756 1613 -1744
rect 1647 -1883 1648 -1755
rect 1710 -1756 1711 -1744
rect 1738 -1883 1739 -1755
rect 107 -1883 108 -1757
rect 1192 -1758 1193 -1744
rect 1199 -1758 1200 -1744
rect 1248 -1883 1249 -1757
rect 1332 -1758 1333 -1744
rect 1367 -1883 1368 -1757
rect 1374 -1758 1375 -1744
rect 1535 -1883 1536 -1757
rect 1605 -1758 1606 -1744
rect 1612 -1883 1613 -1757
rect 1626 -1883 1627 -1757
rect 1640 -1758 1641 -1744
rect 1696 -1758 1697 -1744
rect 1710 -1883 1711 -1757
rect 110 -1883 111 -1759
rect 254 -1883 255 -1759
rect 275 -1883 276 -1759
rect 800 -1760 801 -1744
rect 814 -1760 815 -1744
rect 842 -1883 843 -1759
rect 870 -1760 871 -1744
rect 1059 -1883 1060 -1759
rect 1080 -1760 1081 -1744
rect 1115 -1760 1116 -1744
rect 1160 -1883 1161 -1759
rect 1213 -1760 1214 -1744
rect 1374 -1883 1375 -1759
rect 1493 -1760 1494 -1744
rect 1528 -1760 1529 -1744
rect 1640 -1883 1641 -1759
rect 114 -1762 115 -1744
rect 618 -1883 619 -1761
rect 667 -1762 668 -1744
rect 765 -1883 766 -1761
rect 793 -1762 794 -1744
rect 877 -1883 878 -1761
rect 887 -1762 888 -1744
rect 1318 -1762 1319 -1744
rect 1444 -1762 1445 -1744
rect 1493 -1883 1494 -1761
rect 1528 -1883 1529 -1761
rect 1619 -1762 1620 -1744
rect 1633 -1762 1634 -1744
rect 1696 -1883 1697 -1761
rect 114 -1883 115 -1763
rect 366 -1764 367 -1744
rect 408 -1883 409 -1763
rect 485 -1764 486 -1744
rect 625 -1764 626 -1744
rect 667 -1883 668 -1763
rect 677 -1764 678 -1744
rect 772 -1764 773 -1744
rect 800 -1883 801 -1763
rect 1045 -1764 1046 -1744
rect 1052 -1764 1053 -1744
rect 1052 -1883 1053 -1763
rect 1052 -1764 1053 -1744
rect 1052 -1883 1053 -1763
rect 1073 -1764 1074 -1744
rect 1080 -1883 1081 -1763
rect 1108 -1764 1109 -1744
rect 1199 -1883 1200 -1763
rect 1276 -1764 1277 -1744
rect 1318 -1883 1319 -1763
rect 1430 -1764 1431 -1744
rect 1444 -1883 1445 -1763
rect 1563 -1764 1564 -1744
rect 1605 -1883 1606 -1763
rect 149 -1766 150 -1744
rect 1073 -1883 1074 -1765
rect 1111 -1883 1112 -1765
rect 1668 -1766 1669 -1744
rect 149 -1883 150 -1767
rect 184 -1768 185 -1744
rect 191 -1768 192 -1744
rect 436 -1768 437 -1744
rect 478 -1768 479 -1744
rect 1780 -1883 1781 -1767
rect 170 -1883 171 -1769
rect 810 -1883 811 -1769
rect 821 -1770 822 -1744
rect 870 -1883 871 -1769
rect 891 -1770 892 -1744
rect 1479 -1770 1480 -1744
rect 1549 -1770 1550 -1744
rect 1668 -1883 1669 -1769
rect 180 -1772 181 -1744
rect 422 -1772 423 -1744
rect 436 -1883 437 -1771
rect 443 -1772 444 -1744
rect 625 -1883 626 -1771
rect 726 -1772 727 -1744
rect 733 -1772 734 -1744
rect 1479 -1883 1480 -1771
rect 1584 -1772 1585 -1744
rect 1619 -1883 1620 -1771
rect 180 -1883 181 -1773
rect 1661 -1774 1662 -1744
rect 184 -1883 185 -1775
rect 548 -1776 549 -1744
rect 688 -1776 689 -1744
rect 982 -1776 983 -1744
rect 989 -1883 990 -1775
rect 1031 -1776 1032 -1744
rect 1041 -1883 1042 -1775
rect 1269 -1776 1270 -1744
rect 1279 -1883 1280 -1775
rect 1549 -1883 1550 -1775
rect 1570 -1776 1571 -1744
rect 1661 -1883 1662 -1775
rect 191 -1883 192 -1777
rect 1654 -1778 1655 -1744
rect 208 -1883 209 -1779
rect 541 -1883 542 -1779
rect 548 -1883 549 -1779
rect 1010 -1780 1011 -1744
rect 1017 -1780 1018 -1744
rect 1213 -1883 1214 -1779
rect 1234 -1780 1235 -1744
rect 1430 -1883 1431 -1779
rect 1521 -1780 1522 -1744
rect 1584 -1883 1585 -1779
rect 1591 -1780 1592 -1744
rect 1654 -1883 1655 -1779
rect 233 -1782 234 -1744
rect 341 -1883 342 -1781
rect 348 -1782 349 -1744
rect 835 -1782 836 -1744
rect 849 -1782 850 -1744
rect 891 -1883 892 -1781
rect 915 -1782 916 -1744
rect 1388 -1782 1389 -1744
rect 1507 -1782 1508 -1744
rect 1591 -1883 1592 -1781
rect 233 -1883 234 -1783
rect 432 -1784 433 -1744
rect 576 -1784 577 -1744
rect 688 -1883 689 -1783
rect 695 -1784 696 -1744
rect 786 -1883 787 -1783
rect 821 -1883 822 -1783
rect 1283 -1784 1284 -1744
rect 1381 -1784 1382 -1744
rect 1521 -1883 1522 -1783
rect 1556 -1784 1557 -1744
rect 1570 -1883 1571 -1783
rect 240 -1786 241 -1744
rect 240 -1883 241 -1785
rect 240 -1786 241 -1744
rect 240 -1883 241 -1785
rect 268 -1786 269 -1744
rect 366 -1883 367 -1785
rect 411 -1786 412 -1744
rect 803 -1786 804 -1744
rect 824 -1883 825 -1785
rect 1633 -1883 1634 -1785
rect 268 -1883 269 -1787
rect 569 -1788 570 -1744
rect 576 -1883 577 -1787
rect 894 -1788 895 -1744
rect 919 -1788 920 -1744
rect 1724 -1788 1725 -1744
rect 282 -1790 283 -1744
rect 296 -1883 297 -1789
rect 317 -1790 318 -1744
rect 478 -1883 479 -1789
rect 632 -1790 633 -1744
rect 695 -1883 696 -1789
rect 702 -1790 703 -1744
rect 1171 -1790 1172 -1744
rect 1220 -1790 1221 -1744
rect 1234 -1883 1235 -1789
rect 1269 -1883 1270 -1789
rect 1311 -1790 1312 -1744
rect 1465 -1790 1466 -1744
rect 1507 -1883 1508 -1789
rect 1703 -1790 1704 -1744
rect 1724 -1883 1725 -1789
rect 156 -1792 157 -1744
rect 1465 -1883 1466 -1791
rect 1675 -1792 1676 -1744
rect 1703 -1883 1704 -1791
rect 156 -1883 157 -1793
rect 632 -1883 633 -1793
rect 639 -1794 640 -1744
rect 702 -1883 703 -1793
rect 709 -1794 710 -1744
rect 793 -1883 794 -1793
rect 828 -1794 829 -1744
rect 1157 -1794 1158 -1744
rect 1171 -1883 1172 -1793
rect 1804 -1883 1805 -1793
rect 198 -1796 199 -1744
rect 317 -1883 318 -1795
rect 324 -1883 325 -1795
rect 394 -1796 395 -1744
rect 415 -1883 416 -1795
rect 922 -1796 923 -1744
rect 926 -1796 927 -1744
rect 1136 -1796 1137 -1744
rect 1157 -1883 1158 -1795
rect 1416 -1796 1417 -1744
rect 1675 -1883 1676 -1795
rect 1689 -1796 1690 -1744
rect 198 -1883 199 -1797
rect 513 -1798 514 -1744
rect 639 -1883 640 -1797
rect 646 -1798 647 -1744
rect 709 -1883 710 -1797
rect 1066 -1798 1067 -1744
rect 1115 -1883 1116 -1797
rect 1164 -1798 1165 -1744
rect 1178 -1798 1179 -1744
rect 1220 -1883 1221 -1797
rect 1276 -1883 1277 -1797
rect 1689 -1883 1690 -1797
rect 247 -1800 248 -1744
rect 282 -1883 283 -1799
rect 289 -1800 290 -1744
rect 1136 -1883 1137 -1799
rect 1283 -1883 1284 -1799
rect 1290 -1800 1291 -1744
rect 1416 -1883 1417 -1799
rect 1745 -1800 1746 -1744
rect 121 -1802 122 -1744
rect 289 -1883 290 -1801
rect 310 -1802 311 -1744
rect 394 -1883 395 -1801
rect 422 -1883 423 -1801
rect 674 -1802 675 -1744
rect 716 -1802 717 -1744
rect 1010 -1883 1011 -1801
rect 1017 -1883 1018 -1801
rect 1486 -1802 1487 -1744
rect 1731 -1802 1732 -1744
rect 1745 -1883 1746 -1801
rect 93 -1804 94 -1744
rect 716 -1883 717 -1803
rect 737 -1804 738 -1744
rect 1381 -1883 1382 -1803
rect 1717 -1804 1718 -1744
rect 1731 -1883 1732 -1803
rect 93 -1883 94 -1805
rect 257 -1806 258 -1744
rect 303 -1806 304 -1744
rect 737 -1883 738 -1805
rect 744 -1806 745 -1744
rect 912 -1806 913 -1744
rect 919 -1883 920 -1805
rect 1776 -1883 1777 -1805
rect 79 -1808 80 -1744
rect 303 -1883 304 -1807
rect 331 -1808 332 -1744
rect 352 -1883 353 -1807
rect 359 -1808 360 -1744
rect 485 -1883 486 -1807
rect 674 -1883 675 -1807
rect 1108 -1883 1109 -1807
rect 1153 -1883 1154 -1807
rect 1486 -1883 1487 -1807
rect 79 -1883 80 -1809
rect 380 -1810 381 -1744
rect 446 -1883 447 -1809
rect 1556 -1883 1557 -1809
rect 121 -1883 122 -1811
rect 506 -1812 507 -1744
rect 744 -1883 745 -1811
rect 751 -1812 752 -1744
rect 758 -1812 759 -1744
rect 814 -1883 815 -1811
rect 828 -1883 829 -1811
rect 1787 -1883 1788 -1811
rect 135 -1814 136 -1744
rect 758 -1883 759 -1813
rect 772 -1883 773 -1813
rect 1801 -1883 1802 -1813
rect 100 -1816 101 -1744
rect 135 -1883 136 -1815
rect 205 -1816 206 -1744
rect 310 -1883 311 -1815
rect 331 -1883 332 -1815
rect 443 -1883 444 -1815
rect 464 -1816 465 -1744
rect 513 -1883 514 -1815
rect 611 -1816 612 -1744
rect 751 -1883 752 -1815
rect 789 -1816 790 -1744
rect 1717 -1883 1718 -1815
rect 100 -1883 101 -1817
rect 226 -1818 227 -1744
rect 338 -1818 339 -1744
rect 474 -1883 475 -1817
rect 506 -1883 507 -1817
rect 555 -1818 556 -1744
rect 597 -1818 598 -1744
rect 611 -1883 612 -1817
rect 849 -1883 850 -1817
rect 1087 -1818 1088 -1744
rect 1101 -1818 1102 -1744
rect 1178 -1883 1179 -1817
rect 1290 -1883 1291 -1817
rect 1773 -1818 1774 -1744
rect 86 -1820 87 -1744
rect 555 -1883 556 -1819
rect 597 -1883 598 -1819
rect 779 -1820 780 -1744
rect 863 -1820 864 -1744
rect 1101 -1883 1102 -1819
rect 1542 -1820 1543 -1744
rect 1773 -1883 1774 -1819
rect 72 -1822 73 -1744
rect 86 -1883 87 -1821
rect 205 -1883 206 -1821
rect 1255 -1822 1256 -1744
rect 1458 -1822 1459 -1744
rect 1542 -1883 1543 -1821
rect 44 -1824 45 -1744
rect 72 -1883 73 -1823
rect 212 -1824 213 -1744
rect 779 -1883 780 -1823
rect 863 -1883 864 -1823
rect 1262 -1824 1263 -1744
rect 1423 -1824 1424 -1744
rect 1458 -1883 1459 -1823
rect 44 -1883 45 -1825
rect 163 -1826 164 -1744
rect 212 -1883 213 -1825
rect 492 -1826 493 -1744
rect 912 -1883 913 -1825
rect 954 -1826 955 -1744
rect 982 -1883 983 -1825
rect 1241 -1826 1242 -1744
rect 1339 -1826 1340 -1744
rect 1423 -1883 1424 -1825
rect 163 -1883 164 -1827
rect 831 -1828 832 -1744
rect 926 -1883 927 -1827
rect 1577 -1828 1578 -1744
rect 219 -1830 220 -1744
rect 226 -1883 227 -1829
rect 338 -1883 339 -1829
rect 467 -1883 468 -1829
rect 471 -1830 472 -1744
rect 569 -1883 570 -1829
rect 831 -1883 832 -1829
rect 1332 -1883 1333 -1829
rect 1402 -1830 1403 -1744
rect 1577 -1883 1578 -1829
rect 219 -1883 220 -1831
rect 691 -1832 692 -1744
rect 929 -1832 930 -1744
rect 1500 -1832 1501 -1744
rect 359 -1883 360 -1833
rect 373 -1834 374 -1744
rect 380 -1883 381 -1833
rect 457 -1834 458 -1744
rect 492 -1883 493 -1833
rect 527 -1834 528 -1744
rect 936 -1883 937 -1833
rect 1150 -1834 1151 -1744
rect 1206 -1834 1207 -1744
rect 1255 -1883 1256 -1833
rect 1395 -1834 1396 -1744
rect 1402 -1883 1403 -1833
rect 37 -1836 38 -1744
rect 527 -1883 528 -1835
rect 947 -1836 948 -1744
rect 1388 -1883 1389 -1835
rect 37 -1883 38 -1837
rect 51 -1838 52 -1744
rect 247 -1883 248 -1837
rect 457 -1883 458 -1837
rect 898 -1838 899 -1744
rect 947 -1883 948 -1837
rect 975 -1883 976 -1837
rect 1150 -1883 1151 -1837
rect 1206 -1883 1207 -1837
rect 1304 -1838 1305 -1744
rect 1346 -1838 1347 -1744
rect 1395 -1883 1396 -1837
rect 51 -1883 52 -1839
rect 142 -1840 143 -1744
rect 373 -1883 374 -1839
rect 562 -1840 563 -1744
rect 898 -1883 899 -1839
rect 929 -1883 930 -1839
rect 933 -1840 934 -1744
rect 1346 -1883 1347 -1839
rect 142 -1883 143 -1841
rect 177 -1883 178 -1841
rect 401 -1883 402 -1841
rect 471 -1883 472 -1841
rect 562 -1883 563 -1841
rect 649 -1883 650 -1841
rect 856 -1842 857 -1744
rect 933 -1883 934 -1841
rect 996 -1842 997 -1744
rect 1192 -1883 1193 -1841
rect 1227 -1842 1228 -1744
rect 1262 -1883 1263 -1841
rect 1297 -1842 1298 -1744
rect 1304 -1883 1305 -1841
rect 429 -1883 430 -1843
rect 464 -1883 465 -1843
rect 656 -1883 657 -1843
rect 1227 -1883 1228 -1843
rect 1251 -1844 1252 -1744
rect 1339 -1883 1340 -1843
rect 681 -1846 682 -1744
rect 856 -1883 857 -1845
rect 961 -1846 962 -1744
rect 996 -1883 997 -1845
rect 1003 -1846 1004 -1744
rect 1031 -1883 1032 -1845
rect 1038 -1846 1039 -1744
rect 1087 -1883 1088 -1845
rect 1143 -1846 1144 -1744
rect 1241 -1883 1242 -1845
rect 1297 -1883 1298 -1845
rect 1514 -1846 1515 -1744
rect 345 -1883 346 -1847
rect 1038 -1883 1039 -1847
rect 1045 -1883 1046 -1847
rect 1563 -1883 1564 -1847
rect 583 -1850 584 -1744
rect 681 -1883 682 -1849
rect 835 -1883 836 -1849
rect 1003 -1883 1004 -1849
rect 1024 -1850 1025 -1744
rect 1164 -1883 1165 -1849
rect 1353 -1850 1354 -1744
rect 1514 -1883 1515 -1849
rect 583 -1883 584 -1851
rect 590 -1852 591 -1744
rect 653 -1852 654 -1744
rect 961 -1883 962 -1851
rect 968 -1852 969 -1744
rect 1024 -1883 1025 -1851
rect 1027 -1883 1028 -1851
rect 1598 -1883 1599 -1851
rect 450 -1883 451 -1853
rect 653 -1883 654 -1853
rect 968 -1883 969 -1853
rect 985 -1883 986 -1853
rect 1048 -1883 1049 -1853
rect 1500 -1883 1501 -1853
rect 590 -1883 591 -1855
rect 660 -1856 661 -1744
rect 1066 -1883 1067 -1855
rect 1129 -1856 1130 -1744
rect 1353 -1883 1354 -1855
rect 1472 -1856 1473 -1744
rect 660 -1883 661 -1857
rect 782 -1858 783 -1744
rect 905 -1858 906 -1744
rect 1129 -1883 1130 -1857
rect 1451 -1858 1452 -1744
rect 1472 -1883 1473 -1857
rect 807 -1860 808 -1744
rect 1451 -1883 1452 -1859
rect 905 -1883 906 -1861
rect 1437 -1862 1438 -1744
rect 1094 -1864 1095 -1744
rect 1143 -1883 1144 -1863
rect 1409 -1864 1410 -1744
rect 1437 -1883 1438 -1863
rect 194 -1866 195 -1744
rect 1409 -1883 1410 -1865
rect 1094 -1883 1095 -1867
rect 1122 -1868 1123 -1744
rect 1122 -1883 1123 -1869
rect 1185 -1870 1186 -1744
rect 1185 -1883 1186 -1871
rect 1360 -1872 1361 -1744
rect 1325 -1874 1326 -1744
rect 1360 -1883 1361 -1873
rect 723 -1876 724 -1744
rect 1325 -1883 1326 -1875
rect 387 -1878 388 -1744
rect 723 -1883 724 -1877
rect 387 -1883 388 -1879
rect 520 -1880 521 -1744
rect 250 -1883 251 -1881
rect 520 -1883 521 -1881
rect 51 -1893 52 -1891
rect 215 -2016 216 -1892
rect 233 -1893 234 -1891
rect 887 -2016 888 -1892
rect 905 -1893 906 -1891
rect 1199 -1893 1200 -1891
rect 1216 -2016 1217 -1892
rect 1227 -1893 1228 -1891
rect 1234 -1893 1235 -1891
rect 1234 -2016 1235 -1892
rect 1234 -1893 1235 -1891
rect 1234 -2016 1235 -1892
rect 1276 -1893 1277 -1891
rect 1577 -1893 1578 -1891
rect 1654 -1893 1655 -1891
rect 1804 -1893 1805 -1891
rect 51 -2016 52 -1894
rect 268 -1895 269 -1891
rect 296 -1895 297 -1891
rect 296 -2016 297 -1894
rect 296 -1895 297 -1891
rect 296 -2016 297 -1894
rect 303 -1895 304 -1891
rect 474 -1895 475 -1891
rect 478 -1895 479 -1891
rect 905 -2016 906 -1894
rect 912 -1895 913 -1891
rect 912 -2016 913 -1894
rect 912 -1895 913 -1891
rect 912 -2016 913 -1894
rect 919 -1895 920 -1891
rect 982 -2016 983 -1894
rect 1017 -1895 1018 -1891
rect 1164 -1895 1165 -1891
rect 1171 -1895 1172 -1891
rect 1171 -2016 1172 -1894
rect 1171 -1895 1172 -1891
rect 1171 -2016 1172 -1894
rect 1276 -2016 1277 -1894
rect 1416 -1895 1417 -1891
rect 1668 -1895 1669 -1891
rect 1668 -2016 1669 -1894
rect 1668 -1895 1669 -1891
rect 1668 -2016 1669 -1894
rect 1773 -1895 1774 -1891
rect 1794 -1895 1795 -1891
rect 65 -1897 66 -1891
rect 65 -2016 66 -1896
rect 65 -1897 66 -1891
rect 65 -2016 66 -1896
rect 68 -2016 69 -1896
rect 548 -1897 549 -1891
rect 572 -1897 573 -1891
rect 1346 -1897 1347 -1891
rect 1381 -1897 1382 -1891
rect 1384 -1897 1385 -1891
rect 1409 -1897 1410 -1891
rect 1776 -1897 1777 -1891
rect 1794 -2016 1795 -1896
rect 1808 -1897 1809 -1891
rect 72 -1899 73 -1891
rect 107 -1899 108 -1891
rect 135 -1899 136 -1891
rect 261 -2016 262 -1898
rect 303 -2016 304 -1898
rect 562 -1899 563 -1891
rect 593 -2016 594 -1898
rect 1451 -1899 1452 -1891
rect 1493 -1899 1494 -1891
rect 1808 -2016 1809 -1898
rect 72 -2016 73 -1900
rect 149 -1901 150 -1891
rect 156 -1901 157 -1891
rect 233 -2016 234 -1900
rect 240 -1901 241 -1891
rect 240 -2016 241 -1900
rect 240 -1901 241 -1891
rect 240 -2016 241 -1900
rect 250 -1901 251 -1891
rect 548 -2016 549 -1900
rect 562 -2016 563 -1900
rect 947 -1901 948 -1891
rect 954 -2016 955 -1900
rect 968 -1901 969 -1891
rect 1024 -1901 1025 -1891
rect 1759 -1901 1760 -1891
rect 79 -1903 80 -1891
rect 338 -2016 339 -1902
rect 345 -1903 346 -1891
rect 828 -2016 829 -1902
rect 831 -1903 832 -1891
rect 1101 -1903 1102 -1891
rect 1111 -2016 1112 -1902
rect 1724 -1903 1725 -1891
rect 79 -2016 80 -1904
rect 611 -1905 612 -1891
rect 646 -1905 647 -1891
rect 779 -1905 780 -1891
rect 796 -2016 797 -1904
rect 842 -1905 843 -1891
rect 849 -1905 850 -1891
rect 1199 -2016 1200 -1904
rect 1279 -1905 1280 -1891
rect 1724 -2016 1725 -1904
rect 86 -1907 87 -1891
rect 107 -2016 108 -1906
rect 135 -2016 136 -1906
rect 401 -1907 402 -1891
rect 436 -1907 437 -1891
rect 999 -2016 1000 -1906
rect 1024 -2016 1025 -1906
rect 1143 -1907 1144 -1891
rect 1153 -1907 1154 -1891
rect 1731 -1907 1732 -1891
rect 86 -2016 87 -1908
rect 310 -1909 311 -1891
rect 324 -1909 325 -1891
rect 467 -1909 468 -1891
rect 499 -2016 500 -1908
rect 866 -1909 867 -1891
rect 922 -2016 923 -1908
rect 985 -1909 986 -1891
rect 1031 -1909 1032 -1891
rect 1101 -2016 1102 -1908
rect 1115 -1909 1116 -1891
rect 1227 -2016 1228 -1908
rect 1283 -1909 1284 -1891
rect 1283 -2016 1284 -1908
rect 1283 -1909 1284 -1891
rect 1283 -2016 1284 -1908
rect 1314 -1909 1315 -1891
rect 1633 -1909 1634 -1891
rect 1731 -2016 1732 -1908
rect 1752 -1909 1753 -1891
rect 89 -2016 90 -1910
rect 1164 -2016 1165 -1910
rect 1353 -1911 1354 -1891
rect 1493 -2016 1494 -1910
rect 1633 -2016 1634 -1910
rect 1647 -1911 1648 -1891
rect 1752 -2016 1753 -1910
rect 1780 -1911 1781 -1891
rect 100 -1913 101 -1891
rect 446 -1913 447 -1891
rect 464 -1913 465 -1891
rect 877 -1913 878 -1891
rect 926 -1913 927 -1891
rect 996 -1913 997 -1891
rect 1003 -1913 1004 -1891
rect 1115 -2016 1116 -1912
rect 1139 -2016 1140 -1912
rect 1773 -2016 1774 -1912
rect 1780 -2016 1781 -1912
rect 1801 -1913 1802 -1891
rect 100 -2016 101 -1914
rect 1577 -2016 1578 -1914
rect 1801 -2016 1802 -1914
rect 1815 -1915 1816 -1891
rect 110 -1917 111 -1891
rect 436 -2016 437 -1916
rect 509 -2016 510 -1916
rect 1346 -2016 1347 -1916
rect 1381 -2016 1382 -1916
rect 1507 -1917 1508 -1891
rect 142 -1919 143 -1891
rect 1654 -2016 1655 -1918
rect 142 -2016 143 -1920
rect 1556 -1921 1557 -1891
rect 145 -2016 146 -1922
rect 310 -2016 311 -1922
rect 324 -2016 325 -1922
rect 394 -1923 395 -1891
rect 527 -1923 528 -1891
rect 1689 -1923 1690 -1891
rect 149 -2016 150 -1924
rect 208 -1925 209 -1891
rect 212 -1925 213 -1891
rect 443 -1925 444 -1891
rect 527 -2016 528 -1924
rect 674 -1925 675 -1891
rect 723 -1925 724 -1891
rect 947 -2016 948 -1924
rect 957 -1925 958 -1891
rect 1318 -1925 1319 -1891
rect 1409 -2016 1410 -1924
rect 1521 -1925 1522 -1891
rect 1626 -1925 1627 -1891
rect 1689 -2016 1690 -1924
rect 156 -2016 157 -1926
rect 184 -1927 185 -1891
rect 191 -1927 192 -1891
rect 268 -2016 269 -1926
rect 334 -2016 335 -1926
rect 443 -2016 444 -1926
rect 541 -1927 542 -1891
rect 611 -2016 612 -1926
rect 618 -1927 619 -1891
rect 926 -2016 927 -1926
rect 929 -1927 930 -1891
rect 1003 -2016 1004 -1926
rect 1027 -1927 1028 -1891
rect 1647 -2016 1648 -1926
rect 128 -1929 129 -1891
rect 184 -2016 185 -1928
rect 191 -2016 192 -1928
rect 415 -1929 416 -1891
rect 506 -1929 507 -1891
rect 541 -2016 542 -1928
rect 597 -1929 598 -1891
rect 779 -2016 780 -1928
rect 800 -1929 801 -1891
rect 975 -1929 976 -1891
rect 1031 -2016 1032 -1928
rect 1080 -1929 1081 -1891
rect 1143 -2016 1144 -1928
rect 1248 -1929 1249 -1891
rect 1318 -2016 1319 -1928
rect 1360 -1929 1361 -1891
rect 1374 -1929 1375 -1891
rect 1521 -2016 1522 -1928
rect 1626 -2016 1627 -1928
rect 1675 -1929 1676 -1891
rect 152 -2016 153 -1930
rect 415 -2016 416 -1930
rect 457 -1931 458 -1891
rect 597 -2016 598 -1930
rect 604 -1931 605 -1891
rect 604 -2016 605 -1930
rect 604 -1931 605 -1891
rect 604 -2016 605 -1930
rect 618 -2016 619 -1930
rect 639 -1931 640 -1891
rect 653 -1931 654 -1891
rect 1213 -1931 1214 -1891
rect 1248 -2016 1249 -1930
rect 1262 -1931 1263 -1891
rect 1360 -2016 1361 -1930
rect 1444 -1931 1445 -1891
rect 1675 -2016 1676 -1930
rect 1710 -1931 1711 -1891
rect 37 -1933 38 -1891
rect 457 -2016 458 -1932
rect 506 -2016 507 -1932
rect 1759 -2016 1760 -1932
rect 159 -1935 160 -1891
rect 863 -2016 864 -1934
rect 901 -2016 902 -1934
rect 1556 -2016 1557 -1934
rect 1710 -2016 1711 -1934
rect 1745 -1935 1746 -1891
rect 163 -1937 164 -1891
rect 247 -1937 248 -1891
rect 254 -1937 255 -1891
rect 1048 -1937 1049 -1891
rect 1059 -1937 1060 -1891
rect 1353 -2016 1354 -1936
rect 1374 -2016 1375 -1936
rect 1395 -1937 1396 -1891
rect 1423 -1937 1424 -1891
rect 1444 -2016 1445 -1936
rect 163 -2016 164 -1938
rect 341 -1939 342 -1891
rect 345 -2016 346 -1938
rect 429 -1939 430 -1891
rect 632 -1939 633 -1891
rect 646 -2016 647 -1938
rect 653 -2016 654 -1938
rect 1041 -2016 1042 -1938
rect 1045 -1939 1046 -1891
rect 1297 -1939 1298 -1891
rect 1395 -2016 1396 -1938
rect 1500 -1939 1501 -1891
rect 93 -1941 94 -1891
rect 1500 -2016 1501 -1940
rect 93 -2016 94 -1942
rect 177 -1943 178 -1891
rect 198 -1943 199 -1891
rect 429 -2016 430 -1942
rect 632 -2016 633 -1942
rect 702 -1943 703 -1891
rect 737 -1943 738 -1891
rect 737 -2016 738 -1942
rect 737 -1943 738 -1891
rect 737 -2016 738 -1942
rect 751 -1943 752 -1891
rect 751 -2016 752 -1942
rect 751 -1943 752 -1891
rect 751 -2016 752 -1942
rect 772 -1943 773 -1891
rect 772 -2016 773 -1942
rect 772 -1943 773 -1891
rect 772 -2016 773 -1942
rect 793 -1943 794 -1891
rect 800 -2016 801 -1942
rect 807 -1943 808 -1891
rect 961 -1943 962 -1891
rect 968 -2016 969 -1942
rect 1332 -1943 1333 -1891
rect 1423 -2016 1424 -1942
rect 1514 -1943 1515 -1891
rect 103 -2016 104 -1944
rect 1332 -2016 1333 -1944
rect 1437 -1945 1438 -1891
rect 1451 -2016 1452 -1944
rect 1514 -2016 1515 -1944
rect 1535 -1945 1536 -1891
rect 170 -1947 171 -1891
rect 401 -2016 402 -1946
rect 460 -2016 461 -1946
rect 702 -2016 703 -1946
rect 807 -2016 808 -1946
rect 891 -1947 892 -1891
rect 933 -2016 934 -1946
rect 940 -1947 941 -1891
rect 975 -2016 976 -1946
rect 1339 -1947 1340 -1891
rect 1402 -1947 1403 -1891
rect 1437 -2016 1438 -1946
rect 1535 -2016 1536 -1946
rect 1563 -1947 1564 -1891
rect 110 -2016 111 -1948
rect 1402 -2016 1403 -1948
rect 1563 -2016 1564 -1948
rect 1570 -1949 1571 -1891
rect 170 -2016 171 -1950
rect 226 -1951 227 -1891
rect 247 -2016 248 -1950
rect 275 -1951 276 -1891
rect 373 -1951 374 -1891
rect 376 -1967 377 -1950
rect 380 -1951 381 -1891
rect 478 -2016 479 -1950
rect 639 -2016 640 -1950
rect 821 -1951 822 -1891
rect 824 -1951 825 -1891
rect 884 -1951 885 -1891
rect 891 -2016 892 -1950
rect 1458 -1951 1459 -1891
rect 114 -1953 115 -1891
rect 821 -2016 822 -1952
rect 835 -2016 836 -1952
rect 908 -1953 909 -1891
rect 1010 -1953 1011 -1891
rect 1045 -2016 1046 -1952
rect 1080 -2016 1081 -1952
rect 1108 -1953 1109 -1891
rect 1157 -1953 1158 -1891
rect 1185 -1953 1186 -1891
rect 1206 -1953 1207 -1891
rect 1339 -2016 1340 -1952
rect 1430 -1953 1431 -1891
rect 1458 -2016 1459 -1952
rect 114 -2016 115 -1954
rect 282 -1955 283 -1891
rect 373 -2016 374 -1954
rect 492 -1955 493 -1891
rect 667 -1955 668 -1891
rect 674 -2016 675 -1954
rect 719 -2016 720 -1954
rect 1108 -2016 1109 -1954
rect 1122 -1955 1123 -1891
rect 1430 -2016 1431 -1954
rect 131 -2016 132 -1956
rect 226 -2016 227 -1956
rect 254 -2016 255 -1956
rect 534 -1957 535 -1891
rect 667 -2016 668 -1956
rect 758 -1957 759 -1891
rect 786 -1957 787 -1891
rect 940 -2016 941 -1956
rect 989 -1957 990 -1891
rect 1010 -2016 1011 -1956
rect 1020 -1957 1021 -1891
rect 1059 -2016 1060 -1956
rect 1087 -1957 1088 -1891
rect 1122 -2016 1123 -1956
rect 1129 -1957 1130 -1891
rect 1157 -2016 1158 -1956
rect 1206 -2016 1207 -1956
rect 1241 -1957 1242 -1891
rect 1262 -2016 1263 -1956
rect 1486 -1957 1487 -1891
rect 177 -2016 178 -1958
rect 894 -2016 895 -1958
rect 989 -2016 990 -1958
rect 1584 -1959 1585 -1891
rect 180 -1961 181 -1891
rect 793 -2016 794 -1960
rect 814 -1961 815 -1891
rect 842 -2016 843 -1960
rect 877 -2016 878 -1960
rect 884 -2016 885 -1960
rect 1052 -1961 1053 -1891
rect 1185 -2016 1186 -1960
rect 1241 -2016 1242 -1960
rect 1255 -1961 1256 -1891
rect 1297 -2016 1298 -1960
rect 1325 -1961 1326 -1891
rect 1486 -2016 1487 -1960
rect 1619 -1961 1620 -1891
rect 180 -2016 181 -1962
rect 422 -1963 423 -1891
rect 492 -2016 493 -1962
rect 534 -2016 535 -1962
rect 555 -1963 556 -1891
rect 590 -1963 591 -1891
rect 786 -2016 787 -1962
rect 810 -1963 811 -1891
rect 1325 -2016 1326 -1962
rect 1528 -1963 1529 -1891
rect 1584 -2016 1585 -1962
rect 1619 -2016 1620 -1962
rect 1640 -1963 1641 -1891
rect 58 -1965 59 -1891
rect 555 -2016 556 -1964
rect 758 -2016 759 -1964
rect 1066 -1965 1067 -1891
rect 1073 -1965 1074 -1891
rect 1129 -2016 1130 -1964
rect 1220 -1965 1221 -1891
rect 1255 -2016 1256 -1964
rect 1311 -1965 1312 -1891
rect 1570 -2016 1571 -1964
rect 1640 -2016 1641 -1964
rect 1682 -1965 1683 -1891
rect 58 -2016 59 -1966
rect 709 -1967 710 -1891
rect 814 -2016 815 -1966
rect 856 -1967 857 -1891
rect 1052 -2016 1053 -1966
rect 1136 -1967 1137 -1891
rect 1192 -1967 1193 -1891
rect 1220 -2016 1221 -1966
rect 1269 -1967 1270 -1891
rect 1311 -2016 1312 -1966
rect 1384 -2016 1385 -1966
rect 1507 -2016 1508 -1966
rect 1528 -2016 1529 -1966
rect 1549 -1967 1550 -1891
rect 1682 -2016 1683 -1966
rect 1717 -1967 1718 -1891
rect 198 -2016 199 -1968
rect 761 -2016 762 -1968
rect 838 -1969 839 -1891
rect 1388 -1969 1389 -1891
rect 1542 -1969 1543 -1891
rect 1549 -2016 1550 -1968
rect 205 -2016 206 -1970
rect 289 -1971 290 -1891
rect 387 -1971 388 -1891
rect 464 -2016 465 -1970
rect 649 -1971 650 -1891
rect 1717 -2016 1718 -1970
rect 212 -2016 213 -1972
rect 1598 -1973 1599 -1891
rect 219 -1975 220 -1891
rect 1087 -2016 1088 -1974
rect 1178 -1975 1179 -1891
rect 1269 -2016 1270 -1974
rect 1388 -2016 1389 -1974
rect 1472 -1975 1473 -1891
rect 1598 -2016 1599 -1974
rect 1612 -1975 1613 -1891
rect 219 -2016 220 -1976
rect 380 -2016 381 -1976
rect 394 -2016 395 -1976
rect 716 -1977 717 -1891
rect 856 -2016 857 -1976
rect 870 -1977 871 -1891
rect 1017 -2016 1018 -1976
rect 1136 -2016 1137 -1976
rect 1178 -2016 1179 -1976
rect 1367 -1977 1368 -1891
rect 1465 -1977 1466 -1891
rect 1472 -2016 1473 -1976
rect 1612 -2016 1613 -1976
rect 1661 -1977 1662 -1891
rect 264 -1979 265 -1891
rect 289 -2016 290 -1978
rect 422 -2016 423 -1978
rect 730 -1979 731 -1891
rect 870 -2016 871 -1978
rect 936 -1979 937 -1891
rect 1038 -1979 1039 -1891
rect 1542 -2016 1543 -1978
rect 1661 -2016 1662 -1978
rect 1703 -1979 1704 -1891
rect 275 -2016 276 -1980
rect 359 -1981 360 -1891
rect 709 -2016 710 -1980
rect 898 -1981 899 -1891
rect 1038 -2016 1039 -1980
rect 1696 -1981 1697 -1891
rect 1703 -2016 1704 -1980
rect 1738 -1981 1739 -1891
rect 282 -2016 283 -1982
rect 471 -1983 472 -1891
rect 716 -2016 717 -1982
rect 849 -2016 850 -1982
rect 1066 -2016 1067 -1982
rect 1290 -1983 1291 -1891
rect 1293 -2016 1294 -1982
rect 1696 -2016 1697 -1982
rect 1738 -2016 1739 -1982
rect 1766 -1983 1767 -1891
rect 359 -2016 360 -1984
rect 688 -1985 689 -1891
rect 723 -2016 724 -1984
rect 898 -2016 899 -1984
rect 1073 -2016 1074 -1984
rect 1094 -1985 1095 -1891
rect 1192 -2016 1193 -1984
rect 1416 -2016 1417 -1984
rect 1465 -2016 1466 -1984
rect 1605 -1985 1606 -1891
rect 1766 -2016 1767 -1984
rect 1787 -1985 1788 -1891
rect 366 -1987 367 -1891
rect 471 -2016 472 -1986
rect 583 -1987 584 -1891
rect 1094 -2016 1095 -1986
rect 1304 -1987 1305 -1891
rect 1367 -2016 1368 -1986
rect 1591 -1987 1592 -1891
rect 1605 -2016 1606 -1986
rect 317 -1989 318 -1891
rect 366 -2016 367 -1988
rect 583 -2016 584 -1988
rect 625 -1989 626 -1891
rect 628 -2016 629 -1988
rect 1304 -2016 1305 -1988
rect 317 -2016 318 -1990
rect 408 -1991 409 -1891
rect 625 -2016 626 -1990
rect 695 -1991 696 -1891
rect 730 -2016 731 -1990
rect 1150 -1991 1151 -1891
rect 1160 -1991 1161 -1891
rect 1591 -2016 1592 -1990
rect 352 -1993 353 -1891
rect 408 -2016 409 -1992
rect 576 -1993 577 -1891
rect 695 -2016 696 -1992
rect 919 -2016 920 -1992
rect 1787 -2016 1788 -1992
rect 30 -1995 31 -1891
rect 576 -2016 577 -1994
rect 681 -1995 682 -1891
rect 688 -2016 689 -1994
rect 961 -2016 962 -1994
rect 1150 -2016 1151 -1994
rect 30 -2016 31 -1996
rect 331 -1997 332 -1891
rect 681 -2016 682 -1996
rect 765 -1997 766 -1891
rect 44 -1999 45 -1891
rect 331 -2016 332 -1998
rect 744 -1999 745 -1891
rect 765 -2016 766 -1998
rect 44 -2016 45 -2000
rect 530 -2001 531 -1891
rect 660 -2001 661 -1891
rect 744 -2016 745 -2000
rect 124 -2016 125 -2002
rect 352 -2016 353 -2002
rect 520 -2003 521 -1891
rect 660 -2016 661 -2002
rect 513 -2005 514 -1891
rect 520 -2016 521 -2004
rect 450 -2007 451 -1891
rect 513 -2016 514 -2006
rect 450 -2016 451 -2008
rect 569 -2009 570 -1891
rect 121 -2011 122 -1891
rect 569 -2016 570 -2010
rect 121 -2016 122 -2012
rect 1479 -2013 1480 -1891
rect 656 -2015 657 -1891
rect 1479 -2016 1480 -2014
rect 37 -2171 38 -2025
rect 625 -2026 626 -2024
rect 632 -2026 633 -2024
rect 632 -2171 633 -2025
rect 632 -2026 633 -2024
rect 632 -2171 633 -2025
rect 667 -2026 668 -2024
rect 670 -2046 671 -2025
rect 702 -2026 703 -2024
rect 957 -2026 958 -2024
rect 964 -2026 965 -2024
rect 1052 -2026 1053 -2024
rect 1062 -2171 1063 -2025
rect 1080 -2026 1081 -2024
rect 1139 -2026 1140 -2024
rect 1437 -2026 1438 -2024
rect 1479 -2026 1480 -2024
rect 1748 -2026 1749 -2024
rect 44 -2028 45 -2024
rect 712 -2171 713 -2027
rect 719 -2028 720 -2024
rect 926 -2028 927 -2024
rect 929 -2171 930 -2027
rect 1430 -2028 1431 -2024
rect 1591 -2028 1592 -2024
rect 1594 -2028 1595 -2024
rect 1713 -2171 1714 -2027
rect 1794 -2028 1795 -2024
rect 44 -2171 45 -2029
rect 180 -2030 181 -2024
rect 222 -2030 223 -2024
rect 247 -2030 248 -2024
rect 278 -2171 279 -2029
rect 1164 -2030 1165 -2024
rect 1195 -2030 1196 -2024
rect 1444 -2030 1445 -2024
rect 1591 -2171 1592 -2029
rect 1605 -2030 1606 -2024
rect 1745 -2030 1746 -2024
rect 1780 -2030 1781 -2024
rect 51 -2032 52 -2024
rect 177 -2032 178 -2024
rect 229 -2171 230 -2031
rect 1199 -2032 1200 -2024
rect 1213 -2032 1214 -2024
rect 1682 -2032 1683 -2024
rect 51 -2171 52 -2033
rect 275 -2034 276 -2024
rect 296 -2034 297 -2024
rect 296 -2171 297 -2033
rect 296 -2034 297 -2024
rect 296 -2171 297 -2033
rect 331 -2034 332 -2024
rect 471 -2034 472 -2024
rect 516 -2171 517 -2033
rect 940 -2034 941 -2024
rect 954 -2034 955 -2024
rect 1339 -2034 1340 -2024
rect 1423 -2034 1424 -2024
rect 1437 -2171 1438 -2033
rect 1444 -2171 1445 -2033
rect 1521 -2034 1522 -2024
rect 1682 -2171 1683 -2033
rect 1710 -2034 1711 -2024
rect 61 -2171 62 -2035
rect 1094 -2036 1095 -2024
rect 1157 -2036 1158 -2024
rect 1479 -2171 1480 -2035
rect 72 -2038 73 -2024
rect 201 -2171 202 -2037
rect 240 -2038 241 -2024
rect 250 -2171 251 -2037
rect 331 -2171 332 -2037
rect 460 -2038 461 -2024
rect 464 -2038 465 -2024
rect 506 -2171 507 -2037
rect 520 -2038 521 -2024
rect 523 -2046 524 -2037
rect 555 -2038 556 -2024
rect 586 -2171 587 -2037
rect 590 -2171 591 -2037
rect 597 -2038 598 -2024
rect 614 -2171 615 -2037
rect 975 -2038 976 -2024
rect 996 -2038 997 -2024
rect 1339 -2171 1340 -2037
rect 1395 -2038 1396 -2024
rect 1423 -2171 1424 -2037
rect 1430 -2171 1431 -2037
rect 1514 -2038 1515 -2024
rect 72 -2171 73 -2039
rect 261 -2040 262 -2024
rect 338 -2040 339 -2024
rect 593 -2040 594 -2024
rect 667 -2171 668 -2039
rect 730 -2040 731 -2024
rect 744 -2040 745 -2024
rect 744 -2171 745 -2039
rect 744 -2040 745 -2024
rect 744 -2171 745 -2039
rect 751 -2040 752 -2024
rect 894 -2040 895 -2024
rect 898 -2171 899 -2039
rect 1297 -2040 1298 -2024
rect 1314 -2171 1315 -2039
rect 1703 -2040 1704 -2024
rect 100 -2042 101 -2024
rect 422 -2042 423 -2024
rect 520 -2171 521 -2041
rect 558 -2171 559 -2041
rect 1521 -2171 1522 -2041
rect 1703 -2171 1704 -2041
rect 1724 -2042 1725 -2024
rect 103 -2044 104 -2024
rect 863 -2044 864 -2024
rect 877 -2044 878 -2024
rect 961 -2171 962 -2043
rect 996 -2171 997 -2043
rect 1178 -2044 1179 -2024
rect 1195 -2171 1196 -2043
rect 1668 -2044 1669 -2024
rect 1724 -2171 1725 -2043
rect 1787 -2044 1788 -2024
rect 103 -2171 104 -2045
rect 191 -2046 192 -2024
rect 205 -2046 206 -2024
rect 464 -2171 465 -2045
rect 702 -2171 703 -2045
rect 1451 -2046 1452 -2024
rect 1514 -2171 1515 -2045
rect 1570 -2046 1571 -2024
rect 1594 -2171 1595 -2045
rect 1605 -2171 1606 -2045
rect 1626 -2046 1627 -2024
rect 1668 -2171 1669 -2045
rect 110 -2171 111 -2047
rect 149 -2171 150 -2047
rect 177 -2171 178 -2047
rect 583 -2048 584 -2024
rect 751 -2171 752 -2047
rect 772 -2048 773 -2024
rect 786 -2048 787 -2024
rect 992 -2048 993 -2024
rect 999 -2048 1000 -2024
rect 1738 -2048 1739 -2024
rect 114 -2050 115 -2024
rect 597 -2171 598 -2049
rect 761 -2050 762 -2024
rect 835 -2050 836 -2024
rect 842 -2050 843 -2024
rect 842 -2171 843 -2049
rect 842 -2050 843 -2024
rect 842 -2171 843 -2049
rect 856 -2050 857 -2024
rect 863 -2171 864 -2049
rect 887 -2050 888 -2024
rect 1619 -2050 1620 -2024
rect 1626 -2171 1627 -2049
rect 1661 -2050 1662 -2024
rect 1738 -2171 1739 -2049
rect 1808 -2050 1809 -2024
rect 114 -2171 115 -2051
rect 653 -2052 654 -2024
rect 786 -2171 787 -2051
rect 884 -2052 885 -2024
rect 905 -2052 906 -2024
rect 954 -2171 955 -2051
rect 999 -2171 1000 -2051
rect 1115 -2052 1116 -2024
rect 1157 -2171 1158 -2051
rect 1171 -2052 1172 -2024
rect 1199 -2171 1200 -2051
rect 1332 -2052 1333 -2024
rect 1395 -2171 1396 -2051
rect 1409 -2052 1410 -2024
rect 1451 -2171 1452 -2051
rect 1458 -2052 1459 -2024
rect 1570 -2171 1571 -2051
rect 1577 -2052 1578 -2024
rect 1619 -2171 1620 -2051
rect 1640 -2052 1641 -2024
rect 1661 -2171 1662 -2051
rect 1759 -2052 1760 -2024
rect 121 -2054 122 -2024
rect 1500 -2054 1501 -2024
rect 1507 -2054 1508 -2024
rect 1640 -2171 1641 -2053
rect 121 -2171 122 -2055
rect 457 -2056 458 -2024
rect 572 -2056 573 -2024
rect 653 -2171 654 -2055
rect 695 -2056 696 -2024
rect 884 -2171 885 -2055
rect 912 -2056 913 -2024
rect 940 -2171 941 -2055
rect 1017 -2056 1018 -2024
rect 1038 -2171 1039 -2055
rect 1052 -2171 1053 -2055
rect 1101 -2056 1102 -2024
rect 1164 -2171 1165 -2055
rect 1248 -2056 1249 -2024
rect 1293 -2056 1294 -2024
rect 1367 -2056 1368 -2024
rect 1409 -2171 1410 -2055
rect 1416 -2056 1417 -2024
rect 1458 -2171 1459 -2055
rect 1528 -2056 1529 -2024
rect 1577 -2171 1578 -2055
rect 1598 -2056 1599 -2024
rect 124 -2058 125 -2024
rect 205 -2171 206 -2057
rect 219 -2058 220 -2024
rect 1297 -2171 1298 -2057
rect 1332 -2171 1333 -2057
rect 1388 -2058 1389 -2024
rect 1500 -2171 1501 -2057
rect 1696 -2058 1697 -2024
rect 124 -2171 125 -2059
rect 310 -2060 311 -2024
rect 338 -2171 339 -2059
rect 1108 -2060 1109 -2024
rect 1171 -2171 1172 -2059
rect 1241 -2060 1242 -2024
rect 1283 -2060 1284 -2024
rect 1367 -2171 1368 -2059
rect 1507 -2171 1508 -2059
rect 1563 -2060 1564 -2024
rect 1584 -2060 1585 -2024
rect 1598 -2171 1599 -2059
rect 1689 -2060 1690 -2024
rect 1696 -2171 1697 -2059
rect 131 -2062 132 -2024
rect 562 -2062 563 -2024
rect 569 -2062 570 -2024
rect 1248 -2171 1249 -2061
rect 1283 -2171 1284 -2061
rect 1318 -2062 1319 -2024
rect 1563 -2171 1564 -2061
rect 1612 -2062 1613 -2024
rect 1689 -2171 1690 -2061
rect 1717 -2062 1718 -2024
rect 131 -2171 132 -2063
rect 1654 -2064 1655 -2024
rect 135 -2066 136 -2024
rect 275 -2171 276 -2065
rect 359 -2066 360 -2024
rect 387 -2066 388 -2024
rect 394 -2066 395 -2024
rect 803 -2171 804 -2065
rect 817 -2171 818 -2065
rect 870 -2066 871 -2024
rect 873 -2171 874 -2065
rect 1528 -2171 1529 -2065
rect 1612 -2171 1613 -2065
rect 1647 -2066 1648 -2024
rect 1654 -2171 1655 -2065
rect 1752 -2066 1753 -2024
rect 30 -2068 31 -2024
rect 135 -2171 136 -2067
rect 142 -2068 143 -2024
rect 905 -2171 906 -2067
rect 912 -2171 913 -2067
rect 947 -2068 948 -2024
rect 968 -2068 969 -2024
rect 1108 -2171 1109 -2067
rect 1241 -2171 1242 -2067
rect 1276 -2068 1277 -2024
rect 1318 -2171 1319 -2067
rect 1381 -2068 1382 -2024
rect 1647 -2171 1648 -2067
rect 1731 -2068 1732 -2024
rect 30 -2171 31 -2069
rect 96 -2171 97 -2069
rect 142 -2171 143 -2069
rect 723 -2070 724 -2024
rect 793 -2171 794 -2069
rect 828 -2070 829 -2024
rect 831 -2171 832 -2069
rect 1255 -2070 1256 -2024
rect 1381 -2171 1382 -2069
rect 1542 -2070 1543 -2024
rect 1731 -2171 1732 -2069
rect 1801 -2070 1802 -2024
rect 145 -2072 146 -2024
rect 1003 -2072 1004 -2024
rect 1024 -2072 1025 -2024
rect 1115 -2171 1116 -2071
rect 1255 -2171 1256 -2071
rect 1311 -2072 1312 -2024
rect 184 -2074 185 -2024
rect 310 -2171 311 -2073
rect 317 -2074 318 -2024
rect 359 -2171 360 -2073
rect 366 -2074 367 -2024
rect 509 -2074 510 -2024
rect 548 -2074 549 -2024
rect 1584 -2171 1585 -2073
rect 184 -2171 185 -2075
rect 212 -2076 213 -2024
rect 233 -2076 234 -2024
rect 877 -2171 878 -2075
rect 922 -2076 923 -2024
rect 1185 -2076 1186 -2024
rect 1290 -2076 1291 -2024
rect 1542 -2171 1543 -2075
rect 65 -2078 66 -2024
rect 212 -2171 213 -2077
rect 240 -2171 241 -2077
rect 292 -2171 293 -2077
rect 317 -2171 318 -2077
rect 324 -2078 325 -2024
rect 366 -2171 367 -2077
rect 485 -2078 486 -2024
rect 541 -2078 542 -2024
rect 548 -2171 549 -2077
rect 628 -2078 629 -2024
rect 723 -2171 724 -2077
rect 796 -2078 797 -2024
rect 1213 -2171 1214 -2077
rect 65 -2171 66 -2079
rect 705 -2171 706 -2079
rect 709 -2080 710 -2024
rect 1017 -2171 1018 -2079
rect 1024 -2171 1025 -2079
rect 1143 -2080 1144 -2024
rect 1185 -2171 1186 -2079
rect 1269 -2080 1270 -2024
rect 86 -2082 87 -2024
rect 233 -2171 234 -2081
rect 247 -2171 248 -2081
rect 471 -2171 472 -2081
rect 541 -2171 542 -2081
rect 821 -2082 822 -2024
rect 835 -2171 836 -2081
rect 1027 -2171 1028 -2081
rect 1066 -2082 1067 -2024
rect 1066 -2171 1067 -2081
rect 1066 -2082 1067 -2024
rect 1066 -2171 1067 -2081
rect 1073 -2082 1074 -2024
rect 1136 -2171 1137 -2081
rect 1143 -2171 1144 -2081
rect 1304 -2082 1305 -2024
rect 86 -2171 87 -2083
rect 625 -2171 626 -2083
rect 695 -2171 696 -2083
rect 737 -2084 738 -2024
rect 821 -2171 822 -2083
rect 1472 -2084 1473 -2024
rect 191 -2171 192 -2085
rect 450 -2086 451 -2024
rect 457 -2171 458 -2085
rect 604 -2086 605 -2024
rect 681 -2086 682 -2024
rect 737 -2171 738 -2085
rect 856 -2171 857 -2085
rect 891 -2086 892 -2024
rect 919 -2086 920 -2024
rect 1290 -2171 1291 -2085
rect 1304 -2171 1305 -2085
rect 1360 -2086 1361 -2024
rect 1472 -2171 1473 -2085
rect 1493 -2086 1494 -2024
rect 93 -2088 94 -2024
rect 919 -2171 920 -2087
rect 933 -2088 934 -2024
rect 968 -2171 969 -2087
rect 989 -2088 990 -2024
rect 1276 -2171 1277 -2087
rect 1493 -2171 1494 -2087
rect 1556 -2088 1557 -2024
rect 93 -2171 94 -2089
rect 1633 -2090 1634 -2024
rect 163 -2092 164 -2024
rect 604 -2171 605 -2091
rect 660 -2092 661 -2024
rect 681 -2171 682 -2091
rect 807 -2092 808 -2024
rect 933 -2171 934 -2091
rect 947 -2171 948 -2091
rect 982 -2092 983 -2024
rect 1031 -2092 1032 -2024
rect 1073 -2171 1074 -2091
rect 1080 -2171 1081 -2091
rect 1129 -2092 1130 -2024
rect 1262 -2092 1263 -2024
rect 1360 -2171 1361 -2091
rect 1486 -2092 1487 -2024
rect 1556 -2171 1557 -2091
rect 1633 -2171 1634 -2091
rect 1675 -2092 1676 -2024
rect 163 -2171 164 -2093
rect 975 -2171 976 -2093
rect 978 -2171 979 -2093
rect 1262 -2171 1263 -2093
rect 1269 -2171 1270 -2093
rect 1325 -2094 1326 -2024
rect 1675 -2171 1676 -2093
rect 1766 -2094 1767 -2024
rect 198 -2096 199 -2024
rect 387 -2171 388 -2095
rect 394 -2171 395 -2095
rect 513 -2096 514 -2024
rect 555 -2171 556 -2095
rect 989 -2171 990 -2095
rect 1010 -2096 1011 -2024
rect 1031 -2171 1032 -2095
rect 1087 -2096 1088 -2024
rect 1416 -2171 1417 -2095
rect 198 -2171 199 -2097
rect 219 -2171 220 -2097
rect 254 -2098 255 -2024
rect 562 -2171 563 -2097
rect 583 -2171 584 -2097
rect 1486 -2171 1487 -2097
rect 254 -2171 255 -2099
rect 576 -2100 577 -2024
rect 807 -2171 808 -2099
rect 849 -2100 850 -2024
rect 891 -2171 892 -2099
rect 1132 -2171 1133 -2099
rect 1325 -2171 1326 -2099
rect 1353 -2100 1354 -2024
rect 156 -2102 157 -2024
rect 576 -2171 577 -2101
rect 716 -2102 717 -2024
rect 1353 -2171 1354 -2101
rect 58 -2104 59 -2024
rect 156 -2171 157 -2103
rect 268 -2104 269 -2024
rect 422 -2171 423 -2103
rect 429 -2104 430 -2024
rect 569 -2171 570 -2103
rect 716 -2171 717 -2103
rect 1192 -2171 1193 -2103
rect 226 -2106 227 -2024
rect 268 -2171 269 -2105
rect 282 -2106 283 -2024
rect 485 -2171 486 -2105
rect 814 -2106 815 -2024
rect 849 -2171 850 -2105
rect 982 -2171 983 -2105
rect 1059 -2106 1060 -2024
rect 1087 -2171 1088 -2105
rect 1227 -2106 1228 -2024
rect 226 -2171 227 -2107
rect 1178 -2171 1179 -2107
rect 1227 -2171 1228 -2107
rect 1710 -2171 1711 -2107
rect 282 -2171 283 -2109
rect 527 -2110 528 -2024
rect 1010 -2171 1011 -2109
rect 1374 -2110 1375 -2024
rect 289 -2112 290 -2024
rect 660 -2171 661 -2111
rect 1059 -2171 1060 -2111
rect 1388 -2171 1389 -2111
rect 170 -2114 171 -2024
rect 289 -2171 290 -2113
rect 324 -2171 325 -2113
rect 373 -2114 374 -2024
rect 380 -2114 381 -2024
rect 814 -2171 815 -2113
rect 1094 -2171 1095 -2113
rect 1122 -2114 1123 -2024
rect 1129 -2171 1130 -2113
rect 1773 -2114 1774 -2024
rect 170 -2171 171 -2115
rect 478 -2116 479 -2024
rect 527 -2171 528 -2115
rect 779 -2116 780 -2024
rect 1101 -2171 1102 -2115
rect 1150 -2116 1151 -2024
rect 1374 -2171 1375 -2115
rect 1465 -2116 1466 -2024
rect 107 -2118 108 -2024
rect 1465 -2171 1466 -2117
rect 107 -2171 108 -2119
rect 688 -2120 689 -2024
rect 758 -2120 759 -2024
rect 1150 -2171 1151 -2119
rect 345 -2122 346 -2024
rect 478 -2171 479 -2121
rect 499 -2122 500 -2024
rect 688 -2171 689 -2121
rect 765 -2122 766 -2024
rect 779 -2171 780 -2121
rect 345 -2171 346 -2123
rect 443 -2124 444 -2024
rect 499 -2171 500 -2123
rect 611 -2124 612 -2024
rect 765 -2171 766 -2123
rect 800 -2124 801 -2024
rect 303 -2126 304 -2024
rect 443 -2171 444 -2125
rect 492 -2126 493 -2024
rect 611 -2171 612 -2125
rect 303 -2171 304 -2127
rect 901 -2128 902 -2024
rect 352 -2130 353 -2024
rect 758 -2171 759 -2129
rect 352 -2171 353 -2131
rect 513 -2171 514 -2131
rect 373 -2171 374 -2133
rect 1346 -2134 1347 -2024
rect 128 -2136 129 -2024
rect 1346 -2171 1347 -2135
rect 128 -2171 129 -2137
rect 261 -2171 262 -2137
rect 380 -2171 381 -2137
rect 646 -2138 647 -2024
rect 401 -2140 402 -2024
rect 492 -2171 493 -2139
rect 646 -2171 647 -2139
rect 674 -2140 675 -2024
rect 79 -2142 80 -2024
rect 401 -2171 402 -2141
rect 408 -2142 409 -2024
rect 450 -2171 451 -2141
rect 674 -2171 675 -2141
rect 1125 -2171 1126 -2141
rect 79 -2171 80 -2143
rect 415 -2144 416 -2024
rect 418 -2171 419 -2143
rect 1003 -2171 1004 -2143
rect 408 -2171 409 -2145
rect 628 -2171 629 -2145
rect 429 -2171 430 -2147
rect 1311 -2171 1312 -2147
rect 436 -2150 437 -2024
rect 772 -2171 773 -2149
rect 436 -2171 437 -2151
rect 639 -2152 640 -2024
rect 618 -2154 619 -2024
rect 639 -2171 640 -2153
rect 618 -2171 619 -2155
rect 1045 -2156 1046 -2024
rect 1045 -2171 1046 -2157
rect 1220 -2158 1221 -2024
rect 1206 -2160 1207 -2024
rect 1220 -2171 1221 -2159
rect 1206 -2171 1207 -2161
rect 1234 -2162 1235 -2024
rect 1234 -2171 1235 -2163
rect 1402 -2164 1403 -2024
rect 1402 -2171 1403 -2165
rect 1535 -2166 1536 -2024
rect 1535 -2171 1536 -2167
rect 1549 -2168 1550 -2024
rect 152 -2170 153 -2024
rect 1549 -2171 1550 -2169
rect 51 -2181 52 -2179
rect 415 -2181 416 -2179
rect 418 -2181 419 -2179
rect 800 -2300 801 -2180
rect 803 -2181 804 -2179
rect 1689 -2181 1690 -2179
rect 1696 -2181 1697 -2179
rect 1710 -2181 1711 -2179
rect 58 -2300 59 -2182
rect 135 -2183 136 -2179
rect 145 -2300 146 -2182
rect 905 -2183 906 -2179
rect 940 -2183 941 -2179
rect 1059 -2183 1060 -2179
rect 1125 -2183 1126 -2179
rect 1423 -2183 1424 -2179
rect 1549 -2183 1550 -2179
rect 1549 -2300 1550 -2182
rect 1549 -2183 1550 -2179
rect 1549 -2300 1550 -2182
rect 1563 -2183 1564 -2179
rect 1563 -2300 1564 -2182
rect 1563 -2183 1564 -2179
rect 1563 -2300 1564 -2182
rect 1640 -2183 1641 -2179
rect 1717 -2183 1718 -2179
rect 72 -2185 73 -2179
rect 628 -2185 629 -2179
rect 660 -2185 661 -2179
rect 828 -2300 829 -2184
rect 866 -2300 867 -2184
rect 1339 -2185 1340 -2179
rect 1409 -2185 1410 -2179
rect 1412 -2185 1413 -2179
rect 1650 -2300 1651 -2184
rect 1668 -2185 1669 -2179
rect 1671 -2300 1672 -2184
rect 1738 -2185 1739 -2179
rect 93 -2187 94 -2179
rect 310 -2187 311 -2179
rect 317 -2187 318 -2179
rect 376 -2187 377 -2179
rect 380 -2187 381 -2179
rect 926 -2187 927 -2179
rect 943 -2300 944 -2186
rect 1087 -2187 1088 -2179
rect 1132 -2187 1133 -2179
rect 1682 -2187 1683 -2179
rect 1689 -2300 1690 -2186
rect 1724 -2187 1725 -2179
rect 93 -2300 94 -2188
rect 1202 -2300 1203 -2188
rect 1262 -2189 1263 -2179
rect 1682 -2300 1683 -2188
rect 1696 -2300 1697 -2188
rect 1731 -2189 1732 -2179
rect 100 -2191 101 -2179
rect 1041 -2300 1042 -2190
rect 1059 -2300 1060 -2190
rect 1066 -2191 1067 -2179
rect 1087 -2300 1088 -2190
rect 1122 -2191 1123 -2179
rect 1150 -2191 1151 -2179
rect 1339 -2300 1340 -2190
rect 1388 -2191 1389 -2179
rect 1668 -2300 1669 -2190
rect 61 -2193 62 -2179
rect 100 -2300 101 -2192
rect 107 -2300 108 -2192
rect 408 -2193 409 -2179
rect 492 -2193 493 -2179
rect 583 -2193 584 -2179
rect 586 -2193 587 -2179
rect 933 -2193 934 -2179
rect 975 -2193 976 -2179
rect 1367 -2193 1368 -2179
rect 1388 -2300 1389 -2192
rect 1444 -2193 1445 -2179
rect 110 -2195 111 -2179
rect 198 -2300 199 -2194
rect 201 -2195 202 -2179
rect 422 -2195 423 -2179
rect 499 -2195 500 -2179
rect 824 -2195 825 -2179
rect 873 -2195 874 -2179
rect 1297 -2195 1298 -2179
rect 1311 -2195 1312 -2179
rect 1507 -2195 1508 -2179
rect 72 -2300 73 -2196
rect 873 -2300 874 -2196
rect 877 -2197 878 -2179
rect 926 -2300 927 -2196
rect 933 -2300 934 -2196
rect 982 -2197 983 -2179
rect 999 -2197 1000 -2179
rect 1080 -2197 1081 -2179
rect 1150 -2300 1151 -2196
rect 1720 -2197 1721 -2179
rect 114 -2199 115 -2179
rect 422 -2300 423 -2198
rect 499 -2300 500 -2198
rect 506 -2199 507 -2179
rect 513 -2199 514 -2179
rect 1122 -2300 1123 -2198
rect 1174 -2300 1175 -2198
rect 1248 -2199 1249 -2179
rect 1262 -2300 1263 -2198
rect 1353 -2199 1354 -2179
rect 1409 -2300 1410 -2198
rect 1486 -2199 1487 -2179
rect 1507 -2300 1508 -2198
rect 1542 -2199 1543 -2179
rect 114 -2300 115 -2200
rect 614 -2201 615 -2179
rect 618 -2201 619 -2179
rect 670 -2300 671 -2200
rect 688 -2201 689 -2179
rect 870 -2300 871 -2200
rect 877 -2300 878 -2200
rect 1227 -2201 1228 -2179
rect 1248 -2300 1249 -2200
rect 1269 -2201 1270 -2179
rect 1311 -2300 1312 -2200
rect 1332 -2201 1333 -2179
rect 1353 -2300 1354 -2200
rect 1465 -2201 1466 -2179
rect 1542 -2300 1543 -2200
rect 1598 -2201 1599 -2179
rect 121 -2300 122 -2202
rect 457 -2203 458 -2179
rect 506 -2300 507 -2202
rect 576 -2203 577 -2179
rect 583 -2300 584 -2202
rect 590 -2203 591 -2179
rect 604 -2203 605 -2179
rect 838 -2300 839 -2202
rect 905 -2300 906 -2202
rect 961 -2203 962 -2179
rect 975 -2300 976 -2202
rect 1038 -2203 1039 -2179
rect 1066 -2300 1067 -2202
rect 1108 -2203 1109 -2179
rect 1227 -2300 1228 -2202
rect 1416 -2203 1417 -2179
rect 1444 -2300 1445 -2202
rect 1451 -2203 1452 -2179
rect 1598 -2300 1599 -2202
rect 1633 -2203 1634 -2179
rect 44 -2205 45 -2179
rect 457 -2300 458 -2204
rect 495 -2300 496 -2204
rect 590 -2300 591 -2204
rect 611 -2300 612 -2204
rect 632 -2205 633 -2179
rect 660 -2300 661 -2204
rect 912 -2205 913 -2179
rect 961 -2300 962 -2204
rect 1003 -2205 1004 -2179
rect 1020 -2300 1021 -2204
rect 1297 -2300 1298 -2204
rect 1318 -2205 1319 -2179
rect 1367 -2300 1368 -2204
rect 1374 -2205 1375 -2179
rect 1465 -2300 1466 -2204
rect 44 -2300 45 -2206
rect 96 -2207 97 -2179
rect 128 -2207 129 -2179
rect 135 -2300 136 -2206
rect 156 -2207 157 -2179
rect 408 -2300 409 -2206
rect 513 -2300 514 -2206
rect 520 -2207 521 -2179
rect 534 -2207 535 -2179
rect 558 -2207 559 -2179
rect 618 -2300 619 -2206
rect 646 -2207 647 -2179
rect 688 -2300 689 -2206
rect 807 -2207 808 -2179
rect 817 -2207 818 -2179
rect 1640 -2300 1641 -2206
rect 128 -2300 129 -2208
rect 653 -2209 654 -2179
rect 691 -2300 692 -2208
rect 723 -2209 724 -2179
rect 761 -2300 762 -2208
rect 1017 -2209 1018 -2179
rect 1027 -2209 1028 -2179
rect 1220 -2209 1221 -2179
rect 1314 -2209 1315 -2179
rect 1374 -2300 1375 -2208
rect 1381 -2209 1382 -2179
rect 1416 -2300 1417 -2208
rect 131 -2211 132 -2179
rect 149 -2211 150 -2179
rect 156 -2300 157 -2210
rect 464 -2211 465 -2179
rect 520 -2300 521 -2210
rect 569 -2211 570 -2179
rect 597 -2211 598 -2179
rect 646 -2300 647 -2210
rect 698 -2300 699 -2210
rect 786 -2211 787 -2179
rect 807 -2300 808 -2210
rect 863 -2211 864 -2179
rect 978 -2211 979 -2179
rect 1703 -2211 1704 -2179
rect 65 -2213 66 -2179
rect 863 -2300 864 -2212
rect 982 -2300 983 -2212
rect 1052 -2213 1053 -2179
rect 1062 -2213 1063 -2179
rect 1318 -2300 1319 -2212
rect 1332 -2300 1333 -2212
rect 1430 -2213 1431 -2179
rect 65 -2300 66 -2214
rect 282 -2215 283 -2179
rect 285 -2300 286 -2214
rect 1528 -2215 1529 -2179
rect 124 -2217 125 -2179
rect 1430 -2300 1431 -2216
rect 1528 -2300 1529 -2216
rect 1626 -2217 1627 -2179
rect 138 -2300 139 -2218
rect 653 -2300 654 -2218
rect 709 -2219 710 -2179
rect 1451 -2300 1452 -2218
rect 1626 -2300 1627 -2218
rect 1675 -2219 1676 -2179
rect 163 -2221 164 -2179
rect 247 -2300 248 -2220
rect 254 -2300 255 -2220
rect 338 -2221 339 -2179
rect 359 -2221 360 -2179
rect 380 -2300 381 -2220
rect 394 -2221 395 -2179
rect 579 -2300 580 -2220
rect 600 -2300 601 -2220
rect 1052 -2300 1053 -2220
rect 1080 -2300 1081 -2220
rect 1136 -2221 1137 -2179
rect 1381 -2300 1382 -2220
rect 1395 -2221 1396 -2179
rect 163 -2300 164 -2222
rect 737 -2223 738 -2179
rect 786 -2300 787 -2222
rect 849 -2223 850 -2179
rect 1003 -2300 1004 -2222
rect 1073 -2223 1074 -2179
rect 1108 -2300 1109 -2222
rect 1195 -2223 1196 -2179
rect 1395 -2300 1396 -2222
rect 1437 -2223 1438 -2179
rect 170 -2225 171 -2179
rect 415 -2300 416 -2224
rect 464 -2300 465 -2224
rect 667 -2225 668 -2179
rect 674 -2225 675 -2179
rect 849 -2300 850 -2224
rect 1017 -2300 1018 -2224
rect 1472 -2225 1473 -2179
rect 30 -2227 31 -2179
rect 170 -2300 171 -2226
rect 177 -2227 178 -2179
rect 642 -2300 643 -2226
rect 667 -2300 668 -2226
rect 919 -2227 920 -2179
rect 1024 -2227 1025 -2179
rect 1220 -2300 1221 -2226
rect 1437 -2300 1438 -2226
rect 1556 -2227 1557 -2179
rect 30 -2300 31 -2228
rect 208 -2300 209 -2228
rect 212 -2229 213 -2179
rect 289 -2300 290 -2228
rect 296 -2229 297 -2179
rect 299 -2263 300 -2228
rect 303 -2229 304 -2179
rect 702 -2229 703 -2179
rect 709 -2300 710 -2228
rect 898 -2229 899 -2179
rect 1027 -2300 1028 -2228
rect 1164 -2229 1165 -2179
rect 1556 -2300 1557 -2228
rect 1577 -2229 1578 -2179
rect 177 -2300 178 -2230
rect 695 -2231 696 -2179
rect 716 -2231 717 -2179
rect 919 -2300 920 -2230
rect 1073 -2300 1074 -2230
rect 1178 -2231 1179 -2179
rect 1577 -2300 1578 -2230
rect 1661 -2231 1662 -2179
rect 184 -2233 185 -2179
rect 184 -2300 185 -2232
rect 184 -2233 185 -2179
rect 184 -2300 185 -2232
rect 215 -2300 216 -2232
rect 1010 -2233 1011 -2179
rect 1115 -2233 1116 -2179
rect 1633 -2300 1634 -2232
rect 219 -2235 220 -2179
rect 219 -2300 220 -2234
rect 219 -2235 220 -2179
rect 219 -2300 220 -2234
rect 226 -2235 227 -2179
rect 541 -2235 542 -2179
rect 555 -2235 556 -2179
rect 639 -2235 640 -2179
rect 681 -2235 682 -2179
rect 702 -2300 703 -2234
rect 737 -2300 738 -2234
rect 1024 -2300 1025 -2234
rect 1115 -2300 1116 -2234
rect 1157 -2235 1158 -2179
rect 1178 -2300 1179 -2234
rect 1290 -2235 1291 -2179
rect 1535 -2235 1536 -2179
rect 1661 -2300 1662 -2234
rect 226 -2300 227 -2236
rect 240 -2237 241 -2179
rect 261 -2237 262 -2179
rect 373 -2300 374 -2236
rect 394 -2300 395 -2236
rect 450 -2237 451 -2179
rect 509 -2300 510 -2236
rect 716 -2300 717 -2236
rect 821 -2237 822 -2179
rect 1423 -2300 1424 -2236
rect 229 -2239 230 -2179
rect 1472 -2300 1473 -2238
rect 233 -2241 234 -2179
rect 1136 -2300 1137 -2240
rect 1143 -2241 1144 -2179
rect 1164 -2300 1165 -2240
rect 1199 -2241 1200 -2179
rect 1290 -2300 1291 -2240
rect 233 -2300 234 -2242
rect 912 -2300 913 -2242
rect 989 -2243 990 -2179
rect 1157 -2300 1158 -2242
rect 1206 -2243 1207 -2179
rect 1535 -2300 1536 -2242
rect 240 -2300 241 -2244
rect 597 -2300 598 -2244
rect 625 -2245 626 -2179
rect 1479 -2245 1480 -2179
rect 261 -2300 262 -2246
rect 1192 -2247 1193 -2179
rect 1206 -2300 1207 -2246
rect 1241 -2247 1242 -2179
rect 1479 -2300 1480 -2246
rect 1493 -2247 1494 -2179
rect 268 -2249 269 -2179
rect 275 -2300 276 -2248
rect 282 -2300 283 -2248
rect 954 -2249 955 -2179
rect 989 -2300 990 -2248
rect 1094 -2249 1095 -2179
rect 1143 -2300 1144 -2248
rect 1185 -2249 1186 -2179
rect 1241 -2300 1242 -2248
rect 1276 -2249 1277 -2179
rect 1493 -2300 1494 -2248
rect 1570 -2249 1571 -2179
rect 268 -2300 269 -2250
rect 345 -2251 346 -2179
rect 359 -2300 360 -2250
rect 831 -2251 832 -2179
rect 898 -2300 899 -2250
rect 968 -2251 969 -2179
rect 996 -2251 997 -2179
rect 1185 -2300 1186 -2250
rect 1276 -2300 1277 -2250
rect 1458 -2251 1459 -2179
rect 1570 -2300 1571 -2250
rect 1591 -2251 1592 -2179
rect 79 -2253 80 -2179
rect 345 -2300 346 -2252
rect 401 -2253 402 -2179
rect 569 -2300 570 -2252
rect 628 -2300 629 -2252
rect 1269 -2300 1270 -2252
rect 1591 -2300 1592 -2252
rect 1612 -2253 1613 -2179
rect 79 -2300 80 -2254
rect 1521 -2255 1522 -2179
rect 1605 -2255 1606 -2179
rect 1612 -2300 1613 -2254
rect 103 -2257 104 -2179
rect 1458 -2300 1459 -2256
rect 1521 -2300 1522 -2256
rect 1584 -2257 1585 -2179
rect 1605 -2300 1606 -2256
rect 1647 -2257 1648 -2179
rect 250 -2259 251 -2179
rect 401 -2300 402 -2258
rect 471 -2259 472 -2179
rect 968 -2300 969 -2258
rect 996 -2300 997 -2258
rect 1101 -2259 1102 -2179
rect 1584 -2300 1585 -2258
rect 1619 -2259 1620 -2179
rect 1647 -2300 1648 -2258
rect 1675 -2300 1676 -2258
rect 296 -2300 297 -2260
rect 471 -2300 472 -2260
rect 772 -2261 773 -2179
rect 821 -2300 822 -2260
rect 856 -2261 857 -2179
rect 929 -2261 930 -2179
rect 1192 -2300 1193 -2260
rect 1619 -2300 1620 -2260
rect 1654 -2261 1655 -2179
rect 257 -2263 258 -2179
rect 772 -2300 773 -2262
rect 856 -2300 857 -2262
rect 947 -2263 948 -2179
rect 954 -2300 955 -2262
rect 1213 -2263 1214 -2179
rect 1412 -2300 1413 -2262
rect 1486 -2300 1487 -2262
rect 303 -2300 304 -2264
rect 443 -2265 444 -2179
rect 534 -2300 535 -2264
rect 730 -2265 731 -2179
rect 814 -2265 815 -2179
rect 947 -2300 948 -2264
rect 1010 -2300 1011 -2264
rect 1713 -2265 1714 -2179
rect 191 -2267 192 -2179
rect 443 -2300 444 -2266
rect 541 -2300 542 -2266
rect 842 -2267 843 -2179
rect 1094 -2300 1095 -2266
rect 1171 -2267 1172 -2179
rect 1213 -2300 1214 -2266
rect 1255 -2267 1256 -2179
rect 149 -2300 150 -2268
rect 191 -2300 192 -2268
rect 310 -2300 311 -2268
rect 331 -2269 332 -2179
rect 338 -2300 339 -2268
rect 352 -2269 353 -2179
rect 548 -2269 549 -2179
rect 555 -2300 556 -2268
rect 632 -2300 633 -2268
rect 891 -2269 892 -2179
rect 1255 -2300 1256 -2268
rect 1346 -2269 1347 -2179
rect 86 -2271 87 -2179
rect 352 -2300 353 -2270
rect 681 -2300 682 -2270
rect 751 -2271 752 -2179
rect 758 -2271 759 -2179
rect 842 -2300 843 -2270
rect 1234 -2271 1235 -2179
rect 1346 -2300 1347 -2270
rect 86 -2300 87 -2272
rect 677 -2300 678 -2272
rect 705 -2300 706 -2272
rect 1101 -2300 1102 -2272
rect 1234 -2300 1235 -2272
rect 1325 -2273 1326 -2179
rect 152 -2300 153 -2274
rect 548 -2300 549 -2274
rect 730 -2300 731 -2274
rect 779 -2275 780 -2179
rect 793 -2275 794 -2179
rect 891 -2300 892 -2274
rect 1283 -2275 1284 -2179
rect 1325 -2300 1326 -2274
rect 205 -2277 206 -2179
rect 751 -2300 752 -2276
rect 814 -2300 815 -2276
rect 884 -2277 885 -2179
rect 1283 -2300 1284 -2276
rect 1304 -2277 1305 -2179
rect 317 -2300 318 -2278
rect 366 -2279 367 -2179
rect 527 -2279 528 -2179
rect 758 -2300 759 -2278
rect 884 -2300 885 -2278
rect 1045 -2279 1046 -2179
rect 1304 -2300 1305 -2278
rect 1360 -2279 1361 -2179
rect 142 -2281 143 -2179
rect 527 -2300 528 -2280
rect 604 -2300 605 -2280
rect 779 -2300 780 -2280
rect 1031 -2281 1032 -2179
rect 1045 -2300 1046 -2280
rect 1360 -2300 1361 -2280
rect 1402 -2281 1403 -2179
rect 142 -2300 143 -2282
rect 723 -2300 724 -2282
rect 744 -2283 745 -2179
rect 793 -2300 794 -2282
rect 1031 -2300 1032 -2282
rect 1129 -2283 1130 -2179
rect 1402 -2300 1403 -2282
rect 1500 -2283 1501 -2179
rect 205 -2300 206 -2284
rect 1129 -2300 1130 -2284
rect 1500 -2300 1501 -2284
rect 1514 -2285 1515 -2179
rect 324 -2287 325 -2179
rect 516 -2287 517 -2179
rect 744 -2300 745 -2286
rect 765 -2287 766 -2179
rect 324 -2300 325 -2288
rect 485 -2289 486 -2179
rect 765 -2300 766 -2288
rect 835 -2289 836 -2179
rect 331 -2300 332 -2290
rect 436 -2291 437 -2179
rect 485 -2300 486 -2290
rect 1038 -2300 1039 -2290
rect 366 -2300 367 -2292
rect 387 -2293 388 -2179
rect 436 -2300 437 -2292
rect 562 -2293 563 -2179
rect 835 -2300 836 -2292
rect 1514 -2300 1515 -2292
rect 37 -2295 38 -2179
rect 562 -2300 563 -2294
rect 387 -2300 388 -2296
rect 478 -2297 479 -2179
rect 450 -2300 451 -2298
rect 478 -2300 479 -2298
rect 30 -2310 31 -2308
rect 149 -2310 150 -2308
rect 205 -2421 206 -2309
rect 219 -2310 220 -2308
rect 254 -2310 255 -2308
rect 523 -2421 524 -2309
rect 548 -2310 549 -2308
rect 943 -2310 944 -2308
rect 971 -2421 972 -2309
rect 1094 -2310 1095 -2308
rect 1115 -2310 1116 -2308
rect 1115 -2421 1116 -2309
rect 1115 -2310 1116 -2308
rect 1115 -2421 1116 -2309
rect 1143 -2310 1144 -2308
rect 1143 -2421 1144 -2309
rect 1143 -2310 1144 -2308
rect 1143 -2421 1144 -2309
rect 1174 -2310 1175 -2308
rect 1493 -2310 1494 -2308
rect 1514 -2310 1515 -2308
rect 1514 -2421 1515 -2309
rect 1514 -2310 1515 -2308
rect 1514 -2421 1515 -2309
rect 1622 -2421 1623 -2309
rect 1696 -2310 1697 -2308
rect 51 -2421 52 -2311
rect 359 -2312 360 -2308
rect 387 -2312 388 -2308
rect 548 -2421 549 -2311
rect 576 -2312 577 -2308
rect 828 -2312 829 -2308
rect 835 -2312 836 -2308
rect 1451 -2312 1452 -2308
rect 1465 -2312 1466 -2308
rect 1465 -2421 1466 -2311
rect 1465 -2312 1466 -2308
rect 1465 -2421 1466 -2311
rect 1493 -2421 1494 -2311
rect 1542 -2312 1543 -2308
rect 1647 -2312 1648 -2308
rect 1689 -2312 1690 -2308
rect 65 -2314 66 -2308
rect 68 -2364 69 -2313
rect 79 -2314 80 -2308
rect 562 -2314 563 -2308
rect 597 -2421 598 -2313
rect 761 -2314 762 -2308
rect 779 -2314 780 -2308
rect 1346 -2314 1347 -2308
rect 1437 -2314 1438 -2308
rect 1437 -2421 1438 -2313
rect 1437 -2314 1438 -2308
rect 1437 -2421 1438 -2313
rect 1451 -2421 1452 -2313
rect 1654 -2314 1655 -2308
rect 65 -2421 66 -2315
rect 261 -2316 262 -2308
rect 285 -2421 286 -2315
rect 310 -2316 311 -2308
rect 317 -2316 318 -2308
rect 586 -2421 587 -2315
rect 625 -2316 626 -2308
rect 751 -2316 752 -2308
rect 821 -2316 822 -2308
rect 828 -2421 829 -2315
rect 859 -2421 860 -2315
rect 1430 -2316 1431 -2308
rect 1542 -2421 1543 -2315
rect 1584 -2316 1585 -2308
rect 79 -2421 80 -2317
rect 401 -2318 402 -2308
rect 415 -2318 416 -2308
rect 600 -2318 601 -2308
rect 635 -2421 636 -2317
rect 674 -2421 675 -2317
rect 677 -2318 678 -2308
rect 730 -2318 731 -2308
rect 740 -2421 741 -2317
rect 1633 -2318 1634 -2308
rect 128 -2320 129 -2308
rect 702 -2320 703 -2308
rect 705 -2320 706 -2308
rect 807 -2320 808 -2308
rect 866 -2320 867 -2308
rect 1248 -2320 1249 -2308
rect 1251 -2421 1252 -2319
rect 1325 -2320 1326 -2308
rect 1346 -2421 1347 -2319
rect 1374 -2320 1375 -2308
rect 1430 -2421 1431 -2319
rect 1458 -2320 1459 -2308
rect 1612 -2320 1613 -2308
rect 1633 -2421 1634 -2319
rect 114 -2322 115 -2308
rect 807 -2421 808 -2321
rect 873 -2322 874 -2308
rect 1304 -2322 1305 -2308
rect 1311 -2322 1312 -2308
rect 1311 -2421 1312 -2321
rect 1311 -2322 1312 -2308
rect 1311 -2421 1312 -2321
rect 1374 -2421 1375 -2321
rect 1395 -2322 1396 -2308
rect 1444 -2322 1445 -2308
rect 1458 -2421 1459 -2321
rect 1612 -2421 1613 -2321
rect 1640 -2322 1641 -2308
rect 114 -2421 115 -2323
rect 408 -2324 409 -2308
rect 450 -2324 451 -2308
rect 1136 -2324 1137 -2308
rect 1171 -2324 1172 -2308
rect 1654 -2421 1655 -2323
rect 135 -2421 136 -2325
rect 541 -2326 542 -2308
rect 562 -2421 563 -2325
rect 891 -2326 892 -2308
rect 912 -2326 913 -2308
rect 1290 -2326 1291 -2308
rect 1444 -2421 1445 -2325
rect 1472 -2326 1473 -2308
rect 149 -2421 150 -2327
rect 1066 -2328 1067 -2308
rect 1073 -2328 1074 -2308
rect 1136 -2421 1137 -2327
rect 1164 -2328 1165 -2308
rect 1171 -2421 1172 -2327
rect 1199 -2421 1200 -2327
rect 1535 -2328 1536 -2308
rect 208 -2330 209 -2308
rect 464 -2330 465 -2308
rect 492 -2330 493 -2308
rect 1041 -2330 1042 -2308
rect 1052 -2330 1053 -2308
rect 1094 -2421 1095 -2329
rect 1129 -2330 1130 -2308
rect 1584 -2421 1585 -2329
rect 215 -2332 216 -2308
rect 324 -2332 325 -2308
rect 359 -2421 360 -2331
rect 534 -2332 535 -2308
rect 541 -2421 542 -2331
rect 569 -2332 570 -2308
rect 579 -2332 580 -2308
rect 1052 -2421 1053 -2331
rect 1073 -2421 1074 -2331
rect 1080 -2332 1081 -2308
rect 1087 -2332 1088 -2308
rect 1087 -2421 1088 -2331
rect 1087 -2332 1088 -2308
rect 1087 -2421 1088 -2331
rect 1122 -2332 1123 -2308
rect 1129 -2421 1130 -2331
rect 1157 -2332 1158 -2308
rect 1164 -2421 1165 -2331
rect 1202 -2332 1203 -2308
rect 1381 -2332 1382 -2308
rect 1472 -2421 1473 -2331
rect 1507 -2332 1508 -2308
rect 1535 -2421 1536 -2331
rect 1591 -2332 1592 -2308
rect 86 -2334 87 -2308
rect 569 -2421 570 -2333
rect 590 -2334 591 -2308
rect 625 -2421 626 -2333
rect 639 -2334 640 -2308
rect 842 -2334 843 -2308
rect 891 -2421 892 -2333
rect 898 -2334 899 -2308
rect 912 -2421 913 -2333
rect 1293 -2421 1294 -2333
rect 1591 -2421 1592 -2333
rect 1605 -2334 1606 -2308
rect 72 -2336 73 -2308
rect 590 -2421 591 -2335
rect 639 -2421 640 -2335
rect 681 -2336 682 -2308
rect 684 -2421 685 -2335
rect 821 -2421 822 -2335
rect 842 -2421 843 -2335
rect 905 -2336 906 -2308
rect 915 -2336 916 -2308
rect 1416 -2336 1417 -2308
rect 1605 -2421 1606 -2335
rect 1671 -2336 1672 -2308
rect 72 -2421 73 -2337
rect 632 -2338 633 -2308
rect 667 -2421 668 -2337
rect 856 -2338 857 -2308
rect 919 -2338 920 -2308
rect 919 -2421 920 -2337
rect 919 -2338 920 -2308
rect 919 -2421 920 -2337
rect 989 -2338 990 -2308
rect 992 -2338 993 -2308
rect 1017 -2338 1018 -2308
rect 1108 -2338 1109 -2308
rect 1122 -2421 1123 -2337
rect 1577 -2338 1578 -2308
rect 86 -2421 87 -2339
rect 229 -2421 230 -2339
rect 233 -2340 234 -2308
rect 254 -2421 255 -2339
rect 261 -2421 262 -2339
rect 275 -2340 276 -2308
rect 289 -2340 290 -2308
rect 408 -2421 409 -2339
rect 436 -2340 437 -2308
rect 492 -2421 493 -2339
rect 495 -2340 496 -2308
rect 646 -2340 647 -2308
rect 681 -2421 682 -2339
rect 1157 -2421 1158 -2339
rect 1185 -2340 1186 -2308
rect 1507 -2421 1508 -2339
rect 117 -2421 118 -2341
rect 289 -2421 290 -2341
rect 296 -2342 297 -2308
rect 576 -2421 577 -2341
rect 632 -2421 633 -2341
rect 954 -2342 955 -2308
rect 975 -2342 976 -2308
rect 1108 -2421 1109 -2341
rect 1185 -2421 1186 -2341
rect 1367 -2342 1368 -2308
rect 142 -2344 143 -2308
rect 233 -2421 234 -2343
rect 247 -2344 248 -2308
rect 324 -2421 325 -2343
rect 373 -2344 374 -2308
rect 464 -2421 465 -2343
rect 478 -2344 479 -2308
rect 905 -2421 906 -2343
rect 975 -2421 976 -2343
rect 982 -2344 983 -2308
rect 989 -2421 990 -2343
rect 1003 -2344 1004 -2308
rect 1020 -2344 1021 -2308
rect 1059 -2344 1060 -2308
rect 1206 -2344 1207 -2308
rect 1244 -2344 1245 -2308
rect 1248 -2421 1249 -2343
rect 1626 -2344 1627 -2308
rect 142 -2421 143 -2345
rect 240 -2346 241 -2308
rect 247 -2421 248 -2345
rect 331 -2346 332 -2308
rect 373 -2421 374 -2345
rect 604 -2346 605 -2308
rect 688 -2346 689 -2308
rect 786 -2346 787 -2308
rect 849 -2346 850 -2308
rect 982 -2421 983 -2345
rect 1003 -2421 1004 -2345
rect 1031 -2346 1032 -2308
rect 1038 -2346 1039 -2308
rect 1388 -2346 1389 -2308
rect 1570 -2346 1571 -2308
rect 1626 -2421 1627 -2345
rect 170 -2348 171 -2308
rect 275 -2421 276 -2347
rect 282 -2348 283 -2308
rect 954 -2421 955 -2347
rect 996 -2348 997 -2308
rect 1031 -2421 1032 -2347
rect 1045 -2348 1046 -2308
rect 1080 -2421 1081 -2347
rect 1206 -2421 1207 -2347
rect 1363 -2421 1364 -2347
rect 1367 -2421 1368 -2347
rect 1500 -2348 1501 -2308
rect 170 -2421 171 -2349
rect 191 -2350 192 -2308
rect 219 -2421 220 -2349
rect 226 -2350 227 -2308
rect 240 -2421 241 -2349
rect 366 -2350 367 -2308
rect 380 -2350 381 -2308
rect 401 -2421 402 -2349
rect 422 -2350 423 -2308
rect 646 -2421 647 -2349
rect 691 -2350 692 -2308
rect 779 -2421 780 -2349
rect 786 -2421 787 -2349
rect 1668 -2350 1669 -2308
rect 184 -2352 185 -2308
rect 191 -2421 192 -2351
rect 226 -2421 227 -2351
rect 968 -2352 969 -2308
rect 1059 -2421 1060 -2351
rect 1227 -2352 1228 -2308
rect 1237 -2421 1238 -2351
rect 1486 -2352 1487 -2308
rect 184 -2421 185 -2353
rect 499 -2354 500 -2308
rect 499 -2421 500 -2353
rect 499 -2354 500 -2308
rect 499 -2421 500 -2353
rect 506 -2354 507 -2308
rect 702 -2421 703 -2353
rect 709 -2354 710 -2308
rect 1045 -2421 1046 -2353
rect 1150 -2354 1151 -2308
rect 1227 -2421 1228 -2353
rect 1241 -2354 1242 -2308
rect 1479 -2354 1480 -2308
rect 1486 -2421 1487 -2353
rect 1650 -2354 1651 -2308
rect 268 -2356 269 -2308
rect 415 -2421 416 -2355
rect 422 -2421 423 -2355
rect 457 -2356 458 -2308
rect 506 -2421 507 -2355
rect 555 -2356 556 -2308
rect 604 -2421 605 -2355
rect 611 -2356 612 -2308
rect 621 -2421 622 -2355
rect 1500 -2421 1501 -2355
rect 1650 -2421 1651 -2355
rect 1661 -2356 1662 -2308
rect 268 -2421 269 -2357
rect 835 -2421 836 -2357
rect 838 -2358 839 -2308
rect 1570 -2421 1571 -2357
rect 1661 -2421 1662 -2357
rect 1682 -2358 1683 -2308
rect 282 -2421 283 -2359
rect 1479 -2421 1480 -2359
rect 296 -2421 297 -2361
rect 338 -2362 339 -2308
rect 345 -2362 346 -2308
rect 688 -2421 689 -2361
rect 695 -2362 696 -2308
rect 877 -2362 878 -2308
rect 947 -2362 948 -2308
rect 1038 -2421 1039 -2361
rect 1150 -2421 1151 -2361
rect 1381 -2421 1382 -2361
rect 1388 -2421 1389 -2361
rect 1409 -2362 1410 -2308
rect 100 -2364 101 -2308
rect 695 -2421 696 -2363
rect 709 -2421 710 -2363
rect 793 -2364 794 -2308
rect 800 -2364 801 -2308
rect 877 -2421 878 -2363
rect 947 -2421 948 -2363
rect 961 -2364 962 -2308
rect 992 -2421 993 -2363
rect 996 -2421 997 -2363
rect 1220 -2364 1221 -2308
rect 1220 -2421 1221 -2363
rect 1220 -2364 1221 -2308
rect 1220 -2421 1221 -2363
rect 1241 -2421 1242 -2363
rect 1297 -2364 1298 -2308
rect 1318 -2364 1319 -2308
rect 1416 -2421 1417 -2363
rect 100 -2421 101 -2365
rect 814 -2366 815 -2308
rect 870 -2366 871 -2308
rect 1297 -2421 1298 -2365
rect 1318 -2421 1319 -2365
rect 1332 -2366 1333 -2308
rect 1339 -2366 1340 -2308
rect 1409 -2421 1410 -2365
rect 303 -2368 304 -2308
rect 303 -2421 304 -2367
rect 303 -2368 304 -2308
rect 303 -2421 304 -2367
rect 310 -2421 311 -2367
rect 471 -2368 472 -2308
rect 509 -2368 510 -2308
rect 513 -2368 514 -2308
rect 534 -2421 535 -2367
rect 929 -2421 930 -2367
rect 1269 -2368 1270 -2308
rect 1325 -2421 1326 -2367
rect 1332 -2421 1333 -2367
rect 1353 -2368 1354 -2308
rect 58 -2370 59 -2308
rect 513 -2421 514 -2369
rect 611 -2421 612 -2369
rect 793 -2421 794 -2369
rect 870 -2421 871 -2369
rect 1024 -2370 1025 -2308
rect 1255 -2370 1256 -2308
rect 1269 -2421 1270 -2369
rect 1283 -2370 1284 -2308
rect 1304 -2421 1305 -2369
rect 1339 -2421 1340 -2369
rect 1360 -2370 1361 -2308
rect 44 -2372 45 -2308
rect 58 -2421 59 -2371
rect 317 -2421 318 -2371
rect 670 -2372 671 -2308
rect 716 -2372 717 -2308
rect 800 -2421 801 -2371
rect 926 -2372 927 -2308
rect 961 -2421 962 -2371
rect 1234 -2372 1235 -2308
rect 1255 -2421 1256 -2371
rect 1262 -2372 1263 -2308
rect 1283 -2421 1284 -2371
rect 1290 -2421 1291 -2371
rect 1528 -2372 1529 -2308
rect 44 -2421 45 -2373
rect 782 -2374 783 -2308
rect 898 -2421 899 -2373
rect 926 -2421 927 -2373
rect 1017 -2421 1018 -2373
rect 1234 -2421 1235 -2373
rect 1353 -2421 1354 -2373
rect 1423 -2374 1424 -2308
rect 1528 -2421 1529 -2373
rect 1549 -2374 1550 -2308
rect 331 -2421 332 -2375
rect 649 -2421 650 -2375
rect 653 -2376 654 -2308
rect 1024 -2421 1025 -2375
rect 1192 -2376 1193 -2308
rect 1423 -2421 1424 -2375
rect 1549 -2421 1550 -2375
rect 1556 -2376 1557 -2308
rect 107 -2378 108 -2308
rect 653 -2421 654 -2377
rect 660 -2378 661 -2308
rect 814 -2421 815 -2377
rect 1178 -2378 1179 -2308
rect 1192 -2421 1193 -2377
rect 1213 -2378 1214 -2308
rect 1262 -2421 1263 -2377
rect 1402 -2378 1403 -2308
rect 1556 -2421 1557 -2377
rect 138 -2380 139 -2308
rect 1178 -2421 1179 -2379
rect 1213 -2421 1214 -2379
rect 1521 -2380 1522 -2308
rect 163 -2382 164 -2308
rect 660 -2421 661 -2381
rect 723 -2382 724 -2308
rect 1066 -2421 1067 -2381
rect 1276 -2382 1277 -2308
rect 1402 -2421 1403 -2381
rect 1521 -2421 1522 -2381
rect 1563 -2382 1564 -2308
rect 163 -2421 164 -2383
rect 429 -2384 430 -2308
rect 436 -2421 437 -2383
rect 520 -2384 521 -2308
rect 583 -2384 584 -2308
rect 716 -2421 717 -2383
rect 723 -2421 724 -2383
rect 1675 -2384 1676 -2308
rect 338 -2421 339 -2385
rect 352 -2386 353 -2308
rect 366 -2421 367 -2385
rect 527 -2386 528 -2308
rect 730 -2421 731 -2385
rect 884 -2386 885 -2308
rect 1202 -2421 1203 -2385
rect 1276 -2421 1277 -2385
rect 1563 -2421 1564 -2385
rect 1598 -2386 1599 -2308
rect 156 -2388 157 -2308
rect 352 -2421 353 -2387
rect 380 -2421 381 -2387
rect 1104 -2421 1105 -2387
rect 1598 -2421 1599 -2387
rect 1619 -2388 1620 -2308
rect 156 -2421 157 -2389
rect 733 -2421 734 -2389
rect 747 -2421 748 -2389
rect 1395 -2421 1396 -2389
rect 345 -2421 346 -2391
rect 583 -2421 584 -2391
rect 751 -2421 752 -2391
rect 863 -2392 864 -2308
rect 387 -2421 388 -2393
rect 394 -2394 395 -2308
rect 404 -2421 405 -2393
rect 429 -2421 430 -2393
rect 443 -2394 444 -2308
rect 478 -2421 479 -2393
rect 520 -2421 521 -2393
rect 555 -2421 556 -2393
rect 744 -2394 745 -2308
rect 863 -2421 864 -2393
rect 128 -2421 129 -2395
rect 744 -2421 745 -2395
rect 758 -2396 759 -2308
rect 884 -2421 885 -2395
rect 443 -2421 444 -2397
rect 940 -2398 941 -2308
rect 450 -2421 451 -2399
rect 1619 -2421 1620 -2399
rect 453 -2402 454 -2308
rect 737 -2402 738 -2308
rect 758 -2421 759 -2401
rect 765 -2402 766 -2308
rect 775 -2421 776 -2401
rect 1577 -2421 1578 -2401
rect 394 -2421 395 -2403
rect 737 -2421 738 -2403
rect 765 -2421 766 -2403
rect 772 -2404 773 -2308
rect 933 -2404 934 -2308
rect 940 -2421 941 -2403
rect 457 -2421 458 -2405
rect 1010 -2406 1011 -2308
rect 471 -2421 472 -2407
rect 618 -2408 619 -2308
rect 642 -2408 643 -2308
rect 933 -2421 934 -2407
rect 1010 -2421 1011 -2407
rect 1101 -2408 1102 -2308
rect 121 -2410 122 -2308
rect 618 -2421 619 -2409
rect 121 -2421 122 -2411
rect 212 -2412 213 -2308
rect 527 -2421 528 -2411
rect 772 -2421 773 -2411
rect 198 -2414 199 -2308
rect 212 -2421 213 -2413
rect 93 -2416 94 -2308
rect 198 -2421 199 -2415
rect 93 -2421 94 -2417
rect 177 -2418 178 -2308
rect 152 -2420 153 -2308
rect 177 -2421 178 -2419
rect 44 -2431 45 -2429
rect 530 -2540 531 -2430
rect 562 -2431 563 -2429
rect 1395 -2431 1396 -2429
rect 1444 -2431 1445 -2429
rect 1444 -2540 1445 -2430
rect 1444 -2431 1445 -2429
rect 1444 -2540 1445 -2430
rect 1500 -2431 1501 -2429
rect 1500 -2540 1501 -2430
rect 1500 -2431 1501 -2429
rect 1500 -2540 1501 -2430
rect 1615 -2540 1616 -2430
rect 1633 -2431 1634 -2429
rect 93 -2433 94 -2429
rect 117 -2433 118 -2429
rect 121 -2433 122 -2429
rect 775 -2433 776 -2429
rect 831 -2540 832 -2432
rect 1213 -2433 1214 -2429
rect 1234 -2540 1235 -2432
rect 1587 -2540 1588 -2432
rect 1622 -2433 1623 -2429
rect 1661 -2433 1662 -2429
rect 93 -2540 94 -2434
rect 443 -2435 444 -2429
rect 471 -2435 472 -2429
rect 614 -2435 615 -2429
rect 674 -2435 675 -2429
rect 740 -2435 741 -2429
rect 747 -2435 748 -2429
rect 1577 -2435 1578 -2429
rect 1626 -2435 1627 -2429
rect 1643 -2435 1644 -2429
rect 107 -2437 108 -2429
rect 1514 -2437 1515 -2429
rect 1577 -2540 1578 -2436
rect 1584 -2437 1585 -2429
rect 107 -2540 108 -2438
rect 110 -2439 111 -2429
rect 121 -2540 122 -2438
rect 723 -2439 724 -2429
rect 737 -2439 738 -2429
rect 1227 -2439 1228 -2429
rect 1248 -2540 1249 -2438
rect 1605 -2439 1606 -2429
rect 135 -2441 136 -2429
rect 646 -2441 647 -2429
rect 674 -2540 675 -2440
rect 1027 -2540 1028 -2440
rect 1066 -2441 1067 -2429
rect 1122 -2540 1123 -2440
rect 1185 -2441 1186 -2429
rect 1213 -2540 1214 -2440
rect 1251 -2441 1252 -2429
rect 1409 -2441 1410 -2429
rect 1549 -2441 1550 -2429
rect 1605 -2540 1606 -2440
rect 135 -2540 136 -2442
rect 457 -2443 458 -2429
rect 520 -2443 521 -2429
rect 660 -2443 661 -2429
rect 681 -2443 682 -2429
rect 863 -2443 864 -2429
rect 901 -2540 902 -2442
rect 975 -2443 976 -2429
rect 989 -2443 990 -2429
rect 1066 -2540 1067 -2442
rect 1104 -2443 1105 -2429
rect 1262 -2443 1263 -2429
rect 1290 -2443 1291 -2429
rect 1416 -2443 1417 -2429
rect 1549 -2540 1550 -2442
rect 1570 -2443 1571 -2429
rect 142 -2445 143 -2429
rect 481 -2540 482 -2444
rect 572 -2540 573 -2444
rect 716 -2445 717 -2429
rect 723 -2540 724 -2444
rect 1188 -2445 1189 -2429
rect 1199 -2445 1200 -2429
rect 1437 -2445 1438 -2429
rect 142 -2540 143 -2446
rect 387 -2447 388 -2429
rect 394 -2447 395 -2429
rect 471 -2540 472 -2446
rect 569 -2447 570 -2429
rect 716 -2540 717 -2446
rect 733 -2447 734 -2429
rect 1570 -2540 1571 -2446
rect 163 -2449 164 -2429
rect 810 -2540 811 -2448
rect 821 -2449 822 -2429
rect 989 -2540 990 -2448
rect 1013 -2540 1014 -2448
rect 1528 -2449 1529 -2429
rect 163 -2540 164 -2450
rect 390 -2540 391 -2450
rect 394 -2540 395 -2450
rect 632 -2451 633 -2429
rect 639 -2451 640 -2429
rect 646 -2540 647 -2450
rect 681 -2540 682 -2450
rect 684 -2451 685 -2429
rect 688 -2451 689 -2429
rect 803 -2540 804 -2450
rect 821 -2540 822 -2450
rect 1405 -2540 1406 -2450
rect 1493 -2451 1494 -2429
rect 1528 -2540 1529 -2450
rect 170 -2453 171 -2429
rect 257 -2540 258 -2452
rect 282 -2453 283 -2429
rect 772 -2453 773 -2429
rect 835 -2453 836 -2429
rect 1045 -2453 1046 -2429
rect 1115 -2453 1116 -2429
rect 1115 -2540 1116 -2452
rect 1115 -2453 1116 -2429
rect 1115 -2540 1116 -2452
rect 1164 -2453 1165 -2429
rect 1199 -2540 1200 -2452
rect 1220 -2453 1221 -2429
rect 1290 -2540 1291 -2452
rect 1332 -2453 1333 -2429
rect 1395 -2540 1396 -2452
rect 1486 -2453 1487 -2429
rect 1493 -2540 1494 -2452
rect 51 -2455 52 -2429
rect 170 -2540 171 -2454
rect 219 -2455 220 -2429
rect 226 -2540 227 -2454
rect 229 -2455 230 -2429
rect 1650 -2455 1651 -2429
rect 51 -2540 52 -2456
rect 401 -2457 402 -2429
rect 404 -2457 405 -2429
rect 429 -2457 430 -2429
rect 583 -2457 584 -2429
rect 1486 -2540 1487 -2456
rect 114 -2459 115 -2429
rect 219 -2540 220 -2458
rect 240 -2459 241 -2429
rect 429 -2540 430 -2458
rect 583 -2540 584 -2458
rect 709 -2459 710 -2429
rect 740 -2540 741 -2458
rect 842 -2459 843 -2429
rect 849 -2459 850 -2429
rect 1297 -2459 1298 -2429
rect 1339 -2459 1340 -2429
rect 1409 -2540 1410 -2458
rect 58 -2461 59 -2429
rect 114 -2540 115 -2460
rect 128 -2461 129 -2429
rect 835 -2540 836 -2460
rect 849 -2540 850 -2460
rect 877 -2461 878 -2429
rect 919 -2461 920 -2429
rect 1325 -2461 1326 -2429
rect 1346 -2461 1347 -2429
rect 1416 -2540 1417 -2460
rect 58 -2540 59 -2462
rect 285 -2540 286 -2462
rect 303 -2463 304 -2429
rect 730 -2463 731 -2429
rect 758 -2463 759 -2429
rect 772 -2540 773 -2462
rect 828 -2463 829 -2429
rect 842 -2540 843 -2462
rect 852 -2463 853 -2429
rect 1108 -2463 1109 -2429
rect 1192 -2463 1193 -2429
rect 1297 -2540 1298 -2462
rect 1318 -2463 1319 -2429
rect 1325 -2540 1326 -2462
rect 1353 -2463 1354 -2429
rect 1437 -2540 1438 -2462
rect 79 -2465 80 -2429
rect 758 -2540 759 -2464
rect 856 -2465 857 -2429
rect 1514 -2540 1515 -2464
rect 79 -2540 80 -2466
rect 247 -2467 248 -2429
rect 254 -2467 255 -2429
rect 282 -2540 283 -2466
rect 303 -2540 304 -2466
rect 1125 -2467 1126 -2429
rect 1143 -2467 1144 -2429
rect 1192 -2540 1193 -2466
rect 1206 -2467 1207 -2429
rect 1339 -2540 1340 -2466
rect 1360 -2467 1361 -2429
rect 1563 -2467 1564 -2429
rect 247 -2540 248 -2468
rect 478 -2469 479 -2429
rect 576 -2469 577 -2429
rect 730 -2540 731 -2468
rect 793 -2469 794 -2429
rect 856 -2540 857 -2468
rect 929 -2469 930 -2429
rect 1402 -2469 1403 -2429
rect 1563 -2540 1564 -2468
rect 1612 -2469 1613 -2429
rect 254 -2540 255 -2470
rect 859 -2471 860 -2429
rect 933 -2471 934 -2429
rect 1108 -2540 1109 -2470
rect 1171 -2471 1172 -2429
rect 1360 -2540 1361 -2470
rect 1374 -2471 1375 -2429
rect 1381 -2471 1382 -2429
rect 1384 -2471 1385 -2429
rect 1591 -2471 1592 -2429
rect 338 -2473 339 -2429
rect 457 -2540 458 -2472
rect 523 -2473 524 -2429
rect 576 -2540 577 -2472
rect 586 -2473 587 -2429
rect 1227 -2540 1228 -2472
rect 1241 -2473 1242 -2429
rect 1346 -2540 1347 -2472
rect 324 -2475 325 -2429
rect 338 -2540 339 -2474
rect 359 -2475 360 -2429
rect 478 -2540 479 -2474
rect 590 -2475 591 -2429
rect 590 -2540 591 -2474
rect 590 -2475 591 -2429
rect 590 -2540 591 -2474
rect 600 -2540 601 -2474
rect 961 -2475 962 -2429
rect 1024 -2475 1025 -2429
rect 1101 -2540 1102 -2474
rect 1150 -2475 1151 -2429
rect 1171 -2540 1172 -2474
rect 1202 -2475 1203 -2429
rect 1241 -2540 1242 -2474
rect 1251 -2540 1252 -2474
rect 1262 -2540 1263 -2474
rect 1269 -2475 1270 -2429
rect 1318 -2540 1319 -2474
rect 233 -2477 234 -2429
rect 324 -2540 325 -2476
rect 359 -2540 360 -2476
rect 464 -2477 465 -2429
rect 604 -2477 605 -2429
rect 660 -2540 661 -2476
rect 667 -2477 668 -2429
rect 877 -2540 878 -2476
rect 905 -2477 906 -2429
rect 961 -2540 962 -2476
rect 1024 -2540 1025 -2476
rect 1507 -2477 1508 -2429
rect 233 -2540 234 -2478
rect 373 -2479 374 -2429
rect 380 -2479 381 -2429
rect 863 -2540 864 -2478
rect 898 -2479 899 -2429
rect 905 -2540 906 -2478
rect 940 -2479 941 -2429
rect 940 -2540 941 -2478
rect 940 -2479 941 -2429
rect 940 -2540 941 -2478
rect 947 -2479 948 -2429
rect 975 -2540 976 -2478
rect 1038 -2479 1039 -2429
rect 1185 -2540 1186 -2478
rect 1206 -2540 1207 -2478
rect 1640 -2479 1641 -2429
rect 296 -2481 297 -2429
rect 373 -2540 374 -2480
rect 380 -2540 381 -2480
rect 702 -2481 703 -2429
rect 709 -2540 710 -2480
rect 765 -2481 766 -2429
rect 793 -2540 794 -2480
rect 800 -2481 801 -2429
rect 828 -2540 829 -2480
rect 1381 -2540 1382 -2480
rect 1507 -2540 1508 -2480
rect 1535 -2481 1536 -2429
rect 1640 -2540 1641 -2480
rect 1654 -2481 1655 -2429
rect 173 -2540 174 -2482
rect 296 -2540 297 -2482
rect 366 -2483 367 -2429
rect 562 -2540 563 -2482
rect 618 -2483 619 -2429
rect 919 -2540 920 -2482
rect 947 -2540 948 -2482
rect 1094 -2483 1095 -2429
rect 1178 -2483 1179 -2429
rect 1269 -2540 1270 -2482
rect 1276 -2483 1277 -2429
rect 1591 -2540 1592 -2482
rect 366 -2540 367 -2484
rect 499 -2485 500 -2429
rect 618 -2540 619 -2484
rect 625 -2485 626 -2429
rect 639 -2540 640 -2484
rect 838 -2485 839 -2429
rect 891 -2485 892 -2429
rect 1276 -2540 1277 -2484
rect 1283 -2485 1284 -2429
rect 1332 -2540 1333 -2484
rect 1535 -2540 1536 -2484
rect 1556 -2485 1557 -2429
rect 401 -2540 402 -2486
rect 436 -2487 437 -2429
rect 464 -2540 465 -2486
rect 653 -2487 654 -2429
rect 695 -2487 696 -2429
rect 933 -2540 934 -2486
rect 996 -2487 997 -2429
rect 1038 -2540 1039 -2486
rect 1045 -2540 1046 -2486
rect 1087 -2487 1088 -2429
rect 1129 -2487 1130 -2429
rect 1178 -2540 1179 -2486
rect 1220 -2540 1221 -2486
rect 1237 -2487 1238 -2429
rect 1304 -2487 1305 -2429
rect 1353 -2540 1354 -2486
rect 1556 -2540 1557 -2486
rect 1598 -2487 1599 -2429
rect 128 -2540 129 -2488
rect 996 -2540 997 -2488
rect 1052 -2489 1053 -2429
rect 1150 -2540 1151 -2488
rect 1304 -2540 1305 -2488
rect 1311 -2489 1312 -2429
rect 1458 -2489 1459 -2429
rect 1598 -2540 1599 -2488
rect 408 -2491 409 -2429
rect 443 -2540 444 -2490
rect 485 -2491 486 -2429
rect 604 -2540 605 -2490
rect 621 -2491 622 -2429
rect 688 -2540 689 -2490
rect 702 -2540 703 -2490
rect 807 -2491 808 -2429
rect 870 -2491 871 -2429
rect 891 -2540 892 -2490
rect 926 -2491 927 -2429
rect 1094 -2540 1095 -2490
rect 1146 -2540 1147 -2490
rect 1458 -2540 1459 -2490
rect 65 -2493 66 -2429
rect 485 -2540 486 -2492
rect 499 -2540 500 -2492
rect 541 -2493 542 -2429
rect 569 -2540 570 -2492
rect 1129 -2540 1130 -2492
rect 1255 -2493 1256 -2429
rect 1311 -2540 1312 -2492
rect 65 -2540 66 -2494
rect 1619 -2495 1620 -2429
rect 310 -2497 311 -2429
rect 408 -2540 409 -2496
rect 436 -2540 437 -2496
rect 450 -2497 451 -2429
rect 513 -2497 514 -2429
rect 695 -2540 696 -2496
rect 737 -2540 738 -2496
rect 1612 -2540 1613 -2496
rect 198 -2499 199 -2429
rect 310 -2540 311 -2498
rect 352 -2499 353 -2429
rect 541 -2540 542 -2498
rect 611 -2499 612 -2429
rect 1255 -2540 1256 -2498
rect 89 -2540 90 -2500
rect 352 -2540 353 -2500
rect 450 -2540 451 -2500
rect 565 -2501 566 -2429
rect 625 -2540 626 -2500
rect 912 -2501 913 -2429
rect 1052 -2540 1053 -2500
rect 1080 -2501 1081 -2429
rect 198 -2540 199 -2502
rect 205 -2503 206 -2429
rect 492 -2503 493 -2429
rect 513 -2540 514 -2502
rect 527 -2503 528 -2429
rect 1283 -2540 1284 -2502
rect 205 -2540 206 -2504
rect 212 -2505 213 -2429
rect 345 -2505 346 -2429
rect 527 -2540 528 -2504
rect 548 -2505 549 -2429
rect 611 -2540 612 -2504
rect 649 -2505 650 -2429
rect 1374 -2540 1375 -2504
rect 212 -2540 213 -2506
rect 275 -2507 276 -2429
rect 289 -2507 290 -2429
rect 345 -2540 346 -2506
rect 492 -2540 493 -2506
rect 786 -2507 787 -2429
rect 800 -2540 801 -2506
rect 1451 -2507 1452 -2429
rect 240 -2540 241 -2508
rect 289 -2540 290 -2508
rect 548 -2540 549 -2508
rect 597 -2509 598 -2429
rect 653 -2540 654 -2508
rect 779 -2509 780 -2429
rect 807 -2540 808 -2508
rect 1542 -2509 1543 -2429
rect 275 -2540 276 -2510
rect 422 -2511 423 -2429
rect 506 -2511 507 -2429
rect 597 -2540 598 -2510
rect 744 -2511 745 -2429
rect 1087 -2540 1088 -2510
rect 1367 -2511 1368 -2429
rect 1451 -2540 1452 -2510
rect 1521 -2511 1522 -2429
rect 1542 -2540 1543 -2510
rect 86 -2513 87 -2429
rect 506 -2540 507 -2512
rect 565 -2540 566 -2512
rect 632 -2540 633 -2512
rect 765 -2540 766 -2512
rect 1647 -2513 1648 -2429
rect 86 -2540 87 -2514
rect 520 -2540 521 -2514
rect 779 -2540 780 -2514
rect 1363 -2515 1364 -2429
rect 1479 -2515 1480 -2429
rect 1521 -2540 1522 -2514
rect 156 -2517 157 -2429
rect 422 -2540 423 -2516
rect 814 -2517 815 -2429
rect 870 -2540 871 -2516
rect 884 -2517 885 -2429
rect 926 -2540 927 -2516
rect 1010 -2517 1011 -2429
rect 1080 -2540 1081 -2516
rect 1157 -2517 1158 -2429
rect 1367 -2540 1368 -2516
rect 1472 -2517 1473 -2429
rect 1479 -2540 1480 -2516
rect 100 -2519 101 -2429
rect 156 -2540 157 -2518
rect 268 -2519 269 -2429
rect 814 -2540 815 -2518
rect 884 -2540 885 -2518
rect 1003 -2519 1004 -2429
rect 1073 -2519 1074 -2429
rect 1164 -2540 1165 -2518
rect 1465 -2519 1466 -2429
rect 1472 -2540 1473 -2518
rect 100 -2540 101 -2520
rect 331 -2521 332 -2429
rect 534 -2521 535 -2429
rect 1010 -2540 1011 -2520
rect 1073 -2540 1074 -2520
rect 1136 -2521 1137 -2429
rect 1430 -2521 1431 -2429
rect 1465 -2540 1466 -2520
rect 72 -2523 73 -2429
rect 534 -2540 535 -2522
rect 786 -2540 787 -2522
rect 1157 -2540 1158 -2522
rect 1423 -2523 1424 -2429
rect 1430 -2540 1431 -2522
rect 72 -2540 73 -2524
rect 261 -2525 262 -2429
rect 331 -2540 332 -2524
rect 415 -2525 416 -2429
rect 912 -2540 913 -2524
rect 954 -2525 955 -2429
rect 968 -2525 969 -2429
rect 1003 -2540 1004 -2524
rect 1388 -2525 1389 -2429
rect 1423 -2540 1424 -2524
rect 149 -2527 150 -2429
rect 1136 -2540 1137 -2526
rect 149 -2540 150 -2528
rect 191 -2529 192 -2429
rect 261 -2540 262 -2528
rect 317 -2529 318 -2429
rect 555 -2529 556 -2429
rect 1388 -2540 1389 -2528
rect 184 -2531 185 -2429
rect 268 -2540 269 -2530
rect 278 -2540 279 -2530
rect 555 -2540 556 -2530
rect 751 -2531 752 -2429
rect 954 -2540 955 -2530
rect 968 -2540 969 -2530
rect 982 -2531 983 -2429
rect 177 -2533 178 -2429
rect 184 -2540 185 -2532
rect 191 -2540 192 -2532
rect 744 -2540 745 -2532
rect 982 -2540 983 -2532
rect 1017 -2533 1018 -2429
rect 177 -2540 178 -2534
rect 215 -2540 216 -2534
rect 317 -2540 318 -2534
rect 387 -2540 388 -2534
rect 1017 -2540 1018 -2534
rect 1059 -2535 1060 -2429
rect 1031 -2537 1032 -2429
rect 1059 -2540 1060 -2536
rect 971 -2539 972 -2429
rect 1031 -2540 1032 -2538
rect 44 -2669 45 -2549
rect 303 -2550 304 -2548
rect 387 -2669 388 -2549
rect 639 -2550 640 -2548
rect 656 -2669 657 -2549
rect 1549 -2550 1550 -2548
rect 1556 -2550 1557 -2548
rect 1559 -2556 1560 -2549
rect 1584 -2550 1585 -2548
rect 1605 -2550 1606 -2548
rect 1629 -2669 1630 -2549
rect 1640 -2550 1641 -2548
rect 72 -2552 73 -2548
rect 292 -2552 293 -2548
rect 303 -2669 304 -2551
rect 425 -2669 426 -2551
rect 429 -2552 430 -2548
rect 429 -2669 430 -2551
rect 429 -2552 430 -2548
rect 429 -2669 430 -2551
rect 457 -2552 458 -2548
rect 478 -2669 479 -2551
rect 527 -2669 528 -2551
rect 681 -2552 682 -2548
rect 730 -2552 731 -2548
rect 1465 -2552 1466 -2548
rect 1472 -2552 1473 -2548
rect 1549 -2669 1550 -2551
rect 1556 -2669 1557 -2551
rect 1612 -2552 1613 -2548
rect 72 -2669 73 -2553
rect 618 -2554 619 -2548
rect 625 -2554 626 -2548
rect 807 -2669 808 -2553
rect 849 -2554 850 -2548
rect 898 -2554 899 -2548
rect 950 -2669 951 -2553
rect 1479 -2554 1480 -2548
rect 1514 -2554 1515 -2548
rect 1584 -2669 1585 -2553
rect 1591 -2554 1592 -2548
rect 1619 -2669 1620 -2553
rect 86 -2556 87 -2548
rect 180 -2669 181 -2555
rect 212 -2556 213 -2548
rect 296 -2669 297 -2555
rect 352 -2556 353 -2548
rect 681 -2669 682 -2555
rect 737 -2556 738 -2548
rect 1486 -2556 1487 -2548
rect 1612 -2669 1613 -2555
rect 86 -2669 87 -2557
rect 646 -2558 647 -2548
rect 737 -2669 738 -2557
rect 901 -2558 902 -2548
rect 971 -2669 972 -2557
rect 1122 -2558 1123 -2548
rect 1143 -2558 1144 -2548
rect 1325 -2558 1326 -2548
rect 1405 -2558 1406 -2548
rect 1542 -2558 1543 -2548
rect 1598 -2558 1599 -2548
rect 1626 -2669 1627 -2557
rect 93 -2560 94 -2548
rect 212 -2669 213 -2559
rect 233 -2560 234 -2548
rect 667 -2560 668 -2548
rect 744 -2560 745 -2548
rect 1101 -2560 1102 -2548
rect 1136 -2560 1137 -2548
rect 1143 -2669 1144 -2559
rect 1188 -2669 1189 -2559
rect 1430 -2560 1431 -2548
rect 1444 -2560 1445 -2548
rect 1479 -2669 1480 -2559
rect 1507 -2560 1508 -2548
rect 1542 -2669 1543 -2559
rect 1577 -2560 1578 -2548
rect 1598 -2669 1599 -2559
rect 93 -2669 94 -2561
rect 530 -2562 531 -2548
rect 534 -2562 535 -2548
rect 747 -2562 748 -2548
rect 789 -2562 790 -2548
rect 1276 -2562 1277 -2548
rect 1304 -2562 1305 -2548
rect 1402 -2669 1403 -2561
rect 1409 -2562 1410 -2548
rect 1486 -2669 1487 -2561
rect 121 -2564 122 -2548
rect 831 -2564 832 -2548
rect 835 -2564 836 -2548
rect 849 -2669 850 -2563
rect 887 -2669 888 -2563
rect 1297 -2564 1298 -2548
rect 1304 -2669 1305 -2563
rect 1437 -2564 1438 -2548
rect 1458 -2564 1459 -2548
rect 1514 -2669 1515 -2563
rect 65 -2566 66 -2548
rect 121 -2669 122 -2565
rect 135 -2566 136 -2548
rect 828 -2566 829 -2548
rect 901 -2669 902 -2565
rect 1066 -2566 1067 -2548
rect 1073 -2566 1074 -2548
rect 1465 -2669 1466 -2565
rect 65 -2669 66 -2567
rect 100 -2568 101 -2548
rect 135 -2669 136 -2567
rect 177 -2568 178 -2548
rect 201 -2669 202 -2567
rect 1444 -2669 1445 -2567
rect 100 -2669 101 -2569
rect 107 -2570 108 -2548
rect 142 -2570 143 -2548
rect 415 -2570 416 -2548
rect 422 -2570 423 -2548
rect 646 -2669 647 -2569
rect 667 -2669 668 -2569
rect 716 -2570 717 -2548
rect 730 -2669 731 -2569
rect 744 -2669 745 -2569
rect 758 -2570 759 -2548
rect 835 -2669 836 -2569
rect 954 -2570 955 -2548
rect 1325 -2669 1326 -2569
rect 1388 -2570 1389 -2548
rect 1437 -2669 1438 -2569
rect 107 -2669 108 -2571
rect 131 -2669 132 -2571
rect 142 -2669 143 -2571
rect 205 -2572 206 -2548
rect 215 -2572 216 -2548
rect 422 -2669 423 -2571
rect 450 -2572 451 -2548
rect 1122 -2669 1123 -2571
rect 1129 -2572 1130 -2548
rect 1136 -2669 1137 -2571
rect 1234 -2572 1235 -2548
rect 1591 -2669 1592 -2571
rect 152 -2669 153 -2573
rect 1507 -2669 1508 -2573
rect 163 -2576 164 -2548
rect 236 -2669 237 -2575
rect 254 -2576 255 -2548
rect 961 -2576 962 -2548
rect 978 -2669 979 -2575
rect 1283 -2576 1284 -2548
rect 1346 -2576 1347 -2548
rect 1388 -2669 1389 -2575
rect 1409 -2669 1410 -2575
rect 1570 -2576 1571 -2548
rect 226 -2578 227 -2548
rect 254 -2669 255 -2577
rect 275 -2578 276 -2548
rect 758 -2669 759 -2577
rect 803 -2578 804 -2548
rect 1360 -2578 1361 -2548
rect 1423 -2578 1424 -2548
rect 1458 -2669 1459 -2577
rect 198 -2580 199 -2548
rect 226 -2669 227 -2579
rect 268 -2580 269 -2548
rect 275 -2669 276 -2579
rect 278 -2580 279 -2548
rect 688 -2580 689 -2548
rect 828 -2669 829 -2579
rect 877 -2580 878 -2548
rect 926 -2580 927 -2548
rect 954 -2669 955 -2579
rect 961 -2669 962 -2579
rect 1059 -2580 1060 -2548
rect 1066 -2669 1067 -2579
rect 1087 -2580 1088 -2548
rect 1090 -2669 1091 -2579
rect 1535 -2580 1536 -2548
rect 268 -2669 269 -2581
rect 376 -2669 377 -2581
rect 380 -2582 381 -2548
rect 534 -2669 535 -2581
rect 562 -2582 563 -2548
rect 590 -2582 591 -2548
rect 597 -2582 598 -2548
rect 1577 -2669 1578 -2581
rect 247 -2584 248 -2548
rect 590 -2669 591 -2583
rect 600 -2584 601 -2548
rect 1472 -2669 1473 -2583
rect 247 -2669 248 -2585
rect 310 -2586 311 -2548
rect 317 -2586 318 -2548
rect 352 -2669 353 -2585
rect 390 -2586 391 -2548
rect 408 -2586 409 -2548
rect 450 -2669 451 -2585
rect 957 -2669 958 -2585
rect 996 -2586 997 -2548
rect 1563 -2586 1564 -2548
rect 89 -2588 90 -2548
rect 1563 -2669 1564 -2587
rect 191 -2590 192 -2548
rect 310 -2669 311 -2589
rect 345 -2590 346 -2548
rect 380 -2669 381 -2589
rect 394 -2590 395 -2548
rect 415 -2669 416 -2589
rect 457 -2669 458 -2589
rect 485 -2590 486 -2548
rect 492 -2590 493 -2548
rect 618 -2669 619 -2589
rect 625 -2669 626 -2589
rect 709 -2590 710 -2548
rect 880 -2669 881 -2589
rect 996 -2669 997 -2589
rect 1017 -2590 1018 -2548
rect 1297 -2669 1298 -2589
rect 1318 -2590 1319 -2548
rect 1360 -2669 1361 -2589
rect 1374 -2590 1375 -2548
rect 1423 -2669 1424 -2589
rect 58 -2592 59 -2548
rect 191 -2669 192 -2591
rect 282 -2592 283 -2548
rect 443 -2592 444 -2548
rect 464 -2592 465 -2548
rect 562 -2669 563 -2591
rect 565 -2592 566 -2548
rect 1535 -2669 1536 -2591
rect 58 -2669 59 -2593
rect 324 -2594 325 -2548
rect 345 -2669 346 -2593
rect 373 -2594 374 -2548
rect 401 -2594 402 -2548
rect 408 -2669 409 -2593
rect 464 -2669 465 -2593
rect 821 -2594 822 -2548
rect 905 -2594 906 -2548
rect 1059 -2669 1060 -2593
rect 1073 -2669 1074 -2593
rect 1227 -2594 1228 -2548
rect 1251 -2594 1252 -2548
rect 1528 -2594 1529 -2548
rect 233 -2669 234 -2595
rect 324 -2669 325 -2595
rect 401 -2669 402 -2595
rect 541 -2596 542 -2548
rect 555 -2596 556 -2548
rect 709 -2669 710 -2595
rect 786 -2596 787 -2548
rect 1017 -2669 1018 -2595
rect 1024 -2669 1025 -2595
rect 1521 -2596 1522 -2548
rect 257 -2598 258 -2548
rect 443 -2669 444 -2597
rect 481 -2598 482 -2548
rect 492 -2669 493 -2597
rect 502 -2669 503 -2597
rect 597 -2669 598 -2597
rect 611 -2598 612 -2548
rect 639 -2669 640 -2597
rect 688 -2669 689 -2597
rect 814 -2598 815 -2548
rect 821 -2669 822 -2597
rect 891 -2598 892 -2548
rect 905 -2669 906 -2597
rect 975 -2598 976 -2548
rect 1027 -2669 1028 -2597
rect 1339 -2598 1340 -2548
rect 1493 -2598 1494 -2548
rect 1521 -2669 1522 -2597
rect 156 -2600 157 -2548
rect 611 -2669 612 -2599
rect 614 -2669 615 -2599
rect 1283 -2669 1284 -2599
rect 1339 -2669 1340 -2599
rect 1615 -2600 1616 -2548
rect 156 -2669 157 -2601
rect 205 -2669 206 -2601
rect 261 -2602 262 -2548
rect 282 -2669 283 -2601
rect 289 -2602 290 -2548
rect 317 -2669 318 -2601
rect 485 -2669 486 -2601
rect 674 -2602 675 -2548
rect 786 -2669 787 -2601
rect 793 -2602 794 -2548
rect 814 -2669 815 -2601
rect 842 -2602 843 -2548
rect 877 -2669 878 -2601
rect 891 -2669 892 -2601
rect 912 -2602 913 -2548
rect 926 -2669 927 -2601
rect 1038 -2602 1039 -2548
rect 1101 -2669 1102 -2601
rect 1129 -2669 1130 -2601
rect 1262 -2602 1263 -2548
rect 1269 -2602 1270 -2548
rect 1318 -2669 1319 -2601
rect 1416 -2602 1417 -2548
rect 1493 -2669 1494 -2601
rect 1500 -2602 1501 -2548
rect 1528 -2669 1529 -2601
rect 163 -2669 164 -2603
rect 975 -2669 976 -2603
rect 1038 -2669 1039 -2603
rect 1115 -2604 1116 -2548
rect 1178 -2604 1179 -2548
rect 1374 -2669 1375 -2603
rect 1451 -2604 1452 -2548
rect 1500 -2669 1501 -2603
rect 240 -2606 241 -2548
rect 842 -2669 843 -2605
rect 912 -2669 913 -2605
rect 933 -2606 934 -2548
rect 1045 -2606 1046 -2548
rect 1430 -2669 1431 -2605
rect 219 -2608 220 -2548
rect 240 -2669 241 -2607
rect 261 -2669 262 -2607
rect 604 -2608 605 -2548
rect 632 -2608 633 -2548
rect 632 -2669 633 -2607
rect 632 -2608 633 -2548
rect 632 -2669 633 -2607
rect 733 -2608 734 -2548
rect 1178 -2669 1179 -2607
rect 1220 -2608 1221 -2548
rect 1262 -2669 1263 -2607
rect 1269 -2669 1270 -2607
rect 1636 -2669 1637 -2607
rect 219 -2669 220 -2609
rect 264 -2669 265 -2609
rect 289 -2669 290 -2609
rect 338 -2610 339 -2548
rect 520 -2610 521 -2548
rect 674 -2669 675 -2609
rect 733 -2669 734 -2609
rect 1241 -2610 1242 -2548
rect 1255 -2610 1256 -2548
rect 1346 -2669 1347 -2609
rect 1367 -2610 1368 -2548
rect 1416 -2669 1417 -2609
rect 338 -2669 339 -2611
rect 499 -2612 500 -2548
rect 520 -2669 521 -2611
rect 544 -2612 545 -2548
rect 555 -2669 556 -2611
rect 569 -2612 570 -2548
rect 572 -2612 573 -2548
rect 660 -2612 661 -2548
rect 793 -2669 794 -2611
rect 1010 -2612 1011 -2548
rect 1052 -2612 1053 -2548
rect 1146 -2612 1147 -2548
rect 1171 -2612 1172 -2548
rect 1220 -2669 1221 -2611
rect 1227 -2669 1228 -2611
rect 1248 -2612 1249 -2548
rect 1276 -2669 1277 -2611
rect 1587 -2612 1588 -2548
rect 499 -2669 500 -2613
rect 541 -2669 542 -2613
rect 569 -2669 570 -2613
rect 723 -2614 724 -2548
rect 800 -2614 801 -2548
rect 1045 -2669 1046 -2613
rect 1087 -2669 1088 -2613
rect 1234 -2669 1235 -2613
rect 1241 -2669 1242 -2613
rect 1381 -2614 1382 -2548
rect 1395 -2614 1396 -2548
rect 1451 -2669 1452 -2613
rect 471 -2616 472 -2548
rect 723 -2669 724 -2615
rect 863 -2616 864 -2548
rect 1248 -2669 1249 -2615
rect 1332 -2616 1333 -2548
rect 1367 -2669 1368 -2615
rect 359 -2618 360 -2548
rect 471 -2669 472 -2617
rect 583 -2618 584 -2548
rect 754 -2618 755 -2548
rect 863 -2669 864 -2617
rect 870 -2618 871 -2548
rect 884 -2618 885 -2548
rect 933 -2669 934 -2617
rect 940 -2618 941 -2548
rect 1010 -2669 1011 -2617
rect 1031 -2618 1032 -2548
rect 1052 -2669 1053 -2617
rect 1108 -2618 1109 -2548
rect 1171 -2669 1172 -2617
rect 1213 -2618 1214 -2548
rect 1255 -2669 1256 -2617
rect 1290 -2618 1291 -2548
rect 1332 -2669 1333 -2617
rect 1353 -2618 1354 -2548
rect 1395 -2669 1396 -2617
rect 208 -2669 209 -2619
rect 1108 -2669 1109 -2619
rect 1115 -2669 1116 -2619
rect 1199 -2620 1200 -2548
rect 1311 -2620 1312 -2548
rect 1353 -2669 1354 -2619
rect 359 -2669 360 -2621
rect 418 -2622 419 -2548
rect 583 -2669 584 -2621
rect 653 -2622 654 -2548
rect 660 -2669 661 -2621
rect 947 -2622 948 -2548
rect 1031 -2669 1032 -2621
rect 1206 -2622 1207 -2548
rect 331 -2624 332 -2548
rect 653 -2669 654 -2623
rect 670 -2624 671 -2548
rect 1381 -2669 1382 -2623
rect 79 -2626 80 -2548
rect 331 -2669 332 -2625
rect 604 -2669 605 -2625
rect 702 -2626 703 -2548
rect 740 -2626 741 -2548
rect 1206 -2669 1207 -2625
rect 79 -2669 80 -2627
rect 128 -2628 129 -2548
rect 702 -2669 703 -2627
rect 989 -2628 990 -2548
rect 1080 -2628 1081 -2548
rect 1213 -2669 1214 -2627
rect 803 -2669 804 -2629
rect 1290 -2669 1291 -2629
rect 810 -2632 811 -2548
rect 947 -2669 948 -2631
rect 989 -2669 990 -2631
rect 1003 -2632 1004 -2548
rect 1164 -2632 1165 -2548
rect 1199 -2669 1200 -2631
rect 856 -2634 857 -2548
rect 870 -2669 871 -2633
rect 884 -2669 885 -2633
rect 1094 -2634 1095 -2548
rect 1157 -2634 1158 -2548
rect 1164 -2669 1165 -2633
rect 1192 -2634 1193 -2548
rect 1311 -2669 1312 -2633
rect 170 -2636 171 -2548
rect 1094 -2669 1095 -2635
rect 1150 -2636 1151 -2548
rect 1157 -2669 1158 -2635
rect 170 -2669 171 -2637
rect 184 -2638 185 -2548
rect 751 -2638 752 -2548
rect 1192 -2669 1193 -2637
rect 184 -2669 185 -2639
rect 719 -2669 720 -2639
rect 859 -2669 860 -2639
rect 1080 -2669 1081 -2639
rect 1150 -2669 1151 -2639
rect 1605 -2669 1606 -2639
rect 506 -2642 507 -2548
rect 751 -2669 752 -2641
rect 919 -2642 920 -2548
rect 940 -2669 941 -2641
rect 982 -2642 983 -2548
rect 1003 -2669 1004 -2641
rect 506 -2669 507 -2643
rect 548 -2644 549 -2548
rect 919 -2669 920 -2643
rect 1153 -2669 1154 -2643
rect 436 -2646 437 -2548
rect 548 -2669 549 -2645
rect 968 -2646 969 -2548
rect 982 -2669 983 -2645
rect 436 -2669 437 -2647
rect 513 -2648 514 -2548
rect 968 -2669 969 -2647
rect 1185 -2648 1186 -2548
rect 513 -2669 514 -2649
rect 576 -2650 577 -2548
rect 1185 -2669 1186 -2649
rect 1570 -2669 1571 -2649
rect 576 -2669 577 -2651
rect 765 -2652 766 -2548
rect 765 -2669 766 -2653
rect 772 -2654 773 -2548
rect 695 -2656 696 -2548
rect 772 -2669 773 -2655
rect 695 -2669 696 -2657
rect 779 -2658 780 -2548
rect 51 -2660 52 -2548
rect 779 -2669 780 -2659
rect 51 -2669 52 -2661
rect 149 -2662 150 -2548
rect 114 -2664 115 -2548
rect 149 -2669 150 -2663
rect 114 -2669 115 -2665
rect 366 -2666 367 -2548
rect 366 -2669 367 -2667
rect 898 -2669 899 -2667
rect 44 -2679 45 -2677
rect 747 -2782 748 -2678
rect 782 -2782 783 -2678
rect 1584 -2679 1585 -2677
rect 44 -2782 45 -2680
rect 394 -2681 395 -2677
rect 397 -2681 398 -2677
rect 429 -2681 430 -2677
rect 436 -2681 437 -2677
rect 499 -2681 500 -2677
rect 534 -2681 535 -2677
rect 646 -2782 647 -2680
rect 649 -2681 650 -2677
rect 772 -2681 773 -2677
rect 786 -2681 787 -2677
rect 884 -2681 885 -2677
rect 908 -2782 909 -2680
rect 1297 -2681 1298 -2677
rect 1524 -2782 1525 -2680
rect 1598 -2681 1599 -2677
rect 51 -2683 52 -2677
rect 201 -2683 202 -2677
rect 205 -2683 206 -2677
rect 345 -2683 346 -2677
rect 394 -2782 395 -2682
rect 1188 -2683 1189 -2677
rect 1262 -2683 1263 -2677
rect 1300 -2782 1301 -2682
rect 58 -2685 59 -2677
rect 236 -2685 237 -2677
rect 264 -2685 265 -2677
rect 1283 -2685 1284 -2677
rect 58 -2782 59 -2686
rect 128 -2687 129 -2677
rect 135 -2687 136 -2677
rect 177 -2687 178 -2677
rect 198 -2687 199 -2677
rect 310 -2687 311 -2677
rect 331 -2687 332 -2677
rect 429 -2782 430 -2686
rect 446 -2782 447 -2686
rect 1507 -2687 1508 -2677
rect 72 -2689 73 -2677
rect 677 -2782 678 -2688
rect 681 -2689 682 -2677
rect 772 -2782 773 -2688
rect 786 -2782 787 -2688
rect 1465 -2689 1466 -2677
rect 1507 -2782 1508 -2688
rect 1605 -2689 1606 -2677
rect 72 -2782 73 -2690
rect 170 -2691 171 -2677
rect 177 -2782 178 -2690
rect 443 -2691 444 -2677
rect 499 -2782 500 -2690
rect 793 -2691 794 -2677
rect 800 -2691 801 -2677
rect 1171 -2691 1172 -2677
rect 1185 -2691 1186 -2677
rect 1549 -2691 1550 -2677
rect 79 -2693 80 -2677
rect 373 -2693 374 -2677
rect 408 -2693 409 -2677
rect 422 -2693 423 -2677
rect 534 -2782 535 -2692
rect 807 -2693 808 -2677
rect 817 -2782 818 -2692
rect 1486 -2693 1487 -2677
rect 79 -2782 80 -2694
rect 765 -2695 766 -2677
rect 793 -2782 794 -2694
rect 814 -2695 815 -2677
rect 877 -2695 878 -2677
rect 1010 -2695 1011 -2677
rect 1024 -2695 1025 -2677
rect 1465 -2782 1466 -2694
rect 1486 -2782 1487 -2694
rect 1577 -2695 1578 -2677
rect 86 -2697 87 -2677
rect 565 -2782 566 -2696
rect 576 -2697 577 -2677
rect 716 -2782 717 -2696
rect 730 -2782 731 -2696
rect 1153 -2697 1154 -2677
rect 1185 -2782 1186 -2696
rect 1339 -2697 1340 -2677
rect 86 -2782 87 -2698
rect 100 -2699 101 -2677
rect 114 -2699 115 -2677
rect 331 -2782 332 -2698
rect 345 -2782 346 -2698
rect 352 -2699 353 -2677
rect 373 -2782 374 -2698
rect 415 -2699 416 -2677
rect 422 -2782 423 -2698
rect 541 -2699 542 -2677
rect 576 -2782 577 -2698
rect 695 -2699 696 -2677
rect 709 -2699 710 -2677
rect 733 -2699 734 -2677
rect 737 -2699 738 -2677
rect 898 -2699 899 -2677
rect 940 -2699 941 -2677
rect 950 -2699 951 -2677
rect 957 -2699 958 -2677
rect 1311 -2699 1312 -2677
rect 65 -2701 66 -2677
rect 114 -2782 115 -2700
rect 124 -2782 125 -2700
rect 198 -2782 199 -2700
rect 205 -2782 206 -2700
rect 240 -2701 241 -2677
rect 264 -2782 265 -2700
rect 296 -2701 297 -2677
rect 310 -2782 311 -2700
rect 611 -2701 612 -2677
rect 653 -2701 654 -2677
rect 800 -2782 801 -2700
rect 845 -2782 846 -2700
rect 898 -2782 899 -2700
rect 933 -2701 934 -2677
rect 940 -2782 941 -2700
rect 968 -2782 969 -2700
rect 996 -2701 997 -2677
rect 1010 -2782 1011 -2700
rect 1626 -2701 1627 -2677
rect 65 -2782 66 -2702
rect 152 -2703 153 -2677
rect 156 -2703 157 -2677
rect 618 -2703 619 -2677
rect 653 -2782 654 -2702
rect 1143 -2703 1144 -2677
rect 1150 -2703 1151 -2677
rect 1612 -2703 1613 -2677
rect 93 -2705 94 -2677
rect 159 -2782 160 -2704
rect 170 -2782 171 -2704
rect 450 -2705 451 -2677
rect 464 -2705 465 -2677
rect 541 -2782 542 -2704
rect 569 -2705 570 -2677
rect 618 -2782 619 -2704
rect 656 -2705 657 -2677
rect 1052 -2705 1053 -2677
rect 1073 -2705 1074 -2677
rect 1171 -2782 1172 -2704
rect 1241 -2705 1242 -2677
rect 1339 -2782 1340 -2704
rect 93 -2782 94 -2706
rect 247 -2707 248 -2677
rect 275 -2707 276 -2677
rect 275 -2782 276 -2706
rect 275 -2707 276 -2677
rect 275 -2782 276 -2706
rect 296 -2782 297 -2706
rect 471 -2707 472 -2677
rect 520 -2707 521 -2677
rect 877 -2782 878 -2706
rect 880 -2707 881 -2677
rect 1374 -2707 1375 -2677
rect 100 -2782 101 -2708
rect 208 -2709 209 -2677
rect 212 -2709 213 -2677
rect 247 -2782 248 -2708
rect 352 -2782 353 -2708
rect 401 -2709 402 -2677
rect 415 -2782 416 -2708
rect 555 -2709 556 -2677
rect 569 -2782 570 -2708
rect 590 -2709 591 -2677
rect 604 -2709 605 -2677
rect 737 -2782 738 -2708
rect 744 -2709 745 -2677
rect 761 -2782 762 -2708
rect 765 -2782 766 -2708
rect 821 -2709 822 -2677
rect 880 -2782 881 -2708
rect 1101 -2709 1102 -2677
rect 1150 -2782 1151 -2708
rect 1381 -2709 1382 -2677
rect 128 -2782 129 -2710
rect 436 -2782 437 -2710
rect 450 -2782 451 -2710
rect 506 -2711 507 -2677
rect 555 -2782 556 -2710
rect 723 -2711 724 -2677
rect 744 -2782 745 -2710
rect 1430 -2711 1431 -2677
rect 135 -2782 136 -2712
rect 639 -2713 640 -2677
rect 660 -2713 661 -2677
rect 1090 -2713 1091 -2677
rect 1101 -2782 1102 -2712
rect 1206 -2713 1207 -2677
rect 1241 -2782 1242 -2712
rect 1353 -2713 1354 -2677
rect 1381 -2782 1382 -2712
rect 1542 -2713 1543 -2677
rect 142 -2715 143 -2677
rect 261 -2782 262 -2714
rect 401 -2782 402 -2714
rect 492 -2715 493 -2677
rect 506 -2782 507 -2714
rect 667 -2715 668 -2677
rect 674 -2715 675 -2677
rect 814 -2782 815 -2714
rect 821 -2782 822 -2714
rect 849 -2715 850 -2677
rect 884 -2782 885 -2714
rect 947 -2715 948 -2677
rect 954 -2715 955 -2677
rect 1143 -2782 1144 -2714
rect 1188 -2782 1189 -2714
rect 1374 -2782 1375 -2714
rect 1430 -2782 1431 -2714
rect 1514 -2715 1515 -2677
rect 142 -2782 143 -2716
rect 289 -2717 290 -2677
rect 425 -2717 426 -2677
rect 604 -2782 605 -2716
rect 611 -2782 612 -2716
rect 919 -2717 920 -2677
rect 926 -2717 927 -2677
rect 1052 -2782 1053 -2716
rect 1087 -2782 1088 -2716
rect 1178 -2717 1179 -2677
rect 1262 -2782 1263 -2716
rect 1367 -2717 1368 -2677
rect 1514 -2782 1515 -2716
rect 1619 -2717 1620 -2677
rect 149 -2719 150 -2677
rect 856 -2719 857 -2677
rect 870 -2719 871 -2677
rect 919 -2782 920 -2718
rect 933 -2782 934 -2718
rect 982 -2719 983 -2677
rect 996 -2782 997 -2718
rect 1003 -2719 1004 -2677
rect 1024 -2782 1025 -2718
rect 1108 -2719 1109 -2677
rect 1129 -2719 1130 -2677
rect 1206 -2782 1207 -2718
rect 1283 -2782 1284 -2718
rect 1451 -2719 1452 -2677
rect 149 -2782 150 -2720
rect 268 -2721 269 -2677
rect 464 -2782 465 -2720
rect 597 -2721 598 -2677
rect 625 -2721 626 -2677
rect 723 -2782 724 -2720
rect 779 -2721 780 -2677
rect 1073 -2782 1074 -2720
rect 1108 -2782 1109 -2720
rect 1192 -2721 1193 -2677
rect 1311 -2782 1312 -2720
rect 1395 -2721 1396 -2677
rect 1451 -2782 1452 -2720
rect 1528 -2721 1529 -2677
rect 156 -2782 157 -2722
rect 1269 -2723 1270 -2677
rect 1353 -2782 1354 -2722
rect 1444 -2723 1445 -2677
rect 163 -2725 164 -2677
rect 268 -2782 269 -2724
rect 387 -2725 388 -2677
rect 597 -2782 598 -2724
rect 660 -2782 661 -2724
rect 1591 -2725 1592 -2677
rect 163 -2782 164 -2726
rect 219 -2727 220 -2677
rect 226 -2727 227 -2677
rect 240 -2782 241 -2726
rect 387 -2782 388 -2726
rect 548 -2727 549 -2677
rect 562 -2727 563 -2677
rect 639 -2782 640 -2726
rect 663 -2782 664 -2726
rect 870 -2782 871 -2726
rect 901 -2727 902 -2677
rect 1269 -2782 1270 -2726
rect 1367 -2782 1368 -2726
rect 1458 -2727 1459 -2677
rect 138 -2782 139 -2728
rect 1458 -2782 1459 -2728
rect 215 -2782 216 -2730
rect 254 -2731 255 -2677
rect 408 -2782 409 -2730
rect 562 -2782 563 -2730
rect 681 -2782 682 -2730
rect 751 -2731 752 -2677
rect 849 -2782 850 -2730
rect 989 -2731 990 -2677
rect 1115 -2731 1116 -2677
rect 1129 -2782 1130 -2730
rect 1192 -2782 1193 -2730
rect 1423 -2731 1424 -2677
rect 1444 -2782 1445 -2730
rect 1629 -2731 1630 -2677
rect 219 -2782 220 -2732
rect 303 -2733 304 -2677
rect 366 -2733 367 -2677
rect 751 -2782 752 -2732
rect 856 -2782 857 -2732
rect 863 -2733 864 -2677
rect 905 -2733 906 -2677
rect 1178 -2782 1179 -2732
rect 1395 -2782 1396 -2732
rect 1472 -2733 1473 -2677
rect 226 -2782 227 -2734
rect 233 -2735 234 -2677
rect 254 -2782 255 -2734
rect 282 -2735 283 -2677
rect 303 -2782 304 -2734
rect 338 -2735 339 -2677
rect 471 -2782 472 -2734
rect 485 -2735 486 -2677
rect 492 -2782 493 -2734
rect 614 -2735 615 -2677
rect 691 -2782 692 -2734
rect 1080 -2735 1081 -2677
rect 1115 -2782 1116 -2734
rect 1227 -2735 1228 -2677
rect 1472 -2782 1473 -2734
rect 1556 -2735 1557 -2677
rect 212 -2782 213 -2736
rect 485 -2782 486 -2736
rect 527 -2737 528 -2677
rect 625 -2782 626 -2736
rect 695 -2782 696 -2736
rect 1094 -2737 1095 -2677
rect 1227 -2782 1228 -2736
rect 1325 -2737 1326 -2677
rect 324 -2739 325 -2677
rect 366 -2782 367 -2738
rect 478 -2739 479 -2677
rect 520 -2782 521 -2738
rect 527 -2782 528 -2738
rect 632 -2739 633 -2677
rect 702 -2739 703 -2677
rect 926 -2782 927 -2738
rect 954 -2782 955 -2738
rect 1136 -2739 1137 -2677
rect 1255 -2739 1256 -2677
rect 1325 -2782 1326 -2738
rect 292 -2782 293 -2740
rect 478 -2782 479 -2740
rect 548 -2782 549 -2740
rect 842 -2741 843 -2677
rect 859 -2741 860 -2677
rect 1423 -2782 1424 -2740
rect 324 -2782 325 -2742
rect 513 -2743 514 -2677
rect 583 -2743 584 -2677
rect 632 -2782 633 -2742
rect 702 -2782 703 -2742
rect 758 -2743 759 -2677
rect 842 -2782 843 -2742
rect 1059 -2743 1060 -2677
rect 1080 -2782 1081 -2742
rect 1157 -2743 1158 -2677
rect 1255 -2782 1256 -2742
rect 1360 -2743 1361 -2677
rect 338 -2782 339 -2744
rect 359 -2745 360 -2677
rect 457 -2745 458 -2677
rect 513 -2782 514 -2744
rect 583 -2782 584 -2744
rect 688 -2745 689 -2677
rect 709 -2782 710 -2744
rect 835 -2745 836 -2677
rect 863 -2782 864 -2744
rect 1157 -2782 1158 -2744
rect 1160 -2782 1161 -2744
rect 1360 -2782 1361 -2744
rect 184 -2747 185 -2677
rect 359 -2782 360 -2746
rect 380 -2747 381 -2677
rect 457 -2782 458 -2746
rect 758 -2782 759 -2746
rect 1346 -2747 1347 -2677
rect 184 -2782 185 -2748
rect 803 -2749 804 -2677
rect 828 -2749 829 -2677
rect 835 -2782 836 -2748
rect 891 -2749 892 -2677
rect 905 -2782 906 -2748
rect 961 -2749 962 -2677
rect 982 -2782 983 -2748
rect 989 -2782 990 -2748
rect 1017 -2749 1018 -2677
rect 1059 -2782 1060 -2748
rect 1220 -2749 1221 -2677
rect 1346 -2782 1347 -2748
rect 1437 -2749 1438 -2677
rect 121 -2751 122 -2677
rect 891 -2782 892 -2750
rect 971 -2751 972 -2677
rect 1038 -2751 1039 -2677
rect 1094 -2782 1095 -2750
rect 1164 -2751 1165 -2677
rect 1220 -2782 1221 -2750
rect 1636 -2751 1637 -2677
rect 121 -2782 122 -2752
rect 131 -2753 132 -2677
rect 317 -2753 318 -2677
rect 380 -2782 381 -2752
rect 779 -2782 780 -2752
rect 961 -2782 962 -2752
rect 975 -2753 976 -2677
rect 1045 -2753 1046 -2677
rect 1136 -2782 1137 -2752
rect 1234 -2753 1235 -2677
rect 1437 -2782 1438 -2752
rect 1521 -2753 1522 -2677
rect 107 -2755 108 -2677
rect 131 -2782 132 -2754
rect 191 -2755 192 -2677
rect 317 -2782 318 -2754
rect 828 -2782 829 -2754
rect 912 -2755 913 -2677
rect 947 -2782 948 -2754
rect 1521 -2782 1522 -2754
rect 107 -2782 108 -2756
rect 191 -2782 192 -2756
rect 289 -2782 290 -2756
rect 975 -2782 976 -2756
rect 978 -2757 979 -2677
rect 1493 -2757 1494 -2677
rect 667 -2782 668 -2758
rect 912 -2782 913 -2758
rect 1017 -2782 1018 -2758
rect 1031 -2759 1032 -2677
rect 1038 -2782 1039 -2758
rect 1122 -2759 1123 -2677
rect 1164 -2782 1165 -2758
rect 1248 -2759 1249 -2677
rect 1493 -2782 1494 -2758
rect 1570 -2759 1571 -2677
rect 1031 -2782 1032 -2760
rect 1066 -2761 1067 -2677
rect 1122 -2782 1123 -2760
rect 1276 -2761 1277 -2677
rect 1045 -2782 1046 -2762
rect 1213 -2763 1214 -2677
rect 1234 -2782 1235 -2762
rect 1332 -2763 1333 -2677
rect 1066 -2782 1067 -2764
rect 1199 -2765 1200 -2677
rect 1213 -2782 1214 -2764
rect 1318 -2765 1319 -2677
rect 1332 -2782 1333 -2764
rect 1409 -2765 1410 -2677
rect 1199 -2782 1200 -2766
rect 1290 -2767 1291 -2677
rect 1318 -2782 1319 -2766
rect 1416 -2767 1417 -2677
rect 887 -2769 888 -2677
rect 1416 -2782 1417 -2768
rect 1248 -2782 1249 -2770
rect 1633 -2771 1634 -2677
rect 1276 -2782 1277 -2772
rect 1388 -2773 1389 -2677
rect 1409 -2782 1410 -2772
rect 1500 -2773 1501 -2677
rect 1290 -2782 1291 -2774
rect 1535 -2775 1536 -2677
rect 1304 -2777 1305 -2677
rect 1388 -2782 1389 -2776
rect 1402 -2777 1403 -2677
rect 1500 -2782 1501 -2776
rect 674 -2782 675 -2778
rect 1304 -2782 1305 -2778
rect 1402 -2782 1403 -2778
rect 1479 -2779 1480 -2677
rect 1479 -2782 1480 -2780
rect 1563 -2781 1564 -2677
rect 58 -2792 59 -2790
rect 236 -2792 237 -2790
rect 247 -2792 248 -2790
rect 292 -2792 293 -2790
rect 296 -2792 297 -2790
rect 296 -2907 297 -2791
rect 296 -2792 297 -2790
rect 296 -2907 297 -2791
rect 303 -2792 304 -2790
rect 558 -2907 559 -2791
rect 593 -2792 594 -2790
rect 730 -2792 731 -2790
rect 747 -2792 748 -2790
rect 1143 -2792 1144 -2790
rect 1160 -2792 1161 -2790
rect 1500 -2792 1501 -2790
rect 65 -2794 66 -2790
rect 138 -2794 139 -2790
rect 149 -2794 150 -2790
rect 282 -2794 283 -2790
rect 285 -2907 286 -2793
rect 366 -2794 367 -2790
rect 373 -2794 374 -2790
rect 373 -2907 374 -2793
rect 373 -2794 374 -2790
rect 373 -2907 374 -2793
rect 380 -2794 381 -2790
rect 446 -2794 447 -2790
rect 499 -2794 500 -2790
rect 789 -2794 790 -2790
rect 810 -2794 811 -2790
rect 1479 -2794 1480 -2790
rect 86 -2796 87 -2790
rect 107 -2796 108 -2790
rect 110 -2796 111 -2790
rect 828 -2796 829 -2790
rect 845 -2796 846 -2790
rect 996 -2796 997 -2790
rect 1006 -2796 1007 -2790
rect 1325 -2796 1326 -2790
rect 86 -2907 87 -2797
rect 317 -2798 318 -2790
rect 324 -2798 325 -2790
rect 705 -2907 706 -2797
rect 730 -2907 731 -2797
rect 737 -2798 738 -2790
rect 772 -2798 773 -2790
rect 922 -2907 923 -2797
rect 996 -2907 997 -2797
rect 1136 -2798 1137 -2790
rect 1297 -2798 1298 -2790
rect 1381 -2798 1382 -2790
rect 93 -2800 94 -2790
rect 838 -2907 839 -2799
rect 866 -2907 867 -2799
rect 1486 -2800 1487 -2790
rect 93 -2907 94 -2801
rect 184 -2802 185 -2790
rect 198 -2802 199 -2790
rect 292 -2907 293 -2801
rect 310 -2802 311 -2790
rect 324 -2907 325 -2801
rect 331 -2802 332 -2790
rect 495 -2907 496 -2801
rect 499 -2907 500 -2801
rect 670 -2802 671 -2790
rect 688 -2802 689 -2790
rect 723 -2802 724 -2790
rect 737 -2907 738 -2801
rect 751 -2802 752 -2790
rect 772 -2907 773 -2801
rect 884 -2802 885 -2790
rect 898 -2802 899 -2790
rect 1185 -2802 1186 -2790
rect 1297 -2907 1298 -2801
rect 1395 -2802 1396 -2790
rect 107 -2907 108 -2803
rect 352 -2804 353 -2790
rect 366 -2907 367 -2803
rect 422 -2804 423 -2790
rect 429 -2804 430 -2790
rect 660 -2804 661 -2790
rect 688 -2907 689 -2803
rect 1150 -2804 1151 -2790
rect 1185 -2907 1186 -2803
rect 1255 -2804 1256 -2790
rect 1325 -2907 1326 -2803
rect 1437 -2804 1438 -2790
rect 100 -2806 101 -2790
rect 429 -2907 430 -2805
rect 443 -2806 444 -2790
rect 908 -2806 909 -2790
rect 912 -2806 913 -2790
rect 1157 -2806 1158 -2790
rect 1255 -2907 1256 -2805
rect 1311 -2806 1312 -2790
rect 1363 -2907 1364 -2805
rect 1395 -2907 1396 -2805
rect 114 -2808 115 -2790
rect 117 -2812 118 -2807
rect 121 -2808 122 -2790
rect 653 -2808 654 -2790
rect 723 -2907 724 -2807
rect 1010 -2808 1011 -2790
rect 1020 -2907 1021 -2807
rect 1507 -2808 1508 -2790
rect 114 -2907 115 -2809
rect 275 -2810 276 -2790
rect 310 -2907 311 -2809
rect 408 -2810 409 -2790
rect 443 -2907 444 -2809
rect 492 -2810 493 -2790
rect 506 -2810 507 -2790
rect 779 -2810 780 -2790
rect 828 -2907 829 -2809
rect 849 -2810 850 -2790
rect 898 -2907 899 -2809
rect 954 -2810 955 -2790
rect 1010 -2907 1011 -2809
rect 1164 -2810 1165 -2790
rect 1311 -2907 1312 -2809
rect 1430 -2810 1431 -2790
rect 275 -2907 276 -2811
rect 338 -2812 339 -2790
rect 422 -2907 423 -2811
rect 506 -2907 507 -2811
rect 625 -2812 626 -2790
rect 653 -2907 654 -2811
rect 1003 -2812 1004 -2790
rect 1097 -2907 1098 -2811
rect 1283 -2812 1284 -2790
rect 1381 -2907 1382 -2811
rect 1521 -2812 1522 -2790
rect 124 -2814 125 -2790
rect 331 -2907 332 -2813
rect 345 -2814 346 -2790
rect 590 -2814 591 -2790
rect 597 -2814 598 -2790
rect 807 -2814 808 -2790
rect 842 -2814 843 -2790
rect 884 -2907 885 -2813
rect 1003 -2907 1004 -2813
rect 1101 -2814 1102 -2790
rect 1129 -2814 1130 -2790
rect 1143 -2907 1144 -2813
rect 1150 -2907 1151 -2813
rect 1269 -2814 1270 -2790
rect 1283 -2907 1284 -2813
rect 1374 -2814 1375 -2790
rect 1430 -2907 1431 -2813
rect 1493 -2814 1494 -2790
rect 44 -2816 45 -2790
rect 124 -2907 125 -2815
rect 128 -2816 129 -2790
rect 513 -2816 514 -2790
rect 520 -2816 521 -2790
rect 562 -2816 563 -2790
rect 565 -2816 566 -2790
rect 1269 -2907 1270 -2815
rect 1374 -2907 1375 -2815
rect 1465 -2816 1466 -2790
rect 103 -2907 104 -2817
rect 128 -2907 129 -2817
rect 135 -2818 136 -2790
rect 660 -2907 661 -2817
rect 744 -2818 745 -2790
rect 1157 -2907 1158 -2817
rect 1164 -2907 1165 -2817
rect 1276 -2818 1277 -2790
rect 135 -2907 136 -2819
rect 569 -2820 570 -2790
rect 590 -2907 591 -2819
rect 604 -2820 605 -2790
rect 625 -2907 626 -2819
rect 947 -2820 948 -2790
rect 1101 -2907 1102 -2819
rect 1262 -2820 1263 -2790
rect 1276 -2907 1277 -2819
rect 1367 -2820 1368 -2790
rect 142 -2822 143 -2790
rect 338 -2907 339 -2821
rect 345 -2907 346 -2821
rect 401 -2822 402 -2790
rect 408 -2907 409 -2821
rect 485 -2822 486 -2790
rect 513 -2907 514 -2821
rect 709 -2822 710 -2790
rect 744 -2907 745 -2821
rect 1094 -2822 1095 -2790
rect 1129 -2907 1130 -2821
rect 1213 -2822 1214 -2790
rect 1262 -2907 1263 -2821
rect 1360 -2822 1361 -2790
rect 1367 -2907 1368 -2821
rect 1458 -2822 1459 -2790
rect 142 -2907 143 -2823
rect 149 -2907 150 -2823
rect 156 -2907 157 -2823
rect 555 -2824 556 -2790
rect 597 -2907 598 -2823
rect 681 -2824 682 -2790
rect 709 -2907 710 -2823
rect 880 -2824 881 -2790
rect 1136 -2907 1137 -2823
rect 1300 -2824 1301 -2790
rect 159 -2826 160 -2790
rect 856 -2826 857 -2790
rect 1213 -2907 1214 -2825
rect 1339 -2826 1340 -2790
rect 170 -2828 171 -2790
rect 303 -2907 304 -2827
rect 317 -2907 318 -2827
rect 1094 -2907 1095 -2827
rect 170 -2907 171 -2829
rect 250 -2907 251 -2829
rect 261 -2907 262 -2829
rect 541 -2830 542 -2790
rect 548 -2830 549 -2790
rect 667 -2830 668 -2790
rect 681 -2907 682 -2829
rect 947 -2907 948 -2829
rect 177 -2832 178 -2790
rect 478 -2907 479 -2831
rect 520 -2907 521 -2831
rect 765 -2832 766 -2790
rect 779 -2907 780 -2831
rect 891 -2832 892 -2790
rect 177 -2907 178 -2833
rect 450 -2834 451 -2790
rect 471 -2834 472 -2790
rect 485 -2907 486 -2833
rect 527 -2834 528 -2790
rect 562 -2907 563 -2833
rect 632 -2834 633 -2790
rect 667 -2907 668 -2833
rect 765 -2907 766 -2833
rect 863 -2834 864 -2790
rect 891 -2907 892 -2833
rect 989 -2834 990 -2790
rect 184 -2907 185 -2835
rect 205 -2836 206 -2790
rect 212 -2836 213 -2790
rect 1290 -2836 1291 -2790
rect 72 -2838 73 -2790
rect 205 -2907 206 -2837
rect 212 -2907 213 -2837
rect 282 -2907 283 -2837
rect 352 -2907 353 -2837
rect 457 -2838 458 -2790
rect 527 -2907 528 -2837
rect 957 -2907 958 -2837
rect 989 -2907 990 -2837
rect 1087 -2838 1088 -2790
rect 72 -2907 73 -2839
rect 163 -2840 164 -2790
rect 191 -2840 192 -2790
rect 198 -2907 199 -2839
rect 215 -2840 216 -2790
rect 677 -2840 678 -2790
rect 800 -2840 801 -2790
rect 807 -2907 808 -2839
rect 842 -2907 843 -2839
rect 982 -2840 983 -2790
rect 163 -2907 164 -2841
rect 268 -2842 269 -2790
rect 380 -2907 381 -2841
rect 642 -2907 643 -2841
rect 663 -2842 664 -2790
rect 1339 -2907 1340 -2841
rect 191 -2907 192 -2843
rect 208 -2907 209 -2843
rect 233 -2844 234 -2790
rect 751 -2907 752 -2843
rect 800 -2907 801 -2843
rect 940 -2844 941 -2790
rect 954 -2907 955 -2843
rect 1087 -2907 1088 -2843
rect 226 -2846 227 -2790
rect 233 -2907 234 -2845
rect 247 -2907 248 -2845
rect 695 -2846 696 -2790
rect 845 -2907 846 -2845
rect 940 -2907 941 -2845
rect 982 -2907 983 -2845
rect 1066 -2846 1067 -2790
rect 226 -2907 227 -2847
rect 618 -2848 619 -2790
rect 632 -2907 633 -2847
rect 1024 -2848 1025 -2790
rect 1066 -2907 1067 -2847
rect 1220 -2848 1221 -2790
rect 254 -2850 255 -2790
rect 268 -2907 269 -2849
rect 387 -2850 388 -2790
rect 814 -2850 815 -2790
rect 849 -2907 850 -2849
rect 1073 -2850 1074 -2790
rect 219 -2852 220 -2790
rect 387 -2907 388 -2851
rect 401 -2907 402 -2851
rect 464 -2852 465 -2790
rect 534 -2852 535 -2790
rect 824 -2907 825 -2851
rect 856 -2907 857 -2851
rect 961 -2852 962 -2790
rect 1073 -2907 1074 -2851
rect 1241 -2852 1242 -2790
rect 219 -2907 220 -2853
rect 817 -2854 818 -2790
rect 912 -2907 913 -2853
rect 1290 -2907 1291 -2853
rect 229 -2907 230 -2855
rect 464 -2907 465 -2855
rect 534 -2907 535 -2855
rect 702 -2856 703 -2790
rect 761 -2856 762 -2790
rect 1220 -2907 1221 -2855
rect 1241 -2907 1242 -2855
rect 1353 -2856 1354 -2790
rect 240 -2858 241 -2790
rect 254 -2907 255 -2857
rect 264 -2858 265 -2790
rect 359 -2858 360 -2790
rect 436 -2858 437 -2790
rect 471 -2907 472 -2857
rect 541 -2907 542 -2857
rect 646 -2858 647 -2790
rect 674 -2907 675 -2857
rect 702 -2907 703 -2857
rect 761 -2907 762 -2857
rect 1052 -2858 1053 -2790
rect 1353 -2907 1354 -2857
rect 1472 -2858 1473 -2790
rect 79 -2860 80 -2790
rect 436 -2907 437 -2859
rect 450 -2907 451 -2859
rect 576 -2860 577 -2790
rect 618 -2907 619 -2859
rect 639 -2860 640 -2790
rect 695 -2907 696 -2859
rect 793 -2860 794 -2790
rect 814 -2907 815 -2859
rect 919 -2860 920 -2790
rect 961 -2907 962 -2859
rect 1045 -2860 1046 -2790
rect 1052 -2907 1053 -2859
rect 1227 -2860 1228 -2790
rect 79 -2907 80 -2861
rect 278 -2907 279 -2861
rect 359 -2907 360 -2861
rect 415 -2862 416 -2790
rect 457 -2907 458 -2861
rect 915 -2907 916 -2861
rect 919 -2907 920 -2861
rect 1122 -2862 1123 -2790
rect 121 -2907 122 -2863
rect 646 -2907 647 -2863
rect 793 -2907 794 -2863
rect 835 -2864 836 -2790
rect 877 -2864 878 -2790
rect 1227 -2907 1228 -2863
rect 240 -2907 241 -2865
rect 870 -2866 871 -2790
rect 1045 -2907 1046 -2865
rect 1199 -2866 1200 -2790
rect 394 -2868 395 -2790
rect 415 -2907 416 -2867
rect 548 -2907 549 -2867
rect 716 -2868 717 -2790
rect 786 -2868 787 -2790
rect 877 -2907 878 -2867
rect 1122 -2907 1123 -2867
rect 1318 -2868 1319 -2790
rect 145 -2907 146 -2869
rect 394 -2907 395 -2869
rect 555 -2907 556 -2869
rect 604 -2907 605 -2869
rect 611 -2870 612 -2790
rect 639 -2907 640 -2869
rect 716 -2907 717 -2869
rect 758 -2907 759 -2869
rect 786 -2907 787 -2869
rect 821 -2870 822 -2790
rect 870 -2907 871 -2869
rect 926 -2870 927 -2790
rect 1192 -2870 1193 -2790
rect 1199 -2907 1200 -2869
rect 1318 -2907 1319 -2869
rect 1388 -2870 1389 -2790
rect 569 -2907 570 -2871
rect 835 -2907 836 -2871
rect 926 -2907 927 -2871
rect 933 -2872 934 -2790
rect 1017 -2872 1018 -2790
rect 1192 -2907 1193 -2871
rect 1332 -2872 1333 -2790
rect 1388 -2907 1389 -2871
rect 576 -2907 577 -2873
rect 1038 -2874 1039 -2790
rect 1332 -2907 1333 -2873
rect 1444 -2874 1445 -2790
rect 583 -2876 584 -2790
rect 611 -2907 612 -2875
rect 821 -2907 822 -2875
rect 1108 -2876 1109 -2790
rect 933 -2907 934 -2877
rect 975 -2878 976 -2790
rect 1017 -2907 1018 -2877
rect 1024 -2907 1025 -2877
rect 1038 -2907 1039 -2877
rect 1206 -2878 1207 -2790
rect 975 -2907 976 -2879
rect 1059 -2880 1060 -2790
rect 1108 -2907 1109 -2879
rect 1234 -2880 1235 -2790
rect 1059 -2907 1060 -2881
rect 1080 -2882 1081 -2790
rect 1206 -2907 1207 -2881
rect 1402 -2882 1403 -2790
rect 1080 -2907 1081 -2883
rect 1171 -2884 1172 -2790
rect 1234 -2907 1235 -2883
rect 1346 -2884 1347 -2790
rect 1402 -2907 1403 -2883
rect 1514 -2884 1515 -2790
rect 1171 -2907 1172 -2885
rect 1248 -2886 1249 -2790
rect 1346 -2907 1347 -2885
rect 1451 -2886 1452 -2790
rect 1248 -2907 1249 -2887
rect 1409 -2888 1410 -2790
rect 905 -2890 906 -2790
rect 1409 -2907 1410 -2889
rect 905 -2907 906 -2891
rect 968 -2892 969 -2790
rect 968 -2907 969 -2893
rect 1115 -2894 1116 -2790
rect 1115 -2907 1116 -2895
rect 1178 -2896 1179 -2790
rect 1178 -2907 1179 -2897
rect 1304 -2898 1305 -2790
rect 1304 -2907 1305 -2899
rect 1423 -2900 1424 -2790
rect 1416 -2902 1417 -2790
rect 1423 -2907 1424 -2901
rect 1031 -2904 1032 -2790
rect 1416 -2907 1417 -2903
rect 663 -2907 664 -2905
rect 1031 -2907 1032 -2905
rect 72 -2917 73 -2915
rect 247 -2917 248 -2915
rect 250 -2917 251 -2915
rect 569 -2917 570 -2915
rect 583 -2917 584 -2915
rect 954 -2917 955 -2915
rect 957 -2917 958 -2915
rect 1185 -2917 1186 -2915
rect 1199 -2917 1200 -2915
rect 1199 -3026 1200 -2916
rect 1199 -2917 1200 -2915
rect 1199 -3026 1200 -2916
rect 1227 -2917 1228 -2915
rect 1230 -2917 1231 -2915
rect 1360 -2917 1361 -2915
rect 1430 -2917 1431 -2915
rect 93 -2919 94 -2915
rect 124 -2919 125 -2915
rect 128 -2919 129 -2915
rect 128 -3026 129 -2918
rect 128 -2919 129 -2915
rect 128 -3026 129 -2918
rect 166 -3026 167 -2918
rect 576 -2919 577 -2915
rect 586 -2919 587 -2915
rect 618 -2919 619 -2915
rect 754 -3026 755 -2918
rect 793 -2919 794 -2915
rect 800 -2919 801 -2915
rect 1094 -2919 1095 -2915
rect 1097 -2919 1098 -2915
rect 1248 -2919 1249 -2915
rect 1360 -3026 1361 -2918
rect 1409 -2919 1410 -2915
rect 93 -3026 94 -2920
rect 205 -2921 206 -2915
rect 208 -2921 209 -2915
rect 310 -2921 311 -2915
rect 436 -2921 437 -2915
rect 702 -2921 703 -2915
rect 765 -2921 766 -2915
rect 793 -3026 794 -2920
rect 828 -2921 829 -2915
rect 828 -3026 829 -2920
rect 828 -2921 829 -2915
rect 828 -3026 829 -2920
rect 838 -2921 839 -2915
rect 1192 -2921 1193 -2915
rect 1227 -3026 1228 -2920
rect 1255 -2921 1256 -2915
rect 1409 -3026 1410 -2920
rect 1423 -2921 1424 -2915
rect 100 -3026 101 -2922
rect 149 -2923 150 -2915
rect 184 -2923 185 -2915
rect 285 -2923 286 -2915
rect 289 -2923 290 -2915
rect 296 -2923 297 -2915
rect 310 -3026 311 -2922
rect 324 -2923 325 -2915
rect 457 -2923 458 -2915
rect 824 -2923 825 -2915
rect 838 -3026 839 -2922
rect 884 -2923 885 -2915
rect 891 -2923 892 -2915
rect 894 -2935 895 -2922
rect 912 -2923 913 -2915
rect 1171 -2923 1172 -2915
rect 1178 -2923 1179 -2915
rect 1178 -3026 1179 -2922
rect 1178 -2923 1179 -2915
rect 1178 -3026 1179 -2922
rect 1185 -3026 1186 -2922
rect 1213 -2923 1214 -2915
rect 1248 -3026 1249 -2922
rect 1297 -2923 1298 -2915
rect 103 -2925 104 -2915
rect 744 -2925 745 -2915
rect 768 -3026 769 -2924
rect 1115 -2925 1116 -2915
rect 1136 -2925 1137 -2915
rect 1136 -3026 1137 -2924
rect 1136 -2925 1137 -2915
rect 1136 -3026 1137 -2924
rect 1192 -3026 1193 -2924
rect 1234 -2925 1235 -2915
rect 1276 -2925 1277 -2915
rect 1297 -3026 1298 -2924
rect 121 -2927 122 -2915
rect 849 -2927 850 -2915
rect 884 -3026 885 -2926
rect 926 -2927 927 -2915
rect 947 -2927 948 -2915
rect 982 -2927 983 -2915
rect 996 -2927 997 -2915
rect 996 -3026 997 -2926
rect 996 -2927 997 -2915
rect 996 -3026 997 -2926
rect 1017 -2927 1018 -2915
rect 1059 -2927 1060 -2915
rect 1076 -3026 1077 -2926
rect 1220 -2927 1221 -2915
rect 1234 -3026 1235 -2926
rect 1290 -2927 1291 -2915
rect 121 -3026 122 -2928
rect 212 -2929 213 -2915
rect 219 -2929 220 -2915
rect 576 -3026 577 -2928
rect 604 -2929 605 -2915
rect 618 -3026 619 -2928
rect 667 -2929 668 -2915
rect 702 -3026 703 -2928
rect 744 -3026 745 -2928
rect 751 -2929 752 -2915
rect 789 -3026 790 -2928
rect 1080 -2929 1081 -2915
rect 1087 -2929 1088 -2915
rect 1115 -3026 1116 -2928
rect 1213 -3026 1214 -2928
rect 1241 -2929 1242 -2915
rect 1269 -2929 1270 -2915
rect 1276 -3026 1277 -2928
rect 142 -2931 143 -2915
rect 436 -3026 437 -2930
rect 457 -3026 458 -2930
rect 590 -2931 591 -2915
rect 604 -3026 605 -2930
rect 737 -2931 738 -2915
rect 821 -2931 822 -2915
rect 982 -3026 983 -2930
rect 1024 -2931 1025 -2915
rect 1059 -3026 1060 -2930
rect 1080 -3026 1081 -2930
rect 1129 -2931 1130 -2915
rect 1220 -3026 1221 -2930
rect 1262 -2931 1263 -2915
rect 1269 -3026 1270 -2930
rect 1325 -2931 1326 -2915
rect 107 -2933 108 -2915
rect 590 -3026 591 -2932
rect 611 -2933 612 -2915
rect 642 -2933 643 -2915
rect 646 -2933 647 -2915
rect 667 -3026 668 -2932
rect 681 -2933 682 -2915
rect 849 -3026 850 -2932
rect 891 -3026 892 -2932
rect 912 -3026 913 -2932
rect 989 -2933 990 -2915
rect 1094 -3026 1095 -2932
rect 1157 -2933 1158 -2915
rect 1206 -2933 1207 -2915
rect 1325 -3026 1326 -2932
rect 107 -3026 108 -2934
rect 548 -2935 549 -2915
rect 597 -2935 598 -2915
rect 611 -3026 612 -2934
rect 691 -3026 692 -2934
rect 1087 -3026 1088 -2934
rect 1101 -2935 1102 -2915
rect 1171 -3026 1172 -2934
rect 1230 -3026 1231 -2934
rect 1255 -3026 1256 -2934
rect 1262 -3026 1263 -2934
rect 1311 -2935 1312 -2915
rect 142 -3026 143 -2936
rect 646 -3026 647 -2936
rect 709 -2937 710 -2915
rect 737 -3026 738 -2936
rect 807 -2937 808 -2915
rect 1024 -3026 1025 -2936
rect 1052 -2937 1053 -2915
rect 1157 -3026 1158 -2936
rect 1241 -3026 1242 -2936
rect 1332 -2937 1333 -2915
rect 184 -3026 185 -2938
rect 639 -2939 640 -2915
rect 772 -2939 773 -2915
rect 807 -3026 808 -2938
rect 821 -3026 822 -2938
rect 870 -2939 871 -2915
rect 898 -2939 899 -2915
rect 947 -3026 948 -2938
rect 954 -3026 955 -2938
rect 961 -2939 962 -2915
rect 968 -2939 969 -2915
rect 968 -3026 969 -2938
rect 968 -2939 969 -2915
rect 968 -3026 969 -2938
rect 989 -3026 990 -2938
rect 1045 -2939 1046 -2915
rect 1066 -2939 1067 -2915
rect 1101 -3026 1102 -2938
rect 1129 -3026 1130 -2938
rect 1164 -2939 1165 -2915
rect 1304 -2939 1305 -2915
rect 1332 -3026 1333 -2938
rect 208 -3026 209 -2940
rect 233 -2941 234 -2915
rect 240 -2941 241 -2915
rect 800 -3026 801 -2940
rect 835 -2941 836 -2915
rect 1052 -3026 1053 -2940
rect 1108 -2941 1109 -2915
rect 1164 -3026 1165 -2940
rect 1311 -3026 1312 -2940
rect 1388 -2941 1389 -2915
rect 212 -3026 213 -2942
rect 366 -2943 367 -2915
rect 411 -3026 412 -2942
rect 1290 -3026 1291 -2942
rect 1388 -3026 1389 -2942
rect 1416 -2943 1417 -2915
rect 222 -3026 223 -2944
rect 450 -2945 451 -2915
rect 492 -2945 493 -2915
rect 492 -3026 493 -2944
rect 492 -2945 493 -2915
rect 492 -3026 493 -2944
rect 495 -2945 496 -2915
rect 926 -3026 927 -2944
rect 950 -2945 951 -2915
rect 1045 -3026 1046 -2944
rect 1143 -2945 1144 -2915
rect 1206 -3026 1207 -2944
rect 226 -3026 227 -2946
rect 268 -2947 269 -2915
rect 275 -2947 276 -2915
rect 583 -3026 584 -2946
rect 597 -3026 598 -2946
rect 625 -2947 626 -2915
rect 639 -3026 640 -2946
rect 660 -2947 661 -2915
rect 688 -2947 689 -2915
rect 835 -3026 836 -2946
rect 842 -2947 843 -2915
rect 1395 -2947 1396 -2915
rect 163 -2949 164 -2915
rect 268 -3026 269 -2948
rect 275 -3026 276 -2948
rect 422 -2949 423 -2915
rect 443 -2949 444 -2915
rect 681 -3026 682 -2948
rect 751 -3026 752 -2948
rect 1066 -3026 1067 -2948
rect 1143 -3026 1144 -2948
rect 1150 -2949 1151 -2915
rect 163 -3026 164 -2950
rect 380 -2951 381 -2915
rect 443 -3026 444 -2950
rect 471 -2951 472 -2915
rect 513 -2951 514 -2915
rect 625 -3026 626 -2950
rect 660 -3026 661 -2950
rect 1395 -3026 1396 -2950
rect 135 -2953 136 -2915
rect 471 -3026 472 -2952
rect 520 -2953 521 -2915
rect 649 -3026 650 -2952
rect 772 -3026 773 -2952
rect 786 -2953 787 -2915
rect 842 -3026 843 -2952
rect 856 -2953 857 -2915
rect 870 -3026 871 -2952
rect 1122 -2953 1123 -2915
rect 135 -3026 136 -2954
rect 653 -2955 654 -2915
rect 898 -3026 899 -2954
rect 933 -2955 934 -2915
rect 961 -3026 962 -2954
rect 975 -2955 976 -2915
rect 1017 -3026 1018 -2954
rect 1122 -3026 1123 -2954
rect 149 -3026 150 -2956
rect 856 -3026 857 -2956
rect 915 -2957 916 -2915
rect 1038 -2957 1039 -2915
rect 191 -2959 192 -2915
rect 422 -3026 423 -2958
rect 464 -2959 465 -2915
rect 933 -3026 934 -2958
rect 1031 -2959 1032 -2915
rect 1304 -3026 1305 -2958
rect 191 -3026 192 -2960
rect 198 -2961 199 -2915
rect 229 -2961 230 -2915
rect 632 -2961 633 -2915
rect 786 -3026 787 -2960
rect 975 -3026 976 -2960
rect 1038 -3026 1039 -2960
rect 1073 -2961 1074 -2915
rect 86 -2963 87 -2915
rect 198 -3026 199 -2962
rect 233 -3026 234 -2962
rect 292 -2963 293 -2915
rect 296 -3026 297 -2962
rect 688 -3026 689 -2962
rect 919 -2963 920 -2915
rect 1003 -2963 1004 -2915
rect 1073 -3026 1074 -2962
rect 1318 -2963 1319 -2915
rect 79 -2965 80 -2915
rect 86 -3026 87 -2964
rect 219 -3026 220 -2964
rect 919 -3026 920 -2964
rect 940 -2965 941 -2915
rect 1031 -3026 1032 -2964
rect 1283 -2965 1284 -2915
rect 1318 -3026 1319 -2964
rect 240 -3026 241 -2966
rect 373 -2967 374 -2915
rect 387 -2967 388 -2915
rect 653 -3026 654 -2966
rect 674 -2967 675 -2915
rect 940 -3026 941 -2966
rect 1003 -3026 1004 -2966
rect 1010 -2967 1011 -2915
rect 1283 -3026 1284 -2966
rect 1339 -2967 1340 -2915
rect 170 -2969 171 -2915
rect 387 -3026 388 -2968
rect 401 -2969 402 -2915
rect 513 -3026 514 -2968
rect 520 -3026 521 -2968
rect 866 -2969 867 -2915
rect 1339 -3026 1340 -2968
rect 1346 -2969 1347 -2915
rect 170 -3026 171 -2970
rect 873 -3026 874 -2970
rect 1346 -3026 1347 -2970
rect 1381 -2971 1382 -2915
rect 247 -3026 248 -2972
rect 761 -2973 762 -2915
rect 282 -2975 283 -2915
rect 747 -2975 748 -2915
rect 254 -2977 255 -2915
rect 282 -3026 283 -2976
rect 289 -3026 290 -2976
rect 663 -2977 664 -2915
rect 674 -3026 675 -2976
rect 915 -3026 916 -2976
rect 254 -3026 255 -2978
rect 278 -2979 279 -2915
rect 303 -2979 304 -2915
rect 366 -3026 367 -2978
rect 373 -3026 374 -2978
rect 394 -2979 395 -2915
rect 464 -3026 465 -2978
rect 485 -2979 486 -2915
rect 534 -2979 535 -2915
rect 569 -3026 570 -2978
rect 632 -3026 633 -2978
rect 1108 -3026 1109 -2978
rect 261 -2981 262 -2915
rect 534 -3026 535 -2980
rect 548 -3026 549 -2980
rect 877 -2981 878 -2915
rect 261 -3026 262 -2982
rect 380 -3026 381 -2982
rect 394 -3026 395 -2982
rect 408 -2983 409 -2915
rect 485 -3026 486 -2982
rect 716 -2983 717 -2915
rect 303 -3026 304 -2984
rect 317 -2985 318 -2915
rect 324 -3026 325 -2984
rect 506 -2985 507 -2915
rect 555 -3026 556 -2984
rect 866 -3026 867 -2984
rect 317 -3026 318 -2986
rect 338 -2987 339 -2915
rect 345 -2987 346 -2915
rect 450 -3026 451 -2986
rect 562 -2987 563 -2915
rect 709 -3026 710 -2986
rect 716 -3026 717 -2986
rect 863 -2987 864 -2915
rect 145 -2989 146 -2915
rect 338 -3026 339 -2988
rect 345 -3026 346 -2988
rect 499 -2989 500 -2915
rect 695 -2989 696 -2915
rect 863 -3026 864 -2988
rect 264 -3026 265 -2990
rect 562 -3026 563 -2990
rect 698 -3026 699 -2990
rect 1010 -3026 1011 -2990
rect 359 -2993 360 -2915
rect 401 -3026 402 -2992
rect 408 -3026 409 -2992
rect 877 -3026 878 -2992
rect 359 -3026 360 -2994
rect 478 -2995 479 -2915
rect 499 -3026 500 -2994
rect 635 -3026 636 -2994
rect 705 -2995 706 -2915
rect 1381 -3026 1382 -2994
rect 429 -2997 430 -2915
rect 695 -3026 696 -2996
rect 177 -2999 178 -2915
rect 429 -3026 430 -2998
rect 478 -3026 479 -2998
rect 541 -2999 542 -2915
rect 156 -3001 157 -2915
rect 177 -3026 178 -3000
rect 541 -3026 542 -3000
rect 723 -3001 724 -2915
rect 156 -3026 157 -3002
rect 352 -3003 353 -2915
rect 723 -3026 724 -3002
rect 730 -3003 731 -2915
rect 352 -3026 353 -3004
rect 415 -3005 416 -2915
rect 730 -3026 731 -3004
rect 814 -3005 815 -2915
rect 331 -3007 332 -2915
rect 415 -3026 416 -3006
rect 779 -3007 780 -2915
rect 814 -3026 815 -3006
rect 114 -3009 115 -2915
rect 331 -3026 332 -3008
rect 779 -3026 780 -3008
rect 922 -3009 923 -2915
rect 114 -3026 115 -3010
rect 1020 -3011 1021 -2915
rect 922 -3026 923 -3012
rect 1353 -3013 1354 -2915
rect 1353 -3026 1354 -3014
rect 1367 -3015 1368 -2915
rect 1367 -3026 1368 -3016
rect 1374 -3017 1375 -2915
rect 1374 -3026 1375 -3018
rect 1402 -3019 1403 -2915
rect 758 -3021 759 -2915
rect 1402 -3026 1403 -3020
rect 527 -3023 528 -2915
rect 758 -3026 759 -3022
rect 527 -3026 528 -3024
rect 663 -3026 664 -3024
rect 86 -3036 87 -3034
rect 149 -3036 150 -3034
rect 156 -3036 157 -3034
rect 408 -3036 409 -3034
rect 411 -3036 412 -3034
rect 653 -3036 654 -3034
rect 660 -3036 661 -3034
rect 982 -3036 983 -3034
rect 1017 -3137 1018 -3035
rect 1045 -3036 1046 -3034
rect 1073 -3036 1074 -3034
rect 1402 -3036 1403 -3034
rect 93 -3038 94 -3034
rect 810 -3137 811 -3037
rect 835 -3038 836 -3034
rect 1171 -3038 1172 -3034
rect 1283 -3038 1284 -3034
rect 1283 -3137 1284 -3037
rect 1283 -3038 1284 -3034
rect 1283 -3137 1284 -3037
rect 100 -3040 101 -3034
rect 152 -3040 153 -3034
rect 198 -3040 199 -3034
rect 208 -3040 209 -3034
rect 275 -3040 276 -3034
rect 278 -3074 279 -3039
rect 289 -3040 290 -3034
rect 506 -3137 507 -3039
rect 516 -3137 517 -3039
rect 541 -3040 542 -3034
rect 555 -3040 556 -3034
rect 653 -3137 654 -3039
rect 660 -3137 661 -3039
rect 877 -3040 878 -3034
rect 919 -3040 920 -3034
rect 1332 -3040 1333 -3034
rect 100 -3137 101 -3041
rect 128 -3042 129 -3034
rect 135 -3042 136 -3034
rect 205 -3137 206 -3041
rect 275 -3137 276 -3041
rect 366 -3042 367 -3034
rect 422 -3042 423 -3034
rect 915 -3137 916 -3041
rect 926 -3042 927 -3034
rect 1335 -3137 1336 -3041
rect 107 -3044 108 -3034
rect 222 -3137 223 -3043
rect 310 -3044 311 -3034
rect 411 -3137 412 -3043
rect 450 -3044 451 -3034
rect 450 -3137 451 -3043
rect 450 -3044 451 -3034
rect 450 -3137 451 -3043
rect 471 -3044 472 -3034
rect 541 -3137 542 -3043
rect 569 -3044 570 -3034
rect 569 -3137 570 -3043
rect 569 -3044 570 -3034
rect 569 -3137 570 -3043
rect 576 -3044 577 -3034
rect 632 -3137 633 -3043
rect 681 -3044 682 -3034
rect 695 -3044 696 -3034
rect 698 -3044 699 -3034
rect 989 -3044 990 -3034
rect 1020 -3044 1021 -3034
rect 1276 -3044 1277 -3034
rect 107 -3137 108 -3045
rect 261 -3046 262 -3034
rect 310 -3137 311 -3045
rect 866 -3046 867 -3034
rect 873 -3046 874 -3034
rect 1395 -3046 1396 -3034
rect 114 -3048 115 -3034
rect 114 -3137 115 -3047
rect 114 -3048 115 -3034
rect 114 -3137 115 -3047
rect 128 -3137 129 -3047
rect 233 -3048 234 -3034
rect 324 -3048 325 -3034
rect 838 -3048 839 -3034
rect 863 -3048 864 -3034
rect 1325 -3048 1326 -3034
rect 135 -3137 136 -3049
rect 1209 -3137 1210 -3049
rect 1241 -3050 1242 -3034
rect 1276 -3137 1277 -3049
rect 1325 -3137 1326 -3049
rect 1381 -3050 1382 -3034
rect 142 -3052 143 -3034
rect 142 -3137 143 -3051
rect 142 -3052 143 -3034
rect 142 -3137 143 -3051
rect 149 -3137 150 -3051
rect 922 -3052 923 -3034
rect 926 -3137 927 -3051
rect 996 -3052 997 -3034
rect 1038 -3052 1039 -3034
rect 1073 -3137 1074 -3051
rect 1136 -3052 1137 -3034
rect 1171 -3137 1172 -3051
rect 1241 -3137 1242 -3051
rect 1269 -3052 1270 -3034
rect 170 -3054 171 -3034
rect 198 -3137 199 -3053
rect 229 -3137 230 -3053
rect 261 -3137 262 -3053
rect 327 -3137 328 -3053
rect 646 -3137 647 -3053
rect 691 -3054 692 -3034
rect 1255 -3054 1256 -3034
rect 170 -3137 171 -3055
rect 247 -3137 248 -3055
rect 338 -3056 339 -3034
rect 471 -3137 472 -3055
rect 513 -3056 514 -3034
rect 555 -3137 556 -3055
rect 583 -3056 584 -3034
rect 989 -3137 990 -3055
rect 1038 -3137 1039 -3055
rect 1066 -3056 1067 -3034
rect 1115 -3056 1116 -3034
rect 1136 -3137 1137 -3055
rect 1150 -3056 1151 -3034
rect 1297 -3056 1298 -3034
rect 184 -3058 185 -3034
rect 289 -3137 290 -3057
rect 338 -3137 339 -3057
rect 527 -3058 528 -3034
rect 534 -3058 535 -3034
rect 607 -3137 608 -3057
rect 618 -3058 619 -3034
rect 649 -3058 650 -3034
rect 698 -3137 699 -3057
rect 1178 -3058 1179 -3034
rect 1234 -3058 1235 -3034
rect 1255 -3137 1256 -3057
rect 1297 -3137 1298 -3057
rect 1332 -3137 1333 -3057
rect 184 -3137 185 -3059
rect 226 -3060 227 -3034
rect 233 -3137 234 -3059
rect 254 -3060 255 -3034
rect 345 -3060 346 -3034
rect 509 -3060 510 -3034
rect 527 -3137 528 -3059
rect 590 -3060 591 -3034
rect 618 -3137 619 -3059
rect 765 -3060 766 -3034
rect 789 -3060 790 -3034
rect 870 -3137 871 -3059
rect 877 -3137 878 -3059
rect 1220 -3060 1221 -3034
rect 121 -3062 122 -3034
rect 226 -3137 227 -3061
rect 345 -3137 346 -3061
rect 436 -3062 437 -3034
rect 443 -3062 444 -3034
rect 576 -3137 577 -3061
rect 590 -3137 591 -3061
rect 1087 -3062 1088 -3034
rect 1150 -3137 1151 -3061
rect 1206 -3062 1207 -3034
rect 1220 -3137 1221 -3061
rect 1227 -3062 1228 -3034
rect 121 -3137 122 -3063
rect 219 -3064 220 -3034
rect 331 -3064 332 -3034
rect 436 -3137 437 -3063
rect 464 -3064 465 -3034
rect 513 -3137 514 -3063
rect 534 -3137 535 -3063
rect 597 -3064 598 -3034
rect 625 -3064 626 -3034
rect 625 -3137 626 -3063
rect 625 -3064 626 -3034
rect 625 -3137 626 -3063
rect 635 -3064 636 -3034
rect 681 -3137 682 -3063
rect 730 -3064 731 -3034
rect 733 -3064 734 -3034
rect 740 -3137 741 -3063
rect 947 -3064 948 -3034
rect 982 -3137 983 -3063
rect 1202 -3137 1203 -3063
rect 1213 -3064 1214 -3034
rect 1227 -3137 1228 -3063
rect 166 -3066 167 -3034
rect 331 -3137 332 -3065
rect 352 -3066 353 -3034
rect 366 -3137 367 -3065
rect 380 -3066 381 -3034
rect 464 -3137 465 -3065
rect 478 -3066 479 -3034
rect 583 -3137 584 -3065
rect 597 -3137 598 -3065
rect 667 -3066 668 -3034
rect 730 -3137 731 -3065
rect 793 -3066 794 -3034
rect 796 -3137 797 -3065
rect 1234 -3137 1235 -3065
rect 177 -3068 178 -3034
rect 254 -3137 255 -3067
rect 257 -3137 258 -3067
rect 478 -3137 479 -3067
rect 520 -3068 521 -3034
rect 667 -3137 668 -3067
rect 744 -3068 745 -3034
rect 765 -3137 766 -3067
rect 835 -3137 836 -3067
rect 842 -3068 843 -3034
rect 863 -3137 864 -3067
rect 891 -3068 892 -3034
rect 898 -3068 899 -3034
rect 919 -3137 920 -3067
rect 1045 -3137 1046 -3067
rect 1101 -3068 1102 -3034
rect 1178 -3137 1179 -3067
rect 1367 -3068 1368 -3034
rect 177 -3137 178 -3069
rect 499 -3070 500 -3034
rect 520 -3137 521 -3069
rect 639 -3070 640 -3034
rect 649 -3137 650 -3069
rect 1087 -3137 1088 -3069
rect 1101 -3137 1102 -3069
rect 1122 -3070 1123 -3034
rect 1213 -3137 1214 -3069
rect 1304 -3070 1305 -3034
rect 1367 -3137 1368 -3069
rect 1388 -3070 1389 -3034
rect 352 -3137 353 -3071
rect 380 -3137 381 -3071
rect 457 -3072 458 -3034
rect 499 -3137 500 -3071
rect 604 -3072 605 -3034
rect 611 -3072 612 -3034
rect 639 -3137 640 -3071
rect 744 -3137 745 -3071
rect 1157 -3072 1158 -3034
rect 1304 -3137 1305 -3071
rect 1353 -3072 1354 -3034
rect 394 -3074 395 -3034
rect 422 -3137 423 -3073
rect 429 -3074 430 -3034
rect 457 -3137 458 -3073
rect 548 -3074 549 -3034
rect 611 -3137 612 -3073
rect 733 -3137 734 -3073
rect 793 -3137 794 -3073
rect 842 -3137 843 -3073
rect 905 -3074 906 -3034
rect 933 -3074 934 -3034
rect 1157 -3137 1158 -3073
rect 1353 -3137 1354 -3073
rect 1360 -3074 1361 -3034
rect 303 -3076 304 -3034
rect 548 -3137 549 -3075
rect 747 -3137 748 -3075
rect 1269 -3137 1270 -3075
rect 1360 -3137 1361 -3075
rect 1374 -3076 1375 -3034
rect 303 -3137 304 -3077
rect 387 -3078 388 -3034
rect 394 -3137 395 -3077
rect 761 -3137 762 -3077
rect 887 -3078 888 -3034
rect 947 -3137 948 -3077
rect 1059 -3078 1060 -3034
rect 1066 -3137 1067 -3077
rect 1122 -3137 1123 -3077
rect 1129 -3078 1130 -3034
rect 1374 -3137 1375 -3077
rect 1409 -3078 1410 -3034
rect 401 -3080 402 -3034
rect 429 -3137 430 -3079
rect 751 -3137 752 -3079
rect 779 -3080 780 -3034
rect 891 -3137 892 -3079
rect 954 -3080 955 -3034
rect 1059 -3137 1060 -3079
rect 1080 -3080 1081 -3034
rect 1108 -3080 1109 -3034
rect 1129 -3137 1130 -3079
rect 296 -3082 297 -3034
rect 401 -3137 402 -3081
rect 415 -3082 416 -3034
rect 443 -3137 444 -3081
rect 772 -3082 773 -3034
rect 779 -3137 780 -3081
rect 898 -3137 899 -3081
rect 1199 -3082 1200 -3034
rect 296 -3137 297 -3083
rect 373 -3084 374 -3034
rect 415 -3137 416 -3083
rect 754 -3084 755 -3034
rect 758 -3084 759 -3034
rect 772 -3137 773 -3083
rect 901 -3137 902 -3083
rect 1115 -3137 1116 -3083
rect 373 -3137 374 -3085
rect 688 -3086 689 -3034
rect 905 -3137 906 -3085
rect 1024 -3086 1025 -3034
rect 1080 -3137 1081 -3085
rect 1143 -3086 1144 -3034
rect 688 -3137 689 -3087
rect 723 -3088 724 -3034
rect 933 -3137 934 -3087
rect 961 -3088 962 -3034
rect 1024 -3137 1025 -3087
rect 1052 -3088 1053 -3034
rect 1108 -3137 1109 -3087
rect 1192 -3088 1193 -3034
rect 674 -3090 675 -3034
rect 1052 -3137 1053 -3089
rect 1143 -3137 1144 -3089
rect 1185 -3090 1186 -3034
rect 1192 -3137 1193 -3089
rect 1290 -3090 1291 -3034
rect 674 -3137 675 -3091
rect 702 -3092 703 -3034
rect 716 -3092 717 -3034
rect 723 -3137 724 -3091
rect 940 -3092 941 -3034
rect 961 -3137 962 -3091
rect 1003 -3092 1004 -3034
rect 1185 -3137 1186 -3091
rect 1290 -3137 1291 -3091
rect 1339 -3092 1340 -3034
rect 485 -3094 486 -3034
rect 716 -3137 717 -3093
rect 940 -3137 941 -3093
rect 968 -3094 969 -3034
rect 1003 -3137 1004 -3093
rect 1031 -3094 1032 -3034
rect 1339 -3137 1340 -3093
rect 1346 -3094 1347 -3034
rect 317 -3096 318 -3034
rect 485 -3137 486 -3095
rect 702 -3137 703 -3095
rect 709 -3096 710 -3034
rect 912 -3096 913 -3034
rect 968 -3137 969 -3095
rect 1031 -3137 1032 -3095
rect 1094 -3096 1095 -3034
rect 163 -3098 164 -3034
rect 1094 -3137 1095 -3097
rect 163 -3137 164 -3099
rect 268 -3100 269 -3034
rect 317 -3137 318 -3099
rect 359 -3100 360 -3034
rect 562 -3100 563 -3034
rect 709 -3137 710 -3099
rect 912 -3137 913 -3099
rect 1164 -3100 1165 -3034
rect 212 -3102 213 -3034
rect 268 -3137 269 -3101
rect 324 -3137 325 -3101
rect 562 -3137 563 -3101
rect 954 -3137 955 -3101
rect 975 -3102 976 -3034
rect 1164 -3137 1165 -3101
rect 1262 -3102 1263 -3034
rect 191 -3104 192 -3034
rect 212 -3137 213 -3103
rect 240 -3104 241 -3034
rect 359 -3137 360 -3103
rect 975 -3137 976 -3103
rect 1010 -3104 1011 -3034
rect 1248 -3104 1249 -3034
rect 1262 -3137 1263 -3103
rect 156 -3137 157 -3105
rect 191 -3137 192 -3105
rect 240 -3137 241 -3105
rect 1153 -3106 1154 -3034
rect 695 -3137 696 -3107
rect 1248 -3137 1249 -3107
rect 1010 -3137 1011 -3109
rect 1318 -3110 1319 -3034
rect 1311 -3112 1312 -3034
rect 1318 -3137 1319 -3111
rect 884 -3114 885 -3034
rect 1311 -3137 1312 -3113
rect 856 -3116 857 -3034
rect 884 -3137 885 -3115
rect 849 -3118 850 -3034
rect 856 -3137 857 -3117
rect 828 -3120 829 -3034
rect 849 -3137 850 -3119
rect 814 -3122 815 -3034
rect 828 -3137 829 -3121
rect 814 -3137 815 -3123
rect 821 -3124 822 -3034
rect 737 -3126 738 -3034
rect 821 -3137 822 -3125
rect 492 -3128 493 -3034
rect 737 -3137 738 -3127
rect 492 -3137 493 -3129
rect 786 -3130 787 -3034
rect 786 -3137 787 -3131
rect 800 -3132 801 -3034
rect 800 -3137 801 -3133
rect 807 -3134 808 -3034
rect 807 -3137 808 -3135
rect 996 -3137 997 -3135
rect 100 -3147 101 -3145
rect 159 -3147 160 -3145
rect 184 -3147 185 -3145
rect 324 -3147 325 -3145
rect 331 -3147 332 -3145
rect 390 -3147 391 -3145
rect 394 -3147 395 -3145
rect 754 -3230 755 -3146
rect 758 -3147 759 -3145
rect 814 -3147 815 -3145
rect 842 -3147 843 -3145
rect 842 -3230 843 -3146
rect 842 -3147 843 -3145
rect 842 -3230 843 -3146
rect 863 -3147 864 -3145
rect 863 -3230 864 -3146
rect 863 -3147 864 -3145
rect 863 -3230 864 -3146
rect 898 -3147 899 -3145
rect 1171 -3147 1172 -3145
rect 1199 -3147 1200 -3145
rect 1220 -3147 1221 -3145
rect 1293 -3230 1294 -3146
rect 1339 -3147 1340 -3145
rect 1346 -3230 1347 -3146
rect 1360 -3147 1361 -3145
rect 107 -3149 108 -3145
rect 285 -3230 286 -3148
rect 296 -3149 297 -3145
rect 695 -3149 696 -3145
rect 698 -3149 699 -3145
rect 968 -3149 969 -3145
rect 1045 -3149 1046 -3145
rect 1045 -3230 1046 -3148
rect 1045 -3149 1046 -3145
rect 1045 -3230 1046 -3148
rect 1171 -3230 1172 -3148
rect 1213 -3149 1214 -3145
rect 1297 -3149 1298 -3145
rect 1297 -3230 1298 -3148
rect 1297 -3149 1298 -3145
rect 1297 -3230 1298 -3148
rect 1335 -3149 1336 -3145
rect 1367 -3149 1368 -3145
rect 114 -3151 115 -3145
rect 187 -3230 188 -3150
rect 191 -3151 192 -3145
rect 250 -3151 251 -3145
rect 254 -3230 255 -3150
rect 373 -3151 374 -3145
rect 387 -3151 388 -3145
rect 485 -3151 486 -3145
rect 492 -3151 493 -3145
rect 810 -3151 811 -3145
rect 870 -3151 871 -3145
rect 898 -3230 899 -3150
rect 912 -3230 913 -3150
rect 1199 -3230 1200 -3150
rect 1206 -3151 1207 -3145
rect 1241 -3151 1242 -3145
rect 1353 -3151 1354 -3145
rect 1353 -3230 1354 -3150
rect 1353 -3151 1354 -3145
rect 1353 -3230 1354 -3150
rect 1360 -3230 1361 -3150
rect 1374 -3151 1375 -3145
rect 121 -3153 122 -3145
rect 222 -3153 223 -3145
rect 247 -3153 248 -3145
rect 352 -3153 353 -3145
rect 373 -3230 374 -3152
rect 429 -3153 430 -3145
rect 460 -3230 461 -3152
rect 527 -3153 528 -3145
rect 593 -3153 594 -3145
rect 1286 -3230 1287 -3152
rect 177 -3155 178 -3145
rect 387 -3230 388 -3154
rect 394 -3230 395 -3154
rect 457 -3155 458 -3145
rect 464 -3155 465 -3145
rect 544 -3230 545 -3154
rect 607 -3155 608 -3145
rect 1157 -3155 1158 -3145
rect 1206 -3230 1207 -3154
rect 1276 -3155 1277 -3145
rect 177 -3230 178 -3156
rect 768 -3230 769 -3156
rect 807 -3157 808 -3145
rect 894 -3230 895 -3156
rect 915 -3157 916 -3145
rect 1230 -3230 1231 -3156
rect 1241 -3230 1242 -3156
rect 1318 -3157 1319 -3145
rect 191 -3230 192 -3158
rect 747 -3159 748 -3145
rect 758 -3230 759 -3158
rect 849 -3159 850 -3145
rect 870 -3230 871 -3158
rect 884 -3159 885 -3145
rect 943 -3230 944 -3158
rect 1136 -3159 1137 -3145
rect 1209 -3159 1210 -3145
rect 1220 -3230 1221 -3158
rect 1276 -3230 1277 -3158
rect 1325 -3159 1326 -3145
rect 198 -3161 199 -3145
rect 226 -3230 227 -3160
rect 233 -3161 234 -3145
rect 247 -3230 248 -3160
rect 268 -3161 269 -3145
rect 268 -3230 269 -3160
rect 268 -3161 269 -3145
rect 268 -3230 269 -3160
rect 275 -3161 276 -3145
rect 296 -3230 297 -3160
rect 327 -3161 328 -3145
rect 485 -3230 486 -3160
rect 492 -3230 493 -3160
rect 611 -3161 612 -3145
rect 618 -3161 619 -3145
rect 1010 -3161 1011 -3145
rect 1059 -3161 1060 -3145
rect 1136 -3230 1137 -3160
rect 1213 -3230 1214 -3160
rect 1304 -3161 1305 -3145
rect 128 -3163 129 -3145
rect 198 -3230 199 -3162
rect 212 -3163 213 -3145
rect 212 -3230 213 -3162
rect 212 -3163 213 -3145
rect 212 -3230 213 -3162
rect 219 -3230 220 -3162
rect 289 -3163 290 -3145
rect 331 -3230 332 -3162
rect 380 -3163 381 -3145
rect 401 -3163 402 -3145
rect 618 -3230 619 -3162
rect 635 -3230 636 -3162
rect 828 -3163 829 -3145
rect 849 -3230 850 -3162
rect 975 -3163 976 -3145
rect 1234 -3163 1235 -3145
rect 1304 -3230 1305 -3162
rect 135 -3165 136 -3145
rect 275 -3230 276 -3164
rect 338 -3165 339 -3145
rect 590 -3165 591 -3145
rect 611 -3230 612 -3164
rect 681 -3165 682 -3145
rect 695 -3230 696 -3164
rect 772 -3165 773 -3145
rect 810 -3230 811 -3164
rect 1185 -3165 1186 -3145
rect 1234 -3230 1235 -3164
rect 1290 -3165 1291 -3145
rect 184 -3230 185 -3166
rect 289 -3230 290 -3166
rect 338 -3230 339 -3166
rect 366 -3167 367 -3145
rect 401 -3230 402 -3166
rect 436 -3167 437 -3145
rect 464 -3230 465 -3166
rect 1332 -3167 1333 -3145
rect 233 -3230 234 -3168
rect 282 -3169 283 -3145
rect 345 -3169 346 -3145
rect 747 -3230 748 -3168
rect 772 -3230 773 -3168
rect 786 -3169 787 -3145
rect 877 -3169 878 -3145
rect 1059 -3230 1060 -3168
rect 1108 -3169 1109 -3145
rect 1185 -3230 1186 -3168
rect 282 -3230 283 -3170
rect 324 -3230 325 -3170
rect 345 -3230 346 -3170
rect 450 -3171 451 -3145
rect 506 -3171 507 -3145
rect 744 -3171 745 -3145
rect 761 -3171 762 -3145
rect 786 -3230 787 -3170
rect 877 -3230 878 -3170
rect 954 -3171 955 -3145
rect 968 -3230 969 -3170
rect 982 -3171 983 -3145
rect 1108 -3230 1109 -3170
rect 1227 -3171 1228 -3145
rect 205 -3173 206 -3145
rect 450 -3230 451 -3172
rect 471 -3173 472 -3145
rect 506 -3230 507 -3172
rect 520 -3173 521 -3145
rect 737 -3173 738 -3145
rect 740 -3173 741 -3145
rect 1157 -3230 1158 -3172
rect 205 -3230 206 -3174
rect 261 -3175 262 -3145
rect 352 -3230 353 -3174
rect 534 -3175 535 -3145
rect 590 -3230 591 -3174
rect 744 -3230 745 -3174
rect 884 -3230 885 -3174
rect 891 -3175 892 -3145
rect 905 -3175 906 -3145
rect 954 -3230 955 -3174
rect 975 -3230 976 -3174
rect 1024 -3175 1025 -3145
rect 142 -3177 143 -3145
rect 261 -3230 262 -3176
rect 317 -3177 318 -3145
rect 891 -3230 892 -3176
rect 905 -3230 906 -3176
rect 933 -3177 934 -3145
rect 982 -3230 983 -3176
rect 1017 -3177 1018 -3145
rect 1024 -3230 1025 -3176
rect 1101 -3177 1102 -3145
rect 240 -3179 241 -3145
rect 317 -3230 318 -3178
rect 359 -3179 360 -3145
rect 380 -3230 381 -3178
rect 415 -3179 416 -3145
rect 429 -3230 430 -3178
rect 471 -3230 472 -3178
rect 555 -3179 556 -3145
rect 625 -3179 626 -3145
rect 737 -3230 738 -3178
rect 919 -3179 920 -3145
rect 1010 -3230 1011 -3178
rect 1101 -3230 1102 -3178
rect 1143 -3179 1144 -3145
rect 240 -3230 241 -3180
rect 604 -3181 605 -3145
rect 646 -3181 647 -3145
rect 765 -3181 766 -3145
rect 919 -3230 920 -3180
rect 1202 -3181 1203 -3145
rect 359 -3230 360 -3182
rect 411 -3183 412 -3145
rect 422 -3183 423 -3145
rect 436 -3230 437 -3182
rect 443 -3183 444 -3145
rect 604 -3230 605 -3182
rect 646 -3230 647 -3182
rect 709 -3183 710 -3145
rect 716 -3183 717 -3145
rect 901 -3183 902 -3145
rect 926 -3183 927 -3145
rect 933 -3230 934 -3182
rect 996 -3183 997 -3145
rect 1017 -3230 1018 -3182
rect 1143 -3230 1144 -3182
rect 1262 -3183 1263 -3145
rect 366 -3230 367 -3184
rect 639 -3185 640 -3145
rect 667 -3185 668 -3145
rect 828 -3230 829 -3184
rect 926 -3230 927 -3184
rect 1003 -3185 1004 -3145
rect 1150 -3185 1151 -3145
rect 1202 -3230 1203 -3184
rect 408 -3187 409 -3145
rect 415 -3230 416 -3186
rect 422 -3230 423 -3186
rect 499 -3187 500 -3145
rect 513 -3187 514 -3145
rect 625 -3230 626 -3186
rect 667 -3230 668 -3186
rect 793 -3187 794 -3145
rect 961 -3187 962 -3145
rect 1262 -3230 1263 -3186
rect 163 -3189 164 -3145
rect 408 -3230 409 -3188
rect 443 -3230 444 -3188
rect 457 -3230 458 -3188
rect 513 -3230 514 -3188
rect 653 -3189 654 -3145
rect 681 -3230 682 -3188
rect 751 -3189 752 -3145
rect 765 -3230 766 -3188
rect 1311 -3189 1312 -3145
rect 156 -3191 157 -3145
rect 163 -3230 164 -3190
rect 303 -3191 304 -3145
rect 499 -3230 500 -3190
rect 520 -3230 521 -3190
rect 548 -3191 549 -3145
rect 555 -3230 556 -3190
rect 569 -3191 570 -3145
rect 597 -3191 598 -3145
rect 639 -3230 640 -3190
rect 709 -3230 710 -3190
rect 1178 -3191 1179 -3145
rect 303 -3230 304 -3192
rect 310 -3193 311 -3145
rect 527 -3230 528 -3192
rect 541 -3193 542 -3145
rect 548 -3230 549 -3192
rect 576 -3193 577 -3145
rect 597 -3230 598 -3192
rect 807 -3230 808 -3192
rect 996 -3230 997 -3192
rect 1094 -3193 1095 -3145
rect 1150 -3230 1151 -3192
rect 1269 -3193 1270 -3145
rect 149 -3195 150 -3145
rect 310 -3230 311 -3194
rect 534 -3230 535 -3194
rect 821 -3195 822 -3145
rect 947 -3195 948 -3145
rect 1094 -3230 1095 -3194
rect 562 -3197 563 -3145
rect 653 -3230 654 -3196
rect 716 -3230 717 -3196
rect 730 -3197 731 -3145
rect 751 -3230 752 -3196
rect 1178 -3230 1179 -3196
rect 562 -3230 563 -3198
rect 583 -3199 584 -3145
rect 730 -3230 731 -3198
rect 779 -3199 780 -3145
rect 793 -3230 794 -3198
rect 800 -3199 801 -3145
rect 821 -3230 822 -3198
rect 835 -3199 836 -3145
rect 940 -3199 941 -3145
rect 947 -3230 948 -3198
rect 1003 -3230 1004 -3198
rect 1073 -3199 1074 -3145
rect 170 -3201 171 -3145
rect 800 -3230 801 -3200
rect 835 -3230 836 -3200
rect 856 -3201 857 -3145
rect 940 -3230 941 -3200
rect 1066 -3201 1067 -3145
rect 170 -3230 171 -3202
rect 723 -3203 724 -3145
rect 856 -3230 857 -3202
rect 989 -3203 990 -3145
rect 1031 -3203 1032 -3145
rect 1073 -3230 1074 -3202
rect 478 -3205 479 -3145
rect 779 -3230 780 -3204
rect 989 -3230 990 -3204
rect 1038 -3205 1039 -3145
rect 1066 -3230 1067 -3204
rect 1255 -3205 1256 -3145
rect 478 -3230 479 -3206
rect 1129 -3207 1130 -3145
rect 516 -3209 517 -3145
rect 583 -3230 584 -3208
rect 723 -3230 724 -3208
rect 1087 -3209 1088 -3145
rect 1129 -3230 1130 -3208
rect 1248 -3209 1249 -3145
rect 569 -3230 570 -3210
rect 632 -3211 633 -3145
rect 814 -3230 815 -3210
rect 1255 -3230 1256 -3210
rect 229 -3213 230 -3145
rect 632 -3230 633 -3212
rect 1031 -3230 1032 -3212
rect 1115 -3213 1116 -3145
rect 1248 -3230 1249 -3212
rect 1283 -3213 1284 -3145
rect 576 -3230 577 -3214
rect 702 -3215 703 -3145
rect 961 -3230 962 -3214
rect 1115 -3230 1116 -3214
rect 1269 -3230 1270 -3214
rect 1283 -3230 1284 -3214
rect 688 -3217 689 -3145
rect 702 -3230 703 -3216
rect 1038 -3230 1039 -3216
rect 1052 -3217 1053 -3145
rect 1087 -3230 1088 -3216
rect 1290 -3230 1291 -3216
rect 660 -3219 661 -3145
rect 688 -3230 689 -3218
rect 1052 -3230 1053 -3218
rect 1080 -3219 1081 -3145
rect 660 -3230 661 -3220
rect 674 -3221 675 -3145
rect 1080 -3230 1081 -3220
rect 1122 -3221 1123 -3145
rect 674 -3230 675 -3222
rect 1167 -3230 1168 -3222
rect 1122 -3230 1123 -3224
rect 1164 -3225 1165 -3145
rect 1164 -3230 1165 -3226
rect 1192 -3227 1193 -3145
rect 796 -3229 797 -3145
rect 1192 -3230 1193 -3228
rect 156 -3307 157 -3239
rect 212 -3240 213 -3238
rect 219 -3240 220 -3238
rect 460 -3240 461 -3238
rect 499 -3240 500 -3238
rect 709 -3240 710 -3238
rect 712 -3240 713 -3238
rect 1255 -3240 1256 -3238
rect 1290 -3307 1291 -3239
rect 1304 -3240 1305 -3238
rect 1339 -3307 1340 -3239
rect 1360 -3240 1361 -3238
rect 163 -3242 164 -3238
rect 201 -3307 202 -3241
rect 212 -3307 213 -3241
rect 240 -3242 241 -3238
rect 243 -3307 244 -3241
rect 324 -3242 325 -3238
rect 352 -3242 353 -3238
rect 663 -3307 664 -3241
rect 702 -3242 703 -3238
rect 702 -3307 703 -3241
rect 702 -3242 703 -3238
rect 702 -3307 703 -3241
rect 733 -3307 734 -3241
rect 814 -3242 815 -3238
rect 838 -3307 839 -3241
rect 1192 -3242 1193 -3238
rect 1199 -3307 1200 -3241
rect 1206 -3242 1207 -3238
rect 1227 -3242 1228 -3238
rect 1283 -3242 1284 -3238
rect 1293 -3242 1294 -3238
rect 1297 -3242 1298 -3238
rect 1346 -3242 1347 -3238
rect 1349 -3246 1350 -3241
rect 163 -3307 164 -3243
rect 366 -3244 367 -3238
rect 373 -3244 374 -3238
rect 373 -3307 374 -3243
rect 373 -3244 374 -3238
rect 373 -3307 374 -3243
rect 394 -3244 395 -3238
rect 544 -3244 545 -3238
rect 548 -3244 549 -3238
rect 576 -3307 577 -3243
rect 632 -3307 633 -3243
rect 681 -3244 682 -3238
rect 744 -3244 745 -3238
rect 1066 -3244 1067 -3238
rect 1101 -3244 1102 -3238
rect 1101 -3307 1102 -3243
rect 1101 -3244 1102 -3238
rect 1101 -3307 1102 -3243
rect 1136 -3244 1137 -3238
rect 1255 -3307 1256 -3243
rect 1346 -3307 1347 -3243
rect 1353 -3244 1354 -3238
rect 170 -3246 171 -3238
rect 481 -3246 482 -3238
rect 499 -3307 500 -3245
rect 747 -3246 748 -3238
rect 751 -3246 752 -3238
rect 772 -3246 773 -3238
rect 807 -3246 808 -3238
rect 1227 -3307 1228 -3245
rect 1241 -3246 1242 -3238
rect 1241 -3307 1242 -3245
rect 1241 -3246 1242 -3238
rect 1241 -3307 1242 -3245
rect 1353 -3307 1354 -3245
rect 170 -3307 171 -3247
rect 656 -3307 657 -3247
rect 667 -3248 668 -3238
rect 751 -3307 752 -3247
rect 758 -3248 759 -3238
rect 772 -3307 773 -3247
rect 807 -3307 808 -3247
rect 894 -3307 895 -3247
rect 933 -3248 934 -3238
rect 1066 -3307 1067 -3247
rect 1164 -3248 1165 -3238
rect 1234 -3248 1235 -3238
rect 177 -3250 178 -3238
rect 394 -3307 395 -3249
rect 408 -3250 409 -3238
rect 478 -3250 479 -3238
rect 527 -3250 528 -3238
rect 527 -3307 528 -3249
rect 527 -3250 528 -3238
rect 527 -3307 528 -3249
rect 541 -3250 542 -3238
rect 737 -3250 738 -3238
rect 758 -3307 759 -3249
rect 793 -3250 794 -3238
rect 810 -3250 811 -3238
rect 1038 -3250 1039 -3238
rect 1045 -3250 1046 -3238
rect 1258 -3250 1259 -3238
rect 177 -3307 178 -3251
rect 282 -3252 283 -3238
rect 289 -3252 290 -3238
rect 814 -3307 815 -3251
rect 863 -3252 864 -3238
rect 933 -3307 934 -3251
rect 947 -3252 948 -3238
rect 1038 -3307 1039 -3251
rect 1143 -3252 1144 -3238
rect 1164 -3307 1165 -3251
rect 1178 -3252 1179 -3238
rect 1206 -3307 1207 -3251
rect 1220 -3252 1221 -3238
rect 1234 -3307 1235 -3251
rect 187 -3254 188 -3238
rect 254 -3254 255 -3238
rect 268 -3254 269 -3238
rect 268 -3307 269 -3253
rect 268 -3254 269 -3238
rect 268 -3307 269 -3253
rect 282 -3307 283 -3253
rect 296 -3254 297 -3238
rect 317 -3254 318 -3238
rect 366 -3307 367 -3253
rect 408 -3307 409 -3253
rect 436 -3254 437 -3238
rect 450 -3254 451 -3238
rect 579 -3254 580 -3238
rect 618 -3254 619 -3238
rect 744 -3307 745 -3253
rect 765 -3307 766 -3253
rect 786 -3254 787 -3238
rect 793 -3307 794 -3253
rect 828 -3254 829 -3238
rect 863 -3307 864 -3253
rect 884 -3254 885 -3238
rect 891 -3254 892 -3238
rect 1003 -3254 1004 -3238
rect 1024 -3254 1025 -3238
rect 1192 -3307 1193 -3253
rect 1213 -3254 1214 -3238
rect 1220 -3307 1221 -3253
rect 198 -3256 199 -3238
rect 219 -3307 220 -3255
rect 247 -3256 248 -3238
rect 254 -3307 255 -3255
rect 296 -3307 297 -3255
rect 443 -3256 444 -3238
rect 450 -3307 451 -3255
rect 520 -3256 521 -3238
rect 541 -3307 542 -3255
rect 569 -3256 570 -3238
rect 618 -3307 619 -3255
rect 912 -3256 913 -3238
rect 947 -3307 948 -3255
rect 1087 -3256 1088 -3238
rect 1108 -3256 1109 -3238
rect 1143 -3307 1144 -3255
rect 1213 -3307 1214 -3255
rect 1248 -3256 1249 -3238
rect 205 -3258 206 -3238
rect 289 -3307 290 -3257
rect 303 -3258 304 -3238
rect 317 -3307 318 -3257
rect 324 -3307 325 -3257
rect 345 -3258 346 -3238
rect 352 -3307 353 -3257
rect 513 -3258 514 -3238
rect 548 -3307 549 -3257
rect 562 -3258 563 -3238
rect 709 -3307 710 -3257
rect 1024 -3307 1025 -3257
rect 1059 -3258 1060 -3238
rect 1108 -3307 1109 -3257
rect 205 -3307 206 -3259
rect 226 -3260 227 -3238
rect 247 -3307 248 -3259
rect 646 -3260 647 -3238
rect 737 -3307 738 -3259
rect 1272 -3307 1273 -3259
rect 198 -3307 199 -3261
rect 226 -3307 227 -3261
rect 303 -3307 304 -3261
rect 380 -3262 381 -3238
rect 387 -3262 388 -3238
rect 520 -3307 521 -3261
rect 562 -3307 563 -3261
rect 754 -3262 755 -3238
rect 768 -3262 769 -3238
rect 898 -3262 899 -3238
rect 912 -3307 913 -3261
rect 926 -3262 927 -3238
rect 954 -3262 955 -3238
rect 1178 -3307 1179 -3261
rect 191 -3264 192 -3238
rect 380 -3307 381 -3263
rect 387 -3307 388 -3263
rect 779 -3264 780 -3238
rect 786 -3307 787 -3263
rect 919 -3264 920 -3238
rect 954 -3307 955 -3263
rect 1136 -3307 1137 -3263
rect 191 -3307 192 -3265
rect 275 -3266 276 -3238
rect 331 -3266 332 -3238
rect 345 -3307 346 -3265
rect 415 -3266 416 -3238
rect 670 -3307 671 -3265
rect 779 -3307 780 -3265
rect 842 -3266 843 -3238
rect 870 -3266 871 -3238
rect 961 -3266 962 -3238
rect 964 -3266 965 -3238
rect 1185 -3266 1186 -3238
rect 275 -3307 276 -3267
rect 359 -3268 360 -3238
rect 415 -3307 416 -3267
rect 660 -3268 661 -3238
rect 800 -3268 801 -3238
rect 926 -3307 927 -3267
rect 996 -3268 997 -3238
rect 1045 -3307 1046 -3267
rect 1059 -3307 1060 -3267
rect 1073 -3268 1074 -3238
rect 1171 -3268 1172 -3238
rect 1185 -3307 1186 -3267
rect 331 -3307 332 -3269
rect 464 -3270 465 -3238
rect 478 -3307 479 -3269
rect 639 -3270 640 -3238
rect 646 -3307 647 -3269
rect 695 -3270 696 -3238
rect 828 -3307 829 -3269
rect 849 -3270 850 -3238
rect 856 -3270 857 -3238
rect 961 -3307 962 -3269
rect 996 -3307 997 -3269
rect 1031 -3270 1032 -3238
rect 1052 -3270 1053 -3238
rect 1073 -3307 1074 -3269
rect 1157 -3270 1158 -3238
rect 1171 -3307 1172 -3269
rect 184 -3272 185 -3238
rect 695 -3307 696 -3271
rect 842 -3307 843 -3271
rect 968 -3272 969 -3238
rect 982 -3272 983 -3238
rect 1031 -3307 1032 -3271
rect 1052 -3307 1053 -3271
rect 1150 -3272 1151 -3238
rect 184 -3307 185 -3273
rect 233 -3274 234 -3238
rect 310 -3274 311 -3238
rect 464 -3307 465 -3273
rect 485 -3274 486 -3238
rect 569 -3307 570 -3273
rect 614 -3307 615 -3273
rect 898 -3307 899 -3273
rect 919 -3307 920 -3273
rect 975 -3274 976 -3238
rect 982 -3307 983 -3273
rect 989 -3274 990 -3238
rect 1010 -3274 1011 -3238
rect 1248 -3307 1249 -3273
rect 233 -3307 234 -3275
rect 940 -3276 941 -3238
rect 968 -3307 969 -3275
rect 1122 -3276 1123 -3238
rect 1129 -3276 1130 -3238
rect 1150 -3307 1151 -3275
rect 310 -3307 311 -3277
rect 597 -3278 598 -3238
rect 625 -3278 626 -3238
rect 639 -3307 640 -3277
rect 660 -3307 661 -3277
rect 1129 -3307 1130 -3277
rect 359 -3307 360 -3279
rect 590 -3280 591 -3238
rect 625 -3307 626 -3279
rect 691 -3307 692 -3279
rect 821 -3280 822 -3238
rect 975 -3307 976 -3279
rect 989 -3307 990 -3279
rect 1202 -3280 1203 -3238
rect 422 -3282 423 -3238
rect 488 -3307 489 -3281
rect 513 -3307 514 -3281
rect 653 -3282 654 -3238
rect 667 -3307 668 -3281
rect 800 -3307 801 -3281
rect 884 -3307 885 -3281
rect 905 -3282 906 -3238
rect 940 -3307 941 -3281
rect 1003 -3307 1004 -3281
rect 1017 -3282 1018 -3238
rect 1087 -3307 1088 -3281
rect 1115 -3282 1116 -3238
rect 1122 -3307 1123 -3281
rect 422 -3307 423 -3283
rect 555 -3284 556 -3238
rect 583 -3284 584 -3238
rect 597 -3307 598 -3283
rect 653 -3307 654 -3283
rect 859 -3307 860 -3283
rect 877 -3284 878 -3238
rect 905 -3307 906 -3283
rect 1017 -3307 1018 -3283
rect 1080 -3284 1081 -3238
rect 1094 -3284 1095 -3238
rect 1115 -3307 1116 -3283
rect 429 -3286 430 -3238
rect 555 -3307 556 -3285
rect 583 -3307 584 -3285
rect 611 -3286 612 -3238
rect 681 -3307 682 -3285
rect 821 -3307 822 -3285
rect 877 -3307 878 -3285
rect 1262 -3286 1263 -3238
rect 429 -3307 430 -3287
rect 824 -3307 825 -3287
rect 1006 -3307 1007 -3287
rect 1080 -3307 1081 -3287
rect 1262 -3307 1263 -3287
rect 1276 -3288 1277 -3238
rect 436 -3307 437 -3289
rect 492 -3290 493 -3238
rect 534 -3290 535 -3238
rect 590 -3307 591 -3289
rect 611 -3307 612 -3289
rect 891 -3307 892 -3289
rect 1027 -3307 1028 -3289
rect 1157 -3307 1158 -3289
rect 1269 -3290 1270 -3238
rect 1276 -3307 1277 -3289
rect 261 -3292 262 -3238
rect 492 -3307 493 -3291
rect 688 -3292 689 -3238
rect 849 -3307 850 -3291
rect 261 -3307 262 -3293
rect 401 -3294 402 -3238
rect 443 -3307 444 -3293
rect 506 -3294 507 -3238
rect 688 -3307 689 -3293
rect 1010 -3307 1011 -3293
rect 338 -3296 339 -3238
rect 401 -3307 402 -3295
rect 457 -3296 458 -3238
rect 1094 -3307 1095 -3295
rect 338 -3307 339 -3297
rect 471 -3298 472 -3238
rect 485 -3307 486 -3297
rect 723 -3298 724 -3238
rect 457 -3307 458 -3299
rect 604 -3300 605 -3238
rect 716 -3300 717 -3238
rect 723 -3307 724 -3299
rect 471 -3307 472 -3301
rect 537 -3307 538 -3301
rect 604 -3307 605 -3301
rect 835 -3302 836 -3238
rect 506 -3307 507 -3303
rect 674 -3304 675 -3238
rect 716 -3307 717 -3303
rect 730 -3304 731 -3238
rect 674 -3307 675 -3305
rect 873 -3307 874 -3305
rect 156 -3317 157 -3315
rect 271 -3380 272 -3316
rect 303 -3317 304 -3315
rect 485 -3317 486 -3315
rect 520 -3317 521 -3315
rect 558 -3380 559 -3316
rect 576 -3317 577 -3315
rect 614 -3317 615 -3315
rect 646 -3317 647 -3315
rect 646 -3380 647 -3316
rect 646 -3317 647 -3315
rect 646 -3380 647 -3316
rect 653 -3317 654 -3315
rect 849 -3317 850 -3315
rect 856 -3317 857 -3315
rect 1143 -3317 1144 -3315
rect 1181 -3380 1182 -3316
rect 1262 -3317 1263 -3315
rect 1269 -3317 1270 -3315
rect 1290 -3317 1291 -3315
rect 1339 -3317 1340 -3315
rect 1339 -3380 1340 -3316
rect 1339 -3317 1340 -3315
rect 1339 -3380 1340 -3316
rect 1346 -3317 1347 -3315
rect 1346 -3380 1347 -3316
rect 1346 -3317 1347 -3315
rect 1346 -3380 1347 -3316
rect 1353 -3317 1354 -3315
rect 1353 -3380 1354 -3316
rect 1353 -3317 1354 -3315
rect 1353 -3380 1354 -3316
rect 163 -3319 164 -3315
rect 425 -3380 426 -3318
rect 436 -3319 437 -3315
rect 485 -3380 486 -3318
rect 544 -3380 545 -3318
rect 751 -3319 752 -3315
rect 761 -3319 762 -3315
rect 905 -3319 906 -3315
rect 1003 -3319 1004 -3315
rect 1073 -3319 1074 -3315
rect 1136 -3319 1137 -3315
rect 1241 -3319 1242 -3315
rect 1272 -3319 1273 -3315
rect 1276 -3319 1277 -3315
rect 177 -3321 178 -3315
rect 579 -3380 580 -3320
rect 611 -3380 612 -3320
rect 639 -3321 640 -3315
rect 660 -3321 661 -3315
rect 779 -3321 780 -3315
rect 786 -3321 787 -3315
rect 821 -3380 822 -3320
rect 824 -3321 825 -3315
rect 1066 -3321 1067 -3315
rect 1073 -3380 1074 -3320
rect 1150 -3321 1151 -3315
rect 184 -3323 185 -3315
rect 243 -3323 244 -3315
rect 254 -3323 255 -3315
rect 254 -3380 255 -3322
rect 254 -3323 255 -3315
rect 254 -3380 255 -3322
rect 261 -3323 262 -3315
rect 394 -3323 395 -3315
rect 411 -3380 412 -3322
rect 873 -3323 874 -3315
rect 891 -3323 892 -3315
rect 1031 -3323 1032 -3315
rect 1038 -3323 1039 -3315
rect 1041 -3380 1042 -3322
rect 1055 -3380 1056 -3322
rect 1087 -3323 1088 -3315
rect 1139 -3323 1140 -3315
rect 1157 -3323 1158 -3315
rect 198 -3380 199 -3324
rect 219 -3325 220 -3315
rect 226 -3325 227 -3315
rect 240 -3380 241 -3324
rect 282 -3325 283 -3315
rect 303 -3380 304 -3324
rect 359 -3325 360 -3315
rect 667 -3325 668 -3315
rect 670 -3325 671 -3315
rect 1178 -3325 1179 -3315
rect 205 -3327 206 -3315
rect 205 -3380 206 -3326
rect 205 -3327 206 -3315
rect 205 -3380 206 -3326
rect 212 -3327 213 -3315
rect 212 -3380 213 -3326
rect 212 -3327 213 -3315
rect 212 -3380 213 -3326
rect 226 -3380 227 -3326
rect 310 -3327 311 -3315
rect 387 -3327 388 -3315
rect 859 -3327 860 -3315
rect 870 -3327 871 -3315
rect 1192 -3327 1193 -3315
rect 275 -3329 276 -3315
rect 359 -3380 360 -3328
rect 387 -3380 388 -3328
rect 478 -3329 479 -3315
rect 513 -3329 514 -3315
rect 639 -3380 640 -3328
rect 660 -3380 661 -3328
rect 737 -3329 738 -3315
rect 751 -3380 752 -3328
rect 772 -3329 773 -3315
rect 779 -3380 780 -3328
rect 814 -3329 815 -3315
rect 828 -3329 829 -3315
rect 828 -3380 829 -3328
rect 828 -3329 829 -3315
rect 828 -3380 829 -3328
rect 835 -3329 836 -3315
rect 1248 -3329 1249 -3315
rect 275 -3380 276 -3330
rect 345 -3331 346 -3315
rect 394 -3380 395 -3330
rect 506 -3331 507 -3315
rect 513 -3380 514 -3330
rect 653 -3380 654 -3330
rect 667 -3380 668 -3330
rect 723 -3331 724 -3315
rect 737 -3380 738 -3330
rect 765 -3331 766 -3315
rect 807 -3331 808 -3315
rect 814 -3380 815 -3330
rect 835 -3380 836 -3330
rect 926 -3331 927 -3315
rect 947 -3331 948 -3315
rect 1087 -3380 1088 -3330
rect 1192 -3380 1193 -3330
rect 1213 -3331 1214 -3315
rect 282 -3380 283 -3332
rect 296 -3333 297 -3315
rect 310 -3380 311 -3332
rect 317 -3333 318 -3315
rect 345 -3380 346 -3332
rect 373 -3333 374 -3315
rect 422 -3333 423 -3315
rect 537 -3333 538 -3315
rect 569 -3333 570 -3315
rect 772 -3380 773 -3332
rect 838 -3333 839 -3315
rect 1115 -3333 1116 -3315
rect 219 -3380 220 -3334
rect 569 -3380 570 -3334
rect 572 -3380 573 -3334
rect 723 -3380 724 -3334
rect 761 -3380 762 -3334
rect 1045 -3335 1046 -3315
rect 296 -3380 297 -3336
rect 324 -3337 325 -3315
rect 373 -3380 374 -3336
rect 401 -3337 402 -3315
rect 436 -3380 437 -3336
rect 464 -3337 465 -3315
rect 478 -3380 479 -3336
rect 541 -3337 542 -3315
rect 632 -3337 633 -3315
rect 807 -3380 808 -3336
rect 842 -3337 843 -3315
rect 842 -3380 843 -3336
rect 842 -3337 843 -3315
rect 842 -3380 843 -3336
rect 849 -3380 850 -3336
rect 961 -3337 962 -3315
rect 1003 -3380 1004 -3336
rect 1052 -3337 1053 -3315
rect 317 -3380 318 -3338
rect 408 -3339 409 -3315
rect 506 -3380 507 -3338
rect 541 -3380 542 -3338
rect 632 -3380 633 -3338
rect 730 -3339 731 -3315
rect 765 -3380 766 -3338
rect 793 -3339 794 -3315
rect 856 -3380 857 -3338
rect 940 -3339 941 -3315
rect 947 -3380 948 -3338
rect 968 -3339 969 -3315
rect 1024 -3380 1025 -3338
rect 1234 -3339 1235 -3315
rect 324 -3380 325 -3340
rect 471 -3341 472 -3315
rect 534 -3341 535 -3315
rect 786 -3380 787 -3340
rect 870 -3380 871 -3340
rect 1094 -3341 1095 -3315
rect 170 -3343 171 -3315
rect 471 -3380 472 -3342
rect 534 -3380 535 -3342
rect 548 -3343 549 -3315
rect 681 -3343 682 -3315
rect 968 -3380 969 -3342
rect 1027 -3343 1028 -3315
rect 1185 -3343 1186 -3315
rect 331 -3345 332 -3315
rect 793 -3380 794 -3344
rect 884 -3345 885 -3315
rect 1031 -3380 1032 -3344
rect 1045 -3380 1046 -3344
rect 1108 -3345 1109 -3315
rect 1185 -3380 1186 -3344
rect 1199 -3345 1200 -3315
rect 331 -3380 332 -3346
rect 443 -3347 444 -3315
rect 548 -3380 549 -3346
rect 625 -3347 626 -3315
rect 688 -3347 689 -3315
rect 702 -3347 703 -3315
rect 730 -3380 731 -3346
rect 744 -3347 745 -3315
rect 884 -3380 885 -3346
rect 1010 -3347 1011 -3315
rect 1052 -3380 1053 -3346
rect 1255 -3347 1256 -3315
rect 380 -3349 381 -3315
rect 401 -3380 402 -3348
rect 408 -3380 409 -3348
rect 464 -3380 465 -3348
rect 492 -3349 493 -3315
rect 625 -3380 626 -3348
rect 702 -3380 703 -3348
rect 716 -3349 717 -3315
rect 744 -3380 745 -3348
rect 877 -3349 878 -3315
rect 891 -3380 892 -3348
rect 912 -3349 913 -3315
rect 926 -3380 927 -3348
rect 1227 -3349 1228 -3315
rect 380 -3380 381 -3350
rect 499 -3351 500 -3315
rect 597 -3351 598 -3315
rect 681 -3380 682 -3350
rect 691 -3351 692 -3315
rect 716 -3380 717 -3350
rect 877 -3380 878 -3350
rect 982 -3351 983 -3315
rect 1094 -3380 1095 -3350
rect 1122 -3351 1123 -3315
rect 443 -3380 444 -3352
rect 527 -3353 528 -3315
rect 618 -3353 619 -3315
rect 688 -3380 689 -3352
rect 894 -3353 895 -3315
rect 933 -3353 934 -3315
rect 940 -3380 941 -3352
rect 1080 -3353 1081 -3315
rect 1122 -3380 1123 -3352
rect 1220 -3353 1221 -3315
rect 450 -3355 451 -3315
rect 499 -3380 500 -3354
rect 527 -3380 528 -3354
rect 663 -3355 664 -3315
rect 898 -3355 899 -3315
rect 1069 -3380 1070 -3354
rect 1080 -3380 1081 -3354
rect 1101 -3355 1102 -3315
rect 233 -3357 234 -3315
rect 450 -3380 451 -3356
rect 457 -3357 458 -3315
rect 597 -3380 598 -3356
rect 898 -3380 899 -3356
rect 954 -3357 955 -3315
rect 961 -3380 962 -3356
rect 1206 -3357 1207 -3315
rect 233 -3380 234 -3358
rect 338 -3359 339 -3315
rect 422 -3380 423 -3358
rect 457 -3380 458 -3358
rect 492 -3380 493 -3358
rect 604 -3359 605 -3315
rect 758 -3359 759 -3315
rect 954 -3380 955 -3358
rect 975 -3359 976 -3315
rect 1010 -3380 1011 -3358
rect 1017 -3359 1018 -3315
rect 1101 -3380 1102 -3358
rect 338 -3380 339 -3360
rect 562 -3361 563 -3315
rect 576 -3380 577 -3360
rect 604 -3380 605 -3360
rect 674 -3361 675 -3315
rect 975 -3380 976 -3360
rect 982 -3380 983 -3360
rect 1171 -3361 1172 -3315
rect 247 -3363 248 -3315
rect 674 -3380 675 -3362
rect 905 -3380 906 -3362
rect 919 -3363 920 -3315
rect 933 -3380 934 -3362
rect 989 -3363 990 -3315
rect 1013 -3380 1014 -3362
rect 1017 -3380 1018 -3362
rect 191 -3365 192 -3315
rect 247 -3380 248 -3364
rect 352 -3365 353 -3315
rect 562 -3380 563 -3364
rect 583 -3365 584 -3315
rect 618 -3380 619 -3364
rect 912 -3380 913 -3364
rect 996 -3365 997 -3315
rect 352 -3380 353 -3366
rect 555 -3367 556 -3315
rect 583 -3380 584 -3366
rect 709 -3367 710 -3315
rect 800 -3367 801 -3315
rect 996 -3380 997 -3366
rect 415 -3369 416 -3315
rect 555 -3380 556 -3368
rect 590 -3369 591 -3315
rect 709 -3380 710 -3368
rect 800 -3380 801 -3368
rect 863 -3369 864 -3315
rect 919 -3380 920 -3368
rect 1066 -3380 1067 -3368
rect 404 -3380 405 -3370
rect 590 -3380 591 -3370
rect 695 -3371 696 -3315
rect 863 -3380 864 -3370
rect 989 -3380 990 -3370
rect 1059 -3371 1060 -3315
rect 415 -3380 416 -3372
rect 429 -3373 430 -3315
rect 656 -3373 657 -3315
rect 695 -3380 696 -3372
rect 1059 -3380 1060 -3372
rect 1129 -3373 1130 -3315
rect 366 -3375 367 -3315
rect 429 -3380 430 -3374
rect 520 -3380 521 -3374
rect 656 -3380 657 -3374
rect 1129 -3380 1130 -3374
rect 1164 -3375 1165 -3315
rect 289 -3377 290 -3315
rect 366 -3380 367 -3376
rect 268 -3379 269 -3315
rect 289 -3380 290 -3378
rect 198 -3390 199 -3388
rect 292 -3443 293 -3389
rect 296 -3390 297 -3388
rect 446 -3443 447 -3389
rect 457 -3390 458 -3388
rect 460 -3408 461 -3389
rect 492 -3390 493 -3388
rect 656 -3390 657 -3388
rect 681 -3390 682 -3388
rect 681 -3443 682 -3389
rect 681 -3390 682 -3388
rect 681 -3443 682 -3389
rect 723 -3390 724 -3388
rect 758 -3390 759 -3388
rect 793 -3390 794 -3388
rect 870 -3390 871 -3388
rect 1003 -3390 1004 -3388
rect 1003 -3443 1004 -3389
rect 1003 -3390 1004 -3388
rect 1003 -3443 1004 -3389
rect 1013 -3390 1014 -3388
rect 1087 -3390 1088 -3388
rect 1101 -3390 1102 -3388
rect 1136 -3443 1137 -3389
rect 1178 -3443 1179 -3389
rect 1185 -3390 1186 -3388
rect 1339 -3390 1340 -3388
rect 1339 -3443 1340 -3389
rect 1339 -3390 1340 -3388
rect 1339 -3443 1340 -3389
rect 1346 -3390 1347 -3388
rect 1349 -3390 1350 -3388
rect 205 -3392 206 -3388
rect 278 -3392 279 -3388
rect 317 -3392 318 -3388
rect 408 -3392 409 -3388
rect 422 -3392 423 -3388
rect 723 -3443 724 -3391
rect 737 -3392 738 -3388
rect 793 -3443 794 -3391
rect 807 -3392 808 -3388
rect 810 -3408 811 -3391
rect 824 -3443 825 -3391
rect 898 -3392 899 -3388
rect 1027 -3443 1028 -3391
rect 1122 -3392 1123 -3388
rect 1181 -3392 1182 -3388
rect 1192 -3392 1193 -3388
rect 1346 -3443 1347 -3391
rect 1353 -3392 1354 -3388
rect 212 -3394 213 -3388
rect 268 -3394 269 -3388
rect 271 -3394 272 -3388
rect 691 -3443 692 -3393
rect 737 -3443 738 -3393
rect 975 -3394 976 -3388
rect 1066 -3394 1067 -3388
rect 1080 -3394 1081 -3388
rect 1087 -3443 1088 -3393
rect 1094 -3394 1095 -3388
rect 1115 -3443 1116 -3393
rect 1129 -3394 1130 -3388
rect 219 -3396 220 -3388
rect 502 -3443 503 -3395
rect 530 -3443 531 -3395
rect 576 -3396 577 -3388
rect 579 -3396 580 -3388
rect 646 -3396 647 -3388
rect 649 -3443 650 -3395
rect 961 -3396 962 -3388
rect 1010 -3396 1011 -3388
rect 1094 -3443 1095 -3395
rect 247 -3398 248 -3388
rect 474 -3398 475 -3388
rect 555 -3443 556 -3397
rect 590 -3398 591 -3388
rect 597 -3398 598 -3388
rect 646 -3443 647 -3397
rect 653 -3443 654 -3397
rect 996 -3398 997 -3388
rect 1010 -3443 1011 -3397
rect 1045 -3398 1046 -3388
rect 240 -3400 241 -3388
rect 247 -3443 248 -3399
rect 261 -3400 262 -3388
rect 289 -3400 290 -3388
rect 324 -3400 325 -3388
rect 348 -3443 349 -3399
rect 366 -3400 367 -3388
rect 404 -3400 405 -3388
rect 408 -3443 409 -3399
rect 429 -3400 430 -3388
rect 450 -3400 451 -3388
rect 492 -3443 493 -3399
rect 558 -3400 559 -3388
rect 590 -3443 591 -3399
rect 667 -3400 668 -3388
rect 758 -3443 759 -3399
rect 807 -3443 808 -3399
rect 877 -3400 878 -3388
rect 933 -3400 934 -3388
rect 975 -3443 976 -3399
rect 1031 -3400 1032 -3388
rect 1045 -3443 1046 -3399
rect 226 -3402 227 -3388
rect 366 -3443 367 -3401
rect 387 -3402 388 -3388
rect 429 -3443 430 -3401
rect 450 -3443 451 -3401
rect 611 -3402 612 -3388
rect 667 -3443 668 -3401
rect 786 -3402 787 -3388
rect 859 -3443 860 -3401
rect 873 -3443 874 -3401
rect 877 -3443 878 -3401
rect 891 -3402 892 -3388
rect 961 -3443 962 -3401
rect 1024 -3402 1025 -3388
rect 1031 -3443 1032 -3401
rect 1059 -3402 1060 -3388
rect 254 -3404 255 -3388
rect 261 -3443 262 -3403
rect 282 -3404 283 -3388
rect 317 -3443 318 -3403
rect 359 -3404 360 -3388
rect 387 -3443 388 -3403
rect 401 -3443 402 -3403
rect 478 -3404 479 -3388
rect 485 -3404 486 -3388
rect 597 -3443 598 -3403
rect 716 -3404 717 -3388
rect 933 -3443 934 -3403
rect 968 -3404 969 -3388
rect 1024 -3443 1025 -3403
rect 303 -3406 304 -3388
rect 324 -3443 325 -3405
rect 345 -3406 346 -3388
rect 359 -3443 360 -3405
rect 415 -3406 416 -3388
rect 422 -3443 423 -3405
rect 457 -3443 458 -3405
rect 548 -3406 549 -3388
rect 611 -3443 612 -3405
rect 716 -3443 717 -3405
rect 772 -3406 773 -3388
rect 786 -3443 787 -3405
rect 800 -3406 801 -3388
rect 863 -3406 864 -3388
rect 887 -3443 888 -3405
rect 968 -3443 969 -3405
rect 989 -3406 990 -3388
rect 233 -3408 234 -3388
rect 345 -3443 346 -3407
rect 373 -3408 374 -3388
rect 415 -3443 416 -3407
rect 478 -3443 479 -3407
rect 506 -3408 507 -3388
rect 541 -3408 542 -3388
rect 548 -3443 549 -3407
rect 569 -3408 570 -3388
rect 618 -3408 619 -3388
rect 660 -3408 661 -3388
rect 772 -3443 773 -3407
rect 800 -3443 801 -3407
rect 814 -3408 815 -3388
rect 863 -3443 864 -3407
rect 919 -3408 920 -3388
rect 1349 -3443 1350 -3407
rect 1353 -3443 1354 -3407
rect 373 -3443 374 -3409
rect 796 -3410 797 -3388
rect 919 -3443 920 -3409
rect 947 -3410 948 -3388
rect 394 -3412 395 -3388
rect 569 -3443 570 -3411
rect 572 -3412 573 -3388
rect 957 -3412 958 -3388
rect 338 -3414 339 -3388
rect 394 -3443 395 -3413
rect 485 -3443 486 -3413
rect 499 -3414 500 -3388
rect 506 -3443 507 -3413
rect 604 -3414 605 -3388
rect 618 -3443 619 -3413
rect 695 -3414 696 -3388
rect 940 -3414 941 -3388
rect 947 -3443 948 -3413
rect 310 -3416 311 -3388
rect 338 -3443 339 -3415
rect 436 -3416 437 -3388
rect 604 -3443 605 -3415
rect 632 -3416 633 -3388
rect 695 -3443 696 -3415
rect 905 -3416 906 -3388
rect 940 -3443 941 -3415
rect 310 -3443 311 -3417
rect 331 -3418 332 -3388
rect 380 -3418 381 -3388
rect 436 -3443 437 -3417
rect 499 -3443 500 -3417
rect 779 -3418 780 -3388
rect 856 -3418 857 -3388
rect 905 -3443 906 -3417
rect 331 -3443 332 -3419
rect 513 -3420 514 -3388
rect 541 -3443 542 -3419
rect 639 -3420 640 -3388
rect 674 -3420 675 -3388
rect 814 -3443 815 -3419
rect 380 -3443 381 -3421
rect 464 -3422 465 -3388
rect 513 -3443 514 -3421
rect 520 -3422 521 -3388
rect 562 -3422 563 -3388
rect 660 -3443 661 -3421
rect 674 -3443 675 -3421
rect 751 -3422 752 -3388
rect 352 -3424 353 -3388
rect 562 -3443 563 -3423
rect 576 -3443 577 -3423
rect 625 -3424 626 -3388
rect 632 -3443 633 -3423
rect 835 -3424 836 -3388
rect 352 -3443 353 -3425
rect 411 -3426 412 -3388
rect 443 -3426 444 -3388
rect 520 -3443 521 -3425
rect 625 -3443 626 -3425
rect 709 -3426 710 -3388
rect 835 -3443 836 -3425
rect 842 -3426 843 -3388
rect 464 -3443 465 -3427
rect 471 -3428 472 -3388
rect 639 -3443 640 -3427
rect 765 -3428 766 -3388
rect 842 -3443 843 -3427
rect 926 -3428 927 -3388
rect 471 -3443 472 -3429
rect 534 -3430 535 -3388
rect 688 -3430 689 -3388
rect 779 -3443 780 -3429
rect 912 -3430 913 -3388
rect 926 -3443 927 -3429
rect 534 -3443 535 -3431
rect 583 -3432 584 -3388
rect 702 -3432 703 -3388
rect 751 -3443 752 -3431
rect 765 -3443 766 -3431
rect 828 -3432 829 -3388
rect 912 -3443 913 -3431
rect 982 -3432 983 -3388
rect 583 -3443 584 -3433
rect 744 -3434 745 -3388
rect 828 -3443 829 -3433
rect 884 -3434 885 -3388
rect 982 -3443 983 -3433
rect 1038 -3434 1039 -3388
rect 702 -3443 703 -3435
rect 730 -3436 731 -3388
rect 744 -3443 745 -3435
rect 1017 -3436 1018 -3388
rect 1038 -3443 1039 -3435
rect 1073 -3436 1074 -3388
rect 709 -3443 710 -3437
rect 821 -3438 822 -3388
rect 884 -3443 885 -3437
rect 954 -3443 955 -3437
rect 730 -3443 731 -3439
rect 849 -3440 850 -3388
rect 740 -3443 741 -3441
rect 849 -3443 850 -3441
rect 247 -3453 248 -3451
rect 247 -3500 248 -3452
rect 247 -3453 248 -3451
rect 247 -3500 248 -3452
rect 261 -3453 262 -3451
rect 261 -3500 262 -3452
rect 261 -3453 262 -3451
rect 261 -3500 262 -3452
rect 275 -3500 276 -3452
rect 289 -3453 290 -3451
rect 292 -3453 293 -3451
rect 310 -3453 311 -3451
rect 331 -3453 332 -3451
rect 366 -3500 367 -3452
rect 380 -3453 381 -3451
rect 383 -3469 384 -3452
rect 464 -3453 465 -3451
rect 467 -3500 468 -3452
rect 513 -3453 514 -3451
rect 579 -3500 580 -3452
rect 611 -3453 612 -3451
rect 649 -3453 650 -3451
rect 677 -3500 678 -3452
rect 957 -3500 958 -3452
rect 989 -3500 990 -3452
rect 1010 -3453 1011 -3451
rect 1045 -3453 1046 -3451
rect 1052 -3500 1053 -3452
rect 1080 -3500 1081 -3452
rect 1087 -3453 1088 -3451
rect 1094 -3453 1095 -3451
rect 1122 -3500 1123 -3452
rect 1136 -3453 1137 -3451
rect 1150 -3500 1151 -3452
rect 1178 -3453 1179 -3451
rect 1178 -3500 1179 -3452
rect 1178 -3453 1179 -3451
rect 1178 -3500 1179 -3452
rect 1339 -3453 1340 -3451
rect 1342 -3453 1343 -3451
rect 317 -3455 318 -3451
rect 331 -3500 332 -3454
rect 338 -3455 339 -3451
rect 345 -3500 346 -3454
rect 359 -3455 360 -3451
rect 362 -3469 363 -3454
rect 380 -3500 381 -3454
rect 436 -3455 437 -3451
rect 513 -3500 514 -3454
rect 534 -3455 535 -3451
rect 611 -3500 612 -3454
rect 667 -3455 668 -3451
rect 688 -3455 689 -3451
rect 702 -3455 703 -3451
rect 726 -3500 727 -3454
rect 807 -3455 808 -3451
rect 817 -3500 818 -3454
rect 863 -3455 864 -3451
rect 870 -3455 871 -3451
rect 884 -3455 885 -3451
rect 898 -3455 899 -3451
rect 982 -3455 983 -3451
rect 996 -3500 997 -3454
rect 1038 -3455 1039 -3451
rect 1087 -3500 1088 -3454
rect 1171 -3500 1172 -3454
rect 1339 -3500 1340 -3454
rect 1346 -3455 1347 -3451
rect 324 -3457 325 -3451
rect 338 -3500 339 -3456
rect 359 -3500 360 -3456
rect 408 -3457 409 -3451
rect 464 -3500 465 -3456
rect 478 -3457 479 -3451
rect 534 -3500 535 -3456
rect 604 -3457 605 -3451
rect 667 -3500 668 -3456
rect 681 -3457 682 -3451
rect 688 -3500 689 -3456
rect 691 -3457 692 -3451
rect 842 -3457 843 -3451
rect 849 -3457 850 -3451
rect 901 -3457 902 -3451
rect 905 -3457 906 -3451
rect 999 -3500 1000 -3456
rect 1003 -3457 1004 -3451
rect 1003 -3500 1004 -3456
rect 1003 -3457 1004 -3451
rect 1003 -3500 1004 -3456
rect 1010 -3500 1011 -3456
rect 1031 -3457 1032 -3451
rect 1108 -3500 1109 -3456
rect 1115 -3457 1116 -3451
rect 1346 -3500 1347 -3456
rect 1353 -3457 1354 -3451
rect 408 -3500 409 -3458
rect 450 -3459 451 -3451
rect 478 -3500 479 -3458
rect 548 -3459 549 -3451
rect 597 -3459 598 -3451
rect 604 -3500 605 -3458
rect 628 -3500 629 -3458
rect 1027 -3459 1028 -3451
rect 422 -3461 423 -3451
rect 450 -3500 451 -3460
rect 499 -3461 500 -3451
rect 548 -3500 549 -3460
rect 562 -3461 563 -3451
rect 597 -3500 598 -3460
rect 646 -3500 647 -3460
rect 737 -3461 738 -3451
rect 744 -3461 745 -3451
rect 744 -3500 745 -3460
rect 744 -3461 745 -3451
rect 744 -3500 745 -3460
rect 751 -3461 752 -3451
rect 754 -3469 755 -3460
rect 765 -3461 766 -3451
rect 765 -3500 766 -3460
rect 765 -3461 766 -3451
rect 765 -3500 766 -3460
rect 779 -3461 780 -3451
rect 863 -3500 864 -3460
rect 877 -3461 878 -3451
rect 887 -3461 888 -3451
rect 905 -3500 906 -3460
rect 912 -3461 913 -3451
rect 919 -3461 920 -3451
rect 919 -3500 920 -3460
rect 919 -3461 920 -3451
rect 919 -3500 920 -3460
rect 926 -3461 927 -3451
rect 929 -3469 930 -3460
rect 933 -3461 934 -3451
rect 936 -3461 937 -3451
rect 940 -3461 941 -3451
rect 943 -3461 944 -3451
rect 954 -3461 955 -3451
rect 982 -3500 983 -3460
rect 436 -3500 437 -3462
rect 471 -3463 472 -3451
rect 520 -3463 521 -3451
rect 583 -3463 584 -3451
rect 653 -3463 654 -3451
rect 702 -3500 703 -3462
rect 751 -3500 752 -3462
rect 779 -3500 780 -3462
rect 824 -3463 825 -3451
rect 835 -3463 836 -3451
rect 856 -3463 857 -3451
rect 891 -3463 892 -3451
rect 912 -3500 913 -3462
rect 926 -3500 927 -3462
rect 968 -3463 969 -3451
rect 471 -3500 472 -3464
rect 527 -3465 528 -3451
rect 576 -3465 577 -3451
rect 590 -3465 591 -3451
rect 653 -3500 654 -3464
rect 660 -3465 661 -3451
rect 681 -3500 682 -3464
rect 695 -3465 696 -3451
rect 740 -3465 741 -3451
rect 772 -3465 773 -3451
rect 835 -3500 836 -3464
rect 933 -3500 934 -3464
rect 961 -3465 962 -3451
rect 425 -3500 426 -3466
rect 520 -3500 521 -3466
rect 530 -3467 531 -3451
rect 660 -3500 661 -3466
rect 674 -3467 675 -3451
rect 737 -3500 738 -3466
rect 772 -3500 773 -3466
rect 859 -3467 860 -3451
rect 940 -3500 941 -3466
rect 947 -3467 948 -3451
rect 954 -3500 955 -3466
rect 975 -3467 976 -3451
rect 443 -3469 444 -3451
rect 590 -3500 591 -3468
rect 786 -3469 787 -3451
rect 870 -3500 871 -3468
rect 1342 -3500 1343 -3468
rect 1353 -3500 1354 -3468
rect 443 -3500 444 -3470
rect 457 -3471 458 -3451
rect 506 -3471 507 -3451
rect 527 -3500 528 -3470
rect 562 -3500 563 -3470
rect 618 -3471 619 -3451
rect 793 -3471 794 -3451
rect 821 -3471 822 -3451
rect 828 -3471 829 -3451
rect 856 -3500 857 -3470
rect 422 -3500 423 -3472
rect 506 -3500 507 -3472
rect 618 -3500 619 -3472
rect 625 -3473 626 -3451
rect 723 -3473 724 -3451
rect 821 -3500 822 -3472
rect 446 -3475 447 -3451
rect 499 -3500 500 -3474
rect 583 -3500 584 -3474
rect 625 -3500 626 -3474
rect 800 -3475 801 -3451
rect 842 -3500 843 -3474
rect 457 -3500 458 -3476
rect 485 -3477 486 -3451
rect 709 -3477 710 -3451
rect 800 -3500 801 -3476
rect 807 -3500 808 -3476
rect 1174 -3500 1175 -3476
rect 485 -3500 486 -3478
rect 541 -3479 542 -3451
rect 709 -3500 710 -3478
rect 730 -3479 731 -3451
rect 814 -3479 815 -3451
rect 877 -3500 878 -3478
rect 541 -3500 542 -3480
rect 569 -3481 570 -3451
rect 695 -3500 696 -3480
rect 814 -3500 815 -3480
rect 569 -3500 570 -3482
rect 632 -3483 633 -3451
rect 716 -3483 717 -3451
rect 730 -3500 731 -3482
rect 555 -3485 556 -3451
rect 632 -3500 633 -3484
rect 639 -3485 640 -3451
rect 716 -3500 717 -3484
rect 492 -3487 493 -3451
rect 555 -3500 556 -3486
rect 639 -3500 640 -3486
rect 849 -3500 850 -3486
rect 429 -3489 430 -3451
rect 492 -3500 493 -3488
rect 394 -3491 395 -3451
rect 429 -3500 430 -3490
rect 352 -3493 353 -3451
rect 394 -3500 395 -3492
rect 352 -3500 353 -3494
rect 373 -3495 374 -3451
rect 373 -3500 374 -3496
rect 415 -3497 416 -3451
rect 415 -3500 416 -3498
rect 537 -3500 538 -3498
rect 247 -3510 248 -3508
rect 247 -3541 248 -3509
rect 247 -3510 248 -3508
rect 247 -3541 248 -3509
rect 254 -3541 255 -3509
rect 296 -3541 297 -3509
rect 352 -3510 353 -3508
rect 534 -3510 535 -3508
rect 555 -3510 556 -3508
rect 625 -3510 626 -3508
rect 639 -3510 640 -3508
rect 688 -3510 689 -3508
rect 691 -3541 692 -3509
rect 772 -3510 773 -3508
rect 821 -3510 822 -3508
rect 922 -3541 923 -3509
rect 940 -3510 941 -3508
rect 940 -3541 941 -3509
rect 940 -3510 941 -3508
rect 940 -3541 941 -3509
rect 947 -3510 948 -3508
rect 954 -3510 955 -3508
rect 968 -3510 969 -3508
rect 975 -3541 976 -3509
rect 982 -3510 983 -3508
rect 1006 -3541 1007 -3509
rect 1052 -3510 1053 -3508
rect 1052 -3541 1053 -3509
rect 1052 -3510 1053 -3508
rect 1052 -3541 1053 -3509
rect 1059 -3541 1060 -3509
rect 1087 -3510 1088 -3508
rect 1108 -3510 1109 -3508
rect 1108 -3541 1109 -3509
rect 1108 -3510 1109 -3508
rect 1108 -3541 1109 -3509
rect 1122 -3510 1123 -3508
rect 1160 -3541 1161 -3509
rect 1171 -3510 1172 -3508
rect 1178 -3510 1179 -3508
rect 1339 -3510 1340 -3508
rect 1349 -3510 1350 -3508
rect 261 -3512 262 -3508
rect 261 -3541 262 -3511
rect 261 -3512 262 -3508
rect 261 -3541 262 -3511
rect 268 -3541 269 -3511
rect 275 -3512 276 -3508
rect 401 -3512 402 -3508
rect 425 -3512 426 -3508
rect 429 -3512 430 -3508
rect 562 -3512 563 -3508
rect 576 -3512 577 -3508
rect 604 -3512 605 -3508
rect 611 -3512 612 -3508
rect 611 -3541 612 -3511
rect 611 -3512 612 -3508
rect 611 -3541 612 -3511
rect 618 -3512 619 -3508
rect 625 -3541 626 -3511
rect 653 -3512 654 -3508
rect 688 -3541 689 -3511
rect 702 -3512 703 -3508
rect 702 -3541 703 -3511
rect 702 -3512 703 -3508
rect 702 -3541 703 -3511
rect 709 -3512 710 -3508
rect 709 -3541 710 -3511
rect 709 -3512 710 -3508
rect 709 -3541 710 -3511
rect 730 -3512 731 -3508
rect 733 -3520 734 -3511
rect 751 -3512 752 -3508
rect 751 -3541 752 -3511
rect 751 -3512 752 -3508
rect 751 -3541 752 -3511
rect 758 -3512 759 -3508
rect 758 -3541 759 -3511
rect 758 -3512 759 -3508
rect 758 -3541 759 -3511
rect 765 -3512 766 -3508
rect 765 -3541 766 -3511
rect 765 -3512 766 -3508
rect 765 -3541 766 -3511
rect 849 -3512 850 -3508
rect 898 -3541 899 -3511
rect 905 -3512 906 -3508
rect 905 -3541 906 -3511
rect 905 -3512 906 -3508
rect 905 -3541 906 -3511
rect 933 -3512 934 -3508
rect 947 -3541 948 -3511
rect 961 -3512 962 -3508
rect 968 -3541 969 -3511
rect 989 -3512 990 -3508
rect 989 -3541 990 -3511
rect 989 -3512 990 -3508
rect 989 -3541 990 -3511
rect 996 -3512 997 -3508
rect 1010 -3512 1011 -3508
rect 1080 -3512 1081 -3508
rect 1080 -3541 1081 -3511
rect 1080 -3512 1081 -3508
rect 1080 -3541 1081 -3511
rect 1150 -3512 1151 -3508
rect 1150 -3541 1151 -3511
rect 1150 -3512 1151 -3508
rect 1150 -3541 1151 -3511
rect 1346 -3512 1347 -3508
rect 1353 -3512 1354 -3508
rect 387 -3514 388 -3508
rect 401 -3541 402 -3513
rect 422 -3514 423 -3508
rect 478 -3514 479 -3508
rect 495 -3514 496 -3508
rect 642 -3514 643 -3508
rect 660 -3514 661 -3508
rect 723 -3541 724 -3513
rect 730 -3541 731 -3513
rect 744 -3514 745 -3508
rect 842 -3514 843 -3508
rect 849 -3541 850 -3513
rect 870 -3514 871 -3508
rect 884 -3541 885 -3513
rect 912 -3514 913 -3508
rect 933 -3541 934 -3513
rect 1003 -3514 1004 -3508
rect 1010 -3541 1011 -3513
rect 373 -3516 374 -3508
rect 422 -3541 423 -3515
rect 429 -3541 430 -3515
rect 604 -3541 605 -3515
rect 667 -3516 668 -3508
rect 726 -3516 727 -3508
rect 737 -3516 738 -3508
rect 744 -3541 745 -3515
rect 856 -3516 857 -3508
rect 870 -3541 871 -3515
rect 877 -3516 878 -3508
rect 891 -3541 892 -3515
rect 912 -3541 913 -3515
rect 926 -3516 927 -3508
rect 450 -3518 451 -3508
rect 492 -3518 493 -3508
rect 499 -3518 500 -3508
rect 534 -3541 535 -3517
rect 548 -3518 549 -3508
rect 576 -3541 577 -3517
rect 590 -3518 591 -3508
rect 639 -3541 640 -3517
rect 667 -3541 668 -3517
rect 807 -3518 808 -3508
rect 863 -3518 864 -3508
rect 877 -3541 878 -3517
rect 919 -3518 920 -3508
rect 926 -3541 927 -3517
rect 394 -3520 395 -3508
rect 450 -3541 451 -3519
rect 453 -3541 454 -3519
rect 478 -3541 479 -3519
rect 485 -3520 486 -3508
rect 492 -3541 493 -3519
rect 499 -3541 500 -3519
rect 565 -3520 566 -3508
rect 597 -3520 598 -3508
rect 628 -3541 629 -3519
rect 674 -3520 675 -3508
rect 681 -3520 682 -3508
rect 737 -3541 738 -3519
rect 835 -3520 836 -3508
rect 863 -3541 864 -3519
rect 359 -3522 360 -3508
rect 394 -3541 395 -3521
rect 457 -3522 458 -3508
rect 548 -3541 549 -3521
rect 555 -3541 556 -3521
rect 569 -3522 570 -3508
rect 600 -3541 601 -3521
rect 646 -3522 647 -3508
rect 677 -3522 678 -3508
rect 943 -3541 944 -3521
rect 338 -3524 339 -3508
rect 359 -3541 360 -3523
rect 408 -3524 409 -3508
rect 457 -3541 458 -3523
rect 471 -3524 472 -3508
rect 471 -3541 472 -3523
rect 471 -3524 472 -3508
rect 471 -3541 472 -3523
rect 506 -3524 507 -3508
rect 506 -3541 507 -3523
rect 506 -3524 507 -3508
rect 506 -3541 507 -3523
rect 513 -3524 514 -3508
rect 562 -3541 563 -3523
rect 569 -3541 570 -3523
rect 583 -3524 584 -3508
rect 632 -3524 633 -3508
rect 681 -3541 682 -3523
rect 800 -3524 801 -3508
rect 835 -3541 836 -3523
rect 408 -3541 409 -3525
rect 464 -3526 465 -3508
rect 467 -3526 468 -3508
rect 583 -3541 584 -3525
rect 443 -3528 444 -3508
rect 513 -3541 514 -3527
rect 520 -3528 521 -3508
rect 579 -3528 580 -3508
rect 366 -3530 367 -3508
rect 443 -3541 444 -3529
rect 464 -3541 465 -3529
rect 544 -3541 545 -3529
rect 436 -3532 437 -3508
rect 520 -3541 521 -3531
rect 527 -3532 528 -3508
rect 590 -3541 591 -3531
rect 415 -3534 416 -3508
rect 436 -3541 437 -3533
rect 527 -3541 528 -3533
rect 541 -3534 542 -3508
rect 380 -3536 381 -3508
rect 415 -3541 416 -3535
rect 541 -3541 542 -3535
rect 695 -3536 696 -3508
rect 345 -3538 346 -3508
rect 380 -3541 381 -3537
rect 695 -3541 696 -3537
rect 716 -3538 717 -3508
rect 331 -3540 332 -3508
rect 345 -3541 346 -3539
rect 716 -3541 717 -3539
rect 779 -3540 780 -3508
rect 247 -3551 248 -3549
rect 257 -3551 258 -3549
rect 261 -3551 262 -3549
rect 261 -3578 262 -3550
rect 261 -3551 262 -3549
rect 261 -3578 262 -3550
rect 268 -3551 269 -3549
rect 268 -3578 269 -3550
rect 268 -3551 269 -3549
rect 268 -3578 269 -3550
rect 296 -3551 297 -3549
rect 310 -3578 311 -3550
rect 327 -3578 328 -3550
rect 366 -3578 367 -3550
rect 394 -3551 395 -3549
rect 432 -3551 433 -3549
rect 457 -3551 458 -3549
rect 600 -3551 601 -3549
rect 604 -3551 605 -3549
rect 646 -3578 647 -3550
rect 677 -3578 678 -3550
rect 940 -3578 941 -3550
rect 968 -3551 969 -3549
rect 968 -3578 969 -3550
rect 968 -3551 969 -3549
rect 968 -3578 969 -3550
rect 975 -3551 976 -3549
rect 975 -3578 976 -3550
rect 975 -3551 976 -3549
rect 975 -3578 976 -3550
rect 989 -3551 990 -3549
rect 989 -3578 990 -3550
rect 989 -3551 990 -3549
rect 989 -3578 990 -3550
rect 1006 -3551 1007 -3549
rect 1010 -3551 1011 -3549
rect 1038 -3578 1039 -3550
rect 1059 -3551 1060 -3549
rect 1080 -3551 1081 -3549
rect 1087 -3578 1088 -3550
rect 1108 -3551 1109 -3549
rect 1108 -3578 1109 -3550
rect 1108 -3551 1109 -3549
rect 1108 -3578 1109 -3550
rect 1150 -3551 1151 -3549
rect 1157 -3551 1158 -3549
rect 345 -3553 346 -3549
rect 352 -3578 353 -3552
rect 359 -3553 360 -3549
rect 359 -3578 360 -3552
rect 359 -3553 360 -3549
rect 359 -3578 360 -3552
rect 380 -3553 381 -3549
rect 394 -3578 395 -3552
rect 401 -3553 402 -3549
rect 401 -3578 402 -3552
rect 401 -3553 402 -3549
rect 401 -3578 402 -3552
rect 443 -3578 444 -3552
rect 457 -3578 458 -3552
rect 485 -3578 486 -3552
rect 506 -3553 507 -3549
rect 520 -3553 521 -3549
rect 520 -3578 521 -3552
rect 520 -3553 521 -3549
rect 520 -3578 521 -3552
rect 544 -3553 545 -3549
rect 576 -3553 577 -3549
rect 583 -3553 584 -3549
rect 597 -3578 598 -3552
rect 611 -3553 612 -3549
rect 611 -3578 612 -3552
rect 611 -3553 612 -3549
rect 611 -3578 612 -3552
rect 618 -3578 619 -3552
rect 667 -3553 668 -3549
rect 681 -3553 682 -3549
rect 688 -3578 689 -3552
rect 695 -3553 696 -3549
rect 698 -3565 699 -3552
rect 723 -3553 724 -3549
rect 726 -3553 727 -3549
rect 765 -3553 766 -3549
rect 765 -3578 766 -3552
rect 765 -3553 766 -3549
rect 765 -3578 766 -3552
rect 849 -3553 850 -3549
rect 856 -3578 857 -3552
rect 870 -3553 871 -3549
rect 901 -3578 902 -3552
rect 905 -3553 906 -3549
rect 905 -3578 906 -3552
rect 905 -3553 906 -3549
rect 905 -3578 906 -3552
rect 912 -3553 913 -3549
rect 919 -3553 920 -3549
rect 926 -3553 927 -3549
rect 926 -3578 927 -3552
rect 926 -3553 927 -3549
rect 926 -3578 927 -3552
rect 933 -3553 934 -3549
rect 947 -3553 948 -3549
rect 1052 -3553 1053 -3549
rect 1052 -3578 1053 -3552
rect 1052 -3553 1053 -3549
rect 1052 -3578 1053 -3552
rect 488 -3555 489 -3549
rect 534 -3555 535 -3549
rect 562 -3555 563 -3549
rect 628 -3555 629 -3549
rect 639 -3555 640 -3549
rect 660 -3578 661 -3554
rect 695 -3578 696 -3554
rect 702 -3555 703 -3549
rect 723 -3578 724 -3554
rect 730 -3555 731 -3549
rect 835 -3555 836 -3549
rect 849 -3578 850 -3554
rect 863 -3555 864 -3549
rect 919 -3578 920 -3554
rect 450 -3557 451 -3549
rect 562 -3578 563 -3556
rect 702 -3578 703 -3556
rect 716 -3557 717 -3549
rect 730 -3578 731 -3556
rect 737 -3557 738 -3549
rect 884 -3557 885 -3549
rect 922 -3578 923 -3556
rect 450 -3578 451 -3558
rect 453 -3559 454 -3549
rect 464 -3559 465 -3549
rect 488 -3578 489 -3558
rect 492 -3559 493 -3549
rect 534 -3578 535 -3558
rect 716 -3578 717 -3558
rect 737 -3578 738 -3558
rect 751 -3559 752 -3549
rect 891 -3559 892 -3549
rect 912 -3578 913 -3558
rect 436 -3561 437 -3549
rect 464 -3578 465 -3560
rect 478 -3561 479 -3549
rect 492 -3578 493 -3560
rect 499 -3561 500 -3549
rect 506 -3578 507 -3560
rect 751 -3578 752 -3560
rect 758 -3561 759 -3549
rect 877 -3561 878 -3549
rect 891 -3578 892 -3560
rect 898 -3561 899 -3549
rect 982 -3578 983 -3560
rect 415 -3563 416 -3549
rect 436 -3578 437 -3562
rect 471 -3563 472 -3549
rect 499 -3578 500 -3562
rect 744 -3563 745 -3549
rect 758 -3578 759 -3562
rect 408 -3565 409 -3549
rect 415 -3578 416 -3564
rect 422 -3565 423 -3549
rect 471 -3578 472 -3564
rect 478 -3578 479 -3564
rect 541 -3565 542 -3549
rect 726 -3578 727 -3564
rect 744 -3578 745 -3564
rect 376 -3578 377 -3566
rect 408 -3578 409 -3566
rect 541 -3578 542 -3566
rect 555 -3567 556 -3549
rect 555 -3578 556 -3568
rect 569 -3569 570 -3549
rect 548 -3571 549 -3549
rect 569 -3578 570 -3570
rect 527 -3573 528 -3549
rect 548 -3578 549 -3572
rect 513 -3575 514 -3549
rect 527 -3578 528 -3574
rect 513 -3578 514 -3576
rect 590 -3577 591 -3549
rect 264 -3588 265 -3586
rect 268 -3588 269 -3586
rect 310 -3588 311 -3586
rect 327 -3588 328 -3586
rect 352 -3588 353 -3586
rect 352 -3601 353 -3587
rect 352 -3588 353 -3586
rect 352 -3601 353 -3587
rect 359 -3588 360 -3586
rect 376 -3588 377 -3586
rect 394 -3588 395 -3586
rect 401 -3601 402 -3587
rect 408 -3588 409 -3586
rect 446 -3588 447 -3586
rect 450 -3588 451 -3586
rect 457 -3588 458 -3586
rect 492 -3588 493 -3586
rect 516 -3588 517 -3586
rect 520 -3588 521 -3586
rect 544 -3601 545 -3587
rect 562 -3588 563 -3586
rect 677 -3588 678 -3586
rect 695 -3588 696 -3586
rect 695 -3601 696 -3587
rect 695 -3588 696 -3586
rect 695 -3601 696 -3587
rect 702 -3588 703 -3586
rect 702 -3601 703 -3587
rect 702 -3588 703 -3586
rect 702 -3601 703 -3587
rect 716 -3588 717 -3586
rect 716 -3601 717 -3587
rect 716 -3588 717 -3586
rect 716 -3601 717 -3587
rect 751 -3588 752 -3586
rect 754 -3594 755 -3587
rect 758 -3588 759 -3586
rect 772 -3601 773 -3587
rect 849 -3588 850 -3586
rect 863 -3601 864 -3587
rect 905 -3588 906 -3586
rect 908 -3601 909 -3587
rect 912 -3588 913 -3586
rect 919 -3601 920 -3587
rect 926 -3588 927 -3586
rect 926 -3601 927 -3587
rect 926 -3588 927 -3586
rect 926 -3601 927 -3587
rect 940 -3588 941 -3586
rect 1045 -3601 1046 -3587
rect 1052 -3588 1053 -3586
rect 1052 -3601 1053 -3587
rect 1052 -3588 1053 -3586
rect 1052 -3601 1053 -3587
rect 1083 -3588 1084 -3586
rect 1087 -3588 1088 -3586
rect 1108 -3588 1109 -3586
rect 1108 -3601 1109 -3587
rect 1108 -3588 1109 -3586
rect 1108 -3601 1109 -3587
rect 324 -3590 325 -3586
rect 327 -3601 328 -3589
rect 366 -3590 367 -3586
rect 404 -3590 405 -3586
rect 408 -3601 409 -3589
rect 415 -3590 416 -3586
rect 436 -3590 437 -3586
rect 457 -3601 458 -3589
rect 471 -3590 472 -3586
rect 492 -3601 493 -3589
rect 506 -3590 507 -3586
rect 520 -3601 521 -3589
rect 534 -3590 535 -3586
rect 562 -3601 563 -3589
rect 569 -3590 570 -3586
rect 576 -3601 577 -3589
rect 597 -3590 598 -3586
rect 604 -3601 605 -3589
rect 611 -3590 612 -3586
rect 614 -3601 615 -3589
rect 646 -3590 647 -3586
rect 681 -3601 682 -3589
rect 744 -3590 745 -3586
rect 758 -3601 759 -3589
rect 856 -3590 857 -3586
rect 856 -3601 857 -3589
rect 856 -3590 857 -3586
rect 856 -3601 857 -3589
rect 891 -3590 892 -3586
rect 905 -3601 906 -3589
rect 968 -3590 969 -3586
rect 982 -3590 983 -3586
rect 985 -3590 986 -3586
rect 989 -3590 990 -3586
rect 1031 -3601 1032 -3589
rect 1038 -3590 1039 -3586
rect 443 -3592 444 -3586
rect 478 -3592 479 -3586
rect 499 -3592 500 -3586
rect 506 -3601 507 -3591
rect 516 -3601 517 -3591
rect 541 -3592 542 -3586
rect 548 -3592 549 -3586
rect 569 -3601 570 -3591
rect 597 -3601 598 -3591
rect 618 -3592 619 -3586
rect 660 -3592 661 -3586
rect 674 -3592 675 -3586
rect 737 -3592 738 -3586
rect 744 -3601 745 -3591
rect 751 -3601 752 -3591
rect 765 -3592 766 -3586
rect 975 -3592 976 -3586
rect 982 -3601 983 -3591
rect 464 -3594 465 -3586
rect 471 -3601 472 -3593
rect 548 -3601 549 -3593
rect 555 -3594 556 -3586
rect 730 -3594 731 -3586
rect 737 -3601 738 -3593
rect 765 -3601 766 -3593
rect 901 -3594 902 -3586
rect 975 -3601 976 -3593
rect 527 -3596 528 -3586
rect 555 -3601 556 -3595
rect 723 -3596 724 -3586
rect 730 -3601 731 -3595
rect 709 -3598 710 -3586
rect 723 -3601 724 -3597
rect 688 -3600 689 -3586
rect 709 -3601 710 -3599
rect 401 -3611 402 -3609
rect 404 -3617 405 -3610
rect 457 -3611 458 -3609
rect 464 -3626 465 -3610
rect 471 -3611 472 -3609
rect 471 -3626 472 -3610
rect 471 -3611 472 -3609
rect 471 -3626 472 -3610
rect 492 -3611 493 -3609
rect 513 -3611 514 -3609
rect 520 -3611 521 -3609
rect 527 -3626 528 -3610
rect 541 -3611 542 -3609
rect 548 -3611 549 -3609
rect 555 -3611 556 -3609
rect 583 -3626 584 -3610
rect 590 -3626 591 -3610
rect 597 -3611 598 -3609
rect 604 -3611 605 -3609
rect 611 -3611 612 -3609
rect 684 -3611 685 -3609
rect 800 -3626 801 -3610
rect 856 -3611 857 -3609
rect 856 -3626 857 -3610
rect 856 -3611 857 -3609
rect 856 -3626 857 -3610
rect 863 -3611 864 -3609
rect 863 -3626 864 -3610
rect 863 -3611 864 -3609
rect 863 -3626 864 -3610
rect 926 -3611 927 -3609
rect 933 -3626 934 -3610
rect 975 -3611 976 -3609
rect 1003 -3626 1004 -3610
rect 1031 -3611 1032 -3609
rect 1031 -3626 1032 -3610
rect 1031 -3611 1032 -3609
rect 1031 -3626 1032 -3610
rect 1045 -3611 1046 -3609
rect 1080 -3626 1081 -3610
rect 1108 -3611 1109 -3609
rect 1108 -3626 1109 -3610
rect 1108 -3611 1109 -3609
rect 1108 -3626 1109 -3610
rect 401 -3626 402 -3612
rect 506 -3613 507 -3609
rect 516 -3613 517 -3609
rect 562 -3613 563 -3609
rect 562 -3626 563 -3612
rect 562 -3613 563 -3609
rect 562 -3626 563 -3612
rect 569 -3613 570 -3609
rect 569 -3626 570 -3612
rect 569 -3613 570 -3609
rect 569 -3626 570 -3612
rect 576 -3613 577 -3609
rect 576 -3626 577 -3612
rect 576 -3613 577 -3609
rect 576 -3626 577 -3612
rect 709 -3613 710 -3609
rect 712 -3613 713 -3609
rect 730 -3613 731 -3609
rect 775 -3626 776 -3612
rect 919 -3613 920 -3609
rect 926 -3626 927 -3612
rect 982 -3613 983 -3609
rect 982 -3626 983 -3612
rect 982 -3613 983 -3609
rect 982 -3626 983 -3612
rect 1052 -3613 1053 -3609
rect 1059 -3626 1060 -3612
rect 709 -3626 710 -3614
rect 716 -3615 717 -3609
rect 751 -3615 752 -3609
rect 761 -3615 762 -3609
rect 712 -3626 713 -3616
rect 716 -3626 717 -3616
rect 737 -3617 738 -3609
rect 751 -3626 752 -3616
rect 758 -3617 759 -3609
rect 765 -3617 766 -3609
rect 744 -3619 745 -3609
rect 758 -3626 759 -3618
rect 765 -3626 766 -3618
rect 772 -3619 773 -3609
rect 723 -3621 724 -3609
rect 744 -3626 745 -3620
rect 702 -3623 703 -3609
rect 723 -3626 724 -3622
rect 695 -3625 696 -3609
rect 702 -3626 703 -3624
rect 401 -3636 402 -3634
rect 401 -3641 402 -3635
rect 401 -3636 402 -3634
rect 401 -3641 402 -3635
rect 408 -3636 409 -3634
rect 408 -3641 409 -3635
rect 408 -3636 409 -3634
rect 408 -3641 409 -3635
rect 464 -3636 465 -3634
rect 464 -3641 465 -3635
rect 464 -3636 465 -3634
rect 464 -3641 465 -3635
rect 471 -3636 472 -3634
rect 474 -3641 475 -3635
rect 527 -3636 528 -3634
rect 527 -3641 528 -3635
rect 527 -3636 528 -3634
rect 527 -3641 528 -3635
rect 562 -3636 563 -3634
rect 572 -3641 573 -3635
rect 583 -3636 584 -3634
rect 597 -3641 598 -3635
rect 716 -3636 717 -3634
rect 716 -3641 717 -3635
rect 716 -3636 717 -3634
rect 716 -3641 717 -3635
rect 719 -3641 720 -3635
rect 723 -3636 724 -3634
rect 744 -3636 745 -3634
rect 772 -3636 773 -3634
rect 856 -3636 857 -3634
rect 859 -3641 860 -3635
rect 863 -3636 864 -3634
rect 863 -3641 864 -3635
rect 863 -3636 864 -3634
rect 863 -3641 864 -3635
rect 926 -3636 927 -3634
rect 929 -3641 930 -3635
rect 933 -3636 934 -3634
rect 933 -3641 934 -3635
rect 933 -3636 934 -3634
rect 933 -3641 934 -3635
rect 982 -3636 983 -3634
rect 989 -3641 990 -3635
rect 1031 -3636 1032 -3634
rect 1034 -3641 1035 -3635
rect 1055 -3636 1056 -3634
rect 1059 -3636 1060 -3634
rect 1080 -3636 1081 -3634
rect 1094 -3641 1095 -3635
rect 1108 -3636 1109 -3634
rect 1111 -3641 1112 -3635
rect 576 -3638 577 -3634
rect 583 -3641 584 -3637
rect 590 -3638 591 -3634
rect 590 -3641 591 -3637
rect 590 -3638 591 -3634
rect 590 -3641 591 -3637
rect 709 -3638 710 -3634
rect 723 -3641 724 -3637
rect 751 -3638 752 -3634
rect 751 -3641 752 -3637
rect 751 -3638 752 -3634
rect 751 -3641 752 -3637
rect 758 -3638 759 -3634
rect 758 -3641 759 -3637
rect 758 -3638 759 -3634
rect 758 -3641 759 -3637
rect 765 -3638 766 -3634
rect 765 -3641 766 -3637
rect 765 -3638 766 -3634
rect 765 -3641 766 -3637
rect 800 -3638 801 -3634
rect 926 -3641 927 -3637
rect 985 -3641 986 -3637
rect 1052 -3638 1053 -3634
rect 569 -3640 570 -3634
rect 576 -3641 577 -3639
rect 702 -3640 703 -3634
rect 709 -3641 710 -3639
rect 1003 -3640 1004 -3634
rect 1031 -3641 1032 -3639
rect 401 -3651 402 -3649
rect 401 -3656 402 -3650
rect 401 -3651 402 -3649
rect 401 -3656 402 -3650
rect 408 -3651 409 -3649
rect 408 -3656 409 -3650
rect 408 -3651 409 -3649
rect 408 -3656 409 -3650
rect 464 -3651 465 -3649
rect 474 -3651 475 -3649
rect 527 -3651 528 -3649
rect 534 -3656 535 -3650
rect 569 -3651 570 -3649
rect 576 -3651 577 -3649
rect 583 -3651 584 -3649
rect 590 -3651 591 -3649
rect 709 -3651 710 -3649
rect 719 -3651 720 -3649
rect 765 -3651 766 -3649
rect 772 -3656 773 -3650
rect 856 -3651 857 -3649
rect 863 -3651 864 -3649
rect 929 -3651 930 -3649
rect 933 -3651 934 -3649
rect 985 -3651 986 -3649
rect 989 -3651 990 -3649
rect 1094 -3651 1095 -3649
rect 1108 -3651 1109 -3649
rect 586 -3653 587 -3649
rect 597 -3653 598 -3649
rect 716 -3653 717 -3649
rect 723 -3653 724 -3649
rect 758 -3653 759 -3649
rect 765 -3656 766 -3652
rect 751 -3655 752 -3649
rect 758 -3656 759 -3654
rect 404 -3666 405 -3664
rect 408 -3666 409 -3664
rect 527 -3666 528 -3664
rect 534 -3666 535 -3664
rect 758 -3666 759 -3664
rect 765 -3666 766 -3664
rect 768 -3666 769 -3664
rect 772 -3666 773 -3664
<< labels >>
rlabel pdiffusion 3 -12 3 -12 0 cellNo=80
rlabel pdiffusion 10 -12 10 -12 0 cellNo=1108
rlabel pdiffusion 17 -12 17 -12 0 cellNo=1288
rlabel pdiffusion 24 -12 24 -12 0 cellNo=1173
rlabel pdiffusion 31 -12 31 -12 0 cellNo=688
rlabel pdiffusion 38 -12 38 -12 0 cellNo=1133
rlabel pdiffusion 45 -12 45 -12 0 cellNo=1322
rlabel pdiffusion 52 -12 52 -12 0 cellNo=1379
rlabel pdiffusion 59 -12 59 -12 0 cellNo=1409
rlabel pdiffusion 66 -12 66 -12 0 cellNo=1385
rlabel pdiffusion 73 -12 73 -12 0 cellNo=1132
rlabel pdiffusion 80 -12 80 -12 0 cellNo=1159
rlabel pdiffusion 87 -12 87 -12 0 cellNo=1423
rlabel pdiffusion 94 -12 94 -12 0 cellNo=1157
rlabel pdiffusion 101 -12 101 -12 0 cellNo=1059
rlabel pdiffusion 108 -12 108 -12 0 cellNo=1422
rlabel pdiffusion 115 -12 115 -12 0 cellNo=1126
rlabel pdiffusion 122 -12 122 -12 0 cellNo=1075
rlabel pdiffusion 129 -12 129 -12 0 cellNo=1119
rlabel pdiffusion 136 -12 136 -12 0 cellNo=1175
rlabel pdiffusion 143 -12 143 -12 0 cellNo=1242
rlabel pdiffusion 150 -12 150 -12 0 cellNo=1287
rlabel pdiffusion 157 -12 157 -12 0 cellNo=1330
rlabel pdiffusion 164 -12 164 -12 0 cellNo=1372
rlabel pdiffusion 171 -12 171 -12 0 cellNo=1417
rlabel pdiffusion 227 -12 227 -12 0 feedthrough
rlabel pdiffusion 255 -12 255 -12 0 feedthrough
rlabel pdiffusion 276 -12 276 -12 0 feedthrough
rlabel pdiffusion 318 -12 318 -12 0 feedthrough
rlabel pdiffusion 332 -12 332 -12 0 cellNo=178
rlabel pdiffusion 367 -12 367 -12 0 feedthrough
rlabel pdiffusion 374 -12 374 -12 0 cellNo=743
rlabel pdiffusion 381 -12 381 -12 0 cellNo=474
rlabel pdiffusion 395 -12 395 -12 0 cellNo=234
rlabel pdiffusion 402 -12 402 -12 0 cellNo=931
rlabel pdiffusion 416 -12 416 -12 0 feedthrough
rlabel pdiffusion 430 -12 430 -12 0 cellNo=568
rlabel pdiffusion 437 -12 437 -12 0 feedthrough
rlabel pdiffusion 444 -12 444 -12 0 cellNo=732
rlabel pdiffusion 451 -12 451 -12 0 feedthrough
rlabel pdiffusion 458 -12 458 -12 0 cellNo=964
rlabel pdiffusion 472 -12 472 -12 0 feedthrough
rlabel pdiffusion 493 -12 493 -12 0 feedthrough
rlabel pdiffusion 507 -12 507 -12 0 feedthrough
rlabel pdiffusion 514 -12 514 -12 0 cellNo=446
rlabel pdiffusion 528 -12 528 -12 0 feedthrough
rlabel pdiffusion 535 -12 535 -12 0 cellNo=837
rlabel pdiffusion 542 -12 542 -12 0 cellNo=393
rlabel pdiffusion 563 -12 563 -12 0 cellNo=333
rlabel pdiffusion 570 -12 570 -12 0 feedthrough
rlabel pdiffusion 591 -12 591 -12 0 feedthrough
rlabel pdiffusion 619 -12 619 -12 0 cellNo=678
rlabel pdiffusion 640 -12 640 -12 0 cellNo=420
rlabel pdiffusion 668 -12 668 -12 0 cellNo=626
rlabel pdiffusion 675 -12 675 -12 0 feedthrough
rlabel pdiffusion 703 -12 703 -12 0 cellNo=880
rlabel pdiffusion 766 -12 766 -12 0 feedthrough
rlabel pdiffusion 801 -12 801 -12 0 cellNo=941
rlabel pdiffusion 829 -12 829 -12 0 feedthrough
rlabel pdiffusion 843 -12 843 -12 0 feedthrough
rlabel pdiffusion 3 -41 3 -41 0 cellNo=485
rlabel pdiffusion 10 -41 10 -41 0 cellNo=1369
rlabel pdiffusion 17 -41 17 -41 0 cellNo=1280
rlabel pdiffusion 24 -41 24 -41 0 cellNo=1195
rlabel pdiffusion 31 -41 31 -41 0 cellNo=1377
rlabel pdiffusion 38 -41 38 -41 0 cellNo=1153
rlabel pdiffusion 45 -41 45 -41 0 cellNo=1293
rlabel pdiffusion 52 -41 52 -41 0 cellNo=1092
rlabel pdiffusion 59 -41 59 -41 0 cellNo=1077
rlabel pdiffusion 66 -41 66 -41 0 cellNo=1211
rlabel pdiffusion 73 -41 73 -41 0 cellNo=1418
rlabel pdiffusion 80 -41 80 -41 0 cellNo=1207
rlabel pdiffusion 87 -41 87 -41 0 cellNo=1174
rlabel pdiffusion 94 -41 94 -41 0 cellNo=1078
rlabel pdiffusion 101 -41 101 -41 0 cellNo=1117
rlabel pdiffusion 108 -41 108 -41 0 cellNo=1363
rlabel pdiffusion 115 -41 115 -41 0 cellNo=1156
rlabel pdiffusion 122 -41 122 -41 0 cellNo=1008
rlabel pdiffusion 129 -41 129 -41 0 cellNo=1241
rlabel pdiffusion 136 -41 136 -41 0 feedthrough
rlabel pdiffusion 143 -41 143 -41 0 cellNo=1367
rlabel pdiffusion 150 -41 150 -41 0 cellNo=1258
rlabel pdiffusion 178 -41 178 -41 0 cellNo=659
rlabel pdiffusion 192 -41 192 -41 0 feedthrough
rlabel pdiffusion 206 -41 206 -41 0 feedthrough
rlabel pdiffusion 213 -41 213 -41 0 feedthrough
rlabel pdiffusion 220 -41 220 -41 0 cellNo=452
rlabel pdiffusion 227 -41 227 -41 0 feedthrough
rlabel pdiffusion 234 -41 234 -41 0 cellNo=578
rlabel pdiffusion 255 -41 255 -41 0 feedthrough
rlabel pdiffusion 297 -41 297 -41 0 cellNo=805
rlabel pdiffusion 304 -41 304 -41 0 feedthrough
rlabel pdiffusion 311 -41 311 -41 0 cellNo=857
rlabel pdiffusion 318 -41 318 -41 0 feedthrough
rlabel pdiffusion 325 -41 325 -41 0 cellNo=281
rlabel pdiffusion 332 -41 332 -41 0 feedthrough
rlabel pdiffusion 339 -41 339 -41 0 feedthrough
rlabel pdiffusion 346 -41 346 -41 0 feedthrough
rlabel pdiffusion 353 -41 353 -41 0 feedthrough
rlabel pdiffusion 360 -41 360 -41 0 feedthrough
rlabel pdiffusion 367 -41 367 -41 0 cellNo=502
rlabel pdiffusion 374 -41 374 -41 0 feedthrough
rlabel pdiffusion 381 -41 381 -41 0 feedthrough
rlabel pdiffusion 388 -41 388 -41 0 feedthrough
rlabel pdiffusion 395 -41 395 -41 0 cellNo=252
rlabel pdiffusion 402 -41 402 -41 0 cellNo=146
rlabel pdiffusion 409 -41 409 -41 0 feedthrough
rlabel pdiffusion 416 -41 416 -41 0 feedthrough
rlabel pdiffusion 423 -41 423 -41 0 feedthrough
rlabel pdiffusion 444 -41 444 -41 0 cellNo=694
rlabel pdiffusion 451 -41 451 -41 0 cellNo=799
rlabel pdiffusion 458 -41 458 -41 0 feedthrough
rlabel pdiffusion 465 -41 465 -41 0 cellNo=445
rlabel pdiffusion 472 -41 472 -41 0 feedthrough
rlabel pdiffusion 479 -41 479 -41 0 feedthrough
rlabel pdiffusion 486 -41 486 -41 0 cellNo=309
rlabel pdiffusion 493 -41 493 -41 0 feedthrough
rlabel pdiffusion 514 -41 514 -41 0 feedthrough
rlabel pdiffusion 521 -41 521 -41 0 feedthrough
rlabel pdiffusion 528 -41 528 -41 0 feedthrough
rlabel pdiffusion 535 -41 535 -41 0 feedthrough
rlabel pdiffusion 542 -41 542 -41 0 feedthrough
rlabel pdiffusion 549 -41 549 -41 0 feedthrough
rlabel pdiffusion 556 -41 556 -41 0 feedthrough
rlabel pdiffusion 570 -41 570 -41 0 feedthrough
rlabel pdiffusion 577 -41 577 -41 0 feedthrough
rlabel pdiffusion 584 -41 584 -41 0 feedthrough
rlabel pdiffusion 591 -41 591 -41 0 cellNo=205
rlabel pdiffusion 619 -41 619 -41 0 cellNo=728
rlabel pdiffusion 633 -41 633 -41 0 cellNo=819
rlabel pdiffusion 640 -41 640 -41 0 feedthrough
rlabel pdiffusion 647 -41 647 -41 0 feedthrough
rlabel pdiffusion 654 -41 654 -41 0 feedthrough
rlabel pdiffusion 661 -41 661 -41 0 feedthrough
rlabel pdiffusion 668 -41 668 -41 0 feedthrough
rlabel pdiffusion 682 -41 682 -41 0 cellNo=492
rlabel pdiffusion 696 -41 696 -41 0 feedthrough
rlabel pdiffusion 703 -41 703 -41 0 feedthrough
rlabel pdiffusion 710 -41 710 -41 0 feedthrough
rlabel pdiffusion 759 -41 759 -41 0 cellNo=169
rlabel pdiffusion 766 -41 766 -41 0 feedthrough
rlabel pdiffusion 773 -41 773 -41 0 cellNo=501
rlabel pdiffusion 780 -41 780 -41 0 cellNo=965
rlabel pdiffusion 787 -41 787 -41 0 feedthrough
rlabel pdiffusion 794 -41 794 -41 0 feedthrough
rlabel pdiffusion 801 -41 801 -41 0 feedthrough
rlabel pdiffusion 822 -41 822 -41 0 cellNo=753
rlabel pdiffusion 857 -41 857 -41 0 feedthrough
rlabel pdiffusion 878 -41 878 -41 0 feedthrough
rlabel pdiffusion 920 -41 920 -41 0 feedthrough
rlabel pdiffusion 3 -90 3 -90 0 cellNo=1004
rlabel pdiffusion 10 -90 10 -90 0 cellNo=1022
rlabel pdiffusion 17 -90 17 -90 0 cellNo=1116
rlabel pdiffusion 24 -90 24 -90 0 cellNo=1145
rlabel pdiffusion 31 -90 31 -90 0 cellNo=1110
rlabel pdiffusion 38 -90 38 -90 0 cellNo=1130
rlabel pdiffusion 45 -90 45 -90 0 cellNo=1007
rlabel pdiffusion 52 -90 52 -90 0 cellNo=1081
rlabel pdiffusion 59 -90 59 -90 0 cellNo=1300
rlabel pdiffusion 66 -90 66 -90 0 cellNo=1149
rlabel pdiffusion 73 -90 73 -90 0 cellNo=1169
rlabel pdiffusion 80 -90 80 -90 0 feedthrough
rlabel pdiffusion 87 -90 87 -90 0 cellNo=1206
rlabel pdiffusion 94 -90 94 -90 0 cellNo=1237
rlabel pdiffusion 101 -90 101 -90 0 feedthrough
rlabel pdiffusion 108 -90 108 -90 0 cellNo=1378
rlabel pdiffusion 115 -90 115 -90 0 cellNo=215
rlabel pdiffusion 122 -90 122 -90 0 cellNo=1155
rlabel pdiffusion 129 -90 129 -90 0 feedthrough
rlabel pdiffusion 136 -90 136 -90 0 cellNo=1341
rlabel pdiffusion 143 -90 143 -90 0 cellNo=770
rlabel pdiffusion 150 -90 150 -90 0 feedthrough
rlabel pdiffusion 157 -90 157 -90 0 feedthrough
rlabel pdiffusion 164 -90 164 -90 0 feedthrough
rlabel pdiffusion 171 -90 171 -90 0 feedthrough
rlabel pdiffusion 178 -90 178 -90 0 cellNo=566
rlabel pdiffusion 185 -90 185 -90 0 feedthrough
rlabel pdiffusion 192 -90 192 -90 0 feedthrough
rlabel pdiffusion 199 -90 199 -90 0 feedthrough
rlabel pdiffusion 206 -90 206 -90 0 feedthrough
rlabel pdiffusion 213 -90 213 -90 0 cellNo=930
rlabel pdiffusion 220 -90 220 -90 0 feedthrough
rlabel pdiffusion 227 -90 227 -90 0 cellNo=802
rlabel pdiffusion 234 -90 234 -90 0 cellNo=698
rlabel pdiffusion 241 -90 241 -90 0 cellNo=36
rlabel pdiffusion 248 -90 248 -90 0 cellNo=1089
rlabel pdiffusion 255 -90 255 -90 0 feedthrough
rlabel pdiffusion 262 -90 262 -90 0 feedthrough
rlabel pdiffusion 269 -90 269 -90 0 feedthrough
rlabel pdiffusion 276 -90 276 -90 0 cellNo=479
rlabel pdiffusion 283 -90 283 -90 0 cellNo=894
rlabel pdiffusion 290 -90 290 -90 0 feedthrough
rlabel pdiffusion 297 -90 297 -90 0 cellNo=396
rlabel pdiffusion 304 -90 304 -90 0 feedthrough
rlabel pdiffusion 311 -90 311 -90 0 feedthrough
rlabel pdiffusion 318 -90 318 -90 0 feedthrough
rlabel pdiffusion 325 -90 325 -90 0 feedthrough
rlabel pdiffusion 332 -90 332 -90 0 cellNo=116
rlabel pdiffusion 339 -90 339 -90 0 feedthrough
rlabel pdiffusion 346 -90 346 -90 0 feedthrough
rlabel pdiffusion 353 -90 353 -90 0 feedthrough
rlabel pdiffusion 360 -90 360 -90 0 feedthrough
rlabel pdiffusion 367 -90 367 -90 0 cellNo=308
rlabel pdiffusion 374 -90 374 -90 0 feedthrough
rlabel pdiffusion 381 -90 381 -90 0 feedthrough
rlabel pdiffusion 388 -90 388 -90 0 cellNo=1158
rlabel pdiffusion 395 -90 395 -90 0 cellNo=1080
rlabel pdiffusion 402 -90 402 -90 0 feedthrough
rlabel pdiffusion 409 -90 409 -90 0 feedthrough
rlabel pdiffusion 416 -90 416 -90 0 feedthrough
rlabel pdiffusion 423 -90 423 -90 0 feedthrough
rlabel pdiffusion 430 -90 430 -90 0 feedthrough
rlabel pdiffusion 437 -90 437 -90 0 feedthrough
rlabel pdiffusion 444 -90 444 -90 0 cellNo=159
rlabel pdiffusion 451 -90 451 -90 0 cellNo=179
rlabel pdiffusion 458 -90 458 -90 0 feedthrough
rlabel pdiffusion 465 -90 465 -90 0 feedthrough
rlabel pdiffusion 472 -90 472 -90 0 cellNo=470
rlabel pdiffusion 479 -90 479 -90 0 feedthrough
rlabel pdiffusion 486 -90 486 -90 0 feedthrough
rlabel pdiffusion 493 -90 493 -90 0 feedthrough
rlabel pdiffusion 500 -90 500 -90 0 feedthrough
rlabel pdiffusion 507 -90 507 -90 0 feedthrough
rlabel pdiffusion 514 -90 514 -90 0 feedthrough
rlabel pdiffusion 521 -90 521 -90 0 feedthrough
rlabel pdiffusion 528 -90 528 -90 0 feedthrough
rlabel pdiffusion 535 -90 535 -90 0 feedthrough
rlabel pdiffusion 542 -90 542 -90 0 feedthrough
rlabel pdiffusion 549 -90 549 -90 0 feedthrough
rlabel pdiffusion 556 -90 556 -90 0 feedthrough
rlabel pdiffusion 563 -90 563 -90 0 feedthrough
rlabel pdiffusion 570 -90 570 -90 0 cellNo=636
rlabel pdiffusion 577 -90 577 -90 0 feedthrough
rlabel pdiffusion 584 -90 584 -90 0 feedthrough
rlabel pdiffusion 591 -90 591 -90 0 cellNo=807
rlabel pdiffusion 598 -90 598 -90 0 feedthrough
rlabel pdiffusion 605 -90 605 -90 0 feedthrough
rlabel pdiffusion 612 -90 612 -90 0 feedthrough
rlabel pdiffusion 619 -90 619 -90 0 feedthrough
rlabel pdiffusion 626 -90 626 -90 0 cellNo=200
rlabel pdiffusion 633 -90 633 -90 0 feedthrough
rlabel pdiffusion 640 -90 640 -90 0 cellNo=195
rlabel pdiffusion 647 -90 647 -90 0 feedthrough
rlabel pdiffusion 654 -90 654 -90 0 feedthrough
rlabel pdiffusion 661 -90 661 -90 0 feedthrough
rlabel pdiffusion 668 -90 668 -90 0 feedthrough
rlabel pdiffusion 675 -90 675 -90 0 feedthrough
rlabel pdiffusion 682 -90 682 -90 0 feedthrough
rlabel pdiffusion 689 -90 689 -90 0 feedthrough
rlabel pdiffusion 696 -90 696 -90 0 feedthrough
rlabel pdiffusion 703 -90 703 -90 0 feedthrough
rlabel pdiffusion 710 -90 710 -90 0 feedthrough
rlabel pdiffusion 717 -90 717 -90 0 feedthrough
rlabel pdiffusion 724 -90 724 -90 0 feedthrough
rlabel pdiffusion 731 -90 731 -90 0 cellNo=733
rlabel pdiffusion 738 -90 738 -90 0 cellNo=84
rlabel pdiffusion 745 -90 745 -90 0 feedthrough
rlabel pdiffusion 752 -90 752 -90 0 feedthrough
rlabel pdiffusion 759 -90 759 -90 0 cellNo=808
rlabel pdiffusion 766 -90 766 -90 0 feedthrough
rlabel pdiffusion 773 -90 773 -90 0 feedthrough
rlabel pdiffusion 780 -90 780 -90 0 cellNo=497
rlabel pdiffusion 787 -90 787 -90 0 feedthrough
rlabel pdiffusion 794 -90 794 -90 0 feedthrough
rlabel pdiffusion 801 -90 801 -90 0 feedthrough
rlabel pdiffusion 808 -90 808 -90 0 feedthrough
rlabel pdiffusion 815 -90 815 -90 0 feedthrough
rlabel pdiffusion 822 -90 822 -90 0 feedthrough
rlabel pdiffusion 857 -90 857 -90 0 feedthrough
rlabel pdiffusion 864 -90 864 -90 0 feedthrough
rlabel pdiffusion 871 -90 871 -90 0 feedthrough
rlabel pdiffusion 892 -90 892 -90 0 feedthrough
rlabel pdiffusion 906 -90 906 -90 0 feedthrough
rlabel pdiffusion 969 -90 969 -90 0 feedthrough
rlabel pdiffusion 3 -161 3 -161 0 cellNo=143
rlabel pdiffusion 10 -161 10 -161 0 cellNo=1067
rlabel pdiffusion 17 -161 17 -161 0 cellNo=1002
rlabel pdiffusion 24 -161 24 -161 0 cellNo=1371
rlabel pdiffusion 31 -161 31 -161 0 cellNo=1386
rlabel pdiffusion 38 -161 38 -161 0 cellNo=1006
rlabel pdiffusion 45 -161 45 -161 0 cellNo=1030
rlabel pdiffusion 52 -161 52 -161 0 cellNo=1087
rlabel pdiffusion 59 -161 59 -161 0 cellNo=1205
rlabel pdiffusion 66 -161 66 -161 0 cellNo=1115
rlabel pdiffusion 73 -161 73 -161 0 cellNo=1171
rlabel pdiffusion 80 -161 80 -161 0 cellNo=1125
rlabel pdiffusion 87 -161 87 -161 0 cellNo=1172
rlabel pdiffusion 94 -161 94 -161 0 cellNo=1236
rlabel pdiffusion 101 -161 101 -161 0 cellNo=651
rlabel pdiffusion 108 -161 108 -161 0 cellNo=1252
rlabel pdiffusion 115 -161 115 -161 0 feedthrough
rlabel pdiffusion 122 -161 122 -161 0 cellNo=1416
rlabel pdiffusion 129 -161 129 -161 0 cellNo=1427
rlabel pdiffusion 150 -161 150 -161 0 feedthrough
rlabel pdiffusion 157 -161 157 -161 0 cellNo=926
rlabel pdiffusion 164 -161 164 -161 0 feedthrough
rlabel pdiffusion 171 -161 171 -161 0 feedthrough
rlabel pdiffusion 178 -161 178 -161 0 feedthrough
rlabel pdiffusion 185 -161 185 -161 0 feedthrough
rlabel pdiffusion 192 -161 192 -161 0 feedthrough
rlabel pdiffusion 199 -161 199 -161 0 feedthrough
rlabel pdiffusion 206 -161 206 -161 0 feedthrough
rlabel pdiffusion 213 -161 213 -161 0 feedthrough
rlabel pdiffusion 220 -161 220 -161 0 feedthrough
rlabel pdiffusion 227 -161 227 -161 0 feedthrough
rlabel pdiffusion 234 -161 234 -161 0 feedthrough
rlabel pdiffusion 241 -161 241 -161 0 feedthrough
rlabel pdiffusion 248 -161 248 -161 0 cellNo=640
rlabel pdiffusion 255 -161 255 -161 0 cellNo=284
rlabel pdiffusion 262 -161 262 -161 0 feedthrough
rlabel pdiffusion 269 -161 269 -161 0 cellNo=834
rlabel pdiffusion 276 -161 276 -161 0 cellNo=843
rlabel pdiffusion 283 -161 283 -161 0 cellNo=540
rlabel pdiffusion 290 -161 290 -161 0 cellNo=156
rlabel pdiffusion 297 -161 297 -161 0 cellNo=307
rlabel pdiffusion 304 -161 304 -161 0 feedthrough
rlabel pdiffusion 311 -161 311 -161 0 feedthrough
rlabel pdiffusion 318 -161 318 -161 0 feedthrough
rlabel pdiffusion 325 -161 325 -161 0 feedthrough
rlabel pdiffusion 332 -161 332 -161 0 feedthrough
rlabel pdiffusion 339 -161 339 -161 0 feedthrough
rlabel pdiffusion 346 -161 346 -161 0 feedthrough
rlabel pdiffusion 353 -161 353 -161 0 feedthrough
rlabel pdiffusion 360 -161 360 -161 0 feedthrough
rlabel pdiffusion 367 -161 367 -161 0 feedthrough
rlabel pdiffusion 374 -161 374 -161 0 feedthrough
rlabel pdiffusion 381 -161 381 -161 0 feedthrough
rlabel pdiffusion 388 -161 388 -161 0 cellNo=238
rlabel pdiffusion 395 -161 395 -161 0 feedthrough
rlabel pdiffusion 402 -161 402 -161 0 feedthrough
rlabel pdiffusion 409 -161 409 -161 0 feedthrough
rlabel pdiffusion 416 -161 416 -161 0 cellNo=131
rlabel pdiffusion 423 -161 423 -161 0 feedthrough
rlabel pdiffusion 430 -161 430 -161 0 cellNo=47
rlabel pdiffusion 437 -161 437 -161 0 feedthrough
rlabel pdiffusion 444 -161 444 -161 0 feedthrough
rlabel pdiffusion 451 -161 451 -161 0 feedthrough
rlabel pdiffusion 458 -161 458 -161 0 feedthrough
rlabel pdiffusion 465 -161 465 -161 0 cellNo=55
rlabel pdiffusion 472 -161 472 -161 0 cellNo=533
rlabel pdiffusion 479 -161 479 -161 0 feedthrough
rlabel pdiffusion 486 -161 486 -161 0 cellNo=59
rlabel pdiffusion 493 -161 493 -161 0 feedthrough
rlabel pdiffusion 500 -161 500 -161 0 feedthrough
rlabel pdiffusion 507 -161 507 -161 0 cellNo=296
rlabel pdiffusion 514 -161 514 -161 0 feedthrough
rlabel pdiffusion 521 -161 521 -161 0 feedthrough
rlabel pdiffusion 528 -161 528 -161 0 feedthrough
rlabel pdiffusion 535 -161 535 -161 0 feedthrough
rlabel pdiffusion 542 -161 542 -161 0 feedthrough
rlabel pdiffusion 549 -161 549 -161 0 feedthrough
rlabel pdiffusion 556 -161 556 -161 0 cellNo=993
rlabel pdiffusion 563 -161 563 -161 0 feedthrough
rlabel pdiffusion 570 -161 570 -161 0 feedthrough
rlabel pdiffusion 577 -161 577 -161 0 feedthrough
rlabel pdiffusion 584 -161 584 -161 0 feedthrough
rlabel pdiffusion 591 -161 591 -161 0 feedthrough
rlabel pdiffusion 598 -161 598 -161 0 feedthrough
rlabel pdiffusion 605 -161 605 -161 0 feedthrough
rlabel pdiffusion 612 -161 612 -161 0 feedthrough
rlabel pdiffusion 619 -161 619 -161 0 cellNo=517
rlabel pdiffusion 626 -161 626 -161 0 feedthrough
rlabel pdiffusion 633 -161 633 -161 0 feedthrough
rlabel pdiffusion 640 -161 640 -161 0 feedthrough
rlabel pdiffusion 647 -161 647 -161 0 feedthrough
rlabel pdiffusion 654 -161 654 -161 0 feedthrough
rlabel pdiffusion 661 -161 661 -161 0 feedthrough
rlabel pdiffusion 668 -161 668 -161 0 feedthrough
rlabel pdiffusion 675 -161 675 -161 0 feedthrough
rlabel pdiffusion 682 -161 682 -161 0 cellNo=936
rlabel pdiffusion 689 -161 689 -161 0 feedthrough
rlabel pdiffusion 696 -161 696 -161 0 cellNo=902
rlabel pdiffusion 703 -161 703 -161 0 cellNo=602
rlabel pdiffusion 710 -161 710 -161 0 feedthrough
rlabel pdiffusion 717 -161 717 -161 0 feedthrough
rlabel pdiffusion 724 -161 724 -161 0 feedthrough
rlabel pdiffusion 731 -161 731 -161 0 feedthrough
rlabel pdiffusion 738 -161 738 -161 0 feedthrough
rlabel pdiffusion 745 -161 745 -161 0 feedthrough
rlabel pdiffusion 752 -161 752 -161 0 cellNo=45
rlabel pdiffusion 759 -161 759 -161 0 feedthrough
rlabel pdiffusion 766 -161 766 -161 0 feedthrough
rlabel pdiffusion 773 -161 773 -161 0 feedthrough
rlabel pdiffusion 780 -161 780 -161 0 feedthrough
rlabel pdiffusion 787 -161 787 -161 0 feedthrough
rlabel pdiffusion 794 -161 794 -161 0 feedthrough
rlabel pdiffusion 801 -161 801 -161 0 feedthrough
rlabel pdiffusion 808 -161 808 -161 0 feedthrough
rlabel pdiffusion 815 -161 815 -161 0 feedthrough
rlabel pdiffusion 822 -161 822 -161 0 feedthrough
rlabel pdiffusion 829 -161 829 -161 0 feedthrough
rlabel pdiffusion 836 -161 836 -161 0 feedthrough
rlabel pdiffusion 843 -161 843 -161 0 feedthrough
rlabel pdiffusion 850 -161 850 -161 0 feedthrough
rlabel pdiffusion 857 -161 857 -161 0 feedthrough
rlabel pdiffusion 864 -161 864 -161 0 feedthrough
rlabel pdiffusion 871 -161 871 -161 0 feedthrough
rlabel pdiffusion 878 -161 878 -161 0 feedthrough
rlabel pdiffusion 885 -161 885 -161 0 feedthrough
rlabel pdiffusion 892 -161 892 -161 0 feedthrough
rlabel pdiffusion 899 -161 899 -161 0 feedthrough
rlabel pdiffusion 906 -161 906 -161 0 feedthrough
rlabel pdiffusion 913 -161 913 -161 0 feedthrough
rlabel pdiffusion 920 -161 920 -161 0 feedthrough
rlabel pdiffusion 927 -161 927 -161 0 feedthrough
rlabel pdiffusion 934 -161 934 -161 0 feedthrough
rlabel pdiffusion 941 -161 941 -161 0 cellNo=51
rlabel pdiffusion 948 -161 948 -161 0 cellNo=184
rlabel pdiffusion 955 -161 955 -161 0 feedthrough
rlabel pdiffusion 962 -161 962 -161 0 feedthrough
rlabel pdiffusion 969 -161 969 -161 0 feedthrough
rlabel pdiffusion 976 -161 976 -161 0 feedthrough
rlabel pdiffusion 983 -161 983 -161 0 feedthrough
rlabel pdiffusion 990 -161 990 -161 0 feedthrough
rlabel pdiffusion 997 -161 997 -161 0 cellNo=746
rlabel pdiffusion 1004 -161 1004 -161 0 feedthrough
rlabel pdiffusion 3 -256 3 -256 0 cellNo=1023
rlabel pdiffusion 10 -256 10 -256 0 cellNo=1192
rlabel pdiffusion 17 -256 17 -256 0 cellNo=1200
rlabel pdiffusion 24 -256 24 -256 0 cellNo=1247
rlabel pdiffusion 31 -256 31 -256 0 cellNo=1451
rlabel pdiffusion 38 -256 38 -256 0 cellNo=1334
rlabel pdiffusion 45 -256 45 -256 0 cellNo=1339
rlabel pdiffusion 52 -256 52 -256 0 cellNo=237
rlabel pdiffusion 59 -256 59 -256 0 cellNo=1189
rlabel pdiffusion 66 -256 66 -256 0 cellNo=1276
rlabel pdiffusion 73 -256 73 -256 0 feedthrough
rlabel pdiffusion 80 -256 80 -256 0 cellNo=1294
rlabel pdiffusion 87 -256 87 -256 0 cellNo=1218
rlabel pdiffusion 94 -256 94 -256 0 cellNo=1154
rlabel pdiffusion 101 -256 101 -256 0 feedthrough
rlabel pdiffusion 108 -256 108 -256 0 cellNo=881
rlabel pdiffusion 115 -256 115 -256 0 feedthrough
rlabel pdiffusion 122 -256 122 -256 0 cellNo=565
rlabel pdiffusion 129 -256 129 -256 0 feedthrough
rlabel pdiffusion 136 -256 136 -256 0 feedthrough
rlabel pdiffusion 143 -256 143 -256 0 cellNo=1170
rlabel pdiffusion 150 -256 150 -256 0 cellNo=1204
rlabel pdiffusion 157 -256 157 -256 0 cellNo=1124
rlabel pdiffusion 164 -256 164 -256 0 cellNo=582
rlabel pdiffusion 171 -256 171 -256 0 cellNo=858
rlabel pdiffusion 178 -256 178 -256 0 feedthrough
rlabel pdiffusion 185 -256 185 -256 0 feedthrough
rlabel pdiffusion 192 -256 192 -256 0 feedthrough
rlabel pdiffusion 199 -256 199 -256 0 feedthrough
rlabel pdiffusion 206 -256 206 -256 0 cellNo=448
rlabel pdiffusion 213 -256 213 -256 0 feedthrough
rlabel pdiffusion 220 -256 220 -256 0 cellNo=860
rlabel pdiffusion 227 -256 227 -256 0 feedthrough
rlabel pdiffusion 234 -256 234 -256 0 feedthrough
rlabel pdiffusion 241 -256 241 -256 0 cellNo=1251
rlabel pdiffusion 248 -256 248 -256 0 feedthrough
rlabel pdiffusion 255 -256 255 -256 0 feedthrough
rlabel pdiffusion 262 -256 262 -256 0 feedthrough
rlabel pdiffusion 269 -256 269 -256 0 feedthrough
rlabel pdiffusion 276 -256 276 -256 0 feedthrough
rlabel pdiffusion 283 -256 283 -256 0 cellNo=608
rlabel pdiffusion 290 -256 290 -256 0 feedthrough
rlabel pdiffusion 297 -256 297 -256 0 feedthrough
rlabel pdiffusion 304 -256 304 -256 0 feedthrough
rlabel pdiffusion 311 -256 311 -256 0 feedthrough
rlabel pdiffusion 318 -256 318 -256 0 cellNo=311
rlabel pdiffusion 325 -256 325 -256 0 feedthrough
rlabel pdiffusion 332 -256 332 -256 0 feedthrough
rlabel pdiffusion 339 -256 339 -256 0 cellNo=140
rlabel pdiffusion 346 -256 346 -256 0 feedthrough
rlabel pdiffusion 353 -256 353 -256 0 feedthrough
rlabel pdiffusion 360 -256 360 -256 0 feedthrough
rlabel pdiffusion 367 -256 367 -256 0 feedthrough
rlabel pdiffusion 374 -256 374 -256 0 feedthrough
rlabel pdiffusion 381 -256 381 -256 0 feedthrough
rlabel pdiffusion 388 -256 388 -256 0 feedthrough
rlabel pdiffusion 395 -256 395 -256 0 feedthrough
rlabel pdiffusion 402 -256 402 -256 0 cellNo=527
rlabel pdiffusion 409 -256 409 -256 0 feedthrough
rlabel pdiffusion 416 -256 416 -256 0 feedthrough
rlabel pdiffusion 423 -256 423 -256 0 feedthrough
rlabel pdiffusion 430 -256 430 -256 0 cellNo=835
rlabel pdiffusion 437 -256 437 -256 0 feedthrough
rlabel pdiffusion 444 -256 444 -256 0 cellNo=724
rlabel pdiffusion 451 -256 451 -256 0 cellNo=121
rlabel pdiffusion 458 -256 458 -256 0 feedthrough
rlabel pdiffusion 465 -256 465 -256 0 feedthrough
rlabel pdiffusion 472 -256 472 -256 0 feedthrough
rlabel pdiffusion 479 -256 479 -256 0 cellNo=844
rlabel pdiffusion 486 -256 486 -256 0 cellNo=158
rlabel pdiffusion 493 -256 493 -256 0 cellNo=83
rlabel pdiffusion 500 -256 500 -256 0 feedthrough
rlabel pdiffusion 507 -256 507 -256 0 feedthrough
rlabel pdiffusion 514 -256 514 -256 0 cellNo=551
rlabel pdiffusion 521 -256 521 -256 0 feedthrough
rlabel pdiffusion 528 -256 528 -256 0 feedthrough
rlabel pdiffusion 535 -256 535 -256 0 cellNo=160
rlabel pdiffusion 542 -256 542 -256 0 cellNo=251
rlabel pdiffusion 549 -256 549 -256 0 feedthrough
rlabel pdiffusion 556 -256 556 -256 0 feedthrough
rlabel pdiffusion 563 -256 563 -256 0 feedthrough
rlabel pdiffusion 570 -256 570 -256 0 feedthrough
rlabel pdiffusion 577 -256 577 -256 0 feedthrough
rlabel pdiffusion 584 -256 584 -256 0 cellNo=889
rlabel pdiffusion 591 -256 591 -256 0 feedthrough
rlabel pdiffusion 598 -256 598 -256 0 feedthrough
rlabel pdiffusion 605 -256 605 -256 0 feedthrough
rlabel pdiffusion 612 -256 612 -256 0 cellNo=359
rlabel pdiffusion 619 -256 619 -256 0 feedthrough
rlabel pdiffusion 626 -256 626 -256 0 feedthrough
rlabel pdiffusion 633 -256 633 -256 0 feedthrough
rlabel pdiffusion 640 -256 640 -256 0 feedthrough
rlabel pdiffusion 647 -256 647 -256 0 feedthrough
rlabel pdiffusion 654 -256 654 -256 0 feedthrough
rlabel pdiffusion 661 -256 661 -256 0 feedthrough
rlabel pdiffusion 668 -256 668 -256 0 feedthrough
rlabel pdiffusion 675 -256 675 -256 0 feedthrough
rlabel pdiffusion 682 -256 682 -256 0 cellNo=167
rlabel pdiffusion 689 -256 689 -256 0 feedthrough
rlabel pdiffusion 696 -256 696 -256 0 feedthrough
rlabel pdiffusion 703 -256 703 -256 0 feedthrough
rlabel pdiffusion 710 -256 710 -256 0 feedthrough
rlabel pdiffusion 717 -256 717 -256 0 feedthrough
rlabel pdiffusion 724 -256 724 -256 0 feedthrough
rlabel pdiffusion 731 -256 731 -256 0 feedthrough
rlabel pdiffusion 738 -256 738 -256 0 feedthrough
rlabel pdiffusion 745 -256 745 -256 0 feedthrough
rlabel pdiffusion 752 -256 752 -256 0 feedthrough
rlabel pdiffusion 759 -256 759 -256 0 feedthrough
rlabel pdiffusion 766 -256 766 -256 0 cellNo=561
rlabel pdiffusion 773 -256 773 -256 0 feedthrough
rlabel pdiffusion 780 -256 780 -256 0 feedthrough
rlabel pdiffusion 787 -256 787 -256 0 feedthrough
rlabel pdiffusion 794 -256 794 -256 0 feedthrough
rlabel pdiffusion 801 -256 801 -256 0 feedthrough
rlabel pdiffusion 808 -256 808 -256 0 feedthrough
rlabel pdiffusion 815 -256 815 -256 0 feedthrough
rlabel pdiffusion 822 -256 822 -256 0 feedthrough
rlabel pdiffusion 829 -256 829 -256 0 cellNo=278
rlabel pdiffusion 836 -256 836 -256 0 feedthrough
rlabel pdiffusion 843 -256 843 -256 0 cellNo=469
rlabel pdiffusion 850 -256 850 -256 0 feedthrough
rlabel pdiffusion 857 -256 857 -256 0 feedthrough
rlabel pdiffusion 864 -256 864 -256 0 feedthrough
rlabel pdiffusion 871 -256 871 -256 0 feedthrough
rlabel pdiffusion 878 -256 878 -256 0 feedthrough
rlabel pdiffusion 885 -256 885 -256 0 feedthrough
rlabel pdiffusion 892 -256 892 -256 0 feedthrough
rlabel pdiffusion 899 -256 899 -256 0 feedthrough
rlabel pdiffusion 906 -256 906 -256 0 feedthrough
rlabel pdiffusion 913 -256 913 -256 0 feedthrough
rlabel pdiffusion 920 -256 920 -256 0 feedthrough
rlabel pdiffusion 927 -256 927 -256 0 feedthrough
rlabel pdiffusion 934 -256 934 -256 0 feedthrough
rlabel pdiffusion 941 -256 941 -256 0 feedthrough
rlabel pdiffusion 948 -256 948 -256 0 feedthrough
rlabel pdiffusion 955 -256 955 -256 0 feedthrough
rlabel pdiffusion 962 -256 962 -256 0 feedthrough
rlabel pdiffusion 969 -256 969 -256 0 feedthrough
rlabel pdiffusion 976 -256 976 -256 0 feedthrough
rlabel pdiffusion 983 -256 983 -256 0 feedthrough
rlabel pdiffusion 990 -256 990 -256 0 feedthrough
rlabel pdiffusion 997 -256 997 -256 0 feedthrough
rlabel pdiffusion 1004 -256 1004 -256 0 feedthrough
rlabel pdiffusion 1011 -256 1011 -256 0 feedthrough
rlabel pdiffusion 1018 -256 1018 -256 0 feedthrough
rlabel pdiffusion 1025 -256 1025 -256 0 feedthrough
rlabel pdiffusion 1032 -256 1032 -256 0 feedthrough
rlabel pdiffusion 1039 -256 1039 -256 0 feedthrough
rlabel pdiffusion 1046 -256 1046 -256 0 feedthrough
rlabel pdiffusion 1053 -256 1053 -256 0 feedthrough
rlabel pdiffusion 1060 -256 1060 -256 0 feedthrough
rlabel pdiffusion 1067 -256 1067 -256 0 feedthrough
rlabel pdiffusion 1074 -256 1074 -256 0 feedthrough
rlabel pdiffusion 1081 -256 1081 -256 0 feedthrough
rlabel pdiffusion 1088 -256 1088 -256 0 feedthrough
rlabel pdiffusion 1095 -256 1095 -256 0 feedthrough
rlabel pdiffusion 1102 -256 1102 -256 0 feedthrough
rlabel pdiffusion 1109 -256 1109 -256 0 feedthrough
rlabel pdiffusion 1116 -256 1116 -256 0 feedthrough
rlabel pdiffusion 1123 -256 1123 -256 0 feedthrough
rlabel pdiffusion 1130 -256 1130 -256 0 feedthrough
rlabel pdiffusion 3 -359 3 -359 0 cellNo=1001
rlabel pdiffusion 10 -359 10 -359 0 cellNo=1003
rlabel pdiffusion 17 -359 17 -359 0 cellNo=1279
rlabel pdiffusion 24 -359 24 -359 0 cellNo=1005
rlabel pdiffusion 31 -359 31 -359 0 cellNo=1337
rlabel pdiffusion 38 -359 38 -359 0 cellNo=1013
rlabel pdiffusion 45 -359 45 -359 0 cellNo=1234
rlabel pdiffusion 52 -359 52 -359 0 feedthrough
rlabel pdiffusion 59 -359 59 -359 0 cellNo=57
rlabel pdiffusion 66 -359 66 -359 0 cellNo=1188
rlabel pdiffusion 73 -359 73 -359 0 cellNo=371
rlabel pdiffusion 80 -359 80 -359 0 cellNo=785
rlabel pdiffusion 87 -359 87 -359 0 feedthrough
rlabel pdiffusion 94 -359 94 -359 0 feedthrough
rlabel pdiffusion 101 -359 101 -359 0 feedthrough
rlabel pdiffusion 108 -359 108 -359 0 feedthrough
rlabel pdiffusion 115 -359 115 -359 0 feedthrough
rlabel pdiffusion 122 -359 122 -359 0 cellNo=250
rlabel pdiffusion 129 -359 129 -359 0 feedthrough
rlabel pdiffusion 136 -359 136 -359 0 feedthrough
rlabel pdiffusion 143 -359 143 -359 0 feedthrough
rlabel pdiffusion 150 -359 150 -359 0 feedthrough
rlabel pdiffusion 157 -359 157 -359 0 cellNo=697
rlabel pdiffusion 164 -359 164 -359 0 feedthrough
rlabel pdiffusion 171 -359 171 -359 0 cellNo=35
rlabel pdiffusion 178 -359 178 -359 0 feedthrough
rlabel pdiffusion 185 -359 185 -359 0 feedthrough
rlabel pdiffusion 192 -359 192 -359 0 feedthrough
rlabel pdiffusion 199 -359 199 -359 0 feedthrough
rlabel pdiffusion 206 -359 206 -359 0 feedthrough
rlabel pdiffusion 213 -359 213 -359 0 feedthrough
rlabel pdiffusion 220 -359 220 -359 0 feedthrough
rlabel pdiffusion 227 -359 227 -359 0 feedthrough
rlabel pdiffusion 234 -359 234 -359 0 cellNo=10
rlabel pdiffusion 241 -359 241 -359 0 feedthrough
rlabel pdiffusion 248 -359 248 -359 0 cellNo=1382
rlabel pdiffusion 255 -359 255 -359 0 feedthrough
rlabel pdiffusion 262 -359 262 -359 0 cellNo=1203
rlabel pdiffusion 269 -359 269 -359 0 feedthrough
rlabel pdiffusion 276 -359 276 -359 0 feedthrough
rlabel pdiffusion 283 -359 283 -359 0 cellNo=1428
rlabel pdiffusion 290 -359 290 -359 0 feedthrough
rlabel pdiffusion 297 -359 297 -359 0 feedthrough
rlabel pdiffusion 304 -359 304 -359 0 feedthrough
rlabel pdiffusion 311 -359 311 -359 0 feedthrough
rlabel pdiffusion 318 -359 318 -359 0 feedthrough
rlabel pdiffusion 325 -359 325 -359 0 feedthrough
rlabel pdiffusion 332 -359 332 -359 0 cellNo=1327
rlabel pdiffusion 339 -359 339 -359 0 feedthrough
rlabel pdiffusion 346 -359 346 -359 0 feedthrough
rlabel pdiffusion 353 -359 353 -359 0 feedthrough
rlabel pdiffusion 360 -359 360 -359 0 cellNo=1243
rlabel pdiffusion 367 -359 367 -359 0 cellNo=1260
rlabel pdiffusion 374 -359 374 -359 0 feedthrough
rlabel pdiffusion 381 -359 381 -359 0 feedthrough
rlabel pdiffusion 388 -359 388 -359 0 feedthrough
rlabel pdiffusion 395 -359 395 -359 0 feedthrough
rlabel pdiffusion 402 -359 402 -359 0 feedthrough
rlabel pdiffusion 409 -359 409 -359 0 feedthrough
rlabel pdiffusion 416 -359 416 -359 0 feedthrough
rlabel pdiffusion 423 -359 423 -359 0 feedthrough
rlabel pdiffusion 430 -359 430 -359 0 feedthrough
rlabel pdiffusion 437 -359 437 -359 0 feedthrough
rlabel pdiffusion 444 -359 444 -359 0 feedthrough
rlabel pdiffusion 451 -359 451 -359 0 feedthrough
rlabel pdiffusion 458 -359 458 -359 0 feedthrough
rlabel pdiffusion 465 -359 465 -359 0 cellNo=384
rlabel pdiffusion 472 -359 472 -359 0 cellNo=17
rlabel pdiffusion 479 -359 479 -359 0 cellNo=267
rlabel pdiffusion 486 -359 486 -359 0 cellNo=130
rlabel pdiffusion 493 -359 493 -359 0 cellNo=1383
rlabel pdiffusion 500 -359 500 -359 0 feedthrough
rlabel pdiffusion 507 -359 507 -359 0 feedthrough
rlabel pdiffusion 514 -359 514 -359 0 cellNo=873
rlabel pdiffusion 521 -359 521 -359 0 feedthrough
rlabel pdiffusion 528 -359 528 -359 0 cellNo=93
rlabel pdiffusion 535 -359 535 -359 0 feedthrough
rlabel pdiffusion 542 -359 542 -359 0 feedthrough
rlabel pdiffusion 549 -359 549 -359 0 feedthrough
rlabel pdiffusion 556 -359 556 -359 0 feedthrough
rlabel pdiffusion 563 -359 563 -359 0 cellNo=774
rlabel pdiffusion 570 -359 570 -359 0 cellNo=283
rlabel pdiffusion 577 -359 577 -359 0 cellNo=884
rlabel pdiffusion 584 -359 584 -359 0 cellNo=731
rlabel pdiffusion 591 -359 591 -359 0 cellNo=622
rlabel pdiffusion 598 -359 598 -359 0 feedthrough
rlabel pdiffusion 605 -359 605 -359 0 cellNo=254
rlabel pdiffusion 612 -359 612 -359 0 feedthrough
rlabel pdiffusion 619 -359 619 -359 0 feedthrough
rlabel pdiffusion 626 -359 626 -359 0 feedthrough
rlabel pdiffusion 633 -359 633 -359 0 cellNo=54
rlabel pdiffusion 640 -359 640 -359 0 feedthrough
rlabel pdiffusion 647 -359 647 -359 0 feedthrough
rlabel pdiffusion 654 -359 654 -359 0 feedthrough
rlabel pdiffusion 661 -359 661 -359 0 cellNo=605
rlabel pdiffusion 668 -359 668 -359 0 feedthrough
rlabel pdiffusion 675 -359 675 -359 0 feedthrough
rlabel pdiffusion 682 -359 682 -359 0 cellNo=264
rlabel pdiffusion 689 -359 689 -359 0 feedthrough
rlabel pdiffusion 696 -359 696 -359 0 feedthrough
rlabel pdiffusion 703 -359 703 -359 0 feedthrough
rlabel pdiffusion 710 -359 710 -359 0 feedthrough
rlabel pdiffusion 717 -359 717 -359 0 cellNo=46
rlabel pdiffusion 724 -359 724 -359 0 cellNo=624
rlabel pdiffusion 731 -359 731 -359 0 feedthrough
rlabel pdiffusion 738 -359 738 -359 0 feedthrough
rlabel pdiffusion 745 -359 745 -359 0 feedthrough
rlabel pdiffusion 752 -359 752 -359 0 feedthrough
rlabel pdiffusion 759 -359 759 -359 0 feedthrough
rlabel pdiffusion 766 -359 766 -359 0 feedthrough
rlabel pdiffusion 773 -359 773 -359 0 cellNo=180
rlabel pdiffusion 780 -359 780 -359 0 feedthrough
rlabel pdiffusion 787 -359 787 -359 0 cellNo=233
rlabel pdiffusion 794 -359 794 -359 0 feedthrough
rlabel pdiffusion 801 -359 801 -359 0 feedthrough
rlabel pdiffusion 808 -359 808 -359 0 feedthrough
rlabel pdiffusion 815 -359 815 -359 0 feedthrough
rlabel pdiffusion 822 -359 822 -359 0 feedthrough
rlabel pdiffusion 829 -359 829 -359 0 feedthrough
rlabel pdiffusion 836 -359 836 -359 0 feedthrough
rlabel pdiffusion 843 -359 843 -359 0 feedthrough
rlabel pdiffusion 850 -359 850 -359 0 feedthrough
rlabel pdiffusion 857 -359 857 -359 0 feedthrough
rlabel pdiffusion 864 -359 864 -359 0 feedthrough
rlabel pdiffusion 871 -359 871 -359 0 feedthrough
rlabel pdiffusion 878 -359 878 -359 0 feedthrough
rlabel pdiffusion 885 -359 885 -359 0 feedthrough
rlabel pdiffusion 892 -359 892 -359 0 feedthrough
rlabel pdiffusion 899 -359 899 -359 0 feedthrough
rlabel pdiffusion 906 -359 906 -359 0 feedthrough
rlabel pdiffusion 913 -359 913 -359 0 feedthrough
rlabel pdiffusion 920 -359 920 -359 0 feedthrough
rlabel pdiffusion 927 -359 927 -359 0 feedthrough
rlabel pdiffusion 934 -359 934 -359 0 feedthrough
rlabel pdiffusion 941 -359 941 -359 0 feedthrough
rlabel pdiffusion 948 -359 948 -359 0 feedthrough
rlabel pdiffusion 955 -359 955 -359 0 feedthrough
rlabel pdiffusion 962 -359 962 -359 0 feedthrough
rlabel pdiffusion 969 -359 969 -359 0 feedthrough
rlabel pdiffusion 976 -359 976 -359 0 feedthrough
rlabel pdiffusion 983 -359 983 -359 0 feedthrough
rlabel pdiffusion 990 -359 990 -359 0 feedthrough
rlabel pdiffusion 997 -359 997 -359 0 feedthrough
rlabel pdiffusion 1004 -359 1004 -359 0 feedthrough
rlabel pdiffusion 1011 -359 1011 -359 0 feedthrough
rlabel pdiffusion 1018 -359 1018 -359 0 feedthrough
rlabel pdiffusion 1025 -359 1025 -359 0 feedthrough
rlabel pdiffusion 1032 -359 1032 -359 0 feedthrough
rlabel pdiffusion 1039 -359 1039 -359 0 feedthrough
rlabel pdiffusion 1046 -359 1046 -359 0 feedthrough
rlabel pdiffusion 1053 -359 1053 -359 0 feedthrough
rlabel pdiffusion 1060 -359 1060 -359 0 feedthrough
rlabel pdiffusion 1067 -359 1067 -359 0 feedthrough
rlabel pdiffusion 1074 -359 1074 -359 0 feedthrough
rlabel pdiffusion 1081 -359 1081 -359 0 feedthrough
rlabel pdiffusion 1088 -359 1088 -359 0 feedthrough
rlabel pdiffusion 1095 -359 1095 -359 0 feedthrough
rlabel pdiffusion 1102 -359 1102 -359 0 feedthrough
rlabel pdiffusion 1109 -359 1109 -359 0 feedthrough
rlabel pdiffusion 1116 -359 1116 -359 0 feedthrough
rlabel pdiffusion 1123 -359 1123 -359 0 feedthrough
rlabel pdiffusion 1130 -359 1130 -359 0 feedthrough
rlabel pdiffusion 1137 -359 1137 -359 0 feedthrough
rlabel pdiffusion 1144 -359 1144 -359 0 feedthrough
rlabel pdiffusion 1151 -359 1151 -359 0 feedthrough
rlabel pdiffusion 1158 -359 1158 -359 0 feedthrough
rlabel pdiffusion 1165 -359 1165 -359 0 feedthrough
rlabel pdiffusion 1172 -359 1172 -359 0 feedthrough
rlabel pdiffusion 1179 -359 1179 -359 0 feedthrough
rlabel pdiffusion 1186 -359 1186 -359 0 feedthrough
rlabel pdiffusion 1193 -359 1193 -359 0 feedthrough
rlabel pdiffusion 1200 -359 1200 -359 0 feedthrough
rlabel pdiffusion 1207 -359 1207 -359 0 feedthrough
rlabel pdiffusion 1214 -359 1214 -359 0 feedthrough
rlabel pdiffusion 1221 -359 1221 -359 0 feedthrough
rlabel pdiffusion 1228 -359 1228 -359 0 feedthrough
rlabel pdiffusion 1235 -359 1235 -359 0 feedthrough
rlabel pdiffusion 1242 -359 1242 -359 0 feedthrough
rlabel pdiffusion 1249 -359 1249 -359 0 feedthrough
rlabel pdiffusion 1256 -359 1256 -359 0 feedthrough
rlabel pdiffusion 1263 -359 1263 -359 0 feedthrough
rlabel pdiffusion 1270 -359 1270 -359 0 feedthrough
rlabel pdiffusion 1277 -359 1277 -359 0 feedthrough
rlabel pdiffusion 1284 -359 1284 -359 0 feedthrough
rlabel pdiffusion 1291 -359 1291 -359 0 feedthrough
rlabel pdiffusion 1298 -359 1298 -359 0 cellNo=5
rlabel pdiffusion 3 -484 3 -484 0 cellNo=1010
rlabel pdiffusion 10 -484 10 -484 0 cellNo=1210
rlabel pdiffusion 17 -484 17 -484 0 cellNo=1335
rlabel pdiffusion 24 -484 24 -484 0 cellNo=1217
rlabel pdiffusion 31 -484 31 -484 0 cellNo=1151
rlabel pdiffusion 38 -484 38 -484 0 cellNo=677
rlabel pdiffusion 45 -484 45 -484 0 cellNo=1233
rlabel pdiffusion 52 -484 52 -484 0 cellNo=1494
rlabel pdiffusion 59 -484 59 -484 0 cellNo=1250
rlabel pdiffusion 66 -484 66 -484 0 feedthrough
rlabel pdiffusion 73 -484 73 -484 0 feedthrough
rlabel pdiffusion 80 -484 80 -484 0 feedthrough
rlabel pdiffusion 87 -484 87 -484 0 feedthrough
rlabel pdiffusion 94 -484 94 -484 0 cellNo=944
rlabel pdiffusion 101 -484 101 -484 0 feedthrough
rlabel pdiffusion 108 -484 108 -484 0 feedthrough
rlabel pdiffusion 115 -484 115 -484 0 cellNo=1283
rlabel pdiffusion 122 -484 122 -484 0 cellNo=508
rlabel pdiffusion 129 -484 129 -484 0 cellNo=909
rlabel pdiffusion 136 -484 136 -484 0 feedthrough
rlabel pdiffusion 143 -484 143 -484 0 feedthrough
rlabel pdiffusion 150 -484 150 -484 0 cellNo=809
rlabel pdiffusion 157 -484 157 -484 0 feedthrough
rlabel pdiffusion 164 -484 164 -484 0 feedthrough
rlabel pdiffusion 171 -484 171 -484 0 feedthrough
rlabel pdiffusion 178 -484 178 -484 0 feedthrough
rlabel pdiffusion 185 -484 185 -484 0 feedthrough
rlabel pdiffusion 192 -484 192 -484 0 feedthrough
rlabel pdiffusion 199 -484 199 -484 0 feedthrough
rlabel pdiffusion 206 -484 206 -484 0 feedthrough
rlabel pdiffusion 213 -484 213 -484 0 cellNo=245
rlabel pdiffusion 220 -484 220 -484 0 feedthrough
rlabel pdiffusion 227 -484 227 -484 0 feedthrough
rlabel pdiffusion 234 -484 234 -484 0 feedthrough
rlabel pdiffusion 241 -484 241 -484 0 feedthrough
rlabel pdiffusion 248 -484 248 -484 0 feedthrough
rlabel pdiffusion 255 -484 255 -484 0 feedthrough
rlabel pdiffusion 262 -484 262 -484 0 feedthrough
rlabel pdiffusion 269 -484 269 -484 0 cellNo=758
rlabel pdiffusion 276 -484 276 -484 0 cellNo=1292
rlabel pdiffusion 283 -484 283 -484 0 cellNo=1324
rlabel pdiffusion 290 -484 290 -484 0 cellNo=1365
rlabel pdiffusion 297 -484 297 -484 0 feedthrough
rlabel pdiffusion 304 -484 304 -484 0 feedthrough
rlabel pdiffusion 311 -484 311 -484 0 feedthrough
rlabel pdiffusion 318 -484 318 -484 0 feedthrough
rlabel pdiffusion 325 -484 325 -484 0 feedthrough
rlabel pdiffusion 332 -484 332 -484 0 feedthrough
rlabel pdiffusion 339 -484 339 -484 0 feedthrough
rlabel pdiffusion 346 -484 346 -484 0 feedthrough
rlabel pdiffusion 353 -484 353 -484 0 cellNo=18
rlabel pdiffusion 360 -484 360 -484 0 feedthrough
rlabel pdiffusion 367 -484 367 -484 0 feedthrough
rlabel pdiffusion 374 -484 374 -484 0 feedthrough
rlabel pdiffusion 381 -484 381 -484 0 feedthrough
rlabel pdiffusion 388 -484 388 -484 0 feedthrough
rlabel pdiffusion 395 -484 395 -484 0 feedthrough
rlabel pdiffusion 402 -484 402 -484 0 feedthrough
rlabel pdiffusion 409 -484 409 -484 0 feedthrough
rlabel pdiffusion 416 -484 416 -484 0 feedthrough
rlabel pdiffusion 423 -484 423 -484 0 feedthrough
rlabel pdiffusion 430 -484 430 -484 0 feedthrough
rlabel pdiffusion 437 -484 437 -484 0 feedthrough
rlabel pdiffusion 444 -484 444 -484 0 feedthrough
rlabel pdiffusion 451 -484 451 -484 0 feedthrough
rlabel pdiffusion 458 -484 458 -484 0 cellNo=910
rlabel pdiffusion 465 -484 465 -484 0 feedthrough
rlabel pdiffusion 472 -484 472 -484 0 feedthrough
rlabel pdiffusion 479 -484 479 -484 0 feedthrough
rlabel pdiffusion 486 -484 486 -484 0 feedthrough
rlabel pdiffusion 493 -484 493 -484 0 feedthrough
rlabel pdiffusion 500 -484 500 -484 0 cellNo=342
rlabel pdiffusion 507 -484 507 -484 0 feedthrough
rlabel pdiffusion 514 -484 514 -484 0 cellNo=769
rlabel pdiffusion 521 -484 521 -484 0 feedthrough
rlabel pdiffusion 528 -484 528 -484 0 feedthrough
rlabel pdiffusion 535 -484 535 -484 0 cellNo=313
rlabel pdiffusion 542 -484 542 -484 0 feedthrough
rlabel pdiffusion 549 -484 549 -484 0 feedthrough
rlabel pdiffusion 556 -484 556 -484 0 cellNo=224
rlabel pdiffusion 563 -484 563 -484 0 feedthrough
rlabel pdiffusion 570 -484 570 -484 0 feedthrough
rlabel pdiffusion 577 -484 577 -484 0 cellNo=2
rlabel pdiffusion 584 -484 584 -484 0 feedthrough
rlabel pdiffusion 591 -484 591 -484 0 feedthrough
rlabel pdiffusion 598 -484 598 -484 0 cellNo=66
rlabel pdiffusion 605 -484 605 -484 0 feedthrough
rlabel pdiffusion 612 -484 612 -484 0 cellNo=829
rlabel pdiffusion 619 -484 619 -484 0 feedthrough
rlabel pdiffusion 626 -484 626 -484 0 feedthrough
rlabel pdiffusion 633 -484 633 -484 0 cellNo=227
rlabel pdiffusion 640 -484 640 -484 0 cellNo=586
rlabel pdiffusion 647 -484 647 -484 0 feedthrough
rlabel pdiffusion 654 -484 654 -484 0 feedthrough
rlabel pdiffusion 661 -484 661 -484 0 feedthrough
rlabel pdiffusion 668 -484 668 -484 0 feedthrough
rlabel pdiffusion 675 -484 675 -484 0 cellNo=108
rlabel pdiffusion 682 -484 682 -484 0 cellNo=386
rlabel pdiffusion 689 -484 689 -484 0 cellNo=604
rlabel pdiffusion 696 -484 696 -484 0 cellNo=422
rlabel pdiffusion 703 -484 703 -484 0 feedthrough
rlabel pdiffusion 710 -484 710 -484 0 feedthrough
rlabel pdiffusion 717 -484 717 -484 0 cellNo=176
rlabel pdiffusion 724 -484 724 -484 0 feedthrough
rlabel pdiffusion 731 -484 731 -484 0 feedthrough
rlabel pdiffusion 738 -484 738 -484 0 feedthrough
rlabel pdiffusion 745 -484 745 -484 0 feedthrough
rlabel pdiffusion 752 -484 752 -484 0 cellNo=824
rlabel pdiffusion 759 -484 759 -484 0 cellNo=673
rlabel pdiffusion 766 -484 766 -484 0 feedthrough
rlabel pdiffusion 773 -484 773 -484 0 cellNo=125
rlabel pdiffusion 780 -484 780 -484 0 feedthrough
rlabel pdiffusion 787 -484 787 -484 0 cellNo=414
rlabel pdiffusion 794 -484 794 -484 0 feedthrough
rlabel pdiffusion 801 -484 801 -484 0 feedthrough
rlabel pdiffusion 808 -484 808 -484 0 feedthrough
rlabel pdiffusion 815 -484 815 -484 0 feedthrough
rlabel pdiffusion 822 -484 822 -484 0 feedthrough
rlabel pdiffusion 829 -484 829 -484 0 cellNo=660
rlabel pdiffusion 836 -484 836 -484 0 feedthrough
rlabel pdiffusion 843 -484 843 -484 0 feedthrough
rlabel pdiffusion 850 -484 850 -484 0 feedthrough
rlabel pdiffusion 857 -484 857 -484 0 feedthrough
rlabel pdiffusion 864 -484 864 -484 0 feedthrough
rlabel pdiffusion 871 -484 871 -484 0 feedthrough
rlabel pdiffusion 878 -484 878 -484 0 feedthrough
rlabel pdiffusion 885 -484 885 -484 0 cellNo=295
rlabel pdiffusion 892 -484 892 -484 0 feedthrough
rlabel pdiffusion 899 -484 899 -484 0 feedthrough
rlabel pdiffusion 906 -484 906 -484 0 feedthrough
rlabel pdiffusion 913 -484 913 -484 0 feedthrough
rlabel pdiffusion 920 -484 920 -484 0 feedthrough
rlabel pdiffusion 927 -484 927 -484 0 feedthrough
rlabel pdiffusion 934 -484 934 -484 0 feedthrough
rlabel pdiffusion 941 -484 941 -484 0 feedthrough
rlabel pdiffusion 948 -484 948 -484 0 feedthrough
rlabel pdiffusion 955 -484 955 -484 0 feedthrough
rlabel pdiffusion 962 -484 962 -484 0 feedthrough
rlabel pdiffusion 969 -484 969 -484 0 feedthrough
rlabel pdiffusion 976 -484 976 -484 0 feedthrough
rlabel pdiffusion 983 -484 983 -484 0 feedthrough
rlabel pdiffusion 990 -484 990 -484 0 feedthrough
rlabel pdiffusion 997 -484 997 -484 0 feedthrough
rlabel pdiffusion 1004 -484 1004 -484 0 feedthrough
rlabel pdiffusion 1011 -484 1011 -484 0 feedthrough
rlabel pdiffusion 1018 -484 1018 -484 0 feedthrough
rlabel pdiffusion 1025 -484 1025 -484 0 feedthrough
rlabel pdiffusion 1032 -484 1032 -484 0 feedthrough
rlabel pdiffusion 1039 -484 1039 -484 0 feedthrough
rlabel pdiffusion 1046 -484 1046 -484 0 feedthrough
rlabel pdiffusion 1053 -484 1053 -484 0 feedthrough
rlabel pdiffusion 1060 -484 1060 -484 0 feedthrough
rlabel pdiffusion 1067 -484 1067 -484 0 feedthrough
rlabel pdiffusion 1074 -484 1074 -484 0 feedthrough
rlabel pdiffusion 1081 -484 1081 -484 0 feedthrough
rlabel pdiffusion 1088 -484 1088 -484 0 feedthrough
rlabel pdiffusion 1095 -484 1095 -484 0 feedthrough
rlabel pdiffusion 1102 -484 1102 -484 0 feedthrough
rlabel pdiffusion 1109 -484 1109 -484 0 feedthrough
rlabel pdiffusion 1116 -484 1116 -484 0 feedthrough
rlabel pdiffusion 1123 -484 1123 -484 0 feedthrough
rlabel pdiffusion 1130 -484 1130 -484 0 feedthrough
rlabel pdiffusion 1137 -484 1137 -484 0 feedthrough
rlabel pdiffusion 1144 -484 1144 -484 0 feedthrough
rlabel pdiffusion 1151 -484 1151 -484 0 feedthrough
rlabel pdiffusion 1158 -484 1158 -484 0 feedthrough
rlabel pdiffusion 1165 -484 1165 -484 0 feedthrough
rlabel pdiffusion 1172 -484 1172 -484 0 feedthrough
rlabel pdiffusion 1179 -484 1179 -484 0 feedthrough
rlabel pdiffusion 1186 -484 1186 -484 0 feedthrough
rlabel pdiffusion 1193 -484 1193 -484 0 feedthrough
rlabel pdiffusion 1200 -484 1200 -484 0 feedthrough
rlabel pdiffusion 1207 -484 1207 -484 0 feedthrough
rlabel pdiffusion 1214 -484 1214 -484 0 feedthrough
rlabel pdiffusion 1221 -484 1221 -484 0 feedthrough
rlabel pdiffusion 1228 -484 1228 -484 0 feedthrough
rlabel pdiffusion 1235 -484 1235 -484 0 feedthrough
rlabel pdiffusion 1242 -484 1242 -484 0 feedthrough
rlabel pdiffusion 1249 -484 1249 -484 0 feedthrough
rlabel pdiffusion 1256 -484 1256 -484 0 feedthrough
rlabel pdiffusion 1263 -484 1263 -484 0 feedthrough
rlabel pdiffusion 1270 -484 1270 -484 0 feedthrough
rlabel pdiffusion 1277 -484 1277 -484 0 feedthrough
rlabel pdiffusion 1284 -484 1284 -484 0 feedthrough
rlabel pdiffusion 1291 -484 1291 -484 0 feedthrough
rlabel pdiffusion 1298 -484 1298 -484 0 feedthrough
rlabel pdiffusion 1305 -484 1305 -484 0 feedthrough
rlabel pdiffusion 1312 -484 1312 -484 0 feedthrough
rlabel pdiffusion 1319 -484 1319 -484 0 feedthrough
rlabel pdiffusion 1326 -484 1326 -484 0 feedthrough
rlabel pdiffusion 1333 -484 1333 -484 0 feedthrough
rlabel pdiffusion 1340 -484 1340 -484 0 feedthrough
rlabel pdiffusion 1347 -484 1347 -484 0 feedthrough
rlabel pdiffusion 1354 -484 1354 -484 0 feedthrough
rlabel pdiffusion 1361 -484 1361 -484 0 feedthrough
rlabel pdiffusion 1368 -484 1368 -484 0 feedthrough
rlabel pdiffusion 1375 -484 1375 -484 0 cellNo=175
rlabel pdiffusion 3 -617 3 -617 0 cellNo=1009
rlabel pdiffusion 10 -617 10 -617 0 cellNo=1111
rlabel pdiffusion 17 -617 17 -617 0 cellNo=1282
rlabel pdiffusion 24 -617 24 -617 0 cellNo=1012
rlabel pdiffusion 31 -617 31 -617 0 cellNo=1105
rlabel pdiffusion 38 -617 38 -617 0 cellNo=216
rlabel pdiffusion 45 -617 45 -617 0 cellNo=1275
rlabel pdiffusion 52 -617 52 -617 0 feedthrough
rlabel pdiffusion 59 -617 59 -617 0 feedthrough
rlabel pdiffusion 66 -617 66 -617 0 cellNo=634
rlabel pdiffusion 73 -617 73 -617 0 feedthrough
rlabel pdiffusion 80 -617 80 -617 0 cellNo=761
rlabel pdiffusion 87 -617 87 -617 0 feedthrough
rlabel pdiffusion 94 -617 94 -617 0 cellNo=1129
rlabel pdiffusion 101 -617 101 -617 0 feedthrough
rlabel pdiffusion 108 -617 108 -617 0 feedthrough
rlabel pdiffusion 115 -617 115 -617 0 cellNo=610
rlabel pdiffusion 122 -617 122 -617 0 feedthrough
rlabel pdiffusion 129 -617 129 -617 0 feedthrough
rlabel pdiffusion 136 -617 136 -617 0 cellNo=127
rlabel pdiffusion 143 -617 143 -617 0 feedthrough
rlabel pdiffusion 150 -617 150 -617 0 cellNo=481
rlabel pdiffusion 157 -617 157 -617 0 cellNo=63
rlabel pdiffusion 164 -617 164 -617 0 feedthrough
rlabel pdiffusion 171 -617 171 -617 0 cellNo=1364
rlabel pdiffusion 178 -617 178 -617 0 feedthrough
rlabel pdiffusion 185 -617 185 -617 0 feedthrough
rlabel pdiffusion 192 -617 192 -617 0 feedthrough
rlabel pdiffusion 199 -617 199 -617 0 cellNo=685
rlabel pdiffusion 206 -617 206 -617 0 feedthrough
rlabel pdiffusion 213 -617 213 -617 0 feedthrough
rlabel pdiffusion 220 -617 220 -617 0 cellNo=373
rlabel pdiffusion 227 -617 227 -617 0 feedthrough
rlabel pdiffusion 234 -617 234 -617 0 cellNo=1323
rlabel pdiffusion 241 -617 241 -617 0 cellNo=755
rlabel pdiffusion 248 -617 248 -617 0 cellNo=919
rlabel pdiffusion 255 -617 255 -617 0 cellNo=1289
rlabel pdiffusion 262 -617 262 -617 0 feedthrough
rlabel pdiffusion 269 -617 269 -617 0 feedthrough
rlabel pdiffusion 276 -617 276 -617 0 feedthrough
rlabel pdiffusion 283 -617 283 -617 0 feedthrough
rlabel pdiffusion 290 -617 290 -617 0 feedthrough
rlabel pdiffusion 297 -617 297 -617 0 feedthrough
rlabel pdiffusion 304 -617 304 -617 0 feedthrough
rlabel pdiffusion 311 -617 311 -617 0 feedthrough
rlabel pdiffusion 318 -617 318 -617 0 feedthrough
rlabel pdiffusion 325 -617 325 -617 0 feedthrough
rlabel pdiffusion 332 -617 332 -617 0 feedthrough
rlabel pdiffusion 339 -617 339 -617 0 feedthrough
rlabel pdiffusion 346 -617 346 -617 0 feedthrough
rlabel pdiffusion 353 -617 353 -617 0 feedthrough
rlabel pdiffusion 360 -617 360 -617 0 feedthrough
rlabel pdiffusion 367 -617 367 -617 0 cellNo=1403
rlabel pdiffusion 374 -617 374 -617 0 feedthrough
rlabel pdiffusion 381 -617 381 -617 0 feedthrough
rlabel pdiffusion 388 -617 388 -617 0 feedthrough
rlabel pdiffusion 395 -617 395 -617 0 cellNo=358
rlabel pdiffusion 402 -617 402 -617 0 feedthrough
rlabel pdiffusion 409 -617 409 -617 0 feedthrough
rlabel pdiffusion 416 -617 416 -617 0 feedthrough
rlabel pdiffusion 423 -617 423 -617 0 feedthrough
rlabel pdiffusion 430 -617 430 -617 0 feedthrough
rlabel pdiffusion 437 -617 437 -617 0 feedthrough
rlabel pdiffusion 444 -617 444 -617 0 feedthrough
rlabel pdiffusion 451 -617 451 -617 0 feedthrough
rlabel pdiffusion 458 -617 458 -617 0 feedthrough
rlabel pdiffusion 465 -617 465 -617 0 feedthrough
rlabel pdiffusion 472 -617 472 -617 0 feedthrough
rlabel pdiffusion 479 -617 479 -617 0 feedthrough
rlabel pdiffusion 486 -617 486 -617 0 feedthrough
rlabel pdiffusion 493 -617 493 -617 0 feedthrough
rlabel pdiffusion 500 -617 500 -617 0 cellNo=110
rlabel pdiffusion 507 -617 507 -617 0 feedthrough
rlabel pdiffusion 514 -617 514 -617 0 cellNo=330
rlabel pdiffusion 521 -617 521 -617 0 feedthrough
rlabel pdiffusion 528 -617 528 -617 0 cellNo=583
rlabel pdiffusion 535 -617 535 -617 0 feedthrough
rlabel pdiffusion 542 -617 542 -617 0 cellNo=666
rlabel pdiffusion 549 -617 549 -617 0 feedthrough
rlabel pdiffusion 556 -617 556 -617 0 feedthrough
rlabel pdiffusion 563 -617 563 -617 0 feedthrough
rlabel pdiffusion 570 -617 570 -617 0 feedthrough
rlabel pdiffusion 577 -617 577 -617 0 feedthrough
rlabel pdiffusion 584 -617 584 -617 0 cellNo=825
rlabel pdiffusion 591 -617 591 -617 0 feedthrough
rlabel pdiffusion 598 -617 598 -617 0 feedthrough
rlabel pdiffusion 605 -617 605 -617 0 feedthrough
rlabel pdiffusion 612 -617 612 -617 0 feedthrough
rlabel pdiffusion 619 -617 619 -617 0 feedthrough
rlabel pdiffusion 626 -617 626 -617 0 feedthrough
rlabel pdiffusion 633 -617 633 -617 0 feedthrough
rlabel pdiffusion 640 -617 640 -617 0 feedthrough
rlabel pdiffusion 647 -617 647 -617 0 feedthrough
rlabel pdiffusion 654 -617 654 -617 0 feedthrough
rlabel pdiffusion 661 -617 661 -617 0 feedthrough
rlabel pdiffusion 668 -617 668 -617 0 cellNo=559
rlabel pdiffusion 675 -617 675 -617 0 feedthrough
rlabel pdiffusion 682 -617 682 -617 0 cellNo=193
rlabel pdiffusion 689 -617 689 -617 0 feedthrough
rlabel pdiffusion 696 -617 696 -617 0 cellNo=861
rlabel pdiffusion 703 -617 703 -617 0 cellNo=266
rlabel pdiffusion 710 -617 710 -617 0 feedthrough
rlabel pdiffusion 717 -617 717 -617 0 cellNo=716
rlabel pdiffusion 724 -617 724 -617 0 feedthrough
rlabel pdiffusion 731 -617 731 -617 0 cellNo=783
rlabel pdiffusion 738 -617 738 -617 0 feedthrough
rlabel pdiffusion 745 -617 745 -617 0 feedthrough
rlabel pdiffusion 752 -617 752 -617 0 feedthrough
rlabel pdiffusion 759 -617 759 -617 0 feedthrough
rlabel pdiffusion 766 -617 766 -617 0 cellNo=337
rlabel pdiffusion 773 -617 773 -617 0 cellNo=847
rlabel pdiffusion 780 -617 780 -617 0 cellNo=511
rlabel pdiffusion 787 -617 787 -617 0 feedthrough
rlabel pdiffusion 794 -617 794 -617 0 cellNo=550
rlabel pdiffusion 801 -617 801 -617 0 feedthrough
rlabel pdiffusion 808 -617 808 -617 0 cellNo=554
rlabel pdiffusion 815 -617 815 -617 0 feedthrough
rlabel pdiffusion 822 -617 822 -617 0 feedthrough
rlabel pdiffusion 829 -617 829 -617 0 feedthrough
rlabel pdiffusion 836 -617 836 -617 0 feedthrough
rlabel pdiffusion 843 -617 843 -617 0 feedthrough
rlabel pdiffusion 850 -617 850 -617 0 feedthrough
rlabel pdiffusion 857 -617 857 -617 0 feedthrough
rlabel pdiffusion 864 -617 864 -617 0 feedthrough
rlabel pdiffusion 871 -617 871 -617 0 feedthrough
rlabel pdiffusion 878 -617 878 -617 0 feedthrough
rlabel pdiffusion 885 -617 885 -617 0 feedthrough
rlabel pdiffusion 892 -617 892 -617 0 feedthrough
rlabel pdiffusion 899 -617 899 -617 0 cellNo=377
rlabel pdiffusion 906 -617 906 -617 0 feedthrough
rlabel pdiffusion 913 -617 913 -617 0 feedthrough
rlabel pdiffusion 920 -617 920 -617 0 feedthrough
rlabel pdiffusion 927 -617 927 -617 0 feedthrough
rlabel pdiffusion 934 -617 934 -617 0 feedthrough
rlabel pdiffusion 941 -617 941 -617 0 feedthrough
rlabel pdiffusion 948 -617 948 -617 0 feedthrough
rlabel pdiffusion 955 -617 955 -617 0 feedthrough
rlabel pdiffusion 962 -617 962 -617 0 feedthrough
rlabel pdiffusion 969 -617 969 -617 0 feedthrough
rlabel pdiffusion 976 -617 976 -617 0 cellNo=667
rlabel pdiffusion 983 -617 983 -617 0 feedthrough
rlabel pdiffusion 990 -617 990 -617 0 feedthrough
rlabel pdiffusion 997 -617 997 -617 0 feedthrough
rlabel pdiffusion 1004 -617 1004 -617 0 feedthrough
rlabel pdiffusion 1011 -617 1011 -617 0 feedthrough
rlabel pdiffusion 1018 -617 1018 -617 0 feedthrough
rlabel pdiffusion 1025 -617 1025 -617 0 feedthrough
rlabel pdiffusion 1032 -617 1032 -617 0 feedthrough
rlabel pdiffusion 1039 -617 1039 -617 0 feedthrough
rlabel pdiffusion 1046 -617 1046 -617 0 feedthrough
rlabel pdiffusion 1053 -617 1053 -617 0 feedthrough
rlabel pdiffusion 1060 -617 1060 -617 0 feedthrough
rlabel pdiffusion 1067 -617 1067 -617 0 feedthrough
rlabel pdiffusion 1074 -617 1074 -617 0 feedthrough
rlabel pdiffusion 1081 -617 1081 -617 0 feedthrough
rlabel pdiffusion 1088 -617 1088 -617 0 feedthrough
rlabel pdiffusion 1095 -617 1095 -617 0 feedthrough
rlabel pdiffusion 1102 -617 1102 -617 0 feedthrough
rlabel pdiffusion 1109 -617 1109 -617 0 feedthrough
rlabel pdiffusion 1116 -617 1116 -617 0 feedthrough
rlabel pdiffusion 1123 -617 1123 -617 0 feedthrough
rlabel pdiffusion 1130 -617 1130 -617 0 feedthrough
rlabel pdiffusion 1137 -617 1137 -617 0 feedthrough
rlabel pdiffusion 1144 -617 1144 -617 0 feedthrough
rlabel pdiffusion 1151 -617 1151 -617 0 feedthrough
rlabel pdiffusion 1158 -617 1158 -617 0 feedthrough
rlabel pdiffusion 1165 -617 1165 -617 0 feedthrough
rlabel pdiffusion 1172 -617 1172 -617 0 feedthrough
rlabel pdiffusion 1179 -617 1179 -617 0 feedthrough
rlabel pdiffusion 1186 -617 1186 -617 0 feedthrough
rlabel pdiffusion 1193 -617 1193 -617 0 feedthrough
rlabel pdiffusion 1200 -617 1200 -617 0 feedthrough
rlabel pdiffusion 1207 -617 1207 -617 0 feedthrough
rlabel pdiffusion 1214 -617 1214 -617 0 feedthrough
rlabel pdiffusion 1221 -617 1221 -617 0 feedthrough
rlabel pdiffusion 1228 -617 1228 -617 0 feedthrough
rlabel pdiffusion 1235 -617 1235 -617 0 feedthrough
rlabel pdiffusion 1242 -617 1242 -617 0 feedthrough
rlabel pdiffusion 1249 -617 1249 -617 0 feedthrough
rlabel pdiffusion 1256 -617 1256 -617 0 feedthrough
rlabel pdiffusion 1263 -617 1263 -617 0 feedthrough
rlabel pdiffusion 1270 -617 1270 -617 0 feedthrough
rlabel pdiffusion 1277 -617 1277 -617 0 feedthrough
rlabel pdiffusion 1284 -617 1284 -617 0 feedthrough
rlabel pdiffusion 1291 -617 1291 -617 0 feedthrough
rlabel pdiffusion 1298 -617 1298 -617 0 feedthrough
rlabel pdiffusion 1305 -617 1305 -617 0 feedthrough
rlabel pdiffusion 1312 -617 1312 -617 0 feedthrough
rlabel pdiffusion 1319 -617 1319 -617 0 feedthrough
rlabel pdiffusion 1326 -617 1326 -617 0 feedthrough
rlabel pdiffusion 1333 -617 1333 -617 0 feedthrough
rlabel pdiffusion 1340 -617 1340 -617 0 feedthrough
rlabel pdiffusion 1347 -617 1347 -617 0 feedthrough
rlabel pdiffusion 1354 -617 1354 -617 0 cellNo=4
rlabel pdiffusion 1361 -617 1361 -617 0 feedthrough
rlabel pdiffusion 1368 -617 1368 -617 0 feedthrough
rlabel pdiffusion 1375 -617 1375 -617 0 feedthrough
rlabel pdiffusion 1382 -617 1382 -617 0 feedthrough
rlabel pdiffusion 1389 -617 1389 -617 0 feedthrough
rlabel pdiffusion 1473 -617 1473 -617 0 feedthrough
rlabel pdiffusion 3 -740 3 -740 0 cellNo=1127
rlabel pdiffusion 10 -740 10 -740 0 cellNo=1333
rlabel pdiffusion 17 -740 17 -740 0 cellNo=1291
rlabel pdiffusion 24 -740 24 -740 0 cellNo=1321
rlabel pdiffusion 31 -740 31 -740 0 cellNo=1408
rlabel pdiffusion 38 -740 38 -740 0 cellNo=1285
rlabel pdiffusion 45 -740 45 -740 0 feedthrough
rlabel pdiffusion 52 -740 52 -740 0 feedthrough
rlabel pdiffusion 59 -740 59 -740 0 feedthrough
rlabel pdiffusion 66 -740 66 -740 0 feedthrough
rlabel pdiffusion 73 -740 73 -740 0 feedthrough
rlabel pdiffusion 80 -740 80 -740 0 cellNo=248
rlabel pdiffusion 87 -740 87 -740 0 feedthrough
rlabel pdiffusion 94 -740 94 -740 0 cellNo=81
rlabel pdiffusion 101 -740 101 -740 0 feedthrough
rlabel pdiffusion 108 -740 108 -740 0 feedthrough
rlabel pdiffusion 115 -740 115 -740 0 feedthrough
rlabel pdiffusion 122 -740 122 -740 0 cellNo=407
rlabel pdiffusion 129 -740 129 -740 0 feedthrough
rlabel pdiffusion 136 -740 136 -740 0 feedthrough
rlabel pdiffusion 143 -740 143 -740 0 cellNo=1420
rlabel pdiffusion 150 -740 150 -740 0 feedthrough
rlabel pdiffusion 157 -740 157 -740 0 feedthrough
rlabel pdiffusion 164 -740 164 -740 0 feedthrough
rlabel pdiffusion 171 -740 171 -740 0 feedthrough
rlabel pdiffusion 178 -740 178 -740 0 feedthrough
rlabel pdiffusion 185 -740 185 -740 0 cellNo=32
rlabel pdiffusion 192 -740 192 -740 0 feedthrough
rlabel pdiffusion 199 -740 199 -740 0 feedthrough
rlabel pdiffusion 206 -740 206 -740 0 feedthrough
rlabel pdiffusion 213 -740 213 -740 0 feedthrough
rlabel pdiffusion 220 -740 220 -740 0 feedthrough
rlabel pdiffusion 227 -740 227 -740 0 feedthrough
rlabel pdiffusion 234 -740 234 -740 0 feedthrough
rlabel pdiffusion 241 -740 241 -740 0 feedthrough
rlabel pdiffusion 248 -740 248 -740 0 cellNo=656
rlabel pdiffusion 255 -740 255 -740 0 feedthrough
rlabel pdiffusion 262 -740 262 -740 0 feedthrough
rlabel pdiffusion 269 -740 269 -740 0 feedthrough
rlabel pdiffusion 276 -740 276 -740 0 cellNo=209
rlabel pdiffusion 283 -740 283 -740 0 feedthrough
rlabel pdiffusion 290 -740 290 -740 0 cellNo=639
rlabel pdiffusion 297 -740 297 -740 0 feedthrough
rlabel pdiffusion 304 -740 304 -740 0 feedthrough
rlabel pdiffusion 311 -740 311 -740 0 feedthrough
rlabel pdiffusion 318 -740 318 -740 0 feedthrough
rlabel pdiffusion 325 -740 325 -740 0 feedthrough
rlabel pdiffusion 332 -740 332 -740 0 feedthrough
rlabel pdiffusion 339 -740 339 -740 0 feedthrough
rlabel pdiffusion 346 -740 346 -740 0 feedthrough
rlabel pdiffusion 353 -740 353 -740 0 feedthrough
rlabel pdiffusion 360 -740 360 -740 0 feedthrough
rlabel pdiffusion 367 -740 367 -740 0 feedthrough
rlabel pdiffusion 374 -740 374 -740 0 feedthrough
rlabel pdiffusion 381 -740 381 -740 0 feedthrough
rlabel pdiffusion 388 -740 388 -740 0 feedthrough
rlabel pdiffusion 395 -740 395 -740 0 feedthrough
rlabel pdiffusion 402 -740 402 -740 0 feedthrough
rlabel pdiffusion 409 -740 409 -740 0 feedthrough
rlabel pdiffusion 416 -740 416 -740 0 feedthrough
rlabel pdiffusion 423 -740 423 -740 0 feedthrough
rlabel pdiffusion 430 -740 430 -740 0 cellNo=287
rlabel pdiffusion 437 -740 437 -740 0 cellNo=686
rlabel pdiffusion 444 -740 444 -740 0 feedthrough
rlabel pdiffusion 451 -740 451 -740 0 feedthrough
rlabel pdiffusion 458 -740 458 -740 0 feedthrough
rlabel pdiffusion 465 -740 465 -740 0 feedthrough
rlabel pdiffusion 472 -740 472 -740 0 feedthrough
rlabel pdiffusion 479 -740 479 -740 0 feedthrough
rlabel pdiffusion 486 -740 486 -740 0 cellNo=279
rlabel pdiffusion 493 -740 493 -740 0 feedthrough
rlabel pdiffusion 500 -740 500 -740 0 cellNo=1295
rlabel pdiffusion 507 -740 507 -740 0 feedthrough
rlabel pdiffusion 514 -740 514 -740 0 feedthrough
rlabel pdiffusion 521 -740 521 -740 0 feedthrough
rlabel pdiffusion 528 -740 528 -740 0 feedthrough
rlabel pdiffusion 535 -740 535 -740 0 cellNo=475
rlabel pdiffusion 542 -740 542 -740 0 feedthrough
rlabel pdiffusion 549 -740 549 -740 0 feedthrough
rlabel pdiffusion 556 -740 556 -740 0 cellNo=364
rlabel pdiffusion 563 -740 563 -740 0 cellNo=740
rlabel pdiffusion 570 -740 570 -740 0 feedthrough
rlabel pdiffusion 577 -740 577 -740 0 cellNo=350
rlabel pdiffusion 584 -740 584 -740 0 feedthrough
rlabel pdiffusion 591 -740 591 -740 0 cellNo=138
rlabel pdiffusion 598 -740 598 -740 0 feedthrough
rlabel pdiffusion 605 -740 605 -740 0 cellNo=122
rlabel pdiffusion 612 -740 612 -740 0 feedthrough
rlabel pdiffusion 619 -740 619 -740 0 feedthrough
rlabel pdiffusion 626 -740 626 -740 0 feedthrough
rlabel pdiffusion 633 -740 633 -740 0 cellNo=1384
rlabel pdiffusion 640 -740 640 -740 0 feedthrough
rlabel pdiffusion 647 -740 647 -740 0 cellNo=503
rlabel pdiffusion 654 -740 654 -740 0 cellNo=174
rlabel pdiffusion 661 -740 661 -740 0 feedthrough
rlabel pdiffusion 668 -740 668 -740 0 feedthrough
rlabel pdiffusion 675 -740 675 -740 0 feedthrough
rlabel pdiffusion 682 -740 682 -740 0 feedthrough
rlabel pdiffusion 689 -740 689 -740 0 feedthrough
rlabel pdiffusion 696 -740 696 -740 0 feedthrough
rlabel pdiffusion 703 -740 703 -740 0 feedthrough
rlabel pdiffusion 710 -740 710 -740 0 cellNo=141
rlabel pdiffusion 717 -740 717 -740 0 feedthrough
rlabel pdiffusion 724 -740 724 -740 0 cellNo=58
rlabel pdiffusion 731 -740 731 -740 0 cellNo=869
rlabel pdiffusion 738 -740 738 -740 0 feedthrough
rlabel pdiffusion 745 -740 745 -740 0 feedthrough
rlabel pdiffusion 752 -740 752 -740 0 feedthrough
rlabel pdiffusion 759 -740 759 -740 0 feedthrough
rlabel pdiffusion 766 -740 766 -740 0 feedthrough
rlabel pdiffusion 773 -740 773 -740 0 feedthrough
rlabel pdiffusion 780 -740 780 -740 0 feedthrough
rlabel pdiffusion 787 -740 787 -740 0 feedthrough
rlabel pdiffusion 794 -740 794 -740 0 cellNo=822
rlabel pdiffusion 801 -740 801 -740 0 feedthrough
rlabel pdiffusion 808 -740 808 -740 0 feedthrough
rlabel pdiffusion 815 -740 815 -740 0 feedthrough
rlabel pdiffusion 822 -740 822 -740 0 feedthrough
rlabel pdiffusion 829 -740 829 -740 0 cellNo=494
rlabel pdiffusion 836 -740 836 -740 0 feedthrough
rlabel pdiffusion 843 -740 843 -740 0 feedthrough
rlabel pdiffusion 850 -740 850 -740 0 feedthrough
rlabel pdiffusion 857 -740 857 -740 0 cellNo=464
rlabel pdiffusion 864 -740 864 -740 0 feedthrough
rlabel pdiffusion 871 -740 871 -740 0 cellNo=262
rlabel pdiffusion 878 -740 878 -740 0 feedthrough
rlabel pdiffusion 885 -740 885 -740 0 cellNo=368
rlabel pdiffusion 892 -740 892 -740 0 feedthrough
rlabel pdiffusion 899 -740 899 -740 0 feedthrough
rlabel pdiffusion 906 -740 906 -740 0 cellNo=590
rlabel pdiffusion 913 -740 913 -740 0 cellNo=888
rlabel pdiffusion 920 -740 920 -740 0 cellNo=591
rlabel pdiffusion 927 -740 927 -740 0 feedthrough
rlabel pdiffusion 934 -740 934 -740 0 feedthrough
rlabel pdiffusion 941 -740 941 -740 0 feedthrough
rlabel pdiffusion 948 -740 948 -740 0 feedthrough
rlabel pdiffusion 955 -740 955 -740 0 feedthrough
rlabel pdiffusion 962 -740 962 -740 0 feedthrough
rlabel pdiffusion 969 -740 969 -740 0 feedthrough
rlabel pdiffusion 976 -740 976 -740 0 feedthrough
rlabel pdiffusion 983 -740 983 -740 0 feedthrough
rlabel pdiffusion 990 -740 990 -740 0 cellNo=347
rlabel pdiffusion 997 -740 997 -740 0 feedthrough
rlabel pdiffusion 1004 -740 1004 -740 0 cellNo=947
rlabel pdiffusion 1011 -740 1011 -740 0 feedthrough
rlabel pdiffusion 1018 -740 1018 -740 0 feedthrough
rlabel pdiffusion 1025 -740 1025 -740 0 feedthrough
rlabel pdiffusion 1032 -740 1032 -740 0 feedthrough
rlabel pdiffusion 1039 -740 1039 -740 0 feedthrough
rlabel pdiffusion 1046 -740 1046 -740 0 feedthrough
rlabel pdiffusion 1053 -740 1053 -740 0 feedthrough
rlabel pdiffusion 1060 -740 1060 -740 0 cellNo=690
rlabel pdiffusion 1067 -740 1067 -740 0 feedthrough
rlabel pdiffusion 1074 -740 1074 -740 0 feedthrough
rlabel pdiffusion 1081 -740 1081 -740 0 feedthrough
rlabel pdiffusion 1088 -740 1088 -740 0 feedthrough
rlabel pdiffusion 1095 -740 1095 -740 0 feedthrough
rlabel pdiffusion 1102 -740 1102 -740 0 feedthrough
rlabel pdiffusion 1109 -740 1109 -740 0 feedthrough
rlabel pdiffusion 1116 -740 1116 -740 0 feedthrough
rlabel pdiffusion 1123 -740 1123 -740 0 feedthrough
rlabel pdiffusion 1130 -740 1130 -740 0 feedthrough
rlabel pdiffusion 1137 -740 1137 -740 0 feedthrough
rlabel pdiffusion 1144 -740 1144 -740 0 feedthrough
rlabel pdiffusion 1151 -740 1151 -740 0 feedthrough
rlabel pdiffusion 1158 -740 1158 -740 0 feedthrough
rlabel pdiffusion 1165 -740 1165 -740 0 feedthrough
rlabel pdiffusion 1172 -740 1172 -740 0 feedthrough
rlabel pdiffusion 1179 -740 1179 -740 0 feedthrough
rlabel pdiffusion 1186 -740 1186 -740 0 feedthrough
rlabel pdiffusion 1193 -740 1193 -740 0 feedthrough
rlabel pdiffusion 1200 -740 1200 -740 0 feedthrough
rlabel pdiffusion 1207 -740 1207 -740 0 feedthrough
rlabel pdiffusion 1214 -740 1214 -740 0 feedthrough
rlabel pdiffusion 1221 -740 1221 -740 0 feedthrough
rlabel pdiffusion 1228 -740 1228 -740 0 feedthrough
rlabel pdiffusion 1235 -740 1235 -740 0 feedthrough
rlabel pdiffusion 1242 -740 1242 -740 0 feedthrough
rlabel pdiffusion 1249 -740 1249 -740 0 feedthrough
rlabel pdiffusion 1256 -740 1256 -740 0 feedthrough
rlabel pdiffusion 1263 -740 1263 -740 0 feedthrough
rlabel pdiffusion 1270 -740 1270 -740 0 feedthrough
rlabel pdiffusion 1277 -740 1277 -740 0 feedthrough
rlabel pdiffusion 1284 -740 1284 -740 0 feedthrough
rlabel pdiffusion 1291 -740 1291 -740 0 feedthrough
rlabel pdiffusion 1298 -740 1298 -740 0 feedthrough
rlabel pdiffusion 1305 -740 1305 -740 0 feedthrough
rlabel pdiffusion 1312 -740 1312 -740 0 feedthrough
rlabel pdiffusion 1319 -740 1319 -740 0 feedthrough
rlabel pdiffusion 1326 -740 1326 -740 0 feedthrough
rlabel pdiffusion 1333 -740 1333 -740 0 feedthrough
rlabel pdiffusion 1340 -740 1340 -740 0 feedthrough
rlabel pdiffusion 1347 -740 1347 -740 0 feedthrough
rlabel pdiffusion 1354 -740 1354 -740 0 feedthrough
rlabel pdiffusion 1361 -740 1361 -740 0 feedthrough
rlabel pdiffusion 1368 -740 1368 -740 0 feedthrough
rlabel pdiffusion 1375 -740 1375 -740 0 feedthrough
rlabel pdiffusion 1382 -740 1382 -740 0 feedthrough
rlabel pdiffusion 1389 -740 1389 -740 0 feedthrough
rlabel pdiffusion 1396 -740 1396 -740 0 feedthrough
rlabel pdiffusion 1403 -740 1403 -740 0 feedthrough
rlabel pdiffusion 1410 -740 1410 -740 0 feedthrough
rlabel pdiffusion 1417 -740 1417 -740 0 feedthrough
rlabel pdiffusion 1424 -740 1424 -740 0 cellNo=120
rlabel pdiffusion 1431 -740 1431 -740 0 feedthrough
rlabel pdiffusion 1501 -740 1501 -740 0 feedthrough
rlabel pdiffusion 1522 -740 1522 -740 0 feedthrough
rlabel pdiffusion 1571 -740 1571 -740 0 feedthrough
rlabel pdiffusion 1634 -740 1634 -740 0 feedthrough
rlabel pdiffusion 3 -879 3 -879 0 cellNo=1011
rlabel pdiffusion 10 -879 10 -879 0 cellNo=1202
rlabel pdiffusion 17 -879 17 -879 0 cellNo=1015
rlabel pdiffusion 24 -879 24 -879 0 feedthrough
rlabel pdiffusion 31 -879 31 -879 0 cellNo=628
rlabel pdiffusion 38 -879 38 -879 0 feedthrough
rlabel pdiffusion 45 -879 45 -879 0 feedthrough
rlabel pdiffusion 52 -879 52 -879 0 cellNo=911
rlabel pdiffusion 59 -879 59 -879 0 feedthrough
rlabel pdiffusion 66 -879 66 -879 0 feedthrough
rlabel pdiffusion 73 -879 73 -879 0 feedthrough
rlabel pdiffusion 80 -879 80 -879 0 feedthrough
rlabel pdiffusion 87 -879 87 -879 0 cellNo=642
rlabel pdiffusion 94 -879 94 -879 0 feedthrough
rlabel pdiffusion 101 -879 101 -879 0 cellNo=472
rlabel pdiffusion 108 -879 108 -879 0 cellNo=985
rlabel pdiffusion 115 -879 115 -879 0 feedthrough
rlabel pdiffusion 122 -879 122 -879 0 feedthrough
rlabel pdiffusion 129 -879 129 -879 0 feedthrough
rlabel pdiffusion 136 -879 136 -879 0 cellNo=421
rlabel pdiffusion 143 -879 143 -879 0 feedthrough
rlabel pdiffusion 150 -879 150 -879 0 feedthrough
rlabel pdiffusion 157 -879 157 -879 0 feedthrough
rlabel pdiffusion 164 -879 164 -879 0 cellNo=136
rlabel pdiffusion 171 -879 171 -879 0 feedthrough
rlabel pdiffusion 178 -879 178 -879 0 feedthrough
rlabel pdiffusion 185 -879 185 -879 0 feedthrough
rlabel pdiffusion 192 -879 192 -879 0 feedthrough
rlabel pdiffusion 199 -879 199 -879 0 feedthrough
rlabel pdiffusion 206 -879 206 -879 0 cellNo=275
rlabel pdiffusion 213 -879 213 -879 0 feedthrough
rlabel pdiffusion 220 -879 220 -879 0 feedthrough
rlabel pdiffusion 227 -879 227 -879 0 cellNo=70
rlabel pdiffusion 234 -879 234 -879 0 cellNo=786
rlabel pdiffusion 241 -879 241 -879 0 feedthrough
rlabel pdiffusion 248 -879 248 -879 0 cellNo=203
rlabel pdiffusion 255 -879 255 -879 0 feedthrough
rlabel pdiffusion 262 -879 262 -879 0 feedthrough
rlabel pdiffusion 269 -879 269 -879 0 feedthrough
rlabel pdiffusion 276 -879 276 -879 0 feedthrough
rlabel pdiffusion 283 -879 283 -879 0 feedthrough
rlabel pdiffusion 290 -879 290 -879 0 feedthrough
rlabel pdiffusion 297 -879 297 -879 0 cellNo=1381
rlabel pdiffusion 304 -879 304 -879 0 feedthrough
rlabel pdiffusion 311 -879 311 -879 0 feedthrough
rlabel pdiffusion 318 -879 318 -879 0 cellNo=1361
rlabel pdiffusion 325 -879 325 -879 0 feedthrough
rlabel pdiffusion 332 -879 332 -879 0 feedthrough
rlabel pdiffusion 339 -879 339 -879 0 feedthrough
rlabel pdiffusion 346 -879 346 -879 0 feedthrough
rlabel pdiffusion 353 -879 353 -879 0 feedthrough
rlabel pdiffusion 360 -879 360 -879 0 feedthrough
rlabel pdiffusion 367 -879 367 -879 0 feedthrough
rlabel pdiffusion 374 -879 374 -879 0 feedthrough
rlabel pdiffusion 381 -879 381 -879 0 feedthrough
rlabel pdiffusion 388 -879 388 -879 0 feedthrough
rlabel pdiffusion 395 -879 395 -879 0 feedthrough
rlabel pdiffusion 402 -879 402 -879 0 feedthrough
rlabel pdiffusion 409 -879 409 -879 0 feedthrough
rlabel pdiffusion 416 -879 416 -879 0 feedthrough
rlabel pdiffusion 423 -879 423 -879 0 feedthrough
rlabel pdiffusion 430 -879 430 -879 0 feedthrough
rlabel pdiffusion 437 -879 437 -879 0 feedthrough
rlabel pdiffusion 444 -879 444 -879 0 feedthrough
rlabel pdiffusion 451 -879 451 -879 0 feedthrough
rlabel pdiffusion 458 -879 458 -879 0 feedthrough
rlabel pdiffusion 465 -879 465 -879 0 cellNo=701
rlabel pdiffusion 472 -879 472 -879 0 feedthrough
rlabel pdiffusion 479 -879 479 -879 0 cellNo=199
rlabel pdiffusion 486 -879 486 -879 0 feedthrough
rlabel pdiffusion 493 -879 493 -879 0 feedthrough
rlabel pdiffusion 500 -879 500 -879 0 feedthrough
rlabel pdiffusion 507 -879 507 -879 0 feedthrough
rlabel pdiffusion 514 -879 514 -879 0 feedthrough
rlabel pdiffusion 521 -879 521 -879 0 feedthrough
rlabel pdiffusion 528 -879 528 -879 0 feedthrough
rlabel pdiffusion 535 -879 535 -879 0 feedthrough
rlabel pdiffusion 542 -879 542 -879 0 feedthrough
rlabel pdiffusion 549 -879 549 -879 0 feedthrough
rlabel pdiffusion 556 -879 556 -879 0 feedthrough
rlabel pdiffusion 563 -879 563 -879 0 cellNo=437
rlabel pdiffusion 570 -879 570 -879 0 feedthrough
rlabel pdiffusion 577 -879 577 -879 0 cellNo=345
rlabel pdiffusion 584 -879 584 -879 0 cellNo=29
rlabel pdiffusion 591 -879 591 -879 0 feedthrough
rlabel pdiffusion 598 -879 598 -879 0 feedthrough
rlabel pdiffusion 605 -879 605 -879 0 feedthrough
rlabel pdiffusion 612 -879 612 -879 0 cellNo=367
rlabel pdiffusion 619 -879 619 -879 0 feedthrough
rlabel pdiffusion 626 -879 626 -879 0 cellNo=321
rlabel pdiffusion 633 -879 633 -879 0 feedthrough
rlabel pdiffusion 640 -879 640 -879 0 cellNo=903
rlabel pdiffusion 647 -879 647 -879 0 feedthrough
rlabel pdiffusion 654 -879 654 -879 0 cellNo=1415
rlabel pdiffusion 661 -879 661 -879 0 cellNo=543
rlabel pdiffusion 668 -879 668 -879 0 feedthrough
rlabel pdiffusion 675 -879 675 -879 0 feedthrough
rlabel pdiffusion 682 -879 682 -879 0 feedthrough
rlabel pdiffusion 689 -879 689 -879 0 cellNo=418
rlabel pdiffusion 696 -879 696 -879 0 feedthrough
rlabel pdiffusion 703 -879 703 -879 0 cellNo=556
rlabel pdiffusion 710 -879 710 -879 0 feedthrough
rlabel pdiffusion 717 -879 717 -879 0 feedthrough
rlabel pdiffusion 724 -879 724 -879 0 feedthrough
rlabel pdiffusion 731 -879 731 -879 0 feedthrough
rlabel pdiffusion 738 -879 738 -879 0 cellNo=529
rlabel pdiffusion 745 -879 745 -879 0 feedthrough
rlabel pdiffusion 752 -879 752 -879 0 feedthrough
rlabel pdiffusion 759 -879 759 -879 0 cellNo=72
rlabel pdiffusion 766 -879 766 -879 0 feedthrough
rlabel pdiffusion 773 -879 773 -879 0 feedthrough
rlabel pdiffusion 780 -879 780 -879 0 cellNo=709
rlabel pdiffusion 787 -879 787 -879 0 cellNo=98
rlabel pdiffusion 794 -879 794 -879 0 cellNo=482
rlabel pdiffusion 801 -879 801 -879 0 feedthrough
rlabel pdiffusion 808 -879 808 -879 0 feedthrough
rlabel pdiffusion 815 -879 815 -879 0 feedthrough
rlabel pdiffusion 822 -879 822 -879 0 feedthrough
rlabel pdiffusion 829 -879 829 -879 0 cellNo=804
rlabel pdiffusion 836 -879 836 -879 0 feedthrough
rlabel pdiffusion 843 -879 843 -879 0 feedthrough
rlabel pdiffusion 850 -879 850 -879 0 feedthrough
rlabel pdiffusion 857 -879 857 -879 0 feedthrough
rlabel pdiffusion 864 -879 864 -879 0 feedthrough
rlabel pdiffusion 871 -879 871 -879 0 feedthrough
rlabel pdiffusion 878 -879 878 -879 0 cellNo=620
rlabel pdiffusion 885 -879 885 -879 0 feedthrough
rlabel pdiffusion 892 -879 892 -879 0 feedthrough
rlabel pdiffusion 899 -879 899 -879 0 feedthrough
rlabel pdiffusion 906 -879 906 -879 0 cellNo=759
rlabel pdiffusion 913 -879 913 -879 0 feedthrough
rlabel pdiffusion 920 -879 920 -879 0 feedthrough
rlabel pdiffusion 927 -879 927 -879 0 cellNo=96
rlabel pdiffusion 934 -879 934 -879 0 feedthrough
rlabel pdiffusion 941 -879 941 -879 0 feedthrough
rlabel pdiffusion 948 -879 948 -879 0 feedthrough
rlabel pdiffusion 955 -879 955 -879 0 feedthrough
rlabel pdiffusion 962 -879 962 -879 0 cellNo=320
rlabel pdiffusion 969 -879 969 -879 0 feedthrough
rlabel pdiffusion 976 -879 976 -879 0 feedthrough
rlabel pdiffusion 983 -879 983 -879 0 feedthrough
rlabel pdiffusion 990 -879 990 -879 0 feedthrough
rlabel pdiffusion 997 -879 997 -879 0 feedthrough
rlabel pdiffusion 1004 -879 1004 -879 0 feedthrough
rlabel pdiffusion 1011 -879 1011 -879 0 feedthrough
rlabel pdiffusion 1018 -879 1018 -879 0 feedthrough
rlabel pdiffusion 1025 -879 1025 -879 0 feedthrough
rlabel pdiffusion 1032 -879 1032 -879 0 feedthrough
rlabel pdiffusion 1039 -879 1039 -879 0 feedthrough
rlabel pdiffusion 1046 -879 1046 -879 0 feedthrough
rlabel pdiffusion 1053 -879 1053 -879 0 feedthrough
rlabel pdiffusion 1060 -879 1060 -879 0 cellNo=201
rlabel pdiffusion 1067 -879 1067 -879 0 feedthrough
rlabel pdiffusion 1074 -879 1074 -879 0 feedthrough
rlabel pdiffusion 1081 -879 1081 -879 0 feedthrough
rlabel pdiffusion 1088 -879 1088 -879 0 feedthrough
rlabel pdiffusion 1095 -879 1095 -879 0 feedthrough
rlabel pdiffusion 1102 -879 1102 -879 0 feedthrough
rlabel pdiffusion 1109 -879 1109 -879 0 feedthrough
rlabel pdiffusion 1116 -879 1116 -879 0 feedthrough
rlabel pdiffusion 1123 -879 1123 -879 0 feedthrough
rlabel pdiffusion 1130 -879 1130 -879 0 feedthrough
rlabel pdiffusion 1137 -879 1137 -879 0 feedthrough
rlabel pdiffusion 1144 -879 1144 -879 0 feedthrough
rlabel pdiffusion 1151 -879 1151 -879 0 feedthrough
rlabel pdiffusion 1158 -879 1158 -879 0 feedthrough
rlabel pdiffusion 1165 -879 1165 -879 0 feedthrough
rlabel pdiffusion 1172 -879 1172 -879 0 feedthrough
rlabel pdiffusion 1179 -879 1179 -879 0 feedthrough
rlabel pdiffusion 1186 -879 1186 -879 0 feedthrough
rlabel pdiffusion 1193 -879 1193 -879 0 feedthrough
rlabel pdiffusion 1200 -879 1200 -879 0 feedthrough
rlabel pdiffusion 1207 -879 1207 -879 0 feedthrough
rlabel pdiffusion 1214 -879 1214 -879 0 feedthrough
rlabel pdiffusion 1221 -879 1221 -879 0 feedthrough
rlabel pdiffusion 1228 -879 1228 -879 0 feedthrough
rlabel pdiffusion 1235 -879 1235 -879 0 feedthrough
rlabel pdiffusion 1242 -879 1242 -879 0 feedthrough
rlabel pdiffusion 1249 -879 1249 -879 0 feedthrough
rlabel pdiffusion 1256 -879 1256 -879 0 feedthrough
rlabel pdiffusion 1263 -879 1263 -879 0 feedthrough
rlabel pdiffusion 1270 -879 1270 -879 0 feedthrough
rlabel pdiffusion 1277 -879 1277 -879 0 feedthrough
rlabel pdiffusion 1284 -879 1284 -879 0 feedthrough
rlabel pdiffusion 1291 -879 1291 -879 0 feedthrough
rlabel pdiffusion 1298 -879 1298 -879 0 feedthrough
rlabel pdiffusion 1305 -879 1305 -879 0 feedthrough
rlabel pdiffusion 1312 -879 1312 -879 0 feedthrough
rlabel pdiffusion 1319 -879 1319 -879 0 feedthrough
rlabel pdiffusion 1326 -879 1326 -879 0 feedthrough
rlabel pdiffusion 1333 -879 1333 -879 0 feedthrough
rlabel pdiffusion 1340 -879 1340 -879 0 feedthrough
rlabel pdiffusion 1347 -879 1347 -879 0 feedthrough
rlabel pdiffusion 1354 -879 1354 -879 0 feedthrough
rlabel pdiffusion 1361 -879 1361 -879 0 feedthrough
rlabel pdiffusion 1368 -879 1368 -879 0 feedthrough
rlabel pdiffusion 1375 -879 1375 -879 0 feedthrough
rlabel pdiffusion 1382 -879 1382 -879 0 feedthrough
rlabel pdiffusion 1389 -879 1389 -879 0 feedthrough
rlabel pdiffusion 1396 -879 1396 -879 0 feedthrough
rlabel pdiffusion 1403 -879 1403 -879 0 feedthrough
rlabel pdiffusion 1410 -879 1410 -879 0 feedthrough
rlabel pdiffusion 1417 -879 1417 -879 0 feedthrough
rlabel pdiffusion 1424 -879 1424 -879 0 feedthrough
rlabel pdiffusion 1431 -879 1431 -879 0 feedthrough
rlabel pdiffusion 1438 -879 1438 -879 0 feedthrough
rlabel pdiffusion 1445 -879 1445 -879 0 feedthrough
rlabel pdiffusion 1452 -879 1452 -879 0 feedthrough
rlabel pdiffusion 1459 -879 1459 -879 0 feedthrough
rlabel pdiffusion 1466 -879 1466 -879 0 feedthrough
rlabel pdiffusion 1473 -879 1473 -879 0 feedthrough
rlabel pdiffusion 1480 -879 1480 -879 0 feedthrough
rlabel pdiffusion 1487 -879 1487 -879 0 feedthrough
rlabel pdiffusion 1494 -879 1494 -879 0 feedthrough
rlabel pdiffusion 1501 -879 1501 -879 0 feedthrough
rlabel pdiffusion 1508 -879 1508 -879 0 feedthrough
rlabel pdiffusion 1515 -879 1515 -879 0 feedthrough
rlabel pdiffusion 1522 -879 1522 -879 0 feedthrough
rlabel pdiffusion 1529 -879 1529 -879 0 feedthrough
rlabel pdiffusion 1536 -879 1536 -879 0 feedthrough
rlabel pdiffusion 1543 -879 1543 -879 0 feedthrough
rlabel pdiffusion 1550 -879 1550 -879 0 feedthrough
rlabel pdiffusion 1557 -879 1557 -879 0 feedthrough
rlabel pdiffusion 1564 -879 1564 -879 0 feedthrough
rlabel pdiffusion 1571 -879 1571 -879 0 feedthrough
rlabel pdiffusion 1578 -879 1578 -879 0 feedthrough
rlabel pdiffusion 1585 -879 1585 -879 0 feedthrough
rlabel pdiffusion 1592 -879 1592 -879 0 feedthrough
rlabel pdiffusion 1599 -879 1599 -879 0 cellNo=498
rlabel pdiffusion 1606 -879 1606 -879 0 cellNo=344
rlabel pdiffusion 1613 -879 1613 -879 0 feedthrough
rlabel pdiffusion 1620 -879 1620 -879 0 feedthrough
rlabel pdiffusion 1627 -879 1627 -879 0 feedthrough
rlabel pdiffusion 1634 -879 1634 -879 0 feedthrough
rlabel pdiffusion 1697 -879 1697 -879 0 feedthrough
rlabel pdiffusion 3 -1040 3 -1040 0 cellNo=1014
rlabel pdiffusion 10 -1040 10 -1040 0 cellNo=1413
rlabel pdiffusion 17 -1040 17 -1040 0 cellNo=1018
rlabel pdiffusion 24 -1040 24 -1040 0 cellNo=1297
rlabel pdiffusion 31 -1040 31 -1040 0 feedthrough
rlabel pdiffusion 38 -1040 38 -1040 0 feedthrough
rlabel pdiffusion 45 -1040 45 -1040 0 cellNo=357
rlabel pdiffusion 52 -1040 52 -1040 0 cellNo=375
rlabel pdiffusion 59 -1040 59 -1040 0 feedthrough
rlabel pdiffusion 66 -1040 66 -1040 0 feedthrough
rlabel pdiffusion 73 -1040 73 -1040 0 feedthrough
rlabel pdiffusion 80 -1040 80 -1040 0 feedthrough
rlabel pdiffusion 87 -1040 87 -1040 0 cellNo=687
rlabel pdiffusion 94 -1040 94 -1040 0 feedthrough
rlabel pdiffusion 101 -1040 101 -1040 0 feedthrough
rlabel pdiffusion 108 -1040 108 -1040 0 cellNo=692
rlabel pdiffusion 115 -1040 115 -1040 0 feedthrough
rlabel pdiffusion 122 -1040 122 -1040 0 cellNo=91
rlabel pdiffusion 129 -1040 129 -1040 0 feedthrough
rlabel pdiffusion 136 -1040 136 -1040 0 feedthrough
rlabel pdiffusion 143 -1040 143 -1040 0 feedthrough
rlabel pdiffusion 150 -1040 150 -1040 0 feedthrough
rlabel pdiffusion 157 -1040 157 -1040 0 feedthrough
rlabel pdiffusion 164 -1040 164 -1040 0 feedthrough
rlabel pdiffusion 171 -1040 171 -1040 0 feedthrough
rlabel pdiffusion 178 -1040 178 -1040 0 feedthrough
rlabel pdiffusion 185 -1040 185 -1040 0 feedthrough
rlabel pdiffusion 192 -1040 192 -1040 0 feedthrough
rlabel pdiffusion 199 -1040 199 -1040 0 cellNo=658
rlabel pdiffusion 206 -1040 206 -1040 0 feedthrough
rlabel pdiffusion 213 -1040 213 -1040 0 feedthrough
rlabel pdiffusion 220 -1040 220 -1040 0 cellNo=1414
rlabel pdiffusion 227 -1040 227 -1040 0 feedthrough
rlabel pdiffusion 234 -1040 234 -1040 0 feedthrough
rlabel pdiffusion 241 -1040 241 -1040 0 feedthrough
rlabel pdiffusion 248 -1040 248 -1040 0 feedthrough
rlabel pdiffusion 255 -1040 255 -1040 0 feedthrough
rlabel pdiffusion 262 -1040 262 -1040 0 feedthrough
rlabel pdiffusion 269 -1040 269 -1040 0 feedthrough
rlabel pdiffusion 276 -1040 276 -1040 0 feedthrough
rlabel pdiffusion 283 -1040 283 -1040 0 feedthrough
rlabel pdiffusion 290 -1040 290 -1040 0 cellNo=443
rlabel pdiffusion 297 -1040 297 -1040 0 feedthrough
rlabel pdiffusion 304 -1040 304 -1040 0 feedthrough
rlabel pdiffusion 311 -1040 311 -1040 0 cellNo=893
rlabel pdiffusion 318 -1040 318 -1040 0 feedthrough
rlabel pdiffusion 325 -1040 325 -1040 0 feedthrough
rlabel pdiffusion 332 -1040 332 -1040 0 feedthrough
rlabel pdiffusion 339 -1040 339 -1040 0 feedthrough
rlabel pdiffusion 346 -1040 346 -1040 0 feedthrough
rlabel pdiffusion 353 -1040 353 -1040 0 feedthrough
rlabel pdiffusion 360 -1040 360 -1040 0 feedthrough
rlabel pdiffusion 367 -1040 367 -1040 0 feedthrough
rlabel pdiffusion 374 -1040 374 -1040 0 feedthrough
rlabel pdiffusion 381 -1040 381 -1040 0 feedthrough
rlabel pdiffusion 388 -1040 388 -1040 0 feedthrough
rlabel pdiffusion 395 -1040 395 -1040 0 feedthrough
rlabel pdiffusion 402 -1040 402 -1040 0 feedthrough
rlabel pdiffusion 409 -1040 409 -1040 0 feedthrough
rlabel pdiffusion 416 -1040 416 -1040 0 feedthrough
rlabel pdiffusion 423 -1040 423 -1040 0 feedthrough
rlabel pdiffusion 430 -1040 430 -1040 0 feedthrough
rlabel pdiffusion 437 -1040 437 -1040 0 feedthrough
rlabel pdiffusion 444 -1040 444 -1040 0 feedthrough
rlabel pdiffusion 451 -1040 451 -1040 0 feedthrough
rlabel pdiffusion 458 -1040 458 -1040 0 feedthrough
rlabel pdiffusion 465 -1040 465 -1040 0 cellNo=523
rlabel pdiffusion 472 -1040 472 -1040 0 cellNo=877
rlabel pdiffusion 479 -1040 479 -1040 0 feedthrough
rlabel pdiffusion 486 -1040 486 -1040 0 feedthrough
rlabel pdiffusion 493 -1040 493 -1040 0 feedthrough
rlabel pdiffusion 500 -1040 500 -1040 0 feedthrough
rlabel pdiffusion 507 -1040 507 -1040 0 feedthrough
rlabel pdiffusion 514 -1040 514 -1040 0 feedthrough
rlabel pdiffusion 521 -1040 521 -1040 0 feedthrough
rlabel pdiffusion 528 -1040 528 -1040 0 feedthrough
rlabel pdiffusion 535 -1040 535 -1040 0 cellNo=310
rlabel pdiffusion 542 -1040 542 -1040 0 feedthrough
rlabel pdiffusion 549 -1040 549 -1040 0 cellNo=331
rlabel pdiffusion 556 -1040 556 -1040 0 feedthrough
rlabel pdiffusion 563 -1040 563 -1040 0 feedthrough
rlabel pdiffusion 570 -1040 570 -1040 0 feedthrough
rlabel pdiffusion 577 -1040 577 -1040 0 feedthrough
rlabel pdiffusion 584 -1040 584 -1040 0 feedthrough
rlabel pdiffusion 591 -1040 591 -1040 0 cellNo=381
rlabel pdiffusion 598 -1040 598 -1040 0 cellNo=346
rlabel pdiffusion 605 -1040 605 -1040 0 cellNo=679
rlabel pdiffusion 612 -1040 612 -1040 0 feedthrough
rlabel pdiffusion 619 -1040 619 -1040 0 cellNo=353
rlabel pdiffusion 626 -1040 626 -1040 0 cellNo=473
rlabel pdiffusion 633 -1040 633 -1040 0 cellNo=907
rlabel pdiffusion 640 -1040 640 -1040 0 feedthrough
rlabel pdiffusion 647 -1040 647 -1040 0 feedthrough
rlabel pdiffusion 654 -1040 654 -1040 0 feedthrough
rlabel pdiffusion 661 -1040 661 -1040 0 feedthrough
rlabel pdiffusion 668 -1040 668 -1040 0 feedthrough
rlabel pdiffusion 675 -1040 675 -1040 0 feedthrough
rlabel pdiffusion 682 -1040 682 -1040 0 cellNo=900
rlabel pdiffusion 689 -1040 689 -1040 0 feedthrough
rlabel pdiffusion 696 -1040 696 -1040 0 feedthrough
rlabel pdiffusion 703 -1040 703 -1040 0 feedthrough
rlabel pdiffusion 710 -1040 710 -1040 0 feedthrough
rlabel pdiffusion 717 -1040 717 -1040 0 feedthrough
rlabel pdiffusion 724 -1040 724 -1040 0 cellNo=365
rlabel pdiffusion 731 -1040 731 -1040 0 cellNo=652
rlabel pdiffusion 738 -1040 738 -1040 0 feedthrough
rlabel pdiffusion 745 -1040 745 -1040 0 feedthrough
rlabel pdiffusion 752 -1040 752 -1040 0 feedthrough
rlabel pdiffusion 759 -1040 759 -1040 0 cellNo=778
rlabel pdiffusion 766 -1040 766 -1040 0 cellNo=259
rlabel pdiffusion 773 -1040 773 -1040 0 feedthrough
rlabel pdiffusion 780 -1040 780 -1040 0 feedthrough
rlabel pdiffusion 787 -1040 787 -1040 0 feedthrough
rlabel pdiffusion 794 -1040 794 -1040 0 cellNo=813
rlabel pdiffusion 801 -1040 801 -1040 0 feedthrough
rlabel pdiffusion 808 -1040 808 -1040 0 cellNo=326
rlabel pdiffusion 815 -1040 815 -1040 0 feedthrough
rlabel pdiffusion 822 -1040 822 -1040 0 feedthrough
rlabel pdiffusion 829 -1040 829 -1040 0 cellNo=545
rlabel pdiffusion 836 -1040 836 -1040 0 feedthrough
rlabel pdiffusion 843 -1040 843 -1040 0 cellNo=105
rlabel pdiffusion 850 -1040 850 -1040 0 feedthrough
rlabel pdiffusion 857 -1040 857 -1040 0 cellNo=196
rlabel pdiffusion 864 -1040 864 -1040 0 feedthrough
rlabel pdiffusion 871 -1040 871 -1040 0 cellNo=316
rlabel pdiffusion 878 -1040 878 -1040 0 cellNo=933
rlabel pdiffusion 885 -1040 885 -1040 0 feedthrough
rlabel pdiffusion 892 -1040 892 -1040 0 feedthrough
rlabel pdiffusion 899 -1040 899 -1040 0 cellNo=339
rlabel pdiffusion 906 -1040 906 -1040 0 feedthrough
rlabel pdiffusion 913 -1040 913 -1040 0 feedthrough
rlabel pdiffusion 920 -1040 920 -1040 0 feedthrough
rlabel pdiffusion 927 -1040 927 -1040 0 feedthrough
rlabel pdiffusion 934 -1040 934 -1040 0 feedthrough
rlabel pdiffusion 941 -1040 941 -1040 0 feedthrough
rlabel pdiffusion 948 -1040 948 -1040 0 feedthrough
rlabel pdiffusion 955 -1040 955 -1040 0 cellNo=265
rlabel pdiffusion 962 -1040 962 -1040 0 feedthrough
rlabel pdiffusion 969 -1040 969 -1040 0 feedthrough
rlabel pdiffusion 976 -1040 976 -1040 0 cellNo=516
rlabel pdiffusion 983 -1040 983 -1040 0 feedthrough
rlabel pdiffusion 990 -1040 990 -1040 0 cellNo=867
rlabel pdiffusion 997 -1040 997 -1040 0 feedthrough
rlabel pdiffusion 1004 -1040 1004 -1040 0 feedthrough
rlabel pdiffusion 1011 -1040 1011 -1040 0 feedthrough
rlabel pdiffusion 1018 -1040 1018 -1040 0 feedthrough
rlabel pdiffusion 1025 -1040 1025 -1040 0 feedthrough
rlabel pdiffusion 1032 -1040 1032 -1040 0 feedthrough
rlabel pdiffusion 1039 -1040 1039 -1040 0 feedthrough
rlabel pdiffusion 1046 -1040 1046 -1040 0 feedthrough
rlabel pdiffusion 1053 -1040 1053 -1040 0 feedthrough
rlabel pdiffusion 1060 -1040 1060 -1040 0 cellNo=938
rlabel pdiffusion 1067 -1040 1067 -1040 0 cellNo=88
rlabel pdiffusion 1074 -1040 1074 -1040 0 feedthrough
rlabel pdiffusion 1081 -1040 1081 -1040 0 feedthrough
rlabel pdiffusion 1088 -1040 1088 -1040 0 feedthrough
rlabel pdiffusion 1095 -1040 1095 -1040 0 feedthrough
rlabel pdiffusion 1102 -1040 1102 -1040 0 feedthrough
rlabel pdiffusion 1109 -1040 1109 -1040 0 feedthrough
rlabel pdiffusion 1116 -1040 1116 -1040 0 feedthrough
rlabel pdiffusion 1123 -1040 1123 -1040 0 feedthrough
rlabel pdiffusion 1130 -1040 1130 -1040 0 feedthrough
rlabel pdiffusion 1137 -1040 1137 -1040 0 feedthrough
rlabel pdiffusion 1144 -1040 1144 -1040 0 feedthrough
rlabel pdiffusion 1151 -1040 1151 -1040 0 feedthrough
rlabel pdiffusion 1158 -1040 1158 -1040 0 feedthrough
rlabel pdiffusion 1165 -1040 1165 -1040 0 feedthrough
rlabel pdiffusion 1172 -1040 1172 -1040 0 feedthrough
rlabel pdiffusion 1179 -1040 1179 -1040 0 feedthrough
rlabel pdiffusion 1186 -1040 1186 -1040 0 feedthrough
rlabel pdiffusion 1193 -1040 1193 -1040 0 feedthrough
rlabel pdiffusion 1200 -1040 1200 -1040 0 feedthrough
rlabel pdiffusion 1207 -1040 1207 -1040 0 feedthrough
rlabel pdiffusion 1214 -1040 1214 -1040 0 feedthrough
rlabel pdiffusion 1221 -1040 1221 -1040 0 feedthrough
rlabel pdiffusion 1228 -1040 1228 -1040 0 feedthrough
rlabel pdiffusion 1235 -1040 1235 -1040 0 feedthrough
rlabel pdiffusion 1242 -1040 1242 -1040 0 feedthrough
rlabel pdiffusion 1249 -1040 1249 -1040 0 feedthrough
rlabel pdiffusion 1256 -1040 1256 -1040 0 feedthrough
rlabel pdiffusion 1263 -1040 1263 -1040 0 feedthrough
rlabel pdiffusion 1270 -1040 1270 -1040 0 feedthrough
rlabel pdiffusion 1277 -1040 1277 -1040 0 feedthrough
rlabel pdiffusion 1284 -1040 1284 -1040 0 feedthrough
rlabel pdiffusion 1291 -1040 1291 -1040 0 feedthrough
rlabel pdiffusion 1298 -1040 1298 -1040 0 feedthrough
rlabel pdiffusion 1305 -1040 1305 -1040 0 feedthrough
rlabel pdiffusion 1312 -1040 1312 -1040 0 feedthrough
rlabel pdiffusion 1319 -1040 1319 -1040 0 feedthrough
rlabel pdiffusion 1326 -1040 1326 -1040 0 feedthrough
rlabel pdiffusion 1333 -1040 1333 -1040 0 feedthrough
rlabel pdiffusion 1340 -1040 1340 -1040 0 feedthrough
rlabel pdiffusion 1347 -1040 1347 -1040 0 feedthrough
rlabel pdiffusion 1354 -1040 1354 -1040 0 feedthrough
rlabel pdiffusion 1361 -1040 1361 -1040 0 feedthrough
rlabel pdiffusion 1368 -1040 1368 -1040 0 feedthrough
rlabel pdiffusion 1375 -1040 1375 -1040 0 feedthrough
rlabel pdiffusion 1382 -1040 1382 -1040 0 feedthrough
rlabel pdiffusion 1389 -1040 1389 -1040 0 feedthrough
rlabel pdiffusion 1396 -1040 1396 -1040 0 feedthrough
rlabel pdiffusion 1403 -1040 1403 -1040 0 feedthrough
rlabel pdiffusion 1410 -1040 1410 -1040 0 feedthrough
rlabel pdiffusion 1417 -1040 1417 -1040 0 feedthrough
rlabel pdiffusion 1424 -1040 1424 -1040 0 feedthrough
rlabel pdiffusion 1431 -1040 1431 -1040 0 feedthrough
rlabel pdiffusion 1438 -1040 1438 -1040 0 feedthrough
rlabel pdiffusion 1445 -1040 1445 -1040 0 feedthrough
rlabel pdiffusion 1452 -1040 1452 -1040 0 feedthrough
rlabel pdiffusion 1459 -1040 1459 -1040 0 feedthrough
rlabel pdiffusion 1466 -1040 1466 -1040 0 feedthrough
rlabel pdiffusion 1473 -1040 1473 -1040 0 feedthrough
rlabel pdiffusion 1480 -1040 1480 -1040 0 feedthrough
rlabel pdiffusion 1487 -1040 1487 -1040 0 feedthrough
rlabel pdiffusion 1494 -1040 1494 -1040 0 feedthrough
rlabel pdiffusion 1501 -1040 1501 -1040 0 feedthrough
rlabel pdiffusion 1508 -1040 1508 -1040 0 feedthrough
rlabel pdiffusion 1515 -1040 1515 -1040 0 feedthrough
rlabel pdiffusion 1522 -1040 1522 -1040 0 feedthrough
rlabel pdiffusion 1529 -1040 1529 -1040 0 feedthrough
rlabel pdiffusion 1536 -1040 1536 -1040 0 feedthrough
rlabel pdiffusion 1543 -1040 1543 -1040 0 feedthrough
rlabel pdiffusion 1550 -1040 1550 -1040 0 feedthrough
rlabel pdiffusion 1557 -1040 1557 -1040 0 feedthrough
rlabel pdiffusion 1564 -1040 1564 -1040 0 feedthrough
rlabel pdiffusion 1571 -1040 1571 -1040 0 feedthrough
rlabel pdiffusion 1578 -1040 1578 -1040 0 feedthrough
rlabel pdiffusion 1585 -1040 1585 -1040 0 feedthrough
rlabel pdiffusion 1592 -1040 1592 -1040 0 feedthrough
rlabel pdiffusion 1599 -1040 1599 -1040 0 feedthrough
rlabel pdiffusion 1606 -1040 1606 -1040 0 feedthrough
rlabel pdiffusion 1613 -1040 1613 -1040 0 feedthrough
rlabel pdiffusion 1620 -1040 1620 -1040 0 feedthrough
rlabel pdiffusion 1627 -1040 1627 -1040 0 feedthrough
rlabel pdiffusion 1634 -1040 1634 -1040 0 feedthrough
rlabel pdiffusion 1641 -1040 1641 -1040 0 feedthrough
rlabel pdiffusion 1648 -1040 1648 -1040 0 feedthrough
rlabel pdiffusion 1655 -1040 1655 -1040 0 feedthrough
rlabel pdiffusion 1662 -1040 1662 -1040 0 feedthrough
rlabel pdiffusion 1669 -1040 1669 -1040 0 feedthrough
rlabel pdiffusion 1676 -1040 1676 -1040 0 feedthrough
rlabel pdiffusion 1683 -1040 1683 -1040 0 feedthrough
rlabel pdiffusion 1690 -1040 1690 -1040 0 feedthrough
rlabel pdiffusion 1697 -1040 1697 -1040 0 feedthrough
rlabel pdiffusion 1704 -1040 1704 -1040 0 feedthrough
rlabel pdiffusion 1711 -1040 1711 -1040 0 feedthrough
rlabel pdiffusion 1718 -1040 1718 -1040 0 feedthrough
rlabel pdiffusion 1725 -1040 1725 -1040 0 feedthrough
rlabel pdiffusion 3 -1191 3 -1191 0 cellNo=1017
rlabel pdiffusion 10 -1191 10 -1191 0 cellNo=1328
rlabel pdiffusion 17 -1191 17 -1191 0 cellNo=1019
rlabel pdiffusion 24 -1191 24 -1191 0 cellNo=1020
rlabel pdiffusion 31 -1191 31 -1191 0 feedthrough
rlabel pdiffusion 38 -1191 38 -1191 0 feedthrough
rlabel pdiffusion 45 -1191 45 -1191 0 feedthrough
rlabel pdiffusion 52 -1191 52 -1191 0 feedthrough
rlabel pdiffusion 59 -1191 59 -1191 0 feedthrough
rlabel pdiffusion 66 -1191 66 -1191 0 feedthrough
rlabel pdiffusion 73 -1191 73 -1191 0 cellNo=548
rlabel pdiffusion 80 -1191 80 -1191 0 cellNo=129
rlabel pdiffusion 87 -1191 87 -1191 0 cellNo=181
rlabel pdiffusion 94 -1191 94 -1191 0 feedthrough
rlabel pdiffusion 101 -1191 101 -1191 0 cellNo=906
rlabel pdiffusion 108 -1191 108 -1191 0 feedthrough
rlabel pdiffusion 115 -1191 115 -1191 0 feedthrough
rlabel pdiffusion 122 -1191 122 -1191 0 cellNo=972
rlabel pdiffusion 129 -1191 129 -1191 0 feedthrough
rlabel pdiffusion 136 -1191 136 -1191 0 feedthrough
rlabel pdiffusion 143 -1191 143 -1191 0 feedthrough
rlabel pdiffusion 150 -1191 150 -1191 0 cellNo=432
rlabel pdiffusion 157 -1191 157 -1191 0 feedthrough
rlabel pdiffusion 164 -1191 164 -1191 0 cellNo=206
rlabel pdiffusion 171 -1191 171 -1191 0 feedthrough
rlabel pdiffusion 178 -1191 178 -1191 0 feedthrough
rlabel pdiffusion 185 -1191 185 -1191 0 cellNo=271
rlabel pdiffusion 192 -1191 192 -1191 0 feedthrough
rlabel pdiffusion 199 -1191 199 -1191 0 cellNo=243
rlabel pdiffusion 206 -1191 206 -1191 0 cellNo=33
rlabel pdiffusion 213 -1191 213 -1191 0 feedthrough
rlabel pdiffusion 220 -1191 220 -1191 0 feedthrough
rlabel pdiffusion 227 -1191 227 -1191 0 feedthrough
rlabel pdiffusion 234 -1191 234 -1191 0 cellNo=411
rlabel pdiffusion 241 -1191 241 -1191 0 feedthrough
rlabel pdiffusion 248 -1191 248 -1191 0 feedthrough
rlabel pdiffusion 255 -1191 255 -1191 0 cellNo=27
rlabel pdiffusion 262 -1191 262 -1191 0 feedthrough
rlabel pdiffusion 269 -1191 269 -1191 0 feedthrough
rlabel pdiffusion 276 -1191 276 -1191 0 cellNo=836
rlabel pdiffusion 283 -1191 283 -1191 0 feedthrough
rlabel pdiffusion 290 -1191 290 -1191 0 feedthrough
rlabel pdiffusion 297 -1191 297 -1191 0 feedthrough
rlabel pdiffusion 304 -1191 304 -1191 0 feedthrough
rlabel pdiffusion 311 -1191 311 -1191 0 feedthrough
rlabel pdiffusion 318 -1191 318 -1191 0 feedthrough
rlabel pdiffusion 325 -1191 325 -1191 0 feedthrough
rlabel pdiffusion 332 -1191 332 -1191 0 feedthrough
rlabel pdiffusion 339 -1191 339 -1191 0 feedthrough
rlabel pdiffusion 346 -1191 346 -1191 0 feedthrough
rlabel pdiffusion 353 -1191 353 -1191 0 feedthrough
rlabel pdiffusion 360 -1191 360 -1191 0 feedthrough
rlabel pdiffusion 367 -1191 367 -1191 0 feedthrough
rlabel pdiffusion 374 -1191 374 -1191 0 feedthrough
rlabel pdiffusion 381 -1191 381 -1191 0 feedthrough
rlabel pdiffusion 388 -1191 388 -1191 0 feedthrough
rlabel pdiffusion 395 -1191 395 -1191 0 feedthrough
rlabel pdiffusion 402 -1191 402 -1191 0 feedthrough
rlabel pdiffusion 409 -1191 409 -1191 0 feedthrough
rlabel pdiffusion 416 -1191 416 -1191 0 feedthrough
rlabel pdiffusion 423 -1191 423 -1191 0 feedthrough
rlabel pdiffusion 430 -1191 430 -1191 0 feedthrough
rlabel pdiffusion 437 -1191 437 -1191 0 feedthrough
rlabel pdiffusion 444 -1191 444 -1191 0 feedthrough
rlabel pdiffusion 451 -1191 451 -1191 0 feedthrough
rlabel pdiffusion 458 -1191 458 -1191 0 feedthrough
rlabel pdiffusion 465 -1191 465 -1191 0 cellNo=655
rlabel pdiffusion 472 -1191 472 -1191 0 feedthrough
rlabel pdiffusion 479 -1191 479 -1191 0 feedthrough
rlabel pdiffusion 486 -1191 486 -1191 0 cellNo=940
rlabel pdiffusion 493 -1191 493 -1191 0 feedthrough
rlabel pdiffusion 500 -1191 500 -1191 0 feedthrough
rlabel pdiffusion 507 -1191 507 -1191 0 cellNo=665
rlabel pdiffusion 514 -1191 514 -1191 0 cellNo=343
rlabel pdiffusion 521 -1191 521 -1191 0 feedthrough
rlabel pdiffusion 528 -1191 528 -1191 0 feedthrough
rlabel pdiffusion 535 -1191 535 -1191 0 feedthrough
rlabel pdiffusion 542 -1191 542 -1191 0 cellNo=766
rlabel pdiffusion 549 -1191 549 -1191 0 feedthrough
rlabel pdiffusion 556 -1191 556 -1191 0 feedthrough
rlabel pdiffusion 563 -1191 563 -1191 0 feedthrough
rlabel pdiffusion 570 -1191 570 -1191 0 feedthrough
rlabel pdiffusion 577 -1191 577 -1191 0 cellNo=487
rlabel pdiffusion 584 -1191 584 -1191 0 feedthrough
rlabel pdiffusion 591 -1191 591 -1191 0 feedthrough
rlabel pdiffusion 598 -1191 598 -1191 0 cellNo=410
rlabel pdiffusion 605 -1191 605 -1191 0 feedthrough
rlabel pdiffusion 612 -1191 612 -1191 0 cellNo=263
rlabel pdiffusion 619 -1191 619 -1191 0 cellNo=714
rlabel pdiffusion 626 -1191 626 -1191 0 feedthrough
rlabel pdiffusion 633 -1191 633 -1191 0 feedthrough
rlabel pdiffusion 640 -1191 640 -1191 0 feedthrough
rlabel pdiffusion 647 -1191 647 -1191 0 feedthrough
rlabel pdiffusion 654 -1191 654 -1191 0 feedthrough
rlabel pdiffusion 661 -1191 661 -1191 0 cellNo=668
rlabel pdiffusion 668 -1191 668 -1191 0 feedthrough
rlabel pdiffusion 675 -1191 675 -1191 0 feedthrough
rlabel pdiffusion 682 -1191 682 -1191 0 feedthrough
rlabel pdiffusion 689 -1191 689 -1191 0 feedthrough
rlabel pdiffusion 696 -1191 696 -1191 0 feedthrough
rlabel pdiffusion 703 -1191 703 -1191 0 feedthrough
rlabel pdiffusion 710 -1191 710 -1191 0 feedthrough
rlabel pdiffusion 717 -1191 717 -1191 0 cellNo=618
rlabel pdiffusion 724 -1191 724 -1191 0 cellNo=852
rlabel pdiffusion 731 -1191 731 -1191 0 feedthrough
rlabel pdiffusion 738 -1191 738 -1191 0 feedthrough
rlabel pdiffusion 745 -1191 745 -1191 0 cellNo=794
rlabel pdiffusion 752 -1191 752 -1191 0 cellNo=53
rlabel pdiffusion 759 -1191 759 -1191 0 feedthrough
rlabel pdiffusion 766 -1191 766 -1191 0 feedthrough
rlabel pdiffusion 773 -1191 773 -1191 0 feedthrough
rlabel pdiffusion 780 -1191 780 -1191 0 feedthrough
rlabel pdiffusion 787 -1191 787 -1191 0 feedthrough
rlabel pdiffusion 794 -1191 794 -1191 0 feedthrough
rlabel pdiffusion 801 -1191 801 -1191 0 feedthrough
rlabel pdiffusion 808 -1191 808 -1191 0 feedthrough
rlabel pdiffusion 815 -1191 815 -1191 0 feedthrough
rlabel pdiffusion 822 -1191 822 -1191 0 feedthrough
rlabel pdiffusion 829 -1191 829 -1191 0 cellNo=155
rlabel pdiffusion 836 -1191 836 -1191 0 feedthrough
rlabel pdiffusion 843 -1191 843 -1191 0 feedthrough
rlabel pdiffusion 850 -1191 850 -1191 0 feedthrough
rlabel pdiffusion 857 -1191 857 -1191 0 feedthrough
rlabel pdiffusion 864 -1191 864 -1191 0 feedthrough
rlabel pdiffusion 871 -1191 871 -1191 0 cellNo=348
rlabel pdiffusion 878 -1191 878 -1191 0 feedthrough
rlabel pdiffusion 885 -1191 885 -1191 0 feedthrough
rlabel pdiffusion 892 -1191 892 -1191 0 cellNo=539
rlabel pdiffusion 899 -1191 899 -1191 0 cellNo=595
rlabel pdiffusion 906 -1191 906 -1191 0 feedthrough
rlabel pdiffusion 913 -1191 913 -1191 0 feedthrough
rlabel pdiffusion 920 -1191 920 -1191 0 feedthrough
rlabel pdiffusion 927 -1191 927 -1191 0 feedthrough
rlabel pdiffusion 934 -1191 934 -1191 0 feedthrough
rlabel pdiffusion 941 -1191 941 -1191 0 feedthrough
rlabel pdiffusion 948 -1191 948 -1191 0 feedthrough
rlabel pdiffusion 955 -1191 955 -1191 0 cellNo=890
rlabel pdiffusion 962 -1191 962 -1191 0 feedthrough
rlabel pdiffusion 969 -1191 969 -1191 0 cellNo=536
rlabel pdiffusion 976 -1191 976 -1191 0 feedthrough
rlabel pdiffusion 983 -1191 983 -1191 0 feedthrough
rlabel pdiffusion 990 -1191 990 -1191 0 cellNo=768
rlabel pdiffusion 997 -1191 997 -1191 0 feedthrough
rlabel pdiffusion 1004 -1191 1004 -1191 0 feedthrough
rlabel pdiffusion 1011 -1191 1011 -1191 0 feedthrough
rlabel pdiffusion 1018 -1191 1018 -1191 0 feedthrough
rlabel pdiffusion 1025 -1191 1025 -1191 0 feedthrough
rlabel pdiffusion 1032 -1191 1032 -1191 0 feedthrough
rlabel pdiffusion 1039 -1191 1039 -1191 0 feedthrough
rlabel pdiffusion 1046 -1191 1046 -1191 0 cellNo=164
rlabel pdiffusion 1053 -1191 1053 -1191 0 feedthrough
rlabel pdiffusion 1060 -1191 1060 -1191 0 feedthrough
rlabel pdiffusion 1067 -1191 1067 -1191 0 feedthrough
rlabel pdiffusion 1074 -1191 1074 -1191 0 feedthrough
rlabel pdiffusion 1081 -1191 1081 -1191 0 feedthrough
rlabel pdiffusion 1088 -1191 1088 -1191 0 feedthrough
rlabel pdiffusion 1095 -1191 1095 -1191 0 feedthrough
rlabel pdiffusion 1102 -1191 1102 -1191 0 feedthrough
rlabel pdiffusion 1109 -1191 1109 -1191 0 feedthrough
rlabel pdiffusion 1116 -1191 1116 -1191 0 feedthrough
rlabel pdiffusion 1123 -1191 1123 -1191 0 feedthrough
rlabel pdiffusion 1130 -1191 1130 -1191 0 feedthrough
rlabel pdiffusion 1137 -1191 1137 -1191 0 feedthrough
rlabel pdiffusion 1144 -1191 1144 -1191 0 feedthrough
rlabel pdiffusion 1151 -1191 1151 -1191 0 feedthrough
rlabel pdiffusion 1158 -1191 1158 -1191 0 feedthrough
rlabel pdiffusion 1165 -1191 1165 -1191 0 feedthrough
rlabel pdiffusion 1172 -1191 1172 -1191 0 feedthrough
rlabel pdiffusion 1179 -1191 1179 -1191 0 feedthrough
rlabel pdiffusion 1186 -1191 1186 -1191 0 feedthrough
rlabel pdiffusion 1193 -1191 1193 -1191 0 feedthrough
rlabel pdiffusion 1200 -1191 1200 -1191 0 feedthrough
rlabel pdiffusion 1207 -1191 1207 -1191 0 feedthrough
rlabel pdiffusion 1214 -1191 1214 -1191 0 feedthrough
rlabel pdiffusion 1221 -1191 1221 -1191 0 feedthrough
rlabel pdiffusion 1228 -1191 1228 -1191 0 feedthrough
rlabel pdiffusion 1235 -1191 1235 -1191 0 feedthrough
rlabel pdiffusion 1242 -1191 1242 -1191 0 feedthrough
rlabel pdiffusion 1249 -1191 1249 -1191 0 feedthrough
rlabel pdiffusion 1256 -1191 1256 -1191 0 feedthrough
rlabel pdiffusion 1263 -1191 1263 -1191 0 feedthrough
rlabel pdiffusion 1270 -1191 1270 -1191 0 feedthrough
rlabel pdiffusion 1277 -1191 1277 -1191 0 feedthrough
rlabel pdiffusion 1284 -1191 1284 -1191 0 feedthrough
rlabel pdiffusion 1291 -1191 1291 -1191 0 feedthrough
rlabel pdiffusion 1298 -1191 1298 -1191 0 feedthrough
rlabel pdiffusion 1305 -1191 1305 -1191 0 feedthrough
rlabel pdiffusion 1312 -1191 1312 -1191 0 feedthrough
rlabel pdiffusion 1319 -1191 1319 -1191 0 feedthrough
rlabel pdiffusion 1326 -1191 1326 -1191 0 feedthrough
rlabel pdiffusion 1333 -1191 1333 -1191 0 feedthrough
rlabel pdiffusion 1340 -1191 1340 -1191 0 feedthrough
rlabel pdiffusion 1347 -1191 1347 -1191 0 feedthrough
rlabel pdiffusion 1354 -1191 1354 -1191 0 feedthrough
rlabel pdiffusion 1361 -1191 1361 -1191 0 feedthrough
rlabel pdiffusion 1368 -1191 1368 -1191 0 feedthrough
rlabel pdiffusion 1375 -1191 1375 -1191 0 feedthrough
rlabel pdiffusion 1382 -1191 1382 -1191 0 feedthrough
rlabel pdiffusion 1389 -1191 1389 -1191 0 feedthrough
rlabel pdiffusion 1396 -1191 1396 -1191 0 feedthrough
rlabel pdiffusion 1403 -1191 1403 -1191 0 feedthrough
rlabel pdiffusion 1410 -1191 1410 -1191 0 feedthrough
rlabel pdiffusion 1417 -1191 1417 -1191 0 feedthrough
rlabel pdiffusion 1424 -1191 1424 -1191 0 feedthrough
rlabel pdiffusion 1431 -1191 1431 -1191 0 feedthrough
rlabel pdiffusion 1438 -1191 1438 -1191 0 feedthrough
rlabel pdiffusion 1445 -1191 1445 -1191 0 feedthrough
rlabel pdiffusion 1452 -1191 1452 -1191 0 feedthrough
rlabel pdiffusion 1459 -1191 1459 -1191 0 feedthrough
rlabel pdiffusion 1466 -1191 1466 -1191 0 feedthrough
rlabel pdiffusion 1473 -1191 1473 -1191 0 feedthrough
rlabel pdiffusion 1480 -1191 1480 -1191 0 feedthrough
rlabel pdiffusion 1487 -1191 1487 -1191 0 feedthrough
rlabel pdiffusion 1494 -1191 1494 -1191 0 feedthrough
rlabel pdiffusion 1501 -1191 1501 -1191 0 feedthrough
rlabel pdiffusion 1508 -1191 1508 -1191 0 feedthrough
rlabel pdiffusion 1515 -1191 1515 -1191 0 feedthrough
rlabel pdiffusion 1522 -1191 1522 -1191 0 feedthrough
rlabel pdiffusion 1529 -1191 1529 -1191 0 feedthrough
rlabel pdiffusion 1536 -1191 1536 -1191 0 feedthrough
rlabel pdiffusion 1543 -1191 1543 -1191 0 feedthrough
rlabel pdiffusion 1550 -1191 1550 -1191 0 feedthrough
rlabel pdiffusion 1557 -1191 1557 -1191 0 feedthrough
rlabel pdiffusion 1564 -1191 1564 -1191 0 feedthrough
rlabel pdiffusion 1571 -1191 1571 -1191 0 feedthrough
rlabel pdiffusion 1578 -1191 1578 -1191 0 feedthrough
rlabel pdiffusion 1585 -1191 1585 -1191 0 feedthrough
rlabel pdiffusion 1592 -1191 1592 -1191 0 feedthrough
rlabel pdiffusion 1599 -1191 1599 -1191 0 feedthrough
rlabel pdiffusion 1606 -1191 1606 -1191 0 feedthrough
rlabel pdiffusion 1613 -1191 1613 -1191 0 feedthrough
rlabel pdiffusion 1620 -1191 1620 -1191 0 feedthrough
rlabel pdiffusion 1627 -1191 1627 -1191 0 feedthrough
rlabel pdiffusion 1634 -1191 1634 -1191 0 feedthrough
rlabel pdiffusion 1641 -1191 1641 -1191 0 feedthrough
rlabel pdiffusion 1648 -1191 1648 -1191 0 cellNo=400
rlabel pdiffusion 1655 -1191 1655 -1191 0 feedthrough
rlabel pdiffusion 1662 -1191 1662 -1191 0 cellNo=336
rlabel pdiffusion 1676 -1191 1676 -1191 0 feedthrough
rlabel pdiffusion 1725 -1191 1725 -1191 0 feedthrough
rlabel pdiffusion 1732 -1191 1732 -1191 0 feedthrough
rlabel pdiffusion 3 -1322 3 -1322 0 cellNo=1016
rlabel pdiffusion 10 -1322 10 -1322 0 cellNo=1238
rlabel pdiffusion 17 -1322 17 -1322 0 cellNo=1340
rlabel pdiffusion 24 -1322 24 -1322 0 feedthrough
rlabel pdiffusion 31 -1322 31 -1322 0 feedthrough
rlabel pdiffusion 38 -1322 38 -1322 0 feedthrough
rlabel pdiffusion 45 -1322 45 -1322 0 feedthrough
rlabel pdiffusion 52 -1322 52 -1322 0 feedthrough
rlabel pdiffusion 59 -1322 59 -1322 0 feedthrough
rlabel pdiffusion 66 -1322 66 -1322 0 feedthrough
rlabel pdiffusion 73 -1322 73 -1322 0 cellNo=75
rlabel pdiffusion 80 -1322 80 -1322 0 cellNo=864
rlabel pdiffusion 87 -1322 87 -1322 0 feedthrough
rlabel pdiffusion 94 -1322 94 -1322 0 cellNo=607
rlabel pdiffusion 101 -1322 101 -1322 0 feedthrough
rlabel pdiffusion 108 -1322 108 -1322 0 feedthrough
rlabel pdiffusion 115 -1322 115 -1322 0 feedthrough
rlabel pdiffusion 122 -1322 122 -1322 0 cellNo=496
rlabel pdiffusion 129 -1322 129 -1322 0 feedthrough
rlabel pdiffusion 136 -1322 136 -1322 0 feedthrough
rlabel pdiffusion 143 -1322 143 -1322 0 cellNo=48
rlabel pdiffusion 150 -1322 150 -1322 0 feedthrough
rlabel pdiffusion 157 -1322 157 -1322 0 feedthrough
rlabel pdiffusion 164 -1322 164 -1322 0 cellNo=644
rlabel pdiffusion 171 -1322 171 -1322 0 feedthrough
rlabel pdiffusion 178 -1322 178 -1322 0 feedthrough
rlabel pdiffusion 185 -1322 185 -1322 0 feedthrough
rlabel pdiffusion 192 -1322 192 -1322 0 feedthrough
rlabel pdiffusion 199 -1322 199 -1322 0 feedthrough
rlabel pdiffusion 206 -1322 206 -1322 0 feedthrough
rlabel pdiffusion 213 -1322 213 -1322 0 feedthrough
rlabel pdiffusion 220 -1322 220 -1322 0 feedthrough
rlabel pdiffusion 227 -1322 227 -1322 0 feedthrough
rlabel pdiffusion 234 -1322 234 -1322 0 cellNo=509
rlabel pdiffusion 241 -1322 241 -1322 0 feedthrough
rlabel pdiffusion 248 -1322 248 -1322 0 cellNo=325
rlabel pdiffusion 255 -1322 255 -1322 0 feedthrough
rlabel pdiffusion 262 -1322 262 -1322 0 feedthrough
rlabel pdiffusion 269 -1322 269 -1322 0 feedthrough
rlabel pdiffusion 276 -1322 276 -1322 0 cellNo=612
rlabel pdiffusion 283 -1322 283 -1322 0 feedthrough
rlabel pdiffusion 290 -1322 290 -1322 0 feedthrough
rlabel pdiffusion 297 -1322 297 -1322 0 feedthrough
rlabel pdiffusion 304 -1322 304 -1322 0 feedthrough
rlabel pdiffusion 311 -1322 311 -1322 0 feedthrough
rlabel pdiffusion 318 -1322 318 -1322 0 feedthrough
rlabel pdiffusion 325 -1322 325 -1322 0 feedthrough
rlabel pdiffusion 332 -1322 332 -1322 0 feedthrough
rlabel pdiffusion 339 -1322 339 -1322 0 feedthrough
rlabel pdiffusion 346 -1322 346 -1322 0 feedthrough
rlabel pdiffusion 353 -1322 353 -1322 0 feedthrough
rlabel pdiffusion 360 -1322 360 -1322 0 feedthrough
rlabel pdiffusion 367 -1322 367 -1322 0 feedthrough
rlabel pdiffusion 374 -1322 374 -1322 0 feedthrough
rlabel pdiffusion 381 -1322 381 -1322 0 feedthrough
rlabel pdiffusion 388 -1322 388 -1322 0 feedthrough
rlabel pdiffusion 395 -1322 395 -1322 0 feedthrough
rlabel pdiffusion 402 -1322 402 -1322 0 feedthrough
rlabel pdiffusion 409 -1322 409 -1322 0 feedthrough
rlabel pdiffusion 416 -1322 416 -1322 0 feedthrough
rlabel pdiffusion 423 -1322 423 -1322 0 cellNo=78
rlabel pdiffusion 430 -1322 430 -1322 0 feedthrough
rlabel pdiffusion 437 -1322 437 -1322 0 feedthrough
rlabel pdiffusion 444 -1322 444 -1322 0 feedthrough
rlabel pdiffusion 451 -1322 451 -1322 0 feedthrough
rlabel pdiffusion 458 -1322 458 -1322 0 cellNo=490
rlabel pdiffusion 465 -1322 465 -1322 0 feedthrough
rlabel pdiffusion 472 -1322 472 -1322 0 feedthrough
rlabel pdiffusion 479 -1322 479 -1322 0 cellNo=597
rlabel pdiffusion 486 -1322 486 -1322 0 feedthrough
rlabel pdiffusion 493 -1322 493 -1322 0 feedthrough
rlabel pdiffusion 500 -1322 500 -1322 0 feedthrough
rlabel pdiffusion 507 -1322 507 -1322 0 cellNo=247
rlabel pdiffusion 514 -1322 514 -1322 0 cellNo=820
rlabel pdiffusion 521 -1322 521 -1322 0 feedthrough
rlabel pdiffusion 528 -1322 528 -1322 0 cellNo=30
rlabel pdiffusion 535 -1322 535 -1322 0 feedthrough
rlabel pdiffusion 542 -1322 542 -1322 0 feedthrough
rlabel pdiffusion 549 -1322 549 -1322 0 feedthrough
rlabel pdiffusion 556 -1322 556 -1322 0 feedthrough
rlabel pdiffusion 563 -1322 563 -1322 0 feedthrough
rlabel pdiffusion 570 -1322 570 -1322 0 feedthrough
rlabel pdiffusion 577 -1322 577 -1322 0 cellNo=109
rlabel pdiffusion 584 -1322 584 -1322 0 feedthrough
rlabel pdiffusion 591 -1322 591 -1322 0 cellNo=257
rlabel pdiffusion 598 -1322 598 -1322 0 feedthrough
rlabel pdiffusion 605 -1322 605 -1322 0 feedthrough
rlabel pdiffusion 612 -1322 612 -1322 0 cellNo=230
rlabel pdiffusion 619 -1322 619 -1322 0 feedthrough
rlabel pdiffusion 626 -1322 626 -1322 0 cellNo=507
rlabel pdiffusion 633 -1322 633 -1322 0 feedthrough
rlabel pdiffusion 640 -1322 640 -1322 0 feedthrough
rlabel pdiffusion 647 -1322 647 -1322 0 feedthrough
rlabel pdiffusion 654 -1322 654 -1322 0 feedthrough
rlabel pdiffusion 661 -1322 661 -1322 0 cellNo=77
rlabel pdiffusion 668 -1322 668 -1322 0 feedthrough
rlabel pdiffusion 675 -1322 675 -1322 0 feedthrough
rlabel pdiffusion 682 -1322 682 -1322 0 feedthrough
rlabel pdiffusion 689 -1322 689 -1322 0 cellNo=8
rlabel pdiffusion 696 -1322 696 -1322 0 feedthrough
rlabel pdiffusion 703 -1322 703 -1322 0 feedthrough
rlabel pdiffusion 710 -1322 710 -1322 0 feedthrough
rlabel pdiffusion 717 -1322 717 -1322 0 feedthrough
rlabel pdiffusion 724 -1322 724 -1322 0 feedthrough
rlabel pdiffusion 731 -1322 731 -1322 0 feedthrough
rlabel pdiffusion 738 -1322 738 -1322 0 feedthrough
rlabel pdiffusion 745 -1322 745 -1322 0 feedthrough
rlabel pdiffusion 752 -1322 752 -1322 0 feedthrough
rlabel pdiffusion 759 -1322 759 -1322 0 feedthrough
rlabel pdiffusion 766 -1322 766 -1322 0 cellNo=113
rlabel pdiffusion 773 -1322 773 -1322 0 feedthrough
rlabel pdiffusion 780 -1322 780 -1322 0 feedthrough
rlabel pdiffusion 787 -1322 787 -1322 0 cellNo=273
rlabel pdiffusion 794 -1322 794 -1322 0 cellNo=544
rlabel pdiffusion 801 -1322 801 -1322 0 feedthrough
rlabel pdiffusion 808 -1322 808 -1322 0 cellNo=793
rlabel pdiffusion 815 -1322 815 -1322 0 cellNo=50
rlabel pdiffusion 822 -1322 822 -1322 0 cellNo=157
rlabel pdiffusion 829 -1322 829 -1322 0 cellNo=461
rlabel pdiffusion 836 -1322 836 -1322 0 feedthrough
rlabel pdiffusion 843 -1322 843 -1322 0 feedthrough
rlabel pdiffusion 850 -1322 850 -1322 0 feedthrough
rlabel pdiffusion 857 -1322 857 -1322 0 feedthrough
rlabel pdiffusion 864 -1322 864 -1322 0 feedthrough
rlabel pdiffusion 871 -1322 871 -1322 0 feedthrough
rlabel pdiffusion 878 -1322 878 -1322 0 feedthrough
rlabel pdiffusion 885 -1322 885 -1322 0 feedthrough
rlabel pdiffusion 892 -1322 892 -1322 0 feedthrough
rlabel pdiffusion 899 -1322 899 -1322 0 feedthrough
rlabel pdiffusion 906 -1322 906 -1322 0 feedthrough
rlabel pdiffusion 913 -1322 913 -1322 0 feedthrough
rlabel pdiffusion 920 -1322 920 -1322 0 feedthrough
rlabel pdiffusion 927 -1322 927 -1322 0 feedthrough
rlabel pdiffusion 934 -1322 934 -1322 0 cellNo=12
rlabel pdiffusion 941 -1322 941 -1322 0 feedthrough
rlabel pdiffusion 948 -1322 948 -1322 0 cellNo=589
rlabel pdiffusion 955 -1322 955 -1322 0 feedthrough
rlabel pdiffusion 962 -1322 962 -1322 0 feedthrough
rlabel pdiffusion 969 -1322 969 -1322 0 feedthrough
rlabel pdiffusion 976 -1322 976 -1322 0 cellNo=463
rlabel pdiffusion 983 -1322 983 -1322 0 cellNo=376
rlabel pdiffusion 990 -1322 990 -1322 0 feedthrough
rlabel pdiffusion 997 -1322 997 -1322 0 feedthrough
rlabel pdiffusion 1004 -1322 1004 -1322 0 feedthrough
rlabel pdiffusion 1011 -1322 1011 -1322 0 cellNo=111
rlabel pdiffusion 1018 -1322 1018 -1322 0 feedthrough
rlabel pdiffusion 1025 -1322 1025 -1322 0 feedthrough
rlabel pdiffusion 1032 -1322 1032 -1322 0 feedthrough
rlabel pdiffusion 1039 -1322 1039 -1322 0 feedthrough
rlabel pdiffusion 1046 -1322 1046 -1322 0 feedthrough
rlabel pdiffusion 1053 -1322 1053 -1322 0 cellNo=261
rlabel pdiffusion 1060 -1322 1060 -1322 0 feedthrough
rlabel pdiffusion 1067 -1322 1067 -1322 0 feedthrough
rlabel pdiffusion 1074 -1322 1074 -1322 0 feedthrough
rlabel pdiffusion 1081 -1322 1081 -1322 0 feedthrough
rlabel pdiffusion 1088 -1322 1088 -1322 0 feedthrough
rlabel pdiffusion 1095 -1322 1095 -1322 0 feedthrough
rlabel pdiffusion 1102 -1322 1102 -1322 0 feedthrough
rlabel pdiffusion 1109 -1322 1109 -1322 0 feedthrough
rlabel pdiffusion 1116 -1322 1116 -1322 0 feedthrough
rlabel pdiffusion 1123 -1322 1123 -1322 0 feedthrough
rlabel pdiffusion 1130 -1322 1130 -1322 0 feedthrough
rlabel pdiffusion 1137 -1322 1137 -1322 0 feedthrough
rlabel pdiffusion 1144 -1322 1144 -1322 0 feedthrough
rlabel pdiffusion 1151 -1322 1151 -1322 0 feedthrough
rlabel pdiffusion 1158 -1322 1158 -1322 0 feedthrough
rlabel pdiffusion 1165 -1322 1165 -1322 0 feedthrough
rlabel pdiffusion 1172 -1322 1172 -1322 0 feedthrough
rlabel pdiffusion 1179 -1322 1179 -1322 0 feedthrough
rlabel pdiffusion 1186 -1322 1186 -1322 0 feedthrough
rlabel pdiffusion 1193 -1322 1193 -1322 0 feedthrough
rlabel pdiffusion 1200 -1322 1200 -1322 0 feedthrough
rlabel pdiffusion 1207 -1322 1207 -1322 0 feedthrough
rlabel pdiffusion 1214 -1322 1214 -1322 0 feedthrough
rlabel pdiffusion 1221 -1322 1221 -1322 0 feedthrough
rlabel pdiffusion 1228 -1322 1228 -1322 0 feedthrough
rlabel pdiffusion 1235 -1322 1235 -1322 0 feedthrough
rlabel pdiffusion 1242 -1322 1242 -1322 0 feedthrough
rlabel pdiffusion 1249 -1322 1249 -1322 0 feedthrough
rlabel pdiffusion 1256 -1322 1256 -1322 0 feedthrough
rlabel pdiffusion 1263 -1322 1263 -1322 0 feedthrough
rlabel pdiffusion 1270 -1322 1270 -1322 0 feedthrough
rlabel pdiffusion 1277 -1322 1277 -1322 0 feedthrough
rlabel pdiffusion 1284 -1322 1284 -1322 0 feedthrough
rlabel pdiffusion 1291 -1322 1291 -1322 0 feedthrough
rlabel pdiffusion 1298 -1322 1298 -1322 0 feedthrough
rlabel pdiffusion 1305 -1322 1305 -1322 0 feedthrough
rlabel pdiffusion 1312 -1322 1312 -1322 0 feedthrough
rlabel pdiffusion 1319 -1322 1319 -1322 0 feedthrough
rlabel pdiffusion 1326 -1322 1326 -1322 0 feedthrough
rlabel pdiffusion 1333 -1322 1333 -1322 0 feedthrough
rlabel pdiffusion 1340 -1322 1340 -1322 0 feedthrough
rlabel pdiffusion 1347 -1322 1347 -1322 0 feedthrough
rlabel pdiffusion 1354 -1322 1354 -1322 0 cellNo=269
rlabel pdiffusion 1361 -1322 1361 -1322 0 feedthrough
rlabel pdiffusion 1368 -1322 1368 -1322 0 feedthrough
rlabel pdiffusion 1375 -1322 1375 -1322 0 feedthrough
rlabel pdiffusion 1382 -1322 1382 -1322 0 feedthrough
rlabel pdiffusion 1389 -1322 1389 -1322 0 feedthrough
rlabel pdiffusion 1396 -1322 1396 -1322 0 feedthrough
rlabel pdiffusion 1403 -1322 1403 -1322 0 feedthrough
rlabel pdiffusion 1410 -1322 1410 -1322 0 feedthrough
rlabel pdiffusion 1417 -1322 1417 -1322 0 feedthrough
rlabel pdiffusion 1424 -1322 1424 -1322 0 feedthrough
rlabel pdiffusion 1431 -1322 1431 -1322 0 feedthrough
rlabel pdiffusion 1438 -1322 1438 -1322 0 feedthrough
rlabel pdiffusion 1445 -1322 1445 -1322 0 feedthrough
rlabel pdiffusion 1452 -1322 1452 -1322 0 feedthrough
rlabel pdiffusion 1459 -1322 1459 -1322 0 feedthrough
rlabel pdiffusion 1466 -1322 1466 -1322 0 feedthrough
rlabel pdiffusion 1473 -1322 1473 -1322 0 feedthrough
rlabel pdiffusion 1480 -1322 1480 -1322 0 feedthrough
rlabel pdiffusion 1487 -1322 1487 -1322 0 feedthrough
rlabel pdiffusion 1494 -1322 1494 -1322 0 feedthrough
rlabel pdiffusion 1501 -1322 1501 -1322 0 feedthrough
rlabel pdiffusion 1508 -1322 1508 -1322 0 feedthrough
rlabel pdiffusion 1515 -1322 1515 -1322 0 feedthrough
rlabel pdiffusion 1522 -1322 1522 -1322 0 feedthrough
rlabel pdiffusion 1529 -1322 1529 -1322 0 feedthrough
rlabel pdiffusion 1536 -1322 1536 -1322 0 feedthrough
rlabel pdiffusion 1543 -1322 1543 -1322 0 feedthrough
rlabel pdiffusion 1550 -1322 1550 -1322 0 feedthrough
rlabel pdiffusion 1557 -1322 1557 -1322 0 feedthrough
rlabel pdiffusion 1564 -1322 1564 -1322 0 feedthrough
rlabel pdiffusion 1571 -1322 1571 -1322 0 feedthrough
rlabel pdiffusion 1578 -1322 1578 -1322 0 feedthrough
rlabel pdiffusion 1585 -1322 1585 -1322 0 feedthrough
rlabel pdiffusion 1592 -1322 1592 -1322 0 feedthrough
rlabel pdiffusion 1599 -1322 1599 -1322 0 feedthrough
rlabel pdiffusion 1606 -1322 1606 -1322 0 feedthrough
rlabel pdiffusion 1613 -1322 1613 -1322 0 feedthrough
rlabel pdiffusion 1620 -1322 1620 -1322 0 feedthrough
rlabel pdiffusion 1627 -1322 1627 -1322 0 feedthrough
rlabel pdiffusion 1634 -1322 1634 -1322 0 feedthrough
rlabel pdiffusion 1641 -1322 1641 -1322 0 feedthrough
rlabel pdiffusion 1648 -1322 1648 -1322 0 feedthrough
rlabel pdiffusion 1655 -1322 1655 -1322 0 feedthrough
rlabel pdiffusion 1662 -1322 1662 -1322 0 feedthrough
rlabel pdiffusion 1669 -1322 1669 -1322 0 feedthrough
rlabel pdiffusion 1676 -1322 1676 -1322 0 feedthrough
rlabel pdiffusion 1683 -1322 1683 -1322 0 feedthrough
rlabel pdiffusion 1690 -1322 1690 -1322 0 feedthrough
rlabel pdiffusion 1697 -1322 1697 -1322 0 feedthrough
rlabel pdiffusion 1704 -1322 1704 -1322 0 cellNo=876
rlabel pdiffusion 1711 -1322 1711 -1322 0 cellNo=21
rlabel pdiffusion 1718 -1322 1718 -1322 0 feedthrough
rlabel pdiffusion 1725 -1322 1725 -1322 0 feedthrough
rlabel pdiffusion 1732 -1322 1732 -1322 0 cellNo=797
rlabel pdiffusion 1739 -1322 1739 -1322 0 feedthrough
rlabel pdiffusion 3 -1477 3 -1477 0 cellNo=1281
rlabel pdiffusion 10 -1477 10 -1477 0 cellNo=1286
rlabel pdiffusion 17 -1477 17 -1477 0 feedthrough
rlabel pdiffusion 24 -1477 24 -1477 0 cellNo=277
rlabel pdiffusion 31 -1477 31 -1477 0 feedthrough
rlabel pdiffusion 38 -1477 38 -1477 0 feedthrough
rlabel pdiffusion 45 -1477 45 -1477 0 feedthrough
rlabel pdiffusion 52 -1477 52 -1477 0 feedthrough
rlabel pdiffusion 59 -1477 59 -1477 0 cellNo=745
rlabel pdiffusion 66 -1477 66 -1477 0 feedthrough
rlabel pdiffusion 73 -1477 73 -1477 0 cellNo=800
rlabel pdiffusion 80 -1477 80 -1477 0 cellNo=849
rlabel pdiffusion 87 -1477 87 -1477 0 feedthrough
rlabel pdiffusion 94 -1477 94 -1477 0 cellNo=34
rlabel pdiffusion 101 -1477 101 -1477 0 feedthrough
rlabel pdiffusion 108 -1477 108 -1477 0 cellNo=424
rlabel pdiffusion 115 -1477 115 -1477 0 cellNo=119
rlabel pdiffusion 122 -1477 122 -1477 0 feedthrough
rlabel pdiffusion 129 -1477 129 -1477 0 feedthrough
rlabel pdiffusion 136 -1477 136 -1477 0 feedthrough
rlabel pdiffusion 143 -1477 143 -1477 0 feedthrough
rlabel pdiffusion 150 -1477 150 -1477 0 feedthrough
rlabel pdiffusion 157 -1477 157 -1477 0 cellNo=611
rlabel pdiffusion 164 -1477 164 -1477 0 feedthrough
rlabel pdiffusion 171 -1477 171 -1477 0 feedthrough
rlabel pdiffusion 178 -1477 178 -1477 0 feedthrough
rlabel pdiffusion 185 -1477 185 -1477 0 feedthrough
rlabel pdiffusion 192 -1477 192 -1477 0 feedthrough
rlabel pdiffusion 199 -1477 199 -1477 0 feedthrough
rlabel pdiffusion 206 -1477 206 -1477 0 feedthrough
rlabel pdiffusion 213 -1477 213 -1477 0 feedthrough
rlabel pdiffusion 220 -1477 220 -1477 0 cellNo=24
rlabel pdiffusion 227 -1477 227 -1477 0 cellNo=459
rlabel pdiffusion 234 -1477 234 -1477 0 feedthrough
rlabel pdiffusion 241 -1477 241 -1477 0 feedthrough
rlabel pdiffusion 248 -1477 248 -1477 0 feedthrough
rlabel pdiffusion 255 -1477 255 -1477 0 feedthrough
rlabel pdiffusion 262 -1477 262 -1477 0 cellNo=928
rlabel pdiffusion 269 -1477 269 -1477 0 feedthrough
rlabel pdiffusion 276 -1477 276 -1477 0 feedthrough
rlabel pdiffusion 283 -1477 283 -1477 0 feedthrough
rlabel pdiffusion 290 -1477 290 -1477 0 feedthrough
rlabel pdiffusion 297 -1477 297 -1477 0 cellNo=15
rlabel pdiffusion 304 -1477 304 -1477 0 feedthrough
rlabel pdiffusion 311 -1477 311 -1477 0 feedthrough
rlabel pdiffusion 318 -1477 318 -1477 0 feedthrough
rlabel pdiffusion 325 -1477 325 -1477 0 feedthrough
rlabel pdiffusion 332 -1477 332 -1477 0 feedthrough
rlabel pdiffusion 339 -1477 339 -1477 0 feedthrough
rlabel pdiffusion 346 -1477 346 -1477 0 feedthrough
rlabel pdiffusion 353 -1477 353 -1477 0 feedthrough
rlabel pdiffusion 360 -1477 360 -1477 0 feedthrough
rlabel pdiffusion 367 -1477 367 -1477 0 feedthrough
rlabel pdiffusion 374 -1477 374 -1477 0 feedthrough
rlabel pdiffusion 381 -1477 381 -1477 0 feedthrough
rlabel pdiffusion 388 -1477 388 -1477 0 cellNo=594
rlabel pdiffusion 395 -1477 395 -1477 0 feedthrough
rlabel pdiffusion 402 -1477 402 -1477 0 feedthrough
rlabel pdiffusion 409 -1477 409 -1477 0 cellNo=700
rlabel pdiffusion 416 -1477 416 -1477 0 cellNo=60
rlabel pdiffusion 423 -1477 423 -1477 0 feedthrough
rlabel pdiffusion 430 -1477 430 -1477 0 feedthrough
rlabel pdiffusion 437 -1477 437 -1477 0 feedthrough
rlabel pdiffusion 444 -1477 444 -1477 0 feedthrough
rlabel pdiffusion 451 -1477 451 -1477 0 feedthrough
rlabel pdiffusion 458 -1477 458 -1477 0 feedthrough
rlabel pdiffusion 465 -1477 465 -1477 0 feedthrough
rlabel pdiffusion 472 -1477 472 -1477 0 feedthrough
rlabel pdiffusion 479 -1477 479 -1477 0 feedthrough
rlabel pdiffusion 486 -1477 486 -1477 0 feedthrough
rlabel pdiffusion 493 -1477 493 -1477 0 feedthrough
rlabel pdiffusion 500 -1477 500 -1477 0 cellNo=866
rlabel pdiffusion 507 -1477 507 -1477 0 feedthrough
rlabel pdiffusion 514 -1477 514 -1477 0 feedthrough
rlabel pdiffusion 521 -1477 521 -1477 0 feedthrough
rlabel pdiffusion 528 -1477 528 -1477 0 feedthrough
rlabel pdiffusion 535 -1477 535 -1477 0 feedthrough
rlabel pdiffusion 542 -1477 542 -1477 0 feedthrough
rlabel pdiffusion 549 -1477 549 -1477 0 feedthrough
rlabel pdiffusion 556 -1477 556 -1477 0 cellNo=454
rlabel pdiffusion 563 -1477 563 -1477 0 feedthrough
rlabel pdiffusion 570 -1477 570 -1477 0 feedthrough
rlabel pdiffusion 577 -1477 577 -1477 0 feedthrough
rlabel pdiffusion 584 -1477 584 -1477 0 feedthrough
rlabel pdiffusion 591 -1477 591 -1477 0 cellNo=413
rlabel pdiffusion 598 -1477 598 -1477 0 cellNo=468
rlabel pdiffusion 605 -1477 605 -1477 0 feedthrough
rlabel pdiffusion 612 -1477 612 -1477 0 cellNo=542
rlabel pdiffusion 619 -1477 619 -1477 0 feedthrough
rlabel pdiffusion 626 -1477 626 -1477 0 feedthrough
rlabel pdiffusion 633 -1477 633 -1477 0 cellNo=276
rlabel pdiffusion 640 -1477 640 -1477 0 cellNo=674
rlabel pdiffusion 647 -1477 647 -1477 0 feedthrough
rlabel pdiffusion 654 -1477 654 -1477 0 feedthrough
rlabel pdiffusion 661 -1477 661 -1477 0 feedthrough
rlabel pdiffusion 668 -1477 668 -1477 0 feedthrough
rlabel pdiffusion 675 -1477 675 -1477 0 cellNo=304
rlabel pdiffusion 682 -1477 682 -1477 0 feedthrough
rlabel pdiffusion 689 -1477 689 -1477 0 feedthrough
rlabel pdiffusion 696 -1477 696 -1477 0 feedthrough
rlabel pdiffusion 703 -1477 703 -1477 0 feedthrough
rlabel pdiffusion 710 -1477 710 -1477 0 feedthrough
rlabel pdiffusion 717 -1477 717 -1477 0 cellNo=803
rlabel pdiffusion 724 -1477 724 -1477 0 cellNo=338
rlabel pdiffusion 731 -1477 731 -1477 0 cellNo=456
rlabel pdiffusion 738 -1477 738 -1477 0 feedthrough
rlabel pdiffusion 745 -1477 745 -1477 0 feedthrough
rlabel pdiffusion 752 -1477 752 -1477 0 feedthrough
rlabel pdiffusion 759 -1477 759 -1477 0 feedthrough
rlabel pdiffusion 766 -1477 766 -1477 0 cellNo=978
rlabel pdiffusion 773 -1477 773 -1477 0 feedthrough
rlabel pdiffusion 780 -1477 780 -1477 0 feedthrough
rlabel pdiffusion 787 -1477 787 -1477 0 feedthrough
rlabel pdiffusion 794 -1477 794 -1477 0 feedthrough
rlabel pdiffusion 801 -1477 801 -1477 0 feedthrough
rlabel pdiffusion 808 -1477 808 -1477 0 feedthrough
rlabel pdiffusion 815 -1477 815 -1477 0 feedthrough
rlabel pdiffusion 822 -1477 822 -1477 0 feedthrough
rlabel pdiffusion 829 -1477 829 -1477 0 feedthrough
rlabel pdiffusion 836 -1477 836 -1477 0 feedthrough
rlabel pdiffusion 843 -1477 843 -1477 0 feedthrough
rlabel pdiffusion 850 -1477 850 -1477 0 feedthrough
rlabel pdiffusion 857 -1477 857 -1477 0 feedthrough
rlabel pdiffusion 864 -1477 864 -1477 0 cellNo=773
rlabel pdiffusion 871 -1477 871 -1477 0 cellNo=191
rlabel pdiffusion 878 -1477 878 -1477 0 feedthrough
rlabel pdiffusion 885 -1477 885 -1477 0 feedthrough
rlabel pdiffusion 892 -1477 892 -1477 0 cellNo=286
rlabel pdiffusion 899 -1477 899 -1477 0 cellNo=736
rlabel pdiffusion 906 -1477 906 -1477 0 feedthrough
rlabel pdiffusion 913 -1477 913 -1477 0 feedthrough
rlabel pdiffusion 920 -1477 920 -1477 0 feedthrough
rlabel pdiffusion 927 -1477 927 -1477 0 feedthrough
rlabel pdiffusion 934 -1477 934 -1477 0 cellNo=922
rlabel pdiffusion 941 -1477 941 -1477 0 feedthrough
rlabel pdiffusion 948 -1477 948 -1477 0 feedthrough
rlabel pdiffusion 955 -1477 955 -1477 0 feedthrough
rlabel pdiffusion 962 -1477 962 -1477 0 feedthrough
rlabel pdiffusion 969 -1477 969 -1477 0 feedthrough
rlabel pdiffusion 976 -1477 976 -1477 0 feedthrough
rlabel pdiffusion 983 -1477 983 -1477 0 feedthrough
rlabel pdiffusion 990 -1477 990 -1477 0 feedthrough
rlabel pdiffusion 997 -1477 997 -1477 0 feedthrough
rlabel pdiffusion 1004 -1477 1004 -1477 0 feedthrough
rlabel pdiffusion 1011 -1477 1011 -1477 0 feedthrough
rlabel pdiffusion 1018 -1477 1018 -1477 0 feedthrough
rlabel pdiffusion 1025 -1477 1025 -1477 0 cellNo=821
rlabel pdiffusion 1032 -1477 1032 -1477 0 feedthrough
rlabel pdiffusion 1039 -1477 1039 -1477 0 feedthrough
rlabel pdiffusion 1046 -1477 1046 -1477 0 feedthrough
rlabel pdiffusion 1053 -1477 1053 -1477 0 feedthrough
rlabel pdiffusion 1060 -1477 1060 -1477 0 feedthrough
rlabel pdiffusion 1067 -1477 1067 -1477 0 cellNo=268
rlabel pdiffusion 1074 -1477 1074 -1477 0 feedthrough
rlabel pdiffusion 1081 -1477 1081 -1477 0 feedthrough
rlabel pdiffusion 1088 -1477 1088 -1477 0 feedthrough
rlabel pdiffusion 1095 -1477 1095 -1477 0 feedthrough
rlabel pdiffusion 1102 -1477 1102 -1477 0 feedthrough
rlabel pdiffusion 1109 -1477 1109 -1477 0 feedthrough
rlabel pdiffusion 1116 -1477 1116 -1477 0 feedthrough
rlabel pdiffusion 1123 -1477 1123 -1477 0 cellNo=436
rlabel pdiffusion 1130 -1477 1130 -1477 0 feedthrough
rlabel pdiffusion 1137 -1477 1137 -1477 0 cellNo=341
rlabel pdiffusion 1144 -1477 1144 -1477 0 cellNo=790
rlabel pdiffusion 1151 -1477 1151 -1477 0 feedthrough
rlabel pdiffusion 1158 -1477 1158 -1477 0 feedthrough
rlabel pdiffusion 1165 -1477 1165 -1477 0 feedthrough
rlabel pdiffusion 1172 -1477 1172 -1477 0 feedthrough
rlabel pdiffusion 1179 -1477 1179 -1477 0 feedthrough
rlabel pdiffusion 1186 -1477 1186 -1477 0 feedthrough
rlabel pdiffusion 1193 -1477 1193 -1477 0 feedthrough
rlabel pdiffusion 1200 -1477 1200 -1477 0 feedthrough
rlabel pdiffusion 1207 -1477 1207 -1477 0 feedthrough
rlabel pdiffusion 1214 -1477 1214 -1477 0 feedthrough
rlabel pdiffusion 1221 -1477 1221 -1477 0 feedthrough
rlabel pdiffusion 1228 -1477 1228 -1477 0 feedthrough
rlabel pdiffusion 1235 -1477 1235 -1477 0 feedthrough
rlabel pdiffusion 1242 -1477 1242 -1477 0 feedthrough
rlabel pdiffusion 1249 -1477 1249 -1477 0 feedthrough
rlabel pdiffusion 1256 -1477 1256 -1477 0 feedthrough
rlabel pdiffusion 1263 -1477 1263 -1477 0 feedthrough
rlabel pdiffusion 1270 -1477 1270 -1477 0 feedthrough
rlabel pdiffusion 1277 -1477 1277 -1477 0 feedthrough
rlabel pdiffusion 1284 -1477 1284 -1477 0 feedthrough
rlabel pdiffusion 1291 -1477 1291 -1477 0 feedthrough
rlabel pdiffusion 1298 -1477 1298 -1477 0 feedthrough
rlabel pdiffusion 1305 -1477 1305 -1477 0 feedthrough
rlabel pdiffusion 1312 -1477 1312 -1477 0 feedthrough
rlabel pdiffusion 1319 -1477 1319 -1477 0 feedthrough
rlabel pdiffusion 1326 -1477 1326 -1477 0 feedthrough
rlabel pdiffusion 1333 -1477 1333 -1477 0 feedthrough
rlabel pdiffusion 1340 -1477 1340 -1477 0 feedthrough
rlabel pdiffusion 1347 -1477 1347 -1477 0 feedthrough
rlabel pdiffusion 1354 -1477 1354 -1477 0 feedthrough
rlabel pdiffusion 1361 -1477 1361 -1477 0 feedthrough
rlabel pdiffusion 1368 -1477 1368 -1477 0 feedthrough
rlabel pdiffusion 1375 -1477 1375 -1477 0 feedthrough
rlabel pdiffusion 1382 -1477 1382 -1477 0 feedthrough
rlabel pdiffusion 1389 -1477 1389 -1477 0 feedthrough
rlabel pdiffusion 1396 -1477 1396 -1477 0 feedthrough
rlabel pdiffusion 1403 -1477 1403 -1477 0 feedthrough
rlabel pdiffusion 1410 -1477 1410 -1477 0 feedthrough
rlabel pdiffusion 1417 -1477 1417 -1477 0 feedthrough
rlabel pdiffusion 1424 -1477 1424 -1477 0 feedthrough
rlabel pdiffusion 1431 -1477 1431 -1477 0 feedthrough
rlabel pdiffusion 1438 -1477 1438 -1477 0 feedthrough
rlabel pdiffusion 1445 -1477 1445 -1477 0 feedthrough
rlabel pdiffusion 1452 -1477 1452 -1477 0 feedthrough
rlabel pdiffusion 1459 -1477 1459 -1477 0 feedthrough
rlabel pdiffusion 1466 -1477 1466 -1477 0 feedthrough
rlabel pdiffusion 1473 -1477 1473 -1477 0 feedthrough
rlabel pdiffusion 1480 -1477 1480 -1477 0 feedthrough
rlabel pdiffusion 1487 -1477 1487 -1477 0 feedthrough
rlabel pdiffusion 1494 -1477 1494 -1477 0 feedthrough
rlabel pdiffusion 1501 -1477 1501 -1477 0 feedthrough
rlabel pdiffusion 1508 -1477 1508 -1477 0 feedthrough
rlabel pdiffusion 1515 -1477 1515 -1477 0 feedthrough
rlabel pdiffusion 1522 -1477 1522 -1477 0 feedthrough
rlabel pdiffusion 1529 -1477 1529 -1477 0 feedthrough
rlabel pdiffusion 1536 -1477 1536 -1477 0 feedthrough
rlabel pdiffusion 1543 -1477 1543 -1477 0 feedthrough
rlabel pdiffusion 1550 -1477 1550 -1477 0 feedthrough
rlabel pdiffusion 1557 -1477 1557 -1477 0 feedthrough
rlabel pdiffusion 1564 -1477 1564 -1477 0 feedthrough
rlabel pdiffusion 1571 -1477 1571 -1477 0 feedthrough
rlabel pdiffusion 1578 -1477 1578 -1477 0 feedthrough
rlabel pdiffusion 1585 -1477 1585 -1477 0 feedthrough
rlabel pdiffusion 1592 -1477 1592 -1477 0 feedthrough
rlabel pdiffusion 1599 -1477 1599 -1477 0 feedthrough
rlabel pdiffusion 1606 -1477 1606 -1477 0 feedthrough
rlabel pdiffusion 1613 -1477 1613 -1477 0 feedthrough
rlabel pdiffusion 1620 -1477 1620 -1477 0 feedthrough
rlabel pdiffusion 1627 -1477 1627 -1477 0 feedthrough
rlabel pdiffusion 1634 -1477 1634 -1477 0 feedthrough
rlabel pdiffusion 1641 -1477 1641 -1477 0 feedthrough
rlabel pdiffusion 1648 -1477 1648 -1477 0 feedthrough
rlabel pdiffusion 1655 -1477 1655 -1477 0 feedthrough
rlabel pdiffusion 1662 -1477 1662 -1477 0 feedthrough
rlabel pdiffusion 1669 -1477 1669 -1477 0 feedthrough
rlabel pdiffusion 1676 -1477 1676 -1477 0 feedthrough
rlabel pdiffusion 1683 -1477 1683 -1477 0 feedthrough
rlabel pdiffusion 1690 -1477 1690 -1477 0 feedthrough
rlabel pdiffusion 1697 -1477 1697 -1477 0 cellNo=558
rlabel pdiffusion 1704 -1477 1704 -1477 0 feedthrough
rlabel pdiffusion 1711 -1477 1711 -1477 0 feedthrough
rlabel pdiffusion 1718 -1477 1718 -1477 0 cellNo=653
rlabel pdiffusion 1725 -1477 1725 -1477 0 feedthrough
rlabel pdiffusion 1746 -1477 1746 -1477 0 feedthrough
rlabel pdiffusion 3 -1614 3 -1614 0 cellNo=1021
rlabel pdiffusion 10 -1614 10 -1614 0 cellNo=1088
rlabel pdiffusion 17 -1614 17 -1614 0 cellNo=1144
rlabel pdiffusion 24 -1614 24 -1614 0 feedthrough
rlabel pdiffusion 31 -1614 31 -1614 0 feedthrough
rlabel pdiffusion 38 -1614 38 -1614 0 cellNo=1042
rlabel pdiffusion 45 -1614 45 -1614 0 feedthrough
rlabel pdiffusion 52 -1614 52 -1614 0 feedthrough
rlabel pdiffusion 59 -1614 59 -1614 0 cellNo=772
rlabel pdiffusion 66 -1614 66 -1614 0 cellNo=801
rlabel pdiffusion 73 -1614 73 -1614 0 feedthrough
rlabel pdiffusion 80 -1614 80 -1614 0 feedthrough
rlabel pdiffusion 87 -1614 87 -1614 0 feedthrough
rlabel pdiffusion 94 -1614 94 -1614 0 cellNo=504
rlabel pdiffusion 101 -1614 101 -1614 0 feedthrough
rlabel pdiffusion 108 -1614 108 -1614 0 feedthrough
rlabel pdiffusion 115 -1614 115 -1614 0 feedthrough
rlabel pdiffusion 122 -1614 122 -1614 0 feedthrough
rlabel pdiffusion 129 -1614 129 -1614 0 feedthrough
rlabel pdiffusion 136 -1614 136 -1614 0 feedthrough
rlabel pdiffusion 143 -1614 143 -1614 0 feedthrough
rlabel pdiffusion 150 -1614 150 -1614 0 feedthrough
rlabel pdiffusion 157 -1614 157 -1614 0 feedthrough
rlabel pdiffusion 164 -1614 164 -1614 0 feedthrough
rlabel pdiffusion 171 -1614 171 -1614 0 feedthrough
rlabel pdiffusion 178 -1614 178 -1614 0 feedthrough
rlabel pdiffusion 185 -1614 185 -1614 0 feedthrough
rlabel pdiffusion 192 -1614 192 -1614 0 cellNo=699
rlabel pdiffusion 199 -1614 199 -1614 0 feedthrough
rlabel pdiffusion 206 -1614 206 -1614 0 cellNo=219
rlabel pdiffusion 213 -1614 213 -1614 0 feedthrough
rlabel pdiffusion 220 -1614 220 -1614 0 feedthrough
rlabel pdiffusion 227 -1614 227 -1614 0 feedthrough
rlabel pdiffusion 234 -1614 234 -1614 0 feedthrough
rlabel pdiffusion 241 -1614 241 -1614 0 feedthrough
rlabel pdiffusion 248 -1614 248 -1614 0 feedthrough
rlabel pdiffusion 255 -1614 255 -1614 0 cellNo=404
rlabel pdiffusion 262 -1614 262 -1614 0 feedthrough
rlabel pdiffusion 269 -1614 269 -1614 0 cellNo=615
rlabel pdiffusion 276 -1614 276 -1614 0 feedthrough
rlabel pdiffusion 283 -1614 283 -1614 0 feedthrough
rlabel pdiffusion 290 -1614 290 -1614 0 cellNo=439
rlabel pdiffusion 297 -1614 297 -1614 0 feedthrough
rlabel pdiffusion 304 -1614 304 -1614 0 feedthrough
rlabel pdiffusion 311 -1614 311 -1614 0 feedthrough
rlabel pdiffusion 318 -1614 318 -1614 0 cellNo=211
rlabel pdiffusion 325 -1614 325 -1614 0 feedthrough
rlabel pdiffusion 332 -1614 332 -1614 0 feedthrough
rlabel pdiffusion 339 -1614 339 -1614 0 feedthrough
rlabel pdiffusion 346 -1614 346 -1614 0 feedthrough
rlabel pdiffusion 353 -1614 353 -1614 0 feedthrough
rlabel pdiffusion 360 -1614 360 -1614 0 feedthrough
rlabel pdiffusion 367 -1614 367 -1614 0 cellNo=188
rlabel pdiffusion 374 -1614 374 -1614 0 feedthrough
rlabel pdiffusion 381 -1614 381 -1614 0 cellNo=491
rlabel pdiffusion 388 -1614 388 -1614 0 feedthrough
rlabel pdiffusion 395 -1614 395 -1614 0 feedthrough
rlabel pdiffusion 402 -1614 402 -1614 0 feedthrough
rlabel pdiffusion 409 -1614 409 -1614 0 feedthrough
rlabel pdiffusion 416 -1614 416 -1614 0 feedthrough
rlabel pdiffusion 423 -1614 423 -1614 0 feedthrough
rlabel pdiffusion 430 -1614 430 -1614 0 feedthrough
rlabel pdiffusion 437 -1614 437 -1614 0 feedthrough
rlabel pdiffusion 444 -1614 444 -1614 0 feedthrough
rlabel pdiffusion 451 -1614 451 -1614 0 feedthrough
rlabel pdiffusion 458 -1614 458 -1614 0 feedthrough
rlabel pdiffusion 465 -1614 465 -1614 0 feedthrough
rlabel pdiffusion 472 -1614 472 -1614 0 cellNo=306
rlabel pdiffusion 479 -1614 479 -1614 0 feedthrough
rlabel pdiffusion 486 -1614 486 -1614 0 feedthrough
rlabel pdiffusion 493 -1614 493 -1614 0 cellNo=657
rlabel pdiffusion 500 -1614 500 -1614 0 feedthrough
rlabel pdiffusion 507 -1614 507 -1614 0 feedthrough
rlabel pdiffusion 514 -1614 514 -1614 0 feedthrough
rlabel pdiffusion 521 -1614 521 -1614 0 feedthrough
rlabel pdiffusion 528 -1614 528 -1614 0 cellNo=613
rlabel pdiffusion 535 -1614 535 -1614 0 feedthrough
rlabel pdiffusion 542 -1614 542 -1614 0 cellNo=177
rlabel pdiffusion 549 -1614 549 -1614 0 feedthrough
rlabel pdiffusion 556 -1614 556 -1614 0 feedthrough
rlabel pdiffusion 563 -1614 563 -1614 0 cellNo=455
rlabel pdiffusion 570 -1614 570 -1614 0 feedthrough
rlabel pdiffusion 577 -1614 577 -1614 0 feedthrough
rlabel pdiffusion 584 -1614 584 -1614 0 feedthrough
rlabel pdiffusion 591 -1614 591 -1614 0 feedthrough
rlabel pdiffusion 598 -1614 598 -1614 0 feedthrough
rlabel pdiffusion 605 -1614 605 -1614 0 cellNo=760
rlabel pdiffusion 612 -1614 612 -1614 0 cellNo=771
rlabel pdiffusion 619 -1614 619 -1614 0 cellNo=741
rlabel pdiffusion 626 -1614 626 -1614 0 feedthrough
rlabel pdiffusion 633 -1614 633 -1614 0 feedthrough
rlabel pdiffusion 640 -1614 640 -1614 0 feedthrough
rlabel pdiffusion 647 -1614 647 -1614 0 feedthrough
rlabel pdiffusion 654 -1614 654 -1614 0 feedthrough
rlabel pdiffusion 661 -1614 661 -1614 0 feedthrough
rlabel pdiffusion 668 -1614 668 -1614 0 cellNo=135
rlabel pdiffusion 675 -1614 675 -1614 0 feedthrough
rlabel pdiffusion 682 -1614 682 -1614 0 feedthrough
rlabel pdiffusion 689 -1614 689 -1614 0 feedthrough
rlabel pdiffusion 696 -1614 696 -1614 0 feedthrough
rlabel pdiffusion 703 -1614 703 -1614 0 feedthrough
rlabel pdiffusion 710 -1614 710 -1614 0 cellNo=645
rlabel pdiffusion 717 -1614 717 -1614 0 cellNo=378
rlabel pdiffusion 724 -1614 724 -1614 0 cellNo=406
rlabel pdiffusion 731 -1614 731 -1614 0 feedthrough
rlabel pdiffusion 738 -1614 738 -1614 0 cellNo=1000
rlabel pdiffusion 745 -1614 745 -1614 0 cellNo=564
rlabel pdiffusion 752 -1614 752 -1614 0 feedthrough
rlabel pdiffusion 759 -1614 759 -1614 0 cellNo=684
rlabel pdiffusion 766 -1614 766 -1614 0 feedthrough
rlabel pdiffusion 773 -1614 773 -1614 0 feedthrough
rlabel pdiffusion 780 -1614 780 -1614 0 feedthrough
rlabel pdiffusion 787 -1614 787 -1614 0 feedthrough
rlabel pdiffusion 794 -1614 794 -1614 0 cellNo=285
rlabel pdiffusion 801 -1614 801 -1614 0 feedthrough
rlabel pdiffusion 808 -1614 808 -1614 0 cellNo=62
rlabel pdiffusion 815 -1614 815 -1614 0 feedthrough
rlabel pdiffusion 822 -1614 822 -1614 0 feedthrough
rlabel pdiffusion 829 -1614 829 -1614 0 feedthrough
rlabel pdiffusion 836 -1614 836 -1614 0 feedthrough
rlabel pdiffusion 843 -1614 843 -1614 0 feedthrough
rlabel pdiffusion 850 -1614 850 -1614 0 feedthrough
rlabel pdiffusion 857 -1614 857 -1614 0 feedthrough
rlabel pdiffusion 864 -1614 864 -1614 0 feedthrough
rlabel pdiffusion 871 -1614 871 -1614 0 feedthrough
rlabel pdiffusion 878 -1614 878 -1614 0 feedthrough
rlabel pdiffusion 885 -1614 885 -1614 0 feedthrough
rlabel pdiffusion 892 -1614 892 -1614 0 feedthrough
rlabel pdiffusion 899 -1614 899 -1614 0 feedthrough
rlabel pdiffusion 906 -1614 906 -1614 0 feedthrough
rlabel pdiffusion 913 -1614 913 -1614 0 feedthrough
rlabel pdiffusion 920 -1614 920 -1614 0 feedthrough
rlabel pdiffusion 927 -1614 927 -1614 0 cellNo=532
rlabel pdiffusion 934 -1614 934 -1614 0 feedthrough
rlabel pdiffusion 941 -1614 941 -1614 0 feedthrough
rlabel pdiffusion 948 -1614 948 -1614 0 feedthrough
rlabel pdiffusion 955 -1614 955 -1614 0 feedthrough
rlabel pdiffusion 962 -1614 962 -1614 0 feedthrough
rlabel pdiffusion 969 -1614 969 -1614 0 feedthrough
rlabel pdiffusion 976 -1614 976 -1614 0 feedthrough
rlabel pdiffusion 983 -1614 983 -1614 0 feedthrough
rlabel pdiffusion 990 -1614 990 -1614 0 feedthrough
rlabel pdiffusion 997 -1614 997 -1614 0 feedthrough
rlabel pdiffusion 1004 -1614 1004 -1614 0 feedthrough
rlabel pdiffusion 1011 -1614 1011 -1614 0 feedthrough
rlabel pdiffusion 1018 -1614 1018 -1614 0 cellNo=298
rlabel pdiffusion 1025 -1614 1025 -1614 0 feedthrough
rlabel pdiffusion 1032 -1614 1032 -1614 0 feedthrough
rlabel pdiffusion 1039 -1614 1039 -1614 0 feedthrough
rlabel pdiffusion 1046 -1614 1046 -1614 0 cellNo=833
rlabel pdiffusion 1053 -1614 1053 -1614 0 feedthrough
rlabel pdiffusion 1060 -1614 1060 -1614 0 cellNo=779
rlabel pdiffusion 1067 -1614 1067 -1614 0 feedthrough
rlabel pdiffusion 1074 -1614 1074 -1614 0 feedthrough
rlabel pdiffusion 1081 -1614 1081 -1614 0 feedthrough
rlabel pdiffusion 1088 -1614 1088 -1614 0 feedthrough
rlabel pdiffusion 1095 -1614 1095 -1614 0 feedthrough
rlabel pdiffusion 1102 -1614 1102 -1614 0 cellNo=292
rlabel pdiffusion 1109 -1614 1109 -1614 0 feedthrough
rlabel pdiffusion 1116 -1614 1116 -1614 0 cellNo=280
rlabel pdiffusion 1123 -1614 1123 -1614 0 feedthrough
rlabel pdiffusion 1130 -1614 1130 -1614 0 feedthrough
rlabel pdiffusion 1137 -1614 1137 -1614 0 feedthrough
rlabel pdiffusion 1144 -1614 1144 -1614 0 feedthrough
rlabel pdiffusion 1151 -1614 1151 -1614 0 cellNo=255
rlabel pdiffusion 1158 -1614 1158 -1614 0 feedthrough
rlabel pdiffusion 1165 -1614 1165 -1614 0 feedthrough
rlabel pdiffusion 1172 -1614 1172 -1614 0 feedthrough
rlabel pdiffusion 1179 -1614 1179 -1614 0 feedthrough
rlabel pdiffusion 1186 -1614 1186 -1614 0 feedthrough
rlabel pdiffusion 1193 -1614 1193 -1614 0 feedthrough
rlabel pdiffusion 1200 -1614 1200 -1614 0 feedthrough
rlabel pdiffusion 1207 -1614 1207 -1614 0 feedthrough
rlabel pdiffusion 1214 -1614 1214 -1614 0 feedthrough
rlabel pdiffusion 1221 -1614 1221 -1614 0 feedthrough
rlabel pdiffusion 1228 -1614 1228 -1614 0 feedthrough
rlabel pdiffusion 1235 -1614 1235 -1614 0 feedthrough
rlabel pdiffusion 1242 -1614 1242 -1614 0 feedthrough
rlabel pdiffusion 1249 -1614 1249 -1614 0 feedthrough
rlabel pdiffusion 1256 -1614 1256 -1614 0 cellNo=302
rlabel pdiffusion 1263 -1614 1263 -1614 0 feedthrough
rlabel pdiffusion 1270 -1614 1270 -1614 0 feedthrough
rlabel pdiffusion 1277 -1614 1277 -1614 0 feedthrough
rlabel pdiffusion 1284 -1614 1284 -1614 0 feedthrough
rlabel pdiffusion 1291 -1614 1291 -1614 0 feedthrough
rlabel pdiffusion 1298 -1614 1298 -1614 0 feedthrough
rlabel pdiffusion 1305 -1614 1305 -1614 0 feedthrough
rlabel pdiffusion 1312 -1614 1312 -1614 0 feedthrough
rlabel pdiffusion 1319 -1614 1319 -1614 0 feedthrough
rlabel pdiffusion 1326 -1614 1326 -1614 0 feedthrough
rlabel pdiffusion 1333 -1614 1333 -1614 0 feedthrough
rlabel pdiffusion 1340 -1614 1340 -1614 0 feedthrough
rlabel pdiffusion 1347 -1614 1347 -1614 0 feedthrough
rlabel pdiffusion 1354 -1614 1354 -1614 0 feedthrough
rlabel pdiffusion 1361 -1614 1361 -1614 0 feedthrough
rlabel pdiffusion 1368 -1614 1368 -1614 0 feedthrough
rlabel pdiffusion 1375 -1614 1375 -1614 0 feedthrough
rlabel pdiffusion 1382 -1614 1382 -1614 0 feedthrough
rlabel pdiffusion 1389 -1614 1389 -1614 0 feedthrough
rlabel pdiffusion 1396 -1614 1396 -1614 0 feedthrough
rlabel pdiffusion 1403 -1614 1403 -1614 0 feedthrough
rlabel pdiffusion 1410 -1614 1410 -1614 0 feedthrough
rlabel pdiffusion 1417 -1614 1417 -1614 0 feedthrough
rlabel pdiffusion 1424 -1614 1424 -1614 0 feedthrough
rlabel pdiffusion 1431 -1614 1431 -1614 0 feedthrough
rlabel pdiffusion 1438 -1614 1438 -1614 0 feedthrough
rlabel pdiffusion 1445 -1614 1445 -1614 0 feedthrough
rlabel pdiffusion 1452 -1614 1452 -1614 0 feedthrough
rlabel pdiffusion 1459 -1614 1459 -1614 0 feedthrough
rlabel pdiffusion 1466 -1614 1466 -1614 0 feedthrough
rlabel pdiffusion 1473 -1614 1473 -1614 0 feedthrough
rlabel pdiffusion 1480 -1614 1480 -1614 0 feedthrough
rlabel pdiffusion 1487 -1614 1487 -1614 0 feedthrough
rlabel pdiffusion 1494 -1614 1494 -1614 0 feedthrough
rlabel pdiffusion 1501 -1614 1501 -1614 0 feedthrough
rlabel pdiffusion 1508 -1614 1508 -1614 0 feedthrough
rlabel pdiffusion 1515 -1614 1515 -1614 0 feedthrough
rlabel pdiffusion 1522 -1614 1522 -1614 0 feedthrough
rlabel pdiffusion 1529 -1614 1529 -1614 0 feedthrough
rlabel pdiffusion 1536 -1614 1536 -1614 0 feedthrough
rlabel pdiffusion 1543 -1614 1543 -1614 0 feedthrough
rlabel pdiffusion 1550 -1614 1550 -1614 0 feedthrough
rlabel pdiffusion 1557 -1614 1557 -1614 0 feedthrough
rlabel pdiffusion 1564 -1614 1564 -1614 0 feedthrough
rlabel pdiffusion 1571 -1614 1571 -1614 0 feedthrough
rlabel pdiffusion 1578 -1614 1578 -1614 0 feedthrough
rlabel pdiffusion 1585 -1614 1585 -1614 0 feedthrough
rlabel pdiffusion 1592 -1614 1592 -1614 0 feedthrough
rlabel pdiffusion 1599 -1614 1599 -1614 0 feedthrough
rlabel pdiffusion 1606 -1614 1606 -1614 0 feedthrough
rlabel pdiffusion 1613 -1614 1613 -1614 0 feedthrough
rlabel pdiffusion 1620 -1614 1620 -1614 0 feedthrough
rlabel pdiffusion 1627 -1614 1627 -1614 0 feedthrough
rlabel pdiffusion 1634 -1614 1634 -1614 0 feedthrough
rlabel pdiffusion 1641 -1614 1641 -1614 0 feedthrough
rlabel pdiffusion 1648 -1614 1648 -1614 0 feedthrough
rlabel pdiffusion 1655 -1614 1655 -1614 0 feedthrough
rlabel pdiffusion 1662 -1614 1662 -1614 0 feedthrough
rlabel pdiffusion 1669 -1614 1669 -1614 0 feedthrough
rlabel pdiffusion 1676 -1614 1676 -1614 0 feedthrough
rlabel pdiffusion 1683 -1614 1683 -1614 0 feedthrough
rlabel pdiffusion 1690 -1614 1690 -1614 0 feedthrough
rlabel pdiffusion 1697 -1614 1697 -1614 0 feedthrough
rlabel pdiffusion 1704 -1614 1704 -1614 0 cellNo=165
rlabel pdiffusion 1711 -1614 1711 -1614 0 cellNo=520
rlabel pdiffusion 1718 -1614 1718 -1614 0 feedthrough
rlabel pdiffusion 1753 -1614 1753 -1614 0 feedthrough
rlabel pdiffusion 3 -1741 3 -1741 0 cellNo=1024
rlabel pdiffusion 10 -1741 10 -1741 0 cellNo=1331
rlabel pdiffusion 17 -1741 17 -1741 0 cellNo=848
rlabel pdiffusion 24 -1741 24 -1741 0 cellNo=1113
rlabel pdiffusion 31 -1741 31 -1741 0 cellNo=1025
rlabel pdiffusion 38 -1741 38 -1741 0 feedthrough
rlabel pdiffusion 45 -1741 45 -1741 0 feedthrough
rlabel pdiffusion 52 -1741 52 -1741 0 feedthrough
rlabel pdiffusion 59 -1741 59 -1741 0 cellNo=208
rlabel pdiffusion 66 -1741 66 -1741 0 feedthrough
rlabel pdiffusion 73 -1741 73 -1741 0 feedthrough
rlabel pdiffusion 80 -1741 80 -1741 0 feedthrough
rlabel pdiffusion 87 -1741 87 -1741 0 feedthrough
rlabel pdiffusion 94 -1741 94 -1741 0 feedthrough
rlabel pdiffusion 101 -1741 101 -1741 0 feedthrough
rlabel pdiffusion 108 -1741 108 -1741 0 feedthrough
rlabel pdiffusion 115 -1741 115 -1741 0 feedthrough
rlabel pdiffusion 122 -1741 122 -1741 0 feedthrough
rlabel pdiffusion 129 -1741 129 -1741 0 feedthrough
rlabel pdiffusion 136 -1741 136 -1741 0 feedthrough
rlabel pdiffusion 143 -1741 143 -1741 0 feedthrough
rlabel pdiffusion 150 -1741 150 -1741 0 feedthrough
rlabel pdiffusion 157 -1741 157 -1741 0 cellNo=401
rlabel pdiffusion 164 -1741 164 -1741 0 feedthrough
rlabel pdiffusion 171 -1741 171 -1741 0 cellNo=382
rlabel pdiffusion 178 -1741 178 -1741 0 cellNo=13
rlabel pdiffusion 185 -1741 185 -1741 0 feedthrough
rlabel pdiffusion 192 -1741 192 -1741 0 cellNo=811
rlabel pdiffusion 199 -1741 199 -1741 0 feedthrough
rlabel pdiffusion 206 -1741 206 -1741 0 feedthrough
rlabel pdiffusion 213 -1741 213 -1741 0 feedthrough
rlabel pdiffusion 220 -1741 220 -1741 0 feedthrough
rlabel pdiffusion 227 -1741 227 -1741 0 feedthrough
rlabel pdiffusion 234 -1741 234 -1741 0 feedthrough
rlabel pdiffusion 241 -1741 241 -1741 0 feedthrough
rlabel pdiffusion 248 -1741 248 -1741 0 feedthrough
rlabel pdiffusion 255 -1741 255 -1741 0 cellNo=810
rlabel pdiffusion 262 -1741 262 -1741 0 cellNo=253
rlabel pdiffusion 269 -1741 269 -1741 0 feedthrough
rlabel pdiffusion 276 -1741 276 -1741 0 cellNo=898
rlabel pdiffusion 283 -1741 283 -1741 0 feedthrough
rlabel pdiffusion 290 -1741 290 -1741 0 feedthrough
rlabel pdiffusion 297 -1741 297 -1741 0 feedthrough
rlabel pdiffusion 304 -1741 304 -1741 0 feedthrough
rlabel pdiffusion 311 -1741 311 -1741 0 feedthrough
rlabel pdiffusion 318 -1741 318 -1741 0 feedthrough
rlabel pdiffusion 325 -1741 325 -1741 0 feedthrough
rlabel pdiffusion 332 -1741 332 -1741 0 feedthrough
rlabel pdiffusion 339 -1741 339 -1741 0 feedthrough
rlabel pdiffusion 346 -1741 346 -1741 0 cellNo=727
rlabel pdiffusion 353 -1741 353 -1741 0 feedthrough
rlabel pdiffusion 360 -1741 360 -1741 0 feedthrough
rlabel pdiffusion 367 -1741 367 -1741 0 feedthrough
rlabel pdiffusion 374 -1741 374 -1741 0 feedthrough
rlabel pdiffusion 381 -1741 381 -1741 0 feedthrough
rlabel pdiffusion 388 -1741 388 -1741 0 feedthrough
rlabel pdiffusion 395 -1741 395 -1741 0 feedthrough
rlabel pdiffusion 402 -1741 402 -1741 0 feedthrough
rlabel pdiffusion 409 -1741 409 -1741 0 cellNo=670
rlabel pdiffusion 416 -1741 416 -1741 0 feedthrough
rlabel pdiffusion 423 -1741 423 -1741 0 feedthrough
rlabel pdiffusion 430 -1741 430 -1741 0 cellNo=711
rlabel pdiffusion 437 -1741 437 -1741 0 feedthrough
rlabel pdiffusion 444 -1741 444 -1741 0 feedthrough
rlabel pdiffusion 451 -1741 451 -1741 0 feedthrough
rlabel pdiffusion 458 -1741 458 -1741 0 feedthrough
rlabel pdiffusion 465 -1741 465 -1741 0 feedthrough
rlabel pdiffusion 472 -1741 472 -1741 0 feedthrough
rlabel pdiffusion 479 -1741 479 -1741 0 cellNo=722
rlabel pdiffusion 486 -1741 486 -1741 0 feedthrough
rlabel pdiffusion 493 -1741 493 -1741 0 feedthrough
rlabel pdiffusion 500 -1741 500 -1741 0 feedthrough
rlabel pdiffusion 507 -1741 507 -1741 0 feedthrough
rlabel pdiffusion 514 -1741 514 -1741 0 feedthrough
rlabel pdiffusion 521 -1741 521 -1741 0 feedthrough
rlabel pdiffusion 528 -1741 528 -1741 0 cellNo=299
rlabel pdiffusion 535 -1741 535 -1741 0 feedthrough
rlabel pdiffusion 542 -1741 542 -1741 0 cellNo=549
rlabel pdiffusion 549 -1741 549 -1741 0 feedthrough
rlabel pdiffusion 556 -1741 556 -1741 0 feedthrough
rlabel pdiffusion 563 -1741 563 -1741 0 feedthrough
rlabel pdiffusion 570 -1741 570 -1741 0 feedthrough
rlabel pdiffusion 577 -1741 577 -1741 0 feedthrough
rlabel pdiffusion 584 -1741 584 -1741 0 feedthrough
rlabel pdiffusion 591 -1741 591 -1741 0 feedthrough
rlabel pdiffusion 598 -1741 598 -1741 0 feedthrough
rlabel pdiffusion 605 -1741 605 -1741 0 feedthrough
rlabel pdiffusion 612 -1741 612 -1741 0 feedthrough
rlabel pdiffusion 619 -1741 619 -1741 0 feedthrough
rlabel pdiffusion 626 -1741 626 -1741 0 feedthrough
rlabel pdiffusion 633 -1741 633 -1741 0 feedthrough
rlabel pdiffusion 640 -1741 640 -1741 0 feedthrough
rlabel pdiffusion 647 -1741 647 -1741 0 feedthrough
rlabel pdiffusion 654 -1741 654 -1741 0 feedthrough
rlabel pdiffusion 661 -1741 661 -1741 0 feedthrough
rlabel pdiffusion 668 -1741 668 -1741 0 feedthrough
rlabel pdiffusion 675 -1741 675 -1741 0 cellNo=987
rlabel pdiffusion 682 -1741 682 -1741 0 feedthrough
rlabel pdiffusion 689 -1741 689 -1741 0 cellNo=124
rlabel pdiffusion 696 -1741 696 -1741 0 feedthrough
rlabel pdiffusion 703 -1741 703 -1741 0 cellNo=970
rlabel pdiffusion 710 -1741 710 -1741 0 feedthrough
rlabel pdiffusion 717 -1741 717 -1741 0 feedthrough
rlabel pdiffusion 724 -1741 724 -1741 0 cellNo=577
rlabel pdiffusion 731 -1741 731 -1741 0 cellNo=983
rlabel pdiffusion 738 -1741 738 -1741 0 cellNo=777
rlabel pdiffusion 745 -1741 745 -1741 0 feedthrough
rlabel pdiffusion 752 -1741 752 -1741 0 feedthrough
rlabel pdiffusion 759 -1741 759 -1741 0 feedthrough
rlabel pdiffusion 766 -1741 766 -1741 0 feedthrough
rlabel pdiffusion 773 -1741 773 -1741 0 feedthrough
rlabel pdiffusion 780 -1741 780 -1741 0 cellNo=649
rlabel pdiffusion 787 -1741 787 -1741 0 cellNo=937
rlabel pdiffusion 794 -1741 794 -1741 0 feedthrough
rlabel pdiffusion 801 -1741 801 -1741 0 cellNo=426
rlabel pdiffusion 808 -1741 808 -1741 0 cellNo=104
rlabel pdiffusion 815 -1741 815 -1741 0 feedthrough
rlabel pdiffusion 822 -1741 822 -1741 0 feedthrough
rlabel pdiffusion 829 -1741 829 -1741 0 cellNo=239
rlabel pdiffusion 836 -1741 836 -1741 0 feedthrough
rlabel pdiffusion 843 -1741 843 -1741 0 feedthrough
rlabel pdiffusion 850 -1741 850 -1741 0 feedthrough
rlabel pdiffusion 857 -1741 857 -1741 0 feedthrough
rlabel pdiffusion 864 -1741 864 -1741 0 feedthrough
rlabel pdiffusion 871 -1741 871 -1741 0 cellNo=614
rlabel pdiffusion 878 -1741 878 -1741 0 feedthrough
rlabel pdiffusion 885 -1741 885 -1741 0 cellNo=190
rlabel pdiffusion 892 -1741 892 -1741 0 cellNo=812
rlabel pdiffusion 899 -1741 899 -1741 0 feedthrough
rlabel pdiffusion 906 -1741 906 -1741 0 feedthrough
rlabel pdiffusion 913 -1741 913 -1741 0 cellNo=244
rlabel pdiffusion 920 -1741 920 -1741 0 cellNo=782
rlabel pdiffusion 927 -1741 927 -1741 0 cellNo=442
rlabel pdiffusion 934 -1741 934 -1741 0 feedthrough
rlabel pdiffusion 941 -1741 941 -1741 0 feedthrough
rlabel pdiffusion 948 -1741 948 -1741 0 feedthrough
rlabel pdiffusion 955 -1741 955 -1741 0 feedthrough
rlabel pdiffusion 962 -1741 962 -1741 0 feedthrough
rlabel pdiffusion 969 -1741 969 -1741 0 feedthrough
rlabel pdiffusion 976 -1741 976 -1741 0 cellNo=451
rlabel pdiffusion 983 -1741 983 -1741 0 feedthrough
rlabel pdiffusion 990 -1741 990 -1741 0 cellNo=521
rlabel pdiffusion 997 -1741 997 -1741 0 feedthrough
rlabel pdiffusion 1004 -1741 1004 -1741 0 feedthrough
rlabel pdiffusion 1011 -1741 1011 -1741 0 feedthrough
rlabel pdiffusion 1018 -1741 1018 -1741 0 feedthrough
rlabel pdiffusion 1025 -1741 1025 -1741 0 feedthrough
rlabel pdiffusion 1032 -1741 1032 -1741 0 feedthrough
rlabel pdiffusion 1039 -1741 1039 -1741 0 feedthrough
rlabel pdiffusion 1046 -1741 1046 -1741 0 feedthrough
rlabel pdiffusion 1053 -1741 1053 -1741 0 feedthrough
rlabel pdiffusion 1060 -1741 1060 -1741 0 feedthrough
rlabel pdiffusion 1067 -1741 1067 -1741 0 cellNo=453
rlabel pdiffusion 1074 -1741 1074 -1741 0 feedthrough
rlabel pdiffusion 1081 -1741 1081 -1741 0 feedthrough
rlabel pdiffusion 1088 -1741 1088 -1741 0 feedthrough
rlabel pdiffusion 1095 -1741 1095 -1741 0 feedthrough
rlabel pdiffusion 1102 -1741 1102 -1741 0 feedthrough
rlabel pdiffusion 1109 -1741 1109 -1741 0 feedthrough
rlabel pdiffusion 1116 -1741 1116 -1741 0 cellNo=630
rlabel pdiffusion 1123 -1741 1123 -1741 0 feedthrough
rlabel pdiffusion 1130 -1741 1130 -1741 0 feedthrough
rlabel pdiffusion 1137 -1741 1137 -1741 0 feedthrough
rlabel pdiffusion 1144 -1741 1144 -1741 0 feedthrough
rlabel pdiffusion 1151 -1741 1151 -1741 0 feedthrough
rlabel pdiffusion 1158 -1741 1158 -1741 0 feedthrough
rlabel pdiffusion 1165 -1741 1165 -1741 0 feedthrough
rlabel pdiffusion 1172 -1741 1172 -1741 0 feedthrough
rlabel pdiffusion 1179 -1741 1179 -1741 0 feedthrough
rlabel pdiffusion 1186 -1741 1186 -1741 0 feedthrough
rlabel pdiffusion 1193 -1741 1193 -1741 0 feedthrough
rlabel pdiffusion 1200 -1741 1200 -1741 0 feedthrough
rlabel pdiffusion 1207 -1741 1207 -1741 0 feedthrough
rlabel pdiffusion 1214 -1741 1214 -1741 0 feedthrough
rlabel pdiffusion 1221 -1741 1221 -1741 0 feedthrough
rlabel pdiffusion 1228 -1741 1228 -1741 0 feedthrough
rlabel pdiffusion 1235 -1741 1235 -1741 0 feedthrough
rlabel pdiffusion 1242 -1741 1242 -1741 0 feedthrough
rlabel pdiffusion 1249 -1741 1249 -1741 0 cellNo=742
rlabel pdiffusion 1256 -1741 1256 -1741 0 feedthrough
rlabel pdiffusion 1263 -1741 1263 -1741 0 feedthrough
rlabel pdiffusion 1270 -1741 1270 -1741 0 feedthrough
rlabel pdiffusion 1277 -1741 1277 -1741 0 feedthrough
rlabel pdiffusion 1284 -1741 1284 -1741 0 feedthrough
rlabel pdiffusion 1291 -1741 1291 -1741 0 feedthrough
rlabel pdiffusion 1298 -1741 1298 -1741 0 feedthrough
rlabel pdiffusion 1305 -1741 1305 -1741 0 feedthrough
rlabel pdiffusion 1312 -1741 1312 -1741 0 feedthrough
rlabel pdiffusion 1319 -1741 1319 -1741 0 feedthrough
rlabel pdiffusion 1326 -1741 1326 -1741 0 feedthrough
rlabel pdiffusion 1333 -1741 1333 -1741 0 feedthrough
rlabel pdiffusion 1340 -1741 1340 -1741 0 feedthrough
rlabel pdiffusion 1347 -1741 1347 -1741 0 feedthrough
rlabel pdiffusion 1354 -1741 1354 -1741 0 feedthrough
rlabel pdiffusion 1361 -1741 1361 -1741 0 feedthrough
rlabel pdiffusion 1368 -1741 1368 -1741 0 feedthrough
rlabel pdiffusion 1375 -1741 1375 -1741 0 feedthrough
rlabel pdiffusion 1382 -1741 1382 -1741 0 feedthrough
rlabel pdiffusion 1389 -1741 1389 -1741 0 feedthrough
rlabel pdiffusion 1396 -1741 1396 -1741 0 feedthrough
rlabel pdiffusion 1403 -1741 1403 -1741 0 feedthrough
rlabel pdiffusion 1410 -1741 1410 -1741 0 feedthrough
rlabel pdiffusion 1417 -1741 1417 -1741 0 feedthrough
rlabel pdiffusion 1424 -1741 1424 -1741 0 feedthrough
rlabel pdiffusion 1431 -1741 1431 -1741 0 feedthrough
rlabel pdiffusion 1438 -1741 1438 -1741 0 feedthrough
rlabel pdiffusion 1445 -1741 1445 -1741 0 feedthrough
rlabel pdiffusion 1452 -1741 1452 -1741 0 feedthrough
rlabel pdiffusion 1459 -1741 1459 -1741 0 feedthrough
rlabel pdiffusion 1466 -1741 1466 -1741 0 feedthrough
rlabel pdiffusion 1473 -1741 1473 -1741 0 feedthrough
rlabel pdiffusion 1480 -1741 1480 -1741 0 feedthrough
rlabel pdiffusion 1487 -1741 1487 -1741 0 feedthrough
rlabel pdiffusion 1494 -1741 1494 -1741 0 feedthrough
rlabel pdiffusion 1501 -1741 1501 -1741 0 feedthrough
rlabel pdiffusion 1508 -1741 1508 -1741 0 feedthrough
rlabel pdiffusion 1515 -1741 1515 -1741 0 feedthrough
rlabel pdiffusion 1522 -1741 1522 -1741 0 feedthrough
rlabel pdiffusion 1529 -1741 1529 -1741 0 feedthrough
rlabel pdiffusion 1536 -1741 1536 -1741 0 feedthrough
rlabel pdiffusion 1543 -1741 1543 -1741 0 feedthrough
rlabel pdiffusion 1550 -1741 1550 -1741 0 feedthrough
rlabel pdiffusion 1557 -1741 1557 -1741 0 feedthrough
rlabel pdiffusion 1564 -1741 1564 -1741 0 feedthrough
rlabel pdiffusion 1571 -1741 1571 -1741 0 feedthrough
rlabel pdiffusion 1578 -1741 1578 -1741 0 feedthrough
rlabel pdiffusion 1585 -1741 1585 -1741 0 feedthrough
rlabel pdiffusion 1592 -1741 1592 -1741 0 feedthrough
rlabel pdiffusion 1599 -1741 1599 -1741 0 feedthrough
rlabel pdiffusion 1606 -1741 1606 -1741 0 feedthrough
rlabel pdiffusion 1613 -1741 1613 -1741 0 feedthrough
rlabel pdiffusion 1620 -1741 1620 -1741 0 feedthrough
rlabel pdiffusion 1627 -1741 1627 -1741 0 feedthrough
rlabel pdiffusion 1634 -1741 1634 -1741 0 feedthrough
rlabel pdiffusion 1641 -1741 1641 -1741 0 feedthrough
rlabel pdiffusion 1648 -1741 1648 -1741 0 feedthrough
rlabel pdiffusion 1655 -1741 1655 -1741 0 feedthrough
rlabel pdiffusion 1662 -1741 1662 -1741 0 feedthrough
rlabel pdiffusion 1669 -1741 1669 -1741 0 feedthrough
rlabel pdiffusion 1676 -1741 1676 -1741 0 feedthrough
rlabel pdiffusion 1683 -1741 1683 -1741 0 feedthrough
rlabel pdiffusion 1690 -1741 1690 -1741 0 feedthrough
rlabel pdiffusion 1697 -1741 1697 -1741 0 feedthrough
rlabel pdiffusion 1704 -1741 1704 -1741 0 feedthrough
rlabel pdiffusion 1711 -1741 1711 -1741 0 feedthrough
rlabel pdiffusion 1718 -1741 1718 -1741 0 feedthrough
rlabel pdiffusion 1725 -1741 1725 -1741 0 feedthrough
rlabel pdiffusion 1732 -1741 1732 -1741 0 feedthrough
rlabel pdiffusion 1739 -1741 1739 -1741 0 feedthrough
rlabel pdiffusion 1746 -1741 1746 -1741 0 cellNo=885
rlabel pdiffusion 1753 -1741 1753 -1741 0 feedthrough
rlabel pdiffusion 1760 -1741 1760 -1741 0 feedthrough
rlabel pdiffusion 1767 -1741 1767 -1741 0 feedthrough
rlabel pdiffusion 1774 -1741 1774 -1741 0 feedthrough
rlabel pdiffusion 1781 -1741 1781 -1741 0 feedthrough
rlabel pdiffusion 3 -1888 3 -1888 0 cellNo=1027
rlabel pdiffusion 10 -1888 10 -1888 0 cellNo=1167
rlabel pdiffusion 17 -1888 17 -1888 0 cellNo=1362
rlabel pdiffusion 24 -1888 24 -1888 0 cellNo=1201
rlabel pdiffusion 31 -1888 31 -1888 0 feedthrough
rlabel pdiffusion 38 -1888 38 -1888 0 feedthrough
rlabel pdiffusion 45 -1888 45 -1888 0 feedthrough
rlabel pdiffusion 52 -1888 52 -1888 0 feedthrough
rlabel pdiffusion 59 -1888 59 -1888 0 feedthrough
rlabel pdiffusion 66 -1888 66 -1888 0 feedthrough
rlabel pdiffusion 73 -1888 73 -1888 0 feedthrough
rlabel pdiffusion 80 -1888 80 -1888 0 feedthrough
rlabel pdiffusion 87 -1888 87 -1888 0 feedthrough
rlabel pdiffusion 94 -1888 94 -1888 0 feedthrough
rlabel pdiffusion 101 -1888 101 -1888 0 feedthrough
rlabel pdiffusion 108 -1888 108 -1888 0 cellNo=123
rlabel pdiffusion 115 -1888 115 -1888 0 feedthrough
rlabel pdiffusion 122 -1888 122 -1888 0 feedthrough
rlabel pdiffusion 129 -1888 129 -1888 0 feedthrough
rlabel pdiffusion 136 -1888 136 -1888 0 feedthrough
rlabel pdiffusion 143 -1888 143 -1888 0 feedthrough
rlabel pdiffusion 150 -1888 150 -1888 0 feedthrough
rlabel pdiffusion 157 -1888 157 -1888 0 cellNo=290
rlabel pdiffusion 164 -1888 164 -1888 0 feedthrough
rlabel pdiffusion 171 -1888 171 -1888 0 feedthrough
rlabel pdiffusion 178 -1888 178 -1888 0 cellNo=379
rlabel pdiffusion 185 -1888 185 -1888 0 feedthrough
rlabel pdiffusion 192 -1888 192 -1888 0 cellNo=291
rlabel pdiffusion 199 -1888 199 -1888 0 feedthrough
rlabel pdiffusion 206 -1888 206 -1888 0 cellNo=598
rlabel pdiffusion 213 -1888 213 -1888 0 feedthrough
rlabel pdiffusion 220 -1888 220 -1888 0 feedthrough
rlabel pdiffusion 227 -1888 227 -1888 0 feedthrough
rlabel pdiffusion 234 -1888 234 -1888 0 feedthrough
rlabel pdiffusion 241 -1888 241 -1888 0 feedthrough
rlabel pdiffusion 248 -1888 248 -1888 0 cellNo=989
rlabel pdiffusion 255 -1888 255 -1888 0 feedthrough
rlabel pdiffusion 262 -1888 262 -1888 0 cellNo=387
rlabel pdiffusion 269 -1888 269 -1888 0 feedthrough
rlabel pdiffusion 276 -1888 276 -1888 0 feedthrough
rlabel pdiffusion 283 -1888 283 -1888 0 feedthrough
rlabel pdiffusion 290 -1888 290 -1888 0 feedthrough
rlabel pdiffusion 297 -1888 297 -1888 0 feedthrough
rlabel pdiffusion 304 -1888 304 -1888 0 feedthrough
rlabel pdiffusion 311 -1888 311 -1888 0 feedthrough
rlabel pdiffusion 318 -1888 318 -1888 0 feedthrough
rlabel pdiffusion 325 -1888 325 -1888 0 feedthrough
rlabel pdiffusion 332 -1888 332 -1888 0 feedthrough
rlabel pdiffusion 339 -1888 339 -1888 0 cellNo=842
rlabel pdiffusion 346 -1888 346 -1888 0 feedthrough
rlabel pdiffusion 353 -1888 353 -1888 0 feedthrough
rlabel pdiffusion 360 -1888 360 -1888 0 feedthrough
rlabel pdiffusion 367 -1888 367 -1888 0 feedthrough
rlabel pdiffusion 374 -1888 374 -1888 0 feedthrough
rlabel pdiffusion 381 -1888 381 -1888 0 feedthrough
rlabel pdiffusion 388 -1888 388 -1888 0 feedthrough
rlabel pdiffusion 395 -1888 395 -1888 0 feedthrough
rlabel pdiffusion 402 -1888 402 -1888 0 feedthrough
rlabel pdiffusion 409 -1888 409 -1888 0 feedthrough
rlabel pdiffusion 416 -1888 416 -1888 0 feedthrough
rlabel pdiffusion 423 -1888 423 -1888 0 feedthrough
rlabel pdiffusion 430 -1888 430 -1888 0 feedthrough
rlabel pdiffusion 437 -1888 437 -1888 0 feedthrough
rlabel pdiffusion 444 -1888 444 -1888 0 cellNo=917
rlabel pdiffusion 451 -1888 451 -1888 0 feedthrough
rlabel pdiffusion 458 -1888 458 -1888 0 feedthrough
rlabel pdiffusion 465 -1888 465 -1888 0 cellNo=580
rlabel pdiffusion 472 -1888 472 -1888 0 cellNo=754
rlabel pdiffusion 479 -1888 479 -1888 0 feedthrough
rlabel pdiffusion 486 -1888 486 -1888 0 feedthrough
rlabel pdiffusion 493 -1888 493 -1888 0 feedthrough
rlabel pdiffusion 500 -1888 500 -1888 0 cellNo=28
rlabel pdiffusion 507 -1888 507 -1888 0 feedthrough
rlabel pdiffusion 514 -1888 514 -1888 0 feedthrough
rlabel pdiffusion 521 -1888 521 -1888 0 feedthrough
rlabel pdiffusion 528 -1888 528 -1888 0 cellNo=831
rlabel pdiffusion 535 -1888 535 -1888 0 feedthrough
rlabel pdiffusion 542 -1888 542 -1888 0 feedthrough
rlabel pdiffusion 549 -1888 549 -1888 0 feedthrough
rlabel pdiffusion 556 -1888 556 -1888 0 feedthrough
rlabel pdiffusion 563 -1888 563 -1888 0 feedthrough
rlabel pdiffusion 570 -1888 570 -1888 0 cellNo=744
rlabel pdiffusion 577 -1888 577 -1888 0 feedthrough
rlabel pdiffusion 584 -1888 584 -1888 0 feedthrough
rlabel pdiffusion 591 -1888 591 -1888 0 feedthrough
rlabel pdiffusion 598 -1888 598 -1888 0 feedthrough
rlabel pdiffusion 605 -1888 605 -1888 0 feedthrough
rlabel pdiffusion 612 -1888 612 -1888 0 feedthrough
rlabel pdiffusion 619 -1888 619 -1888 0 feedthrough
rlabel pdiffusion 626 -1888 626 -1888 0 feedthrough
rlabel pdiffusion 633 -1888 633 -1888 0 feedthrough
rlabel pdiffusion 640 -1888 640 -1888 0 feedthrough
rlabel pdiffusion 647 -1888 647 -1888 0 cellNo=61
rlabel pdiffusion 654 -1888 654 -1888 0 cellNo=958
rlabel pdiffusion 661 -1888 661 -1888 0 feedthrough
rlabel pdiffusion 668 -1888 668 -1888 0 feedthrough
rlabel pdiffusion 675 -1888 675 -1888 0 feedthrough
rlabel pdiffusion 682 -1888 682 -1888 0 feedthrough
rlabel pdiffusion 689 -1888 689 -1888 0 feedthrough
rlabel pdiffusion 696 -1888 696 -1888 0 feedthrough
rlabel pdiffusion 703 -1888 703 -1888 0 feedthrough
rlabel pdiffusion 710 -1888 710 -1888 0 feedthrough
rlabel pdiffusion 717 -1888 717 -1888 0 feedthrough
rlabel pdiffusion 724 -1888 724 -1888 0 feedthrough
rlabel pdiffusion 731 -1888 731 -1888 0 feedthrough
rlabel pdiffusion 738 -1888 738 -1888 0 feedthrough
rlabel pdiffusion 745 -1888 745 -1888 0 feedthrough
rlabel pdiffusion 752 -1888 752 -1888 0 feedthrough
rlabel pdiffusion 759 -1888 759 -1888 0 feedthrough
rlabel pdiffusion 766 -1888 766 -1888 0 feedthrough
rlabel pdiffusion 773 -1888 773 -1888 0 feedthrough
rlabel pdiffusion 780 -1888 780 -1888 0 feedthrough
rlabel pdiffusion 787 -1888 787 -1888 0 feedthrough
rlabel pdiffusion 794 -1888 794 -1888 0 feedthrough
rlabel pdiffusion 801 -1888 801 -1888 0 cellNo=369
rlabel pdiffusion 808 -1888 808 -1888 0 cellNo=222
rlabel pdiffusion 815 -1888 815 -1888 0 feedthrough
rlabel pdiffusion 822 -1888 822 -1888 0 cellNo=49
rlabel pdiffusion 829 -1888 829 -1888 0 cellNo=212
rlabel pdiffusion 836 -1888 836 -1888 0 cellNo=663
rlabel pdiffusion 843 -1888 843 -1888 0 feedthrough
rlabel pdiffusion 850 -1888 850 -1888 0 feedthrough
rlabel pdiffusion 857 -1888 857 -1888 0 feedthrough
rlabel pdiffusion 864 -1888 864 -1888 0 cellNo=619
rlabel pdiffusion 871 -1888 871 -1888 0 feedthrough
rlabel pdiffusion 878 -1888 878 -1888 0 feedthrough
rlabel pdiffusion 885 -1888 885 -1888 0 feedthrough
rlabel pdiffusion 892 -1888 892 -1888 0 feedthrough
rlabel pdiffusion 899 -1888 899 -1888 0 feedthrough
rlabel pdiffusion 906 -1888 906 -1888 0 cellNo=19
rlabel pdiffusion 913 -1888 913 -1888 0 feedthrough
rlabel pdiffusion 920 -1888 920 -1888 0 feedthrough
rlabel pdiffusion 927 -1888 927 -1888 0 cellNo=351
rlabel pdiffusion 934 -1888 934 -1888 0 cellNo=360
rlabel pdiffusion 941 -1888 941 -1888 0 feedthrough
rlabel pdiffusion 948 -1888 948 -1888 0 feedthrough
rlabel pdiffusion 955 -1888 955 -1888 0 cellNo=449
rlabel pdiffusion 962 -1888 962 -1888 0 feedthrough
rlabel pdiffusion 969 -1888 969 -1888 0 feedthrough
rlabel pdiffusion 976 -1888 976 -1888 0 feedthrough
rlabel pdiffusion 983 -1888 983 -1888 0 cellNo=522
rlabel pdiffusion 990 -1888 990 -1888 0 feedthrough
rlabel pdiffusion 997 -1888 997 -1888 0 feedthrough
rlabel pdiffusion 1004 -1888 1004 -1888 0 feedthrough
rlabel pdiffusion 1011 -1888 1011 -1888 0 feedthrough
rlabel pdiffusion 1018 -1888 1018 -1888 0 cellNo=726
rlabel pdiffusion 1025 -1888 1025 -1888 0 cellNo=106
rlabel pdiffusion 1032 -1888 1032 -1888 0 feedthrough
rlabel pdiffusion 1039 -1888 1039 -1888 0 cellNo=975
rlabel pdiffusion 1046 -1888 1046 -1888 0 cellNo=593
rlabel pdiffusion 1053 -1888 1053 -1888 0 feedthrough
rlabel pdiffusion 1060 -1888 1060 -1888 0 feedthrough
rlabel pdiffusion 1067 -1888 1067 -1888 0 feedthrough
rlabel pdiffusion 1074 -1888 1074 -1888 0 feedthrough
rlabel pdiffusion 1081 -1888 1081 -1888 0 feedthrough
rlabel pdiffusion 1088 -1888 1088 -1888 0 feedthrough
rlabel pdiffusion 1095 -1888 1095 -1888 0 feedthrough
rlabel pdiffusion 1102 -1888 1102 -1888 0 feedthrough
rlabel pdiffusion 1109 -1888 1109 -1888 0 cellNo=669
rlabel pdiffusion 1116 -1888 1116 -1888 0 feedthrough
rlabel pdiffusion 1123 -1888 1123 -1888 0 feedthrough
rlabel pdiffusion 1130 -1888 1130 -1888 0 feedthrough
rlabel pdiffusion 1137 -1888 1137 -1888 0 feedthrough
rlabel pdiffusion 1144 -1888 1144 -1888 0 feedthrough
rlabel pdiffusion 1151 -1888 1151 -1888 0 cellNo=409
rlabel pdiffusion 1158 -1888 1158 -1888 0 cellNo=505
rlabel pdiffusion 1165 -1888 1165 -1888 0 feedthrough
rlabel pdiffusion 1172 -1888 1172 -1888 0 feedthrough
rlabel pdiffusion 1179 -1888 1179 -1888 0 feedthrough
rlabel pdiffusion 1186 -1888 1186 -1888 0 feedthrough
rlabel pdiffusion 1193 -1888 1193 -1888 0 feedthrough
rlabel pdiffusion 1200 -1888 1200 -1888 0 feedthrough
rlabel pdiffusion 1207 -1888 1207 -1888 0 feedthrough
rlabel pdiffusion 1214 -1888 1214 -1888 0 feedthrough
rlabel pdiffusion 1221 -1888 1221 -1888 0 feedthrough
rlabel pdiffusion 1228 -1888 1228 -1888 0 feedthrough
rlabel pdiffusion 1235 -1888 1235 -1888 0 feedthrough
rlabel pdiffusion 1242 -1888 1242 -1888 0 feedthrough
rlabel pdiffusion 1249 -1888 1249 -1888 0 feedthrough
rlabel pdiffusion 1256 -1888 1256 -1888 0 feedthrough
rlabel pdiffusion 1263 -1888 1263 -1888 0 feedthrough
rlabel pdiffusion 1270 -1888 1270 -1888 0 feedthrough
rlabel pdiffusion 1277 -1888 1277 -1888 0 cellNo=748
rlabel pdiffusion 1284 -1888 1284 -1888 0 feedthrough
rlabel pdiffusion 1291 -1888 1291 -1888 0 feedthrough
rlabel pdiffusion 1298 -1888 1298 -1888 0 feedthrough
rlabel pdiffusion 1305 -1888 1305 -1888 0 feedthrough
rlabel pdiffusion 1312 -1888 1312 -1888 0 cellNo=703
rlabel pdiffusion 1319 -1888 1319 -1888 0 feedthrough
rlabel pdiffusion 1326 -1888 1326 -1888 0 feedthrough
rlabel pdiffusion 1333 -1888 1333 -1888 0 feedthrough
rlabel pdiffusion 1340 -1888 1340 -1888 0 feedthrough
rlabel pdiffusion 1347 -1888 1347 -1888 0 feedthrough
rlabel pdiffusion 1354 -1888 1354 -1888 0 feedthrough
rlabel pdiffusion 1361 -1888 1361 -1888 0 feedthrough
rlabel pdiffusion 1368 -1888 1368 -1888 0 feedthrough
rlabel pdiffusion 1375 -1888 1375 -1888 0 feedthrough
rlabel pdiffusion 1382 -1888 1382 -1888 0 feedthrough
rlabel pdiffusion 1389 -1888 1389 -1888 0 feedthrough
rlabel pdiffusion 1396 -1888 1396 -1888 0 feedthrough
rlabel pdiffusion 1403 -1888 1403 -1888 0 feedthrough
rlabel pdiffusion 1410 -1888 1410 -1888 0 feedthrough
rlabel pdiffusion 1417 -1888 1417 -1888 0 feedthrough
rlabel pdiffusion 1424 -1888 1424 -1888 0 feedthrough
rlabel pdiffusion 1431 -1888 1431 -1888 0 feedthrough
rlabel pdiffusion 1438 -1888 1438 -1888 0 feedthrough
rlabel pdiffusion 1445 -1888 1445 -1888 0 feedthrough
rlabel pdiffusion 1452 -1888 1452 -1888 0 feedthrough
rlabel pdiffusion 1459 -1888 1459 -1888 0 feedthrough
rlabel pdiffusion 1466 -1888 1466 -1888 0 feedthrough
rlabel pdiffusion 1473 -1888 1473 -1888 0 feedthrough
rlabel pdiffusion 1480 -1888 1480 -1888 0 feedthrough
rlabel pdiffusion 1487 -1888 1487 -1888 0 feedthrough
rlabel pdiffusion 1494 -1888 1494 -1888 0 feedthrough
rlabel pdiffusion 1501 -1888 1501 -1888 0 feedthrough
rlabel pdiffusion 1508 -1888 1508 -1888 0 feedthrough
rlabel pdiffusion 1515 -1888 1515 -1888 0 feedthrough
rlabel pdiffusion 1522 -1888 1522 -1888 0 feedthrough
rlabel pdiffusion 1529 -1888 1529 -1888 0 feedthrough
rlabel pdiffusion 1536 -1888 1536 -1888 0 feedthrough
rlabel pdiffusion 1543 -1888 1543 -1888 0 feedthrough
rlabel pdiffusion 1550 -1888 1550 -1888 0 feedthrough
rlabel pdiffusion 1557 -1888 1557 -1888 0 feedthrough
rlabel pdiffusion 1564 -1888 1564 -1888 0 feedthrough
rlabel pdiffusion 1571 -1888 1571 -1888 0 feedthrough
rlabel pdiffusion 1578 -1888 1578 -1888 0 feedthrough
rlabel pdiffusion 1585 -1888 1585 -1888 0 feedthrough
rlabel pdiffusion 1592 -1888 1592 -1888 0 feedthrough
rlabel pdiffusion 1599 -1888 1599 -1888 0 feedthrough
rlabel pdiffusion 1606 -1888 1606 -1888 0 feedthrough
rlabel pdiffusion 1613 -1888 1613 -1888 0 feedthrough
rlabel pdiffusion 1620 -1888 1620 -1888 0 feedthrough
rlabel pdiffusion 1627 -1888 1627 -1888 0 feedthrough
rlabel pdiffusion 1634 -1888 1634 -1888 0 feedthrough
rlabel pdiffusion 1641 -1888 1641 -1888 0 feedthrough
rlabel pdiffusion 1648 -1888 1648 -1888 0 feedthrough
rlabel pdiffusion 1655 -1888 1655 -1888 0 feedthrough
rlabel pdiffusion 1662 -1888 1662 -1888 0 feedthrough
rlabel pdiffusion 1669 -1888 1669 -1888 0 feedthrough
rlabel pdiffusion 1676 -1888 1676 -1888 0 feedthrough
rlabel pdiffusion 1683 -1888 1683 -1888 0 feedthrough
rlabel pdiffusion 1690 -1888 1690 -1888 0 feedthrough
rlabel pdiffusion 1697 -1888 1697 -1888 0 feedthrough
rlabel pdiffusion 1704 -1888 1704 -1888 0 feedthrough
rlabel pdiffusion 1711 -1888 1711 -1888 0 feedthrough
rlabel pdiffusion 1718 -1888 1718 -1888 0 feedthrough
rlabel pdiffusion 1725 -1888 1725 -1888 0 feedthrough
rlabel pdiffusion 1732 -1888 1732 -1888 0 feedthrough
rlabel pdiffusion 1739 -1888 1739 -1888 0 feedthrough
rlabel pdiffusion 1746 -1888 1746 -1888 0 feedthrough
rlabel pdiffusion 1753 -1888 1753 -1888 0 feedthrough
rlabel pdiffusion 1760 -1888 1760 -1888 0 feedthrough
rlabel pdiffusion 1767 -1888 1767 -1888 0 feedthrough
rlabel pdiffusion 1774 -1888 1774 -1888 0 cellNo=980
rlabel pdiffusion 1781 -1888 1781 -1888 0 feedthrough
rlabel pdiffusion 1788 -1888 1788 -1888 0 feedthrough
rlabel pdiffusion 1795 -1888 1795 -1888 0 feedthrough
rlabel pdiffusion 1802 -1888 1802 -1888 0 cellNo=791
rlabel pdiffusion 1809 -1888 1809 -1888 0 feedthrough
rlabel pdiffusion 1816 -1888 1816 -1888 0 feedthrough
rlabel pdiffusion 3 -2021 3 -2021 0 cellNo=1028
rlabel pdiffusion 10 -2021 10 -2021 0 cellNo=1161
rlabel pdiffusion 17 -2021 17 -2021 0 cellNo=1244
rlabel pdiffusion 24 -2021 24 -2021 0 cellNo=1032
rlabel pdiffusion 31 -2021 31 -2021 0 feedthrough
rlabel pdiffusion 38 -2021 38 -2021 0 cellNo=1342
rlabel pdiffusion 45 -2021 45 -2021 0 feedthrough
rlabel pdiffusion 52 -2021 52 -2021 0 feedthrough
rlabel pdiffusion 59 -2021 59 -2021 0 feedthrough
rlabel pdiffusion 66 -2021 66 -2021 0 cellNo=95
rlabel pdiffusion 73 -2021 73 -2021 0 feedthrough
rlabel pdiffusion 80 -2021 80 -2021 0 feedthrough
rlabel pdiffusion 87 -2021 87 -2021 0 cellNo=11
rlabel pdiffusion 94 -2021 94 -2021 0 feedthrough
rlabel pdiffusion 101 -2021 101 -2021 0 cellNo=500
rlabel pdiffusion 108 -2021 108 -2021 0 cellNo=303
rlabel pdiffusion 115 -2021 115 -2021 0 feedthrough
rlabel pdiffusion 122 -2021 122 -2021 0 cellNo=471
rlabel pdiffusion 129 -2021 129 -2021 0 cellNo=403
rlabel pdiffusion 136 -2021 136 -2021 0 feedthrough
rlabel pdiffusion 143 -2021 143 -2021 0 cellNo=395
rlabel pdiffusion 150 -2021 150 -2021 0 cellNo=133
rlabel pdiffusion 157 -2021 157 -2021 0 feedthrough
rlabel pdiffusion 164 -2021 164 -2021 0 feedthrough
rlabel pdiffusion 171 -2021 171 -2021 0 feedthrough
rlabel pdiffusion 178 -2021 178 -2021 0 cellNo=814
rlabel pdiffusion 185 -2021 185 -2021 0 feedthrough
rlabel pdiffusion 192 -2021 192 -2021 0 feedthrough
rlabel pdiffusion 199 -2021 199 -2021 0 feedthrough
rlabel pdiffusion 206 -2021 206 -2021 0 feedthrough
rlabel pdiffusion 213 -2021 213 -2021 0 cellNo=249
rlabel pdiffusion 220 -2021 220 -2021 0 cellNo=385
rlabel pdiffusion 227 -2021 227 -2021 0 feedthrough
rlabel pdiffusion 234 -2021 234 -2021 0 feedthrough
rlabel pdiffusion 241 -2021 241 -2021 0 feedthrough
rlabel pdiffusion 248 -2021 248 -2021 0 feedthrough
rlabel pdiffusion 255 -2021 255 -2021 0 feedthrough
rlabel pdiffusion 262 -2021 262 -2021 0 feedthrough
rlabel pdiffusion 269 -2021 269 -2021 0 feedthrough
rlabel pdiffusion 276 -2021 276 -2021 0 feedthrough
rlabel pdiffusion 283 -2021 283 -2021 0 feedthrough
rlabel pdiffusion 290 -2021 290 -2021 0 feedthrough
rlabel pdiffusion 297 -2021 297 -2021 0 feedthrough
rlabel pdiffusion 304 -2021 304 -2021 0 feedthrough
rlabel pdiffusion 311 -2021 311 -2021 0 feedthrough
rlabel pdiffusion 318 -2021 318 -2021 0 feedthrough
rlabel pdiffusion 325 -2021 325 -2021 0 feedthrough
rlabel pdiffusion 332 -2021 332 -2021 0 cellNo=984
rlabel pdiffusion 339 -2021 339 -2021 0 feedthrough
rlabel pdiffusion 346 -2021 346 -2021 0 feedthrough
rlabel pdiffusion 353 -2021 353 -2021 0 feedthrough
rlabel pdiffusion 360 -2021 360 -2021 0 feedthrough
rlabel pdiffusion 367 -2021 367 -2021 0 feedthrough
rlabel pdiffusion 374 -2021 374 -2021 0 feedthrough
rlabel pdiffusion 381 -2021 381 -2021 0 feedthrough
rlabel pdiffusion 388 -2021 388 -2021 0 cellNo=775
rlabel pdiffusion 395 -2021 395 -2021 0 feedthrough
rlabel pdiffusion 402 -2021 402 -2021 0 feedthrough
rlabel pdiffusion 409 -2021 409 -2021 0 feedthrough
rlabel pdiffusion 416 -2021 416 -2021 0 feedthrough
rlabel pdiffusion 423 -2021 423 -2021 0 feedthrough
rlabel pdiffusion 430 -2021 430 -2021 0 feedthrough
rlabel pdiffusion 437 -2021 437 -2021 0 feedthrough
rlabel pdiffusion 444 -2021 444 -2021 0 feedthrough
rlabel pdiffusion 451 -2021 451 -2021 0 feedthrough
rlabel pdiffusion 458 -2021 458 -2021 0 cellNo=139
rlabel pdiffusion 465 -2021 465 -2021 0 feedthrough
rlabel pdiffusion 472 -2021 472 -2021 0 feedthrough
rlabel pdiffusion 479 -2021 479 -2021 0 feedthrough
rlabel pdiffusion 486 -2021 486 -2021 0 feedthrough
rlabel pdiffusion 493 -2021 493 -2021 0 feedthrough
rlabel pdiffusion 500 -2021 500 -2021 0 feedthrough
rlabel pdiffusion 507 -2021 507 -2021 0 cellNo=767
rlabel pdiffusion 514 -2021 514 -2021 0 feedthrough
rlabel pdiffusion 521 -2021 521 -2021 0 feedthrough
rlabel pdiffusion 528 -2021 528 -2021 0 feedthrough
rlabel pdiffusion 535 -2021 535 -2021 0 feedthrough
rlabel pdiffusion 542 -2021 542 -2021 0 feedthrough
rlabel pdiffusion 549 -2021 549 -2021 0 cellNo=332
rlabel pdiffusion 556 -2021 556 -2021 0 feedthrough
rlabel pdiffusion 563 -2021 563 -2021 0 feedthrough
rlabel pdiffusion 570 -2021 570 -2021 0 cellNo=185
rlabel pdiffusion 577 -2021 577 -2021 0 feedthrough
rlabel pdiffusion 584 -2021 584 -2021 0 feedthrough
rlabel pdiffusion 591 -2021 591 -2021 0 cellNo=20
rlabel pdiffusion 598 -2021 598 -2021 0 feedthrough
rlabel pdiffusion 605 -2021 605 -2021 0 feedthrough
rlabel pdiffusion 612 -2021 612 -2021 0 feedthrough
rlabel pdiffusion 619 -2021 619 -2021 0 feedthrough
rlabel pdiffusion 626 -2021 626 -2021 0 cellNo=939
rlabel pdiffusion 633 -2021 633 -2021 0 feedthrough
rlabel pdiffusion 640 -2021 640 -2021 0 feedthrough
rlabel pdiffusion 647 -2021 647 -2021 0 feedthrough
rlabel pdiffusion 654 -2021 654 -2021 0 feedthrough
rlabel pdiffusion 661 -2021 661 -2021 0 feedthrough
rlabel pdiffusion 668 -2021 668 -2021 0 feedthrough
rlabel pdiffusion 675 -2021 675 -2021 0 feedthrough
rlabel pdiffusion 682 -2021 682 -2021 0 feedthrough
rlabel pdiffusion 689 -2021 689 -2021 0 feedthrough
rlabel pdiffusion 696 -2021 696 -2021 0 feedthrough
rlabel pdiffusion 703 -2021 703 -2021 0 feedthrough
rlabel pdiffusion 710 -2021 710 -2021 0 feedthrough
rlabel pdiffusion 717 -2021 717 -2021 0 cellNo=362
rlabel pdiffusion 724 -2021 724 -2021 0 feedthrough
rlabel pdiffusion 731 -2021 731 -2021 0 feedthrough
rlabel pdiffusion 738 -2021 738 -2021 0 feedthrough
rlabel pdiffusion 745 -2021 745 -2021 0 feedthrough
rlabel pdiffusion 752 -2021 752 -2021 0 feedthrough
rlabel pdiffusion 759 -2021 759 -2021 0 cellNo=423
rlabel pdiffusion 766 -2021 766 -2021 0 feedthrough
rlabel pdiffusion 773 -2021 773 -2021 0 feedthrough
rlabel pdiffusion 780 -2021 780 -2021 0 feedthrough
rlabel pdiffusion 787 -2021 787 -2021 0 feedthrough
rlabel pdiffusion 794 -2021 794 -2021 0 cellNo=430
rlabel pdiffusion 801 -2021 801 -2021 0 feedthrough
rlabel pdiffusion 808 -2021 808 -2021 0 feedthrough
rlabel pdiffusion 815 -2021 815 -2021 0 feedthrough
rlabel pdiffusion 822 -2021 822 -2021 0 feedthrough
rlabel pdiffusion 829 -2021 829 -2021 0 feedthrough
rlabel pdiffusion 836 -2021 836 -2021 0 feedthrough
rlabel pdiffusion 843 -2021 843 -2021 0 feedthrough
rlabel pdiffusion 850 -2021 850 -2021 0 feedthrough
rlabel pdiffusion 857 -2021 857 -2021 0 feedthrough
rlabel pdiffusion 864 -2021 864 -2021 0 feedthrough
rlabel pdiffusion 871 -2021 871 -2021 0 feedthrough
rlabel pdiffusion 878 -2021 878 -2021 0 feedthrough
rlabel pdiffusion 885 -2021 885 -2021 0 cellNo=300
rlabel pdiffusion 892 -2021 892 -2021 0 cellNo=704
rlabel pdiffusion 899 -2021 899 -2021 0 cellNo=603
rlabel pdiffusion 906 -2021 906 -2021 0 feedthrough
rlabel pdiffusion 913 -2021 913 -2021 0 feedthrough
rlabel pdiffusion 920 -2021 920 -2021 0 cellNo=192
rlabel pdiffusion 927 -2021 927 -2021 0 feedthrough
rlabel pdiffusion 934 -2021 934 -2021 0 feedthrough
rlabel pdiffusion 941 -2021 941 -2021 0 feedthrough
rlabel pdiffusion 948 -2021 948 -2021 0 feedthrough
rlabel pdiffusion 955 -2021 955 -2021 0 cellNo=553
rlabel pdiffusion 962 -2021 962 -2021 0 cellNo=798
rlabel pdiffusion 969 -2021 969 -2021 0 feedthrough
rlabel pdiffusion 976 -2021 976 -2021 0 feedthrough
rlabel pdiffusion 983 -2021 983 -2021 0 feedthrough
rlabel pdiffusion 990 -2021 990 -2021 0 cellNo=488
rlabel pdiffusion 997 -2021 997 -2021 0 cellNo=462
rlabel pdiffusion 1004 -2021 1004 -2021 0 feedthrough
rlabel pdiffusion 1011 -2021 1011 -2021 0 feedthrough
rlabel pdiffusion 1018 -2021 1018 -2021 0 feedthrough
rlabel pdiffusion 1025 -2021 1025 -2021 0 feedthrough
rlabel pdiffusion 1032 -2021 1032 -2021 0 feedthrough
rlabel pdiffusion 1039 -2021 1039 -2021 0 cellNo=356
rlabel pdiffusion 1046 -2021 1046 -2021 0 feedthrough
rlabel pdiffusion 1053 -2021 1053 -2021 0 feedthrough
rlabel pdiffusion 1060 -2021 1060 -2021 0 feedthrough
rlabel pdiffusion 1067 -2021 1067 -2021 0 feedthrough
rlabel pdiffusion 1074 -2021 1074 -2021 0 feedthrough
rlabel pdiffusion 1081 -2021 1081 -2021 0 feedthrough
rlabel pdiffusion 1088 -2021 1088 -2021 0 feedthrough
rlabel pdiffusion 1095 -2021 1095 -2021 0 feedthrough
rlabel pdiffusion 1102 -2021 1102 -2021 0 feedthrough
rlabel pdiffusion 1109 -2021 1109 -2021 0 cellNo=101
rlabel pdiffusion 1116 -2021 1116 -2021 0 feedthrough
rlabel pdiffusion 1123 -2021 1123 -2021 0 feedthrough
rlabel pdiffusion 1130 -2021 1130 -2021 0 feedthrough
rlabel pdiffusion 1137 -2021 1137 -2021 0 cellNo=855
rlabel pdiffusion 1144 -2021 1144 -2021 0 feedthrough
rlabel pdiffusion 1151 -2021 1151 -2021 0 feedthrough
rlabel pdiffusion 1158 -2021 1158 -2021 0 feedthrough
rlabel pdiffusion 1165 -2021 1165 -2021 0 feedthrough
rlabel pdiffusion 1172 -2021 1172 -2021 0 feedthrough
rlabel pdiffusion 1179 -2021 1179 -2021 0 feedthrough
rlabel pdiffusion 1186 -2021 1186 -2021 0 feedthrough
rlabel pdiffusion 1193 -2021 1193 -2021 0 cellNo=682
rlabel pdiffusion 1200 -2021 1200 -2021 0 feedthrough
rlabel pdiffusion 1207 -2021 1207 -2021 0 feedthrough
rlabel pdiffusion 1214 -2021 1214 -2021 0 cellNo=721
rlabel pdiffusion 1221 -2021 1221 -2021 0 feedthrough
rlabel pdiffusion 1228 -2021 1228 -2021 0 feedthrough
rlabel pdiffusion 1235 -2021 1235 -2021 0 feedthrough
rlabel pdiffusion 1242 -2021 1242 -2021 0 feedthrough
rlabel pdiffusion 1249 -2021 1249 -2021 0 feedthrough
rlabel pdiffusion 1256 -2021 1256 -2021 0 feedthrough
rlabel pdiffusion 1263 -2021 1263 -2021 0 feedthrough
rlabel pdiffusion 1270 -2021 1270 -2021 0 feedthrough
rlabel pdiffusion 1277 -2021 1277 -2021 0 feedthrough
rlabel pdiffusion 1284 -2021 1284 -2021 0 feedthrough
rlabel pdiffusion 1291 -2021 1291 -2021 0 cellNo=282
rlabel pdiffusion 1298 -2021 1298 -2021 0 feedthrough
rlabel pdiffusion 1305 -2021 1305 -2021 0 feedthrough
rlabel pdiffusion 1312 -2021 1312 -2021 0 feedthrough
rlabel pdiffusion 1319 -2021 1319 -2021 0 feedthrough
rlabel pdiffusion 1326 -2021 1326 -2021 0 feedthrough
rlabel pdiffusion 1333 -2021 1333 -2021 0 feedthrough
rlabel pdiffusion 1340 -2021 1340 -2021 0 feedthrough
rlabel pdiffusion 1347 -2021 1347 -2021 0 feedthrough
rlabel pdiffusion 1354 -2021 1354 -2021 0 feedthrough
rlabel pdiffusion 1361 -2021 1361 -2021 0 feedthrough
rlabel pdiffusion 1368 -2021 1368 -2021 0 feedthrough
rlabel pdiffusion 1375 -2021 1375 -2021 0 feedthrough
rlabel pdiffusion 1382 -2021 1382 -2021 0 feedthrough
rlabel pdiffusion 1389 -2021 1389 -2021 0 feedthrough
rlabel pdiffusion 1396 -2021 1396 -2021 0 feedthrough
rlabel pdiffusion 1403 -2021 1403 -2021 0 feedthrough
rlabel pdiffusion 1410 -2021 1410 -2021 0 feedthrough
rlabel pdiffusion 1417 -2021 1417 -2021 0 feedthrough
rlabel pdiffusion 1424 -2021 1424 -2021 0 feedthrough
rlabel pdiffusion 1431 -2021 1431 -2021 0 feedthrough
rlabel pdiffusion 1438 -2021 1438 -2021 0 feedthrough
rlabel pdiffusion 1445 -2021 1445 -2021 0 feedthrough
rlabel pdiffusion 1452 -2021 1452 -2021 0 feedthrough
rlabel pdiffusion 1459 -2021 1459 -2021 0 feedthrough
rlabel pdiffusion 1466 -2021 1466 -2021 0 feedthrough
rlabel pdiffusion 1473 -2021 1473 -2021 0 feedthrough
rlabel pdiffusion 1480 -2021 1480 -2021 0 feedthrough
rlabel pdiffusion 1487 -2021 1487 -2021 0 feedthrough
rlabel pdiffusion 1494 -2021 1494 -2021 0 feedthrough
rlabel pdiffusion 1501 -2021 1501 -2021 0 feedthrough
rlabel pdiffusion 1508 -2021 1508 -2021 0 feedthrough
rlabel pdiffusion 1515 -2021 1515 -2021 0 feedthrough
rlabel pdiffusion 1522 -2021 1522 -2021 0 feedthrough
rlabel pdiffusion 1529 -2021 1529 -2021 0 feedthrough
rlabel pdiffusion 1536 -2021 1536 -2021 0 feedthrough
rlabel pdiffusion 1543 -2021 1543 -2021 0 feedthrough
rlabel pdiffusion 1550 -2021 1550 -2021 0 feedthrough
rlabel pdiffusion 1557 -2021 1557 -2021 0 feedthrough
rlabel pdiffusion 1564 -2021 1564 -2021 0 feedthrough
rlabel pdiffusion 1571 -2021 1571 -2021 0 feedthrough
rlabel pdiffusion 1578 -2021 1578 -2021 0 feedthrough
rlabel pdiffusion 1585 -2021 1585 -2021 0 feedthrough
rlabel pdiffusion 1592 -2021 1592 -2021 0 feedthrough
rlabel pdiffusion 1599 -2021 1599 -2021 0 feedthrough
rlabel pdiffusion 1606 -2021 1606 -2021 0 feedthrough
rlabel pdiffusion 1613 -2021 1613 -2021 0 feedthrough
rlabel pdiffusion 1620 -2021 1620 -2021 0 feedthrough
rlabel pdiffusion 1627 -2021 1627 -2021 0 feedthrough
rlabel pdiffusion 1634 -2021 1634 -2021 0 feedthrough
rlabel pdiffusion 1641 -2021 1641 -2021 0 feedthrough
rlabel pdiffusion 1648 -2021 1648 -2021 0 feedthrough
rlabel pdiffusion 1655 -2021 1655 -2021 0 feedthrough
rlabel pdiffusion 1662 -2021 1662 -2021 0 feedthrough
rlabel pdiffusion 1669 -2021 1669 -2021 0 feedthrough
rlabel pdiffusion 1676 -2021 1676 -2021 0 feedthrough
rlabel pdiffusion 1683 -2021 1683 -2021 0 feedthrough
rlabel pdiffusion 1690 -2021 1690 -2021 0 feedthrough
rlabel pdiffusion 1697 -2021 1697 -2021 0 feedthrough
rlabel pdiffusion 1704 -2021 1704 -2021 0 feedthrough
rlabel pdiffusion 1711 -2021 1711 -2021 0 feedthrough
rlabel pdiffusion 1718 -2021 1718 -2021 0 feedthrough
rlabel pdiffusion 1725 -2021 1725 -2021 0 feedthrough
rlabel pdiffusion 1732 -2021 1732 -2021 0 feedthrough
rlabel pdiffusion 1739 -2021 1739 -2021 0 feedthrough
rlabel pdiffusion 1746 -2021 1746 -2021 0 cellNo=518
rlabel pdiffusion 1753 -2021 1753 -2021 0 feedthrough
rlabel pdiffusion 1760 -2021 1760 -2021 0 feedthrough
rlabel pdiffusion 1767 -2021 1767 -2021 0 feedthrough
rlabel pdiffusion 1774 -2021 1774 -2021 0 feedthrough
rlabel pdiffusion 1781 -2021 1781 -2021 0 feedthrough
rlabel pdiffusion 1788 -2021 1788 -2021 0 feedthrough
rlabel pdiffusion 1795 -2021 1795 -2021 0 feedthrough
rlabel pdiffusion 1802 -2021 1802 -2021 0 feedthrough
rlabel pdiffusion 1809 -2021 1809 -2021 0 feedthrough
rlabel pdiffusion 3 -2176 3 -2176 0 cellNo=1031
rlabel pdiffusion 10 -2176 10 -2176 0 cellNo=1193
rlabel pdiffusion 17 -2176 17 -2176 0 cellNo=1198
rlabel pdiffusion 24 -2176 24 -2176 0 cellNo=1036
rlabel pdiffusion 31 -2176 31 -2176 0 feedthrough
rlabel pdiffusion 38 -2176 38 -2176 0 feedthrough
rlabel pdiffusion 45 -2176 45 -2176 0 feedthrough
rlabel pdiffusion 52 -2176 52 -2176 0 feedthrough
rlabel pdiffusion 59 -2176 59 -2176 0 cellNo=967
rlabel pdiffusion 66 -2176 66 -2176 0 feedthrough
rlabel pdiffusion 73 -2176 73 -2176 0 feedthrough
rlabel pdiffusion 80 -2176 80 -2176 0 feedthrough
rlabel pdiffusion 87 -2176 87 -2176 0 feedthrough
rlabel pdiffusion 94 -2176 94 -2176 0 cellNo=720
rlabel pdiffusion 101 -2176 101 -2176 0 cellNo=161
rlabel pdiffusion 108 -2176 108 -2176 0 cellNo=765
rlabel pdiffusion 115 -2176 115 -2176 0 feedthrough
rlabel pdiffusion 122 -2176 122 -2176 0 cellNo=514
rlabel pdiffusion 129 -2176 129 -2176 0 cellNo=654
rlabel pdiffusion 136 -2176 136 -2176 0 feedthrough
rlabel pdiffusion 143 -2176 143 -2176 0 feedthrough
rlabel pdiffusion 150 -2176 150 -2176 0 feedthrough
rlabel pdiffusion 157 -2176 157 -2176 0 feedthrough
rlabel pdiffusion 164 -2176 164 -2176 0 feedthrough
rlabel pdiffusion 171 -2176 171 -2176 0 feedthrough
rlabel pdiffusion 178 -2176 178 -2176 0 feedthrough
rlabel pdiffusion 185 -2176 185 -2176 0 feedthrough
rlabel pdiffusion 192 -2176 192 -2176 0 feedthrough
rlabel pdiffusion 199 -2176 199 -2176 0 cellNo=632
rlabel pdiffusion 206 -2176 206 -2176 0 feedthrough
rlabel pdiffusion 213 -2176 213 -2176 0 feedthrough
rlabel pdiffusion 220 -2176 220 -2176 0 feedthrough
rlabel pdiffusion 227 -2176 227 -2176 0 cellNo=90
rlabel pdiffusion 234 -2176 234 -2176 0 feedthrough
rlabel pdiffusion 241 -2176 241 -2176 0 feedthrough
rlabel pdiffusion 248 -2176 248 -2176 0 cellNo=641
rlabel pdiffusion 255 -2176 255 -2176 0 cellNo=323
rlabel pdiffusion 262 -2176 262 -2176 0 feedthrough
rlabel pdiffusion 269 -2176 269 -2176 0 feedthrough
rlabel pdiffusion 276 -2176 276 -2176 0 cellNo=67
rlabel pdiffusion 283 -2176 283 -2176 0 feedthrough
rlabel pdiffusion 290 -2176 290 -2176 0 cellNo=137
rlabel pdiffusion 297 -2176 297 -2176 0 feedthrough
rlabel pdiffusion 304 -2176 304 -2176 0 feedthrough
rlabel pdiffusion 311 -2176 311 -2176 0 feedthrough
rlabel pdiffusion 318 -2176 318 -2176 0 feedthrough
rlabel pdiffusion 325 -2176 325 -2176 0 feedthrough
rlabel pdiffusion 332 -2176 332 -2176 0 feedthrough
rlabel pdiffusion 339 -2176 339 -2176 0 feedthrough
rlabel pdiffusion 346 -2176 346 -2176 0 feedthrough
rlabel pdiffusion 353 -2176 353 -2176 0 feedthrough
rlabel pdiffusion 360 -2176 360 -2176 0 feedthrough
rlabel pdiffusion 367 -2176 367 -2176 0 feedthrough
rlabel pdiffusion 374 -2176 374 -2176 0 cellNo=525
rlabel pdiffusion 381 -2176 381 -2176 0 feedthrough
rlabel pdiffusion 388 -2176 388 -2176 0 feedthrough
rlabel pdiffusion 395 -2176 395 -2176 0 feedthrough
rlabel pdiffusion 402 -2176 402 -2176 0 feedthrough
rlabel pdiffusion 409 -2176 409 -2176 0 feedthrough
rlabel pdiffusion 416 -2176 416 -2176 0 cellNo=107
rlabel pdiffusion 423 -2176 423 -2176 0 feedthrough
rlabel pdiffusion 430 -2176 430 -2176 0 feedthrough
rlabel pdiffusion 437 -2176 437 -2176 0 feedthrough
rlabel pdiffusion 444 -2176 444 -2176 0 feedthrough
rlabel pdiffusion 451 -2176 451 -2176 0 feedthrough
rlabel pdiffusion 458 -2176 458 -2176 0 feedthrough
rlabel pdiffusion 465 -2176 465 -2176 0 feedthrough
rlabel pdiffusion 472 -2176 472 -2176 0 feedthrough
rlabel pdiffusion 479 -2176 479 -2176 0 feedthrough
rlabel pdiffusion 486 -2176 486 -2176 0 feedthrough
rlabel pdiffusion 493 -2176 493 -2176 0 feedthrough
rlabel pdiffusion 500 -2176 500 -2176 0 feedthrough
rlabel pdiffusion 507 -2176 507 -2176 0 feedthrough
rlabel pdiffusion 514 -2176 514 -2176 0 cellNo=466
rlabel pdiffusion 521 -2176 521 -2176 0 feedthrough
rlabel pdiffusion 528 -2176 528 -2176 0 feedthrough
rlabel pdiffusion 535 -2176 535 -2176 0 feedthrough
rlabel pdiffusion 542 -2176 542 -2176 0 feedthrough
rlabel pdiffusion 549 -2176 549 -2176 0 feedthrough
rlabel pdiffusion 556 -2176 556 -2176 0 cellNo=506
rlabel pdiffusion 563 -2176 563 -2176 0 feedthrough
rlabel pdiffusion 570 -2176 570 -2176 0 feedthrough
rlabel pdiffusion 577 -2176 577 -2176 0 feedthrough
rlabel pdiffusion 584 -2176 584 -2176 0 cellNo=815
rlabel pdiffusion 591 -2176 591 -2176 0 feedthrough
rlabel pdiffusion 598 -2176 598 -2176 0 feedthrough
rlabel pdiffusion 605 -2176 605 -2176 0 feedthrough
rlabel pdiffusion 612 -2176 612 -2176 0 cellNo=585
rlabel pdiffusion 619 -2176 619 -2176 0 feedthrough
rlabel pdiffusion 626 -2176 626 -2176 0 cellNo=955
rlabel pdiffusion 633 -2176 633 -2176 0 feedthrough
rlabel pdiffusion 640 -2176 640 -2176 0 feedthrough
rlabel pdiffusion 647 -2176 647 -2176 0 feedthrough
rlabel pdiffusion 654 -2176 654 -2176 0 feedthrough
rlabel pdiffusion 661 -2176 661 -2176 0 feedthrough
rlabel pdiffusion 668 -2176 668 -2176 0 feedthrough
rlabel pdiffusion 675 -2176 675 -2176 0 feedthrough
rlabel pdiffusion 682 -2176 682 -2176 0 feedthrough
rlabel pdiffusion 689 -2176 689 -2176 0 feedthrough
rlabel pdiffusion 696 -2176 696 -2176 0 feedthrough
rlabel pdiffusion 703 -2176 703 -2176 0 cellNo=458
rlabel pdiffusion 710 -2176 710 -2176 0 cellNo=646
rlabel pdiffusion 717 -2176 717 -2176 0 feedthrough
rlabel pdiffusion 724 -2176 724 -2176 0 feedthrough
rlabel pdiffusion 731 -2176 731 -2176 0 feedthrough
rlabel pdiffusion 738 -2176 738 -2176 0 feedthrough
rlabel pdiffusion 745 -2176 745 -2176 0 feedthrough
rlabel pdiffusion 752 -2176 752 -2176 0 feedthrough
rlabel pdiffusion 759 -2176 759 -2176 0 feedthrough
rlabel pdiffusion 766 -2176 766 -2176 0 feedthrough
rlabel pdiffusion 773 -2176 773 -2176 0 feedthrough
rlabel pdiffusion 780 -2176 780 -2176 0 feedthrough
rlabel pdiffusion 787 -2176 787 -2176 0 feedthrough
rlabel pdiffusion 794 -2176 794 -2176 0 feedthrough
rlabel pdiffusion 801 -2176 801 -2176 0 cellNo=480
rlabel pdiffusion 808 -2176 808 -2176 0 feedthrough
rlabel pdiffusion 815 -2176 815 -2176 0 cellNo=301
rlabel pdiffusion 822 -2176 822 -2176 0 cellNo=217
rlabel pdiffusion 829 -2176 829 -2176 0 cellNo=433
rlabel pdiffusion 836 -2176 836 -2176 0 feedthrough
rlabel pdiffusion 843 -2176 843 -2176 0 feedthrough
rlabel pdiffusion 850 -2176 850 -2176 0 feedthrough
rlabel pdiffusion 857 -2176 857 -2176 0 feedthrough
rlabel pdiffusion 864 -2176 864 -2176 0 feedthrough
rlabel pdiffusion 871 -2176 871 -2176 0 cellNo=340
rlabel pdiffusion 878 -2176 878 -2176 0 feedthrough
rlabel pdiffusion 885 -2176 885 -2176 0 feedthrough
rlabel pdiffusion 892 -2176 892 -2176 0 feedthrough
rlabel pdiffusion 899 -2176 899 -2176 0 feedthrough
rlabel pdiffusion 906 -2176 906 -2176 0 feedthrough
rlabel pdiffusion 913 -2176 913 -2176 0 feedthrough
rlabel pdiffusion 920 -2176 920 -2176 0 feedthrough
rlabel pdiffusion 927 -2176 927 -2176 0 cellNo=737
rlabel pdiffusion 934 -2176 934 -2176 0 feedthrough
rlabel pdiffusion 941 -2176 941 -2176 0 feedthrough
rlabel pdiffusion 948 -2176 948 -2176 0 feedthrough
rlabel pdiffusion 955 -2176 955 -2176 0 feedthrough
rlabel pdiffusion 962 -2176 962 -2176 0 feedthrough
rlabel pdiffusion 969 -2176 969 -2176 0 feedthrough
rlabel pdiffusion 976 -2176 976 -2176 0 cellNo=637
rlabel pdiffusion 983 -2176 983 -2176 0 feedthrough
rlabel pdiffusion 990 -2176 990 -2176 0 feedthrough
rlabel pdiffusion 997 -2176 997 -2176 0 cellNo=560
rlabel pdiffusion 1004 -2176 1004 -2176 0 feedthrough
rlabel pdiffusion 1011 -2176 1011 -2176 0 feedthrough
rlabel pdiffusion 1018 -2176 1018 -2176 0 feedthrough
rlabel pdiffusion 1025 -2176 1025 -2176 0 cellNo=434
rlabel pdiffusion 1032 -2176 1032 -2176 0 feedthrough
rlabel pdiffusion 1039 -2176 1039 -2176 0 feedthrough
rlabel pdiffusion 1046 -2176 1046 -2176 0 feedthrough
rlabel pdiffusion 1053 -2176 1053 -2176 0 feedthrough
rlabel pdiffusion 1060 -2176 1060 -2176 0 cellNo=734
rlabel pdiffusion 1067 -2176 1067 -2176 0 feedthrough
rlabel pdiffusion 1074 -2176 1074 -2176 0 feedthrough
rlabel pdiffusion 1081 -2176 1081 -2176 0 feedthrough
rlabel pdiffusion 1088 -2176 1088 -2176 0 feedthrough
rlabel pdiffusion 1095 -2176 1095 -2176 0 feedthrough
rlabel pdiffusion 1102 -2176 1102 -2176 0 feedthrough
rlabel pdiffusion 1109 -2176 1109 -2176 0 feedthrough
rlabel pdiffusion 1116 -2176 1116 -2176 0 feedthrough
rlabel pdiffusion 1123 -2176 1123 -2176 0 cellNo=908
rlabel pdiffusion 1130 -2176 1130 -2176 0 cellNo=534
rlabel pdiffusion 1137 -2176 1137 -2176 0 feedthrough
rlabel pdiffusion 1144 -2176 1144 -2176 0 feedthrough
rlabel pdiffusion 1151 -2176 1151 -2176 0 feedthrough
rlabel pdiffusion 1158 -2176 1158 -2176 0 feedthrough
rlabel pdiffusion 1165 -2176 1165 -2176 0 feedthrough
rlabel pdiffusion 1172 -2176 1172 -2176 0 feedthrough
rlabel pdiffusion 1179 -2176 1179 -2176 0 feedthrough
rlabel pdiffusion 1186 -2176 1186 -2176 0 feedthrough
rlabel pdiffusion 1193 -2176 1193 -2176 0 cellNo=256
rlabel pdiffusion 1200 -2176 1200 -2176 0 feedthrough
rlabel pdiffusion 1207 -2176 1207 -2176 0 feedthrough
rlabel pdiffusion 1214 -2176 1214 -2176 0 feedthrough
rlabel pdiffusion 1221 -2176 1221 -2176 0 feedthrough
rlabel pdiffusion 1228 -2176 1228 -2176 0 feedthrough
rlabel pdiffusion 1235 -2176 1235 -2176 0 feedthrough
rlabel pdiffusion 1242 -2176 1242 -2176 0 feedthrough
rlabel pdiffusion 1249 -2176 1249 -2176 0 feedthrough
rlabel pdiffusion 1256 -2176 1256 -2176 0 feedthrough
rlabel pdiffusion 1263 -2176 1263 -2176 0 feedthrough
rlabel pdiffusion 1270 -2176 1270 -2176 0 feedthrough
rlabel pdiffusion 1277 -2176 1277 -2176 0 feedthrough
rlabel pdiffusion 1284 -2176 1284 -2176 0 feedthrough
rlabel pdiffusion 1291 -2176 1291 -2176 0 feedthrough
rlabel pdiffusion 1298 -2176 1298 -2176 0 feedthrough
rlabel pdiffusion 1305 -2176 1305 -2176 0 feedthrough
rlabel pdiffusion 1312 -2176 1312 -2176 0 cellNo=915
rlabel pdiffusion 1319 -2176 1319 -2176 0 feedthrough
rlabel pdiffusion 1326 -2176 1326 -2176 0 feedthrough
rlabel pdiffusion 1333 -2176 1333 -2176 0 feedthrough
rlabel pdiffusion 1340 -2176 1340 -2176 0 feedthrough
rlabel pdiffusion 1347 -2176 1347 -2176 0 feedthrough
rlabel pdiffusion 1354 -2176 1354 -2176 0 feedthrough
rlabel pdiffusion 1361 -2176 1361 -2176 0 feedthrough
rlabel pdiffusion 1368 -2176 1368 -2176 0 feedthrough
rlabel pdiffusion 1375 -2176 1375 -2176 0 feedthrough
rlabel pdiffusion 1382 -2176 1382 -2176 0 feedthrough
rlabel pdiffusion 1389 -2176 1389 -2176 0 feedthrough
rlabel pdiffusion 1396 -2176 1396 -2176 0 feedthrough
rlabel pdiffusion 1403 -2176 1403 -2176 0 feedthrough
rlabel pdiffusion 1410 -2176 1410 -2176 0 feedthrough
rlabel pdiffusion 1417 -2176 1417 -2176 0 feedthrough
rlabel pdiffusion 1424 -2176 1424 -2176 0 feedthrough
rlabel pdiffusion 1431 -2176 1431 -2176 0 feedthrough
rlabel pdiffusion 1438 -2176 1438 -2176 0 feedthrough
rlabel pdiffusion 1445 -2176 1445 -2176 0 feedthrough
rlabel pdiffusion 1452 -2176 1452 -2176 0 feedthrough
rlabel pdiffusion 1459 -2176 1459 -2176 0 feedthrough
rlabel pdiffusion 1466 -2176 1466 -2176 0 feedthrough
rlabel pdiffusion 1473 -2176 1473 -2176 0 feedthrough
rlabel pdiffusion 1480 -2176 1480 -2176 0 feedthrough
rlabel pdiffusion 1487 -2176 1487 -2176 0 feedthrough
rlabel pdiffusion 1494 -2176 1494 -2176 0 feedthrough
rlabel pdiffusion 1501 -2176 1501 -2176 0 feedthrough
rlabel pdiffusion 1508 -2176 1508 -2176 0 feedthrough
rlabel pdiffusion 1515 -2176 1515 -2176 0 feedthrough
rlabel pdiffusion 1522 -2176 1522 -2176 0 feedthrough
rlabel pdiffusion 1529 -2176 1529 -2176 0 feedthrough
rlabel pdiffusion 1536 -2176 1536 -2176 0 feedthrough
rlabel pdiffusion 1543 -2176 1543 -2176 0 feedthrough
rlabel pdiffusion 1550 -2176 1550 -2176 0 feedthrough
rlabel pdiffusion 1557 -2176 1557 -2176 0 feedthrough
rlabel pdiffusion 1564 -2176 1564 -2176 0 feedthrough
rlabel pdiffusion 1571 -2176 1571 -2176 0 feedthrough
rlabel pdiffusion 1578 -2176 1578 -2176 0 feedthrough
rlabel pdiffusion 1585 -2176 1585 -2176 0 feedthrough
rlabel pdiffusion 1592 -2176 1592 -2176 0 feedthrough
rlabel pdiffusion 1599 -2176 1599 -2176 0 feedthrough
rlabel pdiffusion 1606 -2176 1606 -2176 0 feedthrough
rlabel pdiffusion 1613 -2176 1613 -2176 0 feedthrough
rlabel pdiffusion 1620 -2176 1620 -2176 0 feedthrough
rlabel pdiffusion 1627 -2176 1627 -2176 0 feedthrough
rlabel pdiffusion 1634 -2176 1634 -2176 0 feedthrough
rlabel pdiffusion 1641 -2176 1641 -2176 0 feedthrough
rlabel pdiffusion 1648 -2176 1648 -2176 0 feedthrough
rlabel pdiffusion 1655 -2176 1655 -2176 0 feedthrough
rlabel pdiffusion 1662 -2176 1662 -2176 0 feedthrough
rlabel pdiffusion 1669 -2176 1669 -2176 0 feedthrough
rlabel pdiffusion 1676 -2176 1676 -2176 0 feedthrough
rlabel pdiffusion 1683 -2176 1683 -2176 0 feedthrough
rlabel pdiffusion 1690 -2176 1690 -2176 0 feedthrough
rlabel pdiffusion 1697 -2176 1697 -2176 0 feedthrough
rlabel pdiffusion 1704 -2176 1704 -2176 0 feedthrough
rlabel pdiffusion 1711 -2176 1711 -2176 0 cellNo=756
rlabel pdiffusion 1718 -2176 1718 -2176 0 cellNo=747
rlabel pdiffusion 1725 -2176 1725 -2176 0 feedthrough
rlabel pdiffusion 1732 -2176 1732 -2176 0 feedthrough
rlabel pdiffusion 1739 -2176 1739 -2176 0 feedthrough
rlabel pdiffusion 3 -2305 3 -2305 0 cellNo=1029
rlabel pdiffusion 10 -2305 10 -2305 0 cellNo=1106
rlabel pdiffusion 17 -2305 17 -2305 0 cellNo=1035
rlabel pdiffusion 24 -2305 24 -2305 0 cellNo=1038
rlabel pdiffusion 31 -2305 31 -2305 0 feedthrough
rlabel pdiffusion 38 -2305 38 -2305 0 cellNo=1107
rlabel pdiffusion 45 -2305 45 -2305 0 feedthrough
rlabel pdiffusion 52 -2305 52 -2305 0 cellNo=1235
rlabel pdiffusion 59 -2305 59 -2305 0 feedthrough
rlabel pdiffusion 66 -2305 66 -2305 0 feedthrough
rlabel pdiffusion 73 -2305 73 -2305 0 feedthrough
rlabel pdiffusion 80 -2305 80 -2305 0 cellNo=524
rlabel pdiffusion 87 -2305 87 -2305 0 feedthrough
rlabel pdiffusion 94 -2305 94 -2305 0 feedthrough
rlabel pdiffusion 101 -2305 101 -2305 0 feedthrough
rlabel pdiffusion 108 -2305 108 -2305 0 feedthrough
rlabel pdiffusion 115 -2305 115 -2305 0 feedthrough
rlabel pdiffusion 122 -2305 122 -2305 0 feedthrough
rlabel pdiffusion 129 -2305 129 -2305 0 feedthrough
rlabel pdiffusion 136 -2305 136 -2305 0 cellNo=329
rlabel pdiffusion 143 -2305 143 -2305 0 cellNo=94
rlabel pdiffusion 150 -2305 150 -2305 0 cellNo=1
rlabel pdiffusion 157 -2305 157 -2305 0 feedthrough
rlabel pdiffusion 164 -2305 164 -2305 0 feedthrough
rlabel pdiffusion 171 -2305 171 -2305 0 feedthrough
rlabel pdiffusion 178 -2305 178 -2305 0 feedthrough
rlabel pdiffusion 185 -2305 185 -2305 0 feedthrough
rlabel pdiffusion 192 -2305 192 -2305 0 feedthrough
rlabel pdiffusion 199 -2305 199 -2305 0 feedthrough
rlabel pdiffusion 206 -2305 206 -2305 0 cellNo=25
rlabel pdiffusion 213 -2305 213 -2305 0 cellNo=483
rlabel pdiffusion 220 -2305 220 -2305 0 feedthrough
rlabel pdiffusion 227 -2305 227 -2305 0 feedthrough
rlabel pdiffusion 234 -2305 234 -2305 0 feedthrough
rlabel pdiffusion 241 -2305 241 -2305 0 feedthrough
rlabel pdiffusion 248 -2305 248 -2305 0 feedthrough
rlabel pdiffusion 255 -2305 255 -2305 0 feedthrough
rlabel pdiffusion 262 -2305 262 -2305 0 feedthrough
rlabel pdiffusion 269 -2305 269 -2305 0 feedthrough
rlabel pdiffusion 276 -2305 276 -2305 0 feedthrough
rlabel pdiffusion 283 -2305 283 -2305 0 cellNo=838
rlabel pdiffusion 290 -2305 290 -2305 0 feedthrough
rlabel pdiffusion 297 -2305 297 -2305 0 feedthrough
rlabel pdiffusion 304 -2305 304 -2305 0 feedthrough
rlabel pdiffusion 311 -2305 311 -2305 0 feedthrough
rlabel pdiffusion 318 -2305 318 -2305 0 feedthrough
rlabel pdiffusion 325 -2305 325 -2305 0 feedthrough
rlabel pdiffusion 332 -2305 332 -2305 0 feedthrough
rlabel pdiffusion 339 -2305 339 -2305 0 feedthrough
rlabel pdiffusion 346 -2305 346 -2305 0 feedthrough
rlabel pdiffusion 353 -2305 353 -2305 0 feedthrough
rlabel pdiffusion 360 -2305 360 -2305 0 feedthrough
rlabel pdiffusion 367 -2305 367 -2305 0 feedthrough
rlabel pdiffusion 374 -2305 374 -2305 0 feedthrough
rlabel pdiffusion 381 -2305 381 -2305 0 feedthrough
rlabel pdiffusion 388 -2305 388 -2305 0 feedthrough
rlabel pdiffusion 395 -2305 395 -2305 0 feedthrough
rlabel pdiffusion 402 -2305 402 -2305 0 feedthrough
rlabel pdiffusion 409 -2305 409 -2305 0 feedthrough
rlabel pdiffusion 416 -2305 416 -2305 0 feedthrough
rlabel pdiffusion 423 -2305 423 -2305 0 feedthrough
rlabel pdiffusion 430 -2305 430 -2305 0 feedthrough
rlabel pdiffusion 437 -2305 437 -2305 0 feedthrough
rlabel pdiffusion 444 -2305 444 -2305 0 feedthrough
rlabel pdiffusion 451 -2305 451 -2305 0 cellNo=528
rlabel pdiffusion 458 -2305 458 -2305 0 feedthrough
rlabel pdiffusion 465 -2305 465 -2305 0 feedthrough
rlabel pdiffusion 472 -2305 472 -2305 0 feedthrough
rlabel pdiffusion 479 -2305 479 -2305 0 feedthrough
rlabel pdiffusion 486 -2305 486 -2305 0 feedthrough
rlabel pdiffusion 493 -2305 493 -2305 0 cellNo=878
rlabel pdiffusion 500 -2305 500 -2305 0 feedthrough
rlabel pdiffusion 507 -2305 507 -2305 0 cellNo=69
rlabel pdiffusion 514 -2305 514 -2305 0 feedthrough
rlabel pdiffusion 521 -2305 521 -2305 0 feedthrough
rlabel pdiffusion 528 -2305 528 -2305 0 feedthrough
rlabel pdiffusion 535 -2305 535 -2305 0 feedthrough
rlabel pdiffusion 542 -2305 542 -2305 0 feedthrough
rlabel pdiffusion 549 -2305 549 -2305 0 feedthrough
rlabel pdiffusion 556 -2305 556 -2305 0 feedthrough
rlabel pdiffusion 563 -2305 563 -2305 0 feedthrough
rlabel pdiffusion 570 -2305 570 -2305 0 feedthrough
rlabel pdiffusion 577 -2305 577 -2305 0 cellNo=312
rlabel pdiffusion 584 -2305 584 -2305 0 feedthrough
rlabel pdiffusion 591 -2305 591 -2305 0 feedthrough
rlabel pdiffusion 598 -2305 598 -2305 0 cellNo=126
rlabel pdiffusion 605 -2305 605 -2305 0 feedthrough
rlabel pdiffusion 612 -2305 612 -2305 0 feedthrough
rlabel pdiffusion 619 -2305 619 -2305 0 feedthrough
rlabel pdiffusion 626 -2305 626 -2305 0 cellNo=546
rlabel pdiffusion 633 -2305 633 -2305 0 feedthrough
rlabel pdiffusion 640 -2305 640 -2305 0 cellNo=672
rlabel pdiffusion 647 -2305 647 -2305 0 feedthrough
rlabel pdiffusion 654 -2305 654 -2305 0 feedthrough
rlabel pdiffusion 661 -2305 661 -2305 0 feedthrough
rlabel pdiffusion 668 -2305 668 -2305 0 cellNo=150
rlabel pdiffusion 675 -2305 675 -2305 0 cellNo=352
rlabel pdiffusion 682 -2305 682 -2305 0 feedthrough
rlabel pdiffusion 689 -2305 689 -2305 0 cellNo=708
rlabel pdiffusion 696 -2305 696 -2305 0 cellNo=317
rlabel pdiffusion 703 -2305 703 -2305 0 cellNo=44
rlabel pdiffusion 710 -2305 710 -2305 0 feedthrough
rlabel pdiffusion 717 -2305 717 -2305 0 feedthrough
rlabel pdiffusion 724 -2305 724 -2305 0 feedthrough
rlabel pdiffusion 731 -2305 731 -2305 0 feedthrough
rlabel pdiffusion 738 -2305 738 -2305 0 feedthrough
rlabel pdiffusion 745 -2305 745 -2305 0 feedthrough
rlabel pdiffusion 752 -2305 752 -2305 0 feedthrough
rlabel pdiffusion 759 -2305 759 -2305 0 cellNo=998
rlabel pdiffusion 766 -2305 766 -2305 0 feedthrough
rlabel pdiffusion 773 -2305 773 -2305 0 feedthrough
rlabel pdiffusion 780 -2305 780 -2305 0 cellNo=841
rlabel pdiffusion 787 -2305 787 -2305 0 feedthrough
rlabel pdiffusion 794 -2305 794 -2305 0 feedthrough
rlabel pdiffusion 801 -2305 801 -2305 0 feedthrough
rlabel pdiffusion 808 -2305 808 -2305 0 feedthrough
rlabel pdiffusion 815 -2305 815 -2305 0 feedthrough
rlabel pdiffusion 822 -2305 822 -2305 0 feedthrough
rlabel pdiffusion 829 -2305 829 -2305 0 feedthrough
rlabel pdiffusion 836 -2305 836 -2305 0 cellNo=214
rlabel pdiffusion 843 -2305 843 -2305 0 feedthrough
rlabel pdiffusion 850 -2305 850 -2305 0 feedthrough
rlabel pdiffusion 857 -2305 857 -2305 0 feedthrough
rlabel pdiffusion 864 -2305 864 -2305 0 cellNo=828
rlabel pdiffusion 871 -2305 871 -2305 0 cellNo=314
rlabel pdiffusion 878 -2305 878 -2305 0 feedthrough
rlabel pdiffusion 885 -2305 885 -2305 0 feedthrough
rlabel pdiffusion 892 -2305 892 -2305 0 feedthrough
rlabel pdiffusion 899 -2305 899 -2305 0 feedthrough
rlabel pdiffusion 906 -2305 906 -2305 0 feedthrough
rlabel pdiffusion 913 -2305 913 -2305 0 cellNo=689
rlabel pdiffusion 920 -2305 920 -2305 0 feedthrough
rlabel pdiffusion 927 -2305 927 -2305 0 feedthrough
rlabel pdiffusion 934 -2305 934 -2305 0 feedthrough
rlabel pdiffusion 941 -2305 941 -2305 0 cellNo=394
rlabel pdiffusion 948 -2305 948 -2305 0 feedthrough
rlabel pdiffusion 955 -2305 955 -2305 0 feedthrough
rlabel pdiffusion 962 -2305 962 -2305 0 feedthrough
rlabel pdiffusion 969 -2305 969 -2305 0 feedthrough
rlabel pdiffusion 976 -2305 976 -2305 0 feedthrough
rlabel pdiffusion 983 -2305 983 -2305 0 feedthrough
rlabel pdiffusion 990 -2305 990 -2305 0 feedthrough
rlabel pdiffusion 997 -2305 997 -2305 0 feedthrough
rlabel pdiffusion 1004 -2305 1004 -2305 0 feedthrough
rlabel pdiffusion 1011 -2305 1011 -2305 0 feedthrough
rlabel pdiffusion 1018 -2305 1018 -2305 0 cellNo=961
rlabel pdiffusion 1025 -2305 1025 -2305 0 cellNo=531
rlabel pdiffusion 1032 -2305 1032 -2305 0 feedthrough
rlabel pdiffusion 1039 -2305 1039 -2305 0 cellNo=717
rlabel pdiffusion 1046 -2305 1046 -2305 0 feedthrough
rlabel pdiffusion 1053 -2305 1053 -2305 0 feedthrough
rlabel pdiffusion 1060 -2305 1060 -2305 0 feedthrough
rlabel pdiffusion 1067 -2305 1067 -2305 0 feedthrough
rlabel pdiffusion 1074 -2305 1074 -2305 0 feedthrough
rlabel pdiffusion 1081 -2305 1081 -2305 0 feedthrough
rlabel pdiffusion 1088 -2305 1088 -2305 0 feedthrough
rlabel pdiffusion 1095 -2305 1095 -2305 0 feedthrough
rlabel pdiffusion 1102 -2305 1102 -2305 0 feedthrough
rlabel pdiffusion 1109 -2305 1109 -2305 0 feedthrough
rlabel pdiffusion 1116 -2305 1116 -2305 0 feedthrough
rlabel pdiffusion 1123 -2305 1123 -2305 0 feedthrough
rlabel pdiffusion 1130 -2305 1130 -2305 0 feedthrough
rlabel pdiffusion 1137 -2305 1137 -2305 0 feedthrough
rlabel pdiffusion 1144 -2305 1144 -2305 0 feedthrough
rlabel pdiffusion 1151 -2305 1151 -2305 0 feedthrough
rlabel pdiffusion 1158 -2305 1158 -2305 0 feedthrough
rlabel pdiffusion 1165 -2305 1165 -2305 0 feedthrough
rlabel pdiffusion 1172 -2305 1172 -2305 0 cellNo=830
rlabel pdiffusion 1179 -2305 1179 -2305 0 feedthrough
rlabel pdiffusion 1186 -2305 1186 -2305 0 feedthrough
rlabel pdiffusion 1193 -2305 1193 -2305 0 feedthrough
rlabel pdiffusion 1200 -2305 1200 -2305 0 cellNo=713
rlabel pdiffusion 1207 -2305 1207 -2305 0 feedthrough
rlabel pdiffusion 1214 -2305 1214 -2305 0 feedthrough
rlabel pdiffusion 1221 -2305 1221 -2305 0 feedthrough
rlabel pdiffusion 1228 -2305 1228 -2305 0 feedthrough
rlabel pdiffusion 1235 -2305 1235 -2305 0 feedthrough
rlabel pdiffusion 1242 -2305 1242 -2305 0 cellNo=780
rlabel pdiffusion 1249 -2305 1249 -2305 0 feedthrough
rlabel pdiffusion 1256 -2305 1256 -2305 0 feedthrough
rlabel pdiffusion 1263 -2305 1263 -2305 0 feedthrough
rlabel pdiffusion 1270 -2305 1270 -2305 0 feedthrough
rlabel pdiffusion 1277 -2305 1277 -2305 0 feedthrough
rlabel pdiffusion 1284 -2305 1284 -2305 0 feedthrough
rlabel pdiffusion 1291 -2305 1291 -2305 0 feedthrough
rlabel pdiffusion 1298 -2305 1298 -2305 0 feedthrough
rlabel pdiffusion 1305 -2305 1305 -2305 0 feedthrough
rlabel pdiffusion 1312 -2305 1312 -2305 0 feedthrough
rlabel pdiffusion 1319 -2305 1319 -2305 0 feedthrough
rlabel pdiffusion 1326 -2305 1326 -2305 0 feedthrough
rlabel pdiffusion 1333 -2305 1333 -2305 0 feedthrough
rlabel pdiffusion 1340 -2305 1340 -2305 0 feedthrough
rlabel pdiffusion 1347 -2305 1347 -2305 0 feedthrough
rlabel pdiffusion 1354 -2305 1354 -2305 0 feedthrough
rlabel pdiffusion 1361 -2305 1361 -2305 0 feedthrough
rlabel pdiffusion 1368 -2305 1368 -2305 0 feedthrough
rlabel pdiffusion 1375 -2305 1375 -2305 0 feedthrough
rlabel pdiffusion 1382 -2305 1382 -2305 0 feedthrough
rlabel pdiffusion 1389 -2305 1389 -2305 0 feedthrough
rlabel pdiffusion 1396 -2305 1396 -2305 0 feedthrough
rlabel pdiffusion 1403 -2305 1403 -2305 0 feedthrough
rlabel pdiffusion 1410 -2305 1410 -2305 0 feedthrough
rlabel pdiffusion 1417 -2305 1417 -2305 0 feedthrough
rlabel pdiffusion 1424 -2305 1424 -2305 0 feedthrough
rlabel pdiffusion 1431 -2305 1431 -2305 0 feedthrough
rlabel pdiffusion 1438 -2305 1438 -2305 0 feedthrough
rlabel pdiffusion 1445 -2305 1445 -2305 0 feedthrough
rlabel pdiffusion 1452 -2305 1452 -2305 0 feedthrough
rlabel pdiffusion 1459 -2305 1459 -2305 0 feedthrough
rlabel pdiffusion 1466 -2305 1466 -2305 0 feedthrough
rlabel pdiffusion 1473 -2305 1473 -2305 0 feedthrough
rlabel pdiffusion 1480 -2305 1480 -2305 0 feedthrough
rlabel pdiffusion 1487 -2305 1487 -2305 0 feedthrough
rlabel pdiffusion 1494 -2305 1494 -2305 0 feedthrough
rlabel pdiffusion 1501 -2305 1501 -2305 0 feedthrough
rlabel pdiffusion 1508 -2305 1508 -2305 0 feedthrough
rlabel pdiffusion 1515 -2305 1515 -2305 0 feedthrough
rlabel pdiffusion 1522 -2305 1522 -2305 0 feedthrough
rlabel pdiffusion 1529 -2305 1529 -2305 0 feedthrough
rlabel pdiffusion 1536 -2305 1536 -2305 0 feedthrough
rlabel pdiffusion 1543 -2305 1543 -2305 0 feedthrough
rlabel pdiffusion 1550 -2305 1550 -2305 0 feedthrough
rlabel pdiffusion 1557 -2305 1557 -2305 0 feedthrough
rlabel pdiffusion 1564 -2305 1564 -2305 0 feedthrough
rlabel pdiffusion 1571 -2305 1571 -2305 0 feedthrough
rlabel pdiffusion 1578 -2305 1578 -2305 0 feedthrough
rlabel pdiffusion 1585 -2305 1585 -2305 0 feedthrough
rlabel pdiffusion 1592 -2305 1592 -2305 0 feedthrough
rlabel pdiffusion 1599 -2305 1599 -2305 0 feedthrough
rlabel pdiffusion 1606 -2305 1606 -2305 0 feedthrough
rlabel pdiffusion 1613 -2305 1613 -2305 0 feedthrough
rlabel pdiffusion 1620 -2305 1620 -2305 0 feedthrough
rlabel pdiffusion 1627 -2305 1627 -2305 0 feedthrough
rlabel pdiffusion 1634 -2305 1634 -2305 0 feedthrough
rlabel pdiffusion 1641 -2305 1641 -2305 0 feedthrough
rlabel pdiffusion 1648 -2305 1648 -2305 0 cellNo=929
rlabel pdiffusion 1655 -2305 1655 -2305 0 cellNo=969
rlabel pdiffusion 1662 -2305 1662 -2305 0 feedthrough
rlabel pdiffusion 1669 -2305 1669 -2305 0 cellNo=162
rlabel pdiffusion 1676 -2305 1676 -2305 0 feedthrough
rlabel pdiffusion 1683 -2305 1683 -2305 0 feedthrough
rlabel pdiffusion 1690 -2305 1690 -2305 0 feedthrough
rlabel pdiffusion 1697 -2305 1697 -2305 0 feedthrough
rlabel pdiffusion 3 -2426 3 -2426 0 cellNo=1026
rlabel pdiffusion 10 -2426 10 -2426 0 cellNo=1034
rlabel pdiffusion 17 -2426 17 -2426 0 cellNo=1118
rlabel pdiffusion 24 -2426 24 -2426 0 cellNo=1290
rlabel pdiffusion 31 -2426 31 -2426 0 cellNo=1045
rlabel pdiffusion 38 -2426 38 -2426 0 cellNo=1329
rlabel pdiffusion 45 -2426 45 -2426 0 feedthrough
rlabel pdiffusion 52 -2426 52 -2426 0 feedthrough
rlabel pdiffusion 59 -2426 59 -2426 0 feedthrough
rlabel pdiffusion 66 -2426 66 -2426 0 feedthrough
rlabel pdiffusion 73 -2426 73 -2426 0 feedthrough
rlabel pdiffusion 80 -2426 80 -2426 0 feedthrough
rlabel pdiffusion 87 -2426 87 -2426 0 feedthrough
rlabel pdiffusion 94 -2426 94 -2426 0 feedthrough
rlabel pdiffusion 101 -2426 101 -2426 0 feedthrough
rlabel pdiffusion 108 -2426 108 -2426 0 cellNo=163
rlabel pdiffusion 115 -2426 115 -2426 0 cellNo=623
rlabel pdiffusion 122 -2426 122 -2426 0 feedthrough
rlabel pdiffusion 129 -2426 129 -2426 0 feedthrough
rlabel pdiffusion 136 -2426 136 -2426 0 feedthrough
rlabel pdiffusion 143 -2426 143 -2426 0 feedthrough
rlabel pdiffusion 150 -2426 150 -2426 0 feedthrough
rlabel pdiffusion 157 -2426 157 -2426 0 feedthrough
rlabel pdiffusion 164 -2426 164 -2426 0 feedthrough
rlabel pdiffusion 171 -2426 171 -2426 0 feedthrough
rlabel pdiffusion 178 -2426 178 -2426 0 feedthrough
rlabel pdiffusion 185 -2426 185 -2426 0 feedthrough
rlabel pdiffusion 192 -2426 192 -2426 0 feedthrough
rlabel pdiffusion 199 -2426 199 -2426 0 feedthrough
rlabel pdiffusion 206 -2426 206 -2426 0 feedthrough
rlabel pdiffusion 213 -2426 213 -2426 0 feedthrough
rlabel pdiffusion 220 -2426 220 -2426 0 feedthrough
rlabel pdiffusion 227 -2426 227 -2426 0 cellNo=389
rlabel pdiffusion 234 -2426 234 -2426 0 feedthrough
rlabel pdiffusion 241 -2426 241 -2426 0 feedthrough
rlabel pdiffusion 248 -2426 248 -2426 0 feedthrough
rlabel pdiffusion 255 -2426 255 -2426 0 feedthrough
rlabel pdiffusion 262 -2426 262 -2426 0 feedthrough
rlabel pdiffusion 269 -2426 269 -2426 0 feedthrough
rlabel pdiffusion 276 -2426 276 -2426 0 feedthrough
rlabel pdiffusion 283 -2426 283 -2426 0 cellNo=879
rlabel pdiffusion 290 -2426 290 -2426 0 feedthrough
rlabel pdiffusion 297 -2426 297 -2426 0 feedthrough
rlabel pdiffusion 304 -2426 304 -2426 0 feedthrough
rlabel pdiffusion 311 -2426 311 -2426 0 feedthrough
rlabel pdiffusion 318 -2426 318 -2426 0 feedthrough
rlabel pdiffusion 325 -2426 325 -2426 0 feedthrough
rlabel pdiffusion 332 -2426 332 -2426 0 feedthrough
rlabel pdiffusion 339 -2426 339 -2426 0 feedthrough
rlabel pdiffusion 346 -2426 346 -2426 0 feedthrough
rlabel pdiffusion 353 -2426 353 -2426 0 feedthrough
rlabel pdiffusion 360 -2426 360 -2426 0 feedthrough
rlabel pdiffusion 367 -2426 367 -2426 0 feedthrough
rlabel pdiffusion 374 -2426 374 -2426 0 feedthrough
rlabel pdiffusion 381 -2426 381 -2426 0 feedthrough
rlabel pdiffusion 388 -2426 388 -2426 0 feedthrough
rlabel pdiffusion 395 -2426 395 -2426 0 feedthrough
rlabel pdiffusion 402 -2426 402 -2426 0 cellNo=572
rlabel pdiffusion 409 -2426 409 -2426 0 feedthrough
rlabel pdiffusion 416 -2426 416 -2426 0 feedthrough
rlabel pdiffusion 423 -2426 423 -2426 0 feedthrough
rlabel pdiffusion 430 -2426 430 -2426 0 feedthrough
rlabel pdiffusion 437 -2426 437 -2426 0 feedthrough
rlabel pdiffusion 444 -2426 444 -2426 0 feedthrough
rlabel pdiffusion 451 -2426 451 -2426 0 feedthrough
rlabel pdiffusion 458 -2426 458 -2426 0 feedthrough
rlabel pdiffusion 465 -2426 465 -2426 0 feedthrough
rlabel pdiffusion 472 -2426 472 -2426 0 feedthrough
rlabel pdiffusion 479 -2426 479 -2426 0 feedthrough
rlabel pdiffusion 486 -2426 486 -2426 0 feedthrough
rlabel pdiffusion 493 -2426 493 -2426 0 feedthrough
rlabel pdiffusion 500 -2426 500 -2426 0 feedthrough
rlabel pdiffusion 507 -2426 507 -2426 0 feedthrough
rlabel pdiffusion 514 -2426 514 -2426 0 feedthrough
rlabel pdiffusion 521 -2426 521 -2426 0 cellNo=806
rlabel pdiffusion 528 -2426 528 -2426 0 feedthrough
rlabel pdiffusion 535 -2426 535 -2426 0 feedthrough
rlabel pdiffusion 542 -2426 542 -2426 0 feedthrough
rlabel pdiffusion 549 -2426 549 -2426 0 feedthrough
rlabel pdiffusion 556 -2426 556 -2426 0 feedthrough
rlabel pdiffusion 563 -2426 563 -2426 0 cellNo=493
rlabel pdiffusion 570 -2426 570 -2426 0 feedthrough
rlabel pdiffusion 577 -2426 577 -2426 0 feedthrough
rlabel pdiffusion 584 -2426 584 -2426 0 cellNo=757
rlabel pdiffusion 591 -2426 591 -2426 0 feedthrough
rlabel pdiffusion 598 -2426 598 -2426 0 feedthrough
rlabel pdiffusion 605 -2426 605 -2426 0 feedthrough
rlabel pdiffusion 612 -2426 612 -2426 0 cellNo=991
rlabel pdiffusion 619 -2426 619 -2426 0 cellNo=899
rlabel pdiffusion 626 -2426 626 -2426 0 feedthrough
rlabel pdiffusion 633 -2426 633 -2426 0 cellNo=168
rlabel pdiffusion 640 -2426 640 -2426 0 feedthrough
rlabel pdiffusion 647 -2426 647 -2426 0 cellNo=7
rlabel pdiffusion 654 -2426 654 -2426 0 feedthrough
rlabel pdiffusion 661 -2426 661 -2426 0 feedthrough
rlabel pdiffusion 668 -2426 668 -2426 0 feedthrough
rlabel pdiffusion 675 -2426 675 -2426 0 feedthrough
rlabel pdiffusion 682 -2426 682 -2426 0 cellNo=294
rlabel pdiffusion 689 -2426 689 -2426 0 feedthrough
rlabel pdiffusion 696 -2426 696 -2426 0 feedthrough
rlabel pdiffusion 703 -2426 703 -2426 0 feedthrough
rlabel pdiffusion 710 -2426 710 -2426 0 feedthrough
rlabel pdiffusion 717 -2426 717 -2426 0 feedthrough
rlabel pdiffusion 724 -2426 724 -2426 0 feedthrough
rlabel pdiffusion 731 -2426 731 -2426 0 cellNo=198
rlabel pdiffusion 738 -2426 738 -2426 0 cellNo=557
rlabel pdiffusion 745 -2426 745 -2426 0 cellNo=762
rlabel pdiffusion 752 -2426 752 -2426 0 feedthrough
rlabel pdiffusion 759 -2426 759 -2426 0 feedthrough
rlabel pdiffusion 766 -2426 766 -2426 0 feedthrough
rlabel pdiffusion 773 -2426 773 -2426 0 cellNo=923
rlabel pdiffusion 780 -2426 780 -2426 0 feedthrough
rlabel pdiffusion 787 -2426 787 -2426 0 feedthrough
rlabel pdiffusion 794 -2426 794 -2426 0 feedthrough
rlabel pdiffusion 801 -2426 801 -2426 0 feedthrough
rlabel pdiffusion 808 -2426 808 -2426 0 feedthrough
rlabel pdiffusion 815 -2426 815 -2426 0 feedthrough
rlabel pdiffusion 822 -2426 822 -2426 0 feedthrough
rlabel pdiffusion 829 -2426 829 -2426 0 feedthrough
rlabel pdiffusion 836 -2426 836 -2426 0 cellNo=6
rlabel pdiffusion 843 -2426 843 -2426 0 feedthrough
rlabel pdiffusion 850 -2426 850 -2426 0 cellNo=982
rlabel pdiffusion 857 -2426 857 -2426 0 cellNo=818
rlabel pdiffusion 864 -2426 864 -2426 0 feedthrough
rlabel pdiffusion 871 -2426 871 -2426 0 feedthrough
rlabel pdiffusion 878 -2426 878 -2426 0 feedthrough
rlabel pdiffusion 885 -2426 885 -2426 0 feedthrough
rlabel pdiffusion 892 -2426 892 -2426 0 feedthrough
rlabel pdiffusion 899 -2426 899 -2426 0 feedthrough
rlabel pdiffusion 906 -2426 906 -2426 0 feedthrough
rlabel pdiffusion 913 -2426 913 -2426 0 feedthrough
rlabel pdiffusion 920 -2426 920 -2426 0 cellNo=38
rlabel pdiffusion 927 -2426 927 -2426 0 cellNo=182
rlabel pdiffusion 934 -2426 934 -2426 0 feedthrough
rlabel pdiffusion 941 -2426 941 -2426 0 feedthrough
rlabel pdiffusion 948 -2426 948 -2426 0 feedthrough
rlabel pdiffusion 955 -2426 955 -2426 0 feedthrough
rlabel pdiffusion 962 -2426 962 -2426 0 feedthrough
rlabel pdiffusion 969 -2426 969 -2426 0 cellNo=616
rlabel pdiffusion 976 -2426 976 -2426 0 feedthrough
rlabel pdiffusion 983 -2426 983 -2426 0 feedthrough
rlabel pdiffusion 990 -2426 990 -2426 0 feedthrough
rlabel pdiffusion 997 -2426 997 -2426 0 feedthrough
rlabel pdiffusion 1004 -2426 1004 -2426 0 feedthrough
rlabel pdiffusion 1011 -2426 1011 -2426 0 feedthrough
rlabel pdiffusion 1018 -2426 1018 -2426 0 feedthrough
rlabel pdiffusion 1025 -2426 1025 -2426 0 feedthrough
rlabel pdiffusion 1032 -2426 1032 -2426 0 feedthrough
rlabel pdiffusion 1039 -2426 1039 -2426 0 feedthrough
rlabel pdiffusion 1046 -2426 1046 -2426 0 feedthrough
rlabel pdiffusion 1053 -2426 1053 -2426 0 feedthrough
rlabel pdiffusion 1060 -2426 1060 -2426 0 feedthrough
rlabel pdiffusion 1067 -2426 1067 -2426 0 feedthrough
rlabel pdiffusion 1074 -2426 1074 -2426 0 feedthrough
rlabel pdiffusion 1081 -2426 1081 -2426 0 feedthrough
rlabel pdiffusion 1088 -2426 1088 -2426 0 feedthrough
rlabel pdiffusion 1095 -2426 1095 -2426 0 feedthrough
rlabel pdiffusion 1102 -2426 1102 -2426 0 cellNo=924
rlabel pdiffusion 1109 -2426 1109 -2426 0 feedthrough
rlabel pdiffusion 1116 -2426 1116 -2426 0 feedthrough
rlabel pdiffusion 1123 -2426 1123 -2426 0 cellNo=391
rlabel pdiffusion 1130 -2426 1130 -2426 0 feedthrough
rlabel pdiffusion 1137 -2426 1137 -2426 0 feedthrough
rlabel pdiffusion 1144 -2426 1144 -2426 0 feedthrough
rlabel pdiffusion 1151 -2426 1151 -2426 0 feedthrough
rlabel pdiffusion 1158 -2426 1158 -2426 0 feedthrough
rlabel pdiffusion 1165 -2426 1165 -2426 0 feedthrough
rlabel pdiffusion 1172 -2426 1172 -2426 0 feedthrough
rlabel pdiffusion 1179 -2426 1179 -2426 0 feedthrough
rlabel pdiffusion 1186 -2426 1186 -2426 0 cellNo=996
rlabel pdiffusion 1193 -2426 1193 -2426 0 feedthrough
rlabel pdiffusion 1200 -2426 1200 -2426 0 cellNo=710
rlabel pdiffusion 1207 -2426 1207 -2426 0 feedthrough
rlabel pdiffusion 1214 -2426 1214 -2426 0 feedthrough
rlabel pdiffusion 1221 -2426 1221 -2426 0 feedthrough
rlabel pdiffusion 1228 -2426 1228 -2426 0 feedthrough
rlabel pdiffusion 1235 -2426 1235 -2426 0 cellNo=363
rlabel pdiffusion 1242 -2426 1242 -2426 0 feedthrough
rlabel pdiffusion 1249 -2426 1249 -2426 0 cellNo=56
rlabel pdiffusion 1256 -2426 1256 -2426 0 feedthrough
rlabel pdiffusion 1263 -2426 1263 -2426 0 feedthrough
rlabel pdiffusion 1270 -2426 1270 -2426 0 feedthrough
rlabel pdiffusion 1277 -2426 1277 -2426 0 feedthrough
rlabel pdiffusion 1284 -2426 1284 -2426 0 feedthrough
rlabel pdiffusion 1291 -2426 1291 -2426 0 cellNo=370
rlabel pdiffusion 1298 -2426 1298 -2426 0 feedthrough
rlabel pdiffusion 1305 -2426 1305 -2426 0 feedthrough
rlabel pdiffusion 1312 -2426 1312 -2426 0 feedthrough
rlabel pdiffusion 1319 -2426 1319 -2426 0 feedthrough
rlabel pdiffusion 1326 -2426 1326 -2426 0 feedthrough
rlabel pdiffusion 1333 -2426 1333 -2426 0 feedthrough
rlabel pdiffusion 1340 -2426 1340 -2426 0 feedthrough
rlabel pdiffusion 1347 -2426 1347 -2426 0 feedthrough
rlabel pdiffusion 1354 -2426 1354 -2426 0 feedthrough
rlabel pdiffusion 1361 -2426 1361 -2426 0 cellNo=576
rlabel pdiffusion 1368 -2426 1368 -2426 0 feedthrough
rlabel pdiffusion 1375 -2426 1375 -2426 0 feedthrough
rlabel pdiffusion 1382 -2426 1382 -2426 0 cellNo=242
rlabel pdiffusion 1389 -2426 1389 -2426 0 feedthrough
rlabel pdiffusion 1396 -2426 1396 -2426 0 feedthrough
rlabel pdiffusion 1403 -2426 1403 -2426 0 feedthrough
rlabel pdiffusion 1410 -2426 1410 -2426 0 feedthrough
rlabel pdiffusion 1417 -2426 1417 -2426 0 feedthrough
rlabel pdiffusion 1424 -2426 1424 -2426 0 feedthrough
rlabel pdiffusion 1431 -2426 1431 -2426 0 feedthrough
rlabel pdiffusion 1438 -2426 1438 -2426 0 feedthrough
rlabel pdiffusion 1445 -2426 1445 -2426 0 feedthrough
rlabel pdiffusion 1452 -2426 1452 -2426 0 feedthrough
rlabel pdiffusion 1459 -2426 1459 -2426 0 feedthrough
rlabel pdiffusion 1466 -2426 1466 -2426 0 feedthrough
rlabel pdiffusion 1473 -2426 1473 -2426 0 feedthrough
rlabel pdiffusion 1480 -2426 1480 -2426 0 feedthrough
rlabel pdiffusion 1487 -2426 1487 -2426 0 feedthrough
rlabel pdiffusion 1494 -2426 1494 -2426 0 feedthrough
rlabel pdiffusion 1501 -2426 1501 -2426 0 feedthrough
rlabel pdiffusion 1508 -2426 1508 -2426 0 feedthrough
rlabel pdiffusion 1515 -2426 1515 -2426 0 feedthrough
rlabel pdiffusion 1522 -2426 1522 -2426 0 feedthrough
rlabel pdiffusion 1529 -2426 1529 -2426 0 feedthrough
rlabel pdiffusion 1536 -2426 1536 -2426 0 feedthrough
rlabel pdiffusion 1543 -2426 1543 -2426 0 feedthrough
rlabel pdiffusion 1550 -2426 1550 -2426 0 feedthrough
rlabel pdiffusion 1557 -2426 1557 -2426 0 feedthrough
rlabel pdiffusion 1564 -2426 1564 -2426 0 feedthrough
rlabel pdiffusion 1571 -2426 1571 -2426 0 feedthrough
rlabel pdiffusion 1578 -2426 1578 -2426 0 feedthrough
rlabel pdiffusion 1585 -2426 1585 -2426 0 feedthrough
rlabel pdiffusion 1592 -2426 1592 -2426 0 feedthrough
rlabel pdiffusion 1599 -2426 1599 -2426 0 feedthrough
rlabel pdiffusion 1606 -2426 1606 -2426 0 feedthrough
rlabel pdiffusion 1613 -2426 1613 -2426 0 feedthrough
rlabel pdiffusion 1620 -2426 1620 -2426 0 cellNo=149
rlabel pdiffusion 1627 -2426 1627 -2426 0 feedthrough
rlabel pdiffusion 1634 -2426 1634 -2426 0 feedthrough
rlabel pdiffusion 1641 -2426 1641 -2426 0 cellNo=235
rlabel pdiffusion 1648 -2426 1648 -2426 0 cellNo=579
rlabel pdiffusion 1655 -2426 1655 -2426 0 feedthrough
rlabel pdiffusion 1662 -2426 1662 -2426 0 feedthrough
rlabel pdiffusion 3 -2545 3 -2545 0 cellNo=1033
rlabel pdiffusion 10 -2545 10 -2545 0 cellNo=1091
rlabel pdiffusion 17 -2545 17 -2545 0 cellNo=1041
rlabel pdiffusion 24 -2545 24 -2545 0 cellNo=1455
rlabel pdiffusion 31 -2545 31 -2545 0 cellNo=1049
rlabel pdiffusion 38 -2545 38 -2545 0 cellNo=1054
rlabel pdiffusion 45 -2545 45 -2545 0 cellNo=1255
rlabel pdiffusion 52 -2545 52 -2545 0 feedthrough
rlabel pdiffusion 59 -2545 59 -2545 0 feedthrough
rlabel pdiffusion 66 -2545 66 -2545 0 feedthrough
rlabel pdiffusion 73 -2545 73 -2545 0 feedthrough
rlabel pdiffusion 80 -2545 80 -2545 0 feedthrough
rlabel pdiffusion 87 -2545 87 -2545 0 cellNo=962
rlabel pdiffusion 94 -2545 94 -2545 0 feedthrough
rlabel pdiffusion 101 -2545 101 -2545 0 feedthrough
rlabel pdiffusion 108 -2545 108 -2545 0 feedthrough
rlabel pdiffusion 115 -2545 115 -2545 0 feedthrough
rlabel pdiffusion 122 -2545 122 -2545 0 feedthrough
rlabel pdiffusion 129 -2545 129 -2545 0 feedthrough
rlabel pdiffusion 136 -2545 136 -2545 0 feedthrough
rlabel pdiffusion 143 -2545 143 -2545 0 feedthrough
rlabel pdiffusion 150 -2545 150 -2545 0 feedthrough
rlabel pdiffusion 157 -2545 157 -2545 0 feedthrough
rlabel pdiffusion 164 -2545 164 -2545 0 feedthrough
rlabel pdiffusion 171 -2545 171 -2545 0 cellNo=870
rlabel pdiffusion 178 -2545 178 -2545 0 feedthrough
rlabel pdiffusion 185 -2545 185 -2545 0 feedthrough
rlabel pdiffusion 192 -2545 192 -2545 0 feedthrough
rlabel pdiffusion 199 -2545 199 -2545 0 feedthrough
rlabel pdiffusion 206 -2545 206 -2545 0 feedthrough
rlabel pdiffusion 213 -2545 213 -2545 0 cellNo=258
rlabel pdiffusion 220 -2545 220 -2545 0 feedthrough
rlabel pdiffusion 227 -2545 227 -2545 0 feedthrough
rlabel pdiffusion 234 -2545 234 -2545 0 feedthrough
rlabel pdiffusion 241 -2545 241 -2545 0 feedthrough
rlabel pdiffusion 248 -2545 248 -2545 0 feedthrough
rlabel pdiffusion 255 -2545 255 -2545 0 cellNo=563
rlabel pdiffusion 262 -2545 262 -2545 0 feedthrough
rlabel pdiffusion 269 -2545 269 -2545 0 feedthrough
rlabel pdiffusion 276 -2545 276 -2545 0 cellNo=850
rlabel pdiffusion 283 -2545 283 -2545 0 cellNo=839
rlabel pdiffusion 290 -2545 290 -2545 0 cellNo=187
rlabel pdiffusion 297 -2545 297 -2545 0 cellNo=52
rlabel pdiffusion 304 -2545 304 -2545 0 feedthrough
rlabel pdiffusion 311 -2545 311 -2545 0 feedthrough
rlabel pdiffusion 318 -2545 318 -2545 0 feedthrough
rlabel pdiffusion 325 -2545 325 -2545 0 feedthrough
rlabel pdiffusion 332 -2545 332 -2545 0 feedthrough
rlabel pdiffusion 339 -2545 339 -2545 0 feedthrough
rlabel pdiffusion 346 -2545 346 -2545 0 feedthrough
rlabel pdiffusion 353 -2545 353 -2545 0 feedthrough
rlabel pdiffusion 360 -2545 360 -2545 0 feedthrough
rlabel pdiffusion 367 -2545 367 -2545 0 feedthrough
rlabel pdiffusion 374 -2545 374 -2545 0 feedthrough
rlabel pdiffusion 381 -2545 381 -2545 0 feedthrough
rlabel pdiffusion 388 -2545 388 -2545 0 cellNo=361
rlabel pdiffusion 395 -2545 395 -2545 0 feedthrough
rlabel pdiffusion 402 -2545 402 -2545 0 feedthrough
rlabel pdiffusion 409 -2545 409 -2545 0 feedthrough
rlabel pdiffusion 416 -2545 416 -2545 0 cellNo=374
rlabel pdiffusion 423 -2545 423 -2545 0 feedthrough
rlabel pdiffusion 430 -2545 430 -2545 0 feedthrough
rlabel pdiffusion 437 -2545 437 -2545 0 feedthrough
rlabel pdiffusion 444 -2545 444 -2545 0 feedthrough
rlabel pdiffusion 451 -2545 451 -2545 0 feedthrough
rlabel pdiffusion 458 -2545 458 -2545 0 feedthrough
rlabel pdiffusion 465 -2545 465 -2545 0 feedthrough
rlabel pdiffusion 472 -2545 472 -2545 0 feedthrough
rlabel pdiffusion 479 -2545 479 -2545 0 cellNo=693
rlabel pdiffusion 486 -2545 486 -2545 0 feedthrough
rlabel pdiffusion 493 -2545 493 -2545 0 feedthrough
rlabel pdiffusion 500 -2545 500 -2545 0 feedthrough
rlabel pdiffusion 507 -2545 507 -2545 0 feedthrough
rlabel pdiffusion 514 -2545 514 -2545 0 feedthrough
rlabel pdiffusion 521 -2545 521 -2545 0 feedthrough
rlabel pdiffusion 528 -2545 528 -2545 0 cellNo=225
rlabel pdiffusion 535 -2545 535 -2545 0 feedthrough
rlabel pdiffusion 542 -2545 542 -2545 0 cellNo=134
rlabel pdiffusion 549 -2545 549 -2545 0 feedthrough
rlabel pdiffusion 556 -2545 556 -2545 0 feedthrough
rlabel pdiffusion 563 -2545 563 -2545 0 cellNo=220
rlabel pdiffusion 570 -2545 570 -2545 0 cellNo=327
rlabel pdiffusion 577 -2545 577 -2545 0 feedthrough
rlabel pdiffusion 584 -2545 584 -2545 0 feedthrough
rlabel pdiffusion 591 -2545 591 -2545 0 feedthrough
rlabel pdiffusion 598 -2545 598 -2545 0 cellNo=16
rlabel pdiffusion 605 -2545 605 -2545 0 feedthrough
rlabel pdiffusion 612 -2545 612 -2545 0 feedthrough
rlabel pdiffusion 619 -2545 619 -2545 0 feedthrough
rlabel pdiffusion 626 -2545 626 -2545 0 feedthrough
rlabel pdiffusion 633 -2545 633 -2545 0 feedthrough
rlabel pdiffusion 640 -2545 640 -2545 0 feedthrough
rlabel pdiffusion 647 -2545 647 -2545 0 feedthrough
rlabel pdiffusion 654 -2545 654 -2545 0 feedthrough
rlabel pdiffusion 661 -2545 661 -2545 0 feedthrough
rlabel pdiffusion 668 -2545 668 -2545 0 cellNo=87
rlabel pdiffusion 675 -2545 675 -2545 0 feedthrough
rlabel pdiffusion 682 -2545 682 -2545 0 feedthrough
rlabel pdiffusion 689 -2545 689 -2545 0 feedthrough
rlabel pdiffusion 696 -2545 696 -2545 0 feedthrough
rlabel pdiffusion 703 -2545 703 -2545 0 feedthrough
rlabel pdiffusion 710 -2545 710 -2545 0 feedthrough
rlabel pdiffusion 717 -2545 717 -2545 0 feedthrough
rlabel pdiffusion 724 -2545 724 -2545 0 feedthrough
rlabel pdiffusion 731 -2545 731 -2545 0 cellNo=114
rlabel pdiffusion 738 -2545 738 -2545 0 cellNo=662
rlabel pdiffusion 745 -2545 745 -2545 0 cellNo=683
rlabel pdiffusion 752 -2545 752 -2545 0 cellNo=912
rlabel pdiffusion 759 -2545 759 -2545 0 feedthrough
rlabel pdiffusion 766 -2545 766 -2545 0 feedthrough
rlabel pdiffusion 773 -2545 773 -2545 0 feedthrough
rlabel pdiffusion 780 -2545 780 -2545 0 feedthrough
rlabel pdiffusion 787 -2545 787 -2545 0 cellNo=512
rlabel pdiffusion 794 -2545 794 -2545 0 feedthrough
rlabel pdiffusion 801 -2545 801 -2545 0 cellNo=334
rlabel pdiffusion 808 -2545 808 -2545 0 cellNo=784
rlabel pdiffusion 815 -2545 815 -2545 0 feedthrough
rlabel pdiffusion 822 -2545 822 -2545 0 feedthrough
rlabel pdiffusion 829 -2545 829 -2545 0 cellNo=82
rlabel pdiffusion 836 -2545 836 -2545 0 feedthrough
rlabel pdiffusion 843 -2545 843 -2545 0 feedthrough
rlabel pdiffusion 850 -2545 850 -2545 0 feedthrough
rlabel pdiffusion 857 -2545 857 -2545 0 feedthrough
rlabel pdiffusion 864 -2545 864 -2545 0 feedthrough
rlabel pdiffusion 871 -2545 871 -2545 0 feedthrough
rlabel pdiffusion 878 -2545 878 -2545 0 feedthrough
rlabel pdiffusion 885 -2545 885 -2545 0 feedthrough
rlabel pdiffusion 892 -2545 892 -2545 0 feedthrough
rlabel pdiffusion 899 -2545 899 -2545 0 cellNo=575
rlabel pdiffusion 906 -2545 906 -2545 0 feedthrough
rlabel pdiffusion 913 -2545 913 -2545 0 feedthrough
rlabel pdiffusion 920 -2545 920 -2545 0 feedthrough
rlabel pdiffusion 927 -2545 927 -2545 0 feedthrough
rlabel pdiffusion 934 -2545 934 -2545 0 feedthrough
rlabel pdiffusion 941 -2545 941 -2545 0 feedthrough
rlabel pdiffusion 948 -2545 948 -2545 0 feedthrough
rlabel pdiffusion 955 -2545 955 -2545 0 feedthrough
rlabel pdiffusion 962 -2545 962 -2545 0 feedthrough
rlabel pdiffusion 969 -2545 969 -2545 0 feedthrough
rlabel pdiffusion 976 -2545 976 -2545 0 feedthrough
rlabel pdiffusion 983 -2545 983 -2545 0 feedthrough
rlabel pdiffusion 990 -2545 990 -2545 0 feedthrough
rlabel pdiffusion 997 -2545 997 -2545 0 cellNo=297
rlabel pdiffusion 1004 -2545 1004 -2545 0 feedthrough
rlabel pdiffusion 1011 -2545 1011 -2545 0 cellNo=173
rlabel pdiffusion 1018 -2545 1018 -2545 0 feedthrough
rlabel pdiffusion 1025 -2545 1025 -2545 0 cellNo=601
rlabel pdiffusion 1032 -2545 1032 -2545 0 feedthrough
rlabel pdiffusion 1039 -2545 1039 -2545 0 feedthrough
rlabel pdiffusion 1046 -2545 1046 -2545 0 feedthrough
rlabel pdiffusion 1053 -2545 1053 -2545 0 feedthrough
rlabel pdiffusion 1060 -2545 1060 -2545 0 feedthrough
rlabel pdiffusion 1067 -2545 1067 -2545 0 feedthrough
rlabel pdiffusion 1074 -2545 1074 -2545 0 feedthrough
rlabel pdiffusion 1081 -2545 1081 -2545 0 feedthrough
rlabel pdiffusion 1088 -2545 1088 -2545 0 feedthrough
rlabel pdiffusion 1095 -2545 1095 -2545 0 feedthrough
rlabel pdiffusion 1102 -2545 1102 -2545 0 feedthrough
rlabel pdiffusion 1109 -2545 1109 -2545 0 feedthrough
rlabel pdiffusion 1116 -2545 1116 -2545 0 feedthrough
rlabel pdiffusion 1123 -2545 1123 -2545 0 feedthrough
rlabel pdiffusion 1130 -2545 1130 -2545 0 feedthrough
rlabel pdiffusion 1137 -2545 1137 -2545 0 feedthrough
rlabel pdiffusion 1144 -2545 1144 -2545 0 cellNo=152
rlabel pdiffusion 1151 -2545 1151 -2545 0 feedthrough
rlabel pdiffusion 1158 -2545 1158 -2545 0 feedthrough
rlabel pdiffusion 1165 -2545 1165 -2545 0 feedthrough
rlabel pdiffusion 1172 -2545 1172 -2545 0 feedthrough
rlabel pdiffusion 1179 -2545 1179 -2545 0 feedthrough
rlabel pdiffusion 1186 -2545 1186 -2545 0 feedthrough
rlabel pdiffusion 1193 -2545 1193 -2545 0 feedthrough
rlabel pdiffusion 1200 -2545 1200 -2545 0 feedthrough
rlabel pdiffusion 1207 -2545 1207 -2545 0 feedthrough
rlabel pdiffusion 1214 -2545 1214 -2545 0 feedthrough
rlabel pdiffusion 1221 -2545 1221 -2545 0 feedthrough
rlabel pdiffusion 1228 -2545 1228 -2545 0 feedthrough
rlabel pdiffusion 1235 -2545 1235 -2545 0 feedthrough
rlabel pdiffusion 1242 -2545 1242 -2545 0 feedthrough
rlabel pdiffusion 1249 -2545 1249 -2545 0 cellNo=103
rlabel pdiffusion 1256 -2545 1256 -2545 0 feedthrough
rlabel pdiffusion 1263 -2545 1263 -2545 0 feedthrough
rlabel pdiffusion 1270 -2545 1270 -2545 0 feedthrough
rlabel pdiffusion 1277 -2545 1277 -2545 0 feedthrough
rlabel pdiffusion 1284 -2545 1284 -2545 0 feedthrough
rlabel pdiffusion 1291 -2545 1291 -2545 0 feedthrough
rlabel pdiffusion 1298 -2545 1298 -2545 0 feedthrough
rlabel pdiffusion 1305 -2545 1305 -2545 0 feedthrough
rlabel pdiffusion 1312 -2545 1312 -2545 0 feedthrough
rlabel pdiffusion 1319 -2545 1319 -2545 0 feedthrough
rlabel pdiffusion 1326 -2545 1326 -2545 0 feedthrough
rlabel pdiffusion 1333 -2545 1333 -2545 0 feedthrough
rlabel pdiffusion 1340 -2545 1340 -2545 0 feedthrough
rlabel pdiffusion 1347 -2545 1347 -2545 0 feedthrough
rlabel pdiffusion 1354 -2545 1354 -2545 0 feedthrough
rlabel pdiffusion 1361 -2545 1361 -2545 0 feedthrough
rlabel pdiffusion 1368 -2545 1368 -2545 0 feedthrough
rlabel pdiffusion 1375 -2545 1375 -2545 0 feedthrough
rlabel pdiffusion 1382 -2545 1382 -2545 0 feedthrough
rlabel pdiffusion 1389 -2545 1389 -2545 0 feedthrough
rlabel pdiffusion 1396 -2545 1396 -2545 0 feedthrough
rlabel pdiffusion 1403 -2545 1403 -2545 0 cellNo=465
rlabel pdiffusion 1410 -2545 1410 -2545 0 feedthrough
rlabel pdiffusion 1417 -2545 1417 -2545 0 feedthrough
rlabel pdiffusion 1424 -2545 1424 -2545 0 feedthrough
rlabel pdiffusion 1431 -2545 1431 -2545 0 feedthrough
rlabel pdiffusion 1438 -2545 1438 -2545 0 feedthrough
rlabel pdiffusion 1445 -2545 1445 -2545 0 feedthrough
rlabel pdiffusion 1452 -2545 1452 -2545 0 feedthrough
rlabel pdiffusion 1459 -2545 1459 -2545 0 feedthrough
rlabel pdiffusion 1466 -2545 1466 -2545 0 feedthrough
rlabel pdiffusion 1473 -2545 1473 -2545 0 feedthrough
rlabel pdiffusion 1480 -2545 1480 -2545 0 feedthrough
rlabel pdiffusion 1487 -2545 1487 -2545 0 feedthrough
rlabel pdiffusion 1494 -2545 1494 -2545 0 feedthrough
rlabel pdiffusion 1501 -2545 1501 -2545 0 feedthrough
rlabel pdiffusion 1508 -2545 1508 -2545 0 feedthrough
rlabel pdiffusion 1515 -2545 1515 -2545 0 feedthrough
rlabel pdiffusion 1522 -2545 1522 -2545 0 feedthrough
rlabel pdiffusion 1529 -2545 1529 -2545 0 feedthrough
rlabel pdiffusion 1536 -2545 1536 -2545 0 feedthrough
rlabel pdiffusion 1543 -2545 1543 -2545 0 feedthrough
rlabel pdiffusion 1550 -2545 1550 -2545 0 feedthrough
rlabel pdiffusion 1557 -2545 1557 -2545 0 feedthrough
rlabel pdiffusion 1564 -2545 1564 -2545 0 feedthrough
rlabel pdiffusion 1571 -2545 1571 -2545 0 feedthrough
rlabel pdiffusion 1578 -2545 1578 -2545 0 feedthrough
rlabel pdiffusion 1585 -2545 1585 -2545 0 cellNo=538
rlabel pdiffusion 1592 -2545 1592 -2545 0 feedthrough
rlabel pdiffusion 1599 -2545 1599 -2545 0 feedthrough
rlabel pdiffusion 1606 -2545 1606 -2545 0 feedthrough
rlabel pdiffusion 1613 -2545 1613 -2545 0 cellNo=945
rlabel pdiffusion 1641 -2545 1641 -2545 0 feedthrough
rlabel pdiffusion 3 -2674 3 -2674 0 cellNo=1037
rlabel pdiffusion 10 -2674 10 -2674 0 cellNo=1040
rlabel pdiffusion 17 -2674 17 -2674 0 cellNo=1066
rlabel pdiffusion 24 -2674 24 -2674 0 cellNo=1048
rlabel pdiffusion 31 -2674 31 -2674 0 cellNo=1373
rlabel pdiffusion 38 -2674 38 -2674 0 cellNo=1058
rlabel pdiffusion 45 -2674 45 -2674 0 feedthrough
rlabel pdiffusion 52 -2674 52 -2674 0 feedthrough
rlabel pdiffusion 59 -2674 59 -2674 0 feedthrough
rlabel pdiffusion 66 -2674 66 -2674 0 feedthrough
rlabel pdiffusion 73 -2674 73 -2674 0 feedthrough
rlabel pdiffusion 80 -2674 80 -2674 0 feedthrough
rlabel pdiffusion 87 -2674 87 -2674 0 feedthrough
rlabel pdiffusion 94 -2674 94 -2674 0 feedthrough
rlabel pdiffusion 101 -2674 101 -2674 0 feedthrough
rlabel pdiffusion 108 -2674 108 -2674 0 feedthrough
rlabel pdiffusion 115 -2674 115 -2674 0 feedthrough
rlabel pdiffusion 122 -2674 122 -2674 0 feedthrough
rlabel pdiffusion 129 -2674 129 -2674 0 cellNo=735
rlabel pdiffusion 136 -2674 136 -2674 0 feedthrough
rlabel pdiffusion 143 -2674 143 -2674 0 feedthrough
rlabel pdiffusion 150 -2674 150 -2674 0 cellNo=428
rlabel pdiffusion 157 -2674 157 -2674 0 cellNo=14
rlabel pdiffusion 164 -2674 164 -2674 0 feedthrough
rlabel pdiffusion 171 -2674 171 -2674 0 feedthrough
rlabel pdiffusion 178 -2674 178 -2674 0 cellNo=752
rlabel pdiffusion 185 -2674 185 -2674 0 feedthrough
rlabel pdiffusion 192 -2674 192 -2674 0 feedthrough
rlabel pdiffusion 199 -2674 199 -2674 0 cellNo=476
rlabel pdiffusion 206 -2674 206 -2674 0 cellNo=976
rlabel pdiffusion 213 -2674 213 -2674 0 feedthrough
rlabel pdiffusion 220 -2674 220 -2674 0 feedthrough
rlabel pdiffusion 227 -2674 227 -2674 0 feedthrough
rlabel pdiffusion 234 -2674 234 -2674 0 cellNo=236
rlabel pdiffusion 241 -2674 241 -2674 0 feedthrough
rlabel pdiffusion 248 -2674 248 -2674 0 cellNo=31
rlabel pdiffusion 255 -2674 255 -2674 0 feedthrough
rlabel pdiffusion 262 -2674 262 -2674 0 cellNo=892
rlabel pdiffusion 269 -2674 269 -2674 0 feedthrough
rlabel pdiffusion 276 -2674 276 -2674 0 feedthrough
rlabel pdiffusion 283 -2674 283 -2674 0 feedthrough
rlabel pdiffusion 290 -2674 290 -2674 0 feedthrough
rlabel pdiffusion 297 -2674 297 -2674 0 feedthrough
rlabel pdiffusion 304 -2674 304 -2674 0 feedthrough
rlabel pdiffusion 311 -2674 311 -2674 0 feedthrough
rlabel pdiffusion 318 -2674 318 -2674 0 feedthrough
rlabel pdiffusion 325 -2674 325 -2674 0 feedthrough
rlabel pdiffusion 332 -2674 332 -2674 0 feedthrough
rlabel pdiffusion 339 -2674 339 -2674 0 feedthrough
rlabel pdiffusion 346 -2674 346 -2674 0 feedthrough
rlabel pdiffusion 353 -2674 353 -2674 0 feedthrough
rlabel pdiffusion 360 -2674 360 -2674 0 feedthrough
rlabel pdiffusion 367 -2674 367 -2674 0 feedthrough
rlabel pdiffusion 374 -2674 374 -2674 0 cellNo=412
rlabel pdiffusion 381 -2674 381 -2674 0 feedthrough
rlabel pdiffusion 388 -2674 388 -2674 0 feedthrough
rlabel pdiffusion 395 -2674 395 -2674 0 cellNo=633
rlabel pdiffusion 402 -2674 402 -2674 0 feedthrough
rlabel pdiffusion 409 -2674 409 -2674 0 feedthrough
rlabel pdiffusion 416 -2674 416 -2674 0 feedthrough
rlabel pdiffusion 423 -2674 423 -2674 0 cellNo=552
rlabel pdiffusion 430 -2674 430 -2674 0 feedthrough
rlabel pdiffusion 437 -2674 437 -2674 0 feedthrough
rlabel pdiffusion 444 -2674 444 -2674 0 feedthrough
rlabel pdiffusion 451 -2674 451 -2674 0 feedthrough
rlabel pdiffusion 458 -2674 458 -2674 0 feedthrough
rlabel pdiffusion 465 -2674 465 -2674 0 feedthrough
rlabel pdiffusion 472 -2674 472 -2674 0 feedthrough
rlabel pdiffusion 479 -2674 479 -2674 0 feedthrough
rlabel pdiffusion 486 -2674 486 -2674 0 feedthrough
rlabel pdiffusion 493 -2674 493 -2674 0 feedthrough
rlabel pdiffusion 500 -2674 500 -2674 0 cellNo=272
rlabel pdiffusion 507 -2674 507 -2674 0 feedthrough
rlabel pdiffusion 514 -2674 514 -2674 0 feedthrough
rlabel pdiffusion 521 -2674 521 -2674 0 feedthrough
rlabel pdiffusion 528 -2674 528 -2674 0 feedthrough
rlabel pdiffusion 535 -2674 535 -2674 0 feedthrough
rlabel pdiffusion 542 -2674 542 -2674 0 feedthrough
rlabel pdiffusion 549 -2674 549 -2674 0 feedthrough
rlabel pdiffusion 556 -2674 556 -2674 0 feedthrough
rlabel pdiffusion 563 -2674 563 -2674 0 feedthrough
rlabel pdiffusion 570 -2674 570 -2674 0 feedthrough
rlabel pdiffusion 577 -2674 577 -2674 0 feedthrough
rlabel pdiffusion 584 -2674 584 -2674 0 feedthrough
rlabel pdiffusion 591 -2674 591 -2674 0 feedthrough
rlabel pdiffusion 598 -2674 598 -2674 0 feedthrough
rlabel pdiffusion 605 -2674 605 -2674 0 feedthrough
rlabel pdiffusion 612 -2674 612 -2674 0 cellNo=293
rlabel pdiffusion 619 -2674 619 -2674 0 feedthrough
rlabel pdiffusion 626 -2674 626 -2674 0 feedthrough
rlabel pdiffusion 633 -2674 633 -2674 0 feedthrough
rlabel pdiffusion 640 -2674 640 -2674 0 feedthrough
rlabel pdiffusion 647 -2674 647 -2674 0 cellNo=39
rlabel pdiffusion 654 -2674 654 -2674 0 cellNo=913
rlabel pdiffusion 661 -2674 661 -2674 0 feedthrough
rlabel pdiffusion 668 -2674 668 -2674 0 feedthrough
rlabel pdiffusion 675 -2674 675 -2674 0 feedthrough
rlabel pdiffusion 682 -2674 682 -2674 0 feedthrough
rlabel pdiffusion 689 -2674 689 -2674 0 feedthrough
rlabel pdiffusion 696 -2674 696 -2674 0 feedthrough
rlabel pdiffusion 703 -2674 703 -2674 0 feedthrough
rlabel pdiffusion 710 -2674 710 -2674 0 feedthrough
rlabel pdiffusion 717 -2674 717 -2674 0 cellNo=484
rlabel pdiffusion 724 -2674 724 -2674 0 feedthrough
rlabel pdiffusion 731 -2674 731 -2674 0 cellNo=599
rlabel pdiffusion 738 -2674 738 -2674 0 feedthrough
rlabel pdiffusion 745 -2674 745 -2674 0 feedthrough
rlabel pdiffusion 752 -2674 752 -2674 0 feedthrough
rlabel pdiffusion 759 -2674 759 -2674 0 feedthrough
rlabel pdiffusion 766 -2674 766 -2674 0 feedthrough
rlabel pdiffusion 773 -2674 773 -2674 0 feedthrough
rlabel pdiffusion 780 -2674 780 -2674 0 feedthrough
rlabel pdiffusion 787 -2674 787 -2674 0 feedthrough
rlabel pdiffusion 794 -2674 794 -2674 0 feedthrough
rlabel pdiffusion 801 -2674 801 -2674 0 cellNo=932
rlabel pdiffusion 808 -2674 808 -2674 0 feedthrough
rlabel pdiffusion 815 -2674 815 -2674 0 feedthrough
rlabel pdiffusion 822 -2674 822 -2674 0 feedthrough
rlabel pdiffusion 829 -2674 829 -2674 0 feedthrough
rlabel pdiffusion 836 -2674 836 -2674 0 feedthrough
rlabel pdiffusion 843 -2674 843 -2674 0 feedthrough
rlabel pdiffusion 850 -2674 850 -2674 0 feedthrough
rlabel pdiffusion 857 -2674 857 -2674 0 cellNo=951
rlabel pdiffusion 864 -2674 864 -2674 0 feedthrough
rlabel pdiffusion 871 -2674 871 -2674 0 feedthrough
rlabel pdiffusion 878 -2674 878 -2674 0 cellNo=322
rlabel pdiffusion 885 -2674 885 -2674 0 cellNo=664
rlabel pdiffusion 892 -2674 892 -2674 0 feedthrough
rlabel pdiffusion 899 -2674 899 -2674 0 cellNo=207
rlabel pdiffusion 906 -2674 906 -2674 0 cellNo=949
rlabel pdiffusion 913 -2674 913 -2674 0 feedthrough
rlabel pdiffusion 920 -2674 920 -2674 0 feedthrough
rlabel pdiffusion 927 -2674 927 -2674 0 feedthrough
rlabel pdiffusion 934 -2674 934 -2674 0 feedthrough
rlabel pdiffusion 941 -2674 941 -2674 0 feedthrough
rlabel pdiffusion 948 -2674 948 -2674 0 cellNo=99
rlabel pdiffusion 955 -2674 955 -2674 0 cellNo=526
rlabel pdiffusion 962 -2674 962 -2674 0 feedthrough
rlabel pdiffusion 969 -2674 969 -2674 0 cellNo=335
rlabel pdiffusion 976 -2674 976 -2674 0 cellNo=388
rlabel pdiffusion 983 -2674 983 -2674 0 feedthrough
rlabel pdiffusion 990 -2674 990 -2674 0 feedthrough
rlabel pdiffusion 997 -2674 997 -2674 0 feedthrough
rlabel pdiffusion 1004 -2674 1004 -2674 0 feedthrough
rlabel pdiffusion 1011 -2674 1011 -2674 0 feedthrough
rlabel pdiffusion 1018 -2674 1018 -2674 0 feedthrough
rlabel pdiffusion 1025 -2674 1025 -2674 0 cellNo=763
rlabel pdiffusion 1032 -2674 1032 -2674 0 feedthrough
rlabel pdiffusion 1039 -2674 1039 -2674 0 feedthrough
rlabel pdiffusion 1046 -2674 1046 -2674 0 feedthrough
rlabel pdiffusion 1053 -2674 1053 -2674 0 feedthrough
rlabel pdiffusion 1060 -2674 1060 -2674 0 feedthrough
rlabel pdiffusion 1067 -2674 1067 -2674 0 feedthrough
rlabel pdiffusion 1074 -2674 1074 -2674 0 feedthrough
rlabel pdiffusion 1081 -2674 1081 -2674 0 feedthrough
rlabel pdiffusion 1088 -2674 1088 -2674 0 cellNo=232
rlabel pdiffusion 1095 -2674 1095 -2674 0 feedthrough
rlabel pdiffusion 1102 -2674 1102 -2674 0 feedthrough
rlabel pdiffusion 1109 -2674 1109 -2674 0 feedthrough
rlabel pdiffusion 1116 -2674 1116 -2674 0 feedthrough
rlabel pdiffusion 1123 -2674 1123 -2674 0 feedthrough
rlabel pdiffusion 1130 -2674 1130 -2674 0 feedthrough
rlabel pdiffusion 1137 -2674 1137 -2674 0 feedthrough
rlabel pdiffusion 1144 -2674 1144 -2674 0 feedthrough
rlabel pdiffusion 1151 -2674 1151 -2674 0 cellNo=172
rlabel pdiffusion 1158 -2674 1158 -2674 0 feedthrough
rlabel pdiffusion 1165 -2674 1165 -2674 0 feedthrough
rlabel pdiffusion 1172 -2674 1172 -2674 0 feedthrough
rlabel pdiffusion 1179 -2674 1179 -2674 0 feedthrough
rlabel pdiffusion 1186 -2674 1186 -2674 0 cellNo=315
rlabel pdiffusion 1193 -2674 1193 -2674 0 feedthrough
rlabel pdiffusion 1200 -2674 1200 -2674 0 feedthrough
rlabel pdiffusion 1207 -2674 1207 -2674 0 feedthrough
rlabel pdiffusion 1214 -2674 1214 -2674 0 feedthrough
rlabel pdiffusion 1221 -2674 1221 -2674 0 feedthrough
rlabel pdiffusion 1228 -2674 1228 -2674 0 feedthrough
rlabel pdiffusion 1235 -2674 1235 -2674 0 feedthrough
rlabel pdiffusion 1242 -2674 1242 -2674 0 feedthrough
rlabel pdiffusion 1249 -2674 1249 -2674 0 feedthrough
rlabel pdiffusion 1256 -2674 1256 -2674 0 feedthrough
rlabel pdiffusion 1263 -2674 1263 -2674 0 feedthrough
rlabel pdiffusion 1270 -2674 1270 -2674 0 feedthrough
rlabel pdiffusion 1277 -2674 1277 -2674 0 feedthrough
rlabel pdiffusion 1284 -2674 1284 -2674 0 feedthrough
rlabel pdiffusion 1291 -2674 1291 -2674 0 feedthrough
rlabel pdiffusion 1298 -2674 1298 -2674 0 feedthrough
rlabel pdiffusion 1305 -2674 1305 -2674 0 feedthrough
rlabel pdiffusion 1312 -2674 1312 -2674 0 feedthrough
rlabel pdiffusion 1319 -2674 1319 -2674 0 feedthrough
rlabel pdiffusion 1326 -2674 1326 -2674 0 feedthrough
rlabel pdiffusion 1333 -2674 1333 -2674 0 feedthrough
rlabel pdiffusion 1340 -2674 1340 -2674 0 feedthrough
rlabel pdiffusion 1347 -2674 1347 -2674 0 feedthrough
rlabel pdiffusion 1354 -2674 1354 -2674 0 feedthrough
rlabel pdiffusion 1361 -2674 1361 -2674 0 feedthrough
rlabel pdiffusion 1368 -2674 1368 -2674 0 feedthrough
rlabel pdiffusion 1375 -2674 1375 -2674 0 feedthrough
rlabel pdiffusion 1382 -2674 1382 -2674 0 feedthrough
rlabel pdiffusion 1389 -2674 1389 -2674 0 feedthrough
rlabel pdiffusion 1396 -2674 1396 -2674 0 feedthrough
rlabel pdiffusion 1403 -2674 1403 -2674 0 feedthrough
rlabel pdiffusion 1410 -2674 1410 -2674 0 feedthrough
rlabel pdiffusion 1417 -2674 1417 -2674 0 feedthrough
rlabel pdiffusion 1424 -2674 1424 -2674 0 feedthrough
rlabel pdiffusion 1431 -2674 1431 -2674 0 feedthrough
rlabel pdiffusion 1438 -2674 1438 -2674 0 feedthrough
rlabel pdiffusion 1445 -2674 1445 -2674 0 feedthrough
rlabel pdiffusion 1452 -2674 1452 -2674 0 feedthrough
rlabel pdiffusion 1459 -2674 1459 -2674 0 feedthrough
rlabel pdiffusion 1466 -2674 1466 -2674 0 feedthrough
rlabel pdiffusion 1473 -2674 1473 -2674 0 feedthrough
rlabel pdiffusion 1480 -2674 1480 -2674 0 feedthrough
rlabel pdiffusion 1487 -2674 1487 -2674 0 feedthrough
rlabel pdiffusion 1494 -2674 1494 -2674 0 feedthrough
rlabel pdiffusion 1501 -2674 1501 -2674 0 feedthrough
rlabel pdiffusion 1508 -2674 1508 -2674 0 feedthrough
rlabel pdiffusion 1515 -2674 1515 -2674 0 feedthrough
rlabel pdiffusion 1522 -2674 1522 -2674 0 feedthrough
rlabel pdiffusion 1529 -2674 1529 -2674 0 feedthrough
rlabel pdiffusion 1536 -2674 1536 -2674 0 feedthrough
rlabel pdiffusion 1543 -2674 1543 -2674 0 feedthrough
rlabel pdiffusion 1550 -2674 1550 -2674 0 feedthrough
rlabel pdiffusion 1557 -2674 1557 -2674 0 feedthrough
rlabel pdiffusion 1564 -2674 1564 -2674 0 feedthrough
rlabel pdiffusion 1571 -2674 1571 -2674 0 feedthrough
rlabel pdiffusion 1578 -2674 1578 -2674 0 feedthrough
rlabel pdiffusion 1585 -2674 1585 -2674 0 feedthrough
rlabel pdiffusion 1592 -2674 1592 -2674 0 feedthrough
rlabel pdiffusion 1599 -2674 1599 -2674 0 feedthrough
rlabel pdiffusion 1606 -2674 1606 -2674 0 feedthrough
rlabel pdiffusion 1613 -2674 1613 -2674 0 feedthrough
rlabel pdiffusion 1620 -2674 1620 -2674 0 feedthrough
rlabel pdiffusion 1627 -2674 1627 -2674 0 cellNo=171
rlabel pdiffusion 1634 -2674 1634 -2674 0 cellNo=147
rlabel pdiffusion 3 -2787 3 -2787 0 cellNo=1039
rlabel pdiffusion 10 -2787 10 -2787 0 cellNo=1044
rlabel pdiffusion 17 -2787 17 -2787 0 cellNo=1047
rlabel pdiffusion 24 -2787 24 -2787 0 cellNo=1053
rlabel pdiffusion 31 -2787 31 -2787 0 cellNo=1057
rlabel pdiffusion 38 -2787 38 -2787 0 cellNo=1062
rlabel pdiffusion 45 -2787 45 -2787 0 feedthrough
rlabel pdiffusion 52 -2787 52 -2787 0 cellNo=1090
rlabel pdiffusion 59 -2787 59 -2787 0 feedthrough
rlabel pdiffusion 66 -2787 66 -2787 0 feedthrough
rlabel pdiffusion 73 -2787 73 -2787 0 feedthrough
rlabel pdiffusion 80 -2787 80 -2787 0 feedthrough
rlabel pdiffusion 87 -2787 87 -2787 0 feedthrough
rlabel pdiffusion 94 -2787 94 -2787 0 feedthrough
rlabel pdiffusion 101 -2787 101 -2787 0 feedthrough
rlabel pdiffusion 108 -2787 108 -2787 0 cellNo=438
rlabel pdiffusion 115 -2787 115 -2787 0 feedthrough
rlabel pdiffusion 122 -2787 122 -2787 0 cellNo=974
rlabel pdiffusion 129 -2787 129 -2787 0 cellNo=117
rlabel pdiffusion 136 -2787 136 -2787 0 cellNo=707
rlabel pdiffusion 143 -2787 143 -2787 0 feedthrough
rlabel pdiffusion 150 -2787 150 -2787 0 feedthrough
rlabel pdiffusion 157 -2787 157 -2787 0 cellNo=64
rlabel pdiffusion 164 -2787 164 -2787 0 feedthrough
rlabel pdiffusion 171 -2787 171 -2787 0 feedthrough
rlabel pdiffusion 178 -2787 178 -2787 0 feedthrough
rlabel pdiffusion 185 -2787 185 -2787 0 feedthrough
rlabel pdiffusion 192 -2787 192 -2787 0 feedthrough
rlabel pdiffusion 199 -2787 199 -2787 0 feedthrough
rlabel pdiffusion 206 -2787 206 -2787 0 feedthrough
rlabel pdiffusion 213 -2787 213 -2787 0 cellNo=355
rlabel pdiffusion 220 -2787 220 -2787 0 feedthrough
rlabel pdiffusion 227 -2787 227 -2787 0 feedthrough
rlabel pdiffusion 234 -2787 234 -2787 0 cellNo=144
rlabel pdiffusion 241 -2787 241 -2787 0 feedthrough
rlabel pdiffusion 248 -2787 248 -2787 0 feedthrough
rlabel pdiffusion 255 -2787 255 -2787 0 feedthrough
rlabel pdiffusion 262 -2787 262 -2787 0 cellNo=792
rlabel pdiffusion 269 -2787 269 -2787 0 feedthrough
rlabel pdiffusion 276 -2787 276 -2787 0 feedthrough
rlabel pdiffusion 283 -2787 283 -2787 0 cellNo=874
rlabel pdiffusion 290 -2787 290 -2787 0 cellNo=643
rlabel pdiffusion 297 -2787 297 -2787 0 feedthrough
rlabel pdiffusion 304 -2787 304 -2787 0 feedthrough
rlabel pdiffusion 311 -2787 311 -2787 0 feedthrough
rlabel pdiffusion 318 -2787 318 -2787 0 feedthrough
rlabel pdiffusion 325 -2787 325 -2787 0 feedthrough
rlabel pdiffusion 332 -2787 332 -2787 0 feedthrough
rlabel pdiffusion 339 -2787 339 -2787 0 feedthrough
rlabel pdiffusion 346 -2787 346 -2787 0 feedthrough
rlabel pdiffusion 353 -2787 353 -2787 0 feedthrough
rlabel pdiffusion 360 -2787 360 -2787 0 feedthrough
rlabel pdiffusion 367 -2787 367 -2787 0 feedthrough
rlabel pdiffusion 374 -2787 374 -2787 0 feedthrough
rlabel pdiffusion 381 -2787 381 -2787 0 feedthrough
rlabel pdiffusion 388 -2787 388 -2787 0 feedthrough
rlabel pdiffusion 395 -2787 395 -2787 0 feedthrough
rlabel pdiffusion 402 -2787 402 -2787 0 feedthrough
rlabel pdiffusion 409 -2787 409 -2787 0 feedthrough
rlabel pdiffusion 416 -2787 416 -2787 0 feedthrough
rlabel pdiffusion 423 -2787 423 -2787 0 feedthrough
rlabel pdiffusion 430 -2787 430 -2787 0 feedthrough
rlabel pdiffusion 437 -2787 437 -2787 0 feedthrough
rlabel pdiffusion 444 -2787 444 -2787 0 cellNo=973
rlabel pdiffusion 451 -2787 451 -2787 0 feedthrough
rlabel pdiffusion 458 -2787 458 -2787 0 feedthrough
rlabel pdiffusion 465 -2787 465 -2787 0 feedthrough
rlabel pdiffusion 472 -2787 472 -2787 0 feedthrough
rlabel pdiffusion 479 -2787 479 -2787 0 cellNo=128
rlabel pdiffusion 486 -2787 486 -2787 0 feedthrough
rlabel pdiffusion 493 -2787 493 -2787 0 feedthrough
rlabel pdiffusion 500 -2787 500 -2787 0 feedthrough
rlabel pdiffusion 507 -2787 507 -2787 0 feedthrough
rlabel pdiffusion 514 -2787 514 -2787 0 feedthrough
rlabel pdiffusion 521 -2787 521 -2787 0 feedthrough
rlabel pdiffusion 528 -2787 528 -2787 0 feedthrough
rlabel pdiffusion 535 -2787 535 -2787 0 feedthrough
rlabel pdiffusion 542 -2787 542 -2787 0 feedthrough
rlabel pdiffusion 549 -2787 549 -2787 0 feedthrough
rlabel pdiffusion 556 -2787 556 -2787 0 feedthrough
rlabel pdiffusion 563 -2787 563 -2787 0 cellNo=383
rlabel pdiffusion 570 -2787 570 -2787 0 feedthrough
rlabel pdiffusion 577 -2787 577 -2787 0 feedthrough
rlabel pdiffusion 584 -2787 584 -2787 0 feedthrough
rlabel pdiffusion 591 -2787 591 -2787 0 cellNo=97
rlabel pdiffusion 598 -2787 598 -2787 0 feedthrough
rlabel pdiffusion 605 -2787 605 -2787 0 feedthrough
rlabel pdiffusion 612 -2787 612 -2787 0 feedthrough
rlabel pdiffusion 619 -2787 619 -2787 0 feedthrough
rlabel pdiffusion 626 -2787 626 -2787 0 feedthrough
rlabel pdiffusion 633 -2787 633 -2787 0 feedthrough
rlabel pdiffusion 640 -2787 640 -2787 0 feedthrough
rlabel pdiffusion 647 -2787 647 -2787 0 feedthrough
rlabel pdiffusion 654 -2787 654 -2787 0 feedthrough
rlabel pdiffusion 661 -2787 661 -2787 0 cellNo=274
rlabel pdiffusion 668 -2787 668 -2787 0 cellNo=100
rlabel pdiffusion 675 -2787 675 -2787 0 cellNo=635
rlabel pdiffusion 682 -2787 682 -2787 0 feedthrough
rlabel pdiffusion 689 -2787 689 -2787 0 cellNo=441
rlabel pdiffusion 696 -2787 696 -2787 0 feedthrough
rlabel pdiffusion 703 -2787 703 -2787 0 feedthrough
rlabel pdiffusion 710 -2787 710 -2787 0 feedthrough
rlabel pdiffusion 717 -2787 717 -2787 0 feedthrough
rlabel pdiffusion 724 -2787 724 -2787 0 feedthrough
rlabel pdiffusion 731 -2787 731 -2787 0 feedthrough
rlabel pdiffusion 738 -2787 738 -2787 0 feedthrough
rlabel pdiffusion 745 -2787 745 -2787 0 cellNo=226
rlabel pdiffusion 752 -2787 752 -2787 0 feedthrough
rlabel pdiffusion 759 -2787 759 -2787 0 cellNo=189
rlabel pdiffusion 766 -2787 766 -2787 0 feedthrough
rlabel pdiffusion 773 -2787 773 -2787 0 feedthrough
rlabel pdiffusion 780 -2787 780 -2787 0 cellNo=153
rlabel pdiffusion 787 -2787 787 -2787 0 cellNo=419
rlabel pdiffusion 794 -2787 794 -2787 0 feedthrough
rlabel pdiffusion 801 -2787 801 -2787 0 feedthrough
rlabel pdiffusion 808 -2787 808 -2787 0 cellNo=845
rlabel pdiffusion 815 -2787 815 -2787 0 cellNo=927
rlabel pdiffusion 822 -2787 822 -2787 0 feedthrough
rlabel pdiffusion 829 -2787 829 -2787 0 feedthrough
rlabel pdiffusion 836 -2787 836 -2787 0 feedthrough
rlabel pdiffusion 843 -2787 843 -2787 0 cellNo=954
rlabel pdiffusion 850 -2787 850 -2787 0 feedthrough
rlabel pdiffusion 857 -2787 857 -2787 0 feedthrough
rlabel pdiffusion 864 -2787 864 -2787 0 feedthrough
rlabel pdiffusion 871 -2787 871 -2787 0 feedthrough
rlabel pdiffusion 878 -2787 878 -2787 0 cellNo=328
rlabel pdiffusion 885 -2787 885 -2787 0 feedthrough
rlabel pdiffusion 892 -2787 892 -2787 0 feedthrough
rlabel pdiffusion 899 -2787 899 -2787 0 feedthrough
rlabel pdiffusion 906 -2787 906 -2787 0 cellNo=567
rlabel pdiffusion 913 -2787 913 -2787 0 feedthrough
rlabel pdiffusion 920 -2787 920 -2787 0 feedthrough
rlabel pdiffusion 927 -2787 927 -2787 0 feedthrough
rlabel pdiffusion 934 -2787 934 -2787 0 feedthrough
rlabel pdiffusion 941 -2787 941 -2787 0 feedthrough
rlabel pdiffusion 948 -2787 948 -2787 0 feedthrough
rlabel pdiffusion 955 -2787 955 -2787 0 feedthrough
rlabel pdiffusion 962 -2787 962 -2787 0 feedthrough
rlabel pdiffusion 969 -2787 969 -2787 0 feedthrough
rlabel pdiffusion 976 -2787 976 -2787 0 feedthrough
rlabel pdiffusion 983 -2787 983 -2787 0 feedthrough
rlabel pdiffusion 990 -2787 990 -2787 0 feedthrough
rlabel pdiffusion 997 -2787 997 -2787 0 feedthrough
rlabel pdiffusion 1004 -2787 1004 -2787 0 cellNo=574
rlabel pdiffusion 1011 -2787 1011 -2787 0 feedthrough
rlabel pdiffusion 1018 -2787 1018 -2787 0 feedthrough
rlabel pdiffusion 1025 -2787 1025 -2787 0 feedthrough
rlabel pdiffusion 1032 -2787 1032 -2787 0 feedthrough
rlabel pdiffusion 1039 -2787 1039 -2787 0 feedthrough
rlabel pdiffusion 1046 -2787 1046 -2787 0 feedthrough
rlabel pdiffusion 1053 -2787 1053 -2787 0 feedthrough
rlabel pdiffusion 1060 -2787 1060 -2787 0 feedthrough
rlabel pdiffusion 1067 -2787 1067 -2787 0 feedthrough
rlabel pdiffusion 1074 -2787 1074 -2787 0 feedthrough
rlabel pdiffusion 1081 -2787 1081 -2787 0 feedthrough
rlabel pdiffusion 1088 -2787 1088 -2787 0 feedthrough
rlabel pdiffusion 1095 -2787 1095 -2787 0 feedthrough
rlabel pdiffusion 1102 -2787 1102 -2787 0 feedthrough
rlabel pdiffusion 1109 -2787 1109 -2787 0 feedthrough
rlabel pdiffusion 1116 -2787 1116 -2787 0 feedthrough
rlabel pdiffusion 1123 -2787 1123 -2787 0 feedthrough
rlabel pdiffusion 1130 -2787 1130 -2787 0 feedthrough
rlabel pdiffusion 1137 -2787 1137 -2787 0 feedthrough
rlabel pdiffusion 1144 -2787 1144 -2787 0 feedthrough
rlabel pdiffusion 1151 -2787 1151 -2787 0 feedthrough
rlabel pdiffusion 1158 -2787 1158 -2787 0 cellNo=676
rlabel pdiffusion 1165 -2787 1165 -2787 0 feedthrough
rlabel pdiffusion 1172 -2787 1172 -2787 0 feedthrough
rlabel pdiffusion 1179 -2787 1179 -2787 0 feedthrough
rlabel pdiffusion 1186 -2787 1186 -2787 0 cellNo=895
rlabel pdiffusion 1193 -2787 1193 -2787 0 feedthrough
rlabel pdiffusion 1200 -2787 1200 -2787 0 feedthrough
rlabel pdiffusion 1207 -2787 1207 -2787 0 feedthrough
rlabel pdiffusion 1214 -2787 1214 -2787 0 feedthrough
rlabel pdiffusion 1221 -2787 1221 -2787 0 feedthrough
rlabel pdiffusion 1228 -2787 1228 -2787 0 feedthrough
rlabel pdiffusion 1235 -2787 1235 -2787 0 feedthrough
rlabel pdiffusion 1242 -2787 1242 -2787 0 feedthrough
rlabel pdiffusion 1249 -2787 1249 -2787 0 feedthrough
rlabel pdiffusion 1256 -2787 1256 -2787 0 feedthrough
rlabel pdiffusion 1263 -2787 1263 -2787 0 feedthrough
rlabel pdiffusion 1270 -2787 1270 -2787 0 feedthrough
rlabel pdiffusion 1277 -2787 1277 -2787 0 feedthrough
rlabel pdiffusion 1284 -2787 1284 -2787 0 feedthrough
rlabel pdiffusion 1291 -2787 1291 -2787 0 feedthrough
rlabel pdiffusion 1298 -2787 1298 -2787 0 cellNo=319
rlabel pdiffusion 1305 -2787 1305 -2787 0 feedthrough
rlabel pdiffusion 1312 -2787 1312 -2787 0 feedthrough
rlabel pdiffusion 1319 -2787 1319 -2787 0 feedthrough
rlabel pdiffusion 1326 -2787 1326 -2787 0 feedthrough
rlabel pdiffusion 1333 -2787 1333 -2787 0 feedthrough
rlabel pdiffusion 1340 -2787 1340 -2787 0 feedthrough
rlabel pdiffusion 1347 -2787 1347 -2787 0 feedthrough
rlabel pdiffusion 1354 -2787 1354 -2787 0 feedthrough
rlabel pdiffusion 1361 -2787 1361 -2787 0 feedthrough
rlabel pdiffusion 1368 -2787 1368 -2787 0 feedthrough
rlabel pdiffusion 1375 -2787 1375 -2787 0 feedthrough
rlabel pdiffusion 1382 -2787 1382 -2787 0 feedthrough
rlabel pdiffusion 1389 -2787 1389 -2787 0 feedthrough
rlabel pdiffusion 1396 -2787 1396 -2787 0 feedthrough
rlabel pdiffusion 1403 -2787 1403 -2787 0 feedthrough
rlabel pdiffusion 1410 -2787 1410 -2787 0 feedthrough
rlabel pdiffusion 1417 -2787 1417 -2787 0 feedthrough
rlabel pdiffusion 1424 -2787 1424 -2787 0 feedthrough
rlabel pdiffusion 1431 -2787 1431 -2787 0 feedthrough
rlabel pdiffusion 1438 -2787 1438 -2787 0 feedthrough
rlabel pdiffusion 1445 -2787 1445 -2787 0 feedthrough
rlabel pdiffusion 1452 -2787 1452 -2787 0 feedthrough
rlabel pdiffusion 1459 -2787 1459 -2787 0 feedthrough
rlabel pdiffusion 1466 -2787 1466 -2787 0 feedthrough
rlabel pdiffusion 1473 -2787 1473 -2787 0 feedthrough
rlabel pdiffusion 1480 -2787 1480 -2787 0 feedthrough
rlabel pdiffusion 1487 -2787 1487 -2787 0 feedthrough
rlabel pdiffusion 1494 -2787 1494 -2787 0 feedthrough
rlabel pdiffusion 1501 -2787 1501 -2787 0 feedthrough
rlabel pdiffusion 1508 -2787 1508 -2787 0 feedthrough
rlabel pdiffusion 1515 -2787 1515 -2787 0 feedthrough
rlabel pdiffusion 1522 -2787 1522 -2787 0 cellNo=901
rlabel pdiffusion 3 -2912 3 -2912 0 cellNo=1043
rlabel pdiffusion 10 -2912 10 -2912 0 cellNo=1046
rlabel pdiffusion 17 -2912 17 -2912 0 cellNo=1050
rlabel pdiffusion 24 -2912 24 -2912 0 cellNo=1056
rlabel pdiffusion 31 -2912 31 -2912 0 cellNo=1061
rlabel pdiffusion 38 -2912 38 -2912 0 cellNo=1064
rlabel pdiffusion 45 -2912 45 -2912 0 cellNo=1068
rlabel pdiffusion 52 -2912 52 -2912 0 cellNo=1070
rlabel pdiffusion 59 -2912 59 -2912 0 cellNo=1072
rlabel pdiffusion 66 -2912 66 -2912 0 cellNo=1074
rlabel pdiffusion 73 -2912 73 -2912 0 feedthrough
rlabel pdiffusion 80 -2912 80 -2912 0 feedthrough
rlabel pdiffusion 87 -2912 87 -2912 0 feedthrough
rlabel pdiffusion 94 -2912 94 -2912 0 feedthrough
rlabel pdiffusion 101 -2912 101 -2912 0 cellNo=887
rlabel pdiffusion 108 -2912 108 -2912 0 feedthrough
rlabel pdiffusion 115 -2912 115 -2912 0 feedthrough
rlabel pdiffusion 122 -2912 122 -2912 0 cellNo=499
rlabel pdiffusion 129 -2912 129 -2912 0 feedthrough
rlabel pdiffusion 136 -2912 136 -2912 0 feedthrough
rlabel pdiffusion 143 -2912 143 -2912 0 cellNo=402
rlabel pdiffusion 150 -2912 150 -2912 0 feedthrough
rlabel pdiffusion 157 -2912 157 -2912 0 feedthrough
rlabel pdiffusion 164 -2912 164 -2912 0 feedthrough
rlabel pdiffusion 171 -2912 171 -2912 0 feedthrough
rlabel pdiffusion 178 -2912 178 -2912 0 feedthrough
rlabel pdiffusion 185 -2912 185 -2912 0 feedthrough
rlabel pdiffusion 192 -2912 192 -2912 0 feedthrough
rlabel pdiffusion 199 -2912 199 -2912 0 feedthrough
rlabel pdiffusion 206 -2912 206 -2912 0 cellNo=952
rlabel pdiffusion 213 -2912 213 -2912 0 feedthrough
rlabel pdiffusion 220 -2912 220 -2912 0 feedthrough
rlabel pdiffusion 227 -2912 227 -2912 0 cellNo=288
rlabel pdiffusion 234 -2912 234 -2912 0 feedthrough
rlabel pdiffusion 241 -2912 241 -2912 0 feedthrough
rlabel pdiffusion 248 -2912 248 -2912 0 cellNo=827
rlabel pdiffusion 255 -2912 255 -2912 0 feedthrough
rlabel pdiffusion 262 -2912 262 -2912 0 feedthrough
rlabel pdiffusion 269 -2912 269 -2912 0 feedthrough
rlabel pdiffusion 276 -2912 276 -2912 0 cellNo=541
rlabel pdiffusion 283 -2912 283 -2912 0 cellNo=145
rlabel pdiffusion 290 -2912 290 -2912 0 cellNo=218
rlabel pdiffusion 297 -2912 297 -2912 0 feedthrough
rlabel pdiffusion 304 -2912 304 -2912 0 feedthrough
rlabel pdiffusion 311 -2912 311 -2912 0 feedthrough
rlabel pdiffusion 318 -2912 318 -2912 0 feedthrough
rlabel pdiffusion 325 -2912 325 -2912 0 feedthrough
rlabel pdiffusion 332 -2912 332 -2912 0 feedthrough
rlabel pdiffusion 339 -2912 339 -2912 0 feedthrough
rlabel pdiffusion 346 -2912 346 -2912 0 feedthrough
rlabel pdiffusion 353 -2912 353 -2912 0 feedthrough
rlabel pdiffusion 360 -2912 360 -2912 0 feedthrough
rlabel pdiffusion 367 -2912 367 -2912 0 feedthrough
rlabel pdiffusion 374 -2912 374 -2912 0 feedthrough
rlabel pdiffusion 381 -2912 381 -2912 0 feedthrough
rlabel pdiffusion 388 -2912 388 -2912 0 feedthrough
rlabel pdiffusion 395 -2912 395 -2912 0 feedthrough
rlabel pdiffusion 402 -2912 402 -2912 0 feedthrough
rlabel pdiffusion 409 -2912 409 -2912 0 feedthrough
rlabel pdiffusion 416 -2912 416 -2912 0 feedthrough
rlabel pdiffusion 423 -2912 423 -2912 0 feedthrough
rlabel pdiffusion 430 -2912 430 -2912 0 feedthrough
rlabel pdiffusion 437 -2912 437 -2912 0 feedthrough
rlabel pdiffusion 444 -2912 444 -2912 0 feedthrough
rlabel pdiffusion 451 -2912 451 -2912 0 feedthrough
rlabel pdiffusion 458 -2912 458 -2912 0 feedthrough
rlabel pdiffusion 465 -2912 465 -2912 0 feedthrough
rlabel pdiffusion 472 -2912 472 -2912 0 feedthrough
rlabel pdiffusion 479 -2912 479 -2912 0 feedthrough
rlabel pdiffusion 486 -2912 486 -2912 0 feedthrough
rlabel pdiffusion 493 -2912 493 -2912 0 cellNo=573
rlabel pdiffusion 500 -2912 500 -2912 0 feedthrough
rlabel pdiffusion 507 -2912 507 -2912 0 feedthrough
rlabel pdiffusion 514 -2912 514 -2912 0 feedthrough
rlabel pdiffusion 521 -2912 521 -2912 0 feedthrough
rlabel pdiffusion 528 -2912 528 -2912 0 feedthrough
rlabel pdiffusion 535 -2912 535 -2912 0 feedthrough
rlabel pdiffusion 542 -2912 542 -2912 0 feedthrough
rlabel pdiffusion 549 -2912 549 -2912 0 feedthrough
rlabel pdiffusion 556 -2912 556 -2912 0 cellNo=22
rlabel pdiffusion 563 -2912 563 -2912 0 feedthrough
rlabel pdiffusion 570 -2912 570 -2912 0 feedthrough
rlabel pdiffusion 577 -2912 577 -2912 0 feedthrough
rlabel pdiffusion 584 -2912 584 -2912 0 cellNo=751
rlabel pdiffusion 591 -2912 591 -2912 0 feedthrough
rlabel pdiffusion 598 -2912 598 -2912 0 feedthrough
rlabel pdiffusion 605 -2912 605 -2912 0 feedthrough
rlabel pdiffusion 612 -2912 612 -2912 0 feedthrough
rlabel pdiffusion 619 -2912 619 -2912 0 feedthrough
rlabel pdiffusion 626 -2912 626 -2912 0 feedthrough
rlabel pdiffusion 633 -2912 633 -2912 0 feedthrough
rlabel pdiffusion 640 -2912 640 -2912 0 cellNo=366
rlabel pdiffusion 647 -2912 647 -2912 0 feedthrough
rlabel pdiffusion 654 -2912 654 -2912 0 feedthrough
rlabel pdiffusion 661 -2912 661 -2912 0 cellNo=457
rlabel pdiffusion 668 -2912 668 -2912 0 feedthrough
rlabel pdiffusion 675 -2912 675 -2912 0 feedthrough
rlabel pdiffusion 682 -2912 682 -2912 0 feedthrough
rlabel pdiffusion 689 -2912 689 -2912 0 feedthrough
rlabel pdiffusion 696 -2912 696 -2912 0 feedthrough
rlabel pdiffusion 703 -2912 703 -2912 0 cellNo=89
rlabel pdiffusion 710 -2912 710 -2912 0 feedthrough
rlabel pdiffusion 717 -2912 717 -2912 0 feedthrough
rlabel pdiffusion 724 -2912 724 -2912 0 feedthrough
rlabel pdiffusion 731 -2912 731 -2912 0 feedthrough
rlabel pdiffusion 738 -2912 738 -2912 0 feedthrough
rlabel pdiffusion 745 -2912 745 -2912 0 cellNo=875
rlabel pdiffusion 752 -2912 752 -2912 0 feedthrough
rlabel pdiffusion 759 -2912 759 -2912 0 cellNo=851
rlabel pdiffusion 766 -2912 766 -2912 0 feedthrough
rlabel pdiffusion 773 -2912 773 -2912 0 feedthrough
rlabel pdiffusion 780 -2912 780 -2912 0 feedthrough
rlabel pdiffusion 787 -2912 787 -2912 0 feedthrough
rlabel pdiffusion 794 -2912 794 -2912 0 feedthrough
rlabel pdiffusion 801 -2912 801 -2912 0 feedthrough
rlabel pdiffusion 808 -2912 808 -2912 0 feedthrough
rlabel pdiffusion 815 -2912 815 -2912 0 feedthrough
rlabel pdiffusion 822 -2912 822 -2912 0 cellNo=817
rlabel pdiffusion 829 -2912 829 -2912 0 feedthrough
rlabel pdiffusion 836 -2912 836 -2912 0 cellNo=535
rlabel pdiffusion 843 -2912 843 -2912 0 cellNo=229
rlabel pdiffusion 850 -2912 850 -2912 0 feedthrough
rlabel pdiffusion 857 -2912 857 -2912 0 feedthrough
rlabel pdiffusion 864 -2912 864 -2912 0 cellNo=629
rlabel pdiffusion 871 -2912 871 -2912 0 feedthrough
rlabel pdiffusion 878 -2912 878 -2912 0 feedthrough
rlabel pdiffusion 885 -2912 885 -2912 0 feedthrough
rlabel pdiffusion 892 -2912 892 -2912 0 feedthrough
rlabel pdiffusion 899 -2912 899 -2912 0 feedthrough
rlabel pdiffusion 906 -2912 906 -2912 0 feedthrough
rlabel pdiffusion 913 -2912 913 -2912 0 cellNo=349
rlabel pdiffusion 920 -2912 920 -2912 0 cellNo=194
rlabel pdiffusion 927 -2912 927 -2912 0 feedthrough
rlabel pdiffusion 934 -2912 934 -2912 0 feedthrough
rlabel pdiffusion 941 -2912 941 -2912 0 feedthrough
rlabel pdiffusion 948 -2912 948 -2912 0 cellNo=197
rlabel pdiffusion 955 -2912 955 -2912 0 cellNo=963
rlabel pdiffusion 962 -2912 962 -2912 0 feedthrough
rlabel pdiffusion 969 -2912 969 -2912 0 feedthrough
rlabel pdiffusion 976 -2912 976 -2912 0 feedthrough
rlabel pdiffusion 983 -2912 983 -2912 0 feedthrough
rlabel pdiffusion 990 -2912 990 -2912 0 feedthrough
rlabel pdiffusion 997 -2912 997 -2912 0 feedthrough
rlabel pdiffusion 1004 -2912 1004 -2912 0 feedthrough
rlabel pdiffusion 1011 -2912 1011 -2912 0 feedthrough
rlabel pdiffusion 1018 -2912 1018 -2912 0 cellNo=68
rlabel pdiffusion 1025 -2912 1025 -2912 0 feedthrough
rlabel pdiffusion 1032 -2912 1032 -2912 0 feedthrough
rlabel pdiffusion 1039 -2912 1039 -2912 0 feedthrough
rlabel pdiffusion 1046 -2912 1046 -2912 0 feedthrough
rlabel pdiffusion 1053 -2912 1053 -2912 0 feedthrough
rlabel pdiffusion 1060 -2912 1060 -2912 0 feedthrough
rlabel pdiffusion 1067 -2912 1067 -2912 0 feedthrough
rlabel pdiffusion 1074 -2912 1074 -2912 0 feedthrough
rlabel pdiffusion 1081 -2912 1081 -2912 0 feedthrough
rlabel pdiffusion 1088 -2912 1088 -2912 0 feedthrough
rlabel pdiffusion 1095 -2912 1095 -2912 0 cellNo=994
rlabel pdiffusion 1102 -2912 1102 -2912 0 feedthrough
rlabel pdiffusion 1109 -2912 1109 -2912 0 feedthrough
rlabel pdiffusion 1116 -2912 1116 -2912 0 feedthrough
rlabel pdiffusion 1123 -2912 1123 -2912 0 feedthrough
rlabel pdiffusion 1130 -2912 1130 -2912 0 feedthrough
rlabel pdiffusion 1137 -2912 1137 -2912 0 feedthrough
rlabel pdiffusion 1144 -2912 1144 -2912 0 feedthrough
rlabel pdiffusion 1151 -2912 1151 -2912 0 feedthrough
rlabel pdiffusion 1158 -2912 1158 -2912 0 feedthrough
rlabel pdiffusion 1165 -2912 1165 -2912 0 feedthrough
rlabel pdiffusion 1172 -2912 1172 -2912 0 feedthrough
rlabel pdiffusion 1179 -2912 1179 -2912 0 feedthrough
rlabel pdiffusion 1186 -2912 1186 -2912 0 feedthrough
rlabel pdiffusion 1193 -2912 1193 -2912 0 feedthrough
rlabel pdiffusion 1200 -2912 1200 -2912 0 feedthrough
rlabel pdiffusion 1207 -2912 1207 -2912 0 feedthrough
rlabel pdiffusion 1214 -2912 1214 -2912 0 feedthrough
rlabel pdiffusion 1221 -2912 1221 -2912 0 feedthrough
rlabel pdiffusion 1228 -2912 1228 -2912 0 feedthrough
rlabel pdiffusion 1235 -2912 1235 -2912 0 feedthrough
rlabel pdiffusion 1242 -2912 1242 -2912 0 feedthrough
rlabel pdiffusion 1249 -2912 1249 -2912 0 feedthrough
rlabel pdiffusion 1256 -2912 1256 -2912 0 feedthrough
rlabel pdiffusion 1263 -2912 1263 -2912 0 feedthrough
rlabel pdiffusion 1270 -2912 1270 -2912 0 feedthrough
rlabel pdiffusion 1277 -2912 1277 -2912 0 feedthrough
rlabel pdiffusion 1284 -2912 1284 -2912 0 feedthrough
rlabel pdiffusion 1291 -2912 1291 -2912 0 feedthrough
rlabel pdiffusion 1298 -2912 1298 -2912 0 feedthrough
rlabel pdiffusion 1305 -2912 1305 -2912 0 feedthrough
rlabel pdiffusion 1312 -2912 1312 -2912 0 feedthrough
rlabel pdiffusion 1319 -2912 1319 -2912 0 feedthrough
rlabel pdiffusion 1326 -2912 1326 -2912 0 feedthrough
rlabel pdiffusion 1333 -2912 1333 -2912 0 feedthrough
rlabel pdiffusion 1340 -2912 1340 -2912 0 feedthrough
rlabel pdiffusion 1347 -2912 1347 -2912 0 feedthrough
rlabel pdiffusion 1354 -2912 1354 -2912 0 feedthrough
rlabel pdiffusion 1361 -2912 1361 -2912 0 cellNo=997
rlabel pdiffusion 1368 -2912 1368 -2912 0 feedthrough
rlabel pdiffusion 1375 -2912 1375 -2912 0 feedthrough
rlabel pdiffusion 1382 -2912 1382 -2912 0 feedthrough
rlabel pdiffusion 1389 -2912 1389 -2912 0 feedthrough
rlabel pdiffusion 1396 -2912 1396 -2912 0 feedthrough
rlabel pdiffusion 1403 -2912 1403 -2912 0 feedthrough
rlabel pdiffusion 1410 -2912 1410 -2912 0 feedthrough
rlabel pdiffusion 1417 -2912 1417 -2912 0 feedthrough
rlabel pdiffusion 1424 -2912 1424 -2912 0 feedthrough
rlabel pdiffusion 1431 -2912 1431 -2912 0 feedthrough
rlabel pdiffusion 3 -3031 3 -3031 0 cellNo=1051
rlabel pdiffusion 10 -3031 10 -3031 0 cellNo=1052
rlabel pdiffusion 17 -3031 17 -3031 0 cellNo=1055
rlabel pdiffusion 24 -3031 24 -3031 0 cellNo=1060
rlabel pdiffusion 31 -3031 31 -3031 0 cellNo=1063
rlabel pdiffusion 38 -3031 38 -3031 0 cellNo=1065
rlabel pdiffusion 45 -3031 45 -3031 0 cellNo=1069
rlabel pdiffusion 52 -3031 52 -3031 0 cellNo=1071
rlabel pdiffusion 59 -3031 59 -3031 0 cellNo=1073
rlabel pdiffusion 66 -3031 66 -3031 0 cellNo=1076
rlabel pdiffusion 73 -3031 73 -3031 0 cellNo=1079
rlabel pdiffusion 80 -3031 80 -3031 0 cellNo=1084
rlabel pdiffusion 87 -3031 87 -3031 0 feedthrough
rlabel pdiffusion 94 -3031 94 -3031 0 feedthrough
rlabel pdiffusion 101 -3031 101 -3031 0 feedthrough
rlabel pdiffusion 108 -3031 108 -3031 0 feedthrough
rlabel pdiffusion 115 -3031 115 -3031 0 feedthrough
rlabel pdiffusion 122 -3031 122 -3031 0 feedthrough
rlabel pdiffusion 129 -3031 129 -3031 0 feedthrough
rlabel pdiffusion 136 -3031 136 -3031 0 feedthrough
rlabel pdiffusion 143 -3031 143 -3031 0 feedthrough
rlabel pdiffusion 150 -3031 150 -3031 0 cellNo=675
rlabel pdiffusion 157 -3031 157 -3031 0 feedthrough
rlabel pdiffusion 164 -3031 164 -3031 0 cellNo=86
rlabel pdiffusion 171 -3031 171 -3031 0 feedthrough
rlabel pdiffusion 178 -3031 178 -3031 0 feedthrough
rlabel pdiffusion 185 -3031 185 -3031 0 feedthrough
rlabel pdiffusion 192 -3031 192 -3031 0 feedthrough
rlabel pdiffusion 199 -3031 199 -3031 0 feedthrough
rlabel pdiffusion 206 -3031 206 -3031 0 cellNo=467
rlabel pdiffusion 213 -3031 213 -3031 0 feedthrough
rlabel pdiffusion 220 -3031 220 -3031 0 cellNo=241
rlabel pdiffusion 227 -3031 227 -3031 0 feedthrough
rlabel pdiffusion 234 -3031 234 -3031 0 feedthrough
rlabel pdiffusion 241 -3031 241 -3031 0 feedthrough
rlabel pdiffusion 248 -3031 248 -3031 0 cellNo=696
rlabel pdiffusion 255 -3031 255 -3031 0 feedthrough
rlabel pdiffusion 262 -3031 262 -3031 0 cellNo=416
rlabel pdiffusion 269 -3031 269 -3031 0 feedthrough
rlabel pdiffusion 276 -3031 276 -3031 0 feedthrough
rlabel pdiffusion 283 -3031 283 -3031 0 feedthrough
rlabel pdiffusion 290 -3031 290 -3031 0 feedthrough
rlabel pdiffusion 297 -3031 297 -3031 0 feedthrough
rlabel pdiffusion 304 -3031 304 -3031 0 feedthrough
rlabel pdiffusion 311 -3031 311 -3031 0 feedthrough
rlabel pdiffusion 318 -3031 318 -3031 0 feedthrough
rlabel pdiffusion 325 -3031 325 -3031 0 feedthrough
rlabel pdiffusion 332 -3031 332 -3031 0 feedthrough
rlabel pdiffusion 339 -3031 339 -3031 0 feedthrough
rlabel pdiffusion 346 -3031 346 -3031 0 feedthrough
rlabel pdiffusion 353 -3031 353 -3031 0 feedthrough
rlabel pdiffusion 360 -3031 360 -3031 0 feedthrough
rlabel pdiffusion 367 -3031 367 -3031 0 feedthrough
rlabel pdiffusion 374 -3031 374 -3031 0 feedthrough
rlabel pdiffusion 381 -3031 381 -3031 0 feedthrough
rlabel pdiffusion 388 -3031 388 -3031 0 feedthrough
rlabel pdiffusion 395 -3031 395 -3031 0 feedthrough
rlabel pdiffusion 402 -3031 402 -3031 0 feedthrough
rlabel pdiffusion 409 -3031 409 -3031 0 cellNo=444
rlabel pdiffusion 416 -3031 416 -3031 0 feedthrough
rlabel pdiffusion 423 -3031 423 -3031 0 feedthrough
rlabel pdiffusion 430 -3031 430 -3031 0 feedthrough
rlabel pdiffusion 437 -3031 437 -3031 0 feedthrough
rlabel pdiffusion 444 -3031 444 -3031 0 feedthrough
rlabel pdiffusion 451 -3031 451 -3031 0 feedthrough
rlabel pdiffusion 458 -3031 458 -3031 0 feedthrough
rlabel pdiffusion 465 -3031 465 -3031 0 feedthrough
rlabel pdiffusion 472 -3031 472 -3031 0 feedthrough
rlabel pdiffusion 479 -3031 479 -3031 0 feedthrough
rlabel pdiffusion 486 -3031 486 -3031 0 feedthrough
rlabel pdiffusion 493 -3031 493 -3031 0 feedthrough
rlabel pdiffusion 500 -3031 500 -3031 0 feedthrough
rlabel pdiffusion 507 -3031 507 -3031 0 cellNo=702
rlabel pdiffusion 514 -3031 514 -3031 0 feedthrough
rlabel pdiffusion 521 -3031 521 -3031 0 feedthrough
rlabel pdiffusion 528 -3031 528 -3031 0 feedthrough
rlabel pdiffusion 535 -3031 535 -3031 0 feedthrough
rlabel pdiffusion 542 -3031 542 -3031 0 feedthrough
rlabel pdiffusion 549 -3031 549 -3031 0 feedthrough
rlabel pdiffusion 556 -3031 556 -3031 0 feedthrough
rlabel pdiffusion 563 -3031 563 -3031 0 feedthrough
rlabel pdiffusion 570 -3031 570 -3031 0 feedthrough
rlabel pdiffusion 577 -3031 577 -3031 0 feedthrough
rlabel pdiffusion 584 -3031 584 -3031 0 feedthrough
rlabel pdiffusion 591 -3031 591 -3031 0 feedthrough
rlabel pdiffusion 598 -3031 598 -3031 0 feedthrough
rlabel pdiffusion 605 -3031 605 -3031 0 feedthrough
rlabel pdiffusion 612 -3031 612 -3031 0 feedthrough
rlabel pdiffusion 619 -3031 619 -3031 0 feedthrough
rlabel pdiffusion 626 -3031 626 -3031 0 feedthrough
rlabel pdiffusion 633 -3031 633 -3031 0 cellNo=638
rlabel pdiffusion 640 -3031 640 -3031 0 feedthrough
rlabel pdiffusion 647 -3031 647 -3031 0 cellNo=872
rlabel pdiffusion 654 -3031 654 -3031 0 feedthrough
rlabel pdiffusion 661 -3031 661 -3031 0 cellNo=79
rlabel pdiffusion 668 -3031 668 -3031 0 feedthrough
rlabel pdiffusion 675 -3031 675 -3031 0 feedthrough
rlabel pdiffusion 682 -3031 682 -3031 0 feedthrough
rlabel pdiffusion 689 -3031 689 -3031 0 cellNo=990
rlabel pdiffusion 696 -3031 696 -3031 0 cellNo=289
rlabel pdiffusion 703 -3031 703 -3031 0 feedthrough
rlabel pdiffusion 710 -3031 710 -3031 0 feedthrough
rlabel pdiffusion 717 -3031 717 -3031 0 feedthrough
rlabel pdiffusion 724 -3031 724 -3031 0 feedthrough
rlabel pdiffusion 731 -3031 731 -3031 0 feedthrough
rlabel pdiffusion 738 -3031 738 -3031 0 feedthrough
rlabel pdiffusion 745 -3031 745 -3031 0 feedthrough
rlabel pdiffusion 752 -3031 752 -3031 0 cellNo=547
rlabel pdiffusion 759 -3031 759 -3031 0 feedthrough
rlabel pdiffusion 766 -3031 766 -3031 0 cellNo=988
rlabel pdiffusion 773 -3031 773 -3031 0 feedthrough
rlabel pdiffusion 780 -3031 780 -3031 0 feedthrough
rlabel pdiffusion 787 -3031 787 -3031 0 cellNo=723
rlabel pdiffusion 794 -3031 794 -3031 0 feedthrough
rlabel pdiffusion 801 -3031 801 -3031 0 feedthrough
rlabel pdiffusion 808 -3031 808 -3031 0 feedthrough
rlabel pdiffusion 815 -3031 815 -3031 0 feedthrough
rlabel pdiffusion 822 -3031 822 -3031 0 feedthrough
rlabel pdiffusion 829 -3031 829 -3031 0 feedthrough
rlabel pdiffusion 836 -3031 836 -3031 0 cellNo=896
rlabel pdiffusion 843 -3031 843 -3031 0 feedthrough
rlabel pdiffusion 850 -3031 850 -3031 0 feedthrough
rlabel pdiffusion 857 -3031 857 -3031 0 feedthrough
rlabel pdiffusion 864 -3031 864 -3031 0 cellNo=537
rlabel pdiffusion 871 -3031 871 -3031 0 cellNo=41
rlabel pdiffusion 878 -3031 878 -3031 0 feedthrough
rlabel pdiffusion 885 -3031 885 -3031 0 cellNo=151
rlabel pdiffusion 892 -3031 892 -3031 0 feedthrough
rlabel pdiffusion 899 -3031 899 -3031 0 feedthrough
rlabel pdiffusion 906 -3031 906 -3031 0 feedthrough
rlabel pdiffusion 913 -3031 913 -3031 0 cellNo=935
rlabel pdiffusion 920 -3031 920 -3031 0 cellNo=447
rlabel pdiffusion 927 -3031 927 -3031 0 feedthrough
rlabel pdiffusion 934 -3031 934 -3031 0 feedthrough
rlabel pdiffusion 941 -3031 941 -3031 0 feedthrough
rlabel pdiffusion 948 -3031 948 -3031 0 feedthrough
rlabel pdiffusion 955 -3031 955 -3031 0 feedthrough
rlabel pdiffusion 962 -3031 962 -3031 0 feedthrough
rlabel pdiffusion 969 -3031 969 -3031 0 feedthrough
rlabel pdiffusion 976 -3031 976 -3031 0 feedthrough
rlabel pdiffusion 983 -3031 983 -3031 0 feedthrough
rlabel pdiffusion 990 -3031 990 -3031 0 feedthrough
rlabel pdiffusion 997 -3031 997 -3031 0 feedthrough
rlabel pdiffusion 1004 -3031 1004 -3031 0 feedthrough
rlabel pdiffusion 1011 -3031 1011 -3031 0 feedthrough
rlabel pdiffusion 1018 -3031 1018 -3031 0 cellNo=112
rlabel pdiffusion 1025 -3031 1025 -3031 0 feedthrough
rlabel pdiffusion 1032 -3031 1032 -3031 0 feedthrough
rlabel pdiffusion 1039 -3031 1039 -3031 0 feedthrough
rlabel pdiffusion 1046 -3031 1046 -3031 0 feedthrough
rlabel pdiffusion 1053 -3031 1053 -3031 0 feedthrough
rlabel pdiffusion 1060 -3031 1060 -3031 0 feedthrough
rlabel pdiffusion 1067 -3031 1067 -3031 0 feedthrough
rlabel pdiffusion 1074 -3031 1074 -3031 0 cellNo=571
rlabel pdiffusion 1081 -3031 1081 -3031 0 feedthrough
rlabel pdiffusion 1088 -3031 1088 -3031 0 feedthrough
rlabel pdiffusion 1095 -3031 1095 -3031 0 feedthrough
rlabel pdiffusion 1102 -3031 1102 -3031 0 feedthrough
rlabel pdiffusion 1109 -3031 1109 -3031 0 feedthrough
rlabel pdiffusion 1116 -3031 1116 -3031 0 feedthrough
rlabel pdiffusion 1123 -3031 1123 -3031 0 feedthrough
rlabel pdiffusion 1130 -3031 1130 -3031 0 feedthrough
rlabel pdiffusion 1137 -3031 1137 -3031 0 feedthrough
rlabel pdiffusion 1144 -3031 1144 -3031 0 feedthrough
rlabel pdiffusion 1151 -3031 1151 -3031 0 cellNo=650
rlabel pdiffusion 1158 -3031 1158 -3031 0 feedthrough
rlabel pdiffusion 1165 -3031 1165 -3031 0 feedthrough
rlabel pdiffusion 1172 -3031 1172 -3031 0 feedthrough
rlabel pdiffusion 1179 -3031 1179 -3031 0 feedthrough
rlabel pdiffusion 1186 -3031 1186 -3031 0 feedthrough
rlabel pdiffusion 1193 -3031 1193 -3031 0 feedthrough
rlabel pdiffusion 1200 -3031 1200 -3031 0 feedthrough
rlabel pdiffusion 1207 -3031 1207 -3031 0 feedthrough
rlabel pdiffusion 1214 -3031 1214 -3031 0 feedthrough
rlabel pdiffusion 1221 -3031 1221 -3031 0 feedthrough
rlabel pdiffusion 1228 -3031 1228 -3031 0 feedthrough
rlabel pdiffusion 1235 -3031 1235 -3031 0 feedthrough
rlabel pdiffusion 1242 -3031 1242 -3031 0 feedthrough
rlabel pdiffusion 1249 -3031 1249 -3031 0 feedthrough
rlabel pdiffusion 1256 -3031 1256 -3031 0 feedthrough
rlabel pdiffusion 1263 -3031 1263 -3031 0 feedthrough
rlabel pdiffusion 1270 -3031 1270 -3031 0 feedthrough
rlabel pdiffusion 1277 -3031 1277 -3031 0 feedthrough
rlabel pdiffusion 1284 -3031 1284 -3031 0 feedthrough
rlabel pdiffusion 1291 -3031 1291 -3031 0 feedthrough
rlabel pdiffusion 1298 -3031 1298 -3031 0 feedthrough
rlabel pdiffusion 1305 -3031 1305 -3031 0 feedthrough
rlabel pdiffusion 1312 -3031 1312 -3031 0 feedthrough
rlabel pdiffusion 1319 -3031 1319 -3031 0 feedthrough
rlabel pdiffusion 1326 -3031 1326 -3031 0 feedthrough
rlabel pdiffusion 1333 -3031 1333 -3031 0 feedthrough
rlabel pdiffusion 1340 -3031 1340 -3031 0 feedthrough
rlabel pdiffusion 1347 -3031 1347 -3031 0 feedthrough
rlabel pdiffusion 1354 -3031 1354 -3031 0 feedthrough
rlabel pdiffusion 1361 -3031 1361 -3031 0 feedthrough
rlabel pdiffusion 1368 -3031 1368 -3031 0 feedthrough
rlabel pdiffusion 1375 -3031 1375 -3031 0 feedthrough
rlabel pdiffusion 1382 -3031 1382 -3031 0 feedthrough
rlabel pdiffusion 1389 -3031 1389 -3031 0 feedthrough
rlabel pdiffusion 1396 -3031 1396 -3031 0 feedthrough
rlabel pdiffusion 1403 -3031 1403 -3031 0 feedthrough
rlabel pdiffusion 1410 -3031 1410 -3031 0 feedthrough
rlabel pdiffusion 3 -3142 3 -3142 0 cellNo=1093
rlabel pdiffusion 10 -3142 10 -3142 0 cellNo=1094
rlabel pdiffusion 17 -3142 17 -3142 0 cellNo=1095
rlabel pdiffusion 24 -3142 24 -3142 0 cellNo=1096
rlabel pdiffusion 31 -3142 31 -3142 0 cellNo=1097
rlabel pdiffusion 38 -3142 38 -3142 0 cellNo=1098
rlabel pdiffusion 45 -3142 45 -3142 0 cellNo=1099
rlabel pdiffusion 52 -3142 52 -3142 0 cellNo=1100
rlabel pdiffusion 59 -3142 59 -3142 0 cellNo=1101
rlabel pdiffusion 66 -3142 66 -3142 0 cellNo=1102
rlabel pdiffusion 73 -3142 73 -3142 0 cellNo=1103
rlabel pdiffusion 80 -3142 80 -3142 0 cellNo=1104
rlabel pdiffusion 101 -3142 101 -3142 0 feedthrough
rlabel pdiffusion 108 -3142 108 -3142 0 feedthrough
rlabel pdiffusion 115 -3142 115 -3142 0 feedthrough
rlabel pdiffusion 122 -3142 122 -3142 0 feedthrough
rlabel pdiffusion 129 -3142 129 -3142 0 feedthrough
rlabel pdiffusion 136 -3142 136 -3142 0 feedthrough
rlabel pdiffusion 143 -3142 143 -3142 0 feedthrough
rlabel pdiffusion 150 -3142 150 -3142 0 feedthrough
rlabel pdiffusion 157 -3142 157 -3142 0 cellNo=957
rlabel pdiffusion 164 -3142 164 -3142 0 feedthrough
rlabel pdiffusion 171 -3142 171 -3142 0 feedthrough
rlabel pdiffusion 178 -3142 178 -3142 0 feedthrough
rlabel pdiffusion 185 -3142 185 -3142 0 feedthrough
rlabel pdiffusion 192 -3142 192 -3142 0 feedthrough
rlabel pdiffusion 199 -3142 199 -3142 0 feedthrough
rlabel pdiffusion 206 -3142 206 -3142 0 feedthrough
rlabel pdiffusion 213 -3142 213 -3142 0 feedthrough
rlabel pdiffusion 220 -3142 220 -3142 0 cellNo=581
rlabel pdiffusion 227 -3142 227 -3142 0 cellNo=627
rlabel pdiffusion 234 -3142 234 -3142 0 feedthrough
rlabel pdiffusion 241 -3142 241 -3142 0 feedthrough
rlabel pdiffusion 248 -3142 248 -3142 0 cellNo=23
rlabel pdiffusion 255 -3142 255 -3142 0 cellNo=246
rlabel pdiffusion 262 -3142 262 -3142 0 feedthrough
rlabel pdiffusion 269 -3142 269 -3142 0 feedthrough
rlabel pdiffusion 276 -3142 276 -3142 0 feedthrough
rlabel pdiffusion 283 -3142 283 -3142 0 feedthrough
rlabel pdiffusion 290 -3142 290 -3142 0 feedthrough
rlabel pdiffusion 297 -3142 297 -3142 0 feedthrough
rlabel pdiffusion 304 -3142 304 -3142 0 feedthrough
rlabel pdiffusion 311 -3142 311 -3142 0 feedthrough
rlabel pdiffusion 318 -3142 318 -3142 0 feedthrough
rlabel pdiffusion 325 -3142 325 -3142 0 cellNo=715
rlabel pdiffusion 332 -3142 332 -3142 0 feedthrough
rlabel pdiffusion 339 -3142 339 -3142 0 feedthrough
rlabel pdiffusion 346 -3142 346 -3142 0 feedthrough
rlabel pdiffusion 353 -3142 353 -3142 0 feedthrough
rlabel pdiffusion 360 -3142 360 -3142 0 feedthrough
rlabel pdiffusion 367 -3142 367 -3142 0 feedthrough
rlabel pdiffusion 374 -3142 374 -3142 0 feedthrough
rlabel pdiffusion 381 -3142 381 -3142 0 feedthrough
rlabel pdiffusion 388 -3142 388 -3142 0 cellNo=823
rlabel pdiffusion 395 -3142 395 -3142 0 feedthrough
rlabel pdiffusion 402 -3142 402 -3142 0 feedthrough
rlabel pdiffusion 409 -3142 409 -3142 0 cellNo=204
rlabel pdiffusion 416 -3142 416 -3142 0 feedthrough
rlabel pdiffusion 423 -3142 423 -3142 0 feedthrough
rlabel pdiffusion 430 -3142 430 -3142 0 feedthrough
rlabel pdiffusion 437 -3142 437 -3142 0 feedthrough
rlabel pdiffusion 444 -3142 444 -3142 0 feedthrough
rlabel pdiffusion 451 -3142 451 -3142 0 feedthrough
rlabel pdiffusion 458 -3142 458 -3142 0 feedthrough
rlabel pdiffusion 465 -3142 465 -3142 0 feedthrough
rlabel pdiffusion 472 -3142 472 -3142 0 feedthrough
rlabel pdiffusion 479 -3142 479 -3142 0 feedthrough
rlabel pdiffusion 486 -3142 486 -3142 0 feedthrough
rlabel pdiffusion 493 -3142 493 -3142 0 feedthrough
rlabel pdiffusion 500 -3142 500 -3142 0 feedthrough
rlabel pdiffusion 507 -3142 507 -3142 0 feedthrough
rlabel pdiffusion 514 -3142 514 -3142 0 cellNo=408
rlabel pdiffusion 521 -3142 521 -3142 0 feedthrough
rlabel pdiffusion 528 -3142 528 -3142 0 feedthrough
rlabel pdiffusion 535 -3142 535 -3142 0 feedthrough
rlabel pdiffusion 542 -3142 542 -3142 0 feedthrough
rlabel pdiffusion 549 -3142 549 -3142 0 feedthrough
rlabel pdiffusion 556 -3142 556 -3142 0 feedthrough
rlabel pdiffusion 563 -3142 563 -3142 0 feedthrough
rlabel pdiffusion 570 -3142 570 -3142 0 feedthrough
rlabel pdiffusion 577 -3142 577 -3142 0 feedthrough
rlabel pdiffusion 584 -3142 584 -3142 0 feedthrough
rlabel pdiffusion 591 -3142 591 -3142 0 cellNo=787
rlabel pdiffusion 598 -3142 598 -3142 0 feedthrough
rlabel pdiffusion 605 -3142 605 -3142 0 cellNo=776
rlabel pdiffusion 612 -3142 612 -3142 0 feedthrough
rlabel pdiffusion 619 -3142 619 -3142 0 feedthrough
rlabel pdiffusion 626 -3142 626 -3142 0 feedthrough
rlabel pdiffusion 633 -3142 633 -3142 0 feedthrough
rlabel pdiffusion 640 -3142 640 -3142 0 feedthrough
rlabel pdiffusion 647 -3142 647 -3142 0 cellNo=868
rlabel pdiffusion 654 -3142 654 -3142 0 feedthrough
rlabel pdiffusion 661 -3142 661 -3142 0 feedthrough
rlabel pdiffusion 668 -3142 668 -3142 0 feedthrough
rlabel pdiffusion 675 -3142 675 -3142 0 feedthrough
rlabel pdiffusion 682 -3142 682 -3142 0 feedthrough
rlabel pdiffusion 689 -3142 689 -3142 0 feedthrough
rlabel pdiffusion 696 -3142 696 -3142 0 cellNo=270
rlabel pdiffusion 703 -3142 703 -3142 0 feedthrough
rlabel pdiffusion 710 -3142 710 -3142 0 feedthrough
rlabel pdiffusion 717 -3142 717 -3142 0 feedthrough
rlabel pdiffusion 724 -3142 724 -3142 0 feedthrough
rlabel pdiffusion 731 -3142 731 -3142 0 feedthrough
rlabel pdiffusion 738 -3142 738 -3142 0 cellNo=213
rlabel pdiffusion 745 -3142 745 -3142 0 cellNo=796
rlabel pdiffusion 752 -3142 752 -3142 0 feedthrough
rlabel pdiffusion 759 -3142 759 -3142 0 cellNo=228
rlabel pdiffusion 766 -3142 766 -3142 0 feedthrough
rlabel pdiffusion 773 -3142 773 -3142 0 feedthrough
rlabel pdiffusion 780 -3142 780 -3142 0 feedthrough
rlabel pdiffusion 787 -3142 787 -3142 0 feedthrough
rlabel pdiffusion 794 -3142 794 -3142 0 cellNo=221
rlabel pdiffusion 801 -3142 801 -3142 0 feedthrough
rlabel pdiffusion 808 -3142 808 -3142 0 cellNo=74
rlabel pdiffusion 815 -3142 815 -3142 0 feedthrough
rlabel pdiffusion 822 -3142 822 -3142 0 feedthrough
rlabel pdiffusion 829 -3142 829 -3142 0 feedthrough
rlabel pdiffusion 836 -3142 836 -3142 0 feedthrough
rlabel pdiffusion 843 -3142 843 -3142 0 feedthrough
rlabel pdiffusion 850 -3142 850 -3142 0 feedthrough
rlabel pdiffusion 857 -3142 857 -3142 0 feedthrough
rlabel pdiffusion 864 -3142 864 -3142 0 feedthrough
rlabel pdiffusion 871 -3142 871 -3142 0 feedthrough
rlabel pdiffusion 878 -3142 878 -3142 0 feedthrough
rlabel pdiffusion 885 -3142 885 -3142 0 feedthrough
rlabel pdiffusion 892 -3142 892 -3142 0 feedthrough
rlabel pdiffusion 899 -3142 899 -3142 0 cellNo=570
rlabel pdiffusion 906 -3142 906 -3142 0 feedthrough
rlabel pdiffusion 913 -3142 913 -3142 0 cellNo=495
rlabel pdiffusion 920 -3142 920 -3142 0 feedthrough
rlabel pdiffusion 927 -3142 927 -3142 0 feedthrough
rlabel pdiffusion 934 -3142 934 -3142 0 feedthrough
rlabel pdiffusion 941 -3142 941 -3142 0 feedthrough
rlabel pdiffusion 948 -3142 948 -3142 0 feedthrough
rlabel pdiffusion 955 -3142 955 -3142 0 feedthrough
rlabel pdiffusion 962 -3142 962 -3142 0 feedthrough
rlabel pdiffusion 969 -3142 969 -3142 0 feedthrough
rlabel pdiffusion 976 -3142 976 -3142 0 feedthrough
rlabel pdiffusion 983 -3142 983 -3142 0 feedthrough
rlabel pdiffusion 990 -3142 990 -3142 0 feedthrough
rlabel pdiffusion 997 -3142 997 -3142 0 feedthrough
rlabel pdiffusion 1004 -3142 1004 -3142 0 feedthrough
rlabel pdiffusion 1011 -3142 1011 -3142 0 cellNo=73
rlabel pdiffusion 1018 -3142 1018 -3142 0 feedthrough
rlabel pdiffusion 1025 -3142 1025 -3142 0 feedthrough
rlabel pdiffusion 1032 -3142 1032 -3142 0 feedthrough
rlabel pdiffusion 1039 -3142 1039 -3142 0 feedthrough
rlabel pdiffusion 1046 -3142 1046 -3142 0 feedthrough
rlabel pdiffusion 1053 -3142 1053 -3142 0 feedthrough
rlabel pdiffusion 1060 -3142 1060 -3142 0 feedthrough
rlabel pdiffusion 1067 -3142 1067 -3142 0 feedthrough
rlabel pdiffusion 1074 -3142 1074 -3142 0 feedthrough
rlabel pdiffusion 1081 -3142 1081 -3142 0 feedthrough
rlabel pdiffusion 1088 -3142 1088 -3142 0 feedthrough
rlabel pdiffusion 1095 -3142 1095 -3142 0 feedthrough
rlabel pdiffusion 1102 -3142 1102 -3142 0 feedthrough
rlabel pdiffusion 1109 -3142 1109 -3142 0 feedthrough
rlabel pdiffusion 1116 -3142 1116 -3142 0 feedthrough
rlabel pdiffusion 1123 -3142 1123 -3142 0 feedthrough
rlabel pdiffusion 1130 -3142 1130 -3142 0 feedthrough
rlabel pdiffusion 1137 -3142 1137 -3142 0 feedthrough
rlabel pdiffusion 1144 -3142 1144 -3142 0 feedthrough
rlabel pdiffusion 1151 -3142 1151 -3142 0 feedthrough
rlabel pdiffusion 1158 -3142 1158 -3142 0 feedthrough
rlabel pdiffusion 1165 -3142 1165 -3142 0 feedthrough
rlabel pdiffusion 1172 -3142 1172 -3142 0 feedthrough
rlabel pdiffusion 1179 -3142 1179 -3142 0 feedthrough
rlabel pdiffusion 1186 -3142 1186 -3142 0 feedthrough
rlabel pdiffusion 1193 -3142 1193 -3142 0 feedthrough
rlabel pdiffusion 1200 -3142 1200 -3142 0 cellNo=530
rlabel pdiffusion 1207 -3142 1207 -3142 0 cellNo=519
rlabel pdiffusion 1214 -3142 1214 -3142 0 feedthrough
rlabel pdiffusion 1221 -3142 1221 -3142 0 feedthrough
rlabel pdiffusion 1228 -3142 1228 -3142 0 feedthrough
rlabel pdiffusion 1235 -3142 1235 -3142 0 feedthrough
rlabel pdiffusion 1242 -3142 1242 -3142 0 feedthrough
rlabel pdiffusion 1249 -3142 1249 -3142 0 feedthrough
rlabel pdiffusion 1256 -3142 1256 -3142 0 feedthrough
rlabel pdiffusion 1263 -3142 1263 -3142 0 feedthrough
rlabel pdiffusion 1270 -3142 1270 -3142 0 feedthrough
rlabel pdiffusion 1277 -3142 1277 -3142 0 feedthrough
rlabel pdiffusion 1284 -3142 1284 -3142 0 feedthrough
rlabel pdiffusion 1291 -3142 1291 -3142 0 feedthrough
rlabel pdiffusion 1298 -3142 1298 -3142 0 feedthrough
rlabel pdiffusion 1305 -3142 1305 -3142 0 feedthrough
rlabel pdiffusion 1312 -3142 1312 -3142 0 feedthrough
rlabel pdiffusion 1319 -3142 1319 -3142 0 feedthrough
rlabel pdiffusion 1326 -3142 1326 -3142 0 feedthrough
rlabel pdiffusion 1333 -3142 1333 -3142 0 cellNo=680
rlabel pdiffusion 1340 -3142 1340 -3142 0 feedthrough
rlabel pdiffusion 1354 -3142 1354 -3142 0 feedthrough
rlabel pdiffusion 1361 -3142 1361 -3142 0 feedthrough
rlabel pdiffusion 1368 -3142 1368 -3142 0 feedthrough
rlabel pdiffusion 1375 -3142 1375 -3142 0 feedthrough
rlabel pdiffusion 3 -3235 3 -3235 0 cellNo=1083
rlabel pdiffusion 10 -3235 10 -3235 0 cellNo=1136
rlabel pdiffusion 17 -3235 17 -3235 0 cellNo=1137
rlabel pdiffusion 24 -3235 24 -3235 0 cellNo=1138
rlabel pdiffusion 31 -3235 31 -3235 0 cellNo=1139
rlabel pdiffusion 38 -3235 38 -3235 0 cellNo=1140
rlabel pdiffusion 45 -3235 45 -3235 0 cellNo=1141
rlabel pdiffusion 52 -3235 52 -3235 0 cellNo=1142
rlabel pdiffusion 59 -3235 59 -3235 0 cellNo=1143
rlabel pdiffusion 66 -3235 66 -3235 0 cellNo=1135
rlabel pdiffusion 73 -3235 73 -3235 0 cellNo=1160
rlabel pdiffusion 80 -3235 80 -3235 0 cellNo=1146
rlabel pdiffusion 87 -3235 87 -3235 0 cellNo=1147
rlabel pdiffusion 94 -3235 94 -3235 0 cellNo=1152
rlabel pdiffusion 164 -3235 164 -3235 0 feedthrough
rlabel pdiffusion 171 -3235 171 -3235 0 feedthrough
rlabel pdiffusion 178 -3235 178 -3235 0 feedthrough
rlabel pdiffusion 185 -3235 185 -3235 0 cellNo=999
rlabel pdiffusion 192 -3235 192 -3235 0 feedthrough
rlabel pdiffusion 199 -3235 199 -3235 0 feedthrough
rlabel pdiffusion 206 -3235 206 -3235 0 feedthrough
rlabel pdiffusion 213 -3235 213 -3235 0 feedthrough
rlabel pdiffusion 220 -3235 220 -3235 0 feedthrough
rlabel pdiffusion 227 -3235 227 -3235 0 feedthrough
rlabel pdiffusion 234 -3235 234 -3235 0 feedthrough
rlabel pdiffusion 241 -3235 241 -3235 0 feedthrough
rlabel pdiffusion 248 -3235 248 -3235 0 feedthrough
rlabel pdiffusion 255 -3235 255 -3235 0 feedthrough
rlabel pdiffusion 262 -3235 262 -3235 0 feedthrough
rlabel pdiffusion 269 -3235 269 -3235 0 feedthrough
rlabel pdiffusion 276 -3235 276 -3235 0 feedthrough
rlabel pdiffusion 283 -3235 283 -3235 0 cellNo=695
rlabel pdiffusion 290 -3235 290 -3235 0 feedthrough
rlabel pdiffusion 297 -3235 297 -3235 0 feedthrough
rlabel pdiffusion 304 -3235 304 -3235 0 feedthrough
rlabel pdiffusion 311 -3235 311 -3235 0 feedthrough
rlabel pdiffusion 318 -3235 318 -3235 0 feedthrough
rlabel pdiffusion 325 -3235 325 -3235 0 feedthrough
rlabel pdiffusion 332 -3235 332 -3235 0 feedthrough
rlabel pdiffusion 339 -3235 339 -3235 0 feedthrough
rlabel pdiffusion 346 -3235 346 -3235 0 feedthrough
rlabel pdiffusion 353 -3235 353 -3235 0 feedthrough
rlabel pdiffusion 360 -3235 360 -3235 0 feedthrough
rlabel pdiffusion 367 -3235 367 -3235 0 feedthrough
rlabel pdiffusion 374 -3235 374 -3235 0 feedthrough
rlabel pdiffusion 381 -3235 381 -3235 0 feedthrough
rlabel pdiffusion 388 -3235 388 -3235 0 feedthrough
rlabel pdiffusion 395 -3235 395 -3235 0 feedthrough
rlabel pdiffusion 402 -3235 402 -3235 0 feedthrough
rlabel pdiffusion 409 -3235 409 -3235 0 feedthrough
rlabel pdiffusion 416 -3235 416 -3235 0 feedthrough
rlabel pdiffusion 423 -3235 423 -3235 0 feedthrough
rlabel pdiffusion 430 -3235 430 -3235 0 feedthrough
rlabel pdiffusion 437 -3235 437 -3235 0 feedthrough
rlabel pdiffusion 444 -3235 444 -3235 0 feedthrough
rlabel pdiffusion 451 -3235 451 -3235 0 feedthrough
rlabel pdiffusion 458 -3235 458 -3235 0 cellNo=398
rlabel pdiffusion 465 -3235 465 -3235 0 feedthrough
rlabel pdiffusion 472 -3235 472 -3235 0 feedthrough
rlabel pdiffusion 479 -3235 479 -3235 0 cellNo=584
rlabel pdiffusion 486 -3235 486 -3235 0 feedthrough
rlabel pdiffusion 493 -3235 493 -3235 0 feedthrough
rlabel pdiffusion 500 -3235 500 -3235 0 feedthrough
rlabel pdiffusion 507 -3235 507 -3235 0 feedthrough
rlabel pdiffusion 514 -3235 514 -3235 0 feedthrough
rlabel pdiffusion 521 -3235 521 -3235 0 feedthrough
rlabel pdiffusion 528 -3235 528 -3235 0 feedthrough
rlabel pdiffusion 535 -3235 535 -3235 0 feedthrough
rlabel pdiffusion 542 -3235 542 -3235 0 cellNo=671
rlabel pdiffusion 549 -3235 549 -3235 0 feedthrough
rlabel pdiffusion 556 -3235 556 -3235 0 feedthrough
rlabel pdiffusion 563 -3235 563 -3235 0 feedthrough
rlabel pdiffusion 570 -3235 570 -3235 0 feedthrough
rlabel pdiffusion 577 -3235 577 -3235 0 cellNo=859
rlabel pdiffusion 584 -3235 584 -3235 0 feedthrough
rlabel pdiffusion 591 -3235 591 -3235 0 feedthrough
rlabel pdiffusion 598 -3235 598 -3235 0 feedthrough
rlabel pdiffusion 605 -3235 605 -3235 0 feedthrough
rlabel pdiffusion 612 -3235 612 -3235 0 feedthrough
rlabel pdiffusion 619 -3235 619 -3235 0 feedthrough
rlabel pdiffusion 626 -3235 626 -3235 0 feedthrough
rlabel pdiffusion 633 -3235 633 -3235 0 cellNo=76
rlabel pdiffusion 640 -3235 640 -3235 0 feedthrough
rlabel pdiffusion 647 -3235 647 -3235 0 feedthrough
rlabel pdiffusion 654 -3235 654 -3235 0 feedthrough
rlabel pdiffusion 661 -3235 661 -3235 0 feedthrough
rlabel pdiffusion 668 -3235 668 -3235 0 feedthrough
rlabel pdiffusion 675 -3235 675 -3235 0 feedthrough
rlabel pdiffusion 682 -3235 682 -3235 0 feedthrough
rlabel pdiffusion 689 -3235 689 -3235 0 feedthrough
rlabel pdiffusion 696 -3235 696 -3235 0 feedthrough
rlabel pdiffusion 703 -3235 703 -3235 0 feedthrough
rlabel pdiffusion 710 -3235 710 -3235 0 cellNo=862
rlabel pdiffusion 717 -3235 717 -3235 0 feedthrough
rlabel pdiffusion 724 -3235 724 -3235 0 feedthrough
rlabel pdiffusion 731 -3235 731 -3235 0 feedthrough
rlabel pdiffusion 738 -3235 738 -3235 0 feedthrough
rlabel pdiffusion 745 -3235 745 -3235 0 cellNo=460
rlabel pdiffusion 752 -3235 752 -3235 0 cellNo=986
rlabel pdiffusion 759 -3235 759 -3235 0 feedthrough
rlabel pdiffusion 766 -3235 766 -3235 0 cellNo=606
rlabel pdiffusion 773 -3235 773 -3235 0 feedthrough
rlabel pdiffusion 780 -3235 780 -3235 0 feedthrough
rlabel pdiffusion 787 -3235 787 -3235 0 feedthrough
rlabel pdiffusion 794 -3235 794 -3235 0 feedthrough
rlabel pdiffusion 801 -3235 801 -3235 0 feedthrough
rlabel pdiffusion 808 -3235 808 -3235 0 cellNo=390
rlabel pdiffusion 815 -3235 815 -3235 0 feedthrough
rlabel pdiffusion 822 -3235 822 -3235 0 feedthrough
rlabel pdiffusion 829 -3235 829 -3235 0 feedthrough
rlabel pdiffusion 836 -3235 836 -3235 0 feedthrough
rlabel pdiffusion 843 -3235 843 -3235 0 feedthrough
rlabel pdiffusion 850 -3235 850 -3235 0 feedthrough
rlabel pdiffusion 857 -3235 857 -3235 0 feedthrough
rlabel pdiffusion 864 -3235 864 -3235 0 feedthrough
rlabel pdiffusion 871 -3235 871 -3235 0 feedthrough
rlabel pdiffusion 878 -3235 878 -3235 0 feedthrough
rlabel pdiffusion 885 -3235 885 -3235 0 feedthrough
rlabel pdiffusion 892 -3235 892 -3235 0 cellNo=950
rlabel pdiffusion 899 -3235 899 -3235 0 feedthrough
rlabel pdiffusion 906 -3235 906 -3235 0 feedthrough
rlabel pdiffusion 913 -3235 913 -3235 0 feedthrough
rlabel pdiffusion 920 -3235 920 -3235 0 feedthrough
rlabel pdiffusion 927 -3235 927 -3235 0 feedthrough
rlabel pdiffusion 934 -3235 934 -3235 0 feedthrough
rlabel pdiffusion 941 -3235 941 -3235 0 cellNo=596
rlabel pdiffusion 948 -3235 948 -3235 0 feedthrough
rlabel pdiffusion 955 -3235 955 -3235 0 feedthrough
rlabel pdiffusion 962 -3235 962 -3235 0 cellNo=305
rlabel pdiffusion 969 -3235 969 -3235 0 feedthrough
rlabel pdiffusion 976 -3235 976 -3235 0 feedthrough
rlabel pdiffusion 983 -3235 983 -3235 0 feedthrough
rlabel pdiffusion 990 -3235 990 -3235 0 feedthrough
rlabel pdiffusion 997 -3235 997 -3235 0 feedthrough
rlabel pdiffusion 1004 -3235 1004 -3235 0 feedthrough
rlabel pdiffusion 1011 -3235 1011 -3235 0 feedthrough
rlabel pdiffusion 1018 -3235 1018 -3235 0 feedthrough
rlabel pdiffusion 1025 -3235 1025 -3235 0 feedthrough
rlabel pdiffusion 1032 -3235 1032 -3235 0 feedthrough
rlabel pdiffusion 1039 -3235 1039 -3235 0 feedthrough
rlabel pdiffusion 1046 -3235 1046 -3235 0 feedthrough
rlabel pdiffusion 1053 -3235 1053 -3235 0 feedthrough
rlabel pdiffusion 1060 -3235 1060 -3235 0 feedthrough
rlabel pdiffusion 1067 -3235 1067 -3235 0 feedthrough
rlabel pdiffusion 1074 -3235 1074 -3235 0 feedthrough
rlabel pdiffusion 1081 -3235 1081 -3235 0 feedthrough
rlabel pdiffusion 1088 -3235 1088 -3235 0 feedthrough
rlabel pdiffusion 1095 -3235 1095 -3235 0 feedthrough
rlabel pdiffusion 1102 -3235 1102 -3235 0 feedthrough
rlabel pdiffusion 1109 -3235 1109 -3235 0 feedthrough
rlabel pdiffusion 1116 -3235 1116 -3235 0 feedthrough
rlabel pdiffusion 1123 -3235 1123 -3235 0 feedthrough
rlabel pdiffusion 1130 -3235 1130 -3235 0 feedthrough
rlabel pdiffusion 1137 -3235 1137 -3235 0 feedthrough
rlabel pdiffusion 1144 -3235 1144 -3235 0 feedthrough
rlabel pdiffusion 1151 -3235 1151 -3235 0 feedthrough
rlabel pdiffusion 1158 -3235 1158 -3235 0 feedthrough
rlabel pdiffusion 1165 -3235 1165 -3235 0 cellNo=981
rlabel pdiffusion 1172 -3235 1172 -3235 0 feedthrough
rlabel pdiffusion 1179 -3235 1179 -3235 0 feedthrough
rlabel pdiffusion 1186 -3235 1186 -3235 0 feedthrough
rlabel pdiffusion 1193 -3235 1193 -3235 0 feedthrough
rlabel pdiffusion 1200 -3235 1200 -3235 0 cellNo=730
rlabel pdiffusion 1207 -3235 1207 -3235 0 feedthrough
rlabel pdiffusion 1214 -3235 1214 -3235 0 feedthrough
rlabel pdiffusion 1221 -3235 1221 -3235 0 feedthrough
rlabel pdiffusion 1228 -3235 1228 -3235 0 cellNo=231
rlabel pdiffusion 1235 -3235 1235 -3235 0 feedthrough
rlabel pdiffusion 1242 -3235 1242 -3235 0 feedthrough
rlabel pdiffusion 1249 -3235 1249 -3235 0 feedthrough
rlabel pdiffusion 1256 -3235 1256 -3235 0 cellNo=26
rlabel pdiffusion 1263 -3235 1263 -3235 0 feedthrough
rlabel pdiffusion 1270 -3235 1270 -3235 0 feedthrough
rlabel pdiffusion 1277 -3235 1277 -3235 0 feedthrough
rlabel pdiffusion 1284 -3235 1284 -3235 0 cellNo=569
rlabel pdiffusion 1291 -3235 1291 -3235 0 cellNo=399
rlabel pdiffusion 1298 -3235 1298 -3235 0 feedthrough
rlabel pdiffusion 1305 -3235 1305 -3235 0 feedthrough
rlabel pdiffusion 1347 -3235 1347 -3235 0 feedthrough
rlabel pdiffusion 1354 -3235 1354 -3235 0 feedthrough
rlabel pdiffusion 1361 -3235 1361 -3235 0 feedthrough
rlabel pdiffusion 3 -3312 3 -3312 0 cellNo=1177
rlabel pdiffusion 10 -3312 10 -3312 0 cellNo=1178
rlabel pdiffusion 17 -3312 17 -3312 0 cellNo=1179
rlabel pdiffusion 24 -3312 24 -3312 0 cellNo=1180
rlabel pdiffusion 31 -3312 31 -3312 0 cellNo=1181
rlabel pdiffusion 38 -3312 38 -3312 0 cellNo=1182
rlabel pdiffusion 45 -3312 45 -3312 0 cellNo=1183
rlabel pdiffusion 52 -3312 52 -3312 0 cellNo=1184
rlabel pdiffusion 59 -3312 59 -3312 0 cellNo=1185
rlabel pdiffusion 66 -3312 66 -3312 0 cellNo=1186
rlabel pdiffusion 73 -3312 73 -3312 0 cellNo=1187
rlabel pdiffusion 80 -3312 80 -3312 0 cellNo=1284
rlabel pdiffusion 87 -3312 87 -3312 0 cellNo=1232
rlabel pdiffusion 94 -3312 94 -3312 0 cellNo=1190
rlabel pdiffusion 157 -3312 157 -3312 0 feedthrough
rlabel pdiffusion 164 -3312 164 -3312 0 feedthrough
rlabel pdiffusion 171 -3312 171 -3312 0 feedthrough
rlabel pdiffusion 178 -3312 178 -3312 0 feedthrough
rlabel pdiffusion 185 -3312 185 -3312 0 feedthrough
rlabel pdiffusion 192 -3312 192 -3312 0 feedthrough
rlabel pdiffusion 199 -3312 199 -3312 0 cellNo=415
rlabel pdiffusion 206 -3312 206 -3312 0 feedthrough
rlabel pdiffusion 213 -3312 213 -3312 0 feedthrough
rlabel pdiffusion 220 -3312 220 -3312 0 feedthrough
rlabel pdiffusion 227 -3312 227 -3312 0 feedthrough
rlabel pdiffusion 234 -3312 234 -3312 0 feedthrough
rlabel pdiffusion 241 -3312 241 -3312 0 cellNo=223
rlabel pdiffusion 248 -3312 248 -3312 0 feedthrough
rlabel pdiffusion 255 -3312 255 -3312 0 feedthrough
rlabel pdiffusion 262 -3312 262 -3312 0 feedthrough
rlabel pdiffusion 269 -3312 269 -3312 0 feedthrough
rlabel pdiffusion 276 -3312 276 -3312 0 feedthrough
rlabel pdiffusion 283 -3312 283 -3312 0 feedthrough
rlabel pdiffusion 290 -3312 290 -3312 0 feedthrough
rlabel pdiffusion 297 -3312 297 -3312 0 feedthrough
rlabel pdiffusion 304 -3312 304 -3312 0 feedthrough
rlabel pdiffusion 311 -3312 311 -3312 0 feedthrough
rlabel pdiffusion 318 -3312 318 -3312 0 feedthrough
rlabel pdiffusion 325 -3312 325 -3312 0 feedthrough
rlabel pdiffusion 332 -3312 332 -3312 0 feedthrough
rlabel pdiffusion 339 -3312 339 -3312 0 feedthrough
rlabel pdiffusion 346 -3312 346 -3312 0 feedthrough
rlabel pdiffusion 353 -3312 353 -3312 0 feedthrough
rlabel pdiffusion 360 -3312 360 -3312 0 feedthrough
rlabel pdiffusion 367 -3312 367 -3312 0 feedthrough
rlabel pdiffusion 374 -3312 374 -3312 0 feedthrough
rlabel pdiffusion 381 -3312 381 -3312 0 feedthrough
rlabel pdiffusion 388 -3312 388 -3312 0 feedthrough
rlabel pdiffusion 395 -3312 395 -3312 0 cellNo=856
rlabel pdiffusion 402 -3312 402 -3312 0 feedthrough
rlabel pdiffusion 409 -3312 409 -3312 0 feedthrough
rlabel pdiffusion 416 -3312 416 -3312 0 feedthrough
rlabel pdiffusion 423 -3312 423 -3312 0 feedthrough
rlabel pdiffusion 430 -3312 430 -3312 0 feedthrough
rlabel pdiffusion 437 -3312 437 -3312 0 feedthrough
rlabel pdiffusion 444 -3312 444 -3312 0 feedthrough
rlabel pdiffusion 451 -3312 451 -3312 0 feedthrough
rlabel pdiffusion 458 -3312 458 -3312 0 feedthrough
rlabel pdiffusion 465 -3312 465 -3312 0 feedthrough
rlabel pdiffusion 472 -3312 472 -3312 0 feedthrough
rlabel pdiffusion 479 -3312 479 -3312 0 feedthrough
rlabel pdiffusion 486 -3312 486 -3312 0 cellNo=914
rlabel pdiffusion 493 -3312 493 -3312 0 feedthrough
rlabel pdiffusion 500 -3312 500 -3312 0 feedthrough
rlabel pdiffusion 507 -3312 507 -3312 0 feedthrough
rlabel pdiffusion 514 -3312 514 -3312 0 feedthrough
rlabel pdiffusion 521 -3312 521 -3312 0 feedthrough
rlabel pdiffusion 528 -3312 528 -3312 0 feedthrough
rlabel pdiffusion 535 -3312 535 -3312 0 cellNo=372
rlabel pdiffusion 542 -3312 542 -3312 0 feedthrough
rlabel pdiffusion 549 -3312 549 -3312 0 feedthrough
rlabel pdiffusion 556 -3312 556 -3312 0 feedthrough
rlabel pdiffusion 563 -3312 563 -3312 0 feedthrough
rlabel pdiffusion 570 -3312 570 -3312 0 feedthrough
rlabel pdiffusion 577 -3312 577 -3312 0 feedthrough
rlabel pdiffusion 584 -3312 584 -3312 0 feedthrough
rlabel pdiffusion 591 -3312 591 -3312 0 feedthrough
rlabel pdiffusion 598 -3312 598 -3312 0 feedthrough
rlabel pdiffusion 605 -3312 605 -3312 0 feedthrough
rlabel pdiffusion 612 -3312 612 -3312 0 cellNo=625
rlabel pdiffusion 619 -3312 619 -3312 0 feedthrough
rlabel pdiffusion 626 -3312 626 -3312 0 feedthrough
rlabel pdiffusion 633 -3312 633 -3312 0 feedthrough
rlabel pdiffusion 640 -3312 640 -3312 0 feedthrough
rlabel pdiffusion 647 -3312 647 -3312 0 feedthrough
rlabel pdiffusion 654 -3312 654 -3312 0 cellNo=729
rlabel pdiffusion 661 -3312 661 -3312 0 cellNo=202
rlabel pdiffusion 668 -3312 668 -3312 0 cellNo=154
rlabel pdiffusion 675 -3312 675 -3312 0 feedthrough
rlabel pdiffusion 682 -3312 682 -3312 0 feedthrough
rlabel pdiffusion 689 -3312 689 -3312 0 cellNo=397
rlabel pdiffusion 696 -3312 696 -3312 0 feedthrough
rlabel pdiffusion 703 -3312 703 -3312 0 feedthrough
rlabel pdiffusion 710 -3312 710 -3312 0 feedthrough
rlabel pdiffusion 717 -3312 717 -3312 0 feedthrough
rlabel pdiffusion 724 -3312 724 -3312 0 feedthrough
rlabel pdiffusion 731 -3312 731 -3312 0 cellNo=478
rlabel pdiffusion 738 -3312 738 -3312 0 feedthrough
rlabel pdiffusion 745 -3312 745 -3312 0 feedthrough
rlabel pdiffusion 752 -3312 752 -3312 0 feedthrough
rlabel pdiffusion 759 -3312 759 -3312 0 cellNo=882
rlabel pdiffusion 766 -3312 766 -3312 0 feedthrough
rlabel pdiffusion 773 -3312 773 -3312 0 feedthrough
rlabel pdiffusion 780 -3312 780 -3312 0 feedthrough
rlabel pdiffusion 787 -3312 787 -3312 0 feedthrough
rlabel pdiffusion 794 -3312 794 -3312 0 feedthrough
rlabel pdiffusion 801 -3312 801 -3312 0 feedthrough
rlabel pdiffusion 808 -3312 808 -3312 0 feedthrough
rlabel pdiffusion 815 -3312 815 -3312 0 feedthrough
rlabel pdiffusion 822 -3312 822 -3312 0 cellNo=392
rlabel pdiffusion 829 -3312 829 -3312 0 feedthrough
rlabel pdiffusion 836 -3312 836 -3312 0 cellNo=210
rlabel pdiffusion 843 -3312 843 -3312 0 feedthrough
rlabel pdiffusion 850 -3312 850 -3312 0 feedthrough
rlabel pdiffusion 857 -3312 857 -3312 0 cellNo=781
rlabel pdiffusion 864 -3312 864 -3312 0 feedthrough
rlabel pdiffusion 871 -3312 871 -3312 0 cellNo=966
rlabel pdiffusion 878 -3312 878 -3312 0 feedthrough
rlabel pdiffusion 885 -3312 885 -3312 0 feedthrough
rlabel pdiffusion 892 -3312 892 -3312 0 cellNo=946
rlabel pdiffusion 899 -3312 899 -3312 0 feedthrough
rlabel pdiffusion 906 -3312 906 -3312 0 feedthrough
rlabel pdiffusion 913 -3312 913 -3312 0 feedthrough
rlabel pdiffusion 920 -3312 920 -3312 0 feedthrough
rlabel pdiffusion 927 -3312 927 -3312 0 feedthrough
rlabel pdiffusion 934 -3312 934 -3312 0 feedthrough
rlabel pdiffusion 941 -3312 941 -3312 0 feedthrough
rlabel pdiffusion 948 -3312 948 -3312 0 feedthrough
rlabel pdiffusion 955 -3312 955 -3312 0 feedthrough
rlabel pdiffusion 962 -3312 962 -3312 0 feedthrough
rlabel pdiffusion 969 -3312 969 -3312 0 feedthrough
rlabel pdiffusion 976 -3312 976 -3312 0 feedthrough
rlabel pdiffusion 983 -3312 983 -3312 0 feedthrough
rlabel pdiffusion 990 -3312 990 -3312 0 feedthrough
rlabel pdiffusion 997 -3312 997 -3312 0 feedthrough
rlabel pdiffusion 1004 -3312 1004 -3312 0 cellNo=260
rlabel pdiffusion 1011 -3312 1011 -3312 0 feedthrough
rlabel pdiffusion 1018 -3312 1018 -3312 0 feedthrough
rlabel pdiffusion 1025 -3312 1025 -3312 0 cellNo=691
rlabel pdiffusion 1032 -3312 1032 -3312 0 feedthrough
rlabel pdiffusion 1039 -3312 1039 -3312 0 feedthrough
rlabel pdiffusion 1046 -3312 1046 -3312 0 feedthrough
rlabel pdiffusion 1053 -3312 1053 -3312 0 feedthrough
rlabel pdiffusion 1060 -3312 1060 -3312 0 feedthrough
rlabel pdiffusion 1067 -3312 1067 -3312 0 feedthrough
rlabel pdiffusion 1074 -3312 1074 -3312 0 feedthrough
rlabel pdiffusion 1081 -3312 1081 -3312 0 feedthrough
rlabel pdiffusion 1088 -3312 1088 -3312 0 feedthrough
rlabel pdiffusion 1095 -3312 1095 -3312 0 feedthrough
rlabel pdiffusion 1102 -3312 1102 -3312 0 feedthrough
rlabel pdiffusion 1109 -3312 1109 -3312 0 feedthrough
rlabel pdiffusion 1116 -3312 1116 -3312 0 feedthrough
rlabel pdiffusion 1123 -3312 1123 -3312 0 feedthrough
rlabel pdiffusion 1130 -3312 1130 -3312 0 feedthrough
rlabel pdiffusion 1137 -3312 1137 -3312 0 cellNo=725
rlabel pdiffusion 1144 -3312 1144 -3312 0 feedthrough
rlabel pdiffusion 1151 -3312 1151 -3312 0 feedthrough
rlabel pdiffusion 1158 -3312 1158 -3312 0 feedthrough
rlabel pdiffusion 1165 -3312 1165 -3312 0 feedthrough
rlabel pdiffusion 1172 -3312 1172 -3312 0 feedthrough
rlabel pdiffusion 1179 -3312 1179 -3312 0 feedthrough
rlabel pdiffusion 1186 -3312 1186 -3312 0 feedthrough
rlabel pdiffusion 1193 -3312 1193 -3312 0 feedthrough
rlabel pdiffusion 1200 -3312 1200 -3312 0 feedthrough
rlabel pdiffusion 1207 -3312 1207 -3312 0 feedthrough
rlabel pdiffusion 1214 -3312 1214 -3312 0 feedthrough
rlabel pdiffusion 1221 -3312 1221 -3312 0 feedthrough
rlabel pdiffusion 1228 -3312 1228 -3312 0 feedthrough
rlabel pdiffusion 1235 -3312 1235 -3312 0 feedthrough
rlabel pdiffusion 1242 -3312 1242 -3312 0 feedthrough
rlabel pdiffusion 1249 -3312 1249 -3312 0 feedthrough
rlabel pdiffusion 1256 -3312 1256 -3312 0 feedthrough
rlabel pdiffusion 1263 -3312 1263 -3312 0 feedthrough
rlabel pdiffusion 1270 -3312 1270 -3312 0 cellNo=905
rlabel pdiffusion 1277 -3312 1277 -3312 0 feedthrough
rlabel pdiffusion 1291 -3312 1291 -3312 0 feedthrough
rlabel pdiffusion 1340 -3312 1340 -3312 0 feedthrough
rlabel pdiffusion 1347 -3312 1347 -3312 0 feedthrough
rlabel pdiffusion 1354 -3312 1354 -3312 0 feedthrough
rlabel pdiffusion 3 -3385 3 -3385 0 cellNo=1216
rlabel pdiffusion 10 -3385 10 -3385 0 cellNo=1220
rlabel pdiffusion 17 -3385 17 -3385 0 cellNo=1221
rlabel pdiffusion 24 -3385 24 -3385 0 cellNo=1222
rlabel pdiffusion 31 -3385 31 -3385 0 cellNo=1223
rlabel pdiffusion 38 -3385 38 -3385 0 cellNo=1224
rlabel pdiffusion 45 -3385 45 -3385 0 cellNo=1225
rlabel pdiffusion 52 -3385 52 -3385 0 cellNo=1226
rlabel pdiffusion 59 -3385 59 -3385 0 cellNo=1227
rlabel pdiffusion 66 -3385 66 -3385 0 cellNo=1228
rlabel pdiffusion 73 -3385 73 -3385 0 cellNo=1229
rlabel pdiffusion 80 -3385 80 -3385 0 cellNo=1230
rlabel pdiffusion 87 -3385 87 -3385 0 cellNo=1231
rlabel pdiffusion 94 -3385 94 -3385 0 cellNo=1219
rlabel pdiffusion 199 -3385 199 -3385 0 feedthrough
rlabel pdiffusion 206 -3385 206 -3385 0 feedthrough
rlabel pdiffusion 213 -3385 213 -3385 0 feedthrough
rlabel pdiffusion 220 -3385 220 -3385 0 feedthrough
rlabel pdiffusion 227 -3385 227 -3385 0 feedthrough
rlabel pdiffusion 234 -3385 234 -3385 0 feedthrough
rlabel pdiffusion 241 -3385 241 -3385 0 feedthrough
rlabel pdiffusion 248 -3385 248 -3385 0 feedthrough
rlabel pdiffusion 255 -3385 255 -3385 0 feedthrough
rlabel pdiffusion 262 -3385 262 -3385 0 cellNo=3
rlabel pdiffusion 269 -3385 269 -3385 0 cellNo=977
rlabel pdiffusion 276 -3385 276 -3385 0 cellNo=795
rlabel pdiffusion 283 -3385 283 -3385 0 feedthrough
rlabel pdiffusion 290 -3385 290 -3385 0 feedthrough
rlabel pdiffusion 297 -3385 297 -3385 0 feedthrough
rlabel pdiffusion 304 -3385 304 -3385 0 feedthrough
rlabel pdiffusion 311 -3385 311 -3385 0 feedthrough
rlabel pdiffusion 318 -3385 318 -3385 0 feedthrough
rlabel pdiffusion 325 -3385 325 -3385 0 feedthrough
rlabel pdiffusion 332 -3385 332 -3385 0 feedthrough
rlabel pdiffusion 339 -3385 339 -3385 0 feedthrough
rlabel pdiffusion 346 -3385 346 -3385 0 feedthrough
rlabel pdiffusion 353 -3385 353 -3385 0 feedthrough
rlabel pdiffusion 360 -3385 360 -3385 0 feedthrough
rlabel pdiffusion 367 -3385 367 -3385 0 feedthrough
rlabel pdiffusion 374 -3385 374 -3385 0 feedthrough
rlabel pdiffusion 381 -3385 381 -3385 0 feedthrough
rlabel pdiffusion 388 -3385 388 -3385 0 feedthrough
rlabel pdiffusion 395 -3385 395 -3385 0 feedthrough
rlabel pdiffusion 402 -3385 402 -3385 0 cellNo=738
rlabel pdiffusion 409 -3385 409 -3385 0 cellNo=904
rlabel pdiffusion 416 -3385 416 -3385 0 feedthrough
rlabel pdiffusion 423 -3385 423 -3385 0 cellNo=883
rlabel pdiffusion 430 -3385 430 -3385 0 feedthrough
rlabel pdiffusion 437 -3385 437 -3385 0 feedthrough
rlabel pdiffusion 444 -3385 444 -3385 0 feedthrough
rlabel pdiffusion 451 -3385 451 -3385 0 feedthrough
rlabel pdiffusion 458 -3385 458 -3385 0 feedthrough
rlabel pdiffusion 465 -3385 465 -3385 0 feedthrough
rlabel pdiffusion 472 -3385 472 -3385 0 cellNo=750
rlabel pdiffusion 479 -3385 479 -3385 0 feedthrough
rlabel pdiffusion 486 -3385 486 -3385 0 feedthrough
rlabel pdiffusion 493 -3385 493 -3385 0 feedthrough
rlabel pdiffusion 500 -3385 500 -3385 0 feedthrough
rlabel pdiffusion 507 -3385 507 -3385 0 feedthrough
rlabel pdiffusion 514 -3385 514 -3385 0 feedthrough
rlabel pdiffusion 521 -3385 521 -3385 0 feedthrough
rlabel pdiffusion 528 -3385 528 -3385 0 feedthrough
rlabel pdiffusion 535 -3385 535 -3385 0 feedthrough
rlabel pdiffusion 542 -3385 542 -3385 0 cellNo=115
rlabel pdiffusion 549 -3385 549 -3385 0 feedthrough
rlabel pdiffusion 556 -3385 556 -3385 0 cellNo=959
rlabel pdiffusion 563 -3385 563 -3385 0 feedthrough
rlabel pdiffusion 570 -3385 570 -3385 0 cellNo=186
rlabel pdiffusion 577 -3385 577 -3385 0 cellNo=886
rlabel pdiffusion 584 -3385 584 -3385 0 feedthrough
rlabel pdiffusion 591 -3385 591 -3385 0 feedthrough
rlabel pdiffusion 598 -3385 598 -3385 0 feedthrough
rlabel pdiffusion 605 -3385 605 -3385 0 feedthrough
rlabel pdiffusion 612 -3385 612 -3385 0 feedthrough
rlabel pdiffusion 619 -3385 619 -3385 0 feedthrough
rlabel pdiffusion 626 -3385 626 -3385 0 feedthrough
rlabel pdiffusion 633 -3385 633 -3385 0 feedthrough
rlabel pdiffusion 640 -3385 640 -3385 0 feedthrough
rlabel pdiffusion 647 -3385 647 -3385 0 feedthrough
rlabel pdiffusion 654 -3385 654 -3385 0 cellNo=921
rlabel pdiffusion 661 -3385 661 -3385 0 feedthrough
rlabel pdiffusion 668 -3385 668 -3385 0 feedthrough
rlabel pdiffusion 675 -3385 675 -3385 0 feedthrough
rlabel pdiffusion 682 -3385 682 -3385 0 feedthrough
rlabel pdiffusion 689 -3385 689 -3385 0 feedthrough
rlabel pdiffusion 696 -3385 696 -3385 0 feedthrough
rlabel pdiffusion 703 -3385 703 -3385 0 feedthrough
rlabel pdiffusion 710 -3385 710 -3385 0 feedthrough
rlabel pdiffusion 717 -3385 717 -3385 0 feedthrough
rlabel pdiffusion 724 -3385 724 -3385 0 feedthrough
rlabel pdiffusion 731 -3385 731 -3385 0 feedthrough
rlabel pdiffusion 738 -3385 738 -3385 0 feedthrough
rlabel pdiffusion 745 -3385 745 -3385 0 feedthrough
rlabel pdiffusion 752 -3385 752 -3385 0 feedthrough
rlabel pdiffusion 759 -3385 759 -3385 0 cellNo=170
rlabel pdiffusion 766 -3385 766 -3385 0 feedthrough
rlabel pdiffusion 773 -3385 773 -3385 0 feedthrough
rlabel pdiffusion 780 -3385 780 -3385 0 feedthrough
rlabel pdiffusion 787 -3385 787 -3385 0 feedthrough
rlabel pdiffusion 794 -3385 794 -3385 0 cellNo=631
rlabel pdiffusion 801 -3385 801 -3385 0 feedthrough
rlabel pdiffusion 808 -3385 808 -3385 0 feedthrough
rlabel pdiffusion 815 -3385 815 -3385 0 feedthrough
rlabel pdiffusion 822 -3385 822 -3385 0 feedthrough
rlabel pdiffusion 829 -3385 829 -3385 0 feedthrough
rlabel pdiffusion 836 -3385 836 -3385 0 feedthrough
rlabel pdiffusion 843 -3385 843 -3385 0 feedthrough
rlabel pdiffusion 850 -3385 850 -3385 0 feedthrough
rlabel pdiffusion 857 -3385 857 -3385 0 feedthrough
rlabel pdiffusion 864 -3385 864 -3385 0 feedthrough
rlabel pdiffusion 871 -3385 871 -3385 0 feedthrough
rlabel pdiffusion 878 -3385 878 -3385 0 feedthrough
rlabel pdiffusion 885 -3385 885 -3385 0 feedthrough
rlabel pdiffusion 892 -3385 892 -3385 0 feedthrough
rlabel pdiffusion 899 -3385 899 -3385 0 feedthrough
rlabel pdiffusion 906 -3385 906 -3385 0 feedthrough
rlabel pdiffusion 913 -3385 913 -3385 0 feedthrough
rlabel pdiffusion 920 -3385 920 -3385 0 feedthrough
rlabel pdiffusion 927 -3385 927 -3385 0 feedthrough
rlabel pdiffusion 934 -3385 934 -3385 0 feedthrough
rlabel pdiffusion 941 -3385 941 -3385 0 feedthrough
rlabel pdiffusion 948 -3385 948 -3385 0 feedthrough
rlabel pdiffusion 955 -3385 955 -3385 0 cellNo=440
rlabel pdiffusion 962 -3385 962 -3385 0 feedthrough
rlabel pdiffusion 969 -3385 969 -3385 0 feedthrough
rlabel pdiffusion 976 -3385 976 -3385 0 feedthrough
rlabel pdiffusion 983 -3385 983 -3385 0 feedthrough
rlabel pdiffusion 990 -3385 990 -3385 0 feedthrough
rlabel pdiffusion 997 -3385 997 -3385 0 feedthrough
rlabel pdiffusion 1004 -3385 1004 -3385 0 feedthrough
rlabel pdiffusion 1011 -3385 1011 -3385 0 cellNo=240
rlabel pdiffusion 1018 -3385 1018 -3385 0 feedthrough
rlabel pdiffusion 1025 -3385 1025 -3385 0 feedthrough
rlabel pdiffusion 1032 -3385 1032 -3385 0 feedthrough
rlabel pdiffusion 1039 -3385 1039 -3385 0 cellNo=92
rlabel pdiffusion 1046 -3385 1046 -3385 0 feedthrough
rlabel pdiffusion 1053 -3385 1053 -3385 0 cellNo=587
rlabel pdiffusion 1060 -3385 1060 -3385 0 feedthrough
rlabel pdiffusion 1067 -3385 1067 -3385 0 cellNo=918
rlabel pdiffusion 1074 -3385 1074 -3385 0 feedthrough
rlabel pdiffusion 1081 -3385 1081 -3385 0 feedthrough
rlabel pdiffusion 1088 -3385 1088 -3385 0 feedthrough
rlabel pdiffusion 1095 -3385 1095 -3385 0 feedthrough
rlabel pdiffusion 1102 -3385 1102 -3385 0 feedthrough
rlabel pdiffusion 1123 -3385 1123 -3385 0 feedthrough
rlabel pdiffusion 1130 -3385 1130 -3385 0 feedthrough
rlabel pdiffusion 1179 -3385 1179 -3385 0 cellNo=960
rlabel pdiffusion 1186 -3385 1186 -3385 0 feedthrough
rlabel pdiffusion 1193 -3385 1193 -3385 0 feedthrough
rlabel pdiffusion 1340 -3385 1340 -3385 0 feedthrough
rlabel pdiffusion 1347 -3385 1347 -3385 0 feedthrough
rlabel pdiffusion 1354 -3385 1354 -3385 0 feedthrough
rlabel pdiffusion 3 -3448 3 -3448 0 cellNo=1261
rlabel pdiffusion 10 -3448 10 -3448 0 cellNo=1262
rlabel pdiffusion 17 -3448 17 -3448 0 cellNo=1263
rlabel pdiffusion 24 -3448 24 -3448 0 cellNo=1264
rlabel pdiffusion 31 -3448 31 -3448 0 cellNo=1265
rlabel pdiffusion 38 -3448 38 -3448 0 cellNo=1266
rlabel pdiffusion 45 -3448 45 -3448 0 cellNo=1267
rlabel pdiffusion 52 -3448 52 -3448 0 cellNo=1268
rlabel pdiffusion 59 -3448 59 -3448 0 cellNo=1269
rlabel pdiffusion 66 -3448 66 -3448 0 cellNo=1270
rlabel pdiffusion 73 -3448 73 -3448 0 cellNo=1271
rlabel pdiffusion 80 -3448 80 -3448 0 cellNo=1272
rlabel pdiffusion 87 -3448 87 -3448 0 cellNo=1273
rlabel pdiffusion 94 -3448 94 -3448 0 cellNo=1274
rlabel pdiffusion 101 -3448 101 -3448 0 cellNo=1278
rlabel pdiffusion 108 -3448 108 -3448 0 cellNo=1320
rlabel pdiffusion 248 -3448 248 -3448 0 feedthrough
rlabel pdiffusion 262 -3448 262 -3448 0 feedthrough
rlabel pdiffusion 290 -3448 290 -3448 0 cellNo=85
rlabel pdiffusion 311 -3448 311 -3448 0 feedthrough
rlabel pdiffusion 318 -3448 318 -3448 0 feedthrough
rlabel pdiffusion 325 -3448 325 -3448 0 feedthrough
rlabel pdiffusion 332 -3448 332 -3448 0 feedthrough
rlabel pdiffusion 339 -3448 339 -3448 0 feedthrough
rlabel pdiffusion 346 -3448 346 -3448 0 cellNo=142
rlabel pdiffusion 353 -3448 353 -3448 0 feedthrough
rlabel pdiffusion 360 -3448 360 -3448 0 feedthrough
rlabel pdiffusion 367 -3448 367 -3448 0 cellNo=712
rlabel pdiffusion 374 -3448 374 -3448 0 feedthrough
rlabel pdiffusion 381 -3448 381 -3448 0 feedthrough
rlabel pdiffusion 388 -3448 388 -3448 0 feedthrough
rlabel pdiffusion 395 -3448 395 -3448 0 feedthrough
rlabel pdiffusion 402 -3448 402 -3448 0 feedthrough
rlabel pdiffusion 409 -3448 409 -3448 0 feedthrough
rlabel pdiffusion 416 -3448 416 -3448 0 feedthrough
rlabel pdiffusion 423 -3448 423 -3448 0 feedthrough
rlabel pdiffusion 430 -3448 430 -3448 0 feedthrough
rlabel pdiffusion 437 -3448 437 -3448 0 feedthrough
rlabel pdiffusion 444 -3448 444 -3448 0 cellNo=166
rlabel pdiffusion 451 -3448 451 -3448 0 feedthrough
rlabel pdiffusion 458 -3448 458 -3448 0 feedthrough
rlabel pdiffusion 465 -3448 465 -3448 0 feedthrough
rlabel pdiffusion 472 -3448 472 -3448 0 feedthrough
rlabel pdiffusion 479 -3448 479 -3448 0 feedthrough
rlabel pdiffusion 486 -3448 486 -3448 0 feedthrough
rlabel pdiffusion 493 -3448 493 -3448 0 feedthrough
rlabel pdiffusion 500 -3448 500 -3448 0 cellNo=450
rlabel pdiffusion 507 -3448 507 -3448 0 feedthrough
rlabel pdiffusion 514 -3448 514 -3448 0 feedthrough
rlabel pdiffusion 521 -3448 521 -3448 0 feedthrough
rlabel pdiffusion 528 -3448 528 -3448 0 cellNo=510
rlabel pdiffusion 535 -3448 535 -3448 0 feedthrough
rlabel pdiffusion 542 -3448 542 -3448 0 feedthrough
rlabel pdiffusion 549 -3448 549 -3448 0 cellNo=9
rlabel pdiffusion 556 -3448 556 -3448 0 feedthrough
rlabel pdiffusion 563 -3448 563 -3448 0 feedthrough
rlabel pdiffusion 570 -3448 570 -3448 0 feedthrough
rlabel pdiffusion 577 -3448 577 -3448 0 feedthrough
rlabel pdiffusion 584 -3448 584 -3448 0 cellNo=706
rlabel pdiffusion 591 -3448 591 -3448 0 feedthrough
rlabel pdiffusion 598 -3448 598 -3448 0 feedthrough
rlabel pdiffusion 605 -3448 605 -3448 0 feedthrough
rlabel pdiffusion 612 -3448 612 -3448 0 feedthrough
rlabel pdiffusion 619 -3448 619 -3448 0 feedthrough
rlabel pdiffusion 626 -3448 626 -3448 0 feedthrough
rlabel pdiffusion 633 -3448 633 -3448 0 feedthrough
rlabel pdiffusion 640 -3448 640 -3448 0 feedthrough
rlabel pdiffusion 647 -3448 647 -3448 0 cellNo=37
rlabel pdiffusion 654 -3448 654 -3448 0 feedthrough
rlabel pdiffusion 661 -3448 661 -3448 0 feedthrough
rlabel pdiffusion 668 -3448 668 -3448 0 feedthrough
rlabel pdiffusion 675 -3448 675 -3448 0 feedthrough
rlabel pdiffusion 682 -3448 682 -3448 0 feedthrough
rlabel pdiffusion 689 -3448 689 -3448 0 cellNo=995
rlabel pdiffusion 696 -3448 696 -3448 0 feedthrough
rlabel pdiffusion 703 -3448 703 -3448 0 feedthrough
rlabel pdiffusion 710 -3448 710 -3448 0 feedthrough
rlabel pdiffusion 717 -3448 717 -3448 0 feedthrough
rlabel pdiffusion 724 -3448 724 -3448 0 feedthrough
rlabel pdiffusion 731 -3448 731 -3448 0 feedthrough
rlabel pdiffusion 738 -3448 738 -3448 0 cellNo=425
rlabel pdiffusion 745 -3448 745 -3448 0 feedthrough
rlabel pdiffusion 752 -3448 752 -3448 0 feedthrough
rlabel pdiffusion 759 -3448 759 -3448 0 feedthrough
rlabel pdiffusion 766 -3448 766 -3448 0 feedthrough
rlabel pdiffusion 773 -3448 773 -3448 0 feedthrough
rlabel pdiffusion 780 -3448 780 -3448 0 feedthrough
rlabel pdiffusion 787 -3448 787 -3448 0 feedthrough
rlabel pdiffusion 794 -3448 794 -3448 0 feedthrough
rlabel pdiffusion 801 -3448 801 -3448 0 feedthrough
rlabel pdiffusion 808 -3448 808 -3448 0 feedthrough
rlabel pdiffusion 815 -3448 815 -3448 0 feedthrough
rlabel pdiffusion 822 -3448 822 -3448 0 cellNo=417
rlabel pdiffusion 829 -3448 829 -3448 0 feedthrough
rlabel pdiffusion 836 -3448 836 -3448 0 feedthrough
rlabel pdiffusion 843 -3448 843 -3448 0 feedthrough
rlabel pdiffusion 850 -3448 850 -3448 0 feedthrough
rlabel pdiffusion 857 -3448 857 -3448 0 cellNo=477
rlabel pdiffusion 864 -3448 864 -3448 0 feedthrough
rlabel pdiffusion 871 -3448 871 -3448 0 cellNo=846
rlabel pdiffusion 878 -3448 878 -3448 0 feedthrough
rlabel pdiffusion 885 -3448 885 -3448 0 cellNo=953
rlabel pdiffusion 892 -3448 892 -3448 0 feedthrough
rlabel pdiffusion 899 -3448 899 -3448 0 cellNo=118
rlabel pdiffusion 906 -3448 906 -3448 0 feedthrough
rlabel pdiffusion 913 -3448 913 -3448 0 feedthrough
rlabel pdiffusion 920 -3448 920 -3448 0 feedthrough
rlabel pdiffusion 927 -3448 927 -3448 0 feedthrough
rlabel pdiffusion 934 -3448 934 -3448 0 feedthrough
rlabel pdiffusion 941 -3448 941 -3448 0 feedthrough
rlabel pdiffusion 948 -3448 948 -3448 0 feedthrough
rlabel pdiffusion 955 -3448 955 -3448 0 feedthrough
rlabel pdiffusion 962 -3448 962 -3448 0 feedthrough
rlabel pdiffusion 969 -3448 969 -3448 0 feedthrough
rlabel pdiffusion 976 -3448 976 -3448 0 feedthrough
rlabel pdiffusion 983 -3448 983 -3448 0 feedthrough
rlabel pdiffusion 1004 -3448 1004 -3448 0 feedthrough
rlabel pdiffusion 1011 -3448 1011 -3448 0 feedthrough
rlabel pdiffusion 1025 -3448 1025 -3448 0 cellNo=891
rlabel pdiffusion 1032 -3448 1032 -3448 0 feedthrough
rlabel pdiffusion 1039 -3448 1039 -3448 0 feedthrough
rlabel pdiffusion 1046 -3448 1046 -3448 0 feedthrough
rlabel pdiffusion 1088 -3448 1088 -3448 0 feedthrough
rlabel pdiffusion 1095 -3448 1095 -3448 0 feedthrough
rlabel pdiffusion 1116 -3448 1116 -3448 0 feedthrough
rlabel pdiffusion 1137 -3448 1137 -3448 0 feedthrough
rlabel pdiffusion 1179 -3448 1179 -3448 0 feedthrough
rlabel pdiffusion 1340 -3448 1340 -3448 0 feedthrough
rlabel pdiffusion 1347 -3448 1347 -3448 0 feedthrough
rlabel pdiffusion 1354 -3448 1354 -3448 0 feedthrough
rlabel pdiffusion 3 -3505 3 -3505 0 cellNo=1303
rlabel pdiffusion 10 -3505 10 -3505 0 cellNo=1304
rlabel pdiffusion 17 -3505 17 -3505 0 cellNo=1305
rlabel pdiffusion 24 -3505 24 -3505 0 cellNo=1306
rlabel pdiffusion 31 -3505 31 -3505 0 cellNo=1307
rlabel pdiffusion 38 -3505 38 -3505 0 cellNo=1308
rlabel pdiffusion 45 -3505 45 -3505 0 cellNo=1309
rlabel pdiffusion 52 -3505 52 -3505 0 cellNo=1310
rlabel pdiffusion 59 -3505 59 -3505 0 cellNo=1311
rlabel pdiffusion 66 -3505 66 -3505 0 cellNo=1312
rlabel pdiffusion 73 -3505 73 -3505 0 cellNo=1313
rlabel pdiffusion 80 -3505 80 -3505 0 cellNo=1314
rlabel pdiffusion 87 -3505 87 -3505 0 cellNo=1315
rlabel pdiffusion 94 -3505 94 -3505 0 cellNo=1316
rlabel pdiffusion 101 -3505 101 -3505 0 cellNo=1317
rlabel pdiffusion 108 -3505 108 -3505 0 cellNo=1319
rlabel pdiffusion 115 -3505 115 -3505 0 cellNo=1344
rlabel pdiffusion 248 -3505 248 -3505 0 feedthrough
rlabel pdiffusion 262 -3505 262 -3505 0 feedthrough
rlabel pdiffusion 276 -3505 276 -3505 0 feedthrough
rlabel pdiffusion 332 -3505 332 -3505 0 feedthrough
rlabel pdiffusion 339 -3505 339 -3505 0 feedthrough
rlabel pdiffusion 346 -3505 346 -3505 0 feedthrough
rlabel pdiffusion 353 -3505 353 -3505 0 feedthrough
rlabel pdiffusion 360 -3505 360 -3505 0 feedthrough
rlabel pdiffusion 367 -3505 367 -3505 0 feedthrough
rlabel pdiffusion 374 -3505 374 -3505 0 feedthrough
rlabel pdiffusion 381 -3505 381 -3505 0 feedthrough
rlabel pdiffusion 388 -3505 388 -3505 0 feedthrough
rlabel pdiffusion 395 -3505 395 -3505 0 feedthrough
rlabel pdiffusion 402 -3505 402 -3505 0 feedthrough
rlabel pdiffusion 409 -3505 409 -3505 0 feedthrough
rlabel pdiffusion 416 -3505 416 -3505 0 feedthrough
rlabel pdiffusion 423 -3505 423 -3505 0 cellNo=739
rlabel pdiffusion 430 -3505 430 -3505 0 feedthrough
rlabel pdiffusion 437 -3505 437 -3505 0 feedthrough
rlabel pdiffusion 444 -3505 444 -3505 0 feedthrough
rlabel pdiffusion 451 -3505 451 -3505 0 feedthrough
rlabel pdiffusion 458 -3505 458 -3505 0 feedthrough
rlabel pdiffusion 465 -3505 465 -3505 0 cellNo=749
rlabel pdiffusion 472 -3505 472 -3505 0 feedthrough
rlabel pdiffusion 479 -3505 479 -3505 0 feedthrough
rlabel pdiffusion 486 -3505 486 -3505 0 feedthrough
rlabel pdiffusion 493 -3505 493 -3505 0 cellNo=956
rlabel pdiffusion 500 -3505 500 -3505 0 feedthrough
rlabel pdiffusion 507 -3505 507 -3505 0 feedthrough
rlabel pdiffusion 514 -3505 514 -3505 0 feedthrough
rlabel pdiffusion 521 -3505 521 -3505 0 feedthrough
rlabel pdiffusion 528 -3505 528 -3505 0 feedthrough
rlabel pdiffusion 535 -3505 535 -3505 0 cellNo=132
rlabel pdiffusion 542 -3505 542 -3505 0 feedthrough
rlabel pdiffusion 549 -3505 549 -3505 0 feedthrough
rlabel pdiffusion 556 -3505 556 -3505 0 feedthrough
rlabel pdiffusion 563 -3505 563 -3505 0 cellNo=816
rlabel pdiffusion 570 -3505 570 -3505 0 feedthrough
rlabel pdiffusion 577 -3505 577 -3505 0 cellNo=920
rlabel pdiffusion 584 -3505 584 -3505 0 feedthrough
rlabel pdiffusion 591 -3505 591 -3505 0 feedthrough
rlabel pdiffusion 598 -3505 598 -3505 0 feedthrough
rlabel pdiffusion 605 -3505 605 -3505 0 feedthrough
rlabel pdiffusion 612 -3505 612 -3505 0 feedthrough
rlabel pdiffusion 619 -3505 619 -3505 0 feedthrough
rlabel pdiffusion 626 -3505 626 -3505 0 cellNo=916
rlabel pdiffusion 633 -3505 633 -3505 0 feedthrough
rlabel pdiffusion 640 -3505 640 -3505 0 cellNo=592
rlabel pdiffusion 647 -3505 647 -3505 0 feedthrough
rlabel pdiffusion 654 -3505 654 -3505 0 feedthrough
rlabel pdiffusion 661 -3505 661 -3505 0 feedthrough
rlabel pdiffusion 668 -3505 668 -3505 0 feedthrough
rlabel pdiffusion 675 -3505 675 -3505 0 cellNo=853
rlabel pdiffusion 682 -3505 682 -3505 0 feedthrough
rlabel pdiffusion 689 -3505 689 -3505 0 feedthrough
rlabel pdiffusion 696 -3505 696 -3505 0 feedthrough
rlabel pdiffusion 703 -3505 703 -3505 0 feedthrough
rlabel pdiffusion 710 -3505 710 -3505 0 feedthrough
rlabel pdiffusion 717 -3505 717 -3505 0 feedthrough
rlabel pdiffusion 724 -3505 724 -3505 0 cellNo=71
rlabel pdiffusion 731 -3505 731 -3505 0 feedthrough
rlabel pdiffusion 738 -3505 738 -3505 0 feedthrough
rlabel pdiffusion 745 -3505 745 -3505 0 feedthrough
rlabel pdiffusion 752 -3505 752 -3505 0 feedthrough
rlabel pdiffusion 759 -3505 759 -3505 0 feedthrough
rlabel pdiffusion 766 -3505 766 -3505 0 feedthrough
rlabel pdiffusion 773 -3505 773 -3505 0 feedthrough
rlabel pdiffusion 780 -3505 780 -3505 0 feedthrough
rlabel pdiffusion 801 -3505 801 -3505 0 feedthrough
rlabel pdiffusion 808 -3505 808 -3505 0 feedthrough
rlabel pdiffusion 815 -3505 815 -3505 0 cellNo=40
rlabel pdiffusion 822 -3505 822 -3505 0 feedthrough
rlabel pdiffusion 836 -3505 836 -3505 0 feedthrough
rlabel pdiffusion 843 -3505 843 -3505 0 feedthrough
rlabel pdiffusion 850 -3505 850 -3505 0 feedthrough
rlabel pdiffusion 857 -3505 857 -3505 0 feedthrough
rlabel pdiffusion 864 -3505 864 -3505 0 feedthrough
rlabel pdiffusion 871 -3505 871 -3505 0 feedthrough
rlabel pdiffusion 878 -3505 878 -3505 0 feedthrough
rlabel pdiffusion 906 -3505 906 -3505 0 feedthrough
rlabel pdiffusion 913 -3505 913 -3505 0 feedthrough
rlabel pdiffusion 920 -3505 920 -3505 0 feedthrough
rlabel pdiffusion 927 -3505 927 -3505 0 feedthrough
rlabel pdiffusion 934 -3505 934 -3505 0 feedthrough
rlabel pdiffusion 941 -3505 941 -3505 0 feedthrough
rlabel pdiffusion 948 -3505 948 -3505 0 feedthrough
rlabel pdiffusion 955 -3505 955 -3505 0 cellNo=681
rlabel pdiffusion 962 -3505 962 -3505 0 feedthrough
rlabel pdiffusion 969 -3505 969 -3505 0 feedthrough
rlabel pdiffusion 983 -3505 983 -3505 0 feedthrough
rlabel pdiffusion 990 -3505 990 -3505 0 feedthrough
rlabel pdiffusion 997 -3505 997 -3505 0 cellNo=897
rlabel pdiffusion 1004 -3505 1004 -3505 0 feedthrough
rlabel pdiffusion 1011 -3505 1011 -3505 0 feedthrough
rlabel pdiffusion 1053 -3505 1053 -3505 0 feedthrough
rlabel pdiffusion 1081 -3505 1081 -3505 0 feedthrough
rlabel pdiffusion 1088 -3505 1088 -3505 0 feedthrough
rlabel pdiffusion 1109 -3505 1109 -3505 0 feedthrough
rlabel pdiffusion 1123 -3505 1123 -3505 0 feedthrough
rlabel pdiffusion 1151 -3505 1151 -3505 0 feedthrough
rlabel pdiffusion 1172 -3505 1172 -3505 0 cellNo=513
rlabel pdiffusion 1179 -3505 1179 -3505 0 feedthrough
rlabel pdiffusion 1340 -3505 1340 -3505 0 feedthrough
rlabel pdiffusion 1347 -3505 1347 -3505 0 cellNo=661
rlabel pdiffusion 1354 -3505 1354 -3505 0 feedthrough
rlabel pdiffusion 3 -3546 3 -3546 0 cellNo=1345
rlabel pdiffusion 10 -3546 10 -3546 0 cellNo=1346
rlabel pdiffusion 17 -3546 17 -3546 0 cellNo=1347
rlabel pdiffusion 24 -3546 24 -3546 0 cellNo=1348
rlabel pdiffusion 31 -3546 31 -3546 0 cellNo=1349
rlabel pdiffusion 38 -3546 38 -3546 0 cellNo=1350
rlabel pdiffusion 45 -3546 45 -3546 0 cellNo=1351
rlabel pdiffusion 52 -3546 52 -3546 0 cellNo=1352
rlabel pdiffusion 59 -3546 59 -3546 0 cellNo=1353
rlabel pdiffusion 66 -3546 66 -3546 0 cellNo=1354
rlabel pdiffusion 73 -3546 73 -3546 0 cellNo=1355
rlabel pdiffusion 80 -3546 80 -3546 0 cellNo=1356
rlabel pdiffusion 87 -3546 87 -3546 0 cellNo=1357
rlabel pdiffusion 94 -3546 94 -3546 0 cellNo=1358
rlabel pdiffusion 101 -3546 101 -3546 0 cellNo=1359
rlabel pdiffusion 108 -3546 108 -3546 0 cellNo=1360
rlabel pdiffusion 115 -3546 115 -3546 0 cellNo=1380
rlabel pdiffusion 122 -3546 122 -3546 0 cellNo=1419
rlabel pdiffusion 248 -3546 248 -3546 0 feedthrough
rlabel pdiffusion 255 -3546 255 -3546 0 cellNo=562
rlabel pdiffusion 262 -3546 262 -3546 0 feedthrough
rlabel pdiffusion 269 -3546 269 -3546 0 feedthrough
rlabel pdiffusion 297 -3546 297 -3546 0 feedthrough
rlabel pdiffusion 346 -3546 346 -3546 0 feedthrough
rlabel pdiffusion 360 -3546 360 -3546 0 feedthrough
rlabel pdiffusion 381 -3546 381 -3546 0 feedthrough
rlabel pdiffusion 395 -3546 395 -3546 0 feedthrough
rlabel pdiffusion 402 -3546 402 -3546 0 feedthrough
rlabel pdiffusion 409 -3546 409 -3546 0 feedthrough
rlabel pdiffusion 416 -3546 416 -3546 0 feedthrough
rlabel pdiffusion 423 -3546 423 -3546 0 feedthrough
rlabel pdiffusion 430 -3546 430 -3546 0 cellNo=943
rlabel pdiffusion 437 -3546 437 -3546 0 feedthrough
rlabel pdiffusion 444 -3546 444 -3546 0 cellNo=648
rlabel pdiffusion 451 -3546 451 -3546 0 cellNo=324
rlabel pdiffusion 458 -3546 458 -3546 0 feedthrough
rlabel pdiffusion 465 -3546 465 -3546 0 feedthrough
rlabel pdiffusion 472 -3546 472 -3546 0 feedthrough
rlabel pdiffusion 479 -3546 479 -3546 0 feedthrough
rlabel pdiffusion 486 -3546 486 -3546 0 cellNo=948
rlabel pdiffusion 493 -3546 493 -3546 0 feedthrough
rlabel pdiffusion 500 -3546 500 -3546 0 feedthrough
rlabel pdiffusion 507 -3546 507 -3546 0 feedthrough
rlabel pdiffusion 514 -3546 514 -3546 0 feedthrough
rlabel pdiffusion 521 -3546 521 -3546 0 feedthrough
rlabel pdiffusion 528 -3546 528 -3546 0 feedthrough
rlabel pdiffusion 535 -3546 535 -3546 0 feedthrough
rlabel pdiffusion 542 -3546 542 -3546 0 cellNo=65
rlabel pdiffusion 549 -3546 549 -3546 0 feedthrough
rlabel pdiffusion 556 -3546 556 -3546 0 feedthrough
rlabel pdiffusion 563 -3546 563 -3546 0 feedthrough
rlabel pdiffusion 570 -3546 570 -3546 0 feedthrough
rlabel pdiffusion 577 -3546 577 -3546 0 feedthrough
rlabel pdiffusion 584 -3546 584 -3546 0 feedthrough
rlabel pdiffusion 591 -3546 591 -3546 0 feedthrough
rlabel pdiffusion 598 -3546 598 -3546 0 cellNo=183
rlabel pdiffusion 605 -3546 605 -3546 0 feedthrough
rlabel pdiffusion 612 -3546 612 -3546 0 feedthrough
rlabel pdiffusion 626 -3546 626 -3546 0 cellNo=840
rlabel pdiffusion 640 -3546 640 -3546 0 feedthrough
rlabel pdiffusion 668 -3546 668 -3546 0 feedthrough
rlabel pdiffusion 682 -3546 682 -3546 0 feedthrough
rlabel pdiffusion 689 -3546 689 -3546 0 cellNo=865
rlabel pdiffusion 696 -3546 696 -3546 0 feedthrough
rlabel pdiffusion 703 -3546 703 -3546 0 feedthrough
rlabel pdiffusion 710 -3546 710 -3546 0 feedthrough
rlabel pdiffusion 717 -3546 717 -3546 0 feedthrough
rlabel pdiffusion 724 -3546 724 -3546 0 feedthrough
rlabel pdiffusion 731 -3546 731 -3546 0 feedthrough
rlabel pdiffusion 738 -3546 738 -3546 0 feedthrough
rlabel pdiffusion 745 -3546 745 -3546 0 feedthrough
rlabel pdiffusion 752 -3546 752 -3546 0 feedthrough
rlabel pdiffusion 759 -3546 759 -3546 0 feedthrough
rlabel pdiffusion 766 -3546 766 -3546 0 feedthrough
rlabel pdiffusion 836 -3546 836 -3546 0 feedthrough
rlabel pdiffusion 850 -3546 850 -3546 0 feedthrough
rlabel pdiffusion 864 -3546 864 -3546 0 feedthrough
rlabel pdiffusion 871 -3546 871 -3546 0 feedthrough
rlabel pdiffusion 878 -3546 878 -3546 0 feedthrough
rlabel pdiffusion 885 -3546 885 -3546 0 feedthrough
rlabel pdiffusion 892 -3546 892 -3546 0 feedthrough
rlabel pdiffusion 899 -3546 899 -3546 0 feedthrough
rlabel pdiffusion 906 -3546 906 -3546 0 feedthrough
rlabel pdiffusion 913 -3546 913 -3546 0 feedthrough
rlabel pdiffusion 920 -3546 920 -3546 0 cellNo=42
rlabel pdiffusion 927 -3546 927 -3546 0 feedthrough
rlabel pdiffusion 934 -3546 934 -3546 0 cellNo=380
rlabel pdiffusion 941 -3546 941 -3546 0 cellNo=968
rlabel pdiffusion 948 -3546 948 -3546 0 feedthrough
rlabel pdiffusion 969 -3546 969 -3546 0 feedthrough
rlabel pdiffusion 976 -3546 976 -3546 0 feedthrough
rlabel pdiffusion 990 -3546 990 -3546 0 feedthrough
rlabel pdiffusion 1004 -3546 1004 -3546 0 cellNo=826
rlabel pdiffusion 1011 -3546 1011 -3546 0 feedthrough
rlabel pdiffusion 1053 -3546 1053 -3546 0 feedthrough
rlabel pdiffusion 1060 -3546 1060 -3546 0 feedthrough
rlabel pdiffusion 1081 -3546 1081 -3546 0 feedthrough
rlabel pdiffusion 1109 -3546 1109 -3546 0 feedthrough
rlabel pdiffusion 1151 -3546 1151 -3546 0 feedthrough
rlabel pdiffusion 1158 -3546 1158 -3546 0 cellNo=719
rlabel pdiffusion 3 -3583 3 -3583 0 cellNo=1387
rlabel pdiffusion 10 -3583 10 -3583 0 cellNo=1388
rlabel pdiffusion 17 -3583 17 -3583 0 cellNo=1389
rlabel pdiffusion 24 -3583 24 -3583 0 cellNo=1390
rlabel pdiffusion 31 -3583 31 -3583 0 cellNo=1391
rlabel pdiffusion 38 -3583 38 -3583 0 cellNo=1392
rlabel pdiffusion 45 -3583 45 -3583 0 cellNo=1393
rlabel pdiffusion 52 -3583 52 -3583 0 cellNo=1394
rlabel pdiffusion 59 -3583 59 -3583 0 cellNo=1395
rlabel pdiffusion 66 -3583 66 -3583 0 cellNo=1396
rlabel pdiffusion 73 -3583 73 -3583 0 cellNo=1397
rlabel pdiffusion 80 -3583 80 -3583 0 cellNo=1398
rlabel pdiffusion 87 -3583 87 -3583 0 cellNo=1399
rlabel pdiffusion 94 -3583 94 -3583 0 cellNo=1400
rlabel pdiffusion 101 -3583 101 -3583 0 cellNo=1401
rlabel pdiffusion 108 -3583 108 -3583 0 cellNo=1402
rlabel pdiffusion 115 -3583 115 -3583 0 cellNo=1412
rlabel pdiffusion 122 -3583 122 -3583 0 cellNo=1448
rlabel pdiffusion 262 -3583 262 -3583 0 cellNo=405
rlabel pdiffusion 269 -3583 269 -3583 0 feedthrough
rlabel pdiffusion 311 -3583 311 -3583 0 feedthrough
rlabel pdiffusion 325 -3583 325 -3583 0 cellNo=621
rlabel pdiffusion 353 -3583 353 -3583 0 feedthrough
rlabel pdiffusion 360 -3583 360 -3583 0 feedthrough
rlabel pdiffusion 367 -3583 367 -3583 0 feedthrough
rlabel pdiffusion 374 -3583 374 -3583 0 cellNo=102
rlabel pdiffusion 395 -3583 395 -3583 0 feedthrough
rlabel pdiffusion 402 -3583 402 -3583 0 cellNo=863
rlabel pdiffusion 409 -3583 409 -3583 0 feedthrough
rlabel pdiffusion 416 -3583 416 -3583 0 feedthrough
rlabel pdiffusion 437 -3583 437 -3583 0 feedthrough
rlabel pdiffusion 444 -3583 444 -3583 0 cellNo=43
rlabel pdiffusion 451 -3583 451 -3583 0 cellNo=427
rlabel pdiffusion 458 -3583 458 -3583 0 feedthrough
rlabel pdiffusion 465 -3583 465 -3583 0 feedthrough
rlabel pdiffusion 472 -3583 472 -3583 0 feedthrough
rlabel pdiffusion 479 -3583 479 -3583 0 feedthrough
rlabel pdiffusion 486 -3583 486 -3583 0 cellNo=148
rlabel pdiffusion 493 -3583 493 -3583 0 feedthrough
rlabel pdiffusion 500 -3583 500 -3583 0 feedthrough
rlabel pdiffusion 507 -3583 507 -3583 0 feedthrough
rlabel pdiffusion 514 -3583 514 -3583 0 cellNo=486
rlabel pdiffusion 521 -3583 521 -3583 0 feedthrough
rlabel pdiffusion 528 -3583 528 -3583 0 feedthrough
rlabel pdiffusion 535 -3583 535 -3583 0 feedthrough
rlabel pdiffusion 542 -3583 542 -3583 0 feedthrough
rlabel pdiffusion 549 -3583 549 -3583 0 feedthrough
rlabel pdiffusion 556 -3583 556 -3583 0 feedthrough
rlabel pdiffusion 563 -3583 563 -3583 0 feedthrough
rlabel pdiffusion 570 -3583 570 -3583 0 feedthrough
rlabel pdiffusion 598 -3583 598 -3583 0 feedthrough
rlabel pdiffusion 612 -3583 612 -3583 0 feedthrough
rlabel pdiffusion 619 -3583 619 -3583 0 feedthrough
rlabel pdiffusion 647 -3583 647 -3583 0 feedthrough
rlabel pdiffusion 661 -3583 661 -3583 0 feedthrough
rlabel pdiffusion 675 -3583 675 -3583 0 cellNo=489
rlabel pdiffusion 689 -3583 689 -3583 0 feedthrough
rlabel pdiffusion 696 -3583 696 -3583 0 feedthrough
rlabel pdiffusion 703 -3583 703 -3583 0 feedthrough
rlabel pdiffusion 710 -3583 710 -3583 0 feedthrough
rlabel pdiffusion 717 -3583 717 -3583 0 feedthrough
rlabel pdiffusion 724 -3583 724 -3583 0 feedthrough
rlabel pdiffusion 731 -3583 731 -3583 0 feedthrough
rlabel pdiffusion 738 -3583 738 -3583 0 feedthrough
rlabel pdiffusion 745 -3583 745 -3583 0 feedthrough
rlabel pdiffusion 752 -3583 752 -3583 0 feedthrough
rlabel pdiffusion 759 -3583 759 -3583 0 feedthrough
rlabel pdiffusion 766 -3583 766 -3583 0 feedthrough
rlabel pdiffusion 850 -3583 850 -3583 0 feedthrough
rlabel pdiffusion 857 -3583 857 -3583 0 feedthrough
rlabel pdiffusion 892 -3583 892 -3583 0 feedthrough
rlabel pdiffusion 899 -3583 899 -3583 0 cellNo=788
rlabel pdiffusion 906 -3583 906 -3583 0 feedthrough
rlabel pdiffusion 913 -3583 913 -3583 0 feedthrough
rlabel pdiffusion 920 -3583 920 -3583 0 cellNo=588
rlabel pdiffusion 927 -3583 927 -3583 0 feedthrough
rlabel pdiffusion 941 -3583 941 -3583 0 feedthrough
rlabel pdiffusion 969 -3583 969 -3583 0 feedthrough
rlabel pdiffusion 976 -3583 976 -3583 0 feedthrough
rlabel pdiffusion 983 -3583 983 -3583 0 cellNo=979
rlabel pdiffusion 990 -3583 990 -3583 0 feedthrough
rlabel pdiffusion 1039 -3583 1039 -3583 0 feedthrough
rlabel pdiffusion 1053 -3583 1053 -3583 0 feedthrough
rlabel pdiffusion 1081 -3583 1081 -3583 0 cellNo=435
rlabel pdiffusion 1088 -3583 1088 -3583 0 feedthrough
rlabel pdiffusion 1109 -3583 1109 -3583 0 feedthrough
rlabel pdiffusion 3 -3606 3 -3606 0 cellNo=1429
rlabel pdiffusion 10 -3606 10 -3606 0 cellNo=1430
rlabel pdiffusion 17 -3606 17 -3606 0 cellNo=1431
rlabel pdiffusion 24 -3606 24 -3606 0 cellNo=1432
rlabel pdiffusion 31 -3606 31 -3606 0 cellNo=1433
rlabel pdiffusion 38 -3606 38 -3606 0 cellNo=1434
rlabel pdiffusion 45 -3606 45 -3606 0 cellNo=1435
rlabel pdiffusion 52 -3606 52 -3606 0 cellNo=1436
rlabel pdiffusion 59 -3606 59 -3606 0 cellNo=1437
rlabel pdiffusion 66 -3606 66 -3606 0 cellNo=1438
rlabel pdiffusion 73 -3606 73 -3606 0 cellNo=1439
rlabel pdiffusion 80 -3606 80 -3606 0 cellNo=1440
rlabel pdiffusion 87 -3606 87 -3606 0 cellNo=1441
rlabel pdiffusion 94 -3606 94 -3606 0 cellNo=1442
rlabel pdiffusion 101 -3606 101 -3606 0 cellNo=1443
rlabel pdiffusion 108 -3606 108 -3606 0 cellNo=1444
rlabel pdiffusion 115 -3606 115 -3606 0 cellNo=1447
rlabel pdiffusion 122 -3606 122 -3606 0 cellNo=1466
rlabel pdiffusion 129 -3606 129 -3606 0 cellNo=1465
rlabel pdiffusion 136 -3606 136 -3606 0 cellNo=1452
rlabel pdiffusion 143 -3606 143 -3606 0 cellNo=1453
rlabel pdiffusion 150 -3606 150 -3606 0 cellNo=1456
rlabel pdiffusion 157 -3606 157 -3606 0 cellNo=1457
rlabel pdiffusion 164 -3606 164 -3606 0 cellNo=1458
rlabel pdiffusion 171 -3606 171 -3606 0 cellNo=1459
rlabel pdiffusion 178 -3606 178 -3606 0 cellNo=1460
rlabel pdiffusion 185 -3606 185 -3606 0 cellNo=1461
rlabel pdiffusion 192 -3606 192 -3606 0 cellNo=1462
rlabel pdiffusion 199 -3606 199 -3606 0 cellNo=1463
rlabel pdiffusion 206 -3606 206 -3606 0 cellNo=1464
rlabel pdiffusion 213 -3606 213 -3606 0 cellNo=1467
rlabel pdiffusion 220 -3606 220 -3606 0 cellNo=1468
rlabel pdiffusion 227 -3606 227 -3606 0 cellNo=1469
rlabel pdiffusion 234 -3606 234 -3606 0 cellNo=1470
rlabel pdiffusion 325 -3606 325 -3606 0 cellNo=354
rlabel pdiffusion 353 -3606 353 -3606 0 cellNo=854
rlabel pdiffusion 402 -3606 402 -3606 0 feedthrough
rlabel pdiffusion 409 -3606 409 -3606 0 feedthrough
rlabel pdiffusion 458 -3606 458 -3606 0 feedthrough
rlabel pdiffusion 472 -3606 472 -3606 0 feedthrough
rlabel pdiffusion 493 -3606 493 -3606 0 feedthrough
rlabel pdiffusion 507 -3606 507 -3606 0 feedthrough
rlabel pdiffusion 514 -3606 514 -3606 0 cellNo=871
rlabel pdiffusion 521 -3606 521 -3606 0 feedthrough
rlabel pdiffusion 542 -3606 542 -3606 0 cellNo=942
rlabel pdiffusion 549 -3606 549 -3606 0 feedthrough
rlabel pdiffusion 556 -3606 556 -3606 0 feedthrough
rlabel pdiffusion 563 -3606 563 -3606 0 feedthrough
rlabel pdiffusion 570 -3606 570 -3606 0 feedthrough
rlabel pdiffusion 577 -3606 577 -3606 0 feedthrough
rlabel pdiffusion 598 -3606 598 -3606 0 feedthrough
rlabel pdiffusion 605 -3606 605 -3606 0 feedthrough
rlabel pdiffusion 612 -3606 612 -3606 0 cellNo=971
rlabel pdiffusion 682 -3606 682 -3606 0 cellNo=515
rlabel pdiffusion 696 -3606 696 -3606 0 feedthrough
rlabel pdiffusion 703 -3606 703 -3606 0 feedthrough
rlabel pdiffusion 710 -3606 710 -3606 0 feedthrough
rlabel pdiffusion 717 -3606 717 -3606 0 feedthrough
rlabel pdiffusion 724 -3606 724 -3606 0 feedthrough
rlabel pdiffusion 731 -3606 731 -3606 0 feedthrough
rlabel pdiffusion 738 -3606 738 -3606 0 feedthrough
rlabel pdiffusion 745 -3606 745 -3606 0 feedthrough
rlabel pdiffusion 752 -3606 752 -3606 0 feedthrough
rlabel pdiffusion 759 -3606 759 -3606 0 cellNo=647
rlabel pdiffusion 766 -3606 766 -3606 0 feedthrough
rlabel pdiffusion 773 -3606 773 -3606 0 feedthrough
rlabel pdiffusion 857 -3606 857 -3606 0 feedthrough
rlabel pdiffusion 864 -3606 864 -3606 0 feedthrough
rlabel pdiffusion 906 -3606 906 -3606 0 cellNo=318
rlabel pdiffusion 920 -3606 920 -3606 0 feedthrough
rlabel pdiffusion 927 -3606 927 -3606 0 feedthrough
rlabel pdiffusion 976 -3606 976 -3606 0 feedthrough
rlabel pdiffusion 983 -3606 983 -3606 0 feedthrough
rlabel pdiffusion 1032 -3606 1032 -3606 0 feedthrough
rlabel pdiffusion 1046 -3606 1046 -3606 0 feedthrough
rlabel pdiffusion 1053 -3606 1053 -3606 0 feedthrough
rlabel pdiffusion 1109 -3606 1109 -3606 0 feedthrough
rlabel pdiffusion 3 -3631 3 -3631 0 cellNo=1471
rlabel pdiffusion 10 -3631 10 -3631 0 cellNo=1472
rlabel pdiffusion 17 -3631 17 -3631 0 cellNo=1473
rlabel pdiffusion 24 -3631 24 -3631 0 cellNo=1474
rlabel pdiffusion 31 -3631 31 -3631 0 cellNo=1475
rlabel pdiffusion 38 -3631 38 -3631 0 cellNo=1476
rlabel pdiffusion 45 -3631 45 -3631 0 cellNo=1477
rlabel pdiffusion 52 -3631 52 -3631 0 cellNo=1478
rlabel pdiffusion 59 -3631 59 -3631 0 cellNo=1479
rlabel pdiffusion 66 -3631 66 -3631 0 cellNo=1480
rlabel pdiffusion 73 -3631 73 -3631 0 cellNo=1481
rlabel pdiffusion 80 -3631 80 -3631 0 cellNo=1482
rlabel pdiffusion 87 -3631 87 -3631 0 cellNo=1483
rlabel pdiffusion 94 -3631 94 -3631 0 cellNo=1484
rlabel pdiffusion 101 -3631 101 -3631 0 cellNo=1485
rlabel pdiffusion 108 -3631 108 -3631 0 cellNo=1486
rlabel pdiffusion 115 -3631 115 -3631 0 cellNo=1487
rlabel pdiffusion 122 -3631 122 -3631 0 cellNo=1488
rlabel pdiffusion 129 -3631 129 -3631 0 cellNo=1489
rlabel pdiffusion 136 -3631 136 -3631 0 cellNo=1490
rlabel pdiffusion 143 -3631 143 -3631 0 cellNo=1491
rlabel pdiffusion 150 -3631 150 -3631 0 cellNo=1492
rlabel pdiffusion 157 -3631 157 -3631 0 cellNo=1493
rlabel pdiffusion 164 -3631 164 -3631 0 cellNo=1496
rlabel pdiffusion 171 -3631 171 -3631 0 cellNo=1497
rlabel pdiffusion 178 -3631 178 -3631 0 cellNo=1498
rlabel pdiffusion 185 -3631 185 -3631 0 cellNo=1499
rlabel pdiffusion 192 -3631 192 -3631 0 cellNo=1500
rlabel pdiffusion 402 -3631 402 -3631 0 feedthrough
rlabel pdiffusion 409 -3631 409 -3631 0 feedthrough
rlabel pdiffusion 465 -3631 465 -3631 0 feedthrough
rlabel pdiffusion 472 -3631 472 -3631 0 feedthrough
rlabel pdiffusion 528 -3631 528 -3631 0 feedthrough
rlabel pdiffusion 563 -3631 563 -3631 0 feedthrough
rlabel pdiffusion 570 -3631 570 -3631 0 feedthrough
rlabel pdiffusion 577 -3631 577 -3631 0 feedthrough
rlabel pdiffusion 584 -3631 584 -3631 0 feedthrough
rlabel pdiffusion 591 -3631 591 -3631 0 feedthrough
rlabel pdiffusion 703 -3631 703 -3631 0 feedthrough
rlabel pdiffusion 710 -3631 710 -3631 0 feedthrough
rlabel pdiffusion 717 -3631 717 -3631 0 feedthrough
rlabel pdiffusion 724 -3631 724 -3631 0 feedthrough
rlabel pdiffusion 745 -3631 745 -3631 0 feedthrough
rlabel pdiffusion 752 -3631 752 -3631 0 feedthrough
rlabel pdiffusion 759 -3631 759 -3631 0 feedthrough
rlabel pdiffusion 766 -3631 766 -3631 0 feedthrough
rlabel pdiffusion 773 -3631 773 -3631 0 cellNo=832
rlabel pdiffusion 801 -3631 801 -3631 0 feedthrough
rlabel pdiffusion 857 -3631 857 -3631 0 feedthrough
rlabel pdiffusion 864 -3631 864 -3631 0 feedthrough
rlabel pdiffusion 927 -3631 927 -3631 0 feedthrough
rlabel pdiffusion 934 -3631 934 -3631 0 feedthrough
rlabel pdiffusion 983 -3631 983 -3631 0 feedthrough
rlabel pdiffusion 1004 -3631 1004 -3631 0 feedthrough
rlabel pdiffusion 1032 -3631 1032 -3631 0 feedthrough
rlabel pdiffusion 1053 -3631 1053 -3631 0 cellNo=431
rlabel pdiffusion 1060 -3631 1060 -3631 0 feedthrough
rlabel pdiffusion 1081 -3631 1081 -3631 0 feedthrough
rlabel pdiffusion 1109 -3631 1109 -3631 0 feedthrough
rlabel pdiffusion 3 -3646 3 -3646 0 cellNo=1082
rlabel pdiffusion 10 -3646 10 -3646 0 cellNo=1086
rlabel pdiffusion 17 -3646 17 -3646 0 cellNo=1114
rlabel pdiffusion 24 -3646 24 -3646 0 cellNo=1123
rlabel pdiffusion 31 -3646 31 -3646 0 cellNo=1150
rlabel pdiffusion 38 -3646 38 -3646 0 cellNo=1168
rlabel pdiffusion 45 -3646 45 -3646 0 cellNo=1199
rlabel pdiffusion 52 -3646 52 -3646 0 cellNo=1215
rlabel pdiffusion 59 -3646 59 -3646 0 cellNo=1249
rlabel pdiffusion 66 -3646 66 -3646 0 cellNo=1277
rlabel pdiffusion 73 -3646 73 -3646 0 cellNo=1318
rlabel pdiffusion 80 -3646 80 -3646 0 cellNo=1343
rlabel pdiffusion 87 -3646 87 -3646 0 cellNo=1376
rlabel pdiffusion 94 -3646 94 -3646 0 cellNo=1411
rlabel pdiffusion 101 -3646 101 -3646 0 cellNo=1446
rlabel pdiffusion 402 -3646 402 -3646 0 feedthrough
rlabel pdiffusion 409 -3646 409 -3646 0 feedthrough
rlabel pdiffusion 465 -3646 465 -3646 0 feedthrough
rlabel pdiffusion 472 -3646 472 -3646 0 cellNo=555
rlabel pdiffusion 528 -3646 528 -3646 0 feedthrough
rlabel pdiffusion 570 -3646 570 -3646 0 cellNo=718
rlabel pdiffusion 577 -3646 577 -3646 0 feedthrough
rlabel pdiffusion 584 -3646 584 -3646 0 cellNo=764
rlabel pdiffusion 591 -3646 591 -3646 0 feedthrough
rlabel pdiffusion 598 -3646 598 -3646 0 feedthrough
rlabel pdiffusion 710 -3646 710 -3646 0 feedthrough
rlabel pdiffusion 717 -3646 717 -3646 0 cellNo=609
rlabel pdiffusion 724 -3646 724 -3646 0 feedthrough
rlabel pdiffusion 752 -3646 752 -3646 0 feedthrough
rlabel pdiffusion 759 -3646 759 -3646 0 feedthrough
rlabel pdiffusion 766 -3646 766 -3646 0 feedthrough
rlabel pdiffusion 857 -3646 857 -3646 0 cellNo=934
rlabel pdiffusion 864 -3646 864 -3646 0 feedthrough
rlabel pdiffusion 927 -3646 927 -3646 0 cellNo=429
rlabel pdiffusion 934 -3646 934 -3646 0 feedthrough
rlabel pdiffusion 983 -3646 983 -3646 0 cellNo=705
rlabel pdiffusion 990 -3646 990 -3646 0 feedthrough
rlabel pdiffusion 1032 -3646 1032 -3646 0 cellNo=789
rlabel pdiffusion 1095 -3646 1095 -3646 0 feedthrough
rlabel pdiffusion 1109 -3646 1109 -3646 0 cellNo=925
rlabel pdiffusion 3 -3661 3 -3661 0 cellNo=1085
rlabel pdiffusion 10 -3661 10 -3661 0 cellNo=1112
rlabel pdiffusion 17 -3661 17 -3661 0 cellNo=1122
rlabel pdiffusion 24 -3661 24 -3661 0 cellNo=1148
rlabel pdiffusion 31 -3661 31 -3661 0 cellNo=1166
rlabel pdiffusion 38 -3661 38 -3661 0 cellNo=1197
rlabel pdiffusion 45 -3661 45 -3661 0 cellNo=1214
rlabel pdiffusion 52 -3661 52 -3661 0 cellNo=1248
rlabel pdiffusion 59 -3661 59 -3661 0 cellNo=1259
rlabel pdiffusion 66 -3661 66 -3661 0 cellNo=1302
rlabel pdiffusion 73 -3661 73 -3661 0 cellNo=1338
rlabel pdiffusion 80 -3661 80 -3661 0 cellNo=1375
rlabel pdiffusion 87 -3661 87 -3661 0 cellNo=1410
rlabel pdiffusion 94 -3661 94 -3661 0 cellNo=1445
rlabel pdiffusion 101 -3661 101 -3661 0 cellNo=1449
rlabel pdiffusion 402 -3661 402 -3661 0 cellNo=617
rlabel pdiffusion 409 -3661 409 -3661 0 feedthrough
rlabel pdiffusion 528 -3661 528 -3661 0 cellNo=992
rlabel pdiffusion 535 -3661 535 -3661 0 feedthrough
rlabel pdiffusion 759 -3661 759 -3661 0 feedthrough
rlabel pdiffusion 766 -3661 766 -3661 0 cellNo=600
rlabel pdiffusion 773 -3661 773 -3661 0 feedthrough
rlabel pdiffusion 3 -3672 3 -3672 0 cellNo=1109
rlabel pdiffusion 10 -3672 10 -3672 0 cellNo=1121
rlabel pdiffusion 17 -3672 17 -3672 0 cellNo=1134
rlabel pdiffusion 24 -3672 24 -3672 0 cellNo=1165
rlabel pdiffusion 31 -3672 31 -3672 0 cellNo=1196
rlabel pdiffusion 38 -3672 38 -3672 0 cellNo=1213
rlabel pdiffusion 45 -3672 45 -3672 0 cellNo=1246
rlabel pdiffusion 52 -3672 52 -3672 0 cellNo=1257
rlabel pdiffusion 59 -3672 59 -3672 0 cellNo=1301
rlabel pdiffusion 66 -3672 66 -3672 0 cellNo=1336
rlabel pdiffusion 73 -3672 73 -3672 0 cellNo=1374
rlabel pdiffusion 80 -3672 80 -3672 0 cellNo=1407
rlabel pdiffusion 87 -3672 87 -3672 0 cellNo=1426
rlabel pdiffusion 3 -3681 3 -3681 0 cellNo=1120
rlabel pdiffusion 10 -3681 10 -3681 0 cellNo=1131
rlabel pdiffusion 17 -3681 17 -3681 0 cellNo=1164
rlabel pdiffusion 24 -3681 24 -3681 0 cellNo=1194
rlabel pdiffusion 31 -3681 31 -3681 0 cellNo=1212
rlabel pdiffusion 38 -3681 38 -3681 0 cellNo=1245
rlabel pdiffusion 45 -3681 45 -3681 0 cellNo=1256
rlabel pdiffusion 52 -3681 52 -3681 0 cellNo=1299
rlabel pdiffusion 59 -3681 59 -3681 0 cellNo=1332
rlabel pdiffusion 66 -3681 66 -3681 0 cellNo=1370
rlabel pdiffusion 73 -3681 73 -3681 0 cellNo=1406
rlabel pdiffusion 80 -3681 80 -3681 0 cellNo=1425
rlabel pdiffusion 87 -3681 87 -3681 0 cellNo=1495
rlabel pdiffusion 3 -3690 3 -3690 0 cellNo=1128
rlabel pdiffusion 10 -3690 10 -3690 0 cellNo=1163
rlabel pdiffusion 17 -3690 17 -3690 0 cellNo=1191
rlabel pdiffusion 24 -3690 24 -3690 0 cellNo=1209
rlabel pdiffusion 31 -3690 31 -3690 0 cellNo=1240
rlabel pdiffusion 38 -3690 38 -3690 0 cellNo=1254
rlabel pdiffusion 45 -3690 45 -3690 0 cellNo=1298
rlabel pdiffusion 52 -3690 52 -3690 0 cellNo=1326
rlabel pdiffusion 59 -3690 59 -3690 0 cellNo=1368
rlabel pdiffusion 66 -3690 66 -3690 0 cellNo=1405
rlabel pdiffusion 73 -3690 73 -3690 0 cellNo=1424
rlabel pdiffusion 80 -3690 80 -3690 0 cellNo=1450
rlabel pdiffusion 87 -3690 87 -3690 0 cellNo=1454
rlabel pdiffusion 3 -3699 3 -3699 0 cellNo=1162
rlabel pdiffusion 10 -3699 10 -3699 0 cellNo=1176
rlabel pdiffusion 17 -3699 17 -3699 0 cellNo=1208
rlabel pdiffusion 24 -3699 24 -3699 0 cellNo=1239
rlabel pdiffusion 31 -3699 31 -3699 0 cellNo=1253
rlabel pdiffusion 38 -3699 38 -3699 0 cellNo=1296
rlabel pdiffusion 45 -3699 45 -3699 0 cellNo=1325
rlabel pdiffusion 52 -3699 52 -3699 0 cellNo=1366
rlabel pdiffusion 59 -3699 59 -3699 0 cellNo=1404
rlabel pdiffusion 66 -3699 66 -3699 0 cellNo=1421
rlabel polysilicon 226 -8 226 -8 0 1
rlabel polysilicon 226 -14 226 -14 0 3
rlabel polysilicon 254 -8 254 -8 0 1
rlabel polysilicon 254 -14 254 -14 0 3
rlabel polysilicon 275 -8 275 -8 0 1
rlabel polysilicon 275 -14 275 -14 0 3
rlabel polysilicon 317 -8 317 -8 0 1
rlabel polysilicon 317 -14 317 -14 0 3
rlabel polysilicon 331 -8 331 -8 0 1
rlabel polysilicon 331 -14 331 -14 0 3
rlabel polysilicon 366 -8 366 -8 0 1
rlabel polysilicon 366 -14 366 -14 0 3
rlabel polysilicon 373 -8 373 -8 0 1
rlabel polysilicon 376 -14 376 -14 0 4
rlabel polysilicon 380 -8 380 -8 0 1
rlabel polysilicon 383 -14 383 -14 0 4
rlabel polysilicon 394 -14 394 -14 0 3
rlabel polysilicon 401 -8 401 -8 0 1
rlabel polysilicon 404 -8 404 -8 0 2
rlabel polysilicon 415 -8 415 -8 0 1
rlabel polysilicon 415 -14 415 -14 0 3
rlabel polysilicon 429 -8 429 -8 0 1
rlabel polysilicon 436 -8 436 -8 0 1
rlabel polysilicon 436 -14 436 -14 0 3
rlabel polysilicon 443 -14 443 -14 0 3
rlabel polysilicon 446 -14 446 -14 0 4
rlabel polysilicon 450 -8 450 -8 0 1
rlabel polysilicon 450 -14 450 -14 0 3
rlabel polysilicon 457 -8 457 -8 0 1
rlabel polysilicon 460 -8 460 -8 0 2
rlabel polysilicon 457 -14 457 -14 0 3
rlabel polysilicon 471 -8 471 -8 0 1
rlabel polysilicon 471 -14 471 -14 0 3
rlabel polysilicon 492 -8 492 -8 0 1
rlabel polysilicon 492 -14 492 -14 0 3
rlabel polysilicon 506 -8 506 -8 0 1
rlabel polysilicon 506 -14 506 -14 0 3
rlabel polysilicon 513 -8 513 -8 0 1
rlabel polysilicon 516 -8 516 -8 0 2
rlabel polysilicon 527 -8 527 -8 0 1
rlabel polysilicon 527 -14 527 -14 0 3
rlabel polysilicon 534 -8 534 -8 0 1
rlabel polysilicon 537 -8 537 -8 0 2
rlabel polysilicon 541 -14 541 -14 0 3
rlabel polysilicon 562 -8 562 -8 0 1
rlabel polysilicon 565 -14 565 -14 0 4
rlabel polysilicon 569 -8 569 -8 0 1
rlabel polysilicon 569 -14 569 -14 0 3
rlabel polysilicon 590 -8 590 -8 0 1
rlabel polysilicon 590 -14 590 -14 0 3
rlabel polysilicon 618 -14 618 -14 0 3
rlabel polysilicon 642 -8 642 -8 0 2
rlabel polysilicon 639 -14 639 -14 0 3
rlabel polysilicon 667 -8 667 -8 0 1
rlabel polysilicon 674 -8 674 -8 0 1
rlabel polysilicon 674 -14 674 -14 0 3
rlabel polysilicon 705 -8 705 -8 0 2
rlabel polysilicon 705 -14 705 -14 0 4
rlabel polysilicon 765 -8 765 -8 0 1
rlabel polysilicon 765 -14 765 -14 0 3
rlabel polysilicon 800 -8 800 -8 0 1
rlabel polysilicon 803 -8 803 -8 0 2
rlabel polysilicon 828 -8 828 -8 0 1
rlabel polysilicon 828 -14 828 -14 0 3
rlabel polysilicon 842 -8 842 -8 0 1
rlabel polysilicon 842 -14 842 -14 0 3
rlabel polysilicon 135 -37 135 -37 0 1
rlabel polysilicon 135 -43 135 -43 0 3
rlabel polysilicon 177 -43 177 -43 0 3
rlabel polysilicon 180 -43 180 -43 0 4
rlabel polysilicon 191 -37 191 -37 0 1
rlabel polysilicon 191 -43 191 -43 0 3
rlabel polysilicon 205 -37 205 -37 0 1
rlabel polysilicon 205 -43 205 -43 0 3
rlabel polysilicon 212 -37 212 -37 0 1
rlabel polysilicon 212 -43 212 -43 0 3
rlabel polysilicon 222 -37 222 -37 0 2
rlabel polysilicon 222 -43 222 -43 0 4
rlabel polysilicon 226 -37 226 -37 0 1
rlabel polysilicon 226 -43 226 -43 0 3
rlabel polysilicon 236 -43 236 -43 0 4
rlabel polysilicon 254 -37 254 -37 0 1
rlabel polysilicon 254 -43 254 -43 0 3
rlabel polysilicon 296 -37 296 -37 0 1
rlabel polysilicon 299 -37 299 -37 0 2
rlabel polysilicon 296 -43 296 -43 0 3
rlabel polysilicon 303 -37 303 -37 0 1
rlabel polysilicon 303 -43 303 -43 0 3
rlabel polysilicon 310 -37 310 -37 0 1
rlabel polysilicon 310 -43 310 -43 0 3
rlabel polysilicon 317 -37 317 -37 0 1
rlabel polysilicon 317 -43 317 -43 0 3
rlabel polysilicon 327 -37 327 -37 0 2
rlabel polysilicon 327 -43 327 -43 0 4
rlabel polysilicon 331 -37 331 -37 0 1
rlabel polysilicon 331 -43 331 -43 0 3
rlabel polysilicon 338 -37 338 -37 0 1
rlabel polysilicon 338 -43 338 -43 0 3
rlabel polysilicon 345 -37 345 -37 0 1
rlabel polysilicon 345 -43 345 -43 0 3
rlabel polysilicon 352 -37 352 -37 0 1
rlabel polysilicon 352 -43 352 -43 0 3
rlabel polysilicon 359 -37 359 -37 0 1
rlabel polysilicon 359 -43 359 -43 0 3
rlabel polysilicon 366 -37 366 -37 0 1
rlabel polysilicon 366 -43 366 -43 0 3
rlabel polysilicon 369 -43 369 -43 0 4
rlabel polysilicon 373 -37 373 -37 0 1
rlabel polysilicon 373 -43 373 -43 0 3
rlabel polysilicon 380 -37 380 -37 0 1
rlabel polysilicon 380 -43 380 -43 0 3
rlabel polysilicon 387 -37 387 -37 0 1
rlabel polysilicon 387 -43 387 -43 0 3
rlabel polysilicon 394 -37 394 -37 0 1
rlabel polysilicon 397 -43 397 -43 0 4
rlabel polysilicon 401 -37 401 -37 0 1
rlabel polysilicon 404 -37 404 -37 0 2
rlabel polysilicon 408 -37 408 -37 0 1
rlabel polysilicon 408 -43 408 -43 0 3
rlabel polysilicon 415 -37 415 -37 0 1
rlabel polysilicon 415 -43 415 -43 0 3
rlabel polysilicon 422 -37 422 -37 0 1
rlabel polysilicon 422 -43 422 -43 0 3
rlabel polysilicon 443 -37 443 -37 0 1
rlabel polysilicon 446 -37 446 -37 0 2
rlabel polysilicon 450 -37 450 -37 0 1
rlabel polysilicon 450 -43 450 -43 0 3
rlabel polysilicon 453 -43 453 -43 0 4
rlabel polysilicon 457 -37 457 -37 0 1
rlabel polysilicon 457 -43 457 -43 0 3
rlabel polysilicon 464 -37 464 -37 0 1
rlabel polysilicon 464 -43 464 -43 0 3
rlabel polysilicon 467 -43 467 -43 0 4
rlabel polysilicon 471 -37 471 -37 0 1
rlabel polysilicon 471 -43 471 -43 0 3
rlabel polysilicon 478 -37 478 -37 0 1
rlabel polysilicon 478 -43 478 -43 0 3
rlabel polysilicon 488 -37 488 -37 0 2
rlabel polysilicon 488 -43 488 -43 0 4
rlabel polysilicon 492 -37 492 -37 0 1
rlabel polysilicon 492 -43 492 -43 0 3
rlabel polysilicon 513 -37 513 -37 0 1
rlabel polysilicon 513 -43 513 -43 0 3
rlabel polysilicon 520 -37 520 -37 0 1
rlabel polysilicon 520 -43 520 -43 0 3
rlabel polysilicon 527 -37 527 -37 0 1
rlabel polysilicon 527 -43 527 -43 0 3
rlabel polysilicon 534 -37 534 -37 0 1
rlabel polysilicon 534 -43 534 -43 0 3
rlabel polysilicon 541 -37 541 -37 0 1
rlabel polysilicon 541 -43 541 -43 0 3
rlabel polysilicon 548 -37 548 -37 0 1
rlabel polysilicon 548 -43 548 -43 0 3
rlabel polysilicon 555 -37 555 -37 0 1
rlabel polysilicon 555 -43 555 -43 0 3
rlabel polysilicon 569 -37 569 -37 0 1
rlabel polysilicon 569 -43 569 -43 0 3
rlabel polysilicon 576 -37 576 -37 0 1
rlabel polysilicon 576 -43 576 -43 0 3
rlabel polysilicon 583 -37 583 -37 0 1
rlabel polysilicon 583 -43 583 -43 0 3
rlabel polysilicon 590 -43 590 -43 0 3
rlabel polysilicon 593 -43 593 -43 0 4
rlabel polysilicon 618 -37 618 -37 0 1
rlabel polysilicon 618 -43 618 -43 0 3
rlabel polysilicon 621 -43 621 -43 0 4
rlabel polysilicon 632 -37 632 -37 0 1
rlabel polysilicon 635 -37 635 -37 0 2
rlabel polysilicon 639 -37 639 -37 0 1
rlabel polysilicon 639 -43 639 -43 0 3
rlabel polysilicon 646 -37 646 -37 0 1
rlabel polysilicon 646 -43 646 -43 0 3
rlabel polysilicon 653 -37 653 -37 0 1
rlabel polysilicon 653 -43 653 -43 0 3
rlabel polysilicon 660 -37 660 -37 0 1
rlabel polysilicon 660 -43 660 -43 0 3
rlabel polysilicon 667 -37 667 -37 0 1
rlabel polysilicon 667 -43 667 -43 0 3
rlabel polysilicon 684 -37 684 -37 0 2
rlabel polysilicon 681 -43 681 -43 0 3
rlabel polysilicon 695 -37 695 -37 0 1
rlabel polysilicon 695 -43 695 -43 0 3
rlabel polysilicon 702 -37 702 -37 0 1
rlabel polysilicon 702 -43 702 -43 0 3
rlabel polysilicon 709 -37 709 -37 0 1
rlabel polysilicon 709 -43 709 -43 0 3
rlabel polysilicon 761 -37 761 -37 0 2
rlabel polysilicon 761 -43 761 -43 0 4
rlabel polysilicon 765 -37 765 -37 0 1
rlabel polysilicon 765 -43 765 -43 0 3
rlabel polysilicon 775 -37 775 -37 0 2
rlabel polysilicon 782 -37 782 -37 0 2
rlabel polysilicon 786 -37 786 -37 0 1
rlabel polysilicon 786 -43 786 -43 0 3
rlabel polysilicon 793 -37 793 -37 0 1
rlabel polysilicon 793 -43 793 -43 0 3
rlabel polysilicon 800 -37 800 -37 0 1
rlabel polysilicon 800 -43 800 -43 0 3
rlabel polysilicon 821 -37 821 -37 0 1
rlabel polysilicon 824 -43 824 -43 0 4
rlabel polysilicon 856 -37 856 -37 0 1
rlabel polysilicon 856 -43 856 -43 0 3
rlabel polysilicon 877 -37 877 -37 0 1
rlabel polysilicon 877 -43 877 -43 0 3
rlabel polysilicon 919 -37 919 -37 0 1
rlabel polysilicon 919 -43 919 -43 0 3
rlabel polysilicon 79 -86 79 -86 0 1
rlabel polysilicon 79 -92 79 -92 0 3
rlabel polysilicon 100 -86 100 -86 0 1
rlabel polysilicon 100 -92 100 -92 0 3
rlabel polysilicon 114 -92 114 -92 0 3
rlabel polysilicon 117 -92 117 -92 0 4
rlabel polysilicon 128 -86 128 -86 0 1
rlabel polysilicon 128 -92 128 -92 0 3
rlabel polysilicon 142 -86 142 -86 0 1
rlabel polysilicon 142 -92 142 -92 0 3
rlabel polysilicon 145 -92 145 -92 0 4
rlabel polysilicon 149 -86 149 -86 0 1
rlabel polysilicon 149 -92 149 -92 0 3
rlabel polysilicon 156 -86 156 -86 0 1
rlabel polysilicon 156 -92 156 -92 0 3
rlabel polysilicon 163 -86 163 -86 0 1
rlabel polysilicon 163 -92 163 -92 0 3
rlabel polysilicon 170 -86 170 -86 0 1
rlabel polysilicon 170 -92 170 -92 0 3
rlabel polysilicon 177 -86 177 -86 0 1
rlabel polysilicon 180 -86 180 -86 0 2
rlabel polysilicon 177 -92 177 -92 0 3
rlabel polysilicon 184 -86 184 -86 0 1
rlabel polysilicon 184 -92 184 -92 0 3
rlabel polysilicon 191 -86 191 -86 0 1
rlabel polysilicon 191 -92 191 -92 0 3
rlabel polysilicon 198 -86 198 -86 0 1
rlabel polysilicon 198 -92 198 -92 0 3
rlabel polysilicon 205 -86 205 -86 0 1
rlabel polysilicon 205 -92 205 -92 0 3
rlabel polysilicon 212 -92 212 -92 0 3
rlabel polysilicon 215 -92 215 -92 0 4
rlabel polysilicon 219 -86 219 -86 0 1
rlabel polysilicon 219 -92 219 -92 0 3
rlabel polysilicon 226 -86 226 -86 0 1
rlabel polysilicon 229 -86 229 -86 0 2
rlabel polysilicon 226 -92 226 -92 0 3
rlabel polysilicon 236 -86 236 -86 0 2
rlabel polysilicon 236 -92 236 -92 0 4
rlabel polysilicon 243 -86 243 -86 0 2
rlabel polysilicon 240 -92 240 -92 0 3
rlabel polysilicon 254 -86 254 -86 0 1
rlabel polysilicon 254 -92 254 -92 0 3
rlabel polysilicon 261 -86 261 -86 0 1
rlabel polysilicon 261 -92 261 -92 0 3
rlabel polysilicon 268 -86 268 -86 0 1
rlabel polysilicon 268 -92 268 -92 0 3
rlabel polysilicon 278 -86 278 -86 0 2
rlabel polysilicon 275 -92 275 -92 0 3
rlabel polysilicon 278 -92 278 -92 0 4
rlabel polysilicon 282 -92 282 -92 0 3
rlabel polysilicon 285 -92 285 -92 0 4
rlabel polysilicon 289 -86 289 -86 0 1
rlabel polysilicon 289 -92 289 -92 0 3
rlabel polysilicon 296 -86 296 -86 0 1
rlabel polysilicon 296 -92 296 -92 0 3
rlabel polysilicon 299 -92 299 -92 0 4
rlabel polysilicon 303 -86 303 -86 0 1
rlabel polysilicon 303 -92 303 -92 0 3
rlabel polysilicon 310 -86 310 -86 0 1
rlabel polysilicon 310 -92 310 -92 0 3
rlabel polysilicon 317 -86 317 -86 0 1
rlabel polysilicon 317 -92 317 -92 0 3
rlabel polysilicon 324 -86 324 -86 0 1
rlabel polysilicon 324 -92 324 -92 0 3
rlabel polysilicon 331 -86 331 -86 0 1
rlabel polysilicon 334 -92 334 -92 0 4
rlabel polysilicon 338 -86 338 -86 0 1
rlabel polysilicon 338 -92 338 -92 0 3
rlabel polysilicon 345 -86 345 -86 0 1
rlabel polysilicon 345 -92 345 -92 0 3
rlabel polysilicon 352 -86 352 -86 0 1
rlabel polysilicon 352 -92 352 -92 0 3
rlabel polysilicon 359 -86 359 -86 0 1
rlabel polysilicon 359 -92 359 -92 0 3
rlabel polysilicon 366 -86 366 -86 0 1
rlabel polysilicon 369 -86 369 -86 0 2
rlabel polysilicon 366 -92 366 -92 0 3
rlabel polysilicon 373 -86 373 -86 0 1
rlabel polysilicon 373 -92 373 -92 0 3
rlabel polysilicon 380 -86 380 -86 0 1
rlabel polysilicon 401 -86 401 -86 0 1
rlabel polysilicon 401 -92 401 -92 0 3
rlabel polysilicon 408 -86 408 -86 0 1
rlabel polysilicon 408 -92 408 -92 0 3
rlabel polysilicon 415 -86 415 -86 0 1
rlabel polysilicon 415 -92 415 -92 0 3
rlabel polysilicon 422 -86 422 -86 0 1
rlabel polysilicon 422 -92 422 -92 0 3
rlabel polysilicon 429 -86 429 -86 0 1
rlabel polysilicon 429 -92 429 -92 0 3
rlabel polysilicon 436 -86 436 -86 0 1
rlabel polysilicon 436 -92 436 -92 0 3
rlabel polysilicon 446 -86 446 -86 0 2
rlabel polysilicon 443 -92 443 -92 0 3
rlabel polysilicon 446 -92 446 -92 0 4
rlabel polysilicon 450 -86 450 -86 0 1
rlabel polysilicon 450 -92 450 -92 0 3
rlabel polysilicon 453 -92 453 -92 0 4
rlabel polysilicon 457 -86 457 -86 0 1
rlabel polysilicon 457 -92 457 -92 0 3
rlabel polysilicon 464 -86 464 -86 0 1
rlabel polysilicon 464 -92 464 -92 0 3
rlabel polysilicon 474 -86 474 -86 0 2
rlabel polysilicon 471 -92 471 -92 0 3
rlabel polysilicon 478 -86 478 -86 0 1
rlabel polysilicon 478 -92 478 -92 0 3
rlabel polysilicon 485 -86 485 -86 0 1
rlabel polysilicon 485 -92 485 -92 0 3
rlabel polysilicon 492 -86 492 -86 0 1
rlabel polysilicon 492 -92 492 -92 0 3
rlabel polysilicon 499 -86 499 -86 0 1
rlabel polysilicon 499 -92 499 -92 0 3
rlabel polysilicon 506 -86 506 -86 0 1
rlabel polysilicon 506 -92 506 -92 0 3
rlabel polysilicon 513 -86 513 -86 0 1
rlabel polysilicon 513 -92 513 -92 0 3
rlabel polysilicon 520 -86 520 -86 0 1
rlabel polysilicon 520 -92 520 -92 0 3
rlabel polysilicon 527 -86 527 -86 0 1
rlabel polysilicon 527 -92 527 -92 0 3
rlabel polysilicon 534 -86 534 -86 0 1
rlabel polysilicon 534 -92 534 -92 0 3
rlabel polysilicon 541 -86 541 -86 0 1
rlabel polysilicon 541 -92 541 -92 0 3
rlabel polysilicon 548 -86 548 -86 0 1
rlabel polysilicon 548 -92 548 -92 0 3
rlabel polysilicon 555 -86 555 -86 0 1
rlabel polysilicon 555 -92 555 -92 0 3
rlabel polysilicon 562 -86 562 -86 0 1
rlabel polysilicon 562 -92 562 -92 0 3
rlabel polysilicon 569 -86 569 -86 0 1
rlabel polysilicon 572 -86 572 -86 0 2
rlabel polysilicon 569 -92 569 -92 0 3
rlabel polysilicon 576 -86 576 -86 0 1
rlabel polysilicon 576 -92 576 -92 0 3
rlabel polysilicon 583 -86 583 -86 0 1
rlabel polysilicon 583 -92 583 -92 0 3
rlabel polysilicon 593 -86 593 -86 0 2
rlabel polysilicon 590 -92 590 -92 0 3
rlabel polysilicon 597 -86 597 -86 0 1
rlabel polysilicon 597 -92 597 -92 0 3
rlabel polysilicon 604 -86 604 -86 0 1
rlabel polysilicon 604 -92 604 -92 0 3
rlabel polysilicon 611 -86 611 -86 0 1
rlabel polysilicon 611 -92 611 -92 0 3
rlabel polysilicon 618 -86 618 -86 0 1
rlabel polysilicon 618 -92 618 -92 0 3
rlabel polysilicon 625 -86 625 -86 0 1
rlabel polysilicon 628 -86 628 -86 0 2
rlabel polysilicon 632 -86 632 -86 0 1
rlabel polysilicon 632 -92 632 -92 0 3
rlabel polysilicon 642 -86 642 -86 0 2
rlabel polysilicon 642 -92 642 -92 0 4
rlabel polysilicon 646 -86 646 -86 0 1
rlabel polysilicon 646 -92 646 -92 0 3
rlabel polysilicon 649 -92 649 -92 0 4
rlabel polysilicon 653 -86 653 -86 0 1
rlabel polysilicon 653 -92 653 -92 0 3
rlabel polysilicon 660 -86 660 -86 0 1
rlabel polysilicon 660 -92 660 -92 0 3
rlabel polysilicon 667 -86 667 -86 0 1
rlabel polysilicon 667 -92 667 -92 0 3
rlabel polysilicon 674 -86 674 -86 0 1
rlabel polysilicon 674 -92 674 -92 0 3
rlabel polysilicon 681 -86 681 -86 0 1
rlabel polysilicon 681 -92 681 -92 0 3
rlabel polysilicon 688 -86 688 -86 0 1
rlabel polysilicon 688 -92 688 -92 0 3
rlabel polysilicon 695 -86 695 -86 0 1
rlabel polysilicon 695 -92 695 -92 0 3
rlabel polysilicon 702 -86 702 -86 0 1
rlabel polysilicon 702 -92 702 -92 0 3
rlabel polysilicon 709 -86 709 -86 0 1
rlabel polysilicon 709 -92 709 -92 0 3
rlabel polysilicon 716 -86 716 -86 0 1
rlabel polysilicon 716 -92 716 -92 0 3
rlabel polysilicon 723 -86 723 -86 0 1
rlabel polysilicon 723 -92 723 -92 0 3
rlabel polysilicon 733 -86 733 -86 0 2
rlabel polysilicon 730 -92 730 -92 0 3
rlabel polysilicon 740 -86 740 -86 0 2
rlabel polysilicon 740 -92 740 -92 0 4
rlabel polysilicon 744 -86 744 -86 0 1
rlabel polysilicon 744 -92 744 -92 0 3
rlabel polysilicon 751 -86 751 -86 0 1
rlabel polysilicon 751 -92 751 -92 0 3
rlabel polysilicon 758 -86 758 -86 0 1
rlabel polysilicon 761 -92 761 -92 0 4
rlabel polysilicon 765 -86 765 -86 0 1
rlabel polysilicon 765 -92 765 -92 0 3
rlabel polysilicon 772 -86 772 -86 0 1
rlabel polysilicon 772 -92 772 -92 0 3
rlabel polysilicon 779 -86 779 -86 0 1
rlabel polysilicon 782 -86 782 -86 0 2
rlabel polysilicon 786 -86 786 -86 0 1
rlabel polysilicon 786 -92 786 -92 0 3
rlabel polysilicon 793 -86 793 -86 0 1
rlabel polysilicon 793 -92 793 -92 0 3
rlabel polysilicon 800 -86 800 -86 0 1
rlabel polysilicon 800 -92 800 -92 0 3
rlabel polysilicon 807 -86 807 -86 0 1
rlabel polysilicon 807 -92 807 -92 0 3
rlabel polysilicon 814 -86 814 -86 0 1
rlabel polysilicon 814 -92 814 -92 0 3
rlabel polysilicon 821 -86 821 -86 0 1
rlabel polysilicon 821 -92 821 -92 0 3
rlabel polysilicon 856 -86 856 -86 0 1
rlabel polysilicon 856 -92 856 -92 0 3
rlabel polysilicon 863 -86 863 -86 0 1
rlabel polysilicon 863 -92 863 -92 0 3
rlabel polysilicon 870 -86 870 -86 0 1
rlabel polysilicon 870 -92 870 -92 0 3
rlabel polysilicon 891 -86 891 -86 0 1
rlabel polysilicon 891 -92 891 -92 0 3
rlabel polysilicon 905 -86 905 -86 0 1
rlabel polysilicon 905 -92 905 -92 0 3
rlabel polysilicon 968 -86 968 -86 0 1
rlabel polysilicon 968 -92 968 -92 0 3
rlabel polysilicon 100 -157 100 -157 0 1
rlabel polysilicon 100 -163 100 -163 0 3
rlabel polysilicon 114 -157 114 -157 0 1
rlabel polysilicon 114 -163 114 -163 0 3
rlabel polysilicon 149 -157 149 -157 0 1
rlabel polysilicon 149 -163 149 -163 0 3
rlabel polysilicon 156 -163 156 -163 0 3
rlabel polysilicon 163 -157 163 -157 0 1
rlabel polysilicon 163 -163 163 -163 0 3
rlabel polysilicon 170 -157 170 -157 0 1
rlabel polysilicon 170 -163 170 -163 0 3
rlabel polysilicon 177 -157 177 -157 0 1
rlabel polysilicon 177 -163 177 -163 0 3
rlabel polysilicon 184 -157 184 -157 0 1
rlabel polysilicon 184 -163 184 -163 0 3
rlabel polysilicon 191 -157 191 -157 0 1
rlabel polysilicon 191 -163 191 -163 0 3
rlabel polysilicon 198 -157 198 -157 0 1
rlabel polysilicon 198 -163 198 -163 0 3
rlabel polysilicon 205 -157 205 -157 0 1
rlabel polysilicon 205 -163 205 -163 0 3
rlabel polysilicon 212 -157 212 -157 0 1
rlabel polysilicon 212 -163 212 -163 0 3
rlabel polysilicon 219 -157 219 -157 0 1
rlabel polysilicon 219 -163 219 -163 0 3
rlabel polysilicon 226 -157 226 -157 0 1
rlabel polysilicon 226 -163 226 -163 0 3
rlabel polysilicon 233 -157 233 -157 0 1
rlabel polysilicon 233 -163 233 -163 0 3
rlabel polysilicon 240 -157 240 -157 0 1
rlabel polysilicon 240 -163 240 -163 0 3
rlabel polysilicon 250 -157 250 -157 0 2
rlabel polysilicon 247 -163 247 -163 0 3
rlabel polysilicon 250 -163 250 -163 0 4
rlabel polysilicon 254 -157 254 -157 0 1
rlabel polysilicon 257 -163 257 -163 0 4
rlabel polysilicon 261 -157 261 -157 0 1
rlabel polysilicon 261 -163 261 -163 0 3
rlabel polysilicon 268 -157 268 -157 0 1
rlabel polysilicon 271 -157 271 -157 0 2
rlabel polysilicon 271 -163 271 -163 0 4
rlabel polysilicon 275 -157 275 -157 0 1
rlabel polysilicon 275 -163 275 -163 0 3
rlabel polysilicon 278 -163 278 -163 0 4
rlabel polysilicon 282 -157 282 -157 0 1
rlabel polysilicon 285 -157 285 -157 0 2
rlabel polysilicon 282 -163 282 -163 0 3
rlabel polysilicon 289 -157 289 -157 0 1
rlabel polysilicon 292 -157 292 -157 0 2
rlabel polysilicon 289 -163 289 -163 0 3
rlabel polysilicon 292 -163 292 -163 0 4
rlabel polysilicon 296 -157 296 -157 0 1
rlabel polysilicon 299 -157 299 -157 0 2
rlabel polysilicon 296 -163 296 -163 0 3
rlabel polysilicon 303 -157 303 -157 0 1
rlabel polysilicon 303 -163 303 -163 0 3
rlabel polysilicon 310 -157 310 -157 0 1
rlabel polysilicon 310 -163 310 -163 0 3
rlabel polysilicon 317 -157 317 -157 0 1
rlabel polysilicon 317 -163 317 -163 0 3
rlabel polysilicon 324 -157 324 -157 0 1
rlabel polysilicon 324 -163 324 -163 0 3
rlabel polysilicon 331 -157 331 -157 0 1
rlabel polysilicon 331 -163 331 -163 0 3
rlabel polysilicon 338 -157 338 -157 0 1
rlabel polysilicon 338 -163 338 -163 0 3
rlabel polysilicon 345 -157 345 -157 0 1
rlabel polysilicon 345 -163 345 -163 0 3
rlabel polysilicon 352 -157 352 -157 0 1
rlabel polysilicon 352 -163 352 -163 0 3
rlabel polysilicon 359 -157 359 -157 0 1
rlabel polysilicon 359 -163 359 -163 0 3
rlabel polysilicon 366 -157 366 -157 0 1
rlabel polysilicon 366 -163 366 -163 0 3
rlabel polysilicon 373 -157 373 -157 0 1
rlabel polysilicon 373 -163 373 -163 0 3
rlabel polysilicon 380 -163 380 -163 0 3
rlabel polysilicon 390 -157 390 -157 0 2
rlabel polysilicon 387 -163 387 -163 0 3
rlabel polysilicon 390 -163 390 -163 0 4
rlabel polysilicon 394 -157 394 -157 0 1
rlabel polysilicon 394 -163 394 -163 0 3
rlabel polysilicon 401 -157 401 -157 0 1
rlabel polysilicon 401 -163 401 -163 0 3
rlabel polysilicon 408 -157 408 -157 0 1
rlabel polysilicon 408 -163 408 -163 0 3
rlabel polysilicon 415 -157 415 -157 0 1
rlabel polysilicon 418 -157 418 -157 0 2
rlabel polysilicon 418 -163 418 -163 0 4
rlabel polysilicon 422 -157 422 -157 0 1
rlabel polysilicon 422 -163 422 -163 0 3
rlabel polysilicon 429 -157 429 -157 0 1
rlabel polysilicon 432 -157 432 -157 0 2
rlabel polysilicon 429 -163 429 -163 0 3
rlabel polysilicon 432 -163 432 -163 0 4
rlabel polysilicon 436 -157 436 -157 0 1
rlabel polysilicon 436 -163 436 -163 0 3
rlabel polysilicon 443 -157 443 -157 0 1
rlabel polysilicon 443 -163 443 -163 0 3
rlabel polysilicon 450 -157 450 -157 0 1
rlabel polysilicon 450 -163 450 -163 0 3
rlabel polysilicon 457 -157 457 -157 0 1
rlabel polysilicon 457 -163 457 -163 0 3
rlabel polysilicon 464 -157 464 -157 0 1
rlabel polysilicon 467 -157 467 -157 0 2
rlabel polysilicon 464 -163 464 -163 0 3
rlabel polysilicon 467 -163 467 -163 0 4
rlabel polysilicon 471 -157 471 -157 0 1
rlabel polysilicon 474 -157 474 -157 0 2
rlabel polysilicon 474 -163 474 -163 0 4
rlabel polysilicon 478 -157 478 -157 0 1
rlabel polysilicon 478 -163 478 -163 0 3
rlabel polysilicon 488 -157 488 -157 0 2
rlabel polysilicon 485 -163 485 -163 0 3
rlabel polysilicon 488 -163 488 -163 0 4
rlabel polysilicon 492 -157 492 -157 0 1
rlabel polysilicon 492 -163 492 -163 0 3
rlabel polysilicon 499 -157 499 -157 0 1
rlabel polysilicon 499 -163 499 -163 0 3
rlabel polysilicon 506 -157 506 -157 0 1
rlabel polysilicon 509 -157 509 -157 0 2
rlabel polysilicon 506 -163 506 -163 0 3
rlabel polysilicon 509 -163 509 -163 0 4
rlabel polysilicon 513 -157 513 -157 0 1
rlabel polysilicon 513 -163 513 -163 0 3
rlabel polysilicon 520 -157 520 -157 0 1
rlabel polysilicon 520 -163 520 -163 0 3
rlabel polysilicon 527 -157 527 -157 0 1
rlabel polysilicon 527 -163 527 -163 0 3
rlabel polysilicon 534 -157 534 -157 0 1
rlabel polysilicon 534 -163 534 -163 0 3
rlabel polysilicon 541 -157 541 -157 0 1
rlabel polysilicon 541 -163 541 -163 0 3
rlabel polysilicon 548 -157 548 -157 0 1
rlabel polysilicon 548 -163 548 -163 0 3
rlabel polysilicon 558 -157 558 -157 0 2
rlabel polysilicon 558 -163 558 -163 0 4
rlabel polysilicon 562 -157 562 -157 0 1
rlabel polysilicon 562 -163 562 -163 0 3
rlabel polysilicon 569 -157 569 -157 0 1
rlabel polysilicon 569 -163 569 -163 0 3
rlabel polysilicon 576 -157 576 -157 0 1
rlabel polysilicon 576 -163 576 -163 0 3
rlabel polysilicon 583 -157 583 -157 0 1
rlabel polysilicon 583 -163 583 -163 0 3
rlabel polysilicon 590 -157 590 -157 0 1
rlabel polysilicon 590 -163 590 -163 0 3
rlabel polysilicon 597 -157 597 -157 0 1
rlabel polysilicon 597 -163 597 -163 0 3
rlabel polysilicon 604 -157 604 -157 0 1
rlabel polysilicon 604 -163 604 -163 0 3
rlabel polysilicon 611 -157 611 -157 0 1
rlabel polysilicon 611 -163 611 -163 0 3
rlabel polysilicon 618 -157 618 -157 0 1
rlabel polysilicon 618 -163 618 -163 0 3
rlabel polysilicon 621 -163 621 -163 0 4
rlabel polysilicon 625 -157 625 -157 0 1
rlabel polysilicon 625 -163 625 -163 0 3
rlabel polysilicon 632 -157 632 -157 0 1
rlabel polysilicon 632 -163 632 -163 0 3
rlabel polysilicon 639 -157 639 -157 0 1
rlabel polysilicon 639 -163 639 -163 0 3
rlabel polysilicon 646 -157 646 -157 0 1
rlabel polysilicon 649 -157 649 -157 0 2
rlabel polysilicon 646 -163 646 -163 0 3
rlabel polysilicon 653 -157 653 -157 0 1
rlabel polysilicon 653 -163 653 -163 0 3
rlabel polysilicon 660 -157 660 -157 0 1
rlabel polysilicon 660 -163 660 -163 0 3
rlabel polysilicon 667 -157 667 -157 0 1
rlabel polysilicon 667 -163 667 -163 0 3
rlabel polysilicon 674 -157 674 -157 0 1
rlabel polysilicon 674 -163 674 -163 0 3
rlabel polysilicon 681 -157 681 -157 0 1
rlabel polysilicon 684 -157 684 -157 0 2
rlabel polysilicon 681 -163 681 -163 0 3
rlabel polysilicon 688 -157 688 -157 0 1
rlabel polysilicon 695 -163 695 -163 0 3
rlabel polysilicon 698 -163 698 -163 0 4
rlabel polysilicon 702 -157 702 -157 0 1
rlabel polysilicon 702 -163 702 -163 0 3
rlabel polysilicon 705 -163 705 -163 0 4
rlabel polysilicon 709 -157 709 -157 0 1
rlabel polysilicon 709 -163 709 -163 0 3
rlabel polysilicon 712 -163 712 -163 0 4
rlabel polysilicon 716 -157 716 -157 0 1
rlabel polysilicon 716 -163 716 -163 0 3
rlabel polysilicon 723 -157 723 -157 0 1
rlabel polysilicon 723 -163 723 -163 0 3
rlabel polysilicon 730 -157 730 -157 0 1
rlabel polysilicon 730 -163 730 -163 0 3
rlabel polysilicon 737 -157 737 -157 0 1
rlabel polysilicon 737 -163 737 -163 0 3
rlabel polysilicon 744 -157 744 -157 0 1
rlabel polysilicon 744 -163 744 -163 0 3
rlabel polysilicon 751 -157 751 -157 0 1
rlabel polysilicon 754 -157 754 -157 0 2
rlabel polysilicon 754 -163 754 -163 0 4
rlabel polysilicon 758 -157 758 -157 0 1
rlabel polysilicon 758 -163 758 -163 0 3
rlabel polysilicon 765 -157 765 -157 0 1
rlabel polysilicon 765 -163 765 -163 0 3
rlabel polysilicon 772 -157 772 -157 0 1
rlabel polysilicon 772 -163 772 -163 0 3
rlabel polysilicon 779 -157 779 -157 0 1
rlabel polysilicon 779 -163 779 -163 0 3
rlabel polysilicon 786 -157 786 -157 0 1
rlabel polysilicon 786 -163 786 -163 0 3
rlabel polysilicon 793 -157 793 -157 0 1
rlabel polysilicon 793 -163 793 -163 0 3
rlabel polysilicon 800 -157 800 -157 0 1
rlabel polysilicon 800 -163 800 -163 0 3
rlabel polysilicon 807 -157 807 -157 0 1
rlabel polysilicon 807 -163 807 -163 0 3
rlabel polysilicon 814 -157 814 -157 0 1
rlabel polysilicon 814 -163 814 -163 0 3
rlabel polysilicon 821 -157 821 -157 0 1
rlabel polysilicon 821 -163 821 -163 0 3
rlabel polysilicon 828 -157 828 -157 0 1
rlabel polysilicon 828 -163 828 -163 0 3
rlabel polysilicon 835 -157 835 -157 0 1
rlabel polysilicon 835 -163 835 -163 0 3
rlabel polysilicon 842 -157 842 -157 0 1
rlabel polysilicon 842 -163 842 -163 0 3
rlabel polysilicon 849 -157 849 -157 0 1
rlabel polysilicon 849 -163 849 -163 0 3
rlabel polysilicon 856 -157 856 -157 0 1
rlabel polysilicon 856 -163 856 -163 0 3
rlabel polysilicon 863 -157 863 -157 0 1
rlabel polysilicon 863 -163 863 -163 0 3
rlabel polysilicon 870 -157 870 -157 0 1
rlabel polysilicon 870 -163 870 -163 0 3
rlabel polysilicon 877 -157 877 -157 0 1
rlabel polysilicon 877 -163 877 -163 0 3
rlabel polysilicon 884 -157 884 -157 0 1
rlabel polysilicon 884 -163 884 -163 0 3
rlabel polysilicon 891 -157 891 -157 0 1
rlabel polysilicon 891 -163 891 -163 0 3
rlabel polysilicon 898 -157 898 -157 0 1
rlabel polysilicon 898 -163 898 -163 0 3
rlabel polysilicon 905 -157 905 -157 0 1
rlabel polysilicon 905 -163 905 -163 0 3
rlabel polysilicon 912 -157 912 -157 0 1
rlabel polysilicon 912 -163 912 -163 0 3
rlabel polysilicon 919 -157 919 -157 0 1
rlabel polysilicon 919 -163 919 -163 0 3
rlabel polysilicon 926 -157 926 -157 0 1
rlabel polysilicon 926 -163 926 -163 0 3
rlabel polysilicon 933 -157 933 -157 0 1
rlabel polysilicon 933 -163 933 -163 0 3
rlabel polysilicon 940 -157 940 -157 0 1
rlabel polysilicon 943 -163 943 -163 0 4
rlabel polysilicon 947 -157 947 -157 0 1
rlabel polysilicon 947 -163 947 -163 0 3
rlabel polysilicon 954 -157 954 -157 0 1
rlabel polysilicon 954 -163 954 -163 0 3
rlabel polysilicon 961 -157 961 -157 0 1
rlabel polysilicon 961 -163 961 -163 0 3
rlabel polysilicon 968 -157 968 -157 0 1
rlabel polysilicon 968 -163 968 -163 0 3
rlabel polysilicon 975 -157 975 -157 0 1
rlabel polysilicon 975 -163 975 -163 0 3
rlabel polysilicon 982 -157 982 -157 0 1
rlabel polysilicon 982 -163 982 -163 0 3
rlabel polysilicon 989 -157 989 -157 0 1
rlabel polysilicon 989 -163 989 -163 0 3
rlabel polysilicon 996 -163 996 -163 0 3
rlabel polysilicon 999 -163 999 -163 0 4
rlabel polysilicon 1003 -157 1003 -157 0 1
rlabel polysilicon 1003 -163 1003 -163 0 3
rlabel polysilicon 54 -258 54 -258 0 4
rlabel polysilicon 72 -252 72 -252 0 1
rlabel polysilicon 72 -258 72 -258 0 3
rlabel polysilicon 100 -252 100 -252 0 1
rlabel polysilicon 100 -258 100 -258 0 3
rlabel polysilicon 107 -252 107 -252 0 1
rlabel polysilicon 110 -252 110 -252 0 2
rlabel polysilicon 107 -258 107 -258 0 3
rlabel polysilicon 110 -258 110 -258 0 4
rlabel polysilicon 114 -252 114 -252 0 1
rlabel polysilicon 114 -258 114 -258 0 3
rlabel polysilicon 121 -252 121 -252 0 1
rlabel polysilicon 124 -252 124 -252 0 2
rlabel polysilicon 124 -258 124 -258 0 4
rlabel polysilicon 128 -252 128 -252 0 1
rlabel polysilicon 128 -258 128 -258 0 3
rlabel polysilicon 135 -252 135 -252 0 1
rlabel polysilicon 135 -258 135 -258 0 3
rlabel polysilicon 163 -252 163 -252 0 1
rlabel polysilicon 166 -252 166 -252 0 2
rlabel polysilicon 163 -258 163 -258 0 3
rlabel polysilicon 173 -252 173 -252 0 2
rlabel polysilicon 170 -258 170 -258 0 3
rlabel polysilicon 173 -258 173 -258 0 4
rlabel polysilicon 177 -252 177 -252 0 1
rlabel polysilicon 177 -258 177 -258 0 3
rlabel polysilicon 184 -252 184 -252 0 1
rlabel polysilicon 184 -258 184 -258 0 3
rlabel polysilicon 191 -252 191 -252 0 1
rlabel polysilicon 191 -258 191 -258 0 3
rlabel polysilicon 198 -252 198 -252 0 1
rlabel polysilicon 198 -258 198 -258 0 3
rlabel polysilicon 205 -252 205 -252 0 1
rlabel polysilicon 208 -252 208 -252 0 2
rlabel polysilicon 205 -258 205 -258 0 3
rlabel polysilicon 208 -258 208 -258 0 4
rlabel polysilicon 212 -252 212 -252 0 1
rlabel polysilicon 212 -258 212 -258 0 3
rlabel polysilicon 219 -252 219 -252 0 1
rlabel polysilicon 222 -252 222 -252 0 2
rlabel polysilicon 219 -258 219 -258 0 3
rlabel polysilicon 226 -252 226 -252 0 1
rlabel polysilicon 226 -258 226 -258 0 3
rlabel polysilicon 233 -252 233 -252 0 1
rlabel polysilicon 233 -258 233 -258 0 3
rlabel polysilicon 247 -252 247 -252 0 1
rlabel polysilicon 247 -258 247 -258 0 3
rlabel polysilicon 254 -252 254 -252 0 1
rlabel polysilicon 254 -258 254 -258 0 3
rlabel polysilicon 261 -252 261 -252 0 1
rlabel polysilicon 261 -258 261 -258 0 3
rlabel polysilicon 268 -252 268 -252 0 1
rlabel polysilicon 268 -258 268 -258 0 3
rlabel polysilicon 275 -252 275 -252 0 1
rlabel polysilicon 275 -258 275 -258 0 3
rlabel polysilicon 282 -252 282 -252 0 1
rlabel polysilicon 285 -252 285 -252 0 2
rlabel polysilicon 282 -258 282 -258 0 3
rlabel polysilicon 289 -252 289 -252 0 1
rlabel polysilicon 289 -258 289 -258 0 3
rlabel polysilicon 296 -252 296 -252 0 1
rlabel polysilicon 296 -258 296 -258 0 3
rlabel polysilicon 303 -252 303 -252 0 1
rlabel polysilicon 303 -258 303 -258 0 3
rlabel polysilicon 310 -252 310 -252 0 1
rlabel polysilicon 310 -258 310 -258 0 3
rlabel polysilicon 317 -258 317 -258 0 3
rlabel polysilicon 320 -258 320 -258 0 4
rlabel polysilicon 324 -252 324 -252 0 1
rlabel polysilicon 324 -258 324 -258 0 3
rlabel polysilicon 331 -252 331 -252 0 1
rlabel polysilicon 331 -258 331 -258 0 3
rlabel polysilicon 338 -252 338 -252 0 1
rlabel polysilicon 341 -252 341 -252 0 2
rlabel polysilicon 338 -258 338 -258 0 3
rlabel polysilicon 341 -258 341 -258 0 4
rlabel polysilicon 345 -252 345 -252 0 1
rlabel polysilicon 345 -258 345 -258 0 3
rlabel polysilicon 352 -252 352 -252 0 1
rlabel polysilicon 352 -258 352 -258 0 3
rlabel polysilicon 359 -252 359 -252 0 1
rlabel polysilicon 359 -258 359 -258 0 3
rlabel polysilicon 366 -252 366 -252 0 1
rlabel polysilicon 366 -258 366 -258 0 3
rlabel polysilicon 373 -252 373 -252 0 1
rlabel polysilicon 373 -258 373 -258 0 3
rlabel polysilicon 380 -252 380 -252 0 1
rlabel polysilicon 380 -258 380 -258 0 3
rlabel polysilicon 387 -252 387 -252 0 1
rlabel polysilicon 387 -258 387 -258 0 3
rlabel polysilicon 394 -252 394 -252 0 1
rlabel polysilicon 394 -258 394 -258 0 3
rlabel polysilicon 401 -252 401 -252 0 1
rlabel polysilicon 404 -252 404 -252 0 2
rlabel polysilicon 401 -258 401 -258 0 3
rlabel polysilicon 404 -258 404 -258 0 4
rlabel polysilicon 408 -252 408 -252 0 1
rlabel polysilicon 408 -258 408 -258 0 3
rlabel polysilicon 415 -252 415 -252 0 1
rlabel polysilicon 415 -258 415 -258 0 3
rlabel polysilicon 422 -252 422 -252 0 1
rlabel polysilicon 422 -258 422 -258 0 3
rlabel polysilicon 429 -252 429 -252 0 1
rlabel polysilicon 432 -252 432 -252 0 2
rlabel polysilicon 436 -252 436 -252 0 1
rlabel polysilicon 436 -258 436 -258 0 3
rlabel polysilicon 443 -252 443 -252 0 1
rlabel polysilicon 446 -252 446 -252 0 2
rlabel polysilicon 446 -258 446 -258 0 4
rlabel polysilicon 450 -252 450 -252 0 1
rlabel polysilicon 453 -252 453 -252 0 2
rlabel polysilicon 450 -258 450 -258 0 3
rlabel polysilicon 457 -252 457 -252 0 1
rlabel polysilicon 457 -258 457 -258 0 3
rlabel polysilicon 464 -252 464 -252 0 1
rlabel polysilicon 464 -258 464 -258 0 3
rlabel polysilicon 471 -252 471 -252 0 1
rlabel polysilicon 471 -258 471 -258 0 3
rlabel polysilicon 478 -252 478 -252 0 1
rlabel polysilicon 481 -252 481 -252 0 2
rlabel polysilicon 478 -258 478 -258 0 3
rlabel polysilicon 481 -258 481 -258 0 4
rlabel polysilicon 488 -252 488 -252 0 2
rlabel polysilicon 485 -258 485 -258 0 3
rlabel polysilicon 488 -258 488 -258 0 4
rlabel polysilicon 492 -252 492 -252 0 1
rlabel polysilicon 495 -252 495 -252 0 2
rlabel polysilicon 492 -258 492 -258 0 3
rlabel polysilicon 495 -258 495 -258 0 4
rlabel polysilicon 499 -252 499 -252 0 1
rlabel polysilicon 499 -258 499 -258 0 3
rlabel polysilicon 506 -252 506 -252 0 1
rlabel polysilicon 506 -258 506 -258 0 3
rlabel polysilicon 513 -252 513 -252 0 1
rlabel polysilicon 513 -258 513 -258 0 3
rlabel polysilicon 516 -258 516 -258 0 4
rlabel polysilicon 520 -252 520 -252 0 1
rlabel polysilicon 520 -258 520 -258 0 3
rlabel polysilicon 527 -252 527 -252 0 1
rlabel polysilicon 527 -258 527 -258 0 3
rlabel polysilicon 534 -252 534 -252 0 1
rlabel polysilicon 534 -258 534 -258 0 3
rlabel polysilicon 541 -252 541 -252 0 1
rlabel polysilicon 541 -258 541 -258 0 3
rlabel polysilicon 544 -258 544 -258 0 4
rlabel polysilicon 548 -252 548 -252 0 1
rlabel polysilicon 548 -258 548 -258 0 3
rlabel polysilicon 555 -252 555 -252 0 1
rlabel polysilicon 555 -258 555 -258 0 3
rlabel polysilicon 562 -252 562 -252 0 1
rlabel polysilicon 562 -258 562 -258 0 3
rlabel polysilicon 569 -252 569 -252 0 1
rlabel polysilicon 569 -258 569 -258 0 3
rlabel polysilicon 576 -252 576 -252 0 1
rlabel polysilicon 576 -258 576 -258 0 3
rlabel polysilicon 583 -252 583 -252 0 1
rlabel polysilicon 583 -258 583 -258 0 3
rlabel polysilicon 586 -258 586 -258 0 4
rlabel polysilicon 590 -252 590 -252 0 1
rlabel polysilicon 590 -258 590 -258 0 3
rlabel polysilicon 597 -252 597 -252 0 1
rlabel polysilicon 597 -258 597 -258 0 3
rlabel polysilicon 604 -252 604 -252 0 1
rlabel polysilicon 604 -258 604 -258 0 3
rlabel polysilicon 611 -252 611 -252 0 1
rlabel polysilicon 611 -258 611 -258 0 3
rlabel polysilicon 614 -258 614 -258 0 4
rlabel polysilicon 618 -252 618 -252 0 1
rlabel polysilicon 618 -258 618 -258 0 3
rlabel polysilicon 625 -252 625 -252 0 1
rlabel polysilicon 625 -258 625 -258 0 3
rlabel polysilicon 632 -252 632 -252 0 1
rlabel polysilicon 632 -258 632 -258 0 3
rlabel polysilicon 639 -252 639 -252 0 1
rlabel polysilicon 639 -258 639 -258 0 3
rlabel polysilicon 646 -252 646 -252 0 1
rlabel polysilicon 646 -258 646 -258 0 3
rlabel polysilicon 653 -252 653 -252 0 1
rlabel polysilicon 653 -258 653 -258 0 3
rlabel polysilicon 660 -252 660 -252 0 1
rlabel polysilicon 660 -258 660 -258 0 3
rlabel polysilicon 667 -252 667 -252 0 1
rlabel polysilicon 667 -258 667 -258 0 3
rlabel polysilicon 674 -252 674 -252 0 1
rlabel polysilicon 674 -258 674 -258 0 3
rlabel polysilicon 681 -252 681 -252 0 1
rlabel polysilicon 684 -252 684 -252 0 2
rlabel polysilicon 688 -258 688 -258 0 3
rlabel polysilicon 695 -252 695 -252 0 1
rlabel polysilicon 695 -258 695 -258 0 3
rlabel polysilicon 702 -252 702 -252 0 1
rlabel polysilicon 702 -258 702 -258 0 3
rlabel polysilicon 709 -252 709 -252 0 1
rlabel polysilicon 712 -252 712 -252 0 2
rlabel polysilicon 709 -258 709 -258 0 3
rlabel polysilicon 716 -252 716 -252 0 1
rlabel polysilicon 716 -258 716 -258 0 3
rlabel polysilicon 723 -252 723 -252 0 1
rlabel polysilicon 723 -258 723 -258 0 3
rlabel polysilicon 730 -252 730 -252 0 1
rlabel polysilicon 730 -258 730 -258 0 3
rlabel polysilicon 737 -252 737 -252 0 1
rlabel polysilicon 737 -258 737 -258 0 3
rlabel polysilicon 744 -252 744 -252 0 1
rlabel polysilicon 744 -258 744 -258 0 3
rlabel polysilicon 751 -252 751 -252 0 1
rlabel polysilicon 751 -258 751 -258 0 3
rlabel polysilicon 758 -252 758 -252 0 1
rlabel polysilicon 758 -258 758 -258 0 3
rlabel polysilicon 765 -252 765 -252 0 1
rlabel polysilicon 765 -258 765 -258 0 3
rlabel polysilicon 768 -258 768 -258 0 4
rlabel polysilicon 772 -252 772 -252 0 1
rlabel polysilicon 772 -258 772 -258 0 3
rlabel polysilicon 779 -252 779 -252 0 1
rlabel polysilicon 779 -258 779 -258 0 3
rlabel polysilicon 786 -252 786 -252 0 1
rlabel polysilicon 786 -258 786 -258 0 3
rlabel polysilicon 793 -252 793 -252 0 1
rlabel polysilicon 793 -258 793 -258 0 3
rlabel polysilicon 800 -252 800 -252 0 1
rlabel polysilicon 800 -258 800 -258 0 3
rlabel polysilicon 807 -252 807 -252 0 1
rlabel polysilicon 807 -258 807 -258 0 3
rlabel polysilicon 814 -252 814 -252 0 1
rlabel polysilicon 814 -258 814 -258 0 3
rlabel polysilicon 821 -252 821 -252 0 1
rlabel polysilicon 821 -258 821 -258 0 3
rlabel polysilicon 828 -252 828 -252 0 1
rlabel polysilicon 831 -258 831 -258 0 4
rlabel polysilicon 835 -252 835 -252 0 1
rlabel polysilicon 835 -258 835 -258 0 3
rlabel polysilicon 842 -258 842 -258 0 3
rlabel polysilicon 845 -258 845 -258 0 4
rlabel polysilicon 849 -252 849 -252 0 1
rlabel polysilicon 849 -258 849 -258 0 3
rlabel polysilicon 856 -252 856 -252 0 1
rlabel polysilicon 856 -258 856 -258 0 3
rlabel polysilicon 863 -252 863 -252 0 1
rlabel polysilicon 863 -258 863 -258 0 3
rlabel polysilicon 870 -252 870 -252 0 1
rlabel polysilicon 870 -258 870 -258 0 3
rlabel polysilicon 877 -252 877 -252 0 1
rlabel polysilicon 877 -258 877 -258 0 3
rlabel polysilicon 884 -252 884 -252 0 1
rlabel polysilicon 884 -258 884 -258 0 3
rlabel polysilicon 891 -252 891 -252 0 1
rlabel polysilicon 891 -258 891 -258 0 3
rlabel polysilicon 898 -252 898 -252 0 1
rlabel polysilicon 898 -258 898 -258 0 3
rlabel polysilicon 905 -252 905 -252 0 1
rlabel polysilicon 905 -258 905 -258 0 3
rlabel polysilicon 912 -252 912 -252 0 1
rlabel polysilicon 912 -258 912 -258 0 3
rlabel polysilicon 919 -252 919 -252 0 1
rlabel polysilicon 919 -258 919 -258 0 3
rlabel polysilicon 926 -252 926 -252 0 1
rlabel polysilicon 926 -258 926 -258 0 3
rlabel polysilicon 933 -252 933 -252 0 1
rlabel polysilicon 933 -258 933 -258 0 3
rlabel polysilicon 940 -252 940 -252 0 1
rlabel polysilicon 940 -258 940 -258 0 3
rlabel polysilicon 947 -252 947 -252 0 1
rlabel polysilicon 947 -258 947 -258 0 3
rlabel polysilicon 954 -252 954 -252 0 1
rlabel polysilicon 954 -258 954 -258 0 3
rlabel polysilicon 961 -252 961 -252 0 1
rlabel polysilicon 961 -258 961 -258 0 3
rlabel polysilicon 968 -252 968 -252 0 1
rlabel polysilicon 968 -258 968 -258 0 3
rlabel polysilicon 975 -252 975 -252 0 1
rlabel polysilicon 975 -258 975 -258 0 3
rlabel polysilicon 982 -252 982 -252 0 1
rlabel polysilicon 982 -258 982 -258 0 3
rlabel polysilicon 989 -252 989 -252 0 1
rlabel polysilicon 989 -258 989 -258 0 3
rlabel polysilicon 996 -252 996 -252 0 1
rlabel polysilicon 996 -258 996 -258 0 3
rlabel polysilicon 1003 -252 1003 -252 0 1
rlabel polysilicon 1003 -258 1003 -258 0 3
rlabel polysilicon 1010 -252 1010 -252 0 1
rlabel polysilicon 1010 -258 1010 -258 0 3
rlabel polysilicon 1017 -252 1017 -252 0 1
rlabel polysilicon 1017 -258 1017 -258 0 3
rlabel polysilicon 1024 -252 1024 -252 0 1
rlabel polysilicon 1024 -258 1024 -258 0 3
rlabel polysilicon 1031 -252 1031 -252 0 1
rlabel polysilicon 1031 -258 1031 -258 0 3
rlabel polysilicon 1038 -252 1038 -252 0 1
rlabel polysilicon 1038 -258 1038 -258 0 3
rlabel polysilicon 1045 -252 1045 -252 0 1
rlabel polysilicon 1045 -258 1045 -258 0 3
rlabel polysilicon 1052 -252 1052 -252 0 1
rlabel polysilicon 1052 -258 1052 -258 0 3
rlabel polysilicon 1059 -252 1059 -252 0 1
rlabel polysilicon 1059 -258 1059 -258 0 3
rlabel polysilicon 1066 -252 1066 -252 0 1
rlabel polysilicon 1066 -258 1066 -258 0 3
rlabel polysilicon 1073 -252 1073 -252 0 1
rlabel polysilicon 1073 -258 1073 -258 0 3
rlabel polysilicon 1080 -252 1080 -252 0 1
rlabel polysilicon 1080 -258 1080 -258 0 3
rlabel polysilicon 1087 -252 1087 -252 0 1
rlabel polysilicon 1087 -258 1087 -258 0 3
rlabel polysilicon 1094 -252 1094 -252 0 1
rlabel polysilicon 1094 -258 1094 -258 0 3
rlabel polysilicon 1101 -252 1101 -252 0 1
rlabel polysilicon 1101 -258 1101 -258 0 3
rlabel polysilicon 1108 -252 1108 -252 0 1
rlabel polysilicon 1108 -258 1108 -258 0 3
rlabel polysilicon 1115 -252 1115 -252 0 1
rlabel polysilicon 1115 -258 1115 -258 0 3
rlabel polysilicon 1122 -252 1122 -252 0 1
rlabel polysilicon 1122 -258 1122 -258 0 3
rlabel polysilicon 1129 -252 1129 -252 0 1
rlabel polysilicon 1129 -258 1129 -258 0 3
rlabel polysilicon 51 -355 51 -355 0 1
rlabel polysilicon 51 -361 51 -361 0 3
rlabel polysilicon 58 -355 58 -355 0 1
rlabel polysilicon 58 -361 58 -361 0 3
rlabel polysilicon 72 -355 72 -355 0 1
rlabel polysilicon 72 -361 72 -361 0 3
rlabel polysilicon 79 -355 79 -355 0 1
rlabel polysilicon 82 -355 82 -355 0 2
rlabel polysilicon 82 -361 82 -361 0 4
rlabel polysilicon 86 -355 86 -355 0 1
rlabel polysilicon 86 -361 86 -361 0 3
rlabel polysilicon 93 -355 93 -355 0 1
rlabel polysilicon 93 -361 93 -361 0 3
rlabel polysilicon 100 -355 100 -355 0 1
rlabel polysilicon 100 -361 100 -361 0 3
rlabel polysilicon 107 -355 107 -355 0 1
rlabel polysilicon 107 -361 107 -361 0 3
rlabel polysilicon 114 -355 114 -355 0 1
rlabel polysilicon 114 -361 114 -361 0 3
rlabel polysilicon 121 -355 121 -355 0 1
rlabel polysilicon 124 -355 124 -355 0 2
rlabel polysilicon 124 -361 124 -361 0 4
rlabel polysilicon 128 -355 128 -355 0 1
rlabel polysilicon 128 -361 128 -361 0 3
rlabel polysilicon 135 -355 135 -355 0 1
rlabel polysilicon 135 -361 135 -361 0 3
rlabel polysilicon 142 -355 142 -355 0 1
rlabel polysilicon 142 -361 142 -361 0 3
rlabel polysilicon 149 -355 149 -355 0 1
rlabel polysilicon 149 -361 149 -361 0 3
rlabel polysilicon 156 -355 156 -355 0 1
rlabel polysilicon 156 -361 156 -361 0 3
rlabel polysilicon 159 -361 159 -361 0 4
rlabel polysilicon 163 -355 163 -355 0 1
rlabel polysilicon 163 -361 163 -361 0 3
rlabel polysilicon 170 -355 170 -355 0 1
rlabel polysilicon 170 -361 170 -361 0 3
rlabel polysilicon 173 -361 173 -361 0 4
rlabel polysilicon 177 -355 177 -355 0 1
rlabel polysilicon 177 -361 177 -361 0 3
rlabel polysilicon 184 -355 184 -355 0 1
rlabel polysilicon 184 -361 184 -361 0 3
rlabel polysilicon 191 -355 191 -355 0 1
rlabel polysilicon 191 -361 191 -361 0 3
rlabel polysilicon 198 -355 198 -355 0 1
rlabel polysilicon 198 -361 198 -361 0 3
rlabel polysilicon 205 -355 205 -355 0 1
rlabel polysilicon 205 -361 205 -361 0 3
rlabel polysilicon 212 -355 212 -355 0 1
rlabel polysilicon 212 -361 212 -361 0 3
rlabel polysilicon 219 -355 219 -355 0 1
rlabel polysilicon 219 -361 219 -361 0 3
rlabel polysilicon 226 -355 226 -355 0 1
rlabel polysilicon 226 -361 226 -361 0 3
rlabel polysilicon 236 -355 236 -355 0 2
rlabel polysilicon 233 -361 233 -361 0 3
rlabel polysilicon 240 -355 240 -355 0 1
rlabel polysilicon 240 -361 240 -361 0 3
rlabel polysilicon 254 -355 254 -355 0 1
rlabel polysilicon 254 -361 254 -361 0 3
rlabel polysilicon 268 -355 268 -355 0 1
rlabel polysilicon 268 -361 268 -361 0 3
rlabel polysilicon 275 -355 275 -355 0 1
rlabel polysilicon 275 -361 275 -361 0 3
rlabel polysilicon 289 -355 289 -355 0 1
rlabel polysilicon 289 -361 289 -361 0 3
rlabel polysilicon 296 -355 296 -355 0 1
rlabel polysilicon 296 -361 296 -361 0 3
rlabel polysilicon 303 -355 303 -355 0 1
rlabel polysilicon 303 -361 303 -361 0 3
rlabel polysilicon 310 -355 310 -355 0 1
rlabel polysilicon 310 -361 310 -361 0 3
rlabel polysilicon 317 -355 317 -355 0 1
rlabel polysilicon 317 -361 317 -361 0 3
rlabel polysilicon 324 -355 324 -355 0 1
rlabel polysilicon 324 -361 324 -361 0 3
rlabel polysilicon 338 -355 338 -355 0 1
rlabel polysilicon 338 -361 338 -361 0 3
rlabel polysilicon 345 -355 345 -355 0 1
rlabel polysilicon 345 -361 345 -361 0 3
rlabel polysilicon 352 -355 352 -355 0 1
rlabel polysilicon 352 -361 352 -361 0 3
rlabel polysilicon 373 -355 373 -355 0 1
rlabel polysilicon 373 -361 373 -361 0 3
rlabel polysilicon 380 -355 380 -355 0 1
rlabel polysilicon 380 -361 380 -361 0 3
rlabel polysilicon 387 -355 387 -355 0 1
rlabel polysilicon 387 -361 387 -361 0 3
rlabel polysilicon 394 -355 394 -355 0 1
rlabel polysilicon 394 -361 394 -361 0 3
rlabel polysilicon 401 -355 401 -355 0 1
rlabel polysilicon 401 -361 401 -361 0 3
rlabel polysilicon 408 -355 408 -355 0 1
rlabel polysilicon 408 -361 408 -361 0 3
rlabel polysilicon 415 -355 415 -355 0 1
rlabel polysilicon 415 -361 415 -361 0 3
rlabel polysilicon 422 -355 422 -355 0 1
rlabel polysilicon 422 -361 422 -361 0 3
rlabel polysilicon 429 -355 429 -355 0 1
rlabel polysilicon 429 -361 429 -361 0 3
rlabel polysilicon 436 -355 436 -355 0 1
rlabel polysilicon 436 -361 436 -361 0 3
rlabel polysilicon 443 -355 443 -355 0 1
rlabel polysilicon 443 -361 443 -361 0 3
rlabel polysilicon 450 -355 450 -355 0 1
rlabel polysilicon 450 -361 450 -361 0 3
rlabel polysilicon 457 -355 457 -355 0 1
rlabel polysilicon 457 -361 457 -361 0 3
rlabel polysilicon 467 -355 467 -355 0 2
rlabel polysilicon 467 -361 467 -361 0 4
rlabel polysilicon 471 -355 471 -355 0 1
rlabel polysilicon 471 -361 471 -361 0 3
rlabel polysilicon 474 -361 474 -361 0 4
rlabel polysilicon 478 -355 478 -355 0 1
rlabel polysilicon 481 -355 481 -355 0 2
rlabel polysilicon 478 -361 478 -361 0 3
rlabel polysilicon 481 -361 481 -361 0 4
rlabel polysilicon 485 -355 485 -355 0 1
rlabel polysilicon 488 -355 488 -355 0 2
rlabel polysilicon 485 -361 485 -361 0 3
rlabel polysilicon 488 -361 488 -361 0 4
rlabel polysilicon 499 -355 499 -355 0 1
rlabel polysilicon 499 -361 499 -361 0 3
rlabel polysilicon 506 -355 506 -355 0 1
rlabel polysilicon 506 -361 506 -361 0 3
rlabel polysilicon 513 -355 513 -355 0 1
rlabel polysilicon 513 -361 513 -361 0 3
rlabel polysilicon 516 -361 516 -361 0 4
rlabel polysilicon 520 -355 520 -355 0 1
rlabel polysilicon 520 -361 520 -361 0 3
rlabel polysilicon 527 -355 527 -355 0 1
rlabel polysilicon 530 -355 530 -355 0 2
rlabel polysilicon 527 -361 527 -361 0 3
rlabel polysilicon 530 -361 530 -361 0 4
rlabel polysilicon 534 -355 534 -355 0 1
rlabel polysilicon 534 -361 534 -361 0 3
rlabel polysilicon 541 -355 541 -355 0 1
rlabel polysilicon 541 -361 541 -361 0 3
rlabel polysilicon 548 -355 548 -355 0 1
rlabel polysilicon 548 -361 548 -361 0 3
rlabel polysilicon 555 -355 555 -355 0 1
rlabel polysilicon 555 -361 555 -361 0 3
rlabel polysilicon 562 -355 562 -355 0 1
rlabel polysilicon 562 -361 562 -361 0 3
rlabel polysilicon 565 -361 565 -361 0 4
rlabel polysilicon 569 -355 569 -355 0 1
rlabel polysilicon 569 -361 569 -361 0 3
rlabel polysilicon 572 -361 572 -361 0 4
rlabel polysilicon 576 -355 576 -355 0 1
rlabel polysilicon 579 -355 579 -355 0 2
rlabel polysilicon 576 -361 576 -361 0 3
rlabel polysilicon 579 -361 579 -361 0 4
rlabel polysilicon 583 -355 583 -355 0 1
rlabel polysilicon 586 -355 586 -355 0 2
rlabel polysilicon 583 -361 583 -361 0 3
rlabel polysilicon 586 -361 586 -361 0 4
rlabel polysilicon 590 -355 590 -355 0 1
rlabel polysilicon 593 -355 593 -355 0 2
rlabel polysilicon 590 -361 590 -361 0 3
rlabel polysilicon 597 -355 597 -355 0 1
rlabel polysilicon 597 -361 597 -361 0 3
rlabel polysilicon 604 -355 604 -355 0 1
rlabel polysilicon 607 -355 607 -355 0 2
rlabel polysilicon 604 -361 604 -361 0 3
rlabel polysilicon 607 -361 607 -361 0 4
rlabel polysilicon 611 -355 611 -355 0 1
rlabel polysilicon 611 -361 611 -361 0 3
rlabel polysilicon 618 -355 618 -355 0 1
rlabel polysilicon 618 -361 618 -361 0 3
rlabel polysilicon 625 -355 625 -355 0 1
rlabel polysilicon 625 -361 625 -361 0 3
rlabel polysilicon 632 -355 632 -355 0 1
rlabel polysilicon 635 -355 635 -355 0 2
rlabel polysilicon 632 -361 632 -361 0 3
rlabel polysilicon 635 -361 635 -361 0 4
rlabel polysilicon 639 -355 639 -355 0 1
rlabel polysilicon 639 -361 639 -361 0 3
rlabel polysilicon 646 -355 646 -355 0 1
rlabel polysilicon 646 -361 646 -361 0 3
rlabel polysilicon 653 -355 653 -355 0 1
rlabel polysilicon 653 -361 653 -361 0 3
rlabel polysilicon 663 -355 663 -355 0 2
rlabel polysilicon 660 -361 660 -361 0 3
rlabel polysilicon 663 -361 663 -361 0 4
rlabel polysilicon 667 -355 667 -355 0 1
rlabel polysilicon 667 -361 667 -361 0 3
rlabel polysilicon 674 -355 674 -355 0 1
rlabel polysilicon 674 -361 674 -361 0 3
rlabel polysilicon 684 -355 684 -355 0 2
rlabel polysilicon 681 -361 681 -361 0 3
rlabel polysilicon 684 -361 684 -361 0 4
rlabel polysilicon 688 -355 688 -355 0 1
rlabel polysilicon 688 -361 688 -361 0 3
rlabel polysilicon 695 -355 695 -355 0 1
rlabel polysilicon 695 -361 695 -361 0 3
rlabel polysilicon 702 -355 702 -355 0 1
rlabel polysilicon 702 -361 702 -361 0 3
rlabel polysilicon 709 -355 709 -355 0 1
rlabel polysilicon 709 -361 709 -361 0 3
rlabel polysilicon 719 -355 719 -355 0 2
rlabel polysilicon 716 -361 716 -361 0 3
rlabel polysilicon 726 -355 726 -355 0 2
rlabel polysilicon 723 -361 723 -361 0 3
rlabel polysilicon 726 -361 726 -361 0 4
rlabel polysilicon 730 -355 730 -355 0 1
rlabel polysilicon 730 -361 730 -361 0 3
rlabel polysilicon 737 -355 737 -355 0 1
rlabel polysilicon 737 -361 737 -361 0 3
rlabel polysilicon 744 -355 744 -355 0 1
rlabel polysilicon 744 -361 744 -361 0 3
rlabel polysilicon 751 -355 751 -355 0 1
rlabel polysilicon 751 -361 751 -361 0 3
rlabel polysilicon 758 -355 758 -355 0 1
rlabel polysilicon 758 -361 758 -361 0 3
rlabel polysilicon 765 -355 765 -355 0 1
rlabel polysilicon 765 -361 765 -361 0 3
rlabel polysilicon 772 -361 772 -361 0 3
rlabel polysilicon 775 -361 775 -361 0 4
rlabel polysilicon 779 -355 779 -355 0 1
rlabel polysilicon 779 -361 779 -361 0 3
rlabel polysilicon 786 -355 786 -355 0 1
rlabel polysilicon 789 -361 789 -361 0 4
rlabel polysilicon 793 -355 793 -355 0 1
rlabel polysilicon 793 -361 793 -361 0 3
rlabel polysilicon 800 -355 800 -355 0 1
rlabel polysilicon 800 -361 800 -361 0 3
rlabel polysilicon 807 -355 807 -355 0 1
rlabel polysilicon 807 -361 807 -361 0 3
rlabel polysilicon 814 -355 814 -355 0 1
rlabel polysilicon 814 -361 814 -361 0 3
rlabel polysilicon 821 -355 821 -355 0 1
rlabel polysilicon 821 -361 821 -361 0 3
rlabel polysilicon 828 -355 828 -355 0 1
rlabel polysilicon 828 -361 828 -361 0 3
rlabel polysilicon 835 -355 835 -355 0 1
rlabel polysilicon 835 -361 835 -361 0 3
rlabel polysilicon 842 -355 842 -355 0 1
rlabel polysilicon 842 -361 842 -361 0 3
rlabel polysilicon 849 -355 849 -355 0 1
rlabel polysilicon 849 -361 849 -361 0 3
rlabel polysilicon 856 -355 856 -355 0 1
rlabel polysilicon 856 -361 856 -361 0 3
rlabel polysilicon 863 -355 863 -355 0 1
rlabel polysilicon 863 -361 863 -361 0 3
rlabel polysilicon 870 -355 870 -355 0 1
rlabel polysilicon 870 -361 870 -361 0 3
rlabel polysilicon 877 -355 877 -355 0 1
rlabel polysilicon 877 -361 877 -361 0 3
rlabel polysilicon 884 -355 884 -355 0 1
rlabel polysilicon 884 -361 884 -361 0 3
rlabel polysilicon 891 -355 891 -355 0 1
rlabel polysilicon 891 -361 891 -361 0 3
rlabel polysilicon 898 -355 898 -355 0 1
rlabel polysilicon 898 -361 898 -361 0 3
rlabel polysilicon 905 -355 905 -355 0 1
rlabel polysilicon 905 -361 905 -361 0 3
rlabel polysilicon 912 -355 912 -355 0 1
rlabel polysilicon 912 -361 912 -361 0 3
rlabel polysilicon 919 -355 919 -355 0 1
rlabel polysilicon 919 -361 919 -361 0 3
rlabel polysilicon 926 -355 926 -355 0 1
rlabel polysilicon 926 -361 926 -361 0 3
rlabel polysilicon 933 -355 933 -355 0 1
rlabel polysilicon 933 -361 933 -361 0 3
rlabel polysilicon 940 -355 940 -355 0 1
rlabel polysilicon 940 -361 940 -361 0 3
rlabel polysilicon 947 -355 947 -355 0 1
rlabel polysilicon 947 -361 947 -361 0 3
rlabel polysilicon 954 -355 954 -355 0 1
rlabel polysilicon 954 -361 954 -361 0 3
rlabel polysilicon 961 -355 961 -355 0 1
rlabel polysilicon 961 -361 961 -361 0 3
rlabel polysilicon 968 -355 968 -355 0 1
rlabel polysilicon 968 -361 968 -361 0 3
rlabel polysilicon 975 -355 975 -355 0 1
rlabel polysilicon 975 -361 975 -361 0 3
rlabel polysilicon 982 -355 982 -355 0 1
rlabel polysilicon 982 -361 982 -361 0 3
rlabel polysilicon 989 -355 989 -355 0 1
rlabel polysilicon 989 -361 989 -361 0 3
rlabel polysilicon 996 -355 996 -355 0 1
rlabel polysilicon 996 -361 996 -361 0 3
rlabel polysilicon 1003 -355 1003 -355 0 1
rlabel polysilicon 1003 -361 1003 -361 0 3
rlabel polysilicon 1010 -355 1010 -355 0 1
rlabel polysilicon 1010 -361 1010 -361 0 3
rlabel polysilicon 1017 -355 1017 -355 0 1
rlabel polysilicon 1017 -361 1017 -361 0 3
rlabel polysilicon 1024 -355 1024 -355 0 1
rlabel polysilicon 1024 -361 1024 -361 0 3
rlabel polysilicon 1031 -355 1031 -355 0 1
rlabel polysilicon 1031 -361 1031 -361 0 3
rlabel polysilicon 1038 -355 1038 -355 0 1
rlabel polysilicon 1038 -361 1038 -361 0 3
rlabel polysilicon 1045 -355 1045 -355 0 1
rlabel polysilicon 1045 -361 1045 -361 0 3
rlabel polysilicon 1052 -355 1052 -355 0 1
rlabel polysilicon 1052 -361 1052 -361 0 3
rlabel polysilicon 1059 -355 1059 -355 0 1
rlabel polysilicon 1059 -361 1059 -361 0 3
rlabel polysilicon 1066 -355 1066 -355 0 1
rlabel polysilicon 1066 -361 1066 -361 0 3
rlabel polysilicon 1073 -355 1073 -355 0 1
rlabel polysilicon 1073 -361 1073 -361 0 3
rlabel polysilicon 1080 -355 1080 -355 0 1
rlabel polysilicon 1080 -361 1080 -361 0 3
rlabel polysilicon 1087 -355 1087 -355 0 1
rlabel polysilicon 1087 -361 1087 -361 0 3
rlabel polysilicon 1094 -355 1094 -355 0 1
rlabel polysilicon 1094 -361 1094 -361 0 3
rlabel polysilicon 1101 -355 1101 -355 0 1
rlabel polysilicon 1101 -361 1101 -361 0 3
rlabel polysilicon 1108 -355 1108 -355 0 1
rlabel polysilicon 1108 -361 1108 -361 0 3
rlabel polysilicon 1115 -355 1115 -355 0 1
rlabel polysilicon 1115 -361 1115 -361 0 3
rlabel polysilicon 1122 -355 1122 -355 0 1
rlabel polysilicon 1122 -361 1122 -361 0 3
rlabel polysilicon 1129 -355 1129 -355 0 1
rlabel polysilicon 1129 -361 1129 -361 0 3
rlabel polysilicon 1136 -355 1136 -355 0 1
rlabel polysilicon 1136 -361 1136 -361 0 3
rlabel polysilicon 1143 -355 1143 -355 0 1
rlabel polysilicon 1143 -361 1143 -361 0 3
rlabel polysilicon 1150 -355 1150 -355 0 1
rlabel polysilicon 1150 -361 1150 -361 0 3
rlabel polysilicon 1157 -355 1157 -355 0 1
rlabel polysilicon 1157 -361 1157 -361 0 3
rlabel polysilicon 1164 -355 1164 -355 0 1
rlabel polysilicon 1164 -361 1164 -361 0 3
rlabel polysilicon 1171 -355 1171 -355 0 1
rlabel polysilicon 1171 -361 1171 -361 0 3
rlabel polysilicon 1178 -355 1178 -355 0 1
rlabel polysilicon 1178 -361 1178 -361 0 3
rlabel polysilicon 1185 -355 1185 -355 0 1
rlabel polysilicon 1185 -361 1185 -361 0 3
rlabel polysilicon 1192 -355 1192 -355 0 1
rlabel polysilicon 1192 -361 1192 -361 0 3
rlabel polysilicon 1199 -355 1199 -355 0 1
rlabel polysilicon 1199 -361 1199 -361 0 3
rlabel polysilicon 1206 -355 1206 -355 0 1
rlabel polysilicon 1206 -361 1206 -361 0 3
rlabel polysilicon 1213 -355 1213 -355 0 1
rlabel polysilicon 1213 -361 1213 -361 0 3
rlabel polysilicon 1220 -355 1220 -355 0 1
rlabel polysilicon 1220 -361 1220 -361 0 3
rlabel polysilicon 1227 -355 1227 -355 0 1
rlabel polysilicon 1227 -361 1227 -361 0 3
rlabel polysilicon 1234 -355 1234 -355 0 1
rlabel polysilicon 1234 -361 1234 -361 0 3
rlabel polysilicon 1241 -355 1241 -355 0 1
rlabel polysilicon 1241 -361 1241 -361 0 3
rlabel polysilicon 1248 -355 1248 -355 0 1
rlabel polysilicon 1248 -361 1248 -361 0 3
rlabel polysilicon 1255 -355 1255 -355 0 1
rlabel polysilicon 1255 -361 1255 -361 0 3
rlabel polysilicon 1262 -355 1262 -355 0 1
rlabel polysilicon 1262 -361 1262 -361 0 3
rlabel polysilicon 1269 -355 1269 -355 0 1
rlabel polysilicon 1269 -361 1269 -361 0 3
rlabel polysilicon 1276 -355 1276 -355 0 1
rlabel polysilicon 1276 -361 1276 -361 0 3
rlabel polysilicon 1283 -355 1283 -355 0 1
rlabel polysilicon 1283 -361 1283 -361 0 3
rlabel polysilicon 1290 -355 1290 -355 0 1
rlabel polysilicon 1290 -361 1290 -361 0 3
rlabel polysilicon 1300 -361 1300 -361 0 4
rlabel polysilicon 40 -486 40 -486 0 4
rlabel polysilicon 65 -480 65 -480 0 1
rlabel polysilicon 65 -486 65 -486 0 3
rlabel polysilicon 72 -480 72 -480 0 1
rlabel polysilicon 72 -486 72 -486 0 3
rlabel polysilicon 79 -480 79 -480 0 1
rlabel polysilicon 79 -486 79 -486 0 3
rlabel polysilicon 86 -480 86 -480 0 1
rlabel polysilicon 86 -486 86 -486 0 3
rlabel polysilicon 96 -480 96 -480 0 2
rlabel polysilicon 93 -486 93 -486 0 3
rlabel polysilicon 96 -486 96 -486 0 4
rlabel polysilicon 100 -480 100 -480 0 1
rlabel polysilicon 100 -486 100 -486 0 3
rlabel polysilicon 107 -480 107 -480 0 1
rlabel polysilicon 107 -486 107 -486 0 3
rlabel polysilicon 124 -480 124 -480 0 2
rlabel polysilicon 121 -486 121 -486 0 3
rlabel polysilicon 124 -486 124 -486 0 4
rlabel polysilicon 128 -480 128 -480 0 1
rlabel polysilicon 131 -480 131 -480 0 2
rlabel polysilicon 128 -486 128 -486 0 3
rlabel polysilicon 131 -486 131 -486 0 4
rlabel polysilicon 135 -480 135 -480 0 1
rlabel polysilicon 135 -486 135 -486 0 3
rlabel polysilicon 142 -480 142 -480 0 1
rlabel polysilicon 142 -486 142 -486 0 3
rlabel polysilicon 149 -480 149 -480 0 1
rlabel polysilicon 152 -480 152 -480 0 2
rlabel polysilicon 149 -486 149 -486 0 3
rlabel polysilicon 152 -486 152 -486 0 4
rlabel polysilicon 156 -480 156 -480 0 1
rlabel polysilicon 156 -486 156 -486 0 3
rlabel polysilicon 163 -480 163 -480 0 1
rlabel polysilicon 163 -486 163 -486 0 3
rlabel polysilicon 170 -480 170 -480 0 1
rlabel polysilicon 170 -486 170 -486 0 3
rlabel polysilicon 177 -480 177 -480 0 1
rlabel polysilicon 177 -486 177 -486 0 3
rlabel polysilicon 184 -480 184 -480 0 1
rlabel polysilicon 184 -486 184 -486 0 3
rlabel polysilicon 191 -480 191 -480 0 1
rlabel polysilicon 191 -486 191 -486 0 3
rlabel polysilicon 198 -480 198 -480 0 1
rlabel polysilicon 198 -486 198 -486 0 3
rlabel polysilicon 205 -480 205 -480 0 1
rlabel polysilicon 205 -486 205 -486 0 3
rlabel polysilicon 212 -480 212 -480 0 1
rlabel polysilicon 215 -480 215 -480 0 2
rlabel polysilicon 215 -486 215 -486 0 4
rlabel polysilicon 219 -480 219 -480 0 1
rlabel polysilicon 219 -486 219 -486 0 3
rlabel polysilicon 226 -480 226 -480 0 1
rlabel polysilicon 226 -486 226 -486 0 3
rlabel polysilicon 233 -480 233 -480 0 1
rlabel polysilicon 233 -486 233 -486 0 3
rlabel polysilicon 240 -480 240 -480 0 1
rlabel polysilicon 240 -486 240 -486 0 3
rlabel polysilicon 247 -480 247 -480 0 1
rlabel polysilicon 247 -486 247 -486 0 3
rlabel polysilicon 254 -480 254 -480 0 1
rlabel polysilicon 254 -486 254 -486 0 3
rlabel polysilicon 261 -480 261 -480 0 1
rlabel polysilicon 261 -486 261 -486 0 3
rlabel polysilicon 268 -480 268 -480 0 1
rlabel polysilicon 268 -486 268 -486 0 3
rlabel polysilicon 296 -480 296 -480 0 1
rlabel polysilicon 296 -486 296 -486 0 3
rlabel polysilicon 303 -480 303 -480 0 1
rlabel polysilicon 303 -486 303 -486 0 3
rlabel polysilicon 310 -480 310 -480 0 1
rlabel polysilicon 310 -486 310 -486 0 3
rlabel polysilicon 317 -480 317 -480 0 1
rlabel polysilicon 317 -486 317 -486 0 3
rlabel polysilicon 324 -480 324 -480 0 1
rlabel polysilicon 324 -486 324 -486 0 3
rlabel polysilicon 331 -480 331 -480 0 1
rlabel polysilicon 331 -486 331 -486 0 3
rlabel polysilicon 338 -480 338 -480 0 1
rlabel polysilicon 338 -486 338 -486 0 3
rlabel polysilicon 345 -480 345 -480 0 1
rlabel polysilicon 345 -486 345 -486 0 3
rlabel polysilicon 352 -480 352 -480 0 1
rlabel polysilicon 355 -480 355 -480 0 2
rlabel polysilicon 355 -486 355 -486 0 4
rlabel polysilicon 359 -480 359 -480 0 1
rlabel polysilicon 359 -486 359 -486 0 3
rlabel polysilicon 366 -480 366 -480 0 1
rlabel polysilicon 366 -486 366 -486 0 3
rlabel polysilicon 373 -480 373 -480 0 1
rlabel polysilicon 373 -486 373 -486 0 3
rlabel polysilicon 380 -480 380 -480 0 1
rlabel polysilicon 380 -486 380 -486 0 3
rlabel polysilicon 387 -480 387 -480 0 1
rlabel polysilicon 387 -486 387 -486 0 3
rlabel polysilicon 394 -480 394 -480 0 1
rlabel polysilicon 394 -486 394 -486 0 3
rlabel polysilicon 401 -480 401 -480 0 1
rlabel polysilicon 401 -486 401 -486 0 3
rlabel polysilicon 408 -480 408 -480 0 1
rlabel polysilicon 408 -486 408 -486 0 3
rlabel polysilicon 415 -480 415 -480 0 1
rlabel polysilicon 415 -486 415 -486 0 3
rlabel polysilicon 422 -480 422 -480 0 1
rlabel polysilicon 422 -486 422 -486 0 3
rlabel polysilicon 429 -480 429 -480 0 1
rlabel polysilicon 429 -486 429 -486 0 3
rlabel polysilicon 436 -480 436 -480 0 1
rlabel polysilicon 436 -486 436 -486 0 3
rlabel polysilicon 443 -480 443 -480 0 1
rlabel polysilicon 443 -486 443 -486 0 3
rlabel polysilicon 450 -480 450 -480 0 1
rlabel polysilicon 450 -486 450 -486 0 3
rlabel polysilicon 457 -480 457 -480 0 1
rlabel polysilicon 460 -480 460 -480 0 2
rlabel polysilicon 457 -486 457 -486 0 3
rlabel polysilicon 460 -486 460 -486 0 4
rlabel polysilicon 464 -480 464 -480 0 1
rlabel polysilicon 464 -486 464 -486 0 3
rlabel polysilicon 471 -480 471 -480 0 1
rlabel polysilicon 471 -486 471 -486 0 3
rlabel polysilicon 478 -480 478 -480 0 1
rlabel polysilicon 478 -486 478 -486 0 3
rlabel polysilicon 485 -480 485 -480 0 1
rlabel polysilicon 485 -486 485 -486 0 3
rlabel polysilicon 492 -480 492 -480 0 1
rlabel polysilicon 492 -486 492 -486 0 3
rlabel polysilicon 499 -480 499 -480 0 1
rlabel polysilicon 502 -480 502 -480 0 2
rlabel polysilicon 499 -486 499 -486 0 3
rlabel polysilicon 502 -486 502 -486 0 4
rlabel polysilicon 506 -480 506 -480 0 1
rlabel polysilicon 506 -486 506 -486 0 3
rlabel polysilicon 513 -480 513 -480 0 1
rlabel polysilicon 516 -480 516 -480 0 2
rlabel polysilicon 513 -486 513 -486 0 3
rlabel polysilicon 520 -480 520 -480 0 1
rlabel polysilicon 520 -486 520 -486 0 3
rlabel polysilicon 527 -480 527 -480 0 1
rlabel polysilicon 527 -486 527 -486 0 3
rlabel polysilicon 534 -480 534 -480 0 1
rlabel polysilicon 537 -480 537 -480 0 2
rlabel polysilicon 534 -486 534 -486 0 3
rlabel polysilicon 537 -486 537 -486 0 4
rlabel polysilicon 541 -480 541 -480 0 1
rlabel polysilicon 541 -486 541 -486 0 3
rlabel polysilicon 548 -480 548 -480 0 1
rlabel polysilicon 548 -486 548 -486 0 3
rlabel polysilicon 555 -480 555 -480 0 1
rlabel polysilicon 558 -480 558 -480 0 2
rlabel polysilicon 555 -486 555 -486 0 3
rlabel polysilicon 562 -480 562 -480 0 1
rlabel polysilicon 562 -486 562 -486 0 3
rlabel polysilicon 569 -480 569 -480 0 1
rlabel polysilicon 569 -486 569 -486 0 3
rlabel polysilicon 576 -480 576 -480 0 1
rlabel polysilicon 579 -480 579 -480 0 2
rlabel polysilicon 579 -486 579 -486 0 4
rlabel polysilicon 583 -480 583 -480 0 1
rlabel polysilicon 583 -486 583 -486 0 3
rlabel polysilicon 590 -480 590 -480 0 1
rlabel polysilicon 590 -486 590 -486 0 3
rlabel polysilicon 597 -480 597 -480 0 1
rlabel polysilicon 597 -486 597 -486 0 3
rlabel polysilicon 600 -486 600 -486 0 4
rlabel polysilicon 604 -480 604 -480 0 1
rlabel polysilicon 604 -486 604 -486 0 3
rlabel polysilicon 611 -480 611 -480 0 1
rlabel polysilicon 614 -480 614 -480 0 2
rlabel polysilicon 611 -486 611 -486 0 3
rlabel polysilicon 614 -486 614 -486 0 4
rlabel polysilicon 618 -480 618 -480 0 1
rlabel polysilicon 618 -486 618 -486 0 3
rlabel polysilicon 625 -480 625 -480 0 1
rlabel polysilicon 625 -486 625 -486 0 3
rlabel polysilicon 632 -480 632 -480 0 1
rlabel polysilicon 635 -480 635 -480 0 2
rlabel polysilicon 632 -486 632 -486 0 3
rlabel polysilicon 635 -486 635 -486 0 4
rlabel polysilicon 639 -480 639 -480 0 1
rlabel polysilicon 642 -480 642 -480 0 2
rlabel polysilicon 639 -486 639 -486 0 3
rlabel polysilicon 646 -480 646 -480 0 1
rlabel polysilicon 646 -486 646 -486 0 3
rlabel polysilicon 653 -480 653 -480 0 1
rlabel polysilicon 653 -486 653 -486 0 3
rlabel polysilicon 660 -480 660 -480 0 1
rlabel polysilicon 660 -486 660 -486 0 3
rlabel polysilicon 667 -480 667 -480 0 1
rlabel polysilicon 667 -486 667 -486 0 3
rlabel polysilicon 674 -480 674 -480 0 1
rlabel polysilicon 677 -480 677 -480 0 2
rlabel polysilicon 674 -486 674 -486 0 3
rlabel polysilicon 684 -480 684 -480 0 2
rlabel polysilicon 684 -486 684 -486 0 4
rlabel polysilicon 688 -480 688 -480 0 1
rlabel polysilicon 688 -486 688 -486 0 3
rlabel polysilicon 695 -480 695 -480 0 1
rlabel polysilicon 695 -486 695 -486 0 3
rlabel polysilicon 702 -480 702 -480 0 1
rlabel polysilicon 702 -486 702 -486 0 3
rlabel polysilicon 709 -480 709 -480 0 1
rlabel polysilicon 709 -486 709 -486 0 3
rlabel polysilicon 716 -480 716 -480 0 1
rlabel polysilicon 719 -480 719 -480 0 2
rlabel polysilicon 716 -486 716 -486 0 3
rlabel polysilicon 719 -486 719 -486 0 4
rlabel polysilicon 723 -480 723 -480 0 1
rlabel polysilicon 723 -486 723 -486 0 3
rlabel polysilicon 730 -480 730 -480 0 1
rlabel polysilicon 730 -486 730 -486 0 3
rlabel polysilicon 737 -480 737 -480 0 1
rlabel polysilicon 737 -486 737 -486 0 3
rlabel polysilicon 744 -480 744 -480 0 1
rlabel polysilicon 744 -486 744 -486 0 3
rlabel polysilicon 754 -480 754 -480 0 2
rlabel polysilicon 751 -486 751 -486 0 3
rlabel polysilicon 754 -486 754 -486 0 4
rlabel polysilicon 758 -480 758 -480 0 1
rlabel polysilicon 758 -486 758 -486 0 3
rlabel polysilicon 761 -486 761 -486 0 4
rlabel polysilicon 765 -480 765 -480 0 1
rlabel polysilicon 765 -486 765 -486 0 3
rlabel polysilicon 772 -486 772 -486 0 3
rlabel polysilicon 779 -480 779 -480 0 1
rlabel polysilicon 779 -486 779 -486 0 3
rlabel polysilicon 786 -480 786 -480 0 1
rlabel polysilicon 789 -480 789 -480 0 2
rlabel polysilicon 786 -486 786 -486 0 3
rlabel polysilicon 789 -486 789 -486 0 4
rlabel polysilicon 793 -480 793 -480 0 1
rlabel polysilicon 793 -486 793 -486 0 3
rlabel polysilicon 800 -480 800 -480 0 1
rlabel polysilicon 800 -486 800 -486 0 3
rlabel polysilicon 807 -480 807 -480 0 1
rlabel polysilicon 807 -486 807 -486 0 3
rlabel polysilicon 814 -480 814 -480 0 1
rlabel polysilicon 814 -486 814 -486 0 3
rlabel polysilicon 821 -480 821 -480 0 1
rlabel polysilicon 821 -486 821 -486 0 3
rlabel polysilicon 831 -480 831 -480 0 2
rlabel polysilicon 828 -486 828 -486 0 3
rlabel polysilicon 831 -486 831 -486 0 4
rlabel polysilicon 835 -480 835 -480 0 1
rlabel polysilicon 835 -486 835 -486 0 3
rlabel polysilicon 842 -480 842 -480 0 1
rlabel polysilicon 842 -486 842 -486 0 3
rlabel polysilicon 849 -480 849 -480 0 1
rlabel polysilicon 849 -486 849 -486 0 3
rlabel polysilicon 856 -480 856 -480 0 1
rlabel polysilicon 856 -486 856 -486 0 3
rlabel polysilicon 863 -480 863 -480 0 1
rlabel polysilicon 863 -486 863 -486 0 3
rlabel polysilicon 870 -480 870 -480 0 1
rlabel polysilicon 870 -486 870 -486 0 3
rlabel polysilicon 877 -480 877 -480 0 1
rlabel polysilicon 877 -486 877 -486 0 3
rlabel polysilicon 884 -480 884 -480 0 1
rlabel polysilicon 887 -480 887 -480 0 2
rlabel polysilicon 884 -486 884 -486 0 3
rlabel polysilicon 887 -486 887 -486 0 4
rlabel polysilicon 891 -480 891 -480 0 1
rlabel polysilicon 891 -486 891 -486 0 3
rlabel polysilicon 898 -480 898 -480 0 1
rlabel polysilicon 898 -486 898 -486 0 3
rlabel polysilicon 905 -480 905 -480 0 1
rlabel polysilicon 905 -486 905 -486 0 3
rlabel polysilicon 912 -480 912 -480 0 1
rlabel polysilicon 912 -486 912 -486 0 3
rlabel polysilicon 919 -480 919 -480 0 1
rlabel polysilicon 919 -486 919 -486 0 3
rlabel polysilicon 926 -480 926 -480 0 1
rlabel polysilicon 926 -486 926 -486 0 3
rlabel polysilicon 933 -480 933 -480 0 1
rlabel polysilicon 933 -486 933 -486 0 3
rlabel polysilicon 940 -480 940 -480 0 1
rlabel polysilicon 940 -486 940 -486 0 3
rlabel polysilicon 947 -480 947 -480 0 1
rlabel polysilicon 947 -486 947 -486 0 3
rlabel polysilicon 954 -480 954 -480 0 1
rlabel polysilicon 954 -486 954 -486 0 3
rlabel polysilicon 961 -480 961 -480 0 1
rlabel polysilicon 961 -486 961 -486 0 3
rlabel polysilicon 968 -480 968 -480 0 1
rlabel polysilicon 968 -486 968 -486 0 3
rlabel polysilicon 975 -480 975 -480 0 1
rlabel polysilicon 975 -486 975 -486 0 3
rlabel polysilicon 982 -480 982 -480 0 1
rlabel polysilicon 982 -486 982 -486 0 3
rlabel polysilicon 989 -480 989 -480 0 1
rlabel polysilicon 989 -486 989 -486 0 3
rlabel polysilicon 996 -480 996 -480 0 1
rlabel polysilicon 996 -486 996 -486 0 3
rlabel polysilicon 1003 -480 1003 -480 0 1
rlabel polysilicon 1003 -486 1003 -486 0 3
rlabel polysilicon 1010 -480 1010 -480 0 1
rlabel polysilicon 1010 -486 1010 -486 0 3
rlabel polysilicon 1017 -480 1017 -480 0 1
rlabel polysilicon 1017 -486 1017 -486 0 3
rlabel polysilicon 1024 -480 1024 -480 0 1
rlabel polysilicon 1024 -486 1024 -486 0 3
rlabel polysilicon 1031 -480 1031 -480 0 1
rlabel polysilicon 1031 -486 1031 -486 0 3
rlabel polysilicon 1038 -480 1038 -480 0 1
rlabel polysilicon 1038 -486 1038 -486 0 3
rlabel polysilicon 1045 -480 1045 -480 0 1
rlabel polysilicon 1045 -486 1045 -486 0 3
rlabel polysilicon 1052 -480 1052 -480 0 1
rlabel polysilicon 1052 -486 1052 -486 0 3
rlabel polysilicon 1059 -480 1059 -480 0 1
rlabel polysilicon 1059 -486 1059 -486 0 3
rlabel polysilicon 1066 -480 1066 -480 0 1
rlabel polysilicon 1066 -486 1066 -486 0 3
rlabel polysilicon 1073 -480 1073 -480 0 1
rlabel polysilicon 1073 -486 1073 -486 0 3
rlabel polysilicon 1080 -480 1080 -480 0 1
rlabel polysilicon 1080 -486 1080 -486 0 3
rlabel polysilicon 1087 -480 1087 -480 0 1
rlabel polysilicon 1087 -486 1087 -486 0 3
rlabel polysilicon 1094 -480 1094 -480 0 1
rlabel polysilicon 1094 -486 1094 -486 0 3
rlabel polysilicon 1101 -480 1101 -480 0 1
rlabel polysilicon 1101 -486 1101 -486 0 3
rlabel polysilicon 1108 -480 1108 -480 0 1
rlabel polysilicon 1108 -486 1108 -486 0 3
rlabel polysilicon 1115 -480 1115 -480 0 1
rlabel polysilicon 1115 -486 1115 -486 0 3
rlabel polysilicon 1122 -480 1122 -480 0 1
rlabel polysilicon 1122 -486 1122 -486 0 3
rlabel polysilicon 1129 -480 1129 -480 0 1
rlabel polysilicon 1129 -486 1129 -486 0 3
rlabel polysilicon 1136 -480 1136 -480 0 1
rlabel polysilicon 1136 -486 1136 -486 0 3
rlabel polysilicon 1143 -480 1143 -480 0 1
rlabel polysilicon 1143 -486 1143 -486 0 3
rlabel polysilicon 1150 -480 1150 -480 0 1
rlabel polysilicon 1150 -486 1150 -486 0 3
rlabel polysilicon 1157 -480 1157 -480 0 1
rlabel polysilicon 1157 -486 1157 -486 0 3
rlabel polysilicon 1164 -480 1164 -480 0 1
rlabel polysilicon 1164 -486 1164 -486 0 3
rlabel polysilicon 1171 -480 1171 -480 0 1
rlabel polysilicon 1171 -486 1171 -486 0 3
rlabel polysilicon 1178 -480 1178 -480 0 1
rlabel polysilicon 1178 -486 1178 -486 0 3
rlabel polysilicon 1185 -480 1185 -480 0 1
rlabel polysilicon 1185 -486 1185 -486 0 3
rlabel polysilicon 1192 -480 1192 -480 0 1
rlabel polysilicon 1192 -486 1192 -486 0 3
rlabel polysilicon 1199 -480 1199 -480 0 1
rlabel polysilicon 1199 -486 1199 -486 0 3
rlabel polysilicon 1206 -480 1206 -480 0 1
rlabel polysilicon 1206 -486 1206 -486 0 3
rlabel polysilicon 1213 -480 1213 -480 0 1
rlabel polysilicon 1213 -486 1213 -486 0 3
rlabel polysilicon 1220 -480 1220 -480 0 1
rlabel polysilicon 1220 -486 1220 -486 0 3
rlabel polysilicon 1227 -480 1227 -480 0 1
rlabel polysilicon 1227 -486 1227 -486 0 3
rlabel polysilicon 1234 -480 1234 -480 0 1
rlabel polysilicon 1234 -486 1234 -486 0 3
rlabel polysilicon 1241 -480 1241 -480 0 1
rlabel polysilicon 1241 -486 1241 -486 0 3
rlabel polysilicon 1248 -480 1248 -480 0 1
rlabel polysilicon 1248 -486 1248 -486 0 3
rlabel polysilicon 1255 -480 1255 -480 0 1
rlabel polysilicon 1255 -486 1255 -486 0 3
rlabel polysilicon 1262 -480 1262 -480 0 1
rlabel polysilicon 1262 -486 1262 -486 0 3
rlabel polysilicon 1269 -480 1269 -480 0 1
rlabel polysilicon 1269 -486 1269 -486 0 3
rlabel polysilicon 1276 -480 1276 -480 0 1
rlabel polysilicon 1276 -486 1276 -486 0 3
rlabel polysilicon 1283 -480 1283 -480 0 1
rlabel polysilicon 1283 -486 1283 -486 0 3
rlabel polysilicon 1290 -480 1290 -480 0 1
rlabel polysilicon 1290 -486 1290 -486 0 3
rlabel polysilicon 1297 -480 1297 -480 0 1
rlabel polysilicon 1297 -486 1297 -486 0 3
rlabel polysilicon 1304 -480 1304 -480 0 1
rlabel polysilicon 1304 -486 1304 -486 0 3
rlabel polysilicon 1311 -480 1311 -480 0 1
rlabel polysilicon 1311 -486 1311 -486 0 3
rlabel polysilicon 1318 -480 1318 -480 0 1
rlabel polysilicon 1318 -486 1318 -486 0 3
rlabel polysilicon 1325 -480 1325 -480 0 1
rlabel polysilicon 1325 -486 1325 -486 0 3
rlabel polysilicon 1332 -480 1332 -480 0 1
rlabel polysilicon 1332 -486 1332 -486 0 3
rlabel polysilicon 1339 -480 1339 -480 0 1
rlabel polysilicon 1339 -486 1339 -486 0 3
rlabel polysilicon 1346 -480 1346 -480 0 1
rlabel polysilicon 1346 -486 1346 -486 0 3
rlabel polysilicon 1353 -480 1353 -480 0 1
rlabel polysilicon 1353 -486 1353 -486 0 3
rlabel polysilicon 1360 -480 1360 -480 0 1
rlabel polysilicon 1360 -486 1360 -486 0 3
rlabel polysilicon 1367 -480 1367 -480 0 1
rlabel polysilicon 1367 -486 1367 -486 0 3
rlabel polysilicon 1374 -480 1374 -480 0 1
rlabel polysilicon 1377 -486 1377 -486 0 4
rlabel polysilicon 40 -613 40 -613 0 2
rlabel polysilicon 51 -613 51 -613 0 1
rlabel polysilicon 51 -619 51 -619 0 3
rlabel polysilicon 58 -613 58 -613 0 1
rlabel polysilicon 58 -619 58 -619 0 3
rlabel polysilicon 65 -613 65 -613 0 1
rlabel polysilicon 68 -613 68 -613 0 2
rlabel polysilicon 65 -619 65 -619 0 3
rlabel polysilicon 68 -619 68 -619 0 4
rlabel polysilicon 72 -613 72 -613 0 1
rlabel polysilicon 72 -619 72 -619 0 3
rlabel polysilicon 79 -613 79 -613 0 1
rlabel polysilicon 82 -619 82 -619 0 4
rlabel polysilicon 86 -613 86 -613 0 1
rlabel polysilicon 86 -619 86 -619 0 3
rlabel polysilicon 100 -613 100 -613 0 1
rlabel polysilicon 100 -619 100 -619 0 3
rlabel polysilicon 107 -613 107 -613 0 1
rlabel polysilicon 107 -619 107 -619 0 3
rlabel polysilicon 114 -613 114 -613 0 1
rlabel polysilicon 117 -619 117 -619 0 4
rlabel polysilicon 121 -613 121 -613 0 1
rlabel polysilicon 121 -619 121 -619 0 3
rlabel polysilicon 128 -613 128 -613 0 1
rlabel polysilicon 128 -619 128 -619 0 3
rlabel polysilicon 135 -613 135 -613 0 1
rlabel polysilicon 135 -619 135 -619 0 3
rlabel polysilicon 138 -619 138 -619 0 4
rlabel polysilicon 142 -613 142 -613 0 1
rlabel polysilicon 142 -619 142 -619 0 3
rlabel polysilicon 149 -613 149 -613 0 1
rlabel polysilicon 152 -613 152 -613 0 2
rlabel polysilicon 149 -619 149 -619 0 3
rlabel polysilicon 152 -619 152 -619 0 4
rlabel polysilicon 156 -613 156 -613 0 1
rlabel polysilicon 159 -613 159 -613 0 2
rlabel polysilicon 156 -619 156 -619 0 3
rlabel polysilicon 159 -619 159 -619 0 4
rlabel polysilicon 163 -613 163 -613 0 1
rlabel polysilicon 163 -619 163 -619 0 3
rlabel polysilicon 177 -613 177 -613 0 1
rlabel polysilicon 177 -619 177 -619 0 3
rlabel polysilicon 184 -613 184 -613 0 1
rlabel polysilicon 184 -619 184 -619 0 3
rlabel polysilicon 191 -613 191 -613 0 1
rlabel polysilicon 191 -619 191 -619 0 3
rlabel polysilicon 198 -613 198 -613 0 1
rlabel polysilicon 198 -619 198 -619 0 3
rlabel polysilicon 201 -619 201 -619 0 4
rlabel polysilicon 205 -613 205 -613 0 1
rlabel polysilicon 205 -619 205 -619 0 3
rlabel polysilicon 212 -613 212 -613 0 1
rlabel polysilicon 212 -619 212 -619 0 3
rlabel polysilicon 219 -613 219 -613 0 1
rlabel polysilicon 222 -613 222 -613 0 2
rlabel polysilicon 219 -619 219 -619 0 3
rlabel polysilicon 226 -613 226 -613 0 1
rlabel polysilicon 226 -619 226 -619 0 3
rlabel polysilicon 243 -613 243 -613 0 2
rlabel polysilicon 243 -619 243 -619 0 4
rlabel polysilicon 250 -613 250 -613 0 2
rlabel polysilicon 247 -619 247 -619 0 3
rlabel polysilicon 250 -619 250 -619 0 4
rlabel polysilicon 261 -613 261 -613 0 1
rlabel polysilicon 261 -619 261 -619 0 3
rlabel polysilicon 268 -613 268 -613 0 1
rlabel polysilicon 268 -619 268 -619 0 3
rlabel polysilicon 275 -613 275 -613 0 1
rlabel polysilicon 275 -619 275 -619 0 3
rlabel polysilicon 282 -613 282 -613 0 1
rlabel polysilicon 282 -619 282 -619 0 3
rlabel polysilicon 289 -613 289 -613 0 1
rlabel polysilicon 289 -619 289 -619 0 3
rlabel polysilicon 296 -613 296 -613 0 1
rlabel polysilicon 296 -619 296 -619 0 3
rlabel polysilicon 303 -613 303 -613 0 1
rlabel polysilicon 303 -619 303 -619 0 3
rlabel polysilicon 310 -613 310 -613 0 1
rlabel polysilicon 310 -619 310 -619 0 3
rlabel polysilicon 317 -613 317 -613 0 1
rlabel polysilicon 317 -619 317 -619 0 3
rlabel polysilicon 324 -613 324 -613 0 1
rlabel polysilicon 324 -619 324 -619 0 3
rlabel polysilicon 331 -613 331 -613 0 1
rlabel polysilicon 331 -619 331 -619 0 3
rlabel polysilicon 338 -613 338 -613 0 1
rlabel polysilicon 338 -619 338 -619 0 3
rlabel polysilicon 345 -613 345 -613 0 1
rlabel polysilicon 345 -619 345 -619 0 3
rlabel polysilicon 352 -613 352 -613 0 1
rlabel polysilicon 352 -619 352 -619 0 3
rlabel polysilicon 359 -613 359 -613 0 1
rlabel polysilicon 359 -619 359 -619 0 3
rlabel polysilicon 373 -613 373 -613 0 1
rlabel polysilicon 373 -619 373 -619 0 3
rlabel polysilicon 380 -613 380 -613 0 1
rlabel polysilicon 380 -619 380 -619 0 3
rlabel polysilicon 387 -613 387 -613 0 1
rlabel polysilicon 387 -619 387 -619 0 3
rlabel polysilicon 394 -613 394 -613 0 1
rlabel polysilicon 397 -613 397 -613 0 2
rlabel polysilicon 394 -619 394 -619 0 3
rlabel polysilicon 397 -619 397 -619 0 4
rlabel polysilicon 401 -613 401 -613 0 1
rlabel polysilicon 401 -619 401 -619 0 3
rlabel polysilicon 408 -613 408 -613 0 1
rlabel polysilicon 408 -619 408 -619 0 3
rlabel polysilicon 415 -613 415 -613 0 1
rlabel polysilicon 415 -619 415 -619 0 3
rlabel polysilicon 422 -613 422 -613 0 1
rlabel polysilicon 422 -619 422 -619 0 3
rlabel polysilicon 429 -613 429 -613 0 1
rlabel polysilicon 429 -619 429 -619 0 3
rlabel polysilicon 436 -613 436 -613 0 1
rlabel polysilicon 436 -619 436 -619 0 3
rlabel polysilicon 443 -613 443 -613 0 1
rlabel polysilicon 443 -619 443 -619 0 3
rlabel polysilicon 450 -613 450 -613 0 1
rlabel polysilicon 450 -619 450 -619 0 3
rlabel polysilicon 457 -613 457 -613 0 1
rlabel polysilicon 457 -619 457 -619 0 3
rlabel polysilicon 464 -613 464 -613 0 1
rlabel polysilicon 464 -619 464 -619 0 3
rlabel polysilicon 471 -613 471 -613 0 1
rlabel polysilicon 471 -619 471 -619 0 3
rlabel polysilicon 478 -613 478 -613 0 1
rlabel polysilicon 478 -619 478 -619 0 3
rlabel polysilicon 485 -613 485 -613 0 1
rlabel polysilicon 485 -619 485 -619 0 3
rlabel polysilicon 492 -613 492 -613 0 1
rlabel polysilicon 492 -619 492 -619 0 3
rlabel polysilicon 499 -613 499 -613 0 1
rlabel polysilicon 502 -613 502 -613 0 2
rlabel polysilicon 502 -619 502 -619 0 4
rlabel polysilicon 506 -613 506 -613 0 1
rlabel polysilicon 506 -619 506 -619 0 3
rlabel polysilicon 513 -613 513 -613 0 1
rlabel polysilicon 513 -619 513 -619 0 3
rlabel polysilicon 516 -619 516 -619 0 4
rlabel polysilicon 520 -613 520 -613 0 1
rlabel polysilicon 520 -619 520 -619 0 3
rlabel polysilicon 527 -613 527 -613 0 1
rlabel polysilicon 530 -613 530 -613 0 2
rlabel polysilicon 527 -619 527 -619 0 3
rlabel polysilicon 530 -619 530 -619 0 4
rlabel polysilicon 534 -613 534 -613 0 1
rlabel polysilicon 534 -619 534 -619 0 3
rlabel polysilicon 541 -613 541 -613 0 1
rlabel polysilicon 544 -613 544 -613 0 2
rlabel polysilicon 541 -619 541 -619 0 3
rlabel polysilicon 548 -613 548 -613 0 1
rlabel polysilicon 548 -619 548 -619 0 3
rlabel polysilicon 555 -613 555 -613 0 1
rlabel polysilicon 555 -619 555 -619 0 3
rlabel polysilicon 562 -613 562 -613 0 1
rlabel polysilicon 562 -619 562 -619 0 3
rlabel polysilicon 569 -613 569 -613 0 1
rlabel polysilicon 569 -619 569 -619 0 3
rlabel polysilicon 576 -613 576 -613 0 1
rlabel polysilicon 576 -619 576 -619 0 3
rlabel polysilicon 583 -613 583 -613 0 1
rlabel polysilicon 586 -613 586 -613 0 2
rlabel polysilicon 583 -619 583 -619 0 3
rlabel polysilicon 586 -619 586 -619 0 4
rlabel polysilicon 590 -613 590 -613 0 1
rlabel polysilicon 590 -619 590 -619 0 3
rlabel polysilicon 597 -613 597 -613 0 1
rlabel polysilicon 597 -619 597 -619 0 3
rlabel polysilicon 604 -613 604 -613 0 1
rlabel polysilicon 604 -619 604 -619 0 3
rlabel polysilicon 611 -613 611 -613 0 1
rlabel polysilicon 611 -619 611 -619 0 3
rlabel polysilicon 618 -613 618 -613 0 1
rlabel polysilicon 618 -619 618 -619 0 3
rlabel polysilicon 625 -613 625 -613 0 1
rlabel polysilicon 625 -619 625 -619 0 3
rlabel polysilicon 632 -613 632 -613 0 1
rlabel polysilicon 632 -619 632 -619 0 3
rlabel polysilicon 639 -613 639 -613 0 1
rlabel polysilicon 639 -619 639 -619 0 3
rlabel polysilicon 646 -613 646 -613 0 1
rlabel polysilicon 646 -619 646 -619 0 3
rlabel polysilicon 653 -613 653 -613 0 1
rlabel polysilicon 653 -619 653 -619 0 3
rlabel polysilicon 660 -613 660 -613 0 1
rlabel polysilicon 660 -619 660 -619 0 3
rlabel polysilicon 670 -613 670 -613 0 2
rlabel polysilicon 667 -619 667 -619 0 3
rlabel polysilicon 670 -619 670 -619 0 4
rlabel polysilicon 674 -613 674 -613 0 1
rlabel polysilicon 674 -619 674 -619 0 3
rlabel polysilicon 681 -613 681 -613 0 1
rlabel polysilicon 684 -613 684 -613 0 2
rlabel polysilicon 684 -619 684 -619 0 4
rlabel polysilicon 688 -613 688 -613 0 1
rlabel polysilicon 688 -619 688 -619 0 3
rlabel polysilicon 695 -613 695 -613 0 1
rlabel polysilicon 698 -613 698 -613 0 2
rlabel polysilicon 695 -619 695 -619 0 3
rlabel polysilicon 698 -619 698 -619 0 4
rlabel polysilicon 702 -613 702 -613 0 1
rlabel polysilicon 705 -613 705 -613 0 2
rlabel polysilicon 702 -619 702 -619 0 3
rlabel polysilicon 705 -619 705 -619 0 4
rlabel polysilicon 709 -613 709 -613 0 1
rlabel polysilicon 709 -619 709 -619 0 3
rlabel polysilicon 716 -613 716 -613 0 1
rlabel polysilicon 716 -619 716 -619 0 3
rlabel polysilicon 719 -619 719 -619 0 4
rlabel polysilicon 723 -613 723 -613 0 1
rlabel polysilicon 723 -619 723 -619 0 3
rlabel polysilicon 730 -613 730 -613 0 1
rlabel polysilicon 733 -613 733 -613 0 2
rlabel polysilicon 733 -619 733 -619 0 4
rlabel polysilicon 737 -613 737 -613 0 1
rlabel polysilicon 737 -619 737 -619 0 3
rlabel polysilicon 744 -613 744 -613 0 1
rlabel polysilicon 744 -619 744 -619 0 3
rlabel polysilicon 751 -613 751 -613 0 1
rlabel polysilicon 751 -619 751 -619 0 3
rlabel polysilicon 758 -613 758 -613 0 1
rlabel polysilicon 758 -619 758 -619 0 3
rlabel polysilicon 765 -613 765 -613 0 1
rlabel polysilicon 768 -613 768 -613 0 2
rlabel polysilicon 765 -619 765 -619 0 3
rlabel polysilicon 768 -619 768 -619 0 4
rlabel polysilicon 775 -613 775 -613 0 2
rlabel polysilicon 772 -619 772 -619 0 3
rlabel polysilicon 775 -619 775 -619 0 4
rlabel polysilicon 779 -613 779 -613 0 1
rlabel polysilicon 782 -613 782 -613 0 2
rlabel polysilicon 779 -619 779 -619 0 3
rlabel polysilicon 786 -613 786 -613 0 1
rlabel polysilicon 786 -619 786 -619 0 3
rlabel polysilicon 793 -613 793 -613 0 1
rlabel polysilicon 793 -619 793 -619 0 3
rlabel polysilicon 796 -619 796 -619 0 4
rlabel polysilicon 800 -613 800 -613 0 1
rlabel polysilicon 800 -619 800 -619 0 3
rlabel polysilicon 807 -613 807 -613 0 1
rlabel polysilicon 810 -613 810 -613 0 2
rlabel polysilicon 807 -619 807 -619 0 3
rlabel polysilicon 814 -613 814 -613 0 1
rlabel polysilicon 814 -619 814 -619 0 3
rlabel polysilicon 821 -613 821 -613 0 1
rlabel polysilicon 821 -619 821 -619 0 3
rlabel polysilicon 828 -613 828 -613 0 1
rlabel polysilicon 828 -619 828 -619 0 3
rlabel polysilicon 835 -613 835 -613 0 1
rlabel polysilicon 835 -619 835 -619 0 3
rlabel polysilicon 842 -613 842 -613 0 1
rlabel polysilicon 842 -619 842 -619 0 3
rlabel polysilicon 849 -613 849 -613 0 1
rlabel polysilicon 849 -619 849 -619 0 3
rlabel polysilicon 856 -613 856 -613 0 1
rlabel polysilicon 856 -619 856 -619 0 3
rlabel polysilicon 863 -613 863 -613 0 1
rlabel polysilicon 863 -619 863 -619 0 3
rlabel polysilicon 870 -613 870 -613 0 1
rlabel polysilicon 870 -619 870 -619 0 3
rlabel polysilicon 877 -613 877 -613 0 1
rlabel polysilicon 877 -619 877 -619 0 3
rlabel polysilicon 884 -613 884 -613 0 1
rlabel polysilicon 884 -619 884 -619 0 3
rlabel polysilicon 891 -613 891 -613 0 1
rlabel polysilicon 891 -619 891 -619 0 3
rlabel polysilicon 898 -613 898 -613 0 1
rlabel polysilicon 901 -613 901 -613 0 2
rlabel polysilicon 898 -619 898 -619 0 3
rlabel polysilicon 901 -619 901 -619 0 4
rlabel polysilicon 905 -613 905 -613 0 1
rlabel polysilicon 905 -619 905 -619 0 3
rlabel polysilicon 912 -613 912 -613 0 1
rlabel polysilicon 912 -619 912 -619 0 3
rlabel polysilicon 919 -613 919 -613 0 1
rlabel polysilicon 919 -619 919 -619 0 3
rlabel polysilicon 926 -613 926 -613 0 1
rlabel polysilicon 926 -619 926 -619 0 3
rlabel polysilicon 933 -613 933 -613 0 1
rlabel polysilicon 933 -619 933 -619 0 3
rlabel polysilicon 940 -613 940 -613 0 1
rlabel polysilicon 940 -619 940 -619 0 3
rlabel polysilicon 947 -613 947 -613 0 1
rlabel polysilicon 947 -619 947 -619 0 3
rlabel polysilicon 954 -613 954 -613 0 1
rlabel polysilicon 954 -619 954 -619 0 3
rlabel polysilicon 961 -613 961 -613 0 1
rlabel polysilicon 961 -619 961 -619 0 3
rlabel polysilicon 968 -613 968 -613 0 1
rlabel polysilicon 968 -619 968 -619 0 3
rlabel polysilicon 975 -613 975 -613 0 1
rlabel polysilicon 978 -613 978 -613 0 2
rlabel polysilicon 978 -619 978 -619 0 4
rlabel polysilicon 982 -613 982 -613 0 1
rlabel polysilicon 982 -619 982 -619 0 3
rlabel polysilicon 989 -613 989 -613 0 1
rlabel polysilicon 989 -619 989 -619 0 3
rlabel polysilicon 996 -613 996 -613 0 1
rlabel polysilicon 996 -619 996 -619 0 3
rlabel polysilicon 1003 -613 1003 -613 0 1
rlabel polysilicon 1003 -619 1003 -619 0 3
rlabel polysilicon 1010 -613 1010 -613 0 1
rlabel polysilicon 1010 -619 1010 -619 0 3
rlabel polysilicon 1017 -613 1017 -613 0 1
rlabel polysilicon 1017 -619 1017 -619 0 3
rlabel polysilicon 1024 -613 1024 -613 0 1
rlabel polysilicon 1024 -619 1024 -619 0 3
rlabel polysilicon 1031 -613 1031 -613 0 1
rlabel polysilicon 1031 -619 1031 -619 0 3
rlabel polysilicon 1038 -613 1038 -613 0 1
rlabel polysilicon 1038 -619 1038 -619 0 3
rlabel polysilicon 1045 -613 1045 -613 0 1
rlabel polysilicon 1045 -619 1045 -619 0 3
rlabel polysilicon 1052 -613 1052 -613 0 1
rlabel polysilicon 1052 -619 1052 -619 0 3
rlabel polysilicon 1059 -613 1059 -613 0 1
rlabel polysilicon 1059 -619 1059 -619 0 3
rlabel polysilicon 1066 -613 1066 -613 0 1
rlabel polysilicon 1066 -619 1066 -619 0 3
rlabel polysilicon 1073 -613 1073 -613 0 1
rlabel polysilicon 1073 -619 1073 -619 0 3
rlabel polysilicon 1080 -613 1080 -613 0 1
rlabel polysilicon 1080 -619 1080 -619 0 3
rlabel polysilicon 1087 -613 1087 -613 0 1
rlabel polysilicon 1087 -619 1087 -619 0 3
rlabel polysilicon 1094 -613 1094 -613 0 1
rlabel polysilicon 1094 -619 1094 -619 0 3
rlabel polysilicon 1101 -613 1101 -613 0 1
rlabel polysilicon 1101 -619 1101 -619 0 3
rlabel polysilicon 1108 -613 1108 -613 0 1
rlabel polysilicon 1108 -619 1108 -619 0 3
rlabel polysilicon 1115 -613 1115 -613 0 1
rlabel polysilicon 1115 -619 1115 -619 0 3
rlabel polysilicon 1122 -613 1122 -613 0 1
rlabel polysilicon 1122 -619 1122 -619 0 3
rlabel polysilicon 1129 -613 1129 -613 0 1
rlabel polysilicon 1129 -619 1129 -619 0 3
rlabel polysilicon 1136 -613 1136 -613 0 1
rlabel polysilicon 1136 -619 1136 -619 0 3
rlabel polysilicon 1143 -613 1143 -613 0 1
rlabel polysilicon 1143 -619 1143 -619 0 3
rlabel polysilicon 1150 -613 1150 -613 0 1
rlabel polysilicon 1150 -619 1150 -619 0 3
rlabel polysilicon 1157 -613 1157 -613 0 1
rlabel polysilicon 1157 -619 1157 -619 0 3
rlabel polysilicon 1164 -613 1164 -613 0 1
rlabel polysilicon 1164 -619 1164 -619 0 3
rlabel polysilicon 1171 -613 1171 -613 0 1
rlabel polysilicon 1171 -619 1171 -619 0 3
rlabel polysilicon 1178 -613 1178 -613 0 1
rlabel polysilicon 1178 -619 1178 -619 0 3
rlabel polysilicon 1185 -613 1185 -613 0 1
rlabel polysilicon 1185 -619 1185 -619 0 3
rlabel polysilicon 1192 -613 1192 -613 0 1
rlabel polysilicon 1192 -619 1192 -619 0 3
rlabel polysilicon 1199 -613 1199 -613 0 1
rlabel polysilicon 1199 -619 1199 -619 0 3
rlabel polysilicon 1206 -613 1206 -613 0 1
rlabel polysilicon 1206 -619 1206 -619 0 3
rlabel polysilicon 1213 -613 1213 -613 0 1
rlabel polysilicon 1213 -619 1213 -619 0 3
rlabel polysilicon 1220 -613 1220 -613 0 1
rlabel polysilicon 1220 -619 1220 -619 0 3
rlabel polysilicon 1227 -613 1227 -613 0 1
rlabel polysilicon 1227 -619 1227 -619 0 3
rlabel polysilicon 1234 -613 1234 -613 0 1
rlabel polysilicon 1234 -619 1234 -619 0 3
rlabel polysilicon 1241 -613 1241 -613 0 1
rlabel polysilicon 1241 -619 1241 -619 0 3
rlabel polysilicon 1248 -613 1248 -613 0 1
rlabel polysilicon 1248 -619 1248 -619 0 3
rlabel polysilicon 1255 -613 1255 -613 0 1
rlabel polysilicon 1255 -619 1255 -619 0 3
rlabel polysilicon 1262 -613 1262 -613 0 1
rlabel polysilicon 1262 -619 1262 -619 0 3
rlabel polysilicon 1269 -613 1269 -613 0 1
rlabel polysilicon 1269 -619 1269 -619 0 3
rlabel polysilicon 1276 -613 1276 -613 0 1
rlabel polysilicon 1276 -619 1276 -619 0 3
rlabel polysilicon 1283 -613 1283 -613 0 1
rlabel polysilicon 1283 -619 1283 -619 0 3
rlabel polysilicon 1290 -613 1290 -613 0 1
rlabel polysilicon 1290 -619 1290 -619 0 3
rlabel polysilicon 1297 -613 1297 -613 0 1
rlabel polysilicon 1297 -619 1297 -619 0 3
rlabel polysilicon 1304 -613 1304 -613 0 1
rlabel polysilicon 1304 -619 1304 -619 0 3
rlabel polysilicon 1311 -613 1311 -613 0 1
rlabel polysilicon 1311 -619 1311 -619 0 3
rlabel polysilicon 1318 -613 1318 -613 0 1
rlabel polysilicon 1318 -619 1318 -619 0 3
rlabel polysilicon 1325 -613 1325 -613 0 1
rlabel polysilicon 1325 -619 1325 -619 0 3
rlabel polysilicon 1332 -613 1332 -613 0 1
rlabel polysilicon 1332 -619 1332 -619 0 3
rlabel polysilicon 1339 -613 1339 -613 0 1
rlabel polysilicon 1339 -619 1339 -619 0 3
rlabel polysilicon 1346 -613 1346 -613 0 1
rlabel polysilicon 1346 -619 1346 -619 0 3
rlabel polysilicon 1353 -613 1353 -613 0 1
rlabel polysilicon 1353 -619 1353 -619 0 3
rlabel polysilicon 1356 -619 1356 -619 0 4
rlabel polysilicon 1360 -613 1360 -613 0 1
rlabel polysilicon 1360 -619 1360 -619 0 3
rlabel polysilicon 1367 -613 1367 -613 0 1
rlabel polysilicon 1367 -619 1367 -619 0 3
rlabel polysilicon 1374 -613 1374 -613 0 1
rlabel polysilicon 1374 -619 1374 -619 0 3
rlabel polysilicon 1381 -613 1381 -613 0 1
rlabel polysilicon 1381 -619 1381 -619 0 3
rlabel polysilicon 1388 -613 1388 -613 0 1
rlabel polysilicon 1388 -619 1388 -619 0 3
rlabel polysilicon 1472 -613 1472 -613 0 1
rlabel polysilicon 1472 -619 1472 -619 0 3
rlabel polysilicon 44 -736 44 -736 0 1
rlabel polysilicon 44 -742 44 -742 0 3
rlabel polysilicon 51 -736 51 -736 0 1
rlabel polysilicon 51 -742 51 -742 0 3
rlabel polysilicon 58 -736 58 -736 0 1
rlabel polysilicon 58 -742 58 -742 0 3
rlabel polysilicon 65 -736 65 -736 0 1
rlabel polysilicon 65 -742 65 -742 0 3
rlabel polysilicon 72 -736 72 -736 0 1
rlabel polysilicon 72 -742 72 -742 0 3
rlabel polysilicon 82 -736 82 -736 0 2
rlabel polysilicon 79 -742 79 -742 0 3
rlabel polysilicon 82 -742 82 -742 0 4
rlabel polysilicon 86 -736 86 -736 0 1
rlabel polysilicon 86 -742 86 -742 0 3
rlabel polysilicon 93 -736 93 -736 0 1
rlabel polysilicon 96 -736 96 -736 0 2
rlabel polysilicon 93 -742 93 -742 0 3
rlabel polysilicon 100 -736 100 -736 0 1
rlabel polysilicon 100 -742 100 -742 0 3
rlabel polysilicon 107 -736 107 -736 0 1
rlabel polysilicon 107 -742 107 -742 0 3
rlabel polysilicon 114 -736 114 -736 0 1
rlabel polysilicon 114 -742 114 -742 0 3
rlabel polysilicon 121 -736 121 -736 0 1
rlabel polysilicon 124 -736 124 -736 0 2
rlabel polysilicon 121 -742 121 -742 0 3
rlabel polysilicon 124 -742 124 -742 0 4
rlabel polysilicon 128 -736 128 -736 0 1
rlabel polysilicon 128 -742 128 -742 0 3
rlabel polysilicon 135 -736 135 -736 0 1
rlabel polysilicon 135 -742 135 -742 0 3
rlabel polysilicon 149 -736 149 -736 0 1
rlabel polysilicon 149 -742 149 -742 0 3
rlabel polysilicon 156 -736 156 -736 0 1
rlabel polysilicon 156 -742 156 -742 0 3
rlabel polysilicon 163 -736 163 -736 0 1
rlabel polysilicon 163 -742 163 -742 0 3
rlabel polysilicon 170 -736 170 -736 0 1
rlabel polysilicon 170 -742 170 -742 0 3
rlabel polysilicon 177 -736 177 -736 0 1
rlabel polysilicon 177 -742 177 -742 0 3
rlabel polysilicon 184 -736 184 -736 0 1
rlabel polysilicon 187 -736 187 -736 0 2
rlabel polysilicon 184 -742 184 -742 0 3
rlabel polysilicon 187 -742 187 -742 0 4
rlabel polysilicon 191 -736 191 -736 0 1
rlabel polysilicon 191 -742 191 -742 0 3
rlabel polysilicon 198 -736 198 -736 0 1
rlabel polysilicon 198 -742 198 -742 0 3
rlabel polysilicon 205 -736 205 -736 0 1
rlabel polysilicon 205 -742 205 -742 0 3
rlabel polysilicon 212 -736 212 -736 0 1
rlabel polysilicon 212 -742 212 -742 0 3
rlabel polysilicon 219 -736 219 -736 0 1
rlabel polysilicon 219 -742 219 -742 0 3
rlabel polysilicon 226 -736 226 -736 0 1
rlabel polysilicon 226 -742 226 -742 0 3
rlabel polysilicon 233 -736 233 -736 0 1
rlabel polysilicon 233 -742 233 -742 0 3
rlabel polysilicon 240 -736 240 -736 0 1
rlabel polysilicon 240 -742 240 -742 0 3
rlabel polysilicon 247 -736 247 -736 0 1
rlabel polysilicon 250 -736 250 -736 0 2
rlabel polysilicon 250 -742 250 -742 0 4
rlabel polysilicon 254 -736 254 -736 0 1
rlabel polysilicon 254 -742 254 -742 0 3
rlabel polysilicon 261 -736 261 -736 0 1
rlabel polysilicon 261 -742 261 -742 0 3
rlabel polysilicon 268 -736 268 -736 0 1
rlabel polysilicon 268 -742 268 -742 0 3
rlabel polysilicon 275 -736 275 -736 0 1
rlabel polysilicon 275 -742 275 -742 0 3
rlabel polysilicon 282 -736 282 -736 0 1
rlabel polysilicon 282 -742 282 -742 0 3
rlabel polysilicon 292 -736 292 -736 0 2
rlabel polysilicon 289 -742 289 -742 0 3
rlabel polysilicon 292 -742 292 -742 0 4
rlabel polysilicon 296 -736 296 -736 0 1
rlabel polysilicon 296 -742 296 -742 0 3
rlabel polysilicon 303 -736 303 -736 0 1
rlabel polysilicon 303 -742 303 -742 0 3
rlabel polysilicon 310 -736 310 -736 0 1
rlabel polysilicon 310 -742 310 -742 0 3
rlabel polysilicon 317 -736 317 -736 0 1
rlabel polysilicon 317 -742 317 -742 0 3
rlabel polysilicon 324 -736 324 -736 0 1
rlabel polysilicon 324 -742 324 -742 0 3
rlabel polysilicon 331 -736 331 -736 0 1
rlabel polysilicon 331 -742 331 -742 0 3
rlabel polysilicon 338 -736 338 -736 0 1
rlabel polysilicon 338 -742 338 -742 0 3
rlabel polysilicon 345 -736 345 -736 0 1
rlabel polysilicon 345 -742 345 -742 0 3
rlabel polysilicon 352 -736 352 -736 0 1
rlabel polysilicon 352 -742 352 -742 0 3
rlabel polysilicon 359 -736 359 -736 0 1
rlabel polysilicon 359 -742 359 -742 0 3
rlabel polysilicon 366 -736 366 -736 0 1
rlabel polysilicon 366 -742 366 -742 0 3
rlabel polysilicon 373 -736 373 -736 0 1
rlabel polysilicon 373 -742 373 -742 0 3
rlabel polysilicon 380 -736 380 -736 0 1
rlabel polysilicon 380 -742 380 -742 0 3
rlabel polysilicon 387 -736 387 -736 0 1
rlabel polysilicon 387 -742 387 -742 0 3
rlabel polysilicon 394 -736 394 -736 0 1
rlabel polysilicon 394 -742 394 -742 0 3
rlabel polysilicon 401 -736 401 -736 0 1
rlabel polysilicon 401 -742 401 -742 0 3
rlabel polysilicon 408 -736 408 -736 0 1
rlabel polysilicon 408 -742 408 -742 0 3
rlabel polysilicon 415 -736 415 -736 0 1
rlabel polysilicon 415 -742 415 -742 0 3
rlabel polysilicon 422 -736 422 -736 0 1
rlabel polysilicon 422 -742 422 -742 0 3
rlabel polysilicon 429 -736 429 -736 0 1
rlabel polysilicon 432 -736 432 -736 0 2
rlabel polysilicon 429 -742 429 -742 0 3
rlabel polysilicon 432 -742 432 -742 0 4
rlabel polysilicon 436 -736 436 -736 0 1
rlabel polysilicon 439 -736 439 -736 0 2
rlabel polysilicon 436 -742 436 -742 0 3
rlabel polysilicon 439 -742 439 -742 0 4
rlabel polysilicon 443 -736 443 -736 0 1
rlabel polysilicon 443 -742 443 -742 0 3
rlabel polysilicon 450 -736 450 -736 0 1
rlabel polysilicon 450 -742 450 -742 0 3
rlabel polysilicon 457 -736 457 -736 0 1
rlabel polysilicon 457 -742 457 -742 0 3
rlabel polysilicon 464 -736 464 -736 0 1
rlabel polysilicon 464 -742 464 -742 0 3
rlabel polysilicon 471 -736 471 -736 0 1
rlabel polysilicon 471 -742 471 -742 0 3
rlabel polysilicon 478 -736 478 -736 0 1
rlabel polysilicon 478 -742 478 -742 0 3
rlabel polysilicon 488 -736 488 -736 0 2
rlabel polysilicon 488 -742 488 -742 0 4
rlabel polysilicon 492 -736 492 -736 0 1
rlabel polysilicon 492 -742 492 -742 0 3
rlabel polysilicon 506 -736 506 -736 0 1
rlabel polysilicon 506 -742 506 -742 0 3
rlabel polysilicon 513 -736 513 -736 0 1
rlabel polysilicon 513 -742 513 -742 0 3
rlabel polysilicon 520 -736 520 -736 0 1
rlabel polysilicon 520 -742 520 -742 0 3
rlabel polysilicon 527 -736 527 -736 0 1
rlabel polysilicon 527 -742 527 -742 0 3
rlabel polysilicon 534 -736 534 -736 0 1
rlabel polysilicon 537 -736 537 -736 0 2
rlabel polysilicon 534 -742 534 -742 0 3
rlabel polysilicon 537 -742 537 -742 0 4
rlabel polysilicon 541 -736 541 -736 0 1
rlabel polysilicon 541 -742 541 -742 0 3
rlabel polysilicon 548 -736 548 -736 0 1
rlabel polysilicon 548 -742 548 -742 0 3
rlabel polysilicon 555 -736 555 -736 0 1
rlabel polysilicon 558 -736 558 -736 0 2
rlabel polysilicon 555 -742 555 -742 0 3
rlabel polysilicon 558 -742 558 -742 0 4
rlabel polysilicon 562 -736 562 -736 0 1
rlabel polysilicon 565 -736 565 -736 0 2
rlabel polysilicon 562 -742 562 -742 0 3
rlabel polysilicon 565 -742 565 -742 0 4
rlabel polysilicon 569 -736 569 -736 0 1
rlabel polysilicon 569 -742 569 -742 0 3
rlabel polysilicon 576 -736 576 -736 0 1
rlabel polysilicon 579 -736 579 -736 0 2
rlabel polysilicon 576 -742 576 -742 0 3
rlabel polysilicon 579 -742 579 -742 0 4
rlabel polysilicon 583 -736 583 -736 0 1
rlabel polysilicon 583 -742 583 -742 0 3
rlabel polysilicon 590 -736 590 -736 0 1
rlabel polysilicon 593 -736 593 -736 0 2
rlabel polysilicon 590 -742 590 -742 0 3
rlabel polysilicon 593 -742 593 -742 0 4
rlabel polysilicon 597 -736 597 -736 0 1
rlabel polysilicon 597 -742 597 -742 0 3
rlabel polysilicon 604 -736 604 -736 0 1
rlabel polysilicon 607 -736 607 -736 0 2
rlabel polysilicon 607 -742 607 -742 0 4
rlabel polysilicon 611 -736 611 -736 0 1
rlabel polysilicon 611 -742 611 -742 0 3
rlabel polysilicon 618 -736 618 -736 0 1
rlabel polysilicon 618 -742 618 -742 0 3
rlabel polysilicon 625 -736 625 -736 0 1
rlabel polysilicon 625 -742 625 -742 0 3
rlabel polysilicon 639 -736 639 -736 0 1
rlabel polysilicon 639 -742 639 -742 0 3
rlabel polysilicon 646 -736 646 -736 0 1
rlabel polysilicon 649 -736 649 -736 0 2
rlabel polysilicon 649 -742 649 -742 0 4
rlabel polysilicon 653 -736 653 -736 0 1
rlabel polysilicon 656 -736 656 -736 0 2
rlabel polysilicon 653 -742 653 -742 0 3
rlabel polysilicon 656 -742 656 -742 0 4
rlabel polysilicon 660 -736 660 -736 0 1
rlabel polysilicon 660 -742 660 -742 0 3
rlabel polysilicon 667 -736 667 -736 0 1
rlabel polysilicon 667 -742 667 -742 0 3
rlabel polysilicon 674 -736 674 -736 0 1
rlabel polysilicon 674 -742 674 -742 0 3
rlabel polysilicon 681 -736 681 -736 0 1
rlabel polysilicon 681 -742 681 -742 0 3
rlabel polysilicon 688 -736 688 -736 0 1
rlabel polysilicon 688 -742 688 -742 0 3
rlabel polysilicon 695 -736 695 -736 0 1
rlabel polysilicon 695 -742 695 -742 0 3
rlabel polysilicon 702 -736 702 -736 0 1
rlabel polysilicon 702 -742 702 -742 0 3
rlabel polysilicon 709 -736 709 -736 0 1
rlabel polysilicon 712 -736 712 -736 0 2
rlabel polysilicon 709 -742 709 -742 0 3
rlabel polysilicon 712 -742 712 -742 0 4
rlabel polysilicon 716 -736 716 -736 0 1
rlabel polysilicon 716 -742 716 -742 0 3
rlabel polysilicon 723 -736 723 -736 0 1
rlabel polysilicon 726 -736 726 -736 0 2
rlabel polysilicon 723 -742 723 -742 0 3
rlabel polysilicon 726 -742 726 -742 0 4
rlabel polysilicon 730 -736 730 -736 0 1
rlabel polysilicon 733 -736 733 -736 0 2
rlabel polysilicon 730 -742 730 -742 0 3
rlabel polysilicon 733 -742 733 -742 0 4
rlabel polysilicon 737 -736 737 -736 0 1
rlabel polysilicon 737 -742 737 -742 0 3
rlabel polysilicon 744 -736 744 -736 0 1
rlabel polysilicon 744 -742 744 -742 0 3
rlabel polysilicon 751 -736 751 -736 0 1
rlabel polysilicon 751 -742 751 -742 0 3
rlabel polysilicon 758 -736 758 -736 0 1
rlabel polysilicon 758 -742 758 -742 0 3
rlabel polysilicon 765 -736 765 -736 0 1
rlabel polysilicon 765 -742 765 -742 0 3
rlabel polysilicon 772 -736 772 -736 0 1
rlabel polysilicon 772 -742 772 -742 0 3
rlabel polysilicon 779 -736 779 -736 0 1
rlabel polysilicon 779 -742 779 -742 0 3
rlabel polysilicon 786 -736 786 -736 0 1
rlabel polysilicon 786 -742 786 -742 0 3
rlabel polysilicon 793 -736 793 -736 0 1
rlabel polysilicon 796 -742 796 -742 0 4
rlabel polysilicon 800 -736 800 -736 0 1
rlabel polysilicon 800 -742 800 -742 0 3
rlabel polysilicon 807 -736 807 -736 0 1
rlabel polysilicon 807 -742 807 -742 0 3
rlabel polysilicon 814 -736 814 -736 0 1
rlabel polysilicon 814 -742 814 -742 0 3
rlabel polysilicon 821 -736 821 -736 0 1
rlabel polysilicon 821 -742 821 -742 0 3
rlabel polysilicon 828 -736 828 -736 0 1
rlabel polysilicon 831 -736 831 -736 0 2
rlabel polysilicon 828 -742 828 -742 0 3
rlabel polysilicon 831 -742 831 -742 0 4
rlabel polysilicon 835 -736 835 -736 0 1
rlabel polysilicon 835 -742 835 -742 0 3
rlabel polysilicon 842 -736 842 -736 0 1
rlabel polysilicon 842 -742 842 -742 0 3
rlabel polysilicon 849 -736 849 -736 0 1
rlabel polysilicon 849 -742 849 -742 0 3
rlabel polysilicon 856 -736 856 -736 0 1
rlabel polysilicon 859 -736 859 -736 0 2
rlabel polysilicon 856 -742 856 -742 0 3
rlabel polysilicon 859 -742 859 -742 0 4
rlabel polysilicon 863 -736 863 -736 0 1
rlabel polysilicon 863 -742 863 -742 0 3
rlabel polysilicon 870 -742 870 -742 0 3
rlabel polysilicon 873 -742 873 -742 0 4
rlabel polysilicon 877 -736 877 -736 0 1
rlabel polysilicon 877 -742 877 -742 0 3
rlabel polysilicon 884 -736 884 -736 0 1
rlabel polysilicon 887 -736 887 -736 0 2
rlabel polysilicon 884 -742 884 -742 0 3
rlabel polysilicon 887 -742 887 -742 0 4
rlabel polysilicon 891 -736 891 -736 0 1
rlabel polysilicon 891 -742 891 -742 0 3
rlabel polysilicon 898 -736 898 -736 0 1
rlabel polysilicon 898 -742 898 -742 0 3
rlabel polysilicon 905 -736 905 -736 0 1
rlabel polysilicon 908 -736 908 -736 0 2
rlabel polysilicon 905 -742 905 -742 0 3
rlabel polysilicon 912 -736 912 -736 0 1
rlabel polysilicon 912 -742 912 -742 0 3
rlabel polysilicon 919 -736 919 -736 0 1
rlabel polysilicon 919 -742 919 -742 0 3
rlabel polysilicon 922 -742 922 -742 0 4
rlabel polysilicon 926 -736 926 -736 0 1
rlabel polysilicon 926 -742 926 -742 0 3
rlabel polysilicon 933 -736 933 -736 0 1
rlabel polysilicon 933 -742 933 -742 0 3
rlabel polysilicon 940 -736 940 -736 0 1
rlabel polysilicon 940 -742 940 -742 0 3
rlabel polysilicon 947 -736 947 -736 0 1
rlabel polysilicon 947 -742 947 -742 0 3
rlabel polysilicon 954 -736 954 -736 0 1
rlabel polysilicon 954 -742 954 -742 0 3
rlabel polysilicon 961 -736 961 -736 0 1
rlabel polysilicon 961 -742 961 -742 0 3
rlabel polysilicon 968 -736 968 -736 0 1
rlabel polysilicon 968 -742 968 -742 0 3
rlabel polysilicon 975 -736 975 -736 0 1
rlabel polysilicon 975 -742 975 -742 0 3
rlabel polysilicon 982 -736 982 -736 0 1
rlabel polysilicon 982 -742 982 -742 0 3
rlabel polysilicon 992 -736 992 -736 0 2
rlabel polysilicon 989 -742 989 -742 0 3
rlabel polysilicon 992 -742 992 -742 0 4
rlabel polysilicon 996 -736 996 -736 0 1
rlabel polysilicon 996 -742 996 -742 0 3
rlabel polysilicon 1006 -736 1006 -736 0 2
rlabel polysilicon 1003 -742 1003 -742 0 3
rlabel polysilicon 1006 -742 1006 -742 0 4
rlabel polysilicon 1010 -736 1010 -736 0 1
rlabel polysilicon 1010 -742 1010 -742 0 3
rlabel polysilicon 1017 -736 1017 -736 0 1
rlabel polysilicon 1017 -742 1017 -742 0 3
rlabel polysilicon 1024 -736 1024 -736 0 1
rlabel polysilicon 1024 -742 1024 -742 0 3
rlabel polysilicon 1031 -736 1031 -736 0 1
rlabel polysilicon 1031 -742 1031 -742 0 3
rlabel polysilicon 1038 -736 1038 -736 0 1
rlabel polysilicon 1038 -742 1038 -742 0 3
rlabel polysilicon 1045 -736 1045 -736 0 1
rlabel polysilicon 1045 -742 1045 -742 0 3
rlabel polysilicon 1052 -736 1052 -736 0 1
rlabel polysilicon 1052 -742 1052 -742 0 3
rlabel polysilicon 1059 -736 1059 -736 0 1
rlabel polysilicon 1062 -736 1062 -736 0 2
rlabel polysilicon 1066 -736 1066 -736 0 1
rlabel polysilicon 1066 -742 1066 -742 0 3
rlabel polysilicon 1073 -736 1073 -736 0 1
rlabel polysilicon 1073 -742 1073 -742 0 3
rlabel polysilicon 1080 -736 1080 -736 0 1
rlabel polysilicon 1080 -742 1080 -742 0 3
rlabel polysilicon 1087 -736 1087 -736 0 1
rlabel polysilicon 1087 -742 1087 -742 0 3
rlabel polysilicon 1094 -736 1094 -736 0 1
rlabel polysilicon 1094 -742 1094 -742 0 3
rlabel polysilicon 1101 -736 1101 -736 0 1
rlabel polysilicon 1101 -742 1101 -742 0 3
rlabel polysilicon 1108 -736 1108 -736 0 1
rlabel polysilicon 1108 -742 1108 -742 0 3
rlabel polysilicon 1115 -736 1115 -736 0 1
rlabel polysilicon 1115 -742 1115 -742 0 3
rlabel polysilicon 1122 -736 1122 -736 0 1
rlabel polysilicon 1122 -742 1122 -742 0 3
rlabel polysilicon 1129 -736 1129 -736 0 1
rlabel polysilicon 1129 -742 1129 -742 0 3
rlabel polysilicon 1136 -736 1136 -736 0 1
rlabel polysilicon 1136 -742 1136 -742 0 3
rlabel polysilicon 1143 -736 1143 -736 0 1
rlabel polysilicon 1143 -742 1143 -742 0 3
rlabel polysilicon 1150 -736 1150 -736 0 1
rlabel polysilicon 1150 -742 1150 -742 0 3
rlabel polysilicon 1157 -736 1157 -736 0 1
rlabel polysilicon 1157 -742 1157 -742 0 3
rlabel polysilicon 1164 -736 1164 -736 0 1
rlabel polysilicon 1164 -742 1164 -742 0 3
rlabel polysilicon 1171 -736 1171 -736 0 1
rlabel polysilicon 1171 -742 1171 -742 0 3
rlabel polysilicon 1178 -736 1178 -736 0 1
rlabel polysilicon 1178 -742 1178 -742 0 3
rlabel polysilicon 1185 -736 1185 -736 0 1
rlabel polysilicon 1185 -742 1185 -742 0 3
rlabel polysilicon 1192 -736 1192 -736 0 1
rlabel polysilicon 1192 -742 1192 -742 0 3
rlabel polysilicon 1199 -736 1199 -736 0 1
rlabel polysilicon 1199 -742 1199 -742 0 3
rlabel polysilicon 1206 -736 1206 -736 0 1
rlabel polysilicon 1206 -742 1206 -742 0 3
rlabel polysilicon 1213 -736 1213 -736 0 1
rlabel polysilicon 1213 -742 1213 -742 0 3
rlabel polysilicon 1220 -736 1220 -736 0 1
rlabel polysilicon 1220 -742 1220 -742 0 3
rlabel polysilicon 1227 -736 1227 -736 0 1
rlabel polysilicon 1227 -742 1227 -742 0 3
rlabel polysilicon 1234 -736 1234 -736 0 1
rlabel polysilicon 1234 -742 1234 -742 0 3
rlabel polysilicon 1241 -736 1241 -736 0 1
rlabel polysilicon 1241 -742 1241 -742 0 3
rlabel polysilicon 1248 -736 1248 -736 0 1
rlabel polysilicon 1248 -742 1248 -742 0 3
rlabel polysilicon 1255 -736 1255 -736 0 1
rlabel polysilicon 1255 -742 1255 -742 0 3
rlabel polysilicon 1262 -736 1262 -736 0 1
rlabel polysilicon 1262 -742 1262 -742 0 3
rlabel polysilicon 1269 -736 1269 -736 0 1
rlabel polysilicon 1269 -742 1269 -742 0 3
rlabel polysilicon 1276 -736 1276 -736 0 1
rlabel polysilicon 1276 -742 1276 -742 0 3
rlabel polysilicon 1283 -736 1283 -736 0 1
rlabel polysilicon 1283 -742 1283 -742 0 3
rlabel polysilicon 1290 -736 1290 -736 0 1
rlabel polysilicon 1290 -742 1290 -742 0 3
rlabel polysilicon 1297 -736 1297 -736 0 1
rlabel polysilicon 1297 -742 1297 -742 0 3
rlabel polysilicon 1304 -736 1304 -736 0 1
rlabel polysilicon 1304 -742 1304 -742 0 3
rlabel polysilicon 1311 -736 1311 -736 0 1
rlabel polysilicon 1311 -742 1311 -742 0 3
rlabel polysilicon 1318 -736 1318 -736 0 1
rlabel polysilicon 1318 -742 1318 -742 0 3
rlabel polysilicon 1325 -736 1325 -736 0 1
rlabel polysilicon 1325 -742 1325 -742 0 3
rlabel polysilicon 1332 -736 1332 -736 0 1
rlabel polysilicon 1332 -742 1332 -742 0 3
rlabel polysilicon 1339 -736 1339 -736 0 1
rlabel polysilicon 1339 -742 1339 -742 0 3
rlabel polysilicon 1346 -736 1346 -736 0 1
rlabel polysilicon 1346 -742 1346 -742 0 3
rlabel polysilicon 1353 -736 1353 -736 0 1
rlabel polysilicon 1353 -742 1353 -742 0 3
rlabel polysilicon 1360 -736 1360 -736 0 1
rlabel polysilicon 1360 -742 1360 -742 0 3
rlabel polysilicon 1367 -736 1367 -736 0 1
rlabel polysilicon 1367 -742 1367 -742 0 3
rlabel polysilicon 1374 -736 1374 -736 0 1
rlabel polysilicon 1374 -742 1374 -742 0 3
rlabel polysilicon 1381 -736 1381 -736 0 1
rlabel polysilicon 1381 -742 1381 -742 0 3
rlabel polysilicon 1388 -736 1388 -736 0 1
rlabel polysilicon 1388 -742 1388 -742 0 3
rlabel polysilicon 1395 -736 1395 -736 0 1
rlabel polysilicon 1395 -742 1395 -742 0 3
rlabel polysilicon 1402 -736 1402 -736 0 1
rlabel polysilicon 1402 -742 1402 -742 0 3
rlabel polysilicon 1409 -736 1409 -736 0 1
rlabel polysilicon 1409 -742 1409 -742 0 3
rlabel polysilicon 1416 -736 1416 -736 0 1
rlabel polysilicon 1416 -742 1416 -742 0 3
rlabel polysilicon 1426 -736 1426 -736 0 2
rlabel polysilicon 1423 -742 1423 -742 0 3
rlabel polysilicon 1426 -742 1426 -742 0 4
rlabel polysilicon 1430 -736 1430 -736 0 1
rlabel polysilicon 1430 -742 1430 -742 0 3
rlabel polysilicon 1500 -736 1500 -736 0 1
rlabel polysilicon 1500 -742 1500 -742 0 3
rlabel polysilicon 1521 -736 1521 -736 0 1
rlabel polysilicon 1521 -742 1521 -742 0 3
rlabel polysilicon 1570 -736 1570 -736 0 1
rlabel polysilicon 1570 -742 1570 -742 0 3
rlabel polysilicon 1633 -736 1633 -736 0 1
rlabel polysilicon 1633 -742 1633 -742 0 3
rlabel polysilicon 23 -875 23 -875 0 1
rlabel polysilicon 23 -881 23 -881 0 3
rlabel polysilicon 33 -875 33 -875 0 2
rlabel polysilicon 37 -875 37 -875 0 1
rlabel polysilicon 37 -881 37 -881 0 3
rlabel polysilicon 44 -875 44 -875 0 1
rlabel polysilicon 44 -881 44 -881 0 3
rlabel polysilicon 51 -875 51 -875 0 1
rlabel polysilicon 54 -881 54 -881 0 4
rlabel polysilicon 58 -875 58 -875 0 1
rlabel polysilicon 58 -881 58 -881 0 3
rlabel polysilicon 65 -875 65 -875 0 1
rlabel polysilicon 65 -881 65 -881 0 3
rlabel polysilicon 72 -875 72 -875 0 1
rlabel polysilicon 72 -881 72 -881 0 3
rlabel polysilicon 79 -875 79 -875 0 1
rlabel polysilicon 79 -881 79 -881 0 3
rlabel polysilicon 86 -881 86 -881 0 3
rlabel polysilicon 89 -881 89 -881 0 4
rlabel polysilicon 93 -875 93 -875 0 1
rlabel polysilicon 93 -881 93 -881 0 3
rlabel polysilicon 100 -875 100 -875 0 1
rlabel polysilicon 103 -875 103 -875 0 2
rlabel polysilicon 100 -881 100 -881 0 3
rlabel polysilicon 103 -881 103 -881 0 4
rlabel polysilicon 107 -875 107 -875 0 1
rlabel polysilicon 110 -875 110 -875 0 2
rlabel polysilicon 107 -881 107 -881 0 3
rlabel polysilicon 114 -875 114 -875 0 1
rlabel polysilicon 114 -881 114 -881 0 3
rlabel polysilicon 121 -875 121 -875 0 1
rlabel polysilicon 121 -881 121 -881 0 3
rlabel polysilicon 128 -875 128 -875 0 1
rlabel polysilicon 128 -881 128 -881 0 3
rlabel polysilicon 135 -875 135 -875 0 1
rlabel polysilicon 138 -875 138 -875 0 2
rlabel polysilicon 135 -881 135 -881 0 3
rlabel polysilicon 138 -881 138 -881 0 4
rlabel polysilicon 142 -875 142 -875 0 1
rlabel polysilicon 142 -881 142 -881 0 3
rlabel polysilicon 149 -875 149 -875 0 1
rlabel polysilicon 149 -881 149 -881 0 3
rlabel polysilicon 156 -875 156 -875 0 1
rlabel polysilicon 156 -881 156 -881 0 3
rlabel polysilicon 166 -875 166 -875 0 2
rlabel polysilicon 163 -881 163 -881 0 3
rlabel polysilicon 166 -881 166 -881 0 4
rlabel polysilicon 170 -875 170 -875 0 1
rlabel polysilicon 170 -881 170 -881 0 3
rlabel polysilicon 177 -875 177 -875 0 1
rlabel polysilicon 177 -881 177 -881 0 3
rlabel polysilicon 184 -875 184 -875 0 1
rlabel polysilicon 184 -881 184 -881 0 3
rlabel polysilicon 191 -875 191 -875 0 1
rlabel polysilicon 191 -881 191 -881 0 3
rlabel polysilicon 198 -875 198 -875 0 1
rlabel polysilicon 198 -881 198 -881 0 3
rlabel polysilicon 205 -875 205 -875 0 1
rlabel polysilicon 208 -881 208 -881 0 4
rlabel polysilicon 212 -875 212 -875 0 1
rlabel polysilicon 212 -881 212 -881 0 3
rlabel polysilicon 219 -875 219 -875 0 1
rlabel polysilicon 219 -881 219 -881 0 3
rlabel polysilicon 229 -875 229 -875 0 2
rlabel polysilicon 226 -881 226 -881 0 3
rlabel polysilicon 229 -881 229 -881 0 4
rlabel polysilicon 233 -875 233 -875 0 1
rlabel polysilicon 236 -875 236 -875 0 2
rlabel polysilicon 233 -881 233 -881 0 3
rlabel polysilicon 236 -881 236 -881 0 4
rlabel polysilicon 240 -875 240 -875 0 1
rlabel polysilicon 240 -881 240 -881 0 3
rlabel polysilicon 247 -875 247 -875 0 1
rlabel polysilicon 250 -875 250 -875 0 2
rlabel polysilicon 250 -881 250 -881 0 4
rlabel polysilicon 254 -875 254 -875 0 1
rlabel polysilicon 254 -881 254 -881 0 3
rlabel polysilicon 261 -875 261 -875 0 1
rlabel polysilicon 261 -881 261 -881 0 3
rlabel polysilicon 268 -875 268 -875 0 1
rlabel polysilicon 268 -881 268 -881 0 3
rlabel polysilicon 275 -875 275 -875 0 1
rlabel polysilicon 275 -881 275 -881 0 3
rlabel polysilicon 282 -875 282 -875 0 1
rlabel polysilicon 282 -881 282 -881 0 3
rlabel polysilicon 289 -875 289 -875 0 1
rlabel polysilicon 289 -881 289 -881 0 3
rlabel polysilicon 303 -875 303 -875 0 1
rlabel polysilicon 303 -881 303 -881 0 3
rlabel polysilicon 310 -875 310 -875 0 1
rlabel polysilicon 310 -881 310 -881 0 3
rlabel polysilicon 324 -875 324 -875 0 1
rlabel polysilicon 324 -881 324 -881 0 3
rlabel polysilicon 331 -875 331 -875 0 1
rlabel polysilicon 331 -881 331 -881 0 3
rlabel polysilicon 338 -875 338 -875 0 1
rlabel polysilicon 338 -881 338 -881 0 3
rlabel polysilicon 345 -875 345 -875 0 1
rlabel polysilicon 345 -881 345 -881 0 3
rlabel polysilicon 352 -875 352 -875 0 1
rlabel polysilicon 352 -881 352 -881 0 3
rlabel polysilicon 359 -875 359 -875 0 1
rlabel polysilicon 359 -881 359 -881 0 3
rlabel polysilicon 366 -875 366 -875 0 1
rlabel polysilicon 366 -881 366 -881 0 3
rlabel polysilicon 373 -875 373 -875 0 1
rlabel polysilicon 373 -881 373 -881 0 3
rlabel polysilicon 380 -875 380 -875 0 1
rlabel polysilicon 380 -881 380 -881 0 3
rlabel polysilicon 387 -875 387 -875 0 1
rlabel polysilicon 387 -881 387 -881 0 3
rlabel polysilicon 394 -875 394 -875 0 1
rlabel polysilicon 394 -881 394 -881 0 3
rlabel polysilicon 401 -875 401 -875 0 1
rlabel polysilicon 401 -881 401 -881 0 3
rlabel polysilicon 408 -875 408 -875 0 1
rlabel polysilicon 408 -881 408 -881 0 3
rlabel polysilicon 415 -875 415 -875 0 1
rlabel polysilicon 415 -881 415 -881 0 3
rlabel polysilicon 422 -875 422 -875 0 1
rlabel polysilicon 422 -881 422 -881 0 3
rlabel polysilicon 429 -875 429 -875 0 1
rlabel polysilicon 429 -881 429 -881 0 3
rlabel polysilicon 436 -875 436 -875 0 1
rlabel polysilicon 436 -881 436 -881 0 3
rlabel polysilicon 443 -875 443 -875 0 1
rlabel polysilicon 443 -881 443 -881 0 3
rlabel polysilicon 450 -875 450 -875 0 1
rlabel polysilicon 450 -881 450 -881 0 3
rlabel polysilicon 457 -875 457 -875 0 1
rlabel polysilicon 457 -881 457 -881 0 3
rlabel polysilicon 464 -875 464 -875 0 1
rlabel polysilicon 467 -875 467 -875 0 2
rlabel polysilicon 467 -881 467 -881 0 4
rlabel polysilicon 471 -875 471 -875 0 1
rlabel polysilicon 471 -881 471 -881 0 3
rlabel polysilicon 478 -875 478 -875 0 1
rlabel polysilicon 478 -881 478 -881 0 3
rlabel polysilicon 481 -881 481 -881 0 4
rlabel polysilicon 485 -875 485 -875 0 1
rlabel polysilicon 485 -881 485 -881 0 3
rlabel polysilicon 492 -875 492 -875 0 1
rlabel polysilicon 492 -881 492 -881 0 3
rlabel polysilicon 499 -875 499 -875 0 1
rlabel polysilicon 499 -881 499 -881 0 3
rlabel polysilicon 506 -875 506 -875 0 1
rlabel polysilicon 506 -881 506 -881 0 3
rlabel polysilicon 513 -875 513 -875 0 1
rlabel polysilicon 513 -881 513 -881 0 3
rlabel polysilicon 520 -875 520 -875 0 1
rlabel polysilicon 520 -881 520 -881 0 3
rlabel polysilicon 527 -875 527 -875 0 1
rlabel polysilicon 527 -881 527 -881 0 3
rlabel polysilicon 534 -875 534 -875 0 1
rlabel polysilicon 534 -881 534 -881 0 3
rlabel polysilicon 541 -875 541 -875 0 1
rlabel polysilicon 541 -881 541 -881 0 3
rlabel polysilicon 548 -875 548 -875 0 1
rlabel polysilicon 548 -881 548 -881 0 3
rlabel polysilicon 555 -875 555 -875 0 1
rlabel polysilicon 555 -881 555 -881 0 3
rlabel polysilicon 562 -875 562 -875 0 1
rlabel polysilicon 565 -875 565 -875 0 2
rlabel polysilicon 562 -881 562 -881 0 3
rlabel polysilicon 569 -875 569 -875 0 1
rlabel polysilicon 569 -881 569 -881 0 3
rlabel polysilicon 576 -875 576 -875 0 1
rlabel polysilicon 576 -881 576 -881 0 3
rlabel polysilicon 579 -881 579 -881 0 4
rlabel polysilicon 583 -875 583 -875 0 1
rlabel polysilicon 586 -875 586 -875 0 2
rlabel polysilicon 583 -881 583 -881 0 3
rlabel polysilicon 586 -881 586 -881 0 4
rlabel polysilicon 590 -875 590 -875 0 1
rlabel polysilicon 590 -881 590 -881 0 3
rlabel polysilicon 597 -875 597 -875 0 1
rlabel polysilicon 597 -881 597 -881 0 3
rlabel polysilicon 604 -875 604 -875 0 1
rlabel polysilicon 604 -881 604 -881 0 3
rlabel polysilicon 611 -875 611 -875 0 1
rlabel polysilicon 611 -881 611 -881 0 3
rlabel polysilicon 614 -881 614 -881 0 4
rlabel polysilicon 618 -875 618 -875 0 1
rlabel polysilicon 618 -881 618 -881 0 3
rlabel polysilicon 625 -875 625 -875 0 1
rlabel polysilicon 628 -875 628 -875 0 2
rlabel polysilicon 625 -881 625 -881 0 3
rlabel polysilicon 628 -881 628 -881 0 4
rlabel polysilicon 632 -875 632 -875 0 1
rlabel polysilicon 632 -881 632 -881 0 3
rlabel polysilicon 639 -875 639 -875 0 1
rlabel polysilicon 642 -875 642 -875 0 2
rlabel polysilicon 639 -881 639 -881 0 3
rlabel polysilicon 646 -875 646 -875 0 1
rlabel polysilicon 646 -881 646 -881 0 3
rlabel polysilicon 660 -875 660 -875 0 1
rlabel polysilicon 660 -881 660 -881 0 3
rlabel polysilicon 663 -881 663 -881 0 4
rlabel polysilicon 667 -875 667 -875 0 1
rlabel polysilicon 667 -881 667 -881 0 3
rlabel polysilicon 674 -875 674 -875 0 1
rlabel polysilicon 674 -881 674 -881 0 3
rlabel polysilicon 681 -875 681 -875 0 1
rlabel polysilicon 681 -881 681 -881 0 3
rlabel polysilicon 688 -875 688 -875 0 1
rlabel polysilicon 691 -875 691 -875 0 2
rlabel polysilicon 691 -881 691 -881 0 4
rlabel polysilicon 695 -875 695 -875 0 1
rlabel polysilicon 695 -881 695 -881 0 3
rlabel polysilicon 702 -875 702 -875 0 1
rlabel polysilicon 705 -881 705 -881 0 4
rlabel polysilicon 709 -875 709 -875 0 1
rlabel polysilicon 709 -881 709 -881 0 3
rlabel polysilicon 716 -875 716 -875 0 1
rlabel polysilicon 716 -881 716 -881 0 3
rlabel polysilicon 723 -875 723 -875 0 1
rlabel polysilicon 723 -881 723 -881 0 3
rlabel polysilicon 730 -875 730 -875 0 1
rlabel polysilicon 730 -881 730 -881 0 3
rlabel polysilicon 737 -875 737 -875 0 1
rlabel polysilicon 740 -875 740 -875 0 2
rlabel polysilicon 737 -881 737 -881 0 3
rlabel polysilicon 740 -881 740 -881 0 4
rlabel polysilicon 744 -875 744 -875 0 1
rlabel polysilicon 744 -881 744 -881 0 3
rlabel polysilicon 751 -875 751 -875 0 1
rlabel polysilicon 751 -881 751 -881 0 3
rlabel polysilicon 758 -875 758 -875 0 1
rlabel polysilicon 758 -881 758 -881 0 3
rlabel polysilicon 761 -881 761 -881 0 4
rlabel polysilicon 765 -875 765 -875 0 1
rlabel polysilicon 765 -881 765 -881 0 3
rlabel polysilicon 772 -875 772 -875 0 1
rlabel polysilicon 772 -881 772 -881 0 3
rlabel polysilicon 782 -875 782 -875 0 2
rlabel polysilicon 779 -881 779 -881 0 3
rlabel polysilicon 786 -875 786 -875 0 1
rlabel polysilicon 789 -875 789 -875 0 2
rlabel polysilicon 786 -881 786 -881 0 3
rlabel polysilicon 789 -881 789 -881 0 4
rlabel polysilicon 793 -875 793 -875 0 1
rlabel polysilicon 793 -881 793 -881 0 3
rlabel polysilicon 796 -881 796 -881 0 4
rlabel polysilicon 800 -875 800 -875 0 1
rlabel polysilicon 800 -881 800 -881 0 3
rlabel polysilicon 807 -875 807 -875 0 1
rlabel polysilicon 807 -881 807 -881 0 3
rlabel polysilicon 814 -875 814 -875 0 1
rlabel polysilicon 814 -881 814 -881 0 3
rlabel polysilicon 821 -875 821 -875 0 1
rlabel polysilicon 821 -881 821 -881 0 3
rlabel polysilicon 828 -875 828 -875 0 1
rlabel polysilicon 831 -875 831 -875 0 2
rlabel polysilicon 828 -881 828 -881 0 3
rlabel polysilicon 835 -875 835 -875 0 1
rlabel polysilicon 835 -881 835 -881 0 3
rlabel polysilicon 842 -875 842 -875 0 1
rlabel polysilicon 842 -881 842 -881 0 3
rlabel polysilicon 849 -875 849 -875 0 1
rlabel polysilicon 849 -881 849 -881 0 3
rlabel polysilicon 856 -875 856 -875 0 1
rlabel polysilicon 856 -881 856 -881 0 3
rlabel polysilicon 863 -875 863 -875 0 1
rlabel polysilicon 863 -881 863 -881 0 3
rlabel polysilicon 870 -875 870 -875 0 1
rlabel polysilicon 870 -881 870 -881 0 3
rlabel polysilicon 877 -875 877 -875 0 1
rlabel polysilicon 877 -881 877 -881 0 3
rlabel polysilicon 880 -881 880 -881 0 4
rlabel polysilicon 884 -875 884 -875 0 1
rlabel polysilicon 884 -881 884 -881 0 3
rlabel polysilicon 891 -875 891 -875 0 1
rlabel polysilicon 891 -881 891 -881 0 3
rlabel polysilicon 898 -875 898 -875 0 1
rlabel polysilicon 898 -881 898 -881 0 3
rlabel polysilicon 905 -875 905 -875 0 1
rlabel polysilicon 908 -875 908 -875 0 2
rlabel polysilicon 905 -881 905 -881 0 3
rlabel polysilicon 908 -881 908 -881 0 4
rlabel polysilicon 912 -875 912 -875 0 1
rlabel polysilicon 912 -881 912 -881 0 3
rlabel polysilicon 919 -875 919 -875 0 1
rlabel polysilicon 919 -881 919 -881 0 3
rlabel polysilicon 929 -875 929 -875 0 2
rlabel polysilicon 926 -881 926 -881 0 3
rlabel polysilicon 929 -881 929 -881 0 4
rlabel polysilicon 933 -875 933 -875 0 1
rlabel polysilicon 933 -881 933 -881 0 3
rlabel polysilicon 940 -875 940 -875 0 1
rlabel polysilicon 940 -881 940 -881 0 3
rlabel polysilicon 947 -875 947 -875 0 1
rlabel polysilicon 947 -881 947 -881 0 3
rlabel polysilicon 954 -875 954 -875 0 1
rlabel polysilicon 954 -881 954 -881 0 3
rlabel polysilicon 961 -881 961 -881 0 3
rlabel polysilicon 964 -881 964 -881 0 4
rlabel polysilicon 968 -875 968 -875 0 1
rlabel polysilicon 968 -881 968 -881 0 3
rlabel polysilicon 975 -875 975 -875 0 1
rlabel polysilicon 975 -881 975 -881 0 3
rlabel polysilicon 982 -875 982 -875 0 1
rlabel polysilicon 982 -881 982 -881 0 3
rlabel polysilicon 989 -875 989 -875 0 1
rlabel polysilicon 989 -881 989 -881 0 3
rlabel polysilicon 996 -875 996 -875 0 1
rlabel polysilicon 996 -881 996 -881 0 3
rlabel polysilicon 1003 -875 1003 -875 0 1
rlabel polysilicon 1003 -881 1003 -881 0 3
rlabel polysilicon 1010 -875 1010 -875 0 1
rlabel polysilicon 1010 -881 1010 -881 0 3
rlabel polysilicon 1017 -875 1017 -875 0 1
rlabel polysilicon 1017 -881 1017 -881 0 3
rlabel polysilicon 1024 -875 1024 -875 0 1
rlabel polysilicon 1024 -881 1024 -881 0 3
rlabel polysilicon 1031 -875 1031 -875 0 1
rlabel polysilicon 1031 -881 1031 -881 0 3
rlabel polysilicon 1038 -875 1038 -875 0 1
rlabel polysilicon 1038 -881 1038 -881 0 3
rlabel polysilicon 1045 -875 1045 -875 0 1
rlabel polysilicon 1045 -881 1045 -881 0 3
rlabel polysilicon 1052 -875 1052 -875 0 1
rlabel polysilicon 1052 -881 1052 -881 0 3
rlabel polysilicon 1059 -875 1059 -875 0 1
rlabel polysilicon 1059 -881 1059 -881 0 3
rlabel polysilicon 1062 -881 1062 -881 0 4
rlabel polysilicon 1066 -875 1066 -875 0 1
rlabel polysilicon 1066 -881 1066 -881 0 3
rlabel polysilicon 1073 -875 1073 -875 0 1
rlabel polysilicon 1073 -881 1073 -881 0 3
rlabel polysilicon 1080 -875 1080 -875 0 1
rlabel polysilicon 1080 -881 1080 -881 0 3
rlabel polysilicon 1087 -875 1087 -875 0 1
rlabel polysilicon 1087 -881 1087 -881 0 3
rlabel polysilicon 1094 -875 1094 -875 0 1
rlabel polysilicon 1094 -881 1094 -881 0 3
rlabel polysilicon 1101 -875 1101 -875 0 1
rlabel polysilicon 1101 -881 1101 -881 0 3
rlabel polysilicon 1108 -875 1108 -875 0 1
rlabel polysilicon 1108 -881 1108 -881 0 3
rlabel polysilicon 1115 -875 1115 -875 0 1
rlabel polysilicon 1115 -881 1115 -881 0 3
rlabel polysilicon 1122 -875 1122 -875 0 1
rlabel polysilicon 1122 -881 1122 -881 0 3
rlabel polysilicon 1129 -875 1129 -875 0 1
rlabel polysilicon 1129 -881 1129 -881 0 3
rlabel polysilicon 1136 -875 1136 -875 0 1
rlabel polysilicon 1136 -881 1136 -881 0 3
rlabel polysilicon 1143 -875 1143 -875 0 1
rlabel polysilicon 1143 -881 1143 -881 0 3
rlabel polysilicon 1150 -875 1150 -875 0 1
rlabel polysilicon 1150 -881 1150 -881 0 3
rlabel polysilicon 1157 -875 1157 -875 0 1
rlabel polysilicon 1157 -881 1157 -881 0 3
rlabel polysilicon 1164 -875 1164 -875 0 1
rlabel polysilicon 1164 -881 1164 -881 0 3
rlabel polysilicon 1171 -875 1171 -875 0 1
rlabel polysilicon 1171 -881 1171 -881 0 3
rlabel polysilicon 1178 -875 1178 -875 0 1
rlabel polysilicon 1178 -881 1178 -881 0 3
rlabel polysilicon 1185 -875 1185 -875 0 1
rlabel polysilicon 1185 -881 1185 -881 0 3
rlabel polysilicon 1192 -875 1192 -875 0 1
rlabel polysilicon 1192 -881 1192 -881 0 3
rlabel polysilicon 1199 -875 1199 -875 0 1
rlabel polysilicon 1199 -881 1199 -881 0 3
rlabel polysilicon 1206 -875 1206 -875 0 1
rlabel polysilicon 1206 -881 1206 -881 0 3
rlabel polysilicon 1213 -875 1213 -875 0 1
rlabel polysilicon 1213 -881 1213 -881 0 3
rlabel polysilicon 1220 -875 1220 -875 0 1
rlabel polysilicon 1220 -881 1220 -881 0 3
rlabel polysilicon 1227 -875 1227 -875 0 1
rlabel polysilicon 1227 -881 1227 -881 0 3
rlabel polysilicon 1234 -875 1234 -875 0 1
rlabel polysilicon 1234 -881 1234 -881 0 3
rlabel polysilicon 1241 -875 1241 -875 0 1
rlabel polysilicon 1241 -881 1241 -881 0 3
rlabel polysilicon 1248 -875 1248 -875 0 1
rlabel polysilicon 1248 -881 1248 -881 0 3
rlabel polysilicon 1255 -875 1255 -875 0 1
rlabel polysilicon 1255 -881 1255 -881 0 3
rlabel polysilicon 1262 -875 1262 -875 0 1
rlabel polysilicon 1262 -881 1262 -881 0 3
rlabel polysilicon 1269 -875 1269 -875 0 1
rlabel polysilicon 1269 -881 1269 -881 0 3
rlabel polysilicon 1276 -875 1276 -875 0 1
rlabel polysilicon 1276 -881 1276 -881 0 3
rlabel polysilicon 1283 -875 1283 -875 0 1
rlabel polysilicon 1283 -881 1283 -881 0 3
rlabel polysilicon 1290 -875 1290 -875 0 1
rlabel polysilicon 1290 -881 1290 -881 0 3
rlabel polysilicon 1297 -875 1297 -875 0 1
rlabel polysilicon 1297 -881 1297 -881 0 3
rlabel polysilicon 1304 -875 1304 -875 0 1
rlabel polysilicon 1304 -881 1304 -881 0 3
rlabel polysilicon 1311 -875 1311 -875 0 1
rlabel polysilicon 1311 -881 1311 -881 0 3
rlabel polysilicon 1318 -875 1318 -875 0 1
rlabel polysilicon 1318 -881 1318 -881 0 3
rlabel polysilicon 1325 -875 1325 -875 0 1
rlabel polysilicon 1325 -881 1325 -881 0 3
rlabel polysilicon 1332 -875 1332 -875 0 1
rlabel polysilicon 1332 -881 1332 -881 0 3
rlabel polysilicon 1339 -875 1339 -875 0 1
rlabel polysilicon 1339 -881 1339 -881 0 3
rlabel polysilicon 1346 -875 1346 -875 0 1
rlabel polysilicon 1346 -881 1346 -881 0 3
rlabel polysilicon 1353 -875 1353 -875 0 1
rlabel polysilicon 1353 -881 1353 -881 0 3
rlabel polysilicon 1360 -875 1360 -875 0 1
rlabel polysilicon 1360 -881 1360 -881 0 3
rlabel polysilicon 1367 -875 1367 -875 0 1
rlabel polysilicon 1367 -881 1367 -881 0 3
rlabel polysilicon 1374 -875 1374 -875 0 1
rlabel polysilicon 1374 -881 1374 -881 0 3
rlabel polysilicon 1381 -875 1381 -875 0 1
rlabel polysilicon 1381 -881 1381 -881 0 3
rlabel polysilicon 1388 -875 1388 -875 0 1
rlabel polysilicon 1388 -881 1388 -881 0 3
rlabel polysilicon 1395 -875 1395 -875 0 1
rlabel polysilicon 1395 -881 1395 -881 0 3
rlabel polysilicon 1402 -875 1402 -875 0 1
rlabel polysilicon 1402 -881 1402 -881 0 3
rlabel polysilicon 1409 -875 1409 -875 0 1
rlabel polysilicon 1409 -881 1409 -881 0 3
rlabel polysilicon 1416 -875 1416 -875 0 1
rlabel polysilicon 1416 -881 1416 -881 0 3
rlabel polysilicon 1423 -875 1423 -875 0 1
rlabel polysilicon 1423 -881 1423 -881 0 3
rlabel polysilicon 1430 -875 1430 -875 0 1
rlabel polysilicon 1430 -881 1430 -881 0 3
rlabel polysilicon 1437 -875 1437 -875 0 1
rlabel polysilicon 1437 -881 1437 -881 0 3
rlabel polysilicon 1444 -875 1444 -875 0 1
rlabel polysilicon 1444 -881 1444 -881 0 3
rlabel polysilicon 1451 -875 1451 -875 0 1
rlabel polysilicon 1451 -881 1451 -881 0 3
rlabel polysilicon 1458 -875 1458 -875 0 1
rlabel polysilicon 1458 -881 1458 -881 0 3
rlabel polysilicon 1465 -875 1465 -875 0 1
rlabel polysilicon 1465 -881 1465 -881 0 3
rlabel polysilicon 1472 -875 1472 -875 0 1
rlabel polysilicon 1472 -881 1472 -881 0 3
rlabel polysilicon 1479 -875 1479 -875 0 1
rlabel polysilicon 1479 -881 1479 -881 0 3
rlabel polysilicon 1486 -875 1486 -875 0 1
rlabel polysilicon 1486 -881 1486 -881 0 3
rlabel polysilicon 1493 -875 1493 -875 0 1
rlabel polysilicon 1493 -881 1493 -881 0 3
rlabel polysilicon 1500 -875 1500 -875 0 1
rlabel polysilicon 1500 -881 1500 -881 0 3
rlabel polysilicon 1507 -875 1507 -875 0 1
rlabel polysilicon 1507 -881 1507 -881 0 3
rlabel polysilicon 1514 -875 1514 -875 0 1
rlabel polysilicon 1514 -881 1514 -881 0 3
rlabel polysilicon 1521 -875 1521 -875 0 1
rlabel polysilicon 1521 -881 1521 -881 0 3
rlabel polysilicon 1528 -875 1528 -875 0 1
rlabel polysilicon 1528 -881 1528 -881 0 3
rlabel polysilicon 1535 -875 1535 -875 0 1
rlabel polysilicon 1535 -881 1535 -881 0 3
rlabel polysilicon 1542 -875 1542 -875 0 1
rlabel polysilicon 1542 -881 1542 -881 0 3
rlabel polysilicon 1549 -875 1549 -875 0 1
rlabel polysilicon 1549 -881 1549 -881 0 3
rlabel polysilicon 1556 -875 1556 -875 0 1
rlabel polysilicon 1556 -881 1556 -881 0 3
rlabel polysilicon 1563 -875 1563 -875 0 1
rlabel polysilicon 1563 -881 1563 -881 0 3
rlabel polysilicon 1570 -875 1570 -875 0 1
rlabel polysilicon 1570 -881 1570 -881 0 3
rlabel polysilicon 1577 -875 1577 -875 0 1
rlabel polysilicon 1577 -881 1577 -881 0 3
rlabel polysilicon 1584 -875 1584 -875 0 1
rlabel polysilicon 1584 -881 1584 -881 0 3
rlabel polysilicon 1591 -875 1591 -875 0 1
rlabel polysilicon 1591 -881 1591 -881 0 3
rlabel polysilicon 1601 -881 1601 -881 0 4
rlabel polysilicon 1605 -875 1605 -875 0 1
rlabel polysilicon 1608 -875 1608 -875 0 2
rlabel polysilicon 1608 -881 1608 -881 0 4
rlabel polysilicon 1612 -875 1612 -875 0 1
rlabel polysilicon 1612 -881 1612 -881 0 3
rlabel polysilicon 1619 -875 1619 -875 0 1
rlabel polysilicon 1619 -881 1619 -881 0 3
rlabel polysilicon 1626 -875 1626 -875 0 1
rlabel polysilicon 1626 -881 1626 -881 0 3
rlabel polysilicon 1633 -875 1633 -875 0 1
rlabel polysilicon 1633 -881 1633 -881 0 3
rlabel polysilicon 1696 -875 1696 -875 0 1
rlabel polysilicon 1696 -881 1696 -881 0 3
rlabel polysilicon 30 -1036 30 -1036 0 1
rlabel polysilicon 30 -1042 30 -1042 0 3
rlabel polysilicon 37 -1036 37 -1036 0 1
rlabel polysilicon 37 -1042 37 -1042 0 3
rlabel polysilicon 44 -1036 44 -1036 0 1
rlabel polysilicon 47 -1042 47 -1042 0 4
rlabel polysilicon 54 -1036 54 -1036 0 2
rlabel polysilicon 51 -1042 51 -1042 0 3
rlabel polysilicon 54 -1042 54 -1042 0 4
rlabel polysilicon 58 -1036 58 -1036 0 1
rlabel polysilicon 58 -1042 58 -1042 0 3
rlabel polysilicon 65 -1036 65 -1036 0 1
rlabel polysilicon 65 -1042 65 -1042 0 3
rlabel polysilicon 72 -1036 72 -1036 0 1
rlabel polysilicon 72 -1042 72 -1042 0 3
rlabel polysilicon 79 -1036 79 -1036 0 1
rlabel polysilicon 79 -1042 79 -1042 0 3
rlabel polysilicon 86 -1036 86 -1036 0 1
rlabel polysilicon 89 -1036 89 -1036 0 2
rlabel polysilicon 86 -1042 86 -1042 0 3
rlabel polysilicon 89 -1042 89 -1042 0 4
rlabel polysilicon 93 -1036 93 -1036 0 1
rlabel polysilicon 93 -1042 93 -1042 0 3
rlabel polysilicon 100 -1036 100 -1036 0 1
rlabel polysilicon 100 -1042 100 -1042 0 3
rlabel polysilicon 107 -1036 107 -1036 0 1
rlabel polysilicon 110 -1036 110 -1036 0 2
rlabel polysilicon 107 -1042 107 -1042 0 3
rlabel polysilicon 110 -1042 110 -1042 0 4
rlabel polysilicon 114 -1036 114 -1036 0 1
rlabel polysilicon 114 -1042 114 -1042 0 3
rlabel polysilicon 121 -1036 121 -1036 0 1
rlabel polysilicon 124 -1036 124 -1036 0 2
rlabel polysilicon 121 -1042 121 -1042 0 3
rlabel polysilicon 128 -1036 128 -1036 0 1
rlabel polysilicon 128 -1042 128 -1042 0 3
rlabel polysilicon 135 -1036 135 -1036 0 1
rlabel polysilicon 135 -1042 135 -1042 0 3
rlabel polysilicon 142 -1036 142 -1036 0 1
rlabel polysilicon 142 -1042 142 -1042 0 3
rlabel polysilicon 149 -1036 149 -1036 0 1
rlabel polysilicon 149 -1042 149 -1042 0 3
rlabel polysilicon 156 -1036 156 -1036 0 1
rlabel polysilicon 156 -1042 156 -1042 0 3
rlabel polysilicon 163 -1036 163 -1036 0 1
rlabel polysilicon 163 -1042 163 -1042 0 3
rlabel polysilicon 170 -1036 170 -1036 0 1
rlabel polysilicon 170 -1042 170 -1042 0 3
rlabel polysilicon 177 -1036 177 -1036 0 1
rlabel polysilicon 177 -1042 177 -1042 0 3
rlabel polysilicon 184 -1036 184 -1036 0 1
rlabel polysilicon 184 -1042 184 -1042 0 3
rlabel polysilicon 191 -1036 191 -1036 0 1
rlabel polysilicon 191 -1042 191 -1042 0 3
rlabel polysilicon 198 -1036 198 -1036 0 1
rlabel polysilicon 201 -1036 201 -1036 0 2
rlabel polysilicon 198 -1042 198 -1042 0 3
rlabel polysilicon 201 -1042 201 -1042 0 4
rlabel polysilicon 205 -1036 205 -1036 0 1
rlabel polysilicon 205 -1042 205 -1042 0 3
rlabel polysilicon 212 -1036 212 -1036 0 1
rlabel polysilicon 212 -1042 212 -1042 0 3
rlabel polysilicon 226 -1036 226 -1036 0 1
rlabel polysilicon 226 -1042 226 -1042 0 3
rlabel polysilicon 233 -1036 233 -1036 0 1
rlabel polysilicon 233 -1042 233 -1042 0 3
rlabel polysilicon 240 -1036 240 -1036 0 1
rlabel polysilicon 240 -1042 240 -1042 0 3
rlabel polysilicon 247 -1036 247 -1036 0 1
rlabel polysilicon 247 -1042 247 -1042 0 3
rlabel polysilicon 254 -1036 254 -1036 0 1
rlabel polysilicon 254 -1042 254 -1042 0 3
rlabel polysilicon 261 -1036 261 -1036 0 1
rlabel polysilicon 261 -1042 261 -1042 0 3
rlabel polysilicon 268 -1036 268 -1036 0 1
rlabel polysilicon 268 -1042 268 -1042 0 3
rlabel polysilicon 275 -1036 275 -1036 0 1
rlabel polysilicon 275 -1042 275 -1042 0 3
rlabel polysilicon 282 -1036 282 -1036 0 1
rlabel polysilicon 282 -1042 282 -1042 0 3
rlabel polysilicon 289 -1036 289 -1036 0 1
rlabel polysilicon 292 -1036 292 -1036 0 2
rlabel polysilicon 289 -1042 289 -1042 0 3
rlabel polysilicon 292 -1042 292 -1042 0 4
rlabel polysilicon 296 -1036 296 -1036 0 1
rlabel polysilicon 296 -1042 296 -1042 0 3
rlabel polysilicon 303 -1036 303 -1036 0 1
rlabel polysilicon 303 -1042 303 -1042 0 3
rlabel polysilicon 313 -1036 313 -1036 0 2
rlabel polysilicon 317 -1036 317 -1036 0 1
rlabel polysilicon 317 -1042 317 -1042 0 3
rlabel polysilicon 324 -1036 324 -1036 0 1
rlabel polysilicon 324 -1042 324 -1042 0 3
rlabel polysilicon 331 -1036 331 -1036 0 1
rlabel polysilicon 331 -1042 331 -1042 0 3
rlabel polysilicon 338 -1036 338 -1036 0 1
rlabel polysilicon 338 -1042 338 -1042 0 3
rlabel polysilicon 345 -1036 345 -1036 0 1
rlabel polysilicon 345 -1042 345 -1042 0 3
rlabel polysilicon 352 -1036 352 -1036 0 1
rlabel polysilicon 352 -1042 352 -1042 0 3
rlabel polysilicon 359 -1036 359 -1036 0 1
rlabel polysilicon 359 -1042 359 -1042 0 3
rlabel polysilicon 366 -1036 366 -1036 0 1
rlabel polysilicon 366 -1042 366 -1042 0 3
rlabel polysilicon 373 -1036 373 -1036 0 1
rlabel polysilicon 373 -1042 373 -1042 0 3
rlabel polysilicon 380 -1036 380 -1036 0 1
rlabel polysilicon 380 -1042 380 -1042 0 3
rlabel polysilicon 387 -1036 387 -1036 0 1
rlabel polysilicon 387 -1042 387 -1042 0 3
rlabel polysilicon 394 -1036 394 -1036 0 1
rlabel polysilicon 394 -1042 394 -1042 0 3
rlabel polysilicon 401 -1036 401 -1036 0 1
rlabel polysilicon 401 -1042 401 -1042 0 3
rlabel polysilicon 408 -1036 408 -1036 0 1
rlabel polysilicon 408 -1042 408 -1042 0 3
rlabel polysilicon 415 -1036 415 -1036 0 1
rlabel polysilicon 415 -1042 415 -1042 0 3
rlabel polysilicon 422 -1036 422 -1036 0 1
rlabel polysilicon 422 -1042 422 -1042 0 3
rlabel polysilicon 429 -1036 429 -1036 0 1
rlabel polysilicon 429 -1042 429 -1042 0 3
rlabel polysilicon 436 -1036 436 -1036 0 1
rlabel polysilicon 436 -1042 436 -1042 0 3
rlabel polysilicon 443 -1036 443 -1036 0 1
rlabel polysilicon 443 -1042 443 -1042 0 3
rlabel polysilicon 450 -1036 450 -1036 0 1
rlabel polysilicon 450 -1042 450 -1042 0 3
rlabel polysilicon 457 -1036 457 -1036 0 1
rlabel polysilicon 457 -1042 457 -1042 0 3
rlabel polysilicon 467 -1036 467 -1036 0 2
rlabel polysilicon 467 -1042 467 -1042 0 4
rlabel polysilicon 471 -1036 471 -1036 0 1
rlabel polysilicon 474 -1036 474 -1036 0 2
rlabel polysilicon 471 -1042 471 -1042 0 3
rlabel polysilicon 474 -1042 474 -1042 0 4
rlabel polysilicon 478 -1036 478 -1036 0 1
rlabel polysilicon 478 -1042 478 -1042 0 3
rlabel polysilicon 485 -1036 485 -1036 0 1
rlabel polysilicon 485 -1042 485 -1042 0 3
rlabel polysilicon 492 -1036 492 -1036 0 1
rlabel polysilicon 492 -1042 492 -1042 0 3
rlabel polysilicon 499 -1036 499 -1036 0 1
rlabel polysilicon 499 -1042 499 -1042 0 3
rlabel polysilicon 506 -1036 506 -1036 0 1
rlabel polysilicon 506 -1042 506 -1042 0 3
rlabel polysilicon 513 -1036 513 -1036 0 1
rlabel polysilicon 513 -1042 513 -1042 0 3
rlabel polysilicon 520 -1036 520 -1036 0 1
rlabel polysilicon 520 -1042 520 -1042 0 3
rlabel polysilicon 527 -1036 527 -1036 0 1
rlabel polysilicon 527 -1042 527 -1042 0 3
rlabel polysilicon 534 -1036 534 -1036 0 1
rlabel polysilicon 537 -1036 537 -1036 0 2
rlabel polysilicon 534 -1042 534 -1042 0 3
rlabel polysilicon 537 -1042 537 -1042 0 4
rlabel polysilicon 541 -1036 541 -1036 0 1
rlabel polysilicon 541 -1042 541 -1042 0 3
rlabel polysilicon 548 -1036 548 -1036 0 1
rlabel polysilicon 551 -1036 551 -1036 0 2
rlabel polysilicon 548 -1042 548 -1042 0 3
rlabel polysilicon 551 -1042 551 -1042 0 4
rlabel polysilicon 555 -1036 555 -1036 0 1
rlabel polysilicon 555 -1042 555 -1042 0 3
rlabel polysilicon 562 -1036 562 -1036 0 1
rlabel polysilicon 562 -1042 562 -1042 0 3
rlabel polysilicon 569 -1036 569 -1036 0 1
rlabel polysilicon 569 -1042 569 -1042 0 3
rlabel polysilicon 576 -1036 576 -1036 0 1
rlabel polysilicon 576 -1042 576 -1042 0 3
rlabel polysilicon 583 -1036 583 -1036 0 1
rlabel polysilicon 583 -1042 583 -1042 0 3
rlabel polysilicon 593 -1036 593 -1036 0 2
rlabel polysilicon 590 -1042 590 -1042 0 3
rlabel polysilicon 593 -1042 593 -1042 0 4
rlabel polysilicon 597 -1036 597 -1036 0 1
rlabel polysilicon 600 -1036 600 -1036 0 2
rlabel polysilicon 597 -1042 597 -1042 0 3
rlabel polysilicon 600 -1042 600 -1042 0 4
rlabel polysilicon 604 -1036 604 -1036 0 1
rlabel polysilicon 607 -1036 607 -1036 0 2
rlabel polysilicon 604 -1042 604 -1042 0 3
rlabel polysilicon 607 -1042 607 -1042 0 4
rlabel polysilicon 611 -1036 611 -1036 0 1
rlabel polysilicon 611 -1042 611 -1042 0 3
rlabel polysilicon 618 -1036 618 -1036 0 1
rlabel polysilicon 621 -1036 621 -1036 0 2
rlabel polysilicon 621 -1042 621 -1042 0 4
rlabel polysilicon 625 -1036 625 -1036 0 1
rlabel polysilicon 625 -1042 625 -1042 0 3
rlabel polysilicon 628 -1042 628 -1042 0 4
rlabel polysilicon 632 -1036 632 -1036 0 1
rlabel polysilicon 635 -1036 635 -1036 0 2
rlabel polysilicon 632 -1042 632 -1042 0 3
rlabel polysilicon 635 -1042 635 -1042 0 4
rlabel polysilicon 639 -1036 639 -1036 0 1
rlabel polysilicon 639 -1042 639 -1042 0 3
rlabel polysilicon 646 -1036 646 -1036 0 1
rlabel polysilicon 646 -1042 646 -1042 0 3
rlabel polysilicon 653 -1036 653 -1036 0 1
rlabel polysilicon 653 -1042 653 -1042 0 3
rlabel polysilicon 660 -1036 660 -1036 0 1
rlabel polysilicon 660 -1042 660 -1042 0 3
rlabel polysilicon 667 -1036 667 -1036 0 1
rlabel polysilicon 667 -1042 667 -1042 0 3
rlabel polysilicon 674 -1036 674 -1036 0 1
rlabel polysilicon 674 -1042 674 -1042 0 3
rlabel polysilicon 681 -1036 681 -1036 0 1
rlabel polysilicon 681 -1042 681 -1042 0 3
rlabel polysilicon 688 -1036 688 -1036 0 1
rlabel polysilicon 688 -1042 688 -1042 0 3
rlabel polysilicon 695 -1036 695 -1036 0 1
rlabel polysilicon 695 -1042 695 -1042 0 3
rlabel polysilicon 702 -1036 702 -1036 0 1
rlabel polysilicon 702 -1042 702 -1042 0 3
rlabel polysilicon 709 -1036 709 -1036 0 1
rlabel polysilicon 709 -1042 709 -1042 0 3
rlabel polysilicon 716 -1036 716 -1036 0 1
rlabel polysilicon 716 -1042 716 -1042 0 3
rlabel polysilicon 723 -1036 723 -1036 0 1
rlabel polysilicon 723 -1042 723 -1042 0 3
rlabel polysilicon 726 -1042 726 -1042 0 4
rlabel polysilicon 730 -1036 730 -1036 0 1
rlabel polysilicon 733 -1036 733 -1036 0 2
rlabel polysilicon 730 -1042 730 -1042 0 3
rlabel polysilicon 733 -1042 733 -1042 0 4
rlabel polysilicon 737 -1036 737 -1036 0 1
rlabel polysilicon 737 -1042 737 -1042 0 3
rlabel polysilicon 744 -1036 744 -1036 0 1
rlabel polysilicon 744 -1042 744 -1042 0 3
rlabel polysilicon 751 -1036 751 -1036 0 1
rlabel polysilicon 751 -1042 751 -1042 0 3
rlabel polysilicon 761 -1036 761 -1036 0 2
rlabel polysilicon 758 -1042 758 -1042 0 3
rlabel polysilicon 761 -1042 761 -1042 0 4
rlabel polysilicon 765 -1036 765 -1036 0 1
rlabel polysilicon 768 -1036 768 -1036 0 2
rlabel polysilicon 765 -1042 765 -1042 0 3
rlabel polysilicon 768 -1042 768 -1042 0 4
rlabel polysilicon 772 -1036 772 -1036 0 1
rlabel polysilicon 772 -1042 772 -1042 0 3
rlabel polysilicon 779 -1036 779 -1036 0 1
rlabel polysilicon 779 -1042 779 -1042 0 3
rlabel polysilicon 786 -1036 786 -1036 0 1
rlabel polysilicon 786 -1042 786 -1042 0 3
rlabel polysilicon 793 -1036 793 -1036 0 1
rlabel polysilicon 796 -1036 796 -1036 0 2
rlabel polysilicon 793 -1042 793 -1042 0 3
rlabel polysilicon 800 -1036 800 -1036 0 1
rlabel polysilicon 800 -1042 800 -1042 0 3
rlabel polysilicon 807 -1036 807 -1036 0 1
rlabel polysilicon 810 -1036 810 -1036 0 2
rlabel polysilicon 807 -1042 807 -1042 0 3
rlabel polysilicon 810 -1042 810 -1042 0 4
rlabel polysilicon 814 -1036 814 -1036 0 1
rlabel polysilicon 814 -1042 814 -1042 0 3
rlabel polysilicon 821 -1036 821 -1036 0 1
rlabel polysilicon 821 -1042 821 -1042 0 3
rlabel polysilicon 828 -1036 828 -1036 0 1
rlabel polysilicon 831 -1042 831 -1042 0 4
rlabel polysilicon 835 -1036 835 -1036 0 1
rlabel polysilicon 835 -1042 835 -1042 0 3
rlabel polysilicon 842 -1036 842 -1036 0 1
rlabel polysilicon 845 -1036 845 -1036 0 2
rlabel polysilicon 842 -1042 842 -1042 0 3
rlabel polysilicon 845 -1042 845 -1042 0 4
rlabel polysilicon 849 -1036 849 -1036 0 1
rlabel polysilicon 849 -1042 849 -1042 0 3
rlabel polysilicon 856 -1036 856 -1036 0 1
rlabel polysilicon 856 -1042 856 -1042 0 3
rlabel polysilicon 859 -1042 859 -1042 0 4
rlabel polysilicon 863 -1036 863 -1036 0 1
rlabel polysilicon 863 -1042 863 -1042 0 3
rlabel polysilicon 870 -1036 870 -1036 0 1
rlabel polysilicon 873 -1036 873 -1036 0 2
rlabel polysilicon 870 -1042 870 -1042 0 3
rlabel polysilicon 873 -1042 873 -1042 0 4
rlabel polysilicon 877 -1036 877 -1036 0 1
rlabel polysilicon 880 -1036 880 -1036 0 2
rlabel polysilicon 877 -1042 877 -1042 0 3
rlabel polysilicon 880 -1042 880 -1042 0 4
rlabel polysilicon 884 -1036 884 -1036 0 1
rlabel polysilicon 884 -1042 884 -1042 0 3
rlabel polysilicon 891 -1036 891 -1036 0 1
rlabel polysilicon 891 -1042 891 -1042 0 3
rlabel polysilicon 898 -1036 898 -1036 0 1
rlabel polysilicon 901 -1036 901 -1036 0 2
rlabel polysilicon 898 -1042 898 -1042 0 3
rlabel polysilicon 905 -1036 905 -1036 0 1
rlabel polysilicon 905 -1042 905 -1042 0 3
rlabel polysilicon 912 -1036 912 -1036 0 1
rlabel polysilicon 912 -1042 912 -1042 0 3
rlabel polysilicon 919 -1036 919 -1036 0 1
rlabel polysilicon 919 -1042 919 -1042 0 3
rlabel polysilicon 926 -1036 926 -1036 0 1
rlabel polysilicon 926 -1042 926 -1042 0 3
rlabel polysilicon 933 -1036 933 -1036 0 1
rlabel polysilicon 933 -1042 933 -1042 0 3
rlabel polysilicon 940 -1036 940 -1036 0 1
rlabel polysilicon 940 -1042 940 -1042 0 3
rlabel polysilicon 947 -1036 947 -1036 0 1
rlabel polysilicon 947 -1042 947 -1042 0 3
rlabel polysilicon 954 -1036 954 -1036 0 1
rlabel polysilicon 957 -1036 957 -1036 0 2
rlabel polysilicon 954 -1042 954 -1042 0 3
rlabel polysilicon 957 -1042 957 -1042 0 4
rlabel polysilicon 961 -1036 961 -1036 0 1
rlabel polysilicon 961 -1042 961 -1042 0 3
rlabel polysilicon 968 -1036 968 -1036 0 1
rlabel polysilicon 968 -1042 968 -1042 0 3
rlabel polysilicon 975 -1036 975 -1036 0 1
rlabel polysilicon 978 -1036 978 -1036 0 2
rlabel polysilicon 978 -1042 978 -1042 0 4
rlabel polysilicon 982 -1036 982 -1036 0 1
rlabel polysilicon 982 -1042 982 -1042 0 3
rlabel polysilicon 989 -1036 989 -1036 0 1
rlabel polysilicon 992 -1036 992 -1036 0 2
rlabel polysilicon 989 -1042 989 -1042 0 3
rlabel polysilicon 992 -1042 992 -1042 0 4
rlabel polysilicon 996 -1036 996 -1036 0 1
rlabel polysilicon 996 -1042 996 -1042 0 3
rlabel polysilicon 1003 -1036 1003 -1036 0 1
rlabel polysilicon 1003 -1042 1003 -1042 0 3
rlabel polysilicon 1010 -1036 1010 -1036 0 1
rlabel polysilicon 1010 -1042 1010 -1042 0 3
rlabel polysilicon 1017 -1036 1017 -1036 0 1
rlabel polysilicon 1017 -1042 1017 -1042 0 3
rlabel polysilicon 1024 -1036 1024 -1036 0 1
rlabel polysilicon 1024 -1042 1024 -1042 0 3
rlabel polysilicon 1031 -1036 1031 -1036 0 1
rlabel polysilicon 1031 -1042 1031 -1042 0 3
rlabel polysilicon 1038 -1036 1038 -1036 0 1
rlabel polysilicon 1038 -1042 1038 -1042 0 3
rlabel polysilicon 1045 -1036 1045 -1036 0 1
rlabel polysilicon 1045 -1042 1045 -1042 0 3
rlabel polysilicon 1052 -1036 1052 -1036 0 1
rlabel polysilicon 1052 -1042 1052 -1042 0 3
rlabel polysilicon 1062 -1036 1062 -1036 0 2
rlabel polysilicon 1062 -1042 1062 -1042 0 4
rlabel polysilicon 1066 -1036 1066 -1036 0 1
rlabel polysilicon 1066 -1042 1066 -1042 0 3
rlabel polysilicon 1069 -1042 1069 -1042 0 4
rlabel polysilicon 1073 -1036 1073 -1036 0 1
rlabel polysilicon 1073 -1042 1073 -1042 0 3
rlabel polysilicon 1080 -1036 1080 -1036 0 1
rlabel polysilicon 1080 -1042 1080 -1042 0 3
rlabel polysilicon 1087 -1036 1087 -1036 0 1
rlabel polysilicon 1087 -1042 1087 -1042 0 3
rlabel polysilicon 1094 -1036 1094 -1036 0 1
rlabel polysilicon 1094 -1042 1094 -1042 0 3
rlabel polysilicon 1101 -1036 1101 -1036 0 1
rlabel polysilicon 1101 -1042 1101 -1042 0 3
rlabel polysilicon 1108 -1036 1108 -1036 0 1
rlabel polysilicon 1108 -1042 1108 -1042 0 3
rlabel polysilicon 1115 -1036 1115 -1036 0 1
rlabel polysilicon 1115 -1042 1115 -1042 0 3
rlabel polysilicon 1122 -1036 1122 -1036 0 1
rlabel polysilicon 1122 -1042 1122 -1042 0 3
rlabel polysilicon 1129 -1036 1129 -1036 0 1
rlabel polysilicon 1129 -1042 1129 -1042 0 3
rlabel polysilicon 1136 -1036 1136 -1036 0 1
rlabel polysilicon 1136 -1042 1136 -1042 0 3
rlabel polysilicon 1143 -1036 1143 -1036 0 1
rlabel polysilicon 1143 -1042 1143 -1042 0 3
rlabel polysilicon 1150 -1036 1150 -1036 0 1
rlabel polysilicon 1150 -1042 1150 -1042 0 3
rlabel polysilicon 1157 -1036 1157 -1036 0 1
rlabel polysilicon 1157 -1042 1157 -1042 0 3
rlabel polysilicon 1164 -1036 1164 -1036 0 1
rlabel polysilicon 1164 -1042 1164 -1042 0 3
rlabel polysilicon 1171 -1036 1171 -1036 0 1
rlabel polysilicon 1171 -1042 1171 -1042 0 3
rlabel polysilicon 1178 -1036 1178 -1036 0 1
rlabel polysilicon 1178 -1042 1178 -1042 0 3
rlabel polysilicon 1185 -1036 1185 -1036 0 1
rlabel polysilicon 1185 -1042 1185 -1042 0 3
rlabel polysilicon 1192 -1036 1192 -1036 0 1
rlabel polysilicon 1192 -1042 1192 -1042 0 3
rlabel polysilicon 1199 -1036 1199 -1036 0 1
rlabel polysilicon 1199 -1042 1199 -1042 0 3
rlabel polysilicon 1206 -1036 1206 -1036 0 1
rlabel polysilicon 1206 -1042 1206 -1042 0 3
rlabel polysilicon 1213 -1036 1213 -1036 0 1
rlabel polysilicon 1213 -1042 1213 -1042 0 3
rlabel polysilicon 1220 -1036 1220 -1036 0 1
rlabel polysilicon 1220 -1042 1220 -1042 0 3
rlabel polysilicon 1227 -1036 1227 -1036 0 1
rlabel polysilicon 1227 -1042 1227 -1042 0 3
rlabel polysilicon 1234 -1036 1234 -1036 0 1
rlabel polysilicon 1234 -1042 1234 -1042 0 3
rlabel polysilicon 1241 -1036 1241 -1036 0 1
rlabel polysilicon 1241 -1042 1241 -1042 0 3
rlabel polysilicon 1248 -1036 1248 -1036 0 1
rlabel polysilicon 1248 -1042 1248 -1042 0 3
rlabel polysilicon 1255 -1036 1255 -1036 0 1
rlabel polysilicon 1255 -1042 1255 -1042 0 3
rlabel polysilicon 1262 -1036 1262 -1036 0 1
rlabel polysilicon 1262 -1042 1262 -1042 0 3
rlabel polysilicon 1269 -1036 1269 -1036 0 1
rlabel polysilicon 1269 -1042 1269 -1042 0 3
rlabel polysilicon 1276 -1036 1276 -1036 0 1
rlabel polysilicon 1276 -1042 1276 -1042 0 3
rlabel polysilicon 1283 -1036 1283 -1036 0 1
rlabel polysilicon 1283 -1042 1283 -1042 0 3
rlabel polysilicon 1290 -1036 1290 -1036 0 1
rlabel polysilicon 1290 -1042 1290 -1042 0 3
rlabel polysilicon 1297 -1036 1297 -1036 0 1
rlabel polysilicon 1297 -1042 1297 -1042 0 3
rlabel polysilicon 1304 -1036 1304 -1036 0 1
rlabel polysilicon 1304 -1042 1304 -1042 0 3
rlabel polysilicon 1311 -1036 1311 -1036 0 1
rlabel polysilicon 1311 -1042 1311 -1042 0 3
rlabel polysilicon 1318 -1036 1318 -1036 0 1
rlabel polysilicon 1318 -1042 1318 -1042 0 3
rlabel polysilicon 1325 -1036 1325 -1036 0 1
rlabel polysilicon 1325 -1042 1325 -1042 0 3
rlabel polysilicon 1332 -1036 1332 -1036 0 1
rlabel polysilicon 1332 -1042 1332 -1042 0 3
rlabel polysilicon 1339 -1036 1339 -1036 0 1
rlabel polysilicon 1339 -1042 1339 -1042 0 3
rlabel polysilicon 1346 -1036 1346 -1036 0 1
rlabel polysilicon 1346 -1042 1346 -1042 0 3
rlabel polysilicon 1353 -1036 1353 -1036 0 1
rlabel polysilicon 1353 -1042 1353 -1042 0 3
rlabel polysilicon 1360 -1036 1360 -1036 0 1
rlabel polysilicon 1360 -1042 1360 -1042 0 3
rlabel polysilicon 1367 -1036 1367 -1036 0 1
rlabel polysilicon 1367 -1042 1367 -1042 0 3
rlabel polysilicon 1374 -1036 1374 -1036 0 1
rlabel polysilicon 1374 -1042 1374 -1042 0 3
rlabel polysilicon 1381 -1036 1381 -1036 0 1
rlabel polysilicon 1381 -1042 1381 -1042 0 3
rlabel polysilicon 1388 -1036 1388 -1036 0 1
rlabel polysilicon 1388 -1042 1388 -1042 0 3
rlabel polysilicon 1395 -1036 1395 -1036 0 1
rlabel polysilicon 1395 -1042 1395 -1042 0 3
rlabel polysilicon 1402 -1036 1402 -1036 0 1
rlabel polysilicon 1402 -1042 1402 -1042 0 3
rlabel polysilicon 1409 -1036 1409 -1036 0 1
rlabel polysilicon 1409 -1042 1409 -1042 0 3
rlabel polysilicon 1416 -1036 1416 -1036 0 1
rlabel polysilicon 1416 -1042 1416 -1042 0 3
rlabel polysilicon 1423 -1036 1423 -1036 0 1
rlabel polysilicon 1423 -1042 1423 -1042 0 3
rlabel polysilicon 1430 -1036 1430 -1036 0 1
rlabel polysilicon 1430 -1042 1430 -1042 0 3
rlabel polysilicon 1437 -1036 1437 -1036 0 1
rlabel polysilicon 1437 -1042 1437 -1042 0 3
rlabel polysilicon 1444 -1036 1444 -1036 0 1
rlabel polysilicon 1444 -1042 1444 -1042 0 3
rlabel polysilicon 1451 -1036 1451 -1036 0 1
rlabel polysilicon 1451 -1042 1451 -1042 0 3
rlabel polysilicon 1458 -1036 1458 -1036 0 1
rlabel polysilicon 1458 -1042 1458 -1042 0 3
rlabel polysilicon 1465 -1036 1465 -1036 0 1
rlabel polysilicon 1465 -1042 1465 -1042 0 3
rlabel polysilicon 1472 -1036 1472 -1036 0 1
rlabel polysilicon 1472 -1042 1472 -1042 0 3
rlabel polysilicon 1479 -1036 1479 -1036 0 1
rlabel polysilicon 1479 -1042 1479 -1042 0 3
rlabel polysilicon 1486 -1036 1486 -1036 0 1
rlabel polysilicon 1486 -1042 1486 -1042 0 3
rlabel polysilicon 1493 -1036 1493 -1036 0 1
rlabel polysilicon 1493 -1042 1493 -1042 0 3
rlabel polysilicon 1500 -1036 1500 -1036 0 1
rlabel polysilicon 1500 -1042 1500 -1042 0 3
rlabel polysilicon 1507 -1036 1507 -1036 0 1
rlabel polysilicon 1507 -1042 1507 -1042 0 3
rlabel polysilicon 1514 -1036 1514 -1036 0 1
rlabel polysilicon 1514 -1042 1514 -1042 0 3
rlabel polysilicon 1521 -1036 1521 -1036 0 1
rlabel polysilicon 1521 -1042 1521 -1042 0 3
rlabel polysilicon 1528 -1036 1528 -1036 0 1
rlabel polysilicon 1528 -1042 1528 -1042 0 3
rlabel polysilicon 1535 -1036 1535 -1036 0 1
rlabel polysilicon 1535 -1042 1535 -1042 0 3
rlabel polysilicon 1542 -1036 1542 -1036 0 1
rlabel polysilicon 1542 -1042 1542 -1042 0 3
rlabel polysilicon 1549 -1036 1549 -1036 0 1
rlabel polysilicon 1549 -1042 1549 -1042 0 3
rlabel polysilicon 1556 -1036 1556 -1036 0 1
rlabel polysilicon 1556 -1042 1556 -1042 0 3
rlabel polysilicon 1563 -1036 1563 -1036 0 1
rlabel polysilicon 1563 -1042 1563 -1042 0 3
rlabel polysilicon 1570 -1036 1570 -1036 0 1
rlabel polysilicon 1570 -1042 1570 -1042 0 3
rlabel polysilicon 1577 -1036 1577 -1036 0 1
rlabel polysilicon 1577 -1042 1577 -1042 0 3
rlabel polysilicon 1584 -1036 1584 -1036 0 1
rlabel polysilicon 1584 -1042 1584 -1042 0 3
rlabel polysilicon 1591 -1036 1591 -1036 0 1
rlabel polysilicon 1591 -1042 1591 -1042 0 3
rlabel polysilicon 1598 -1036 1598 -1036 0 1
rlabel polysilicon 1598 -1042 1598 -1042 0 3
rlabel polysilicon 1605 -1036 1605 -1036 0 1
rlabel polysilicon 1605 -1042 1605 -1042 0 3
rlabel polysilicon 1612 -1036 1612 -1036 0 1
rlabel polysilicon 1612 -1042 1612 -1042 0 3
rlabel polysilicon 1619 -1036 1619 -1036 0 1
rlabel polysilicon 1619 -1042 1619 -1042 0 3
rlabel polysilicon 1626 -1036 1626 -1036 0 1
rlabel polysilicon 1626 -1042 1626 -1042 0 3
rlabel polysilicon 1633 -1036 1633 -1036 0 1
rlabel polysilicon 1633 -1042 1633 -1042 0 3
rlabel polysilicon 1640 -1036 1640 -1036 0 1
rlabel polysilicon 1640 -1042 1640 -1042 0 3
rlabel polysilicon 1647 -1036 1647 -1036 0 1
rlabel polysilicon 1647 -1042 1647 -1042 0 3
rlabel polysilicon 1654 -1036 1654 -1036 0 1
rlabel polysilicon 1654 -1042 1654 -1042 0 3
rlabel polysilicon 1661 -1036 1661 -1036 0 1
rlabel polysilicon 1661 -1042 1661 -1042 0 3
rlabel polysilicon 1668 -1036 1668 -1036 0 1
rlabel polysilicon 1668 -1042 1668 -1042 0 3
rlabel polysilicon 1675 -1036 1675 -1036 0 1
rlabel polysilicon 1675 -1042 1675 -1042 0 3
rlabel polysilicon 1682 -1036 1682 -1036 0 1
rlabel polysilicon 1682 -1042 1682 -1042 0 3
rlabel polysilicon 1689 -1036 1689 -1036 0 1
rlabel polysilicon 1689 -1042 1689 -1042 0 3
rlabel polysilicon 1696 -1036 1696 -1036 0 1
rlabel polysilicon 1696 -1042 1696 -1042 0 3
rlabel polysilicon 1703 -1036 1703 -1036 0 1
rlabel polysilicon 1703 -1042 1703 -1042 0 3
rlabel polysilicon 1710 -1036 1710 -1036 0 1
rlabel polysilicon 1710 -1042 1710 -1042 0 3
rlabel polysilicon 1717 -1036 1717 -1036 0 1
rlabel polysilicon 1717 -1042 1717 -1042 0 3
rlabel polysilicon 1724 -1036 1724 -1036 0 1
rlabel polysilicon 1724 -1042 1724 -1042 0 3
rlabel polysilicon 30 -1187 30 -1187 0 1
rlabel polysilicon 30 -1193 30 -1193 0 3
rlabel polysilicon 37 -1187 37 -1187 0 1
rlabel polysilicon 37 -1193 37 -1193 0 3
rlabel polysilicon 44 -1187 44 -1187 0 1
rlabel polysilicon 44 -1193 44 -1193 0 3
rlabel polysilicon 51 -1187 51 -1187 0 1
rlabel polysilicon 51 -1193 51 -1193 0 3
rlabel polysilicon 58 -1187 58 -1187 0 1
rlabel polysilicon 58 -1193 58 -1193 0 3
rlabel polysilicon 65 -1187 65 -1187 0 1
rlabel polysilicon 65 -1193 65 -1193 0 3
rlabel polysilicon 75 -1187 75 -1187 0 2
rlabel polysilicon 75 -1193 75 -1193 0 4
rlabel polysilicon 79 -1187 79 -1187 0 1
rlabel polysilicon 82 -1193 82 -1193 0 4
rlabel polysilicon 89 -1187 89 -1187 0 2
rlabel polysilicon 86 -1193 86 -1193 0 3
rlabel polysilicon 89 -1193 89 -1193 0 4
rlabel polysilicon 93 -1187 93 -1187 0 1
rlabel polysilicon 93 -1193 93 -1193 0 3
rlabel polysilicon 100 -1187 100 -1187 0 1
rlabel polysilicon 103 -1187 103 -1187 0 2
rlabel polysilicon 107 -1187 107 -1187 0 1
rlabel polysilicon 107 -1193 107 -1193 0 3
rlabel polysilicon 114 -1187 114 -1187 0 1
rlabel polysilicon 114 -1193 114 -1193 0 3
rlabel polysilicon 121 -1187 121 -1187 0 1
rlabel polysilicon 124 -1187 124 -1187 0 2
rlabel polysilicon 121 -1193 121 -1193 0 3
rlabel polysilicon 124 -1193 124 -1193 0 4
rlabel polysilicon 128 -1187 128 -1187 0 1
rlabel polysilicon 128 -1193 128 -1193 0 3
rlabel polysilicon 135 -1187 135 -1187 0 1
rlabel polysilicon 135 -1193 135 -1193 0 3
rlabel polysilicon 142 -1187 142 -1187 0 1
rlabel polysilicon 142 -1193 142 -1193 0 3
rlabel polysilicon 149 -1187 149 -1187 0 1
rlabel polysilicon 149 -1193 149 -1193 0 3
rlabel polysilicon 152 -1193 152 -1193 0 4
rlabel polysilicon 156 -1187 156 -1187 0 1
rlabel polysilicon 156 -1193 156 -1193 0 3
rlabel polysilicon 163 -1187 163 -1187 0 1
rlabel polysilicon 166 -1187 166 -1187 0 2
rlabel polysilicon 163 -1193 163 -1193 0 3
rlabel polysilicon 166 -1193 166 -1193 0 4
rlabel polysilicon 170 -1187 170 -1187 0 1
rlabel polysilicon 170 -1193 170 -1193 0 3
rlabel polysilicon 177 -1187 177 -1187 0 1
rlabel polysilicon 177 -1193 177 -1193 0 3
rlabel polysilicon 184 -1187 184 -1187 0 1
rlabel polysilicon 187 -1187 187 -1187 0 2
rlabel polysilicon 184 -1193 184 -1193 0 3
rlabel polysilicon 191 -1187 191 -1187 0 1
rlabel polysilicon 191 -1193 191 -1193 0 3
rlabel polysilicon 198 -1187 198 -1187 0 1
rlabel polysilicon 201 -1187 201 -1187 0 2
rlabel polysilicon 198 -1193 198 -1193 0 3
rlabel polysilicon 201 -1193 201 -1193 0 4
rlabel polysilicon 205 -1187 205 -1187 0 1
rlabel polysilicon 208 -1187 208 -1187 0 2
rlabel polysilicon 205 -1193 205 -1193 0 3
rlabel polysilicon 208 -1193 208 -1193 0 4
rlabel polysilicon 212 -1187 212 -1187 0 1
rlabel polysilicon 212 -1193 212 -1193 0 3
rlabel polysilicon 219 -1187 219 -1187 0 1
rlabel polysilicon 219 -1193 219 -1193 0 3
rlabel polysilicon 226 -1187 226 -1187 0 1
rlabel polysilicon 226 -1193 226 -1193 0 3
rlabel polysilicon 236 -1187 236 -1187 0 2
rlabel polysilicon 233 -1193 233 -1193 0 3
rlabel polysilicon 236 -1193 236 -1193 0 4
rlabel polysilicon 240 -1187 240 -1187 0 1
rlabel polysilicon 240 -1193 240 -1193 0 3
rlabel polysilicon 247 -1187 247 -1187 0 1
rlabel polysilicon 247 -1193 247 -1193 0 3
rlabel polysilicon 254 -1187 254 -1187 0 1
rlabel polysilicon 257 -1193 257 -1193 0 4
rlabel polysilicon 261 -1187 261 -1187 0 1
rlabel polysilicon 261 -1193 261 -1193 0 3
rlabel polysilicon 268 -1187 268 -1187 0 1
rlabel polysilicon 268 -1193 268 -1193 0 3
rlabel polysilicon 275 -1187 275 -1187 0 1
rlabel polysilicon 278 -1193 278 -1193 0 4
rlabel polysilicon 282 -1187 282 -1187 0 1
rlabel polysilicon 282 -1193 282 -1193 0 3
rlabel polysilicon 289 -1187 289 -1187 0 1
rlabel polysilicon 289 -1193 289 -1193 0 3
rlabel polysilicon 296 -1187 296 -1187 0 1
rlabel polysilicon 296 -1193 296 -1193 0 3
rlabel polysilicon 303 -1187 303 -1187 0 1
rlabel polysilicon 303 -1193 303 -1193 0 3
rlabel polysilicon 310 -1187 310 -1187 0 1
rlabel polysilicon 310 -1193 310 -1193 0 3
rlabel polysilicon 317 -1187 317 -1187 0 1
rlabel polysilicon 317 -1193 317 -1193 0 3
rlabel polysilicon 324 -1187 324 -1187 0 1
rlabel polysilicon 324 -1193 324 -1193 0 3
rlabel polysilicon 331 -1187 331 -1187 0 1
rlabel polysilicon 331 -1193 331 -1193 0 3
rlabel polysilicon 338 -1187 338 -1187 0 1
rlabel polysilicon 338 -1193 338 -1193 0 3
rlabel polysilicon 345 -1187 345 -1187 0 1
rlabel polysilicon 345 -1193 345 -1193 0 3
rlabel polysilicon 352 -1187 352 -1187 0 1
rlabel polysilicon 352 -1193 352 -1193 0 3
rlabel polysilicon 359 -1187 359 -1187 0 1
rlabel polysilicon 359 -1193 359 -1193 0 3
rlabel polysilicon 366 -1187 366 -1187 0 1
rlabel polysilicon 366 -1193 366 -1193 0 3
rlabel polysilicon 373 -1187 373 -1187 0 1
rlabel polysilicon 373 -1193 373 -1193 0 3
rlabel polysilicon 380 -1187 380 -1187 0 1
rlabel polysilicon 380 -1193 380 -1193 0 3
rlabel polysilicon 387 -1187 387 -1187 0 1
rlabel polysilicon 387 -1193 387 -1193 0 3
rlabel polysilicon 394 -1187 394 -1187 0 1
rlabel polysilicon 394 -1193 394 -1193 0 3
rlabel polysilicon 401 -1187 401 -1187 0 1
rlabel polysilicon 401 -1193 401 -1193 0 3
rlabel polysilicon 408 -1187 408 -1187 0 1
rlabel polysilicon 408 -1193 408 -1193 0 3
rlabel polysilicon 415 -1187 415 -1187 0 1
rlabel polysilicon 415 -1193 415 -1193 0 3
rlabel polysilicon 422 -1187 422 -1187 0 1
rlabel polysilicon 422 -1193 422 -1193 0 3
rlabel polysilicon 429 -1187 429 -1187 0 1
rlabel polysilicon 429 -1193 429 -1193 0 3
rlabel polysilicon 436 -1187 436 -1187 0 1
rlabel polysilicon 436 -1193 436 -1193 0 3
rlabel polysilicon 443 -1187 443 -1187 0 1
rlabel polysilicon 443 -1193 443 -1193 0 3
rlabel polysilicon 450 -1187 450 -1187 0 1
rlabel polysilicon 450 -1193 450 -1193 0 3
rlabel polysilicon 457 -1187 457 -1187 0 1
rlabel polysilicon 457 -1193 457 -1193 0 3
rlabel polysilicon 464 -1187 464 -1187 0 1
rlabel polysilicon 467 -1187 467 -1187 0 2
rlabel polysilicon 464 -1193 464 -1193 0 3
rlabel polysilicon 467 -1193 467 -1193 0 4
rlabel polysilicon 471 -1187 471 -1187 0 1
rlabel polysilicon 471 -1193 471 -1193 0 3
rlabel polysilicon 478 -1187 478 -1187 0 1
rlabel polysilicon 478 -1193 478 -1193 0 3
rlabel polysilicon 485 -1187 485 -1187 0 1
rlabel polysilicon 488 -1187 488 -1187 0 2
rlabel polysilicon 488 -1193 488 -1193 0 4
rlabel polysilicon 492 -1187 492 -1187 0 1
rlabel polysilicon 492 -1193 492 -1193 0 3
rlabel polysilicon 499 -1187 499 -1187 0 1
rlabel polysilicon 499 -1193 499 -1193 0 3
rlabel polysilicon 506 -1187 506 -1187 0 1
rlabel polysilicon 509 -1193 509 -1193 0 4
rlabel polysilicon 513 -1187 513 -1187 0 1
rlabel polysilicon 516 -1187 516 -1187 0 2
rlabel polysilicon 513 -1193 513 -1193 0 3
rlabel polysilicon 516 -1193 516 -1193 0 4
rlabel polysilicon 520 -1187 520 -1187 0 1
rlabel polysilicon 527 -1187 527 -1187 0 1
rlabel polysilicon 527 -1193 527 -1193 0 3
rlabel polysilicon 534 -1187 534 -1187 0 1
rlabel polysilicon 534 -1193 534 -1193 0 3
rlabel polysilicon 541 -1187 541 -1187 0 1
rlabel polysilicon 544 -1187 544 -1187 0 2
rlabel polysilicon 544 -1193 544 -1193 0 4
rlabel polysilicon 548 -1187 548 -1187 0 1
rlabel polysilicon 548 -1193 548 -1193 0 3
rlabel polysilicon 555 -1187 555 -1187 0 1
rlabel polysilicon 555 -1193 555 -1193 0 3
rlabel polysilicon 562 -1187 562 -1187 0 1
rlabel polysilicon 562 -1193 562 -1193 0 3
rlabel polysilicon 569 -1187 569 -1187 0 1
rlabel polysilicon 569 -1193 569 -1193 0 3
rlabel polysilicon 579 -1187 579 -1187 0 2
rlabel polysilicon 576 -1193 576 -1193 0 3
rlabel polysilicon 583 -1187 583 -1187 0 1
rlabel polysilicon 583 -1193 583 -1193 0 3
rlabel polysilicon 590 -1187 590 -1187 0 1
rlabel polysilicon 590 -1193 590 -1193 0 3
rlabel polysilicon 597 -1187 597 -1187 0 1
rlabel polysilicon 600 -1187 600 -1187 0 2
rlabel polysilicon 597 -1193 597 -1193 0 3
rlabel polysilicon 604 -1187 604 -1187 0 1
rlabel polysilicon 604 -1193 604 -1193 0 3
rlabel polysilicon 611 -1187 611 -1187 0 1
rlabel polysilicon 614 -1187 614 -1187 0 2
rlabel polysilicon 611 -1193 611 -1193 0 3
rlabel polysilicon 614 -1193 614 -1193 0 4
rlabel polysilicon 621 -1187 621 -1187 0 2
rlabel polysilicon 618 -1193 618 -1193 0 3
rlabel polysilicon 621 -1193 621 -1193 0 4
rlabel polysilicon 625 -1187 625 -1187 0 1
rlabel polysilicon 625 -1193 625 -1193 0 3
rlabel polysilicon 632 -1187 632 -1187 0 1
rlabel polysilicon 632 -1193 632 -1193 0 3
rlabel polysilicon 639 -1187 639 -1187 0 1
rlabel polysilicon 639 -1193 639 -1193 0 3
rlabel polysilicon 646 -1187 646 -1187 0 1
rlabel polysilicon 646 -1193 646 -1193 0 3
rlabel polysilicon 653 -1187 653 -1187 0 1
rlabel polysilicon 653 -1193 653 -1193 0 3
rlabel polysilicon 660 -1187 660 -1187 0 1
rlabel polysilicon 663 -1187 663 -1187 0 2
rlabel polysilicon 660 -1193 660 -1193 0 3
rlabel polysilicon 663 -1193 663 -1193 0 4
rlabel polysilicon 667 -1187 667 -1187 0 1
rlabel polysilicon 667 -1193 667 -1193 0 3
rlabel polysilicon 674 -1187 674 -1187 0 1
rlabel polysilicon 674 -1193 674 -1193 0 3
rlabel polysilicon 681 -1187 681 -1187 0 1
rlabel polysilicon 681 -1193 681 -1193 0 3
rlabel polysilicon 688 -1187 688 -1187 0 1
rlabel polysilicon 688 -1193 688 -1193 0 3
rlabel polysilicon 695 -1187 695 -1187 0 1
rlabel polysilicon 695 -1193 695 -1193 0 3
rlabel polysilicon 702 -1187 702 -1187 0 1
rlabel polysilicon 702 -1193 702 -1193 0 3
rlabel polysilicon 709 -1187 709 -1187 0 1
rlabel polysilicon 709 -1193 709 -1193 0 3
rlabel polysilicon 716 -1187 716 -1187 0 1
rlabel polysilicon 719 -1187 719 -1187 0 2
rlabel polysilicon 719 -1193 719 -1193 0 4
rlabel polysilicon 723 -1187 723 -1187 0 1
rlabel polysilicon 726 -1187 726 -1187 0 2
rlabel polysilicon 723 -1193 723 -1193 0 3
rlabel polysilicon 726 -1193 726 -1193 0 4
rlabel polysilicon 730 -1187 730 -1187 0 1
rlabel polysilicon 730 -1193 730 -1193 0 3
rlabel polysilicon 737 -1187 737 -1187 0 1
rlabel polysilicon 737 -1193 737 -1193 0 3
rlabel polysilicon 744 -1187 744 -1187 0 1
rlabel polysilicon 747 -1187 747 -1187 0 2
rlabel polysilicon 744 -1193 744 -1193 0 3
rlabel polysilicon 747 -1193 747 -1193 0 4
rlabel polysilicon 751 -1187 751 -1187 0 1
rlabel polysilicon 754 -1187 754 -1187 0 2
rlabel polysilicon 751 -1193 751 -1193 0 3
rlabel polysilicon 758 -1187 758 -1187 0 1
rlabel polysilicon 758 -1193 758 -1193 0 3
rlabel polysilicon 765 -1187 765 -1187 0 1
rlabel polysilicon 765 -1193 765 -1193 0 3
rlabel polysilicon 772 -1187 772 -1187 0 1
rlabel polysilicon 772 -1193 772 -1193 0 3
rlabel polysilicon 779 -1187 779 -1187 0 1
rlabel polysilicon 779 -1193 779 -1193 0 3
rlabel polysilicon 786 -1187 786 -1187 0 1
rlabel polysilicon 786 -1193 786 -1193 0 3
rlabel polysilicon 793 -1187 793 -1187 0 1
rlabel polysilicon 793 -1193 793 -1193 0 3
rlabel polysilicon 800 -1187 800 -1187 0 1
rlabel polysilicon 800 -1193 800 -1193 0 3
rlabel polysilicon 807 -1187 807 -1187 0 1
rlabel polysilicon 807 -1193 807 -1193 0 3
rlabel polysilicon 814 -1187 814 -1187 0 1
rlabel polysilicon 814 -1193 814 -1193 0 3
rlabel polysilicon 821 -1187 821 -1187 0 1
rlabel polysilicon 821 -1193 821 -1193 0 3
rlabel polysilicon 828 -1187 828 -1187 0 1
rlabel polysilicon 828 -1193 828 -1193 0 3
rlabel polysilicon 831 -1193 831 -1193 0 4
rlabel polysilicon 835 -1187 835 -1187 0 1
rlabel polysilicon 835 -1193 835 -1193 0 3
rlabel polysilicon 842 -1187 842 -1187 0 1
rlabel polysilicon 842 -1193 842 -1193 0 3
rlabel polysilicon 849 -1187 849 -1187 0 1
rlabel polysilicon 849 -1193 849 -1193 0 3
rlabel polysilicon 856 -1187 856 -1187 0 1
rlabel polysilicon 856 -1193 856 -1193 0 3
rlabel polysilicon 863 -1187 863 -1187 0 1
rlabel polysilicon 863 -1193 863 -1193 0 3
rlabel polysilicon 870 -1187 870 -1187 0 1
rlabel polysilicon 870 -1193 870 -1193 0 3
rlabel polysilicon 873 -1193 873 -1193 0 4
rlabel polysilicon 877 -1187 877 -1187 0 1
rlabel polysilicon 877 -1193 877 -1193 0 3
rlabel polysilicon 884 -1187 884 -1187 0 1
rlabel polysilicon 884 -1193 884 -1193 0 3
rlabel polysilicon 894 -1187 894 -1187 0 2
rlabel polysilicon 891 -1193 891 -1193 0 3
rlabel polysilicon 894 -1193 894 -1193 0 4
rlabel polysilicon 898 -1187 898 -1187 0 1
rlabel polysilicon 901 -1187 901 -1187 0 2
rlabel polysilicon 898 -1193 898 -1193 0 3
rlabel polysilicon 901 -1193 901 -1193 0 4
rlabel polysilicon 905 -1187 905 -1187 0 1
rlabel polysilicon 905 -1193 905 -1193 0 3
rlabel polysilicon 912 -1187 912 -1187 0 1
rlabel polysilicon 912 -1193 912 -1193 0 3
rlabel polysilicon 919 -1187 919 -1187 0 1
rlabel polysilicon 919 -1193 919 -1193 0 3
rlabel polysilicon 926 -1187 926 -1187 0 1
rlabel polysilicon 926 -1193 926 -1193 0 3
rlabel polysilicon 933 -1187 933 -1187 0 1
rlabel polysilicon 933 -1193 933 -1193 0 3
rlabel polysilicon 940 -1187 940 -1187 0 1
rlabel polysilicon 940 -1193 940 -1193 0 3
rlabel polysilicon 947 -1187 947 -1187 0 1
rlabel polysilicon 947 -1193 947 -1193 0 3
rlabel polysilicon 954 -1187 954 -1187 0 1
rlabel polysilicon 957 -1187 957 -1187 0 2
rlabel polysilicon 954 -1193 954 -1193 0 3
rlabel polysilicon 957 -1193 957 -1193 0 4
rlabel polysilicon 961 -1187 961 -1187 0 1
rlabel polysilicon 961 -1193 961 -1193 0 3
rlabel polysilicon 968 -1187 968 -1187 0 1
rlabel polysilicon 971 -1187 971 -1187 0 2
rlabel polysilicon 968 -1193 968 -1193 0 3
rlabel polysilicon 971 -1193 971 -1193 0 4
rlabel polysilicon 975 -1187 975 -1187 0 1
rlabel polysilicon 975 -1193 975 -1193 0 3
rlabel polysilicon 982 -1187 982 -1187 0 1
rlabel polysilicon 982 -1193 982 -1193 0 3
rlabel polysilicon 989 -1187 989 -1187 0 1
rlabel polysilicon 992 -1187 992 -1187 0 2
rlabel polysilicon 989 -1193 989 -1193 0 3
rlabel polysilicon 992 -1193 992 -1193 0 4
rlabel polysilicon 996 -1187 996 -1187 0 1
rlabel polysilicon 996 -1193 996 -1193 0 3
rlabel polysilicon 999 -1193 999 -1193 0 4
rlabel polysilicon 1003 -1187 1003 -1187 0 1
rlabel polysilicon 1003 -1193 1003 -1193 0 3
rlabel polysilicon 1010 -1187 1010 -1187 0 1
rlabel polysilicon 1010 -1193 1010 -1193 0 3
rlabel polysilicon 1017 -1187 1017 -1187 0 1
rlabel polysilicon 1017 -1193 1017 -1193 0 3
rlabel polysilicon 1024 -1187 1024 -1187 0 1
rlabel polysilicon 1024 -1193 1024 -1193 0 3
rlabel polysilicon 1031 -1187 1031 -1187 0 1
rlabel polysilicon 1031 -1193 1031 -1193 0 3
rlabel polysilicon 1038 -1187 1038 -1187 0 1
rlabel polysilicon 1038 -1193 1038 -1193 0 3
rlabel polysilicon 1045 -1187 1045 -1187 0 1
rlabel polysilicon 1048 -1187 1048 -1187 0 2
rlabel polysilicon 1045 -1193 1045 -1193 0 3
rlabel polysilicon 1048 -1193 1048 -1193 0 4
rlabel polysilicon 1052 -1187 1052 -1187 0 1
rlabel polysilicon 1052 -1193 1052 -1193 0 3
rlabel polysilicon 1059 -1187 1059 -1187 0 1
rlabel polysilicon 1059 -1193 1059 -1193 0 3
rlabel polysilicon 1066 -1187 1066 -1187 0 1
rlabel polysilicon 1066 -1193 1066 -1193 0 3
rlabel polysilicon 1073 -1187 1073 -1187 0 1
rlabel polysilicon 1073 -1193 1073 -1193 0 3
rlabel polysilicon 1080 -1187 1080 -1187 0 1
rlabel polysilicon 1080 -1193 1080 -1193 0 3
rlabel polysilicon 1087 -1187 1087 -1187 0 1
rlabel polysilicon 1087 -1193 1087 -1193 0 3
rlabel polysilicon 1094 -1187 1094 -1187 0 1
rlabel polysilicon 1094 -1193 1094 -1193 0 3
rlabel polysilicon 1101 -1187 1101 -1187 0 1
rlabel polysilicon 1101 -1193 1101 -1193 0 3
rlabel polysilicon 1108 -1187 1108 -1187 0 1
rlabel polysilicon 1108 -1193 1108 -1193 0 3
rlabel polysilicon 1115 -1187 1115 -1187 0 1
rlabel polysilicon 1115 -1193 1115 -1193 0 3
rlabel polysilicon 1122 -1187 1122 -1187 0 1
rlabel polysilicon 1122 -1193 1122 -1193 0 3
rlabel polysilicon 1129 -1187 1129 -1187 0 1
rlabel polysilicon 1129 -1193 1129 -1193 0 3
rlabel polysilicon 1136 -1187 1136 -1187 0 1
rlabel polysilicon 1136 -1193 1136 -1193 0 3
rlabel polysilicon 1143 -1187 1143 -1187 0 1
rlabel polysilicon 1143 -1193 1143 -1193 0 3
rlabel polysilicon 1150 -1187 1150 -1187 0 1
rlabel polysilicon 1150 -1193 1150 -1193 0 3
rlabel polysilicon 1157 -1187 1157 -1187 0 1
rlabel polysilicon 1157 -1193 1157 -1193 0 3
rlabel polysilicon 1164 -1187 1164 -1187 0 1
rlabel polysilicon 1164 -1193 1164 -1193 0 3
rlabel polysilicon 1171 -1187 1171 -1187 0 1
rlabel polysilicon 1171 -1193 1171 -1193 0 3
rlabel polysilicon 1178 -1187 1178 -1187 0 1
rlabel polysilicon 1178 -1193 1178 -1193 0 3
rlabel polysilicon 1185 -1187 1185 -1187 0 1
rlabel polysilicon 1185 -1193 1185 -1193 0 3
rlabel polysilicon 1192 -1187 1192 -1187 0 1
rlabel polysilicon 1192 -1193 1192 -1193 0 3
rlabel polysilicon 1199 -1187 1199 -1187 0 1
rlabel polysilicon 1199 -1193 1199 -1193 0 3
rlabel polysilicon 1206 -1187 1206 -1187 0 1
rlabel polysilicon 1206 -1193 1206 -1193 0 3
rlabel polysilicon 1213 -1187 1213 -1187 0 1
rlabel polysilicon 1213 -1193 1213 -1193 0 3
rlabel polysilicon 1220 -1187 1220 -1187 0 1
rlabel polysilicon 1220 -1193 1220 -1193 0 3
rlabel polysilicon 1227 -1187 1227 -1187 0 1
rlabel polysilicon 1227 -1193 1227 -1193 0 3
rlabel polysilicon 1234 -1187 1234 -1187 0 1
rlabel polysilicon 1234 -1193 1234 -1193 0 3
rlabel polysilicon 1241 -1187 1241 -1187 0 1
rlabel polysilicon 1241 -1193 1241 -1193 0 3
rlabel polysilicon 1248 -1187 1248 -1187 0 1
rlabel polysilicon 1248 -1193 1248 -1193 0 3
rlabel polysilicon 1255 -1187 1255 -1187 0 1
rlabel polysilicon 1255 -1193 1255 -1193 0 3
rlabel polysilicon 1262 -1187 1262 -1187 0 1
rlabel polysilicon 1262 -1193 1262 -1193 0 3
rlabel polysilicon 1269 -1187 1269 -1187 0 1
rlabel polysilicon 1269 -1193 1269 -1193 0 3
rlabel polysilicon 1276 -1187 1276 -1187 0 1
rlabel polysilicon 1276 -1193 1276 -1193 0 3
rlabel polysilicon 1283 -1187 1283 -1187 0 1
rlabel polysilicon 1283 -1193 1283 -1193 0 3
rlabel polysilicon 1290 -1187 1290 -1187 0 1
rlabel polysilicon 1290 -1193 1290 -1193 0 3
rlabel polysilicon 1297 -1187 1297 -1187 0 1
rlabel polysilicon 1297 -1193 1297 -1193 0 3
rlabel polysilicon 1304 -1187 1304 -1187 0 1
rlabel polysilicon 1304 -1193 1304 -1193 0 3
rlabel polysilicon 1311 -1187 1311 -1187 0 1
rlabel polysilicon 1311 -1193 1311 -1193 0 3
rlabel polysilicon 1318 -1187 1318 -1187 0 1
rlabel polysilicon 1318 -1193 1318 -1193 0 3
rlabel polysilicon 1325 -1187 1325 -1187 0 1
rlabel polysilicon 1325 -1193 1325 -1193 0 3
rlabel polysilicon 1332 -1187 1332 -1187 0 1
rlabel polysilicon 1332 -1193 1332 -1193 0 3
rlabel polysilicon 1339 -1187 1339 -1187 0 1
rlabel polysilicon 1339 -1193 1339 -1193 0 3
rlabel polysilicon 1346 -1187 1346 -1187 0 1
rlabel polysilicon 1346 -1193 1346 -1193 0 3
rlabel polysilicon 1353 -1187 1353 -1187 0 1
rlabel polysilicon 1353 -1193 1353 -1193 0 3
rlabel polysilicon 1360 -1187 1360 -1187 0 1
rlabel polysilicon 1360 -1193 1360 -1193 0 3
rlabel polysilicon 1367 -1187 1367 -1187 0 1
rlabel polysilicon 1367 -1193 1367 -1193 0 3
rlabel polysilicon 1374 -1187 1374 -1187 0 1
rlabel polysilicon 1374 -1193 1374 -1193 0 3
rlabel polysilicon 1381 -1187 1381 -1187 0 1
rlabel polysilicon 1381 -1193 1381 -1193 0 3
rlabel polysilicon 1388 -1187 1388 -1187 0 1
rlabel polysilicon 1388 -1193 1388 -1193 0 3
rlabel polysilicon 1395 -1187 1395 -1187 0 1
rlabel polysilicon 1395 -1193 1395 -1193 0 3
rlabel polysilicon 1402 -1187 1402 -1187 0 1
rlabel polysilicon 1402 -1193 1402 -1193 0 3
rlabel polysilicon 1409 -1187 1409 -1187 0 1
rlabel polysilicon 1409 -1193 1409 -1193 0 3
rlabel polysilicon 1416 -1187 1416 -1187 0 1
rlabel polysilicon 1416 -1193 1416 -1193 0 3
rlabel polysilicon 1423 -1187 1423 -1187 0 1
rlabel polysilicon 1423 -1193 1423 -1193 0 3
rlabel polysilicon 1430 -1187 1430 -1187 0 1
rlabel polysilicon 1430 -1193 1430 -1193 0 3
rlabel polysilicon 1437 -1187 1437 -1187 0 1
rlabel polysilicon 1437 -1193 1437 -1193 0 3
rlabel polysilicon 1444 -1187 1444 -1187 0 1
rlabel polysilicon 1444 -1193 1444 -1193 0 3
rlabel polysilicon 1451 -1187 1451 -1187 0 1
rlabel polysilicon 1451 -1193 1451 -1193 0 3
rlabel polysilicon 1458 -1187 1458 -1187 0 1
rlabel polysilicon 1458 -1193 1458 -1193 0 3
rlabel polysilicon 1465 -1187 1465 -1187 0 1
rlabel polysilicon 1465 -1193 1465 -1193 0 3
rlabel polysilicon 1472 -1187 1472 -1187 0 1
rlabel polysilicon 1472 -1193 1472 -1193 0 3
rlabel polysilicon 1479 -1187 1479 -1187 0 1
rlabel polysilicon 1479 -1193 1479 -1193 0 3
rlabel polysilicon 1486 -1187 1486 -1187 0 1
rlabel polysilicon 1486 -1193 1486 -1193 0 3
rlabel polysilicon 1493 -1187 1493 -1187 0 1
rlabel polysilicon 1493 -1193 1493 -1193 0 3
rlabel polysilicon 1500 -1187 1500 -1187 0 1
rlabel polysilicon 1500 -1193 1500 -1193 0 3
rlabel polysilicon 1507 -1187 1507 -1187 0 1
rlabel polysilicon 1507 -1193 1507 -1193 0 3
rlabel polysilicon 1514 -1187 1514 -1187 0 1
rlabel polysilicon 1514 -1193 1514 -1193 0 3
rlabel polysilicon 1521 -1187 1521 -1187 0 1
rlabel polysilicon 1521 -1193 1521 -1193 0 3
rlabel polysilicon 1528 -1187 1528 -1187 0 1
rlabel polysilicon 1528 -1193 1528 -1193 0 3
rlabel polysilicon 1535 -1187 1535 -1187 0 1
rlabel polysilicon 1535 -1193 1535 -1193 0 3
rlabel polysilicon 1542 -1187 1542 -1187 0 1
rlabel polysilicon 1542 -1193 1542 -1193 0 3
rlabel polysilicon 1549 -1187 1549 -1187 0 1
rlabel polysilicon 1549 -1193 1549 -1193 0 3
rlabel polysilicon 1556 -1187 1556 -1187 0 1
rlabel polysilicon 1556 -1193 1556 -1193 0 3
rlabel polysilicon 1563 -1187 1563 -1187 0 1
rlabel polysilicon 1563 -1193 1563 -1193 0 3
rlabel polysilicon 1570 -1187 1570 -1187 0 1
rlabel polysilicon 1570 -1193 1570 -1193 0 3
rlabel polysilicon 1577 -1187 1577 -1187 0 1
rlabel polysilicon 1577 -1193 1577 -1193 0 3
rlabel polysilicon 1584 -1187 1584 -1187 0 1
rlabel polysilicon 1584 -1193 1584 -1193 0 3
rlabel polysilicon 1591 -1187 1591 -1187 0 1
rlabel polysilicon 1591 -1193 1591 -1193 0 3
rlabel polysilicon 1598 -1187 1598 -1187 0 1
rlabel polysilicon 1598 -1193 1598 -1193 0 3
rlabel polysilicon 1605 -1187 1605 -1187 0 1
rlabel polysilicon 1605 -1193 1605 -1193 0 3
rlabel polysilicon 1612 -1187 1612 -1187 0 1
rlabel polysilicon 1612 -1193 1612 -1193 0 3
rlabel polysilicon 1619 -1187 1619 -1187 0 1
rlabel polysilicon 1619 -1193 1619 -1193 0 3
rlabel polysilicon 1626 -1187 1626 -1187 0 1
rlabel polysilicon 1626 -1193 1626 -1193 0 3
rlabel polysilicon 1633 -1187 1633 -1187 0 1
rlabel polysilicon 1633 -1193 1633 -1193 0 3
rlabel polysilicon 1640 -1187 1640 -1187 0 1
rlabel polysilicon 1640 -1193 1640 -1193 0 3
rlabel polysilicon 1647 -1187 1647 -1187 0 1
rlabel polysilicon 1650 -1187 1650 -1187 0 2
rlabel polysilicon 1647 -1193 1647 -1193 0 3
rlabel polysilicon 1654 -1187 1654 -1187 0 1
rlabel polysilicon 1654 -1193 1654 -1193 0 3
rlabel polysilicon 1664 -1187 1664 -1187 0 2
rlabel polysilicon 1661 -1193 1661 -1193 0 3
rlabel polysilicon 1664 -1193 1664 -1193 0 4
rlabel polysilicon 1675 -1187 1675 -1187 0 1
rlabel polysilicon 1675 -1193 1675 -1193 0 3
rlabel polysilicon 1724 -1187 1724 -1187 0 1
rlabel polysilicon 1724 -1193 1724 -1193 0 3
rlabel polysilicon 1731 -1187 1731 -1187 0 1
rlabel polysilicon 1731 -1193 1731 -1193 0 3
rlabel polysilicon 23 -1318 23 -1318 0 1
rlabel polysilicon 23 -1324 23 -1324 0 3
rlabel polysilicon 30 -1318 30 -1318 0 1
rlabel polysilicon 30 -1324 30 -1324 0 3
rlabel polysilicon 37 -1318 37 -1318 0 1
rlabel polysilicon 37 -1324 37 -1324 0 3
rlabel polysilicon 44 -1318 44 -1318 0 1
rlabel polysilicon 44 -1324 44 -1324 0 3
rlabel polysilicon 51 -1318 51 -1318 0 1
rlabel polysilicon 51 -1324 51 -1324 0 3
rlabel polysilicon 58 -1318 58 -1318 0 1
rlabel polysilicon 58 -1324 58 -1324 0 3
rlabel polysilicon 65 -1318 65 -1318 0 1
rlabel polysilicon 65 -1324 65 -1324 0 3
rlabel polysilicon 75 -1318 75 -1318 0 2
rlabel polysilicon 72 -1324 72 -1324 0 3
rlabel polysilicon 79 -1318 79 -1318 0 1
rlabel polysilicon 82 -1318 82 -1318 0 2
rlabel polysilicon 82 -1324 82 -1324 0 4
rlabel polysilicon 86 -1318 86 -1318 0 1
rlabel polysilicon 86 -1324 86 -1324 0 3
rlabel polysilicon 93 -1318 93 -1318 0 1
rlabel polysilicon 96 -1318 96 -1318 0 2
rlabel polysilicon 93 -1324 93 -1324 0 3
rlabel polysilicon 96 -1324 96 -1324 0 4
rlabel polysilicon 100 -1318 100 -1318 0 1
rlabel polysilicon 100 -1324 100 -1324 0 3
rlabel polysilicon 107 -1318 107 -1318 0 1
rlabel polysilicon 107 -1324 107 -1324 0 3
rlabel polysilicon 114 -1318 114 -1318 0 1
rlabel polysilicon 114 -1324 114 -1324 0 3
rlabel polysilicon 121 -1318 121 -1318 0 1
rlabel polysilicon 124 -1318 124 -1318 0 2
rlabel polysilicon 121 -1324 121 -1324 0 3
rlabel polysilicon 124 -1324 124 -1324 0 4
rlabel polysilicon 128 -1318 128 -1318 0 1
rlabel polysilicon 128 -1324 128 -1324 0 3
rlabel polysilicon 135 -1318 135 -1318 0 1
rlabel polysilicon 135 -1324 135 -1324 0 3
rlabel polysilicon 142 -1318 142 -1318 0 1
rlabel polysilicon 145 -1318 145 -1318 0 2
rlabel polysilicon 142 -1324 142 -1324 0 3
rlabel polysilicon 145 -1324 145 -1324 0 4
rlabel polysilicon 149 -1318 149 -1318 0 1
rlabel polysilicon 149 -1324 149 -1324 0 3
rlabel polysilicon 156 -1318 156 -1318 0 1
rlabel polysilicon 156 -1324 156 -1324 0 3
rlabel polysilicon 163 -1318 163 -1318 0 1
rlabel polysilicon 166 -1318 166 -1318 0 2
rlabel polysilicon 163 -1324 163 -1324 0 3
rlabel polysilicon 170 -1318 170 -1318 0 1
rlabel polysilicon 170 -1324 170 -1324 0 3
rlabel polysilicon 177 -1318 177 -1318 0 1
rlabel polysilicon 177 -1324 177 -1324 0 3
rlabel polysilicon 184 -1318 184 -1318 0 1
rlabel polysilicon 184 -1324 184 -1324 0 3
rlabel polysilicon 191 -1318 191 -1318 0 1
rlabel polysilicon 191 -1324 191 -1324 0 3
rlabel polysilicon 198 -1318 198 -1318 0 1
rlabel polysilicon 198 -1324 198 -1324 0 3
rlabel polysilicon 205 -1318 205 -1318 0 1
rlabel polysilicon 205 -1324 205 -1324 0 3
rlabel polysilicon 212 -1318 212 -1318 0 1
rlabel polysilicon 212 -1324 212 -1324 0 3
rlabel polysilicon 219 -1318 219 -1318 0 1
rlabel polysilicon 219 -1324 219 -1324 0 3
rlabel polysilicon 226 -1318 226 -1318 0 1
rlabel polysilicon 226 -1324 226 -1324 0 3
rlabel polysilicon 233 -1318 233 -1318 0 1
rlabel polysilicon 236 -1324 236 -1324 0 4
rlabel polysilicon 240 -1318 240 -1318 0 1
rlabel polysilicon 240 -1324 240 -1324 0 3
rlabel polysilicon 250 -1318 250 -1318 0 2
rlabel polysilicon 247 -1324 247 -1324 0 3
rlabel polysilicon 250 -1324 250 -1324 0 4
rlabel polysilicon 254 -1318 254 -1318 0 1
rlabel polysilicon 254 -1324 254 -1324 0 3
rlabel polysilicon 261 -1318 261 -1318 0 1
rlabel polysilicon 261 -1324 261 -1324 0 3
rlabel polysilicon 268 -1318 268 -1318 0 1
rlabel polysilicon 268 -1324 268 -1324 0 3
rlabel polysilicon 275 -1324 275 -1324 0 3
rlabel polysilicon 278 -1324 278 -1324 0 4
rlabel polysilicon 282 -1318 282 -1318 0 1
rlabel polysilicon 282 -1324 282 -1324 0 3
rlabel polysilicon 289 -1318 289 -1318 0 1
rlabel polysilicon 289 -1324 289 -1324 0 3
rlabel polysilicon 296 -1318 296 -1318 0 1
rlabel polysilicon 296 -1324 296 -1324 0 3
rlabel polysilicon 303 -1318 303 -1318 0 1
rlabel polysilicon 303 -1324 303 -1324 0 3
rlabel polysilicon 310 -1318 310 -1318 0 1
rlabel polysilicon 310 -1324 310 -1324 0 3
rlabel polysilicon 317 -1318 317 -1318 0 1
rlabel polysilicon 317 -1324 317 -1324 0 3
rlabel polysilicon 324 -1318 324 -1318 0 1
rlabel polysilicon 324 -1324 324 -1324 0 3
rlabel polysilicon 331 -1318 331 -1318 0 1
rlabel polysilicon 331 -1324 331 -1324 0 3
rlabel polysilicon 338 -1318 338 -1318 0 1
rlabel polysilicon 338 -1324 338 -1324 0 3
rlabel polysilicon 345 -1318 345 -1318 0 1
rlabel polysilicon 345 -1324 345 -1324 0 3
rlabel polysilicon 352 -1318 352 -1318 0 1
rlabel polysilicon 352 -1324 352 -1324 0 3
rlabel polysilicon 359 -1318 359 -1318 0 1
rlabel polysilicon 359 -1324 359 -1324 0 3
rlabel polysilicon 366 -1318 366 -1318 0 1
rlabel polysilicon 366 -1324 366 -1324 0 3
rlabel polysilicon 373 -1318 373 -1318 0 1
rlabel polysilicon 373 -1324 373 -1324 0 3
rlabel polysilicon 380 -1318 380 -1318 0 1
rlabel polysilicon 380 -1324 380 -1324 0 3
rlabel polysilicon 387 -1318 387 -1318 0 1
rlabel polysilicon 387 -1324 387 -1324 0 3
rlabel polysilicon 394 -1318 394 -1318 0 1
rlabel polysilicon 394 -1324 394 -1324 0 3
rlabel polysilicon 401 -1318 401 -1318 0 1
rlabel polysilicon 401 -1324 401 -1324 0 3
rlabel polysilicon 408 -1318 408 -1318 0 1
rlabel polysilicon 408 -1324 408 -1324 0 3
rlabel polysilicon 415 -1318 415 -1318 0 1
rlabel polysilicon 415 -1324 415 -1324 0 3
rlabel polysilicon 422 -1318 422 -1318 0 1
rlabel polysilicon 425 -1318 425 -1318 0 2
rlabel polysilicon 422 -1324 422 -1324 0 3
rlabel polysilicon 429 -1318 429 -1318 0 1
rlabel polysilicon 429 -1324 429 -1324 0 3
rlabel polysilicon 436 -1318 436 -1318 0 1
rlabel polysilicon 436 -1324 436 -1324 0 3
rlabel polysilicon 443 -1318 443 -1318 0 1
rlabel polysilicon 443 -1324 443 -1324 0 3
rlabel polysilicon 450 -1318 450 -1318 0 1
rlabel polysilicon 450 -1324 450 -1324 0 3
rlabel polysilicon 460 -1318 460 -1318 0 2
rlabel polysilicon 457 -1324 457 -1324 0 3
rlabel polysilicon 460 -1324 460 -1324 0 4
rlabel polysilicon 464 -1318 464 -1318 0 1
rlabel polysilicon 464 -1324 464 -1324 0 3
rlabel polysilicon 471 -1318 471 -1318 0 1
rlabel polysilicon 471 -1324 471 -1324 0 3
rlabel polysilicon 478 -1318 478 -1318 0 1
rlabel polysilicon 481 -1318 481 -1318 0 2
rlabel polysilicon 478 -1324 478 -1324 0 3
rlabel polysilicon 485 -1318 485 -1318 0 1
rlabel polysilicon 485 -1324 485 -1324 0 3
rlabel polysilicon 492 -1318 492 -1318 0 1
rlabel polysilicon 492 -1324 492 -1324 0 3
rlabel polysilicon 499 -1318 499 -1318 0 1
rlabel polysilicon 499 -1324 499 -1324 0 3
rlabel polysilicon 506 -1318 506 -1318 0 1
rlabel polysilicon 509 -1318 509 -1318 0 2
rlabel polysilicon 506 -1324 506 -1324 0 3
rlabel polysilicon 509 -1324 509 -1324 0 4
rlabel polysilicon 513 -1318 513 -1318 0 1
rlabel polysilicon 516 -1318 516 -1318 0 2
rlabel polysilicon 520 -1324 520 -1324 0 3
rlabel polysilicon 527 -1318 527 -1318 0 1
rlabel polysilicon 530 -1318 530 -1318 0 2
rlabel polysilicon 527 -1324 527 -1324 0 3
rlabel polysilicon 530 -1324 530 -1324 0 4
rlabel polysilicon 534 -1318 534 -1318 0 1
rlabel polysilicon 534 -1324 534 -1324 0 3
rlabel polysilicon 541 -1318 541 -1318 0 1
rlabel polysilicon 541 -1324 541 -1324 0 3
rlabel polysilicon 548 -1318 548 -1318 0 1
rlabel polysilicon 548 -1324 548 -1324 0 3
rlabel polysilicon 555 -1318 555 -1318 0 1
rlabel polysilicon 555 -1324 555 -1324 0 3
rlabel polysilicon 562 -1318 562 -1318 0 1
rlabel polysilicon 562 -1324 562 -1324 0 3
rlabel polysilicon 569 -1318 569 -1318 0 1
rlabel polysilicon 569 -1324 569 -1324 0 3
rlabel polysilicon 576 -1318 576 -1318 0 1
rlabel polysilicon 576 -1324 576 -1324 0 3
rlabel polysilicon 579 -1324 579 -1324 0 4
rlabel polysilicon 583 -1318 583 -1318 0 1
rlabel polysilicon 583 -1324 583 -1324 0 3
rlabel polysilicon 593 -1318 593 -1318 0 2
rlabel polysilicon 590 -1324 590 -1324 0 3
rlabel polysilicon 597 -1318 597 -1318 0 1
rlabel polysilicon 597 -1324 597 -1324 0 3
rlabel polysilicon 604 -1318 604 -1318 0 1
rlabel polysilicon 604 -1324 604 -1324 0 3
rlabel polysilicon 614 -1318 614 -1318 0 2
rlabel polysilicon 611 -1324 611 -1324 0 3
rlabel polysilicon 614 -1324 614 -1324 0 4
rlabel polysilicon 618 -1318 618 -1318 0 1
rlabel polysilicon 618 -1324 618 -1324 0 3
rlabel polysilicon 625 -1318 625 -1318 0 1
rlabel polysilicon 628 -1318 628 -1318 0 2
rlabel polysilicon 625 -1324 625 -1324 0 3
rlabel polysilicon 628 -1324 628 -1324 0 4
rlabel polysilicon 632 -1318 632 -1318 0 1
rlabel polysilicon 632 -1324 632 -1324 0 3
rlabel polysilicon 639 -1318 639 -1318 0 1
rlabel polysilicon 639 -1324 639 -1324 0 3
rlabel polysilicon 646 -1318 646 -1318 0 1
rlabel polysilicon 646 -1324 646 -1324 0 3
rlabel polysilicon 653 -1318 653 -1318 0 1
rlabel polysilicon 653 -1324 653 -1324 0 3
rlabel polysilicon 660 -1318 660 -1318 0 1
rlabel polysilicon 660 -1324 660 -1324 0 3
rlabel polysilicon 663 -1324 663 -1324 0 4
rlabel polysilicon 667 -1318 667 -1318 0 1
rlabel polysilicon 667 -1324 667 -1324 0 3
rlabel polysilicon 674 -1318 674 -1318 0 1
rlabel polysilicon 674 -1324 674 -1324 0 3
rlabel polysilicon 681 -1318 681 -1318 0 1
rlabel polysilicon 681 -1324 681 -1324 0 3
rlabel polysilicon 688 -1318 688 -1318 0 1
rlabel polysilicon 691 -1318 691 -1318 0 2
rlabel polysilicon 688 -1324 688 -1324 0 3
rlabel polysilicon 691 -1324 691 -1324 0 4
rlabel polysilicon 695 -1318 695 -1318 0 1
rlabel polysilicon 695 -1324 695 -1324 0 3
rlabel polysilicon 702 -1318 702 -1318 0 1
rlabel polysilicon 702 -1324 702 -1324 0 3
rlabel polysilicon 709 -1318 709 -1318 0 1
rlabel polysilicon 709 -1324 709 -1324 0 3
rlabel polysilicon 716 -1318 716 -1318 0 1
rlabel polysilicon 716 -1324 716 -1324 0 3
rlabel polysilicon 723 -1318 723 -1318 0 1
rlabel polysilicon 723 -1324 723 -1324 0 3
rlabel polysilicon 730 -1318 730 -1318 0 1
rlabel polysilicon 730 -1324 730 -1324 0 3
rlabel polysilicon 737 -1318 737 -1318 0 1
rlabel polysilicon 737 -1324 737 -1324 0 3
rlabel polysilicon 744 -1318 744 -1318 0 1
rlabel polysilicon 744 -1324 744 -1324 0 3
rlabel polysilicon 751 -1318 751 -1318 0 1
rlabel polysilicon 751 -1324 751 -1324 0 3
rlabel polysilicon 758 -1318 758 -1318 0 1
rlabel polysilicon 758 -1324 758 -1324 0 3
rlabel polysilicon 765 -1318 765 -1318 0 1
rlabel polysilicon 768 -1318 768 -1318 0 2
rlabel polysilicon 765 -1324 765 -1324 0 3
rlabel polysilicon 768 -1324 768 -1324 0 4
rlabel polysilicon 772 -1318 772 -1318 0 1
rlabel polysilicon 772 -1324 772 -1324 0 3
rlabel polysilicon 779 -1318 779 -1318 0 1
rlabel polysilicon 779 -1324 779 -1324 0 3
rlabel polysilicon 786 -1318 786 -1318 0 1
rlabel polysilicon 786 -1324 786 -1324 0 3
rlabel polysilicon 789 -1324 789 -1324 0 4
rlabel polysilicon 793 -1324 793 -1324 0 3
rlabel polysilicon 796 -1324 796 -1324 0 4
rlabel polysilicon 800 -1318 800 -1318 0 1
rlabel polysilicon 800 -1324 800 -1324 0 3
rlabel polysilicon 807 -1318 807 -1318 0 1
rlabel polysilicon 810 -1318 810 -1318 0 2
rlabel polysilicon 814 -1318 814 -1318 0 1
rlabel polysilicon 817 -1318 817 -1318 0 2
rlabel polysilicon 814 -1324 814 -1324 0 3
rlabel polysilicon 817 -1324 817 -1324 0 4
rlabel polysilicon 821 -1318 821 -1318 0 1
rlabel polysilicon 821 -1324 821 -1324 0 3
rlabel polysilicon 824 -1324 824 -1324 0 4
rlabel polysilicon 828 -1318 828 -1318 0 1
rlabel polysilicon 831 -1318 831 -1318 0 2
rlabel polysilicon 828 -1324 828 -1324 0 3
rlabel polysilicon 831 -1324 831 -1324 0 4
rlabel polysilicon 835 -1318 835 -1318 0 1
rlabel polysilicon 835 -1324 835 -1324 0 3
rlabel polysilicon 842 -1318 842 -1318 0 1
rlabel polysilicon 842 -1324 842 -1324 0 3
rlabel polysilicon 849 -1318 849 -1318 0 1
rlabel polysilicon 849 -1324 849 -1324 0 3
rlabel polysilicon 856 -1318 856 -1318 0 1
rlabel polysilicon 856 -1324 856 -1324 0 3
rlabel polysilicon 863 -1318 863 -1318 0 1
rlabel polysilicon 863 -1324 863 -1324 0 3
rlabel polysilicon 870 -1318 870 -1318 0 1
rlabel polysilicon 870 -1324 870 -1324 0 3
rlabel polysilicon 877 -1318 877 -1318 0 1
rlabel polysilicon 877 -1324 877 -1324 0 3
rlabel polysilicon 884 -1318 884 -1318 0 1
rlabel polysilicon 884 -1324 884 -1324 0 3
rlabel polysilicon 891 -1318 891 -1318 0 1
rlabel polysilicon 891 -1324 891 -1324 0 3
rlabel polysilicon 898 -1318 898 -1318 0 1
rlabel polysilicon 898 -1324 898 -1324 0 3
rlabel polysilicon 905 -1318 905 -1318 0 1
rlabel polysilicon 905 -1324 905 -1324 0 3
rlabel polysilicon 912 -1318 912 -1318 0 1
rlabel polysilicon 912 -1324 912 -1324 0 3
rlabel polysilicon 919 -1318 919 -1318 0 1
rlabel polysilicon 919 -1324 919 -1324 0 3
rlabel polysilicon 926 -1318 926 -1318 0 1
rlabel polysilicon 926 -1324 926 -1324 0 3
rlabel polysilicon 933 -1318 933 -1318 0 1
rlabel polysilicon 936 -1318 936 -1318 0 2
rlabel polysilicon 933 -1324 933 -1324 0 3
rlabel polysilicon 936 -1324 936 -1324 0 4
rlabel polysilicon 940 -1318 940 -1318 0 1
rlabel polysilicon 940 -1324 940 -1324 0 3
rlabel polysilicon 947 -1318 947 -1318 0 1
rlabel polysilicon 950 -1318 950 -1318 0 2
rlabel polysilicon 947 -1324 947 -1324 0 3
rlabel polysilicon 954 -1318 954 -1318 0 1
rlabel polysilicon 954 -1324 954 -1324 0 3
rlabel polysilicon 961 -1318 961 -1318 0 1
rlabel polysilicon 961 -1324 961 -1324 0 3
rlabel polysilicon 968 -1318 968 -1318 0 1
rlabel polysilicon 968 -1324 968 -1324 0 3
rlabel polysilicon 975 -1318 975 -1318 0 1
rlabel polysilicon 978 -1318 978 -1318 0 2
rlabel polysilicon 975 -1324 975 -1324 0 3
rlabel polysilicon 978 -1324 978 -1324 0 4
rlabel polysilicon 982 -1318 982 -1318 0 1
rlabel polysilicon 985 -1318 985 -1318 0 2
rlabel polysilicon 982 -1324 982 -1324 0 3
rlabel polysilicon 985 -1324 985 -1324 0 4
rlabel polysilicon 989 -1318 989 -1318 0 1
rlabel polysilicon 989 -1324 989 -1324 0 3
rlabel polysilicon 996 -1318 996 -1318 0 1
rlabel polysilicon 999 -1318 999 -1318 0 2
rlabel polysilicon 996 -1324 996 -1324 0 3
rlabel polysilicon 1003 -1318 1003 -1318 0 1
rlabel polysilicon 1003 -1324 1003 -1324 0 3
rlabel polysilicon 1010 -1318 1010 -1318 0 1
rlabel polysilicon 1013 -1318 1013 -1318 0 2
rlabel polysilicon 1010 -1324 1010 -1324 0 3
rlabel polysilicon 1013 -1324 1013 -1324 0 4
rlabel polysilicon 1017 -1318 1017 -1318 0 1
rlabel polysilicon 1017 -1324 1017 -1324 0 3
rlabel polysilicon 1024 -1318 1024 -1318 0 1
rlabel polysilicon 1024 -1324 1024 -1324 0 3
rlabel polysilicon 1031 -1318 1031 -1318 0 1
rlabel polysilicon 1031 -1324 1031 -1324 0 3
rlabel polysilicon 1038 -1318 1038 -1318 0 1
rlabel polysilicon 1038 -1324 1038 -1324 0 3
rlabel polysilicon 1045 -1318 1045 -1318 0 1
rlabel polysilicon 1045 -1324 1045 -1324 0 3
rlabel polysilicon 1052 -1318 1052 -1318 0 1
rlabel polysilicon 1055 -1318 1055 -1318 0 2
rlabel polysilicon 1052 -1324 1052 -1324 0 3
rlabel polysilicon 1055 -1324 1055 -1324 0 4
rlabel polysilicon 1059 -1318 1059 -1318 0 1
rlabel polysilicon 1059 -1324 1059 -1324 0 3
rlabel polysilicon 1066 -1318 1066 -1318 0 1
rlabel polysilicon 1066 -1324 1066 -1324 0 3
rlabel polysilicon 1073 -1318 1073 -1318 0 1
rlabel polysilicon 1073 -1324 1073 -1324 0 3
rlabel polysilicon 1080 -1318 1080 -1318 0 1
rlabel polysilicon 1080 -1324 1080 -1324 0 3
rlabel polysilicon 1087 -1318 1087 -1318 0 1
rlabel polysilicon 1087 -1324 1087 -1324 0 3
rlabel polysilicon 1094 -1318 1094 -1318 0 1
rlabel polysilicon 1094 -1324 1094 -1324 0 3
rlabel polysilicon 1101 -1318 1101 -1318 0 1
rlabel polysilicon 1101 -1324 1101 -1324 0 3
rlabel polysilicon 1108 -1318 1108 -1318 0 1
rlabel polysilicon 1108 -1324 1108 -1324 0 3
rlabel polysilicon 1115 -1318 1115 -1318 0 1
rlabel polysilicon 1115 -1324 1115 -1324 0 3
rlabel polysilicon 1122 -1318 1122 -1318 0 1
rlabel polysilicon 1122 -1324 1122 -1324 0 3
rlabel polysilicon 1129 -1318 1129 -1318 0 1
rlabel polysilicon 1129 -1324 1129 -1324 0 3
rlabel polysilicon 1136 -1318 1136 -1318 0 1
rlabel polysilicon 1136 -1324 1136 -1324 0 3
rlabel polysilicon 1143 -1318 1143 -1318 0 1
rlabel polysilicon 1143 -1324 1143 -1324 0 3
rlabel polysilicon 1150 -1318 1150 -1318 0 1
rlabel polysilicon 1150 -1324 1150 -1324 0 3
rlabel polysilicon 1157 -1318 1157 -1318 0 1
rlabel polysilicon 1157 -1324 1157 -1324 0 3
rlabel polysilicon 1164 -1318 1164 -1318 0 1
rlabel polysilicon 1164 -1324 1164 -1324 0 3
rlabel polysilicon 1171 -1318 1171 -1318 0 1
rlabel polysilicon 1171 -1324 1171 -1324 0 3
rlabel polysilicon 1178 -1318 1178 -1318 0 1
rlabel polysilicon 1178 -1324 1178 -1324 0 3
rlabel polysilicon 1185 -1318 1185 -1318 0 1
rlabel polysilicon 1185 -1324 1185 -1324 0 3
rlabel polysilicon 1192 -1318 1192 -1318 0 1
rlabel polysilicon 1192 -1324 1192 -1324 0 3
rlabel polysilicon 1199 -1318 1199 -1318 0 1
rlabel polysilicon 1199 -1324 1199 -1324 0 3
rlabel polysilicon 1206 -1318 1206 -1318 0 1
rlabel polysilicon 1206 -1324 1206 -1324 0 3
rlabel polysilicon 1213 -1318 1213 -1318 0 1
rlabel polysilicon 1213 -1324 1213 -1324 0 3
rlabel polysilicon 1220 -1318 1220 -1318 0 1
rlabel polysilicon 1220 -1324 1220 -1324 0 3
rlabel polysilicon 1227 -1318 1227 -1318 0 1
rlabel polysilicon 1227 -1324 1227 -1324 0 3
rlabel polysilicon 1234 -1318 1234 -1318 0 1
rlabel polysilicon 1234 -1324 1234 -1324 0 3
rlabel polysilicon 1241 -1318 1241 -1318 0 1
rlabel polysilicon 1241 -1324 1241 -1324 0 3
rlabel polysilicon 1248 -1318 1248 -1318 0 1
rlabel polysilicon 1248 -1324 1248 -1324 0 3
rlabel polysilicon 1255 -1318 1255 -1318 0 1
rlabel polysilicon 1255 -1324 1255 -1324 0 3
rlabel polysilicon 1262 -1318 1262 -1318 0 1
rlabel polysilicon 1262 -1324 1262 -1324 0 3
rlabel polysilicon 1269 -1318 1269 -1318 0 1
rlabel polysilicon 1269 -1324 1269 -1324 0 3
rlabel polysilicon 1276 -1318 1276 -1318 0 1
rlabel polysilicon 1276 -1324 1276 -1324 0 3
rlabel polysilicon 1283 -1318 1283 -1318 0 1
rlabel polysilicon 1283 -1324 1283 -1324 0 3
rlabel polysilicon 1290 -1318 1290 -1318 0 1
rlabel polysilicon 1290 -1324 1290 -1324 0 3
rlabel polysilicon 1297 -1318 1297 -1318 0 1
rlabel polysilicon 1297 -1324 1297 -1324 0 3
rlabel polysilicon 1304 -1318 1304 -1318 0 1
rlabel polysilicon 1304 -1324 1304 -1324 0 3
rlabel polysilicon 1311 -1318 1311 -1318 0 1
rlabel polysilicon 1311 -1324 1311 -1324 0 3
rlabel polysilicon 1318 -1318 1318 -1318 0 1
rlabel polysilicon 1318 -1324 1318 -1324 0 3
rlabel polysilicon 1325 -1318 1325 -1318 0 1
rlabel polysilicon 1325 -1324 1325 -1324 0 3
rlabel polysilicon 1332 -1318 1332 -1318 0 1
rlabel polysilicon 1332 -1324 1332 -1324 0 3
rlabel polysilicon 1339 -1318 1339 -1318 0 1
rlabel polysilicon 1339 -1324 1339 -1324 0 3
rlabel polysilicon 1346 -1318 1346 -1318 0 1
rlabel polysilicon 1346 -1324 1346 -1324 0 3
rlabel polysilicon 1353 -1318 1353 -1318 0 1
rlabel polysilicon 1356 -1318 1356 -1318 0 2
rlabel polysilicon 1353 -1324 1353 -1324 0 3
rlabel polysilicon 1360 -1318 1360 -1318 0 1
rlabel polysilicon 1360 -1324 1360 -1324 0 3
rlabel polysilicon 1367 -1318 1367 -1318 0 1
rlabel polysilicon 1367 -1324 1367 -1324 0 3
rlabel polysilicon 1374 -1318 1374 -1318 0 1
rlabel polysilicon 1374 -1324 1374 -1324 0 3
rlabel polysilicon 1381 -1318 1381 -1318 0 1
rlabel polysilicon 1381 -1324 1381 -1324 0 3
rlabel polysilicon 1388 -1318 1388 -1318 0 1
rlabel polysilicon 1388 -1324 1388 -1324 0 3
rlabel polysilicon 1395 -1318 1395 -1318 0 1
rlabel polysilicon 1395 -1324 1395 -1324 0 3
rlabel polysilicon 1402 -1318 1402 -1318 0 1
rlabel polysilicon 1402 -1324 1402 -1324 0 3
rlabel polysilicon 1409 -1318 1409 -1318 0 1
rlabel polysilicon 1409 -1324 1409 -1324 0 3
rlabel polysilicon 1416 -1318 1416 -1318 0 1
rlabel polysilicon 1416 -1324 1416 -1324 0 3
rlabel polysilicon 1423 -1318 1423 -1318 0 1
rlabel polysilicon 1423 -1324 1423 -1324 0 3
rlabel polysilicon 1430 -1318 1430 -1318 0 1
rlabel polysilicon 1430 -1324 1430 -1324 0 3
rlabel polysilicon 1437 -1318 1437 -1318 0 1
rlabel polysilicon 1437 -1324 1437 -1324 0 3
rlabel polysilicon 1444 -1318 1444 -1318 0 1
rlabel polysilicon 1444 -1324 1444 -1324 0 3
rlabel polysilicon 1451 -1318 1451 -1318 0 1
rlabel polysilicon 1451 -1324 1451 -1324 0 3
rlabel polysilicon 1458 -1318 1458 -1318 0 1
rlabel polysilicon 1458 -1324 1458 -1324 0 3
rlabel polysilicon 1465 -1318 1465 -1318 0 1
rlabel polysilicon 1465 -1324 1465 -1324 0 3
rlabel polysilicon 1472 -1318 1472 -1318 0 1
rlabel polysilicon 1472 -1324 1472 -1324 0 3
rlabel polysilicon 1479 -1318 1479 -1318 0 1
rlabel polysilicon 1479 -1324 1479 -1324 0 3
rlabel polysilicon 1486 -1318 1486 -1318 0 1
rlabel polysilicon 1486 -1324 1486 -1324 0 3
rlabel polysilicon 1493 -1318 1493 -1318 0 1
rlabel polysilicon 1493 -1324 1493 -1324 0 3
rlabel polysilicon 1500 -1318 1500 -1318 0 1
rlabel polysilicon 1500 -1324 1500 -1324 0 3
rlabel polysilicon 1507 -1318 1507 -1318 0 1
rlabel polysilicon 1507 -1324 1507 -1324 0 3
rlabel polysilicon 1514 -1318 1514 -1318 0 1
rlabel polysilicon 1514 -1324 1514 -1324 0 3
rlabel polysilicon 1521 -1318 1521 -1318 0 1
rlabel polysilicon 1521 -1324 1521 -1324 0 3
rlabel polysilicon 1528 -1318 1528 -1318 0 1
rlabel polysilicon 1528 -1324 1528 -1324 0 3
rlabel polysilicon 1535 -1318 1535 -1318 0 1
rlabel polysilicon 1535 -1324 1535 -1324 0 3
rlabel polysilicon 1542 -1318 1542 -1318 0 1
rlabel polysilicon 1542 -1324 1542 -1324 0 3
rlabel polysilicon 1549 -1318 1549 -1318 0 1
rlabel polysilicon 1549 -1324 1549 -1324 0 3
rlabel polysilicon 1556 -1318 1556 -1318 0 1
rlabel polysilicon 1556 -1324 1556 -1324 0 3
rlabel polysilicon 1563 -1318 1563 -1318 0 1
rlabel polysilicon 1563 -1324 1563 -1324 0 3
rlabel polysilicon 1570 -1318 1570 -1318 0 1
rlabel polysilicon 1570 -1324 1570 -1324 0 3
rlabel polysilicon 1577 -1318 1577 -1318 0 1
rlabel polysilicon 1577 -1324 1577 -1324 0 3
rlabel polysilicon 1584 -1318 1584 -1318 0 1
rlabel polysilicon 1584 -1324 1584 -1324 0 3
rlabel polysilicon 1591 -1318 1591 -1318 0 1
rlabel polysilicon 1591 -1324 1591 -1324 0 3
rlabel polysilicon 1598 -1318 1598 -1318 0 1
rlabel polysilicon 1598 -1324 1598 -1324 0 3
rlabel polysilicon 1605 -1318 1605 -1318 0 1
rlabel polysilicon 1605 -1324 1605 -1324 0 3
rlabel polysilicon 1612 -1318 1612 -1318 0 1
rlabel polysilicon 1612 -1324 1612 -1324 0 3
rlabel polysilicon 1619 -1318 1619 -1318 0 1
rlabel polysilicon 1619 -1324 1619 -1324 0 3
rlabel polysilicon 1626 -1318 1626 -1318 0 1
rlabel polysilicon 1626 -1324 1626 -1324 0 3
rlabel polysilicon 1633 -1318 1633 -1318 0 1
rlabel polysilicon 1633 -1324 1633 -1324 0 3
rlabel polysilicon 1640 -1318 1640 -1318 0 1
rlabel polysilicon 1640 -1324 1640 -1324 0 3
rlabel polysilicon 1647 -1318 1647 -1318 0 1
rlabel polysilicon 1647 -1324 1647 -1324 0 3
rlabel polysilicon 1654 -1318 1654 -1318 0 1
rlabel polysilicon 1654 -1324 1654 -1324 0 3
rlabel polysilicon 1661 -1318 1661 -1318 0 1
rlabel polysilicon 1661 -1324 1661 -1324 0 3
rlabel polysilicon 1668 -1318 1668 -1318 0 1
rlabel polysilicon 1668 -1324 1668 -1324 0 3
rlabel polysilicon 1675 -1318 1675 -1318 0 1
rlabel polysilicon 1675 -1324 1675 -1324 0 3
rlabel polysilicon 1682 -1318 1682 -1318 0 1
rlabel polysilicon 1682 -1324 1682 -1324 0 3
rlabel polysilicon 1689 -1318 1689 -1318 0 1
rlabel polysilicon 1689 -1324 1689 -1324 0 3
rlabel polysilicon 1696 -1318 1696 -1318 0 1
rlabel polysilicon 1696 -1324 1696 -1324 0 3
rlabel polysilicon 1706 -1324 1706 -1324 0 4
rlabel polysilicon 1713 -1318 1713 -1318 0 2
rlabel polysilicon 1717 -1318 1717 -1318 0 1
rlabel polysilicon 1717 -1324 1717 -1324 0 3
rlabel polysilicon 1724 -1318 1724 -1318 0 1
rlabel polysilicon 1724 -1324 1724 -1324 0 3
rlabel polysilicon 1731 -1318 1731 -1318 0 1
rlabel polysilicon 1734 -1318 1734 -1318 0 2
rlabel polysilicon 1731 -1324 1731 -1324 0 3
rlabel polysilicon 1734 -1324 1734 -1324 0 4
rlabel polysilicon 1738 -1318 1738 -1318 0 1
rlabel polysilicon 1738 -1324 1738 -1324 0 3
rlabel polysilicon 16 -1473 16 -1473 0 1
rlabel polysilicon 16 -1479 16 -1479 0 3
rlabel polysilicon 26 -1473 26 -1473 0 2
rlabel polysilicon 30 -1473 30 -1473 0 1
rlabel polysilicon 30 -1479 30 -1479 0 3
rlabel polysilicon 37 -1473 37 -1473 0 1
rlabel polysilicon 37 -1479 37 -1479 0 3
rlabel polysilicon 44 -1473 44 -1473 0 1
rlabel polysilicon 44 -1479 44 -1479 0 3
rlabel polysilicon 51 -1473 51 -1473 0 1
rlabel polysilicon 51 -1479 51 -1479 0 3
rlabel polysilicon 58 -1473 58 -1473 0 1
rlabel polysilicon 61 -1473 61 -1473 0 2
rlabel polysilicon 65 -1473 65 -1473 0 1
rlabel polysilicon 65 -1479 65 -1479 0 3
rlabel polysilicon 75 -1473 75 -1473 0 2
rlabel polysilicon 72 -1479 72 -1479 0 3
rlabel polysilicon 75 -1479 75 -1479 0 4
rlabel polysilicon 79 -1473 79 -1473 0 1
rlabel polysilicon 82 -1473 82 -1473 0 2
rlabel polysilicon 79 -1479 79 -1479 0 3
rlabel polysilicon 82 -1479 82 -1479 0 4
rlabel polysilicon 86 -1473 86 -1473 0 1
rlabel polysilicon 86 -1479 86 -1479 0 3
rlabel polysilicon 93 -1473 93 -1473 0 1
rlabel polysilicon 96 -1473 96 -1473 0 2
rlabel polysilicon 93 -1479 93 -1479 0 3
rlabel polysilicon 100 -1473 100 -1473 0 1
rlabel polysilicon 100 -1479 100 -1479 0 3
rlabel polysilicon 107 -1473 107 -1473 0 1
rlabel polysilicon 110 -1473 110 -1473 0 2
rlabel polysilicon 107 -1479 107 -1479 0 3
rlabel polysilicon 117 -1473 117 -1473 0 2
rlabel polysilicon 114 -1479 114 -1479 0 3
rlabel polysilicon 117 -1479 117 -1479 0 4
rlabel polysilicon 121 -1473 121 -1473 0 1
rlabel polysilicon 121 -1479 121 -1479 0 3
rlabel polysilicon 128 -1473 128 -1473 0 1
rlabel polysilicon 128 -1479 128 -1479 0 3
rlabel polysilicon 135 -1473 135 -1473 0 1
rlabel polysilicon 135 -1479 135 -1479 0 3
rlabel polysilicon 142 -1473 142 -1473 0 1
rlabel polysilicon 142 -1479 142 -1479 0 3
rlabel polysilicon 149 -1473 149 -1473 0 1
rlabel polysilicon 149 -1479 149 -1479 0 3
rlabel polysilicon 156 -1473 156 -1473 0 1
rlabel polysilicon 156 -1479 156 -1479 0 3
rlabel polysilicon 159 -1479 159 -1479 0 4
rlabel polysilicon 163 -1473 163 -1473 0 1
rlabel polysilicon 163 -1479 163 -1479 0 3
rlabel polysilicon 170 -1473 170 -1473 0 1
rlabel polysilicon 170 -1479 170 -1479 0 3
rlabel polysilicon 177 -1473 177 -1473 0 1
rlabel polysilicon 177 -1479 177 -1479 0 3
rlabel polysilicon 184 -1473 184 -1473 0 1
rlabel polysilicon 184 -1479 184 -1479 0 3
rlabel polysilicon 191 -1473 191 -1473 0 1
rlabel polysilicon 191 -1479 191 -1479 0 3
rlabel polysilicon 198 -1473 198 -1473 0 1
rlabel polysilicon 198 -1479 198 -1479 0 3
rlabel polysilicon 205 -1473 205 -1473 0 1
rlabel polysilicon 205 -1479 205 -1479 0 3
rlabel polysilicon 212 -1473 212 -1473 0 1
rlabel polysilicon 212 -1479 212 -1479 0 3
rlabel polysilicon 219 -1473 219 -1473 0 1
rlabel polysilicon 222 -1473 222 -1473 0 2
rlabel polysilicon 219 -1479 219 -1479 0 3
rlabel polysilicon 226 -1473 226 -1473 0 1
rlabel polysilicon 229 -1473 229 -1473 0 2
rlabel polysilicon 226 -1479 226 -1479 0 3
rlabel polysilicon 229 -1479 229 -1479 0 4
rlabel polysilicon 233 -1473 233 -1473 0 1
rlabel polysilicon 233 -1479 233 -1479 0 3
rlabel polysilicon 240 -1473 240 -1473 0 1
rlabel polysilicon 240 -1479 240 -1479 0 3
rlabel polysilicon 247 -1473 247 -1473 0 1
rlabel polysilicon 247 -1479 247 -1479 0 3
rlabel polysilicon 254 -1473 254 -1473 0 1
rlabel polysilicon 254 -1479 254 -1479 0 3
rlabel polysilicon 261 -1473 261 -1473 0 1
rlabel polysilicon 264 -1473 264 -1473 0 2
rlabel polysilicon 264 -1479 264 -1479 0 4
rlabel polysilicon 268 -1473 268 -1473 0 1
rlabel polysilicon 268 -1479 268 -1479 0 3
rlabel polysilicon 275 -1473 275 -1473 0 1
rlabel polysilicon 275 -1479 275 -1479 0 3
rlabel polysilicon 282 -1473 282 -1473 0 1
rlabel polysilicon 282 -1479 282 -1479 0 3
rlabel polysilicon 289 -1473 289 -1473 0 1
rlabel polysilicon 289 -1479 289 -1479 0 3
rlabel polysilicon 299 -1479 299 -1479 0 4
rlabel polysilicon 303 -1473 303 -1473 0 1
rlabel polysilicon 303 -1479 303 -1479 0 3
rlabel polysilicon 310 -1473 310 -1473 0 1
rlabel polysilicon 310 -1479 310 -1479 0 3
rlabel polysilicon 317 -1473 317 -1473 0 1
rlabel polysilicon 317 -1479 317 -1479 0 3
rlabel polysilicon 324 -1473 324 -1473 0 1
rlabel polysilicon 324 -1479 324 -1479 0 3
rlabel polysilicon 331 -1473 331 -1473 0 1
rlabel polysilicon 331 -1479 331 -1479 0 3
rlabel polysilicon 338 -1473 338 -1473 0 1
rlabel polysilicon 338 -1479 338 -1479 0 3
rlabel polysilicon 345 -1473 345 -1473 0 1
rlabel polysilicon 345 -1479 345 -1479 0 3
rlabel polysilicon 352 -1473 352 -1473 0 1
rlabel polysilicon 352 -1479 352 -1479 0 3
rlabel polysilicon 359 -1473 359 -1473 0 1
rlabel polysilicon 359 -1479 359 -1479 0 3
rlabel polysilicon 366 -1473 366 -1473 0 1
rlabel polysilicon 366 -1479 366 -1479 0 3
rlabel polysilicon 373 -1473 373 -1473 0 1
rlabel polysilicon 373 -1479 373 -1479 0 3
rlabel polysilicon 380 -1473 380 -1473 0 1
rlabel polysilicon 380 -1479 380 -1479 0 3
rlabel polysilicon 387 -1473 387 -1473 0 1
rlabel polysilicon 387 -1479 387 -1479 0 3
rlabel polysilicon 390 -1479 390 -1479 0 4
rlabel polysilicon 394 -1473 394 -1473 0 1
rlabel polysilicon 394 -1479 394 -1479 0 3
rlabel polysilicon 401 -1473 401 -1473 0 1
rlabel polysilicon 401 -1479 401 -1479 0 3
rlabel polysilicon 408 -1473 408 -1473 0 1
rlabel polysilicon 408 -1479 408 -1479 0 3
rlabel polysilicon 411 -1479 411 -1479 0 4
rlabel polysilicon 415 -1473 415 -1473 0 1
rlabel polysilicon 418 -1473 418 -1473 0 2
rlabel polysilicon 415 -1479 415 -1479 0 3
rlabel polysilicon 418 -1479 418 -1479 0 4
rlabel polysilicon 422 -1473 422 -1473 0 1
rlabel polysilicon 422 -1479 422 -1479 0 3
rlabel polysilicon 429 -1473 429 -1473 0 1
rlabel polysilicon 429 -1479 429 -1479 0 3
rlabel polysilicon 436 -1473 436 -1473 0 1
rlabel polysilicon 436 -1479 436 -1479 0 3
rlabel polysilicon 443 -1473 443 -1473 0 1
rlabel polysilicon 443 -1479 443 -1479 0 3
rlabel polysilicon 450 -1473 450 -1473 0 1
rlabel polysilicon 450 -1479 450 -1479 0 3
rlabel polysilicon 457 -1473 457 -1473 0 1
rlabel polysilicon 457 -1479 457 -1479 0 3
rlabel polysilicon 464 -1473 464 -1473 0 1
rlabel polysilicon 464 -1479 464 -1479 0 3
rlabel polysilicon 471 -1473 471 -1473 0 1
rlabel polysilicon 471 -1479 471 -1479 0 3
rlabel polysilicon 478 -1473 478 -1473 0 1
rlabel polysilicon 478 -1479 478 -1479 0 3
rlabel polysilicon 485 -1473 485 -1473 0 1
rlabel polysilicon 485 -1479 485 -1479 0 3
rlabel polysilicon 492 -1473 492 -1473 0 1
rlabel polysilicon 492 -1479 492 -1479 0 3
rlabel polysilicon 499 -1473 499 -1473 0 1
rlabel polysilicon 502 -1473 502 -1473 0 2
rlabel polysilicon 502 -1479 502 -1479 0 4
rlabel polysilicon 506 -1473 506 -1473 0 1
rlabel polysilicon 506 -1479 506 -1479 0 3
rlabel polysilicon 513 -1473 513 -1473 0 1
rlabel polysilicon 513 -1479 513 -1479 0 3
rlabel polysilicon 520 -1473 520 -1473 0 1
rlabel polysilicon 520 -1479 520 -1479 0 3
rlabel polysilicon 527 -1473 527 -1473 0 1
rlabel polysilicon 527 -1479 527 -1479 0 3
rlabel polysilicon 534 -1473 534 -1473 0 1
rlabel polysilicon 534 -1479 534 -1479 0 3
rlabel polysilicon 541 -1473 541 -1473 0 1
rlabel polysilicon 541 -1479 541 -1479 0 3
rlabel polysilicon 548 -1473 548 -1473 0 1
rlabel polysilicon 548 -1479 548 -1479 0 3
rlabel polysilicon 555 -1473 555 -1473 0 1
rlabel polysilicon 555 -1479 555 -1479 0 3
rlabel polysilicon 558 -1479 558 -1479 0 4
rlabel polysilicon 562 -1473 562 -1473 0 1
rlabel polysilicon 562 -1479 562 -1479 0 3
rlabel polysilicon 569 -1473 569 -1473 0 1
rlabel polysilicon 569 -1479 569 -1479 0 3
rlabel polysilicon 576 -1473 576 -1473 0 1
rlabel polysilicon 576 -1479 576 -1479 0 3
rlabel polysilicon 583 -1473 583 -1473 0 1
rlabel polysilicon 583 -1479 583 -1479 0 3
rlabel polysilicon 590 -1473 590 -1473 0 1
rlabel polysilicon 593 -1473 593 -1473 0 2
rlabel polysilicon 590 -1479 590 -1479 0 3
rlabel polysilicon 593 -1479 593 -1479 0 4
rlabel polysilicon 597 -1473 597 -1473 0 1
rlabel polysilicon 600 -1473 600 -1473 0 2
rlabel polysilicon 597 -1479 597 -1479 0 3
rlabel polysilicon 604 -1473 604 -1473 0 1
rlabel polysilicon 604 -1479 604 -1479 0 3
rlabel polysilicon 611 -1473 611 -1473 0 1
rlabel polysilicon 614 -1473 614 -1473 0 2
rlabel polysilicon 614 -1479 614 -1479 0 4
rlabel polysilicon 618 -1473 618 -1473 0 1
rlabel polysilicon 618 -1479 618 -1479 0 3
rlabel polysilicon 625 -1473 625 -1473 0 1
rlabel polysilicon 625 -1479 625 -1479 0 3
rlabel polysilicon 632 -1473 632 -1473 0 1
rlabel polysilicon 635 -1473 635 -1473 0 2
rlabel polysilicon 632 -1479 632 -1479 0 3
rlabel polysilicon 635 -1479 635 -1479 0 4
rlabel polysilicon 639 -1473 639 -1473 0 1
rlabel polysilicon 642 -1473 642 -1473 0 2
rlabel polysilicon 639 -1479 639 -1479 0 3
rlabel polysilicon 642 -1479 642 -1479 0 4
rlabel polysilicon 646 -1473 646 -1473 0 1
rlabel polysilicon 646 -1479 646 -1479 0 3
rlabel polysilicon 653 -1473 653 -1473 0 1
rlabel polysilicon 653 -1479 653 -1479 0 3
rlabel polysilicon 660 -1473 660 -1473 0 1
rlabel polysilicon 660 -1479 660 -1479 0 3
rlabel polysilicon 667 -1473 667 -1473 0 1
rlabel polysilicon 667 -1479 667 -1479 0 3
rlabel polysilicon 674 -1473 674 -1473 0 1
rlabel polysilicon 677 -1473 677 -1473 0 2
rlabel polysilicon 674 -1479 674 -1479 0 3
rlabel polysilicon 677 -1479 677 -1479 0 4
rlabel polysilicon 681 -1473 681 -1473 0 1
rlabel polysilicon 681 -1479 681 -1479 0 3
rlabel polysilicon 688 -1473 688 -1473 0 1
rlabel polysilicon 688 -1479 688 -1479 0 3
rlabel polysilicon 695 -1473 695 -1473 0 1
rlabel polysilicon 695 -1479 695 -1479 0 3
rlabel polysilicon 702 -1473 702 -1473 0 1
rlabel polysilicon 702 -1479 702 -1479 0 3
rlabel polysilicon 709 -1473 709 -1473 0 1
rlabel polysilicon 709 -1479 709 -1479 0 3
rlabel polysilicon 716 -1473 716 -1473 0 1
rlabel polysilicon 719 -1473 719 -1473 0 2
rlabel polysilicon 716 -1479 716 -1479 0 3
rlabel polysilicon 719 -1479 719 -1479 0 4
rlabel polysilicon 723 -1473 723 -1473 0 1
rlabel polysilicon 726 -1473 726 -1473 0 2
rlabel polysilicon 723 -1479 723 -1479 0 3
rlabel polysilicon 726 -1479 726 -1479 0 4
rlabel polysilicon 730 -1473 730 -1473 0 1
rlabel polysilicon 733 -1473 733 -1473 0 2
rlabel polysilicon 730 -1479 730 -1479 0 3
rlabel polysilicon 733 -1479 733 -1479 0 4
rlabel polysilicon 737 -1473 737 -1473 0 1
rlabel polysilicon 737 -1479 737 -1479 0 3
rlabel polysilicon 744 -1473 744 -1473 0 1
rlabel polysilicon 744 -1479 744 -1479 0 3
rlabel polysilicon 751 -1473 751 -1473 0 1
rlabel polysilicon 751 -1479 751 -1479 0 3
rlabel polysilicon 758 -1473 758 -1473 0 1
rlabel polysilicon 758 -1479 758 -1479 0 3
rlabel polysilicon 765 -1473 765 -1473 0 1
rlabel polysilicon 765 -1479 765 -1479 0 3
rlabel polysilicon 768 -1479 768 -1479 0 4
rlabel polysilicon 772 -1473 772 -1473 0 1
rlabel polysilicon 772 -1479 772 -1479 0 3
rlabel polysilicon 779 -1473 779 -1473 0 1
rlabel polysilicon 779 -1479 779 -1479 0 3
rlabel polysilicon 786 -1473 786 -1473 0 1
rlabel polysilicon 786 -1479 786 -1479 0 3
rlabel polysilicon 793 -1473 793 -1473 0 1
rlabel polysilicon 793 -1479 793 -1479 0 3
rlabel polysilicon 800 -1473 800 -1473 0 1
rlabel polysilicon 800 -1479 800 -1479 0 3
rlabel polysilicon 807 -1473 807 -1473 0 1
rlabel polysilicon 807 -1479 807 -1479 0 3
rlabel polysilicon 814 -1473 814 -1473 0 1
rlabel polysilicon 814 -1479 814 -1479 0 3
rlabel polysilicon 821 -1473 821 -1473 0 1
rlabel polysilicon 821 -1479 821 -1479 0 3
rlabel polysilicon 828 -1473 828 -1473 0 1
rlabel polysilicon 828 -1479 828 -1479 0 3
rlabel polysilicon 835 -1473 835 -1473 0 1
rlabel polysilicon 835 -1479 835 -1479 0 3
rlabel polysilicon 842 -1473 842 -1473 0 1
rlabel polysilicon 842 -1479 842 -1479 0 3
rlabel polysilicon 849 -1473 849 -1473 0 1
rlabel polysilicon 849 -1479 849 -1479 0 3
rlabel polysilicon 856 -1473 856 -1473 0 1
rlabel polysilicon 856 -1479 856 -1479 0 3
rlabel polysilicon 863 -1473 863 -1473 0 1
rlabel polysilicon 866 -1473 866 -1473 0 2
rlabel polysilicon 863 -1479 863 -1479 0 3
rlabel polysilicon 866 -1479 866 -1479 0 4
rlabel polysilicon 870 -1473 870 -1473 0 1
rlabel polysilicon 873 -1473 873 -1473 0 2
rlabel polysilicon 870 -1479 870 -1479 0 3
rlabel polysilicon 873 -1479 873 -1479 0 4
rlabel polysilicon 877 -1473 877 -1473 0 1
rlabel polysilicon 877 -1479 877 -1479 0 3
rlabel polysilicon 884 -1473 884 -1473 0 1
rlabel polysilicon 884 -1479 884 -1479 0 3
rlabel polysilicon 891 -1473 891 -1473 0 1
rlabel polysilicon 894 -1473 894 -1473 0 2
rlabel polysilicon 891 -1479 891 -1479 0 3
rlabel polysilicon 898 -1473 898 -1473 0 1
rlabel polysilicon 901 -1473 901 -1473 0 2
rlabel polysilicon 901 -1479 901 -1479 0 4
rlabel polysilicon 905 -1473 905 -1473 0 1
rlabel polysilicon 905 -1479 905 -1479 0 3
rlabel polysilicon 912 -1473 912 -1473 0 1
rlabel polysilicon 912 -1479 912 -1479 0 3
rlabel polysilicon 919 -1473 919 -1473 0 1
rlabel polysilicon 919 -1479 919 -1479 0 3
rlabel polysilicon 926 -1473 926 -1473 0 1
rlabel polysilicon 926 -1479 926 -1479 0 3
rlabel polysilicon 933 -1473 933 -1473 0 1
rlabel polysilicon 936 -1473 936 -1473 0 2
rlabel polysilicon 933 -1479 933 -1479 0 3
rlabel polysilicon 936 -1479 936 -1479 0 4
rlabel polysilicon 940 -1473 940 -1473 0 1
rlabel polysilicon 940 -1479 940 -1479 0 3
rlabel polysilicon 947 -1473 947 -1473 0 1
rlabel polysilicon 947 -1479 947 -1479 0 3
rlabel polysilicon 954 -1473 954 -1473 0 1
rlabel polysilicon 954 -1479 954 -1479 0 3
rlabel polysilicon 961 -1473 961 -1473 0 1
rlabel polysilicon 961 -1479 961 -1479 0 3
rlabel polysilicon 968 -1473 968 -1473 0 1
rlabel polysilicon 968 -1479 968 -1479 0 3
rlabel polysilicon 975 -1473 975 -1473 0 1
rlabel polysilicon 975 -1479 975 -1479 0 3
rlabel polysilicon 982 -1473 982 -1473 0 1
rlabel polysilicon 982 -1479 982 -1479 0 3
rlabel polysilicon 989 -1473 989 -1473 0 1
rlabel polysilicon 989 -1479 989 -1479 0 3
rlabel polysilicon 996 -1473 996 -1473 0 1
rlabel polysilicon 996 -1479 996 -1479 0 3
rlabel polysilicon 1003 -1473 1003 -1473 0 1
rlabel polysilicon 1003 -1479 1003 -1479 0 3
rlabel polysilicon 1010 -1473 1010 -1473 0 1
rlabel polysilicon 1010 -1479 1010 -1479 0 3
rlabel polysilicon 1017 -1473 1017 -1473 0 1
rlabel polysilicon 1017 -1479 1017 -1479 0 3
rlabel polysilicon 1027 -1473 1027 -1473 0 2
rlabel polysilicon 1024 -1479 1024 -1479 0 3
rlabel polysilicon 1031 -1473 1031 -1473 0 1
rlabel polysilicon 1031 -1479 1031 -1479 0 3
rlabel polysilicon 1038 -1473 1038 -1473 0 1
rlabel polysilicon 1038 -1479 1038 -1479 0 3
rlabel polysilicon 1045 -1473 1045 -1473 0 1
rlabel polysilicon 1045 -1479 1045 -1479 0 3
rlabel polysilicon 1052 -1473 1052 -1473 0 1
rlabel polysilicon 1052 -1479 1052 -1479 0 3
rlabel polysilicon 1059 -1473 1059 -1473 0 1
rlabel polysilicon 1059 -1479 1059 -1479 0 3
rlabel polysilicon 1066 -1473 1066 -1473 0 1
rlabel polysilicon 1069 -1473 1069 -1473 0 2
rlabel polysilicon 1066 -1479 1066 -1479 0 3
rlabel polysilicon 1073 -1473 1073 -1473 0 1
rlabel polysilicon 1073 -1479 1073 -1479 0 3
rlabel polysilicon 1080 -1473 1080 -1473 0 1
rlabel polysilicon 1080 -1479 1080 -1479 0 3
rlabel polysilicon 1087 -1473 1087 -1473 0 1
rlabel polysilicon 1087 -1479 1087 -1479 0 3
rlabel polysilicon 1094 -1473 1094 -1473 0 1
rlabel polysilicon 1094 -1479 1094 -1479 0 3
rlabel polysilicon 1101 -1473 1101 -1473 0 1
rlabel polysilicon 1101 -1479 1101 -1479 0 3
rlabel polysilicon 1108 -1473 1108 -1473 0 1
rlabel polysilicon 1108 -1479 1108 -1479 0 3
rlabel polysilicon 1115 -1473 1115 -1473 0 1
rlabel polysilicon 1115 -1479 1115 -1479 0 3
rlabel polysilicon 1122 -1473 1122 -1473 0 1
rlabel polysilicon 1125 -1473 1125 -1473 0 2
rlabel polysilicon 1122 -1479 1122 -1479 0 3
rlabel polysilicon 1125 -1479 1125 -1479 0 4
rlabel polysilicon 1129 -1473 1129 -1473 0 1
rlabel polysilicon 1129 -1479 1129 -1479 0 3
rlabel polysilicon 1139 -1473 1139 -1473 0 2
rlabel polysilicon 1139 -1479 1139 -1479 0 4
rlabel polysilicon 1143 -1473 1143 -1473 0 1
rlabel polysilicon 1146 -1473 1146 -1473 0 2
rlabel polysilicon 1143 -1479 1143 -1479 0 3
rlabel polysilicon 1146 -1479 1146 -1479 0 4
rlabel polysilicon 1150 -1473 1150 -1473 0 1
rlabel polysilicon 1150 -1479 1150 -1479 0 3
rlabel polysilicon 1157 -1473 1157 -1473 0 1
rlabel polysilicon 1157 -1479 1157 -1479 0 3
rlabel polysilicon 1164 -1473 1164 -1473 0 1
rlabel polysilicon 1164 -1479 1164 -1479 0 3
rlabel polysilicon 1171 -1473 1171 -1473 0 1
rlabel polysilicon 1171 -1479 1171 -1479 0 3
rlabel polysilicon 1178 -1473 1178 -1473 0 1
rlabel polysilicon 1178 -1479 1178 -1479 0 3
rlabel polysilicon 1185 -1473 1185 -1473 0 1
rlabel polysilicon 1185 -1479 1185 -1479 0 3
rlabel polysilicon 1192 -1473 1192 -1473 0 1
rlabel polysilicon 1192 -1479 1192 -1479 0 3
rlabel polysilicon 1199 -1473 1199 -1473 0 1
rlabel polysilicon 1199 -1479 1199 -1479 0 3
rlabel polysilicon 1206 -1473 1206 -1473 0 1
rlabel polysilicon 1206 -1479 1206 -1479 0 3
rlabel polysilicon 1213 -1473 1213 -1473 0 1
rlabel polysilicon 1213 -1479 1213 -1479 0 3
rlabel polysilicon 1220 -1473 1220 -1473 0 1
rlabel polysilicon 1220 -1479 1220 -1479 0 3
rlabel polysilicon 1227 -1473 1227 -1473 0 1
rlabel polysilicon 1227 -1479 1227 -1479 0 3
rlabel polysilicon 1234 -1473 1234 -1473 0 1
rlabel polysilicon 1234 -1479 1234 -1479 0 3
rlabel polysilicon 1241 -1473 1241 -1473 0 1
rlabel polysilicon 1241 -1479 1241 -1479 0 3
rlabel polysilicon 1248 -1473 1248 -1473 0 1
rlabel polysilicon 1248 -1479 1248 -1479 0 3
rlabel polysilicon 1255 -1473 1255 -1473 0 1
rlabel polysilicon 1255 -1479 1255 -1479 0 3
rlabel polysilicon 1262 -1473 1262 -1473 0 1
rlabel polysilicon 1262 -1479 1262 -1479 0 3
rlabel polysilicon 1269 -1473 1269 -1473 0 1
rlabel polysilicon 1269 -1479 1269 -1479 0 3
rlabel polysilicon 1276 -1473 1276 -1473 0 1
rlabel polysilicon 1276 -1479 1276 -1479 0 3
rlabel polysilicon 1283 -1473 1283 -1473 0 1
rlabel polysilicon 1283 -1479 1283 -1479 0 3
rlabel polysilicon 1290 -1473 1290 -1473 0 1
rlabel polysilicon 1290 -1479 1290 -1479 0 3
rlabel polysilicon 1297 -1473 1297 -1473 0 1
rlabel polysilicon 1297 -1479 1297 -1479 0 3
rlabel polysilicon 1304 -1473 1304 -1473 0 1
rlabel polysilicon 1304 -1479 1304 -1479 0 3
rlabel polysilicon 1311 -1473 1311 -1473 0 1
rlabel polysilicon 1311 -1479 1311 -1479 0 3
rlabel polysilicon 1318 -1473 1318 -1473 0 1
rlabel polysilicon 1318 -1479 1318 -1479 0 3
rlabel polysilicon 1325 -1473 1325 -1473 0 1
rlabel polysilicon 1325 -1479 1325 -1479 0 3
rlabel polysilicon 1332 -1473 1332 -1473 0 1
rlabel polysilicon 1332 -1479 1332 -1479 0 3
rlabel polysilicon 1339 -1473 1339 -1473 0 1
rlabel polysilicon 1339 -1479 1339 -1479 0 3
rlabel polysilicon 1346 -1473 1346 -1473 0 1
rlabel polysilicon 1346 -1479 1346 -1479 0 3
rlabel polysilicon 1353 -1473 1353 -1473 0 1
rlabel polysilicon 1353 -1479 1353 -1479 0 3
rlabel polysilicon 1360 -1473 1360 -1473 0 1
rlabel polysilicon 1360 -1479 1360 -1479 0 3
rlabel polysilicon 1367 -1473 1367 -1473 0 1
rlabel polysilicon 1367 -1479 1367 -1479 0 3
rlabel polysilicon 1374 -1473 1374 -1473 0 1
rlabel polysilicon 1374 -1479 1374 -1479 0 3
rlabel polysilicon 1381 -1473 1381 -1473 0 1
rlabel polysilicon 1381 -1479 1381 -1479 0 3
rlabel polysilicon 1388 -1473 1388 -1473 0 1
rlabel polysilicon 1388 -1479 1388 -1479 0 3
rlabel polysilicon 1395 -1473 1395 -1473 0 1
rlabel polysilicon 1395 -1479 1395 -1479 0 3
rlabel polysilicon 1402 -1473 1402 -1473 0 1
rlabel polysilicon 1402 -1479 1402 -1479 0 3
rlabel polysilicon 1409 -1473 1409 -1473 0 1
rlabel polysilicon 1409 -1479 1409 -1479 0 3
rlabel polysilicon 1416 -1473 1416 -1473 0 1
rlabel polysilicon 1416 -1479 1416 -1479 0 3
rlabel polysilicon 1423 -1473 1423 -1473 0 1
rlabel polysilicon 1423 -1479 1423 -1479 0 3
rlabel polysilicon 1430 -1473 1430 -1473 0 1
rlabel polysilicon 1430 -1479 1430 -1479 0 3
rlabel polysilicon 1437 -1473 1437 -1473 0 1
rlabel polysilicon 1437 -1479 1437 -1479 0 3
rlabel polysilicon 1444 -1473 1444 -1473 0 1
rlabel polysilicon 1444 -1479 1444 -1479 0 3
rlabel polysilicon 1451 -1473 1451 -1473 0 1
rlabel polysilicon 1451 -1479 1451 -1479 0 3
rlabel polysilicon 1458 -1473 1458 -1473 0 1
rlabel polysilicon 1458 -1479 1458 -1479 0 3
rlabel polysilicon 1465 -1473 1465 -1473 0 1
rlabel polysilicon 1465 -1479 1465 -1479 0 3
rlabel polysilicon 1472 -1473 1472 -1473 0 1
rlabel polysilicon 1472 -1479 1472 -1479 0 3
rlabel polysilicon 1479 -1473 1479 -1473 0 1
rlabel polysilicon 1479 -1479 1479 -1479 0 3
rlabel polysilicon 1486 -1473 1486 -1473 0 1
rlabel polysilicon 1486 -1479 1486 -1479 0 3
rlabel polysilicon 1493 -1473 1493 -1473 0 1
rlabel polysilicon 1493 -1479 1493 -1479 0 3
rlabel polysilicon 1500 -1473 1500 -1473 0 1
rlabel polysilicon 1500 -1479 1500 -1479 0 3
rlabel polysilicon 1507 -1473 1507 -1473 0 1
rlabel polysilicon 1507 -1479 1507 -1479 0 3
rlabel polysilicon 1514 -1473 1514 -1473 0 1
rlabel polysilicon 1514 -1479 1514 -1479 0 3
rlabel polysilicon 1521 -1473 1521 -1473 0 1
rlabel polysilicon 1521 -1479 1521 -1479 0 3
rlabel polysilicon 1528 -1473 1528 -1473 0 1
rlabel polysilicon 1528 -1479 1528 -1479 0 3
rlabel polysilicon 1535 -1473 1535 -1473 0 1
rlabel polysilicon 1535 -1479 1535 -1479 0 3
rlabel polysilicon 1542 -1473 1542 -1473 0 1
rlabel polysilicon 1542 -1479 1542 -1479 0 3
rlabel polysilicon 1549 -1473 1549 -1473 0 1
rlabel polysilicon 1549 -1479 1549 -1479 0 3
rlabel polysilicon 1556 -1473 1556 -1473 0 1
rlabel polysilicon 1556 -1479 1556 -1479 0 3
rlabel polysilicon 1563 -1473 1563 -1473 0 1
rlabel polysilicon 1563 -1479 1563 -1479 0 3
rlabel polysilicon 1570 -1473 1570 -1473 0 1
rlabel polysilicon 1570 -1479 1570 -1479 0 3
rlabel polysilicon 1577 -1473 1577 -1473 0 1
rlabel polysilicon 1577 -1479 1577 -1479 0 3
rlabel polysilicon 1584 -1473 1584 -1473 0 1
rlabel polysilicon 1584 -1479 1584 -1479 0 3
rlabel polysilicon 1591 -1473 1591 -1473 0 1
rlabel polysilicon 1591 -1479 1591 -1479 0 3
rlabel polysilicon 1598 -1473 1598 -1473 0 1
rlabel polysilicon 1598 -1479 1598 -1479 0 3
rlabel polysilicon 1605 -1473 1605 -1473 0 1
rlabel polysilicon 1605 -1479 1605 -1479 0 3
rlabel polysilicon 1612 -1473 1612 -1473 0 1
rlabel polysilicon 1612 -1479 1612 -1479 0 3
rlabel polysilicon 1619 -1473 1619 -1473 0 1
rlabel polysilicon 1619 -1479 1619 -1479 0 3
rlabel polysilicon 1626 -1473 1626 -1473 0 1
rlabel polysilicon 1626 -1479 1626 -1479 0 3
rlabel polysilicon 1633 -1473 1633 -1473 0 1
rlabel polysilicon 1633 -1479 1633 -1479 0 3
rlabel polysilicon 1640 -1473 1640 -1473 0 1
rlabel polysilicon 1640 -1479 1640 -1479 0 3
rlabel polysilicon 1647 -1473 1647 -1473 0 1
rlabel polysilicon 1647 -1479 1647 -1479 0 3
rlabel polysilicon 1654 -1473 1654 -1473 0 1
rlabel polysilicon 1654 -1479 1654 -1479 0 3
rlabel polysilicon 1661 -1473 1661 -1473 0 1
rlabel polysilicon 1661 -1479 1661 -1479 0 3
rlabel polysilicon 1668 -1473 1668 -1473 0 1
rlabel polysilicon 1668 -1479 1668 -1479 0 3
rlabel polysilicon 1675 -1473 1675 -1473 0 1
rlabel polysilicon 1675 -1479 1675 -1479 0 3
rlabel polysilicon 1682 -1473 1682 -1473 0 1
rlabel polysilicon 1682 -1479 1682 -1479 0 3
rlabel polysilicon 1689 -1473 1689 -1473 0 1
rlabel polysilicon 1689 -1479 1689 -1479 0 3
rlabel polysilicon 1699 -1473 1699 -1473 0 2
rlabel polysilicon 1703 -1473 1703 -1473 0 1
rlabel polysilicon 1703 -1479 1703 -1479 0 3
rlabel polysilicon 1710 -1473 1710 -1473 0 1
rlabel polysilicon 1710 -1479 1710 -1479 0 3
rlabel polysilicon 1717 -1473 1717 -1473 0 1
rlabel polysilicon 1720 -1473 1720 -1473 0 2
rlabel polysilicon 1717 -1479 1717 -1479 0 3
rlabel polysilicon 1720 -1479 1720 -1479 0 4
rlabel polysilicon 1724 -1473 1724 -1473 0 1
rlabel polysilicon 1724 -1479 1724 -1479 0 3
rlabel polysilicon 1745 -1473 1745 -1473 0 1
rlabel polysilicon 1745 -1479 1745 -1479 0 3
rlabel polysilicon 23 -1610 23 -1610 0 1
rlabel polysilicon 23 -1616 23 -1616 0 3
rlabel polysilicon 30 -1610 30 -1610 0 1
rlabel polysilicon 30 -1616 30 -1616 0 3
rlabel polysilicon 44 -1610 44 -1610 0 1
rlabel polysilicon 44 -1616 44 -1616 0 3
rlabel polysilicon 51 -1610 51 -1610 0 1
rlabel polysilicon 51 -1616 51 -1616 0 3
rlabel polysilicon 58 -1610 58 -1610 0 1
rlabel polysilicon 61 -1610 61 -1610 0 2
rlabel polysilicon 65 -1610 65 -1610 0 1
rlabel polysilicon 68 -1610 68 -1610 0 2
rlabel polysilicon 72 -1610 72 -1610 0 1
rlabel polysilicon 72 -1616 72 -1616 0 3
rlabel polysilicon 79 -1610 79 -1610 0 1
rlabel polysilicon 79 -1616 79 -1616 0 3
rlabel polysilicon 86 -1610 86 -1610 0 1
rlabel polysilicon 86 -1616 86 -1616 0 3
rlabel polysilicon 93 -1610 93 -1610 0 1
rlabel polysilicon 96 -1610 96 -1610 0 2
rlabel polysilicon 93 -1616 93 -1616 0 3
rlabel polysilicon 96 -1616 96 -1616 0 4
rlabel polysilicon 100 -1610 100 -1610 0 1
rlabel polysilicon 100 -1616 100 -1616 0 3
rlabel polysilicon 107 -1610 107 -1610 0 1
rlabel polysilicon 107 -1616 107 -1616 0 3
rlabel polysilicon 114 -1610 114 -1610 0 1
rlabel polysilicon 114 -1616 114 -1616 0 3
rlabel polysilicon 121 -1610 121 -1610 0 1
rlabel polysilicon 121 -1616 121 -1616 0 3
rlabel polysilicon 128 -1610 128 -1610 0 1
rlabel polysilicon 128 -1616 128 -1616 0 3
rlabel polysilicon 135 -1610 135 -1610 0 1
rlabel polysilicon 135 -1616 135 -1616 0 3
rlabel polysilicon 142 -1610 142 -1610 0 1
rlabel polysilicon 142 -1616 142 -1616 0 3
rlabel polysilicon 149 -1610 149 -1610 0 1
rlabel polysilicon 149 -1616 149 -1616 0 3
rlabel polysilicon 156 -1610 156 -1610 0 1
rlabel polysilicon 156 -1616 156 -1616 0 3
rlabel polysilicon 163 -1610 163 -1610 0 1
rlabel polysilicon 163 -1616 163 -1616 0 3
rlabel polysilicon 170 -1610 170 -1610 0 1
rlabel polysilicon 170 -1616 170 -1616 0 3
rlabel polysilicon 177 -1610 177 -1610 0 1
rlabel polysilicon 177 -1616 177 -1616 0 3
rlabel polysilicon 184 -1610 184 -1610 0 1
rlabel polysilicon 184 -1616 184 -1616 0 3
rlabel polysilicon 191 -1610 191 -1610 0 1
rlabel polysilicon 194 -1610 194 -1610 0 2
rlabel polysilicon 191 -1616 191 -1616 0 3
rlabel polysilicon 194 -1616 194 -1616 0 4
rlabel polysilicon 198 -1610 198 -1610 0 1
rlabel polysilicon 198 -1616 198 -1616 0 3
rlabel polysilicon 205 -1610 205 -1610 0 1
rlabel polysilicon 208 -1610 208 -1610 0 2
rlabel polysilicon 205 -1616 205 -1616 0 3
rlabel polysilicon 208 -1616 208 -1616 0 4
rlabel polysilicon 212 -1610 212 -1610 0 1
rlabel polysilicon 212 -1616 212 -1616 0 3
rlabel polysilicon 219 -1610 219 -1610 0 1
rlabel polysilicon 219 -1616 219 -1616 0 3
rlabel polysilicon 226 -1610 226 -1610 0 1
rlabel polysilicon 226 -1616 226 -1616 0 3
rlabel polysilicon 233 -1610 233 -1610 0 1
rlabel polysilicon 233 -1616 233 -1616 0 3
rlabel polysilicon 240 -1610 240 -1610 0 1
rlabel polysilicon 240 -1616 240 -1616 0 3
rlabel polysilicon 247 -1610 247 -1610 0 1
rlabel polysilicon 247 -1616 247 -1616 0 3
rlabel polysilicon 257 -1610 257 -1610 0 2
rlabel polysilicon 254 -1616 254 -1616 0 3
rlabel polysilicon 261 -1610 261 -1610 0 1
rlabel polysilicon 261 -1616 261 -1616 0 3
rlabel polysilicon 268 -1616 268 -1616 0 3
rlabel polysilicon 271 -1616 271 -1616 0 4
rlabel polysilicon 275 -1610 275 -1610 0 1
rlabel polysilicon 275 -1616 275 -1616 0 3
rlabel polysilicon 282 -1610 282 -1610 0 1
rlabel polysilicon 282 -1616 282 -1616 0 3
rlabel polysilicon 289 -1610 289 -1610 0 1
rlabel polysilicon 292 -1610 292 -1610 0 2
rlabel polysilicon 289 -1616 289 -1616 0 3
rlabel polysilicon 296 -1610 296 -1610 0 1
rlabel polysilicon 296 -1616 296 -1616 0 3
rlabel polysilicon 303 -1610 303 -1610 0 1
rlabel polysilicon 303 -1616 303 -1616 0 3
rlabel polysilicon 310 -1610 310 -1610 0 1
rlabel polysilicon 310 -1616 310 -1616 0 3
rlabel polysilicon 320 -1616 320 -1616 0 4
rlabel polysilicon 324 -1610 324 -1610 0 1
rlabel polysilicon 324 -1616 324 -1616 0 3
rlabel polysilicon 331 -1610 331 -1610 0 1
rlabel polysilicon 331 -1616 331 -1616 0 3
rlabel polysilicon 338 -1610 338 -1610 0 1
rlabel polysilicon 338 -1616 338 -1616 0 3
rlabel polysilicon 345 -1610 345 -1610 0 1
rlabel polysilicon 345 -1616 345 -1616 0 3
rlabel polysilicon 352 -1610 352 -1610 0 1
rlabel polysilicon 352 -1616 352 -1616 0 3
rlabel polysilicon 359 -1610 359 -1610 0 1
rlabel polysilicon 359 -1616 359 -1616 0 3
rlabel polysilicon 366 -1610 366 -1610 0 1
rlabel polysilicon 369 -1610 369 -1610 0 2
rlabel polysilicon 366 -1616 366 -1616 0 3
rlabel polysilicon 369 -1616 369 -1616 0 4
rlabel polysilicon 373 -1610 373 -1610 0 1
rlabel polysilicon 373 -1616 373 -1616 0 3
rlabel polysilicon 380 -1610 380 -1610 0 1
rlabel polysilicon 383 -1610 383 -1610 0 2
rlabel polysilicon 380 -1616 380 -1616 0 3
rlabel polysilicon 383 -1616 383 -1616 0 4
rlabel polysilicon 387 -1610 387 -1610 0 1
rlabel polysilicon 387 -1616 387 -1616 0 3
rlabel polysilicon 394 -1610 394 -1610 0 1
rlabel polysilicon 394 -1616 394 -1616 0 3
rlabel polysilicon 401 -1610 401 -1610 0 1
rlabel polysilicon 401 -1616 401 -1616 0 3
rlabel polysilicon 408 -1610 408 -1610 0 1
rlabel polysilicon 408 -1616 408 -1616 0 3
rlabel polysilicon 415 -1610 415 -1610 0 1
rlabel polysilicon 415 -1616 415 -1616 0 3
rlabel polysilicon 422 -1610 422 -1610 0 1
rlabel polysilicon 422 -1616 422 -1616 0 3
rlabel polysilicon 429 -1610 429 -1610 0 1
rlabel polysilicon 429 -1616 429 -1616 0 3
rlabel polysilicon 436 -1610 436 -1610 0 1
rlabel polysilicon 436 -1616 436 -1616 0 3
rlabel polysilicon 443 -1610 443 -1610 0 1
rlabel polysilicon 443 -1616 443 -1616 0 3
rlabel polysilicon 450 -1610 450 -1610 0 1
rlabel polysilicon 450 -1616 450 -1616 0 3
rlabel polysilicon 457 -1610 457 -1610 0 1
rlabel polysilicon 457 -1616 457 -1616 0 3
rlabel polysilicon 464 -1610 464 -1610 0 1
rlabel polysilicon 464 -1616 464 -1616 0 3
rlabel polysilicon 471 -1610 471 -1610 0 1
rlabel polysilicon 474 -1610 474 -1610 0 2
rlabel polysilicon 471 -1616 471 -1616 0 3
rlabel polysilicon 478 -1610 478 -1610 0 1
rlabel polysilicon 478 -1616 478 -1616 0 3
rlabel polysilicon 485 -1610 485 -1610 0 1
rlabel polysilicon 485 -1616 485 -1616 0 3
rlabel polysilicon 492 -1610 492 -1610 0 1
rlabel polysilicon 492 -1616 492 -1616 0 3
rlabel polysilicon 495 -1616 495 -1616 0 4
rlabel polysilicon 499 -1610 499 -1610 0 1
rlabel polysilicon 499 -1616 499 -1616 0 3
rlabel polysilicon 506 -1610 506 -1610 0 1
rlabel polysilicon 506 -1616 506 -1616 0 3
rlabel polysilicon 513 -1610 513 -1610 0 1
rlabel polysilicon 513 -1616 513 -1616 0 3
rlabel polysilicon 520 -1610 520 -1610 0 1
rlabel polysilicon 520 -1616 520 -1616 0 3
rlabel polysilicon 527 -1610 527 -1610 0 1
rlabel polysilicon 527 -1616 527 -1616 0 3
rlabel polysilicon 530 -1616 530 -1616 0 4
rlabel polysilicon 534 -1610 534 -1610 0 1
rlabel polysilicon 534 -1616 534 -1616 0 3
rlabel polysilicon 541 -1610 541 -1610 0 1
rlabel polysilicon 544 -1610 544 -1610 0 2
rlabel polysilicon 541 -1616 541 -1616 0 3
rlabel polysilicon 544 -1616 544 -1616 0 4
rlabel polysilicon 548 -1610 548 -1610 0 1
rlabel polysilicon 548 -1616 548 -1616 0 3
rlabel polysilicon 555 -1610 555 -1610 0 1
rlabel polysilicon 555 -1616 555 -1616 0 3
rlabel polysilicon 562 -1610 562 -1610 0 1
rlabel polysilicon 562 -1616 562 -1616 0 3
rlabel polysilicon 565 -1616 565 -1616 0 4
rlabel polysilicon 569 -1610 569 -1610 0 1
rlabel polysilicon 569 -1616 569 -1616 0 3
rlabel polysilicon 576 -1610 576 -1610 0 1
rlabel polysilicon 576 -1616 576 -1616 0 3
rlabel polysilicon 583 -1610 583 -1610 0 1
rlabel polysilicon 583 -1616 583 -1616 0 3
rlabel polysilicon 590 -1610 590 -1610 0 1
rlabel polysilicon 590 -1616 590 -1616 0 3
rlabel polysilicon 597 -1610 597 -1610 0 1
rlabel polysilicon 597 -1616 597 -1616 0 3
rlabel polysilicon 604 -1610 604 -1610 0 1
rlabel polysilicon 607 -1610 607 -1610 0 2
rlabel polysilicon 604 -1616 604 -1616 0 3
rlabel polysilicon 607 -1616 607 -1616 0 4
rlabel polysilicon 611 -1610 611 -1610 0 1
rlabel polysilicon 614 -1610 614 -1610 0 2
rlabel polysilicon 611 -1616 611 -1616 0 3
rlabel polysilicon 614 -1616 614 -1616 0 4
rlabel polysilicon 618 -1610 618 -1610 0 1
rlabel polysilicon 621 -1610 621 -1610 0 2
rlabel polysilicon 618 -1616 618 -1616 0 3
rlabel polysilicon 621 -1616 621 -1616 0 4
rlabel polysilicon 625 -1610 625 -1610 0 1
rlabel polysilicon 632 -1610 632 -1610 0 1
rlabel polysilicon 632 -1616 632 -1616 0 3
rlabel polysilicon 639 -1610 639 -1610 0 1
rlabel polysilicon 639 -1616 639 -1616 0 3
rlabel polysilicon 646 -1610 646 -1610 0 1
rlabel polysilicon 646 -1616 646 -1616 0 3
rlabel polysilicon 653 -1610 653 -1610 0 1
rlabel polysilicon 653 -1616 653 -1616 0 3
rlabel polysilicon 660 -1610 660 -1610 0 1
rlabel polysilicon 660 -1616 660 -1616 0 3
rlabel polysilicon 667 -1610 667 -1610 0 1
rlabel polysilicon 670 -1610 670 -1610 0 2
rlabel polysilicon 667 -1616 667 -1616 0 3
rlabel polysilicon 670 -1616 670 -1616 0 4
rlabel polysilicon 674 -1610 674 -1610 0 1
rlabel polysilicon 674 -1616 674 -1616 0 3
rlabel polysilicon 681 -1610 681 -1610 0 1
rlabel polysilicon 681 -1616 681 -1616 0 3
rlabel polysilicon 688 -1610 688 -1610 0 1
rlabel polysilicon 688 -1616 688 -1616 0 3
rlabel polysilicon 695 -1610 695 -1610 0 1
rlabel polysilicon 695 -1616 695 -1616 0 3
rlabel polysilicon 702 -1610 702 -1610 0 1
rlabel polysilicon 702 -1616 702 -1616 0 3
rlabel polysilicon 709 -1610 709 -1610 0 1
rlabel polysilicon 712 -1610 712 -1610 0 2
rlabel polysilicon 709 -1616 709 -1616 0 3
rlabel polysilicon 712 -1616 712 -1616 0 4
rlabel polysilicon 716 -1610 716 -1610 0 1
rlabel polysilicon 719 -1610 719 -1610 0 2
rlabel polysilicon 716 -1616 716 -1616 0 3
rlabel polysilicon 719 -1616 719 -1616 0 4
rlabel polysilicon 723 -1610 723 -1610 0 1
rlabel polysilicon 726 -1610 726 -1610 0 2
rlabel polysilicon 723 -1616 723 -1616 0 3
rlabel polysilicon 726 -1616 726 -1616 0 4
rlabel polysilicon 730 -1610 730 -1610 0 1
rlabel polysilicon 730 -1616 730 -1616 0 3
rlabel polysilicon 737 -1610 737 -1610 0 1
rlabel polysilicon 740 -1610 740 -1610 0 2
rlabel polysilicon 737 -1616 737 -1616 0 3
rlabel polysilicon 740 -1616 740 -1616 0 4
rlabel polysilicon 744 -1610 744 -1610 0 1
rlabel polysilicon 747 -1610 747 -1610 0 2
rlabel polysilicon 747 -1616 747 -1616 0 4
rlabel polysilicon 751 -1610 751 -1610 0 1
rlabel polysilicon 751 -1616 751 -1616 0 3
rlabel polysilicon 758 -1610 758 -1610 0 1
rlabel polysilicon 761 -1610 761 -1610 0 2
rlabel polysilicon 758 -1616 758 -1616 0 3
rlabel polysilicon 761 -1616 761 -1616 0 4
rlabel polysilicon 765 -1610 765 -1610 0 1
rlabel polysilicon 765 -1616 765 -1616 0 3
rlabel polysilicon 772 -1610 772 -1610 0 1
rlabel polysilicon 772 -1616 772 -1616 0 3
rlabel polysilicon 779 -1610 779 -1610 0 1
rlabel polysilicon 779 -1616 779 -1616 0 3
rlabel polysilicon 786 -1610 786 -1610 0 1
rlabel polysilicon 786 -1616 786 -1616 0 3
rlabel polysilicon 793 -1610 793 -1610 0 1
rlabel polysilicon 796 -1610 796 -1610 0 2
rlabel polysilicon 793 -1616 793 -1616 0 3
rlabel polysilicon 796 -1616 796 -1616 0 4
rlabel polysilicon 800 -1610 800 -1610 0 1
rlabel polysilicon 800 -1616 800 -1616 0 3
rlabel polysilicon 807 -1610 807 -1610 0 1
rlabel polysilicon 807 -1616 807 -1616 0 3
rlabel polysilicon 814 -1610 814 -1610 0 1
rlabel polysilicon 814 -1616 814 -1616 0 3
rlabel polysilicon 821 -1610 821 -1610 0 1
rlabel polysilicon 821 -1616 821 -1616 0 3
rlabel polysilicon 828 -1610 828 -1610 0 1
rlabel polysilicon 828 -1616 828 -1616 0 3
rlabel polysilicon 835 -1610 835 -1610 0 1
rlabel polysilicon 835 -1616 835 -1616 0 3
rlabel polysilicon 842 -1610 842 -1610 0 1
rlabel polysilicon 842 -1616 842 -1616 0 3
rlabel polysilicon 849 -1610 849 -1610 0 1
rlabel polysilicon 849 -1616 849 -1616 0 3
rlabel polysilicon 856 -1610 856 -1610 0 1
rlabel polysilicon 856 -1616 856 -1616 0 3
rlabel polysilicon 863 -1610 863 -1610 0 1
rlabel polysilicon 863 -1616 863 -1616 0 3
rlabel polysilicon 870 -1610 870 -1610 0 1
rlabel polysilicon 870 -1616 870 -1616 0 3
rlabel polysilicon 877 -1610 877 -1610 0 1
rlabel polysilicon 877 -1616 877 -1616 0 3
rlabel polysilicon 884 -1610 884 -1610 0 1
rlabel polysilicon 884 -1616 884 -1616 0 3
rlabel polysilicon 891 -1610 891 -1610 0 1
rlabel polysilicon 891 -1616 891 -1616 0 3
rlabel polysilicon 898 -1610 898 -1610 0 1
rlabel polysilicon 898 -1616 898 -1616 0 3
rlabel polysilicon 905 -1610 905 -1610 0 1
rlabel polysilicon 905 -1616 905 -1616 0 3
rlabel polysilicon 912 -1610 912 -1610 0 1
rlabel polysilicon 912 -1616 912 -1616 0 3
rlabel polysilicon 919 -1610 919 -1610 0 1
rlabel polysilicon 919 -1616 919 -1616 0 3
rlabel polysilicon 926 -1610 926 -1610 0 1
rlabel polysilicon 929 -1610 929 -1610 0 2
rlabel polysilicon 926 -1616 926 -1616 0 3
rlabel polysilicon 929 -1616 929 -1616 0 4
rlabel polysilicon 933 -1610 933 -1610 0 1
rlabel polysilicon 933 -1616 933 -1616 0 3
rlabel polysilicon 940 -1610 940 -1610 0 1
rlabel polysilicon 940 -1616 940 -1616 0 3
rlabel polysilicon 947 -1610 947 -1610 0 1
rlabel polysilicon 947 -1616 947 -1616 0 3
rlabel polysilicon 954 -1610 954 -1610 0 1
rlabel polysilicon 954 -1616 954 -1616 0 3
rlabel polysilicon 961 -1610 961 -1610 0 1
rlabel polysilicon 961 -1616 961 -1616 0 3
rlabel polysilicon 968 -1610 968 -1610 0 1
rlabel polysilicon 968 -1616 968 -1616 0 3
rlabel polysilicon 975 -1610 975 -1610 0 1
rlabel polysilicon 975 -1616 975 -1616 0 3
rlabel polysilicon 982 -1610 982 -1610 0 1
rlabel polysilicon 982 -1616 982 -1616 0 3
rlabel polysilicon 989 -1610 989 -1610 0 1
rlabel polysilicon 989 -1616 989 -1616 0 3
rlabel polysilicon 996 -1610 996 -1610 0 1
rlabel polysilicon 996 -1616 996 -1616 0 3
rlabel polysilicon 1003 -1610 1003 -1610 0 1
rlabel polysilicon 1003 -1616 1003 -1616 0 3
rlabel polysilicon 1010 -1610 1010 -1610 0 1
rlabel polysilicon 1010 -1616 1010 -1616 0 3
rlabel polysilicon 1017 -1610 1017 -1610 0 1
rlabel polysilicon 1020 -1610 1020 -1610 0 2
rlabel polysilicon 1017 -1616 1017 -1616 0 3
rlabel polysilicon 1020 -1616 1020 -1616 0 4
rlabel polysilicon 1024 -1610 1024 -1610 0 1
rlabel polysilicon 1024 -1616 1024 -1616 0 3
rlabel polysilicon 1031 -1610 1031 -1610 0 1
rlabel polysilicon 1031 -1616 1031 -1616 0 3
rlabel polysilicon 1038 -1610 1038 -1610 0 1
rlabel polysilicon 1038 -1616 1038 -1616 0 3
rlabel polysilicon 1045 -1610 1045 -1610 0 1
rlabel polysilicon 1048 -1610 1048 -1610 0 2
rlabel polysilicon 1045 -1616 1045 -1616 0 3
rlabel polysilicon 1048 -1616 1048 -1616 0 4
rlabel polysilicon 1052 -1610 1052 -1610 0 1
rlabel polysilicon 1052 -1616 1052 -1616 0 3
rlabel polysilicon 1062 -1610 1062 -1610 0 2
rlabel polysilicon 1059 -1616 1059 -1616 0 3
rlabel polysilicon 1066 -1610 1066 -1610 0 1
rlabel polysilicon 1066 -1616 1066 -1616 0 3
rlabel polysilicon 1073 -1610 1073 -1610 0 1
rlabel polysilicon 1073 -1616 1073 -1616 0 3
rlabel polysilicon 1080 -1610 1080 -1610 0 1
rlabel polysilicon 1080 -1616 1080 -1616 0 3
rlabel polysilicon 1087 -1610 1087 -1610 0 1
rlabel polysilicon 1087 -1616 1087 -1616 0 3
rlabel polysilicon 1094 -1610 1094 -1610 0 1
rlabel polysilicon 1094 -1616 1094 -1616 0 3
rlabel polysilicon 1101 -1610 1101 -1610 0 1
rlabel polysilicon 1104 -1610 1104 -1610 0 2
rlabel polysilicon 1101 -1616 1101 -1616 0 3
rlabel polysilicon 1104 -1616 1104 -1616 0 4
rlabel polysilicon 1108 -1610 1108 -1610 0 1
rlabel polysilicon 1108 -1616 1108 -1616 0 3
rlabel polysilicon 1115 -1610 1115 -1610 0 1
rlabel polysilicon 1118 -1610 1118 -1610 0 2
rlabel polysilicon 1115 -1616 1115 -1616 0 3
rlabel polysilicon 1118 -1616 1118 -1616 0 4
rlabel polysilicon 1122 -1610 1122 -1610 0 1
rlabel polysilicon 1122 -1616 1122 -1616 0 3
rlabel polysilicon 1129 -1610 1129 -1610 0 1
rlabel polysilicon 1129 -1616 1129 -1616 0 3
rlabel polysilicon 1136 -1610 1136 -1610 0 1
rlabel polysilicon 1136 -1616 1136 -1616 0 3
rlabel polysilicon 1143 -1610 1143 -1610 0 1
rlabel polysilicon 1143 -1616 1143 -1616 0 3
rlabel polysilicon 1153 -1610 1153 -1610 0 2
rlabel polysilicon 1150 -1616 1150 -1616 0 3
rlabel polysilicon 1153 -1616 1153 -1616 0 4
rlabel polysilicon 1157 -1610 1157 -1610 0 1
rlabel polysilicon 1157 -1616 1157 -1616 0 3
rlabel polysilicon 1164 -1610 1164 -1610 0 1
rlabel polysilicon 1164 -1616 1164 -1616 0 3
rlabel polysilicon 1171 -1610 1171 -1610 0 1
rlabel polysilicon 1171 -1616 1171 -1616 0 3
rlabel polysilicon 1178 -1610 1178 -1610 0 1
rlabel polysilicon 1178 -1616 1178 -1616 0 3
rlabel polysilicon 1185 -1610 1185 -1610 0 1
rlabel polysilicon 1185 -1616 1185 -1616 0 3
rlabel polysilicon 1192 -1610 1192 -1610 0 1
rlabel polysilicon 1192 -1616 1192 -1616 0 3
rlabel polysilicon 1199 -1610 1199 -1610 0 1
rlabel polysilicon 1199 -1616 1199 -1616 0 3
rlabel polysilicon 1206 -1610 1206 -1610 0 1
rlabel polysilicon 1206 -1616 1206 -1616 0 3
rlabel polysilicon 1213 -1610 1213 -1610 0 1
rlabel polysilicon 1213 -1616 1213 -1616 0 3
rlabel polysilicon 1220 -1610 1220 -1610 0 1
rlabel polysilicon 1220 -1616 1220 -1616 0 3
rlabel polysilicon 1227 -1610 1227 -1610 0 1
rlabel polysilicon 1227 -1616 1227 -1616 0 3
rlabel polysilicon 1234 -1610 1234 -1610 0 1
rlabel polysilicon 1234 -1616 1234 -1616 0 3
rlabel polysilicon 1241 -1610 1241 -1610 0 1
rlabel polysilicon 1241 -1616 1241 -1616 0 3
rlabel polysilicon 1248 -1610 1248 -1610 0 1
rlabel polysilicon 1248 -1616 1248 -1616 0 3
rlabel polysilicon 1255 -1610 1255 -1610 0 1
rlabel polysilicon 1258 -1610 1258 -1610 0 2
rlabel polysilicon 1255 -1616 1255 -1616 0 3
rlabel polysilicon 1262 -1610 1262 -1610 0 1
rlabel polysilicon 1262 -1616 1262 -1616 0 3
rlabel polysilicon 1269 -1610 1269 -1610 0 1
rlabel polysilicon 1269 -1616 1269 -1616 0 3
rlabel polysilicon 1276 -1610 1276 -1610 0 1
rlabel polysilicon 1276 -1616 1276 -1616 0 3
rlabel polysilicon 1283 -1610 1283 -1610 0 1
rlabel polysilicon 1283 -1616 1283 -1616 0 3
rlabel polysilicon 1290 -1610 1290 -1610 0 1
rlabel polysilicon 1290 -1616 1290 -1616 0 3
rlabel polysilicon 1297 -1610 1297 -1610 0 1
rlabel polysilicon 1297 -1616 1297 -1616 0 3
rlabel polysilicon 1304 -1610 1304 -1610 0 1
rlabel polysilicon 1304 -1616 1304 -1616 0 3
rlabel polysilicon 1311 -1610 1311 -1610 0 1
rlabel polysilicon 1311 -1616 1311 -1616 0 3
rlabel polysilicon 1318 -1610 1318 -1610 0 1
rlabel polysilicon 1318 -1616 1318 -1616 0 3
rlabel polysilicon 1325 -1610 1325 -1610 0 1
rlabel polysilicon 1325 -1616 1325 -1616 0 3
rlabel polysilicon 1332 -1610 1332 -1610 0 1
rlabel polysilicon 1332 -1616 1332 -1616 0 3
rlabel polysilicon 1339 -1610 1339 -1610 0 1
rlabel polysilicon 1339 -1616 1339 -1616 0 3
rlabel polysilicon 1346 -1610 1346 -1610 0 1
rlabel polysilicon 1346 -1616 1346 -1616 0 3
rlabel polysilicon 1353 -1610 1353 -1610 0 1
rlabel polysilicon 1353 -1616 1353 -1616 0 3
rlabel polysilicon 1360 -1610 1360 -1610 0 1
rlabel polysilicon 1360 -1616 1360 -1616 0 3
rlabel polysilicon 1367 -1610 1367 -1610 0 1
rlabel polysilicon 1367 -1616 1367 -1616 0 3
rlabel polysilicon 1374 -1610 1374 -1610 0 1
rlabel polysilicon 1374 -1616 1374 -1616 0 3
rlabel polysilicon 1381 -1610 1381 -1610 0 1
rlabel polysilicon 1381 -1616 1381 -1616 0 3
rlabel polysilicon 1384 -1616 1384 -1616 0 4
rlabel polysilicon 1388 -1610 1388 -1610 0 1
rlabel polysilicon 1388 -1616 1388 -1616 0 3
rlabel polysilicon 1395 -1610 1395 -1610 0 1
rlabel polysilicon 1395 -1616 1395 -1616 0 3
rlabel polysilicon 1402 -1610 1402 -1610 0 1
rlabel polysilicon 1402 -1616 1402 -1616 0 3
rlabel polysilicon 1409 -1610 1409 -1610 0 1
rlabel polysilicon 1409 -1616 1409 -1616 0 3
rlabel polysilicon 1416 -1610 1416 -1610 0 1
rlabel polysilicon 1416 -1616 1416 -1616 0 3
rlabel polysilicon 1423 -1610 1423 -1610 0 1
rlabel polysilicon 1423 -1616 1423 -1616 0 3
rlabel polysilicon 1430 -1610 1430 -1610 0 1
rlabel polysilicon 1430 -1616 1430 -1616 0 3
rlabel polysilicon 1437 -1610 1437 -1610 0 1
rlabel polysilicon 1437 -1616 1437 -1616 0 3
rlabel polysilicon 1444 -1610 1444 -1610 0 1
rlabel polysilicon 1444 -1616 1444 -1616 0 3
rlabel polysilicon 1451 -1610 1451 -1610 0 1
rlabel polysilicon 1451 -1616 1451 -1616 0 3
rlabel polysilicon 1458 -1610 1458 -1610 0 1
rlabel polysilicon 1458 -1616 1458 -1616 0 3
rlabel polysilicon 1465 -1610 1465 -1610 0 1
rlabel polysilicon 1465 -1616 1465 -1616 0 3
rlabel polysilicon 1472 -1610 1472 -1610 0 1
rlabel polysilicon 1472 -1616 1472 -1616 0 3
rlabel polysilicon 1479 -1610 1479 -1610 0 1
rlabel polysilicon 1479 -1616 1479 -1616 0 3
rlabel polysilicon 1486 -1610 1486 -1610 0 1
rlabel polysilicon 1486 -1616 1486 -1616 0 3
rlabel polysilicon 1493 -1610 1493 -1610 0 1
rlabel polysilicon 1493 -1616 1493 -1616 0 3
rlabel polysilicon 1500 -1610 1500 -1610 0 1
rlabel polysilicon 1500 -1616 1500 -1616 0 3
rlabel polysilicon 1507 -1610 1507 -1610 0 1
rlabel polysilicon 1507 -1616 1507 -1616 0 3
rlabel polysilicon 1514 -1610 1514 -1610 0 1
rlabel polysilicon 1514 -1616 1514 -1616 0 3
rlabel polysilicon 1521 -1610 1521 -1610 0 1
rlabel polysilicon 1521 -1616 1521 -1616 0 3
rlabel polysilicon 1528 -1610 1528 -1610 0 1
rlabel polysilicon 1528 -1616 1528 -1616 0 3
rlabel polysilicon 1535 -1610 1535 -1610 0 1
rlabel polysilicon 1535 -1616 1535 -1616 0 3
rlabel polysilicon 1542 -1610 1542 -1610 0 1
rlabel polysilicon 1542 -1616 1542 -1616 0 3
rlabel polysilicon 1549 -1610 1549 -1610 0 1
rlabel polysilicon 1549 -1616 1549 -1616 0 3
rlabel polysilicon 1556 -1610 1556 -1610 0 1
rlabel polysilicon 1556 -1616 1556 -1616 0 3
rlabel polysilicon 1563 -1610 1563 -1610 0 1
rlabel polysilicon 1563 -1616 1563 -1616 0 3
rlabel polysilicon 1570 -1610 1570 -1610 0 1
rlabel polysilicon 1570 -1616 1570 -1616 0 3
rlabel polysilicon 1577 -1610 1577 -1610 0 1
rlabel polysilicon 1577 -1616 1577 -1616 0 3
rlabel polysilicon 1584 -1610 1584 -1610 0 1
rlabel polysilicon 1584 -1616 1584 -1616 0 3
rlabel polysilicon 1591 -1610 1591 -1610 0 1
rlabel polysilicon 1591 -1616 1591 -1616 0 3
rlabel polysilicon 1598 -1610 1598 -1610 0 1
rlabel polysilicon 1598 -1616 1598 -1616 0 3
rlabel polysilicon 1605 -1610 1605 -1610 0 1
rlabel polysilicon 1605 -1616 1605 -1616 0 3
rlabel polysilicon 1612 -1610 1612 -1610 0 1
rlabel polysilicon 1612 -1616 1612 -1616 0 3
rlabel polysilicon 1619 -1610 1619 -1610 0 1
rlabel polysilicon 1619 -1616 1619 -1616 0 3
rlabel polysilicon 1626 -1610 1626 -1610 0 1
rlabel polysilicon 1626 -1616 1626 -1616 0 3
rlabel polysilicon 1633 -1610 1633 -1610 0 1
rlabel polysilicon 1633 -1616 1633 -1616 0 3
rlabel polysilicon 1640 -1610 1640 -1610 0 1
rlabel polysilicon 1640 -1616 1640 -1616 0 3
rlabel polysilicon 1647 -1610 1647 -1610 0 1
rlabel polysilicon 1647 -1616 1647 -1616 0 3
rlabel polysilicon 1654 -1610 1654 -1610 0 1
rlabel polysilicon 1654 -1616 1654 -1616 0 3
rlabel polysilicon 1661 -1610 1661 -1610 0 1
rlabel polysilicon 1661 -1616 1661 -1616 0 3
rlabel polysilicon 1668 -1610 1668 -1610 0 1
rlabel polysilicon 1668 -1616 1668 -1616 0 3
rlabel polysilicon 1675 -1610 1675 -1610 0 1
rlabel polysilicon 1675 -1616 1675 -1616 0 3
rlabel polysilicon 1682 -1610 1682 -1610 0 1
rlabel polysilicon 1682 -1616 1682 -1616 0 3
rlabel polysilicon 1689 -1610 1689 -1610 0 1
rlabel polysilicon 1689 -1616 1689 -1616 0 3
rlabel polysilicon 1696 -1610 1696 -1610 0 1
rlabel polysilicon 1696 -1616 1696 -1616 0 3
rlabel polysilicon 1703 -1610 1703 -1610 0 1
rlabel polysilicon 1706 -1610 1706 -1610 0 2
rlabel polysilicon 1703 -1616 1703 -1616 0 3
rlabel polysilicon 1706 -1616 1706 -1616 0 4
rlabel polysilicon 1710 -1610 1710 -1610 0 1
rlabel polysilicon 1713 -1610 1713 -1610 0 2
rlabel polysilicon 1710 -1616 1710 -1616 0 3
rlabel polysilicon 1717 -1610 1717 -1610 0 1
rlabel polysilicon 1717 -1616 1717 -1616 0 3
rlabel polysilicon 1752 -1610 1752 -1610 0 1
rlabel polysilicon 1752 -1616 1752 -1616 0 3
rlabel polysilicon 16 -1737 16 -1737 0 1
rlabel polysilicon 37 -1737 37 -1737 0 1
rlabel polysilicon 37 -1743 37 -1743 0 3
rlabel polysilicon 44 -1737 44 -1737 0 1
rlabel polysilicon 44 -1743 44 -1743 0 3
rlabel polysilicon 51 -1737 51 -1737 0 1
rlabel polysilicon 51 -1743 51 -1743 0 3
rlabel polysilicon 58 -1737 58 -1737 0 1
rlabel polysilicon 61 -1737 61 -1737 0 2
rlabel polysilicon 61 -1743 61 -1743 0 4
rlabel polysilicon 65 -1737 65 -1737 0 1
rlabel polysilicon 65 -1743 65 -1743 0 3
rlabel polysilicon 72 -1737 72 -1737 0 1
rlabel polysilicon 72 -1743 72 -1743 0 3
rlabel polysilicon 79 -1737 79 -1737 0 1
rlabel polysilicon 79 -1743 79 -1743 0 3
rlabel polysilicon 86 -1737 86 -1737 0 1
rlabel polysilicon 86 -1743 86 -1743 0 3
rlabel polysilicon 93 -1737 93 -1737 0 1
rlabel polysilicon 93 -1743 93 -1743 0 3
rlabel polysilicon 100 -1737 100 -1737 0 1
rlabel polysilicon 100 -1743 100 -1743 0 3
rlabel polysilicon 107 -1737 107 -1737 0 1
rlabel polysilicon 107 -1743 107 -1743 0 3
rlabel polysilicon 114 -1737 114 -1737 0 1
rlabel polysilicon 114 -1743 114 -1743 0 3
rlabel polysilicon 121 -1737 121 -1737 0 1
rlabel polysilicon 121 -1743 121 -1743 0 3
rlabel polysilicon 128 -1737 128 -1737 0 1
rlabel polysilicon 128 -1743 128 -1743 0 3
rlabel polysilicon 135 -1737 135 -1737 0 1
rlabel polysilicon 135 -1743 135 -1743 0 3
rlabel polysilicon 142 -1737 142 -1737 0 1
rlabel polysilicon 142 -1743 142 -1743 0 3
rlabel polysilicon 149 -1737 149 -1737 0 1
rlabel polysilicon 149 -1743 149 -1743 0 3
rlabel polysilicon 156 -1737 156 -1737 0 1
rlabel polysilicon 159 -1737 159 -1737 0 2
rlabel polysilicon 156 -1743 156 -1743 0 3
rlabel polysilicon 159 -1743 159 -1743 0 4
rlabel polysilicon 163 -1737 163 -1737 0 1
rlabel polysilicon 163 -1743 163 -1743 0 3
rlabel polysilicon 170 -1737 170 -1737 0 1
rlabel polysilicon 173 -1737 173 -1737 0 2
rlabel polysilicon 170 -1743 170 -1743 0 3
rlabel polysilicon 177 -1737 177 -1737 0 1
rlabel polysilicon 177 -1743 177 -1743 0 3
rlabel polysilicon 180 -1743 180 -1743 0 4
rlabel polysilicon 184 -1737 184 -1737 0 1
rlabel polysilicon 184 -1743 184 -1743 0 3
rlabel polysilicon 191 -1737 191 -1737 0 1
rlabel polysilicon 191 -1743 191 -1743 0 3
rlabel polysilicon 194 -1743 194 -1743 0 4
rlabel polysilicon 198 -1737 198 -1737 0 1
rlabel polysilicon 198 -1743 198 -1743 0 3
rlabel polysilicon 205 -1737 205 -1737 0 1
rlabel polysilicon 205 -1743 205 -1743 0 3
rlabel polysilicon 212 -1737 212 -1737 0 1
rlabel polysilicon 212 -1743 212 -1743 0 3
rlabel polysilicon 219 -1737 219 -1737 0 1
rlabel polysilicon 219 -1743 219 -1743 0 3
rlabel polysilicon 226 -1737 226 -1737 0 1
rlabel polysilicon 226 -1743 226 -1743 0 3
rlabel polysilicon 233 -1737 233 -1737 0 1
rlabel polysilicon 233 -1743 233 -1743 0 3
rlabel polysilicon 240 -1737 240 -1737 0 1
rlabel polysilicon 240 -1743 240 -1743 0 3
rlabel polysilicon 247 -1737 247 -1737 0 1
rlabel polysilicon 247 -1743 247 -1743 0 3
rlabel polysilicon 257 -1737 257 -1737 0 2
rlabel polysilicon 254 -1743 254 -1743 0 3
rlabel polysilicon 257 -1743 257 -1743 0 4
rlabel polysilicon 264 -1737 264 -1737 0 2
rlabel polysilicon 264 -1743 264 -1743 0 4
rlabel polysilicon 268 -1737 268 -1737 0 1
rlabel polysilicon 268 -1743 268 -1743 0 3
rlabel polysilicon 275 -1737 275 -1737 0 1
rlabel polysilicon 278 -1737 278 -1737 0 2
rlabel polysilicon 275 -1743 275 -1743 0 3
rlabel polysilicon 282 -1737 282 -1737 0 1
rlabel polysilicon 282 -1743 282 -1743 0 3
rlabel polysilicon 289 -1737 289 -1737 0 1
rlabel polysilicon 289 -1743 289 -1743 0 3
rlabel polysilicon 296 -1737 296 -1737 0 1
rlabel polysilicon 296 -1743 296 -1743 0 3
rlabel polysilicon 303 -1737 303 -1737 0 1
rlabel polysilicon 303 -1743 303 -1743 0 3
rlabel polysilicon 310 -1737 310 -1737 0 1
rlabel polysilicon 310 -1743 310 -1743 0 3
rlabel polysilicon 317 -1737 317 -1737 0 1
rlabel polysilicon 317 -1743 317 -1743 0 3
rlabel polysilicon 324 -1737 324 -1737 0 1
rlabel polysilicon 324 -1743 324 -1743 0 3
rlabel polysilicon 331 -1737 331 -1737 0 1
rlabel polysilicon 331 -1743 331 -1743 0 3
rlabel polysilicon 338 -1737 338 -1737 0 1
rlabel polysilicon 338 -1743 338 -1743 0 3
rlabel polysilicon 345 -1737 345 -1737 0 1
rlabel polysilicon 348 -1737 348 -1737 0 2
rlabel polysilicon 348 -1743 348 -1743 0 4
rlabel polysilicon 352 -1737 352 -1737 0 1
rlabel polysilicon 352 -1743 352 -1743 0 3
rlabel polysilicon 359 -1737 359 -1737 0 1
rlabel polysilicon 359 -1743 359 -1743 0 3
rlabel polysilicon 366 -1737 366 -1737 0 1
rlabel polysilicon 366 -1743 366 -1743 0 3
rlabel polysilicon 373 -1737 373 -1737 0 1
rlabel polysilicon 373 -1743 373 -1743 0 3
rlabel polysilicon 380 -1737 380 -1737 0 1
rlabel polysilicon 380 -1743 380 -1743 0 3
rlabel polysilicon 387 -1737 387 -1737 0 1
rlabel polysilicon 387 -1743 387 -1743 0 3
rlabel polysilicon 394 -1737 394 -1737 0 1
rlabel polysilicon 394 -1743 394 -1743 0 3
rlabel polysilicon 401 -1737 401 -1737 0 1
rlabel polysilicon 401 -1743 401 -1743 0 3
rlabel polysilicon 411 -1737 411 -1737 0 2
rlabel polysilicon 411 -1743 411 -1743 0 4
rlabel polysilicon 415 -1737 415 -1737 0 1
rlabel polysilicon 415 -1743 415 -1743 0 3
rlabel polysilicon 422 -1737 422 -1737 0 1
rlabel polysilicon 422 -1743 422 -1743 0 3
rlabel polysilicon 429 -1737 429 -1737 0 1
rlabel polysilicon 432 -1737 432 -1737 0 2
rlabel polysilicon 432 -1743 432 -1743 0 4
rlabel polysilicon 436 -1737 436 -1737 0 1
rlabel polysilicon 436 -1743 436 -1743 0 3
rlabel polysilicon 443 -1737 443 -1737 0 1
rlabel polysilicon 443 -1743 443 -1743 0 3
rlabel polysilicon 450 -1737 450 -1737 0 1
rlabel polysilicon 450 -1743 450 -1743 0 3
rlabel polysilicon 457 -1737 457 -1737 0 1
rlabel polysilicon 457 -1743 457 -1743 0 3
rlabel polysilicon 464 -1737 464 -1737 0 1
rlabel polysilicon 464 -1743 464 -1743 0 3
rlabel polysilicon 471 -1737 471 -1737 0 1
rlabel polysilicon 471 -1743 471 -1743 0 3
rlabel polysilicon 478 -1737 478 -1737 0 1
rlabel polysilicon 481 -1737 481 -1737 0 2
rlabel polysilicon 478 -1743 478 -1743 0 3
rlabel polysilicon 481 -1743 481 -1743 0 4
rlabel polysilicon 485 -1737 485 -1737 0 1
rlabel polysilicon 485 -1743 485 -1743 0 3
rlabel polysilicon 492 -1737 492 -1737 0 1
rlabel polysilicon 492 -1743 492 -1743 0 3
rlabel polysilicon 499 -1737 499 -1737 0 1
rlabel polysilicon 499 -1743 499 -1743 0 3
rlabel polysilicon 506 -1737 506 -1737 0 1
rlabel polysilicon 506 -1743 506 -1743 0 3
rlabel polysilicon 513 -1737 513 -1737 0 1
rlabel polysilicon 513 -1743 513 -1743 0 3
rlabel polysilicon 520 -1737 520 -1737 0 1
rlabel polysilicon 520 -1743 520 -1743 0 3
rlabel polysilicon 527 -1737 527 -1737 0 1
rlabel polysilicon 530 -1737 530 -1737 0 2
rlabel polysilicon 527 -1743 527 -1743 0 3
rlabel polysilicon 530 -1743 530 -1743 0 4
rlabel polysilicon 534 -1737 534 -1737 0 1
rlabel polysilicon 534 -1743 534 -1743 0 3
rlabel polysilicon 541 -1737 541 -1737 0 1
rlabel polysilicon 544 -1737 544 -1737 0 2
rlabel polysilicon 541 -1743 541 -1743 0 3
rlabel polysilicon 548 -1737 548 -1737 0 1
rlabel polysilicon 548 -1743 548 -1743 0 3
rlabel polysilicon 555 -1737 555 -1737 0 1
rlabel polysilicon 555 -1743 555 -1743 0 3
rlabel polysilicon 562 -1737 562 -1737 0 1
rlabel polysilicon 562 -1743 562 -1743 0 3
rlabel polysilicon 569 -1737 569 -1737 0 1
rlabel polysilicon 569 -1743 569 -1743 0 3
rlabel polysilicon 576 -1737 576 -1737 0 1
rlabel polysilicon 576 -1743 576 -1743 0 3
rlabel polysilicon 583 -1737 583 -1737 0 1
rlabel polysilicon 583 -1743 583 -1743 0 3
rlabel polysilicon 590 -1737 590 -1737 0 1
rlabel polysilicon 590 -1743 590 -1743 0 3
rlabel polysilicon 597 -1737 597 -1737 0 1
rlabel polysilicon 597 -1743 597 -1743 0 3
rlabel polysilicon 604 -1737 604 -1737 0 1
rlabel polysilicon 604 -1743 604 -1743 0 3
rlabel polysilicon 611 -1737 611 -1737 0 1
rlabel polysilicon 611 -1743 611 -1743 0 3
rlabel polysilicon 618 -1737 618 -1737 0 1
rlabel polysilicon 618 -1743 618 -1743 0 3
rlabel polysilicon 625 -1743 625 -1743 0 3
rlabel polysilicon 632 -1737 632 -1737 0 1
rlabel polysilicon 632 -1743 632 -1743 0 3
rlabel polysilicon 639 -1737 639 -1737 0 1
rlabel polysilicon 639 -1743 639 -1743 0 3
rlabel polysilicon 646 -1737 646 -1737 0 1
rlabel polysilicon 646 -1743 646 -1743 0 3
rlabel polysilicon 653 -1737 653 -1737 0 1
rlabel polysilicon 653 -1743 653 -1743 0 3
rlabel polysilicon 660 -1737 660 -1737 0 1
rlabel polysilicon 660 -1743 660 -1743 0 3
rlabel polysilicon 667 -1737 667 -1737 0 1
rlabel polysilicon 667 -1743 667 -1743 0 3
rlabel polysilicon 677 -1737 677 -1737 0 2
rlabel polysilicon 674 -1743 674 -1743 0 3
rlabel polysilicon 677 -1743 677 -1743 0 4
rlabel polysilicon 681 -1737 681 -1737 0 1
rlabel polysilicon 681 -1743 681 -1743 0 3
rlabel polysilicon 688 -1737 688 -1737 0 1
rlabel polysilicon 688 -1743 688 -1743 0 3
rlabel polysilicon 691 -1743 691 -1743 0 4
rlabel polysilicon 695 -1737 695 -1737 0 1
rlabel polysilicon 695 -1743 695 -1743 0 3
rlabel polysilicon 702 -1743 702 -1743 0 3
rlabel polysilicon 709 -1737 709 -1737 0 1
rlabel polysilicon 709 -1743 709 -1743 0 3
rlabel polysilicon 716 -1737 716 -1737 0 1
rlabel polysilicon 716 -1743 716 -1743 0 3
rlabel polysilicon 723 -1737 723 -1737 0 1
rlabel polysilicon 726 -1737 726 -1737 0 2
rlabel polysilicon 723 -1743 723 -1743 0 3
rlabel polysilicon 726 -1743 726 -1743 0 4
rlabel polysilicon 730 -1737 730 -1737 0 1
rlabel polysilicon 733 -1737 733 -1737 0 2
rlabel polysilicon 733 -1743 733 -1743 0 4
rlabel polysilicon 740 -1737 740 -1737 0 2
rlabel polysilicon 737 -1743 737 -1743 0 3
rlabel polysilicon 740 -1743 740 -1743 0 4
rlabel polysilicon 744 -1737 744 -1737 0 1
rlabel polysilicon 744 -1743 744 -1743 0 3
rlabel polysilicon 751 -1737 751 -1737 0 1
rlabel polysilicon 751 -1743 751 -1743 0 3
rlabel polysilicon 758 -1737 758 -1737 0 1
rlabel polysilicon 758 -1743 758 -1743 0 3
rlabel polysilicon 765 -1737 765 -1737 0 1
rlabel polysilicon 765 -1743 765 -1743 0 3
rlabel polysilicon 772 -1737 772 -1737 0 1
rlabel polysilicon 772 -1743 772 -1743 0 3
rlabel polysilicon 779 -1737 779 -1737 0 1
rlabel polysilicon 782 -1737 782 -1737 0 2
rlabel polysilicon 779 -1743 779 -1743 0 3
rlabel polysilicon 782 -1743 782 -1743 0 4
rlabel polysilicon 789 -1737 789 -1737 0 2
rlabel polysilicon 789 -1743 789 -1743 0 4
rlabel polysilicon 793 -1737 793 -1737 0 1
rlabel polysilicon 793 -1743 793 -1743 0 3
rlabel polysilicon 800 -1737 800 -1737 0 1
rlabel polysilicon 803 -1737 803 -1737 0 2
rlabel polysilicon 800 -1743 800 -1743 0 3
rlabel polysilicon 803 -1743 803 -1743 0 4
rlabel polysilicon 807 -1737 807 -1737 0 1
rlabel polysilicon 807 -1743 807 -1743 0 3
rlabel polysilicon 810 -1743 810 -1743 0 4
rlabel polysilicon 814 -1737 814 -1737 0 1
rlabel polysilicon 814 -1743 814 -1743 0 3
rlabel polysilicon 821 -1737 821 -1737 0 1
rlabel polysilicon 821 -1743 821 -1743 0 3
rlabel polysilicon 828 -1737 828 -1737 0 1
rlabel polysilicon 828 -1743 828 -1743 0 3
rlabel polysilicon 831 -1743 831 -1743 0 4
rlabel polysilicon 835 -1737 835 -1737 0 1
rlabel polysilicon 835 -1743 835 -1743 0 3
rlabel polysilicon 842 -1737 842 -1737 0 1
rlabel polysilicon 842 -1743 842 -1743 0 3
rlabel polysilicon 849 -1737 849 -1737 0 1
rlabel polysilicon 849 -1743 849 -1743 0 3
rlabel polysilicon 856 -1737 856 -1737 0 1
rlabel polysilicon 856 -1743 856 -1743 0 3
rlabel polysilicon 863 -1737 863 -1737 0 1
rlabel polysilicon 863 -1743 863 -1743 0 3
rlabel polysilicon 870 -1737 870 -1737 0 1
rlabel polysilicon 873 -1737 873 -1737 0 2
rlabel polysilicon 870 -1743 870 -1743 0 3
rlabel polysilicon 877 -1737 877 -1737 0 1
rlabel polysilicon 877 -1743 877 -1743 0 3
rlabel polysilicon 884 -1737 884 -1737 0 1
rlabel polysilicon 887 -1737 887 -1737 0 2
rlabel polysilicon 887 -1743 887 -1743 0 4
rlabel polysilicon 894 -1737 894 -1737 0 2
rlabel polysilicon 891 -1743 891 -1743 0 3
rlabel polysilicon 894 -1743 894 -1743 0 4
rlabel polysilicon 898 -1737 898 -1737 0 1
rlabel polysilicon 898 -1743 898 -1743 0 3
rlabel polysilicon 905 -1737 905 -1737 0 1
rlabel polysilicon 905 -1743 905 -1743 0 3
rlabel polysilicon 915 -1737 915 -1737 0 2
rlabel polysilicon 912 -1743 912 -1743 0 3
rlabel polysilicon 915 -1743 915 -1743 0 4
rlabel polysilicon 919 -1737 919 -1737 0 1
rlabel polysilicon 922 -1737 922 -1737 0 2
rlabel polysilicon 919 -1743 919 -1743 0 3
rlabel polysilicon 922 -1743 922 -1743 0 4
rlabel polysilicon 926 -1737 926 -1737 0 1
rlabel polysilicon 929 -1737 929 -1737 0 2
rlabel polysilicon 926 -1743 926 -1743 0 3
rlabel polysilicon 929 -1743 929 -1743 0 4
rlabel polysilicon 933 -1737 933 -1737 0 1
rlabel polysilicon 933 -1743 933 -1743 0 3
rlabel polysilicon 940 -1737 940 -1737 0 1
rlabel polysilicon 940 -1743 940 -1743 0 3
rlabel polysilicon 947 -1737 947 -1737 0 1
rlabel polysilicon 947 -1743 947 -1743 0 3
rlabel polysilicon 954 -1737 954 -1737 0 1
rlabel polysilicon 954 -1743 954 -1743 0 3
rlabel polysilicon 961 -1737 961 -1737 0 1
rlabel polysilicon 961 -1743 961 -1743 0 3
rlabel polysilicon 968 -1737 968 -1737 0 1
rlabel polysilicon 968 -1743 968 -1743 0 3
rlabel polysilicon 975 -1737 975 -1737 0 1
rlabel polysilicon 978 -1737 978 -1737 0 2
rlabel polysilicon 978 -1743 978 -1743 0 4
rlabel polysilicon 982 -1737 982 -1737 0 1
rlabel polysilicon 982 -1743 982 -1743 0 3
rlabel polysilicon 989 -1737 989 -1737 0 1
rlabel polysilicon 992 -1737 992 -1737 0 2
rlabel polysilicon 989 -1743 989 -1743 0 3
rlabel polysilicon 996 -1737 996 -1737 0 1
rlabel polysilicon 996 -1743 996 -1743 0 3
rlabel polysilicon 1003 -1737 1003 -1737 0 1
rlabel polysilicon 1003 -1743 1003 -1743 0 3
rlabel polysilicon 1010 -1737 1010 -1737 0 1
rlabel polysilicon 1010 -1743 1010 -1743 0 3
rlabel polysilicon 1017 -1737 1017 -1737 0 1
rlabel polysilicon 1017 -1743 1017 -1743 0 3
rlabel polysilicon 1024 -1737 1024 -1737 0 1
rlabel polysilicon 1024 -1743 1024 -1743 0 3
rlabel polysilicon 1031 -1737 1031 -1737 0 1
rlabel polysilicon 1031 -1743 1031 -1743 0 3
rlabel polysilicon 1038 -1737 1038 -1737 0 1
rlabel polysilicon 1038 -1743 1038 -1743 0 3
rlabel polysilicon 1045 -1737 1045 -1737 0 1
rlabel polysilicon 1045 -1743 1045 -1743 0 3
rlabel polysilicon 1052 -1737 1052 -1737 0 1
rlabel polysilicon 1052 -1743 1052 -1743 0 3
rlabel polysilicon 1059 -1737 1059 -1737 0 1
rlabel polysilicon 1059 -1743 1059 -1743 0 3
rlabel polysilicon 1066 -1737 1066 -1737 0 1
rlabel polysilicon 1066 -1743 1066 -1743 0 3
rlabel polysilicon 1069 -1743 1069 -1743 0 4
rlabel polysilicon 1073 -1737 1073 -1737 0 1
rlabel polysilicon 1073 -1743 1073 -1743 0 3
rlabel polysilicon 1080 -1737 1080 -1737 0 1
rlabel polysilicon 1080 -1743 1080 -1743 0 3
rlabel polysilicon 1087 -1737 1087 -1737 0 1
rlabel polysilicon 1087 -1743 1087 -1743 0 3
rlabel polysilicon 1094 -1737 1094 -1737 0 1
rlabel polysilicon 1094 -1743 1094 -1743 0 3
rlabel polysilicon 1101 -1737 1101 -1737 0 1
rlabel polysilicon 1101 -1743 1101 -1743 0 3
rlabel polysilicon 1108 -1737 1108 -1737 0 1
rlabel polysilicon 1108 -1743 1108 -1743 0 3
rlabel polysilicon 1115 -1737 1115 -1737 0 1
rlabel polysilicon 1118 -1737 1118 -1737 0 2
rlabel polysilicon 1115 -1743 1115 -1743 0 3
rlabel polysilicon 1122 -1737 1122 -1737 0 1
rlabel polysilicon 1122 -1743 1122 -1743 0 3
rlabel polysilicon 1129 -1737 1129 -1737 0 1
rlabel polysilicon 1129 -1743 1129 -1743 0 3
rlabel polysilicon 1136 -1737 1136 -1737 0 1
rlabel polysilicon 1136 -1743 1136 -1743 0 3
rlabel polysilicon 1143 -1737 1143 -1737 0 1
rlabel polysilicon 1143 -1743 1143 -1743 0 3
rlabel polysilicon 1150 -1737 1150 -1737 0 1
rlabel polysilicon 1150 -1743 1150 -1743 0 3
rlabel polysilicon 1157 -1737 1157 -1737 0 1
rlabel polysilicon 1157 -1743 1157 -1743 0 3
rlabel polysilicon 1164 -1737 1164 -1737 0 1
rlabel polysilicon 1164 -1743 1164 -1743 0 3
rlabel polysilicon 1171 -1737 1171 -1737 0 1
rlabel polysilicon 1171 -1743 1171 -1743 0 3
rlabel polysilicon 1178 -1737 1178 -1737 0 1
rlabel polysilicon 1178 -1743 1178 -1743 0 3
rlabel polysilicon 1185 -1737 1185 -1737 0 1
rlabel polysilicon 1185 -1743 1185 -1743 0 3
rlabel polysilicon 1192 -1737 1192 -1737 0 1
rlabel polysilicon 1192 -1743 1192 -1743 0 3
rlabel polysilicon 1199 -1737 1199 -1737 0 1
rlabel polysilicon 1199 -1743 1199 -1743 0 3
rlabel polysilicon 1206 -1737 1206 -1737 0 1
rlabel polysilicon 1206 -1743 1206 -1743 0 3
rlabel polysilicon 1213 -1737 1213 -1737 0 1
rlabel polysilicon 1213 -1743 1213 -1743 0 3
rlabel polysilicon 1220 -1737 1220 -1737 0 1
rlabel polysilicon 1220 -1743 1220 -1743 0 3
rlabel polysilicon 1227 -1737 1227 -1737 0 1
rlabel polysilicon 1227 -1743 1227 -1743 0 3
rlabel polysilicon 1234 -1737 1234 -1737 0 1
rlabel polysilicon 1234 -1743 1234 -1743 0 3
rlabel polysilicon 1241 -1737 1241 -1737 0 1
rlabel polysilicon 1241 -1743 1241 -1743 0 3
rlabel polysilicon 1251 -1737 1251 -1737 0 2
rlabel polysilicon 1248 -1743 1248 -1743 0 3
rlabel polysilicon 1251 -1743 1251 -1743 0 4
rlabel polysilicon 1255 -1737 1255 -1737 0 1
rlabel polysilicon 1255 -1743 1255 -1743 0 3
rlabel polysilicon 1262 -1737 1262 -1737 0 1
rlabel polysilicon 1262 -1743 1262 -1743 0 3
rlabel polysilicon 1269 -1737 1269 -1737 0 1
rlabel polysilicon 1269 -1743 1269 -1743 0 3
rlabel polysilicon 1276 -1737 1276 -1737 0 1
rlabel polysilicon 1276 -1743 1276 -1743 0 3
rlabel polysilicon 1283 -1737 1283 -1737 0 1
rlabel polysilicon 1283 -1743 1283 -1743 0 3
rlabel polysilicon 1290 -1737 1290 -1737 0 1
rlabel polysilicon 1290 -1743 1290 -1743 0 3
rlabel polysilicon 1297 -1737 1297 -1737 0 1
rlabel polysilicon 1297 -1743 1297 -1743 0 3
rlabel polysilicon 1304 -1737 1304 -1737 0 1
rlabel polysilicon 1304 -1743 1304 -1743 0 3
rlabel polysilicon 1311 -1737 1311 -1737 0 1
rlabel polysilicon 1311 -1743 1311 -1743 0 3
rlabel polysilicon 1318 -1737 1318 -1737 0 1
rlabel polysilicon 1318 -1743 1318 -1743 0 3
rlabel polysilicon 1325 -1737 1325 -1737 0 1
rlabel polysilicon 1325 -1743 1325 -1743 0 3
rlabel polysilicon 1332 -1737 1332 -1737 0 1
rlabel polysilicon 1332 -1743 1332 -1743 0 3
rlabel polysilicon 1339 -1737 1339 -1737 0 1
rlabel polysilicon 1339 -1743 1339 -1743 0 3
rlabel polysilicon 1346 -1737 1346 -1737 0 1
rlabel polysilicon 1346 -1743 1346 -1743 0 3
rlabel polysilicon 1353 -1737 1353 -1737 0 1
rlabel polysilicon 1353 -1743 1353 -1743 0 3
rlabel polysilicon 1360 -1737 1360 -1737 0 1
rlabel polysilicon 1360 -1743 1360 -1743 0 3
rlabel polysilicon 1367 -1737 1367 -1737 0 1
rlabel polysilicon 1367 -1743 1367 -1743 0 3
rlabel polysilicon 1374 -1737 1374 -1737 0 1
rlabel polysilicon 1374 -1743 1374 -1743 0 3
rlabel polysilicon 1381 -1737 1381 -1737 0 1
rlabel polysilicon 1384 -1737 1384 -1737 0 2
rlabel polysilicon 1381 -1743 1381 -1743 0 3
rlabel polysilicon 1388 -1737 1388 -1737 0 1
rlabel polysilicon 1388 -1743 1388 -1743 0 3
rlabel polysilicon 1395 -1737 1395 -1737 0 1
rlabel polysilicon 1395 -1743 1395 -1743 0 3
rlabel polysilicon 1402 -1737 1402 -1737 0 1
rlabel polysilicon 1402 -1743 1402 -1743 0 3
rlabel polysilicon 1409 -1737 1409 -1737 0 1
rlabel polysilicon 1409 -1743 1409 -1743 0 3
rlabel polysilicon 1416 -1737 1416 -1737 0 1
rlabel polysilicon 1416 -1743 1416 -1743 0 3
rlabel polysilicon 1423 -1737 1423 -1737 0 1
rlabel polysilicon 1423 -1743 1423 -1743 0 3
rlabel polysilicon 1430 -1737 1430 -1737 0 1
rlabel polysilicon 1430 -1743 1430 -1743 0 3
rlabel polysilicon 1437 -1737 1437 -1737 0 1
rlabel polysilicon 1437 -1743 1437 -1743 0 3
rlabel polysilicon 1444 -1737 1444 -1737 0 1
rlabel polysilicon 1444 -1743 1444 -1743 0 3
rlabel polysilicon 1451 -1737 1451 -1737 0 1
rlabel polysilicon 1451 -1743 1451 -1743 0 3
rlabel polysilicon 1458 -1737 1458 -1737 0 1
rlabel polysilicon 1458 -1743 1458 -1743 0 3
rlabel polysilicon 1465 -1737 1465 -1737 0 1
rlabel polysilicon 1465 -1743 1465 -1743 0 3
rlabel polysilicon 1472 -1737 1472 -1737 0 1
rlabel polysilicon 1472 -1743 1472 -1743 0 3
rlabel polysilicon 1479 -1737 1479 -1737 0 1
rlabel polysilicon 1479 -1743 1479 -1743 0 3
rlabel polysilicon 1486 -1737 1486 -1737 0 1
rlabel polysilicon 1486 -1743 1486 -1743 0 3
rlabel polysilicon 1493 -1737 1493 -1737 0 1
rlabel polysilicon 1493 -1743 1493 -1743 0 3
rlabel polysilicon 1500 -1737 1500 -1737 0 1
rlabel polysilicon 1500 -1743 1500 -1743 0 3
rlabel polysilicon 1507 -1737 1507 -1737 0 1
rlabel polysilicon 1507 -1743 1507 -1743 0 3
rlabel polysilicon 1514 -1737 1514 -1737 0 1
rlabel polysilicon 1514 -1743 1514 -1743 0 3
rlabel polysilicon 1521 -1737 1521 -1737 0 1
rlabel polysilicon 1521 -1743 1521 -1743 0 3
rlabel polysilicon 1528 -1737 1528 -1737 0 1
rlabel polysilicon 1528 -1743 1528 -1743 0 3
rlabel polysilicon 1535 -1737 1535 -1737 0 1
rlabel polysilicon 1535 -1743 1535 -1743 0 3
rlabel polysilicon 1542 -1737 1542 -1737 0 1
rlabel polysilicon 1542 -1743 1542 -1743 0 3
rlabel polysilicon 1549 -1737 1549 -1737 0 1
rlabel polysilicon 1549 -1743 1549 -1743 0 3
rlabel polysilicon 1556 -1737 1556 -1737 0 1
rlabel polysilicon 1556 -1743 1556 -1743 0 3
rlabel polysilicon 1563 -1737 1563 -1737 0 1
rlabel polysilicon 1563 -1743 1563 -1743 0 3
rlabel polysilicon 1570 -1737 1570 -1737 0 1
rlabel polysilicon 1570 -1743 1570 -1743 0 3
rlabel polysilicon 1577 -1737 1577 -1737 0 1
rlabel polysilicon 1577 -1743 1577 -1743 0 3
rlabel polysilicon 1584 -1737 1584 -1737 0 1
rlabel polysilicon 1584 -1743 1584 -1743 0 3
rlabel polysilicon 1591 -1737 1591 -1737 0 1
rlabel polysilicon 1591 -1743 1591 -1743 0 3
rlabel polysilicon 1598 -1737 1598 -1737 0 1
rlabel polysilicon 1598 -1743 1598 -1743 0 3
rlabel polysilicon 1605 -1737 1605 -1737 0 1
rlabel polysilicon 1605 -1743 1605 -1743 0 3
rlabel polysilicon 1612 -1737 1612 -1737 0 1
rlabel polysilicon 1612 -1743 1612 -1743 0 3
rlabel polysilicon 1619 -1737 1619 -1737 0 1
rlabel polysilicon 1619 -1743 1619 -1743 0 3
rlabel polysilicon 1626 -1737 1626 -1737 0 1
rlabel polysilicon 1626 -1743 1626 -1743 0 3
rlabel polysilicon 1633 -1737 1633 -1737 0 1
rlabel polysilicon 1633 -1743 1633 -1743 0 3
rlabel polysilicon 1640 -1737 1640 -1737 0 1
rlabel polysilicon 1640 -1743 1640 -1743 0 3
rlabel polysilicon 1647 -1737 1647 -1737 0 1
rlabel polysilicon 1647 -1743 1647 -1743 0 3
rlabel polysilicon 1654 -1737 1654 -1737 0 1
rlabel polysilicon 1654 -1743 1654 -1743 0 3
rlabel polysilicon 1661 -1737 1661 -1737 0 1
rlabel polysilicon 1661 -1743 1661 -1743 0 3
rlabel polysilicon 1668 -1737 1668 -1737 0 1
rlabel polysilicon 1668 -1743 1668 -1743 0 3
rlabel polysilicon 1675 -1737 1675 -1737 0 1
rlabel polysilicon 1675 -1743 1675 -1743 0 3
rlabel polysilicon 1682 -1737 1682 -1737 0 1
rlabel polysilicon 1682 -1743 1682 -1743 0 3
rlabel polysilicon 1689 -1737 1689 -1737 0 1
rlabel polysilicon 1689 -1743 1689 -1743 0 3
rlabel polysilicon 1696 -1737 1696 -1737 0 1
rlabel polysilicon 1696 -1743 1696 -1743 0 3
rlabel polysilicon 1703 -1737 1703 -1737 0 1
rlabel polysilicon 1703 -1743 1703 -1743 0 3
rlabel polysilicon 1710 -1737 1710 -1737 0 1
rlabel polysilicon 1710 -1743 1710 -1743 0 3
rlabel polysilicon 1717 -1737 1717 -1737 0 1
rlabel polysilicon 1717 -1743 1717 -1743 0 3
rlabel polysilicon 1724 -1737 1724 -1737 0 1
rlabel polysilicon 1724 -1743 1724 -1743 0 3
rlabel polysilicon 1731 -1737 1731 -1737 0 1
rlabel polysilicon 1731 -1743 1731 -1743 0 3
rlabel polysilicon 1738 -1737 1738 -1737 0 1
rlabel polysilicon 1738 -1743 1738 -1743 0 3
rlabel polysilicon 1748 -1737 1748 -1737 0 2
rlabel polysilicon 1745 -1743 1745 -1743 0 3
rlabel polysilicon 1748 -1743 1748 -1743 0 4
rlabel polysilicon 1752 -1737 1752 -1737 0 1
rlabel polysilicon 1752 -1743 1752 -1743 0 3
rlabel polysilicon 1759 -1737 1759 -1737 0 1
rlabel polysilicon 1759 -1743 1759 -1743 0 3
rlabel polysilicon 1766 -1737 1766 -1737 0 1
rlabel polysilicon 1766 -1743 1766 -1743 0 3
rlabel polysilicon 1773 -1737 1773 -1737 0 1
rlabel polysilicon 1773 -1743 1773 -1743 0 3
rlabel polysilicon 1780 -1737 1780 -1737 0 1
rlabel polysilicon 1780 -1743 1780 -1743 0 3
rlabel polysilicon 30 -1884 30 -1884 0 1
rlabel polysilicon 30 -1890 30 -1890 0 3
rlabel polysilicon 37 -1884 37 -1884 0 1
rlabel polysilicon 37 -1890 37 -1890 0 3
rlabel polysilicon 44 -1884 44 -1884 0 1
rlabel polysilicon 44 -1890 44 -1890 0 3
rlabel polysilicon 51 -1884 51 -1884 0 1
rlabel polysilicon 51 -1890 51 -1890 0 3
rlabel polysilicon 58 -1884 58 -1884 0 1
rlabel polysilicon 58 -1890 58 -1890 0 3
rlabel polysilicon 65 -1884 65 -1884 0 1
rlabel polysilicon 65 -1890 65 -1890 0 3
rlabel polysilicon 72 -1884 72 -1884 0 1
rlabel polysilicon 72 -1890 72 -1890 0 3
rlabel polysilicon 79 -1884 79 -1884 0 1
rlabel polysilicon 79 -1890 79 -1890 0 3
rlabel polysilicon 86 -1884 86 -1884 0 1
rlabel polysilicon 86 -1890 86 -1890 0 3
rlabel polysilicon 93 -1884 93 -1884 0 1
rlabel polysilicon 93 -1890 93 -1890 0 3
rlabel polysilicon 100 -1884 100 -1884 0 1
rlabel polysilicon 100 -1890 100 -1890 0 3
rlabel polysilicon 107 -1884 107 -1884 0 1
rlabel polysilicon 110 -1884 110 -1884 0 2
rlabel polysilicon 107 -1890 107 -1890 0 3
rlabel polysilicon 110 -1890 110 -1890 0 4
rlabel polysilicon 114 -1884 114 -1884 0 1
rlabel polysilicon 114 -1890 114 -1890 0 3
rlabel polysilicon 121 -1884 121 -1884 0 1
rlabel polysilicon 121 -1890 121 -1890 0 3
rlabel polysilicon 128 -1884 128 -1884 0 1
rlabel polysilicon 128 -1890 128 -1890 0 3
rlabel polysilicon 135 -1884 135 -1884 0 1
rlabel polysilicon 135 -1890 135 -1890 0 3
rlabel polysilicon 142 -1884 142 -1884 0 1
rlabel polysilicon 142 -1890 142 -1890 0 3
rlabel polysilicon 149 -1884 149 -1884 0 1
rlabel polysilicon 149 -1890 149 -1890 0 3
rlabel polysilicon 156 -1884 156 -1884 0 1
rlabel polysilicon 159 -1884 159 -1884 0 2
rlabel polysilicon 156 -1890 156 -1890 0 3
rlabel polysilicon 159 -1890 159 -1890 0 4
rlabel polysilicon 163 -1884 163 -1884 0 1
rlabel polysilicon 163 -1890 163 -1890 0 3
rlabel polysilicon 170 -1884 170 -1884 0 1
rlabel polysilicon 170 -1890 170 -1890 0 3
rlabel polysilicon 177 -1884 177 -1884 0 1
rlabel polysilicon 180 -1884 180 -1884 0 2
rlabel polysilicon 177 -1890 177 -1890 0 3
rlabel polysilicon 180 -1890 180 -1890 0 4
rlabel polysilicon 184 -1884 184 -1884 0 1
rlabel polysilicon 184 -1890 184 -1890 0 3
rlabel polysilicon 191 -1884 191 -1884 0 1
rlabel polysilicon 191 -1890 191 -1890 0 3
rlabel polysilicon 198 -1884 198 -1884 0 1
rlabel polysilicon 198 -1890 198 -1890 0 3
rlabel polysilicon 205 -1884 205 -1884 0 1
rlabel polysilicon 208 -1884 208 -1884 0 2
rlabel polysilicon 208 -1890 208 -1890 0 4
rlabel polysilicon 212 -1884 212 -1884 0 1
rlabel polysilicon 212 -1890 212 -1890 0 3
rlabel polysilicon 219 -1884 219 -1884 0 1
rlabel polysilicon 219 -1890 219 -1890 0 3
rlabel polysilicon 226 -1884 226 -1884 0 1
rlabel polysilicon 226 -1890 226 -1890 0 3
rlabel polysilicon 233 -1884 233 -1884 0 1
rlabel polysilicon 233 -1890 233 -1890 0 3
rlabel polysilicon 240 -1884 240 -1884 0 1
rlabel polysilicon 240 -1890 240 -1890 0 3
rlabel polysilicon 247 -1884 247 -1884 0 1
rlabel polysilicon 250 -1884 250 -1884 0 2
rlabel polysilicon 247 -1890 247 -1890 0 3
rlabel polysilicon 250 -1890 250 -1890 0 4
rlabel polysilicon 254 -1884 254 -1884 0 1
rlabel polysilicon 254 -1890 254 -1890 0 3
rlabel polysilicon 264 -1884 264 -1884 0 2
rlabel polysilicon 264 -1890 264 -1890 0 4
rlabel polysilicon 268 -1884 268 -1884 0 1
rlabel polysilicon 268 -1890 268 -1890 0 3
rlabel polysilicon 275 -1884 275 -1884 0 1
rlabel polysilicon 275 -1890 275 -1890 0 3
rlabel polysilicon 282 -1884 282 -1884 0 1
rlabel polysilicon 282 -1890 282 -1890 0 3
rlabel polysilicon 289 -1884 289 -1884 0 1
rlabel polysilicon 289 -1890 289 -1890 0 3
rlabel polysilicon 296 -1884 296 -1884 0 1
rlabel polysilicon 296 -1890 296 -1890 0 3
rlabel polysilicon 303 -1884 303 -1884 0 1
rlabel polysilicon 303 -1890 303 -1890 0 3
rlabel polysilicon 310 -1884 310 -1884 0 1
rlabel polysilicon 310 -1890 310 -1890 0 3
rlabel polysilicon 317 -1884 317 -1884 0 1
rlabel polysilicon 317 -1890 317 -1890 0 3
rlabel polysilicon 324 -1884 324 -1884 0 1
rlabel polysilicon 324 -1890 324 -1890 0 3
rlabel polysilicon 331 -1884 331 -1884 0 1
rlabel polysilicon 331 -1890 331 -1890 0 3
rlabel polysilicon 338 -1884 338 -1884 0 1
rlabel polysilicon 341 -1884 341 -1884 0 2
rlabel polysilicon 341 -1890 341 -1890 0 4
rlabel polysilicon 345 -1884 345 -1884 0 1
rlabel polysilicon 345 -1890 345 -1890 0 3
rlabel polysilicon 352 -1884 352 -1884 0 1
rlabel polysilicon 352 -1890 352 -1890 0 3
rlabel polysilicon 359 -1884 359 -1884 0 1
rlabel polysilicon 359 -1890 359 -1890 0 3
rlabel polysilicon 366 -1884 366 -1884 0 1
rlabel polysilicon 366 -1890 366 -1890 0 3
rlabel polysilicon 373 -1884 373 -1884 0 1
rlabel polysilicon 373 -1890 373 -1890 0 3
rlabel polysilicon 380 -1884 380 -1884 0 1
rlabel polysilicon 380 -1890 380 -1890 0 3
rlabel polysilicon 387 -1884 387 -1884 0 1
rlabel polysilicon 387 -1890 387 -1890 0 3
rlabel polysilicon 394 -1884 394 -1884 0 1
rlabel polysilicon 394 -1890 394 -1890 0 3
rlabel polysilicon 401 -1884 401 -1884 0 1
rlabel polysilicon 401 -1890 401 -1890 0 3
rlabel polysilicon 408 -1884 408 -1884 0 1
rlabel polysilicon 408 -1890 408 -1890 0 3
rlabel polysilicon 415 -1884 415 -1884 0 1
rlabel polysilicon 415 -1890 415 -1890 0 3
rlabel polysilicon 422 -1884 422 -1884 0 1
rlabel polysilicon 422 -1890 422 -1890 0 3
rlabel polysilicon 429 -1884 429 -1884 0 1
rlabel polysilicon 429 -1890 429 -1890 0 3
rlabel polysilicon 436 -1884 436 -1884 0 1
rlabel polysilicon 436 -1890 436 -1890 0 3
rlabel polysilicon 443 -1884 443 -1884 0 1
rlabel polysilicon 446 -1884 446 -1884 0 2
rlabel polysilicon 443 -1890 443 -1890 0 3
rlabel polysilicon 446 -1890 446 -1890 0 4
rlabel polysilicon 450 -1884 450 -1884 0 1
rlabel polysilicon 450 -1890 450 -1890 0 3
rlabel polysilicon 457 -1884 457 -1884 0 1
rlabel polysilicon 457 -1890 457 -1890 0 3
rlabel polysilicon 464 -1884 464 -1884 0 1
rlabel polysilicon 467 -1884 467 -1884 0 2
rlabel polysilicon 464 -1890 464 -1890 0 3
rlabel polysilicon 467 -1890 467 -1890 0 4
rlabel polysilicon 471 -1884 471 -1884 0 1
rlabel polysilicon 474 -1884 474 -1884 0 2
rlabel polysilicon 471 -1890 471 -1890 0 3
rlabel polysilicon 474 -1890 474 -1890 0 4
rlabel polysilicon 478 -1884 478 -1884 0 1
rlabel polysilicon 478 -1890 478 -1890 0 3
rlabel polysilicon 485 -1884 485 -1884 0 1
rlabel polysilicon 492 -1884 492 -1884 0 1
rlabel polysilicon 492 -1890 492 -1890 0 3
rlabel polysilicon 502 -1884 502 -1884 0 2
rlabel polysilicon 506 -1884 506 -1884 0 1
rlabel polysilicon 506 -1890 506 -1890 0 3
rlabel polysilicon 513 -1884 513 -1884 0 1
rlabel polysilicon 513 -1890 513 -1890 0 3
rlabel polysilicon 520 -1884 520 -1884 0 1
rlabel polysilicon 520 -1890 520 -1890 0 3
rlabel polysilicon 527 -1884 527 -1884 0 1
rlabel polysilicon 527 -1890 527 -1890 0 3
rlabel polysilicon 530 -1890 530 -1890 0 4
rlabel polysilicon 534 -1884 534 -1884 0 1
rlabel polysilicon 534 -1890 534 -1890 0 3
rlabel polysilicon 541 -1884 541 -1884 0 1
rlabel polysilicon 541 -1890 541 -1890 0 3
rlabel polysilicon 548 -1884 548 -1884 0 1
rlabel polysilicon 548 -1890 548 -1890 0 3
rlabel polysilicon 555 -1884 555 -1884 0 1
rlabel polysilicon 555 -1890 555 -1890 0 3
rlabel polysilicon 562 -1884 562 -1884 0 1
rlabel polysilicon 562 -1890 562 -1890 0 3
rlabel polysilicon 569 -1884 569 -1884 0 1
rlabel polysilicon 569 -1890 569 -1890 0 3
rlabel polysilicon 572 -1890 572 -1890 0 4
rlabel polysilicon 576 -1884 576 -1884 0 1
rlabel polysilicon 576 -1890 576 -1890 0 3
rlabel polysilicon 583 -1884 583 -1884 0 1
rlabel polysilicon 583 -1890 583 -1890 0 3
rlabel polysilicon 590 -1884 590 -1884 0 1
rlabel polysilicon 590 -1890 590 -1890 0 3
rlabel polysilicon 597 -1884 597 -1884 0 1
rlabel polysilicon 597 -1890 597 -1890 0 3
rlabel polysilicon 604 -1884 604 -1884 0 1
rlabel polysilicon 604 -1890 604 -1890 0 3
rlabel polysilicon 611 -1884 611 -1884 0 1
rlabel polysilicon 611 -1890 611 -1890 0 3
rlabel polysilicon 618 -1884 618 -1884 0 1
rlabel polysilicon 618 -1890 618 -1890 0 3
rlabel polysilicon 625 -1884 625 -1884 0 1
rlabel polysilicon 625 -1890 625 -1890 0 3
rlabel polysilicon 632 -1884 632 -1884 0 1
rlabel polysilicon 632 -1890 632 -1890 0 3
rlabel polysilicon 639 -1884 639 -1884 0 1
rlabel polysilicon 639 -1890 639 -1890 0 3
rlabel polysilicon 649 -1884 649 -1884 0 2
rlabel polysilicon 646 -1890 646 -1890 0 3
rlabel polysilicon 649 -1890 649 -1890 0 4
rlabel polysilicon 653 -1884 653 -1884 0 1
rlabel polysilicon 656 -1884 656 -1884 0 2
rlabel polysilicon 653 -1890 653 -1890 0 3
rlabel polysilicon 656 -1890 656 -1890 0 4
rlabel polysilicon 660 -1884 660 -1884 0 1
rlabel polysilicon 660 -1890 660 -1890 0 3
rlabel polysilicon 667 -1884 667 -1884 0 1
rlabel polysilicon 667 -1890 667 -1890 0 3
rlabel polysilicon 674 -1884 674 -1884 0 1
rlabel polysilicon 674 -1890 674 -1890 0 3
rlabel polysilicon 681 -1884 681 -1884 0 1
rlabel polysilicon 681 -1890 681 -1890 0 3
rlabel polysilicon 688 -1884 688 -1884 0 1
rlabel polysilicon 688 -1890 688 -1890 0 3
rlabel polysilicon 695 -1884 695 -1884 0 1
rlabel polysilicon 695 -1890 695 -1890 0 3
rlabel polysilicon 702 -1884 702 -1884 0 1
rlabel polysilicon 702 -1890 702 -1890 0 3
rlabel polysilicon 709 -1884 709 -1884 0 1
rlabel polysilicon 709 -1890 709 -1890 0 3
rlabel polysilicon 716 -1884 716 -1884 0 1
rlabel polysilicon 716 -1890 716 -1890 0 3
rlabel polysilicon 723 -1884 723 -1884 0 1
rlabel polysilicon 723 -1890 723 -1890 0 3
rlabel polysilicon 730 -1884 730 -1884 0 1
rlabel polysilicon 730 -1890 730 -1890 0 3
rlabel polysilicon 737 -1884 737 -1884 0 1
rlabel polysilicon 737 -1890 737 -1890 0 3
rlabel polysilicon 744 -1884 744 -1884 0 1
rlabel polysilicon 744 -1890 744 -1890 0 3
rlabel polysilicon 751 -1884 751 -1884 0 1
rlabel polysilicon 751 -1890 751 -1890 0 3
rlabel polysilicon 758 -1884 758 -1884 0 1
rlabel polysilicon 758 -1890 758 -1890 0 3
rlabel polysilicon 765 -1884 765 -1884 0 1
rlabel polysilicon 765 -1890 765 -1890 0 3
rlabel polysilicon 772 -1884 772 -1884 0 1
rlabel polysilicon 772 -1890 772 -1890 0 3
rlabel polysilicon 779 -1884 779 -1884 0 1
rlabel polysilicon 779 -1890 779 -1890 0 3
rlabel polysilicon 786 -1884 786 -1884 0 1
rlabel polysilicon 786 -1890 786 -1890 0 3
rlabel polysilicon 793 -1884 793 -1884 0 1
rlabel polysilicon 793 -1890 793 -1890 0 3
rlabel polysilicon 800 -1884 800 -1884 0 1
rlabel polysilicon 800 -1890 800 -1890 0 3
rlabel polysilicon 810 -1884 810 -1884 0 2
rlabel polysilicon 807 -1890 807 -1890 0 3
rlabel polysilicon 810 -1890 810 -1890 0 4
rlabel polysilicon 814 -1884 814 -1884 0 1
rlabel polysilicon 814 -1890 814 -1890 0 3
rlabel polysilicon 821 -1884 821 -1884 0 1
rlabel polysilicon 824 -1884 824 -1884 0 2
rlabel polysilicon 821 -1890 821 -1890 0 3
rlabel polysilicon 824 -1890 824 -1890 0 4
rlabel polysilicon 828 -1884 828 -1884 0 1
rlabel polysilicon 831 -1884 831 -1884 0 2
rlabel polysilicon 831 -1890 831 -1890 0 4
rlabel polysilicon 835 -1884 835 -1884 0 1
rlabel polysilicon 838 -1890 838 -1890 0 4
rlabel polysilicon 842 -1884 842 -1884 0 1
rlabel polysilicon 842 -1890 842 -1890 0 3
rlabel polysilicon 849 -1884 849 -1884 0 1
rlabel polysilicon 849 -1890 849 -1890 0 3
rlabel polysilicon 856 -1884 856 -1884 0 1
rlabel polysilicon 856 -1890 856 -1890 0 3
rlabel polysilicon 863 -1884 863 -1884 0 1
rlabel polysilicon 866 -1884 866 -1884 0 2
rlabel polysilicon 866 -1890 866 -1890 0 4
rlabel polysilicon 870 -1884 870 -1884 0 1
rlabel polysilicon 870 -1890 870 -1890 0 3
rlabel polysilicon 877 -1884 877 -1884 0 1
rlabel polysilicon 877 -1890 877 -1890 0 3
rlabel polysilicon 884 -1884 884 -1884 0 1
rlabel polysilicon 884 -1890 884 -1890 0 3
rlabel polysilicon 891 -1884 891 -1884 0 1
rlabel polysilicon 891 -1890 891 -1890 0 3
rlabel polysilicon 898 -1884 898 -1884 0 1
rlabel polysilicon 898 -1890 898 -1890 0 3
rlabel polysilicon 905 -1884 905 -1884 0 1
rlabel polysilicon 905 -1890 905 -1890 0 3
rlabel polysilicon 908 -1890 908 -1890 0 4
rlabel polysilicon 912 -1884 912 -1884 0 1
rlabel polysilicon 912 -1890 912 -1890 0 3
rlabel polysilicon 919 -1884 919 -1884 0 1
rlabel polysilicon 919 -1890 919 -1890 0 3
rlabel polysilicon 926 -1884 926 -1884 0 1
rlabel polysilicon 929 -1884 929 -1884 0 2
rlabel polysilicon 926 -1890 926 -1890 0 3
rlabel polysilicon 929 -1890 929 -1890 0 4
rlabel polysilicon 933 -1884 933 -1884 0 1
rlabel polysilicon 936 -1884 936 -1884 0 2
rlabel polysilicon 936 -1890 936 -1890 0 4
rlabel polysilicon 940 -1884 940 -1884 0 1
rlabel polysilicon 940 -1890 940 -1890 0 3
rlabel polysilicon 947 -1884 947 -1884 0 1
rlabel polysilicon 947 -1890 947 -1890 0 3
rlabel polysilicon 957 -1890 957 -1890 0 4
rlabel polysilicon 961 -1884 961 -1884 0 1
rlabel polysilicon 961 -1890 961 -1890 0 3
rlabel polysilicon 968 -1884 968 -1884 0 1
rlabel polysilicon 968 -1890 968 -1890 0 3
rlabel polysilicon 975 -1884 975 -1884 0 1
rlabel polysilicon 975 -1890 975 -1890 0 3
rlabel polysilicon 982 -1884 982 -1884 0 1
rlabel polysilicon 985 -1884 985 -1884 0 2
rlabel polysilicon 985 -1890 985 -1890 0 4
rlabel polysilicon 989 -1884 989 -1884 0 1
rlabel polysilicon 989 -1890 989 -1890 0 3
rlabel polysilicon 996 -1884 996 -1884 0 1
rlabel polysilicon 996 -1890 996 -1890 0 3
rlabel polysilicon 1003 -1884 1003 -1884 0 1
rlabel polysilicon 1003 -1890 1003 -1890 0 3
rlabel polysilicon 1010 -1884 1010 -1884 0 1
rlabel polysilicon 1010 -1890 1010 -1890 0 3
rlabel polysilicon 1017 -1884 1017 -1884 0 1
rlabel polysilicon 1017 -1890 1017 -1890 0 3
rlabel polysilicon 1020 -1890 1020 -1890 0 4
rlabel polysilicon 1024 -1884 1024 -1884 0 1
rlabel polysilicon 1027 -1884 1027 -1884 0 2
rlabel polysilicon 1024 -1890 1024 -1890 0 3
rlabel polysilicon 1027 -1890 1027 -1890 0 4
rlabel polysilicon 1031 -1884 1031 -1884 0 1
rlabel polysilicon 1031 -1890 1031 -1890 0 3
rlabel polysilicon 1038 -1884 1038 -1884 0 1
rlabel polysilicon 1041 -1884 1041 -1884 0 2
rlabel polysilicon 1038 -1890 1038 -1890 0 3
rlabel polysilicon 1045 -1884 1045 -1884 0 1
rlabel polysilicon 1048 -1884 1048 -1884 0 2
rlabel polysilicon 1045 -1890 1045 -1890 0 3
rlabel polysilicon 1048 -1890 1048 -1890 0 4
rlabel polysilicon 1052 -1884 1052 -1884 0 1
rlabel polysilicon 1052 -1890 1052 -1890 0 3
rlabel polysilicon 1059 -1884 1059 -1884 0 1
rlabel polysilicon 1059 -1890 1059 -1890 0 3
rlabel polysilicon 1066 -1884 1066 -1884 0 1
rlabel polysilicon 1066 -1890 1066 -1890 0 3
rlabel polysilicon 1073 -1884 1073 -1884 0 1
rlabel polysilicon 1073 -1890 1073 -1890 0 3
rlabel polysilicon 1080 -1884 1080 -1884 0 1
rlabel polysilicon 1080 -1890 1080 -1890 0 3
rlabel polysilicon 1087 -1884 1087 -1884 0 1
rlabel polysilicon 1087 -1890 1087 -1890 0 3
rlabel polysilicon 1094 -1884 1094 -1884 0 1
rlabel polysilicon 1094 -1890 1094 -1890 0 3
rlabel polysilicon 1101 -1884 1101 -1884 0 1
rlabel polysilicon 1101 -1890 1101 -1890 0 3
rlabel polysilicon 1108 -1884 1108 -1884 0 1
rlabel polysilicon 1111 -1884 1111 -1884 0 2
rlabel polysilicon 1108 -1890 1108 -1890 0 3
rlabel polysilicon 1115 -1884 1115 -1884 0 1
rlabel polysilicon 1115 -1890 1115 -1890 0 3
rlabel polysilicon 1122 -1884 1122 -1884 0 1
rlabel polysilicon 1122 -1890 1122 -1890 0 3
rlabel polysilicon 1129 -1884 1129 -1884 0 1
rlabel polysilicon 1129 -1890 1129 -1890 0 3
rlabel polysilicon 1136 -1884 1136 -1884 0 1
rlabel polysilicon 1136 -1890 1136 -1890 0 3
rlabel polysilicon 1143 -1884 1143 -1884 0 1
rlabel polysilicon 1143 -1890 1143 -1890 0 3
rlabel polysilicon 1150 -1884 1150 -1884 0 1
rlabel polysilicon 1153 -1884 1153 -1884 0 2
rlabel polysilicon 1150 -1890 1150 -1890 0 3
rlabel polysilicon 1153 -1890 1153 -1890 0 4
rlabel polysilicon 1157 -1884 1157 -1884 0 1
rlabel polysilicon 1160 -1884 1160 -1884 0 2
rlabel polysilicon 1157 -1890 1157 -1890 0 3
rlabel polysilicon 1160 -1890 1160 -1890 0 4
rlabel polysilicon 1164 -1884 1164 -1884 0 1
rlabel polysilicon 1164 -1890 1164 -1890 0 3
rlabel polysilicon 1171 -1884 1171 -1884 0 1
rlabel polysilicon 1171 -1890 1171 -1890 0 3
rlabel polysilicon 1178 -1884 1178 -1884 0 1
rlabel polysilicon 1178 -1890 1178 -1890 0 3
rlabel polysilicon 1185 -1884 1185 -1884 0 1
rlabel polysilicon 1185 -1890 1185 -1890 0 3
rlabel polysilicon 1192 -1884 1192 -1884 0 1
rlabel polysilicon 1192 -1890 1192 -1890 0 3
rlabel polysilicon 1199 -1884 1199 -1884 0 1
rlabel polysilicon 1199 -1890 1199 -1890 0 3
rlabel polysilicon 1206 -1884 1206 -1884 0 1
rlabel polysilicon 1206 -1890 1206 -1890 0 3
rlabel polysilicon 1213 -1884 1213 -1884 0 1
rlabel polysilicon 1213 -1890 1213 -1890 0 3
rlabel polysilicon 1220 -1884 1220 -1884 0 1
rlabel polysilicon 1220 -1890 1220 -1890 0 3
rlabel polysilicon 1227 -1884 1227 -1884 0 1
rlabel polysilicon 1227 -1890 1227 -1890 0 3
rlabel polysilicon 1234 -1884 1234 -1884 0 1
rlabel polysilicon 1234 -1890 1234 -1890 0 3
rlabel polysilicon 1241 -1884 1241 -1884 0 1
rlabel polysilicon 1241 -1890 1241 -1890 0 3
rlabel polysilicon 1248 -1884 1248 -1884 0 1
rlabel polysilicon 1248 -1890 1248 -1890 0 3
rlabel polysilicon 1255 -1884 1255 -1884 0 1
rlabel polysilicon 1255 -1890 1255 -1890 0 3
rlabel polysilicon 1262 -1884 1262 -1884 0 1
rlabel polysilicon 1262 -1890 1262 -1890 0 3
rlabel polysilicon 1269 -1884 1269 -1884 0 1
rlabel polysilicon 1269 -1890 1269 -1890 0 3
rlabel polysilicon 1276 -1884 1276 -1884 0 1
rlabel polysilicon 1279 -1884 1279 -1884 0 2
rlabel polysilicon 1276 -1890 1276 -1890 0 3
rlabel polysilicon 1279 -1890 1279 -1890 0 4
rlabel polysilicon 1283 -1884 1283 -1884 0 1
rlabel polysilicon 1283 -1890 1283 -1890 0 3
rlabel polysilicon 1290 -1884 1290 -1884 0 1
rlabel polysilicon 1290 -1890 1290 -1890 0 3
rlabel polysilicon 1297 -1884 1297 -1884 0 1
rlabel polysilicon 1297 -1890 1297 -1890 0 3
rlabel polysilicon 1304 -1884 1304 -1884 0 1
rlabel polysilicon 1304 -1890 1304 -1890 0 3
rlabel polysilicon 1311 -1890 1311 -1890 0 3
rlabel polysilicon 1314 -1890 1314 -1890 0 4
rlabel polysilicon 1318 -1884 1318 -1884 0 1
rlabel polysilicon 1318 -1890 1318 -1890 0 3
rlabel polysilicon 1325 -1884 1325 -1884 0 1
rlabel polysilicon 1325 -1890 1325 -1890 0 3
rlabel polysilicon 1332 -1884 1332 -1884 0 1
rlabel polysilicon 1332 -1890 1332 -1890 0 3
rlabel polysilicon 1339 -1884 1339 -1884 0 1
rlabel polysilicon 1339 -1890 1339 -1890 0 3
rlabel polysilicon 1346 -1884 1346 -1884 0 1
rlabel polysilicon 1346 -1890 1346 -1890 0 3
rlabel polysilicon 1353 -1884 1353 -1884 0 1
rlabel polysilicon 1353 -1890 1353 -1890 0 3
rlabel polysilicon 1360 -1884 1360 -1884 0 1
rlabel polysilicon 1360 -1890 1360 -1890 0 3
rlabel polysilicon 1367 -1884 1367 -1884 0 1
rlabel polysilicon 1367 -1890 1367 -1890 0 3
rlabel polysilicon 1374 -1884 1374 -1884 0 1
rlabel polysilicon 1374 -1890 1374 -1890 0 3
rlabel polysilicon 1381 -1884 1381 -1884 0 1
rlabel polysilicon 1381 -1890 1381 -1890 0 3
rlabel polysilicon 1384 -1890 1384 -1890 0 4
rlabel polysilicon 1388 -1884 1388 -1884 0 1
rlabel polysilicon 1388 -1890 1388 -1890 0 3
rlabel polysilicon 1395 -1884 1395 -1884 0 1
rlabel polysilicon 1395 -1890 1395 -1890 0 3
rlabel polysilicon 1402 -1884 1402 -1884 0 1
rlabel polysilicon 1402 -1890 1402 -1890 0 3
rlabel polysilicon 1409 -1884 1409 -1884 0 1
rlabel polysilicon 1409 -1890 1409 -1890 0 3
rlabel polysilicon 1416 -1884 1416 -1884 0 1
rlabel polysilicon 1416 -1890 1416 -1890 0 3
rlabel polysilicon 1423 -1884 1423 -1884 0 1
rlabel polysilicon 1423 -1890 1423 -1890 0 3
rlabel polysilicon 1430 -1884 1430 -1884 0 1
rlabel polysilicon 1430 -1890 1430 -1890 0 3
rlabel polysilicon 1437 -1884 1437 -1884 0 1
rlabel polysilicon 1437 -1890 1437 -1890 0 3
rlabel polysilicon 1444 -1884 1444 -1884 0 1
rlabel polysilicon 1444 -1890 1444 -1890 0 3
rlabel polysilicon 1451 -1884 1451 -1884 0 1
rlabel polysilicon 1451 -1890 1451 -1890 0 3
rlabel polysilicon 1458 -1884 1458 -1884 0 1
rlabel polysilicon 1458 -1890 1458 -1890 0 3
rlabel polysilicon 1465 -1884 1465 -1884 0 1
rlabel polysilicon 1465 -1890 1465 -1890 0 3
rlabel polysilicon 1472 -1884 1472 -1884 0 1
rlabel polysilicon 1472 -1890 1472 -1890 0 3
rlabel polysilicon 1479 -1884 1479 -1884 0 1
rlabel polysilicon 1479 -1890 1479 -1890 0 3
rlabel polysilicon 1486 -1884 1486 -1884 0 1
rlabel polysilicon 1486 -1890 1486 -1890 0 3
rlabel polysilicon 1493 -1884 1493 -1884 0 1
rlabel polysilicon 1493 -1890 1493 -1890 0 3
rlabel polysilicon 1500 -1884 1500 -1884 0 1
rlabel polysilicon 1500 -1890 1500 -1890 0 3
rlabel polysilicon 1507 -1884 1507 -1884 0 1
rlabel polysilicon 1507 -1890 1507 -1890 0 3
rlabel polysilicon 1514 -1884 1514 -1884 0 1
rlabel polysilicon 1514 -1890 1514 -1890 0 3
rlabel polysilicon 1521 -1884 1521 -1884 0 1
rlabel polysilicon 1521 -1890 1521 -1890 0 3
rlabel polysilicon 1528 -1884 1528 -1884 0 1
rlabel polysilicon 1528 -1890 1528 -1890 0 3
rlabel polysilicon 1535 -1884 1535 -1884 0 1
rlabel polysilicon 1535 -1890 1535 -1890 0 3
rlabel polysilicon 1542 -1884 1542 -1884 0 1
rlabel polysilicon 1542 -1890 1542 -1890 0 3
rlabel polysilicon 1549 -1884 1549 -1884 0 1
rlabel polysilicon 1549 -1890 1549 -1890 0 3
rlabel polysilicon 1556 -1884 1556 -1884 0 1
rlabel polysilicon 1556 -1890 1556 -1890 0 3
rlabel polysilicon 1563 -1884 1563 -1884 0 1
rlabel polysilicon 1563 -1890 1563 -1890 0 3
rlabel polysilicon 1570 -1884 1570 -1884 0 1
rlabel polysilicon 1570 -1890 1570 -1890 0 3
rlabel polysilicon 1577 -1884 1577 -1884 0 1
rlabel polysilicon 1577 -1890 1577 -1890 0 3
rlabel polysilicon 1584 -1884 1584 -1884 0 1
rlabel polysilicon 1584 -1890 1584 -1890 0 3
rlabel polysilicon 1591 -1884 1591 -1884 0 1
rlabel polysilicon 1591 -1890 1591 -1890 0 3
rlabel polysilicon 1598 -1884 1598 -1884 0 1
rlabel polysilicon 1598 -1890 1598 -1890 0 3
rlabel polysilicon 1605 -1884 1605 -1884 0 1
rlabel polysilicon 1605 -1890 1605 -1890 0 3
rlabel polysilicon 1612 -1884 1612 -1884 0 1
rlabel polysilicon 1612 -1890 1612 -1890 0 3
rlabel polysilicon 1619 -1884 1619 -1884 0 1
rlabel polysilicon 1619 -1890 1619 -1890 0 3
rlabel polysilicon 1626 -1884 1626 -1884 0 1
rlabel polysilicon 1626 -1890 1626 -1890 0 3
rlabel polysilicon 1633 -1884 1633 -1884 0 1
rlabel polysilicon 1633 -1890 1633 -1890 0 3
rlabel polysilicon 1640 -1884 1640 -1884 0 1
rlabel polysilicon 1640 -1890 1640 -1890 0 3
rlabel polysilicon 1647 -1884 1647 -1884 0 1
rlabel polysilicon 1647 -1890 1647 -1890 0 3
rlabel polysilicon 1654 -1884 1654 -1884 0 1
rlabel polysilicon 1654 -1890 1654 -1890 0 3
rlabel polysilicon 1661 -1884 1661 -1884 0 1
rlabel polysilicon 1661 -1890 1661 -1890 0 3
rlabel polysilicon 1668 -1884 1668 -1884 0 1
rlabel polysilicon 1668 -1890 1668 -1890 0 3
rlabel polysilicon 1675 -1884 1675 -1884 0 1
rlabel polysilicon 1675 -1890 1675 -1890 0 3
rlabel polysilicon 1682 -1884 1682 -1884 0 1
rlabel polysilicon 1682 -1890 1682 -1890 0 3
rlabel polysilicon 1689 -1884 1689 -1884 0 1
rlabel polysilicon 1689 -1890 1689 -1890 0 3
rlabel polysilicon 1696 -1884 1696 -1884 0 1
rlabel polysilicon 1696 -1890 1696 -1890 0 3
rlabel polysilicon 1703 -1884 1703 -1884 0 1
rlabel polysilicon 1703 -1890 1703 -1890 0 3
rlabel polysilicon 1710 -1884 1710 -1884 0 1
rlabel polysilicon 1710 -1890 1710 -1890 0 3
rlabel polysilicon 1717 -1884 1717 -1884 0 1
rlabel polysilicon 1717 -1890 1717 -1890 0 3
rlabel polysilicon 1724 -1884 1724 -1884 0 1
rlabel polysilicon 1724 -1890 1724 -1890 0 3
rlabel polysilicon 1731 -1884 1731 -1884 0 1
rlabel polysilicon 1731 -1890 1731 -1890 0 3
rlabel polysilicon 1738 -1884 1738 -1884 0 1
rlabel polysilicon 1738 -1890 1738 -1890 0 3
rlabel polysilicon 1745 -1884 1745 -1884 0 1
rlabel polysilicon 1745 -1890 1745 -1890 0 3
rlabel polysilicon 1752 -1884 1752 -1884 0 1
rlabel polysilicon 1752 -1890 1752 -1890 0 3
rlabel polysilicon 1759 -1884 1759 -1884 0 1
rlabel polysilicon 1759 -1890 1759 -1890 0 3
rlabel polysilicon 1766 -1884 1766 -1884 0 1
rlabel polysilicon 1766 -1890 1766 -1890 0 3
rlabel polysilicon 1773 -1884 1773 -1884 0 1
rlabel polysilicon 1776 -1884 1776 -1884 0 2
rlabel polysilicon 1773 -1890 1773 -1890 0 3
rlabel polysilicon 1776 -1890 1776 -1890 0 4
rlabel polysilicon 1780 -1884 1780 -1884 0 1
rlabel polysilicon 1780 -1890 1780 -1890 0 3
rlabel polysilicon 1787 -1884 1787 -1884 0 1
rlabel polysilicon 1787 -1890 1787 -1890 0 3
rlabel polysilicon 1794 -1884 1794 -1884 0 1
rlabel polysilicon 1794 -1890 1794 -1890 0 3
rlabel polysilicon 1801 -1884 1801 -1884 0 1
rlabel polysilicon 1804 -1884 1804 -1884 0 2
rlabel polysilicon 1801 -1890 1801 -1890 0 3
rlabel polysilicon 1804 -1890 1804 -1890 0 4
rlabel polysilicon 1808 -1884 1808 -1884 0 1
rlabel polysilicon 1808 -1890 1808 -1890 0 3
rlabel polysilicon 1815 -1884 1815 -1884 0 1
rlabel polysilicon 1815 -1890 1815 -1890 0 3
rlabel polysilicon 30 -2017 30 -2017 0 1
rlabel polysilicon 30 -2023 30 -2023 0 3
rlabel polysilicon 44 -2017 44 -2017 0 1
rlabel polysilicon 44 -2023 44 -2023 0 3
rlabel polysilicon 51 -2017 51 -2017 0 1
rlabel polysilicon 51 -2023 51 -2023 0 3
rlabel polysilicon 58 -2017 58 -2017 0 1
rlabel polysilicon 58 -2023 58 -2023 0 3
rlabel polysilicon 65 -2017 65 -2017 0 1
rlabel polysilicon 68 -2017 68 -2017 0 2
rlabel polysilicon 65 -2023 65 -2023 0 3
rlabel polysilicon 72 -2017 72 -2017 0 1
rlabel polysilicon 72 -2023 72 -2023 0 3
rlabel polysilicon 79 -2017 79 -2017 0 1
rlabel polysilicon 79 -2023 79 -2023 0 3
rlabel polysilicon 86 -2017 86 -2017 0 1
rlabel polysilicon 89 -2017 89 -2017 0 2
rlabel polysilicon 86 -2023 86 -2023 0 3
rlabel polysilicon 93 -2017 93 -2017 0 1
rlabel polysilicon 93 -2023 93 -2023 0 3
rlabel polysilicon 100 -2017 100 -2017 0 1
rlabel polysilicon 103 -2017 103 -2017 0 2
rlabel polysilicon 100 -2023 100 -2023 0 3
rlabel polysilicon 103 -2023 103 -2023 0 4
rlabel polysilicon 107 -2017 107 -2017 0 1
rlabel polysilicon 110 -2017 110 -2017 0 2
rlabel polysilicon 107 -2023 107 -2023 0 3
rlabel polysilicon 114 -2017 114 -2017 0 1
rlabel polysilicon 114 -2023 114 -2023 0 3
rlabel polysilicon 121 -2017 121 -2017 0 1
rlabel polysilicon 124 -2017 124 -2017 0 2
rlabel polysilicon 121 -2023 121 -2023 0 3
rlabel polysilicon 124 -2023 124 -2023 0 4
rlabel polysilicon 131 -2017 131 -2017 0 2
rlabel polysilicon 128 -2023 128 -2023 0 3
rlabel polysilicon 131 -2023 131 -2023 0 4
rlabel polysilicon 135 -2017 135 -2017 0 1
rlabel polysilicon 135 -2023 135 -2023 0 3
rlabel polysilicon 142 -2017 142 -2017 0 1
rlabel polysilicon 145 -2017 145 -2017 0 2
rlabel polysilicon 142 -2023 142 -2023 0 3
rlabel polysilicon 145 -2023 145 -2023 0 4
rlabel polysilicon 149 -2017 149 -2017 0 1
rlabel polysilicon 152 -2017 152 -2017 0 2
rlabel polysilicon 152 -2023 152 -2023 0 4
rlabel polysilicon 156 -2017 156 -2017 0 1
rlabel polysilicon 156 -2023 156 -2023 0 3
rlabel polysilicon 163 -2017 163 -2017 0 1
rlabel polysilicon 163 -2023 163 -2023 0 3
rlabel polysilicon 170 -2017 170 -2017 0 1
rlabel polysilicon 170 -2023 170 -2023 0 3
rlabel polysilicon 177 -2017 177 -2017 0 1
rlabel polysilicon 180 -2017 180 -2017 0 2
rlabel polysilicon 177 -2023 177 -2023 0 3
rlabel polysilicon 180 -2023 180 -2023 0 4
rlabel polysilicon 184 -2017 184 -2017 0 1
rlabel polysilicon 184 -2023 184 -2023 0 3
rlabel polysilicon 191 -2017 191 -2017 0 1
rlabel polysilicon 191 -2023 191 -2023 0 3
rlabel polysilicon 198 -2017 198 -2017 0 1
rlabel polysilicon 198 -2023 198 -2023 0 3
rlabel polysilicon 205 -2017 205 -2017 0 1
rlabel polysilicon 205 -2023 205 -2023 0 3
rlabel polysilicon 212 -2017 212 -2017 0 1
rlabel polysilicon 215 -2017 215 -2017 0 2
rlabel polysilicon 212 -2023 212 -2023 0 3
rlabel polysilicon 219 -2017 219 -2017 0 1
rlabel polysilicon 219 -2023 219 -2023 0 3
rlabel polysilicon 222 -2023 222 -2023 0 4
rlabel polysilicon 226 -2017 226 -2017 0 1
rlabel polysilicon 226 -2023 226 -2023 0 3
rlabel polysilicon 233 -2017 233 -2017 0 1
rlabel polysilicon 233 -2023 233 -2023 0 3
rlabel polysilicon 240 -2017 240 -2017 0 1
rlabel polysilicon 240 -2023 240 -2023 0 3
rlabel polysilicon 247 -2017 247 -2017 0 1
rlabel polysilicon 247 -2023 247 -2023 0 3
rlabel polysilicon 254 -2017 254 -2017 0 1
rlabel polysilicon 254 -2023 254 -2023 0 3
rlabel polysilicon 261 -2017 261 -2017 0 1
rlabel polysilicon 261 -2023 261 -2023 0 3
rlabel polysilicon 268 -2017 268 -2017 0 1
rlabel polysilicon 268 -2023 268 -2023 0 3
rlabel polysilicon 275 -2017 275 -2017 0 1
rlabel polysilicon 275 -2023 275 -2023 0 3
rlabel polysilicon 282 -2017 282 -2017 0 1
rlabel polysilicon 282 -2023 282 -2023 0 3
rlabel polysilicon 289 -2017 289 -2017 0 1
rlabel polysilicon 289 -2023 289 -2023 0 3
rlabel polysilicon 296 -2017 296 -2017 0 1
rlabel polysilicon 296 -2023 296 -2023 0 3
rlabel polysilicon 303 -2017 303 -2017 0 1
rlabel polysilicon 303 -2023 303 -2023 0 3
rlabel polysilicon 310 -2017 310 -2017 0 1
rlabel polysilicon 310 -2023 310 -2023 0 3
rlabel polysilicon 317 -2017 317 -2017 0 1
rlabel polysilicon 317 -2023 317 -2023 0 3
rlabel polysilicon 324 -2017 324 -2017 0 1
rlabel polysilicon 324 -2023 324 -2023 0 3
rlabel polysilicon 331 -2017 331 -2017 0 1
rlabel polysilicon 334 -2017 334 -2017 0 2
rlabel polysilicon 331 -2023 331 -2023 0 3
rlabel polysilicon 338 -2017 338 -2017 0 1
rlabel polysilicon 338 -2023 338 -2023 0 3
rlabel polysilicon 345 -2017 345 -2017 0 1
rlabel polysilicon 345 -2023 345 -2023 0 3
rlabel polysilicon 352 -2017 352 -2017 0 1
rlabel polysilicon 352 -2023 352 -2023 0 3
rlabel polysilicon 359 -2017 359 -2017 0 1
rlabel polysilicon 359 -2023 359 -2023 0 3
rlabel polysilicon 366 -2017 366 -2017 0 1
rlabel polysilicon 366 -2023 366 -2023 0 3
rlabel polysilicon 373 -2017 373 -2017 0 1
rlabel polysilicon 373 -2023 373 -2023 0 3
rlabel polysilicon 380 -2017 380 -2017 0 1
rlabel polysilicon 380 -2023 380 -2023 0 3
rlabel polysilicon 387 -2023 387 -2023 0 3
rlabel polysilicon 394 -2017 394 -2017 0 1
rlabel polysilicon 394 -2023 394 -2023 0 3
rlabel polysilicon 401 -2017 401 -2017 0 1
rlabel polysilicon 401 -2023 401 -2023 0 3
rlabel polysilicon 408 -2017 408 -2017 0 1
rlabel polysilicon 408 -2023 408 -2023 0 3
rlabel polysilicon 415 -2017 415 -2017 0 1
rlabel polysilicon 415 -2023 415 -2023 0 3
rlabel polysilicon 422 -2017 422 -2017 0 1
rlabel polysilicon 422 -2023 422 -2023 0 3
rlabel polysilicon 429 -2017 429 -2017 0 1
rlabel polysilicon 429 -2023 429 -2023 0 3
rlabel polysilicon 436 -2017 436 -2017 0 1
rlabel polysilicon 436 -2023 436 -2023 0 3
rlabel polysilicon 443 -2017 443 -2017 0 1
rlabel polysilicon 443 -2023 443 -2023 0 3
rlabel polysilicon 450 -2017 450 -2017 0 1
rlabel polysilicon 450 -2023 450 -2023 0 3
rlabel polysilicon 457 -2017 457 -2017 0 1
rlabel polysilicon 460 -2017 460 -2017 0 2
rlabel polysilicon 457 -2023 457 -2023 0 3
rlabel polysilicon 460 -2023 460 -2023 0 4
rlabel polysilicon 464 -2017 464 -2017 0 1
rlabel polysilicon 464 -2023 464 -2023 0 3
rlabel polysilicon 471 -2017 471 -2017 0 1
rlabel polysilicon 471 -2023 471 -2023 0 3
rlabel polysilicon 478 -2017 478 -2017 0 1
rlabel polysilicon 478 -2023 478 -2023 0 3
rlabel polysilicon 485 -2023 485 -2023 0 3
rlabel polysilicon 492 -2017 492 -2017 0 1
rlabel polysilicon 492 -2023 492 -2023 0 3
rlabel polysilicon 499 -2017 499 -2017 0 1
rlabel polysilicon 499 -2023 499 -2023 0 3
rlabel polysilicon 506 -2017 506 -2017 0 1
rlabel polysilicon 509 -2017 509 -2017 0 2
rlabel polysilicon 509 -2023 509 -2023 0 4
rlabel polysilicon 513 -2017 513 -2017 0 1
rlabel polysilicon 513 -2023 513 -2023 0 3
rlabel polysilicon 520 -2017 520 -2017 0 1
rlabel polysilicon 520 -2023 520 -2023 0 3
rlabel polysilicon 527 -2017 527 -2017 0 1
rlabel polysilicon 527 -2023 527 -2023 0 3
rlabel polysilicon 534 -2017 534 -2017 0 1
rlabel polysilicon 541 -2017 541 -2017 0 1
rlabel polysilicon 541 -2023 541 -2023 0 3
rlabel polysilicon 548 -2017 548 -2017 0 1
rlabel polysilicon 548 -2023 548 -2023 0 3
rlabel polysilicon 555 -2017 555 -2017 0 1
rlabel polysilicon 555 -2023 555 -2023 0 3
rlabel polysilicon 562 -2017 562 -2017 0 1
rlabel polysilicon 562 -2023 562 -2023 0 3
rlabel polysilicon 569 -2017 569 -2017 0 1
rlabel polysilicon 569 -2023 569 -2023 0 3
rlabel polysilicon 572 -2023 572 -2023 0 4
rlabel polysilicon 576 -2017 576 -2017 0 1
rlabel polysilicon 576 -2023 576 -2023 0 3
rlabel polysilicon 583 -2017 583 -2017 0 1
rlabel polysilicon 583 -2023 583 -2023 0 3
rlabel polysilicon 593 -2017 593 -2017 0 2
rlabel polysilicon 593 -2023 593 -2023 0 4
rlabel polysilicon 597 -2017 597 -2017 0 1
rlabel polysilicon 597 -2023 597 -2023 0 3
rlabel polysilicon 604 -2017 604 -2017 0 1
rlabel polysilicon 604 -2023 604 -2023 0 3
rlabel polysilicon 611 -2017 611 -2017 0 1
rlabel polysilicon 611 -2023 611 -2023 0 3
rlabel polysilicon 618 -2017 618 -2017 0 1
rlabel polysilicon 618 -2023 618 -2023 0 3
rlabel polysilicon 625 -2017 625 -2017 0 1
rlabel polysilicon 628 -2017 628 -2017 0 2
rlabel polysilicon 625 -2023 625 -2023 0 3
rlabel polysilicon 628 -2023 628 -2023 0 4
rlabel polysilicon 632 -2017 632 -2017 0 1
rlabel polysilicon 632 -2023 632 -2023 0 3
rlabel polysilicon 639 -2017 639 -2017 0 1
rlabel polysilicon 639 -2023 639 -2023 0 3
rlabel polysilicon 646 -2017 646 -2017 0 1
rlabel polysilicon 646 -2023 646 -2023 0 3
rlabel polysilicon 653 -2017 653 -2017 0 1
rlabel polysilicon 653 -2023 653 -2023 0 3
rlabel polysilicon 660 -2017 660 -2017 0 1
rlabel polysilicon 660 -2023 660 -2023 0 3
rlabel polysilicon 667 -2017 667 -2017 0 1
rlabel polysilicon 667 -2023 667 -2023 0 3
rlabel polysilicon 674 -2017 674 -2017 0 1
rlabel polysilicon 674 -2023 674 -2023 0 3
rlabel polysilicon 681 -2017 681 -2017 0 1
rlabel polysilicon 681 -2023 681 -2023 0 3
rlabel polysilicon 688 -2017 688 -2017 0 1
rlabel polysilicon 688 -2023 688 -2023 0 3
rlabel polysilicon 695 -2017 695 -2017 0 1
rlabel polysilicon 695 -2023 695 -2023 0 3
rlabel polysilicon 702 -2017 702 -2017 0 1
rlabel polysilicon 702 -2023 702 -2023 0 3
rlabel polysilicon 709 -2017 709 -2017 0 1
rlabel polysilicon 709 -2023 709 -2023 0 3
rlabel polysilicon 716 -2017 716 -2017 0 1
rlabel polysilicon 719 -2017 719 -2017 0 2
rlabel polysilicon 716 -2023 716 -2023 0 3
rlabel polysilicon 719 -2023 719 -2023 0 4
rlabel polysilicon 723 -2017 723 -2017 0 1
rlabel polysilicon 723 -2023 723 -2023 0 3
rlabel polysilicon 730 -2017 730 -2017 0 1
rlabel polysilicon 730 -2023 730 -2023 0 3
rlabel polysilicon 737 -2017 737 -2017 0 1
rlabel polysilicon 737 -2023 737 -2023 0 3
rlabel polysilicon 744 -2017 744 -2017 0 1
rlabel polysilicon 744 -2023 744 -2023 0 3
rlabel polysilicon 751 -2017 751 -2017 0 1
rlabel polysilicon 751 -2023 751 -2023 0 3
rlabel polysilicon 758 -2017 758 -2017 0 1
rlabel polysilicon 761 -2017 761 -2017 0 2
rlabel polysilicon 758 -2023 758 -2023 0 3
rlabel polysilicon 761 -2023 761 -2023 0 4
rlabel polysilicon 765 -2017 765 -2017 0 1
rlabel polysilicon 765 -2023 765 -2023 0 3
rlabel polysilicon 772 -2017 772 -2017 0 1
rlabel polysilicon 772 -2023 772 -2023 0 3
rlabel polysilicon 779 -2017 779 -2017 0 1
rlabel polysilicon 779 -2023 779 -2023 0 3
rlabel polysilicon 786 -2017 786 -2017 0 1
rlabel polysilicon 786 -2023 786 -2023 0 3
rlabel polysilicon 793 -2017 793 -2017 0 1
rlabel polysilicon 796 -2017 796 -2017 0 2
rlabel polysilicon 796 -2023 796 -2023 0 4
rlabel polysilicon 800 -2017 800 -2017 0 1
rlabel polysilicon 800 -2023 800 -2023 0 3
rlabel polysilicon 807 -2017 807 -2017 0 1
rlabel polysilicon 807 -2023 807 -2023 0 3
rlabel polysilicon 814 -2017 814 -2017 0 1
rlabel polysilicon 814 -2023 814 -2023 0 3
rlabel polysilicon 821 -2017 821 -2017 0 1
rlabel polysilicon 821 -2023 821 -2023 0 3
rlabel polysilicon 828 -2017 828 -2017 0 1
rlabel polysilicon 828 -2023 828 -2023 0 3
rlabel polysilicon 835 -2017 835 -2017 0 1
rlabel polysilicon 835 -2023 835 -2023 0 3
rlabel polysilicon 842 -2017 842 -2017 0 1
rlabel polysilicon 842 -2023 842 -2023 0 3
rlabel polysilicon 849 -2017 849 -2017 0 1
rlabel polysilicon 849 -2023 849 -2023 0 3
rlabel polysilicon 856 -2017 856 -2017 0 1
rlabel polysilicon 856 -2023 856 -2023 0 3
rlabel polysilicon 863 -2017 863 -2017 0 1
rlabel polysilicon 863 -2023 863 -2023 0 3
rlabel polysilicon 870 -2017 870 -2017 0 1
rlabel polysilicon 870 -2023 870 -2023 0 3
rlabel polysilicon 877 -2017 877 -2017 0 1
rlabel polysilicon 877 -2023 877 -2023 0 3
rlabel polysilicon 884 -2017 884 -2017 0 1
rlabel polysilicon 887 -2017 887 -2017 0 2
rlabel polysilicon 884 -2023 884 -2023 0 3
rlabel polysilicon 887 -2023 887 -2023 0 4
rlabel polysilicon 891 -2017 891 -2017 0 1
rlabel polysilicon 894 -2017 894 -2017 0 2
rlabel polysilicon 891 -2023 891 -2023 0 3
rlabel polysilicon 894 -2023 894 -2023 0 4
rlabel polysilicon 898 -2017 898 -2017 0 1
rlabel polysilicon 901 -2017 901 -2017 0 2
rlabel polysilicon 901 -2023 901 -2023 0 4
rlabel polysilicon 905 -2017 905 -2017 0 1
rlabel polysilicon 905 -2023 905 -2023 0 3
rlabel polysilicon 912 -2017 912 -2017 0 1
rlabel polysilicon 912 -2023 912 -2023 0 3
rlabel polysilicon 919 -2017 919 -2017 0 1
rlabel polysilicon 922 -2017 922 -2017 0 2
rlabel polysilicon 919 -2023 919 -2023 0 3
rlabel polysilicon 922 -2023 922 -2023 0 4
rlabel polysilicon 926 -2017 926 -2017 0 1
rlabel polysilicon 926 -2023 926 -2023 0 3
rlabel polysilicon 933 -2017 933 -2017 0 1
rlabel polysilicon 933 -2023 933 -2023 0 3
rlabel polysilicon 940 -2017 940 -2017 0 1
rlabel polysilicon 940 -2023 940 -2023 0 3
rlabel polysilicon 947 -2017 947 -2017 0 1
rlabel polysilicon 947 -2023 947 -2023 0 3
rlabel polysilicon 954 -2017 954 -2017 0 1
rlabel polysilicon 954 -2023 954 -2023 0 3
rlabel polysilicon 957 -2023 957 -2023 0 4
rlabel polysilicon 961 -2017 961 -2017 0 1
rlabel polysilicon 964 -2023 964 -2023 0 4
rlabel polysilicon 968 -2017 968 -2017 0 1
rlabel polysilicon 968 -2023 968 -2023 0 3
rlabel polysilicon 975 -2017 975 -2017 0 1
rlabel polysilicon 975 -2023 975 -2023 0 3
rlabel polysilicon 982 -2017 982 -2017 0 1
rlabel polysilicon 982 -2023 982 -2023 0 3
rlabel polysilicon 989 -2017 989 -2017 0 1
rlabel polysilicon 989 -2023 989 -2023 0 3
rlabel polysilicon 992 -2023 992 -2023 0 4
rlabel polysilicon 999 -2017 999 -2017 0 2
rlabel polysilicon 996 -2023 996 -2023 0 3
rlabel polysilicon 999 -2023 999 -2023 0 4
rlabel polysilicon 1003 -2017 1003 -2017 0 1
rlabel polysilicon 1003 -2023 1003 -2023 0 3
rlabel polysilicon 1010 -2017 1010 -2017 0 1
rlabel polysilicon 1010 -2023 1010 -2023 0 3
rlabel polysilicon 1017 -2017 1017 -2017 0 1
rlabel polysilicon 1017 -2023 1017 -2023 0 3
rlabel polysilicon 1024 -2017 1024 -2017 0 1
rlabel polysilicon 1024 -2023 1024 -2023 0 3
rlabel polysilicon 1031 -2017 1031 -2017 0 1
rlabel polysilicon 1031 -2023 1031 -2023 0 3
rlabel polysilicon 1038 -2017 1038 -2017 0 1
rlabel polysilicon 1041 -2017 1041 -2017 0 2
rlabel polysilicon 1045 -2017 1045 -2017 0 1
rlabel polysilicon 1045 -2023 1045 -2023 0 3
rlabel polysilicon 1052 -2017 1052 -2017 0 1
rlabel polysilicon 1052 -2023 1052 -2023 0 3
rlabel polysilicon 1059 -2017 1059 -2017 0 1
rlabel polysilicon 1059 -2023 1059 -2023 0 3
rlabel polysilicon 1066 -2017 1066 -2017 0 1
rlabel polysilicon 1066 -2023 1066 -2023 0 3
rlabel polysilicon 1073 -2017 1073 -2017 0 1
rlabel polysilicon 1073 -2023 1073 -2023 0 3
rlabel polysilicon 1080 -2017 1080 -2017 0 1
rlabel polysilicon 1080 -2023 1080 -2023 0 3
rlabel polysilicon 1087 -2017 1087 -2017 0 1
rlabel polysilicon 1087 -2023 1087 -2023 0 3
rlabel polysilicon 1094 -2017 1094 -2017 0 1
rlabel polysilicon 1094 -2023 1094 -2023 0 3
rlabel polysilicon 1101 -2017 1101 -2017 0 1
rlabel polysilicon 1101 -2023 1101 -2023 0 3
rlabel polysilicon 1108 -2017 1108 -2017 0 1
rlabel polysilicon 1111 -2017 1111 -2017 0 2
rlabel polysilicon 1108 -2023 1108 -2023 0 3
rlabel polysilicon 1115 -2017 1115 -2017 0 1
rlabel polysilicon 1115 -2023 1115 -2023 0 3
rlabel polysilicon 1122 -2017 1122 -2017 0 1
rlabel polysilicon 1122 -2023 1122 -2023 0 3
rlabel polysilicon 1129 -2017 1129 -2017 0 1
rlabel polysilicon 1129 -2023 1129 -2023 0 3
rlabel polysilicon 1136 -2017 1136 -2017 0 1
rlabel polysilicon 1139 -2017 1139 -2017 0 2
rlabel polysilicon 1139 -2023 1139 -2023 0 4
rlabel polysilicon 1143 -2017 1143 -2017 0 1
rlabel polysilicon 1143 -2023 1143 -2023 0 3
rlabel polysilicon 1150 -2017 1150 -2017 0 1
rlabel polysilicon 1150 -2023 1150 -2023 0 3
rlabel polysilicon 1157 -2017 1157 -2017 0 1
rlabel polysilicon 1157 -2023 1157 -2023 0 3
rlabel polysilicon 1164 -2017 1164 -2017 0 1
rlabel polysilicon 1164 -2023 1164 -2023 0 3
rlabel polysilicon 1171 -2017 1171 -2017 0 1
rlabel polysilicon 1171 -2023 1171 -2023 0 3
rlabel polysilicon 1178 -2017 1178 -2017 0 1
rlabel polysilicon 1178 -2023 1178 -2023 0 3
rlabel polysilicon 1185 -2017 1185 -2017 0 1
rlabel polysilicon 1185 -2023 1185 -2023 0 3
rlabel polysilicon 1192 -2017 1192 -2017 0 1
rlabel polysilicon 1195 -2023 1195 -2023 0 4
rlabel polysilicon 1199 -2017 1199 -2017 0 1
rlabel polysilicon 1199 -2023 1199 -2023 0 3
rlabel polysilicon 1206 -2017 1206 -2017 0 1
rlabel polysilicon 1206 -2023 1206 -2023 0 3
rlabel polysilicon 1216 -2017 1216 -2017 0 2
rlabel polysilicon 1213 -2023 1213 -2023 0 3
rlabel polysilicon 1220 -2017 1220 -2017 0 1
rlabel polysilicon 1220 -2023 1220 -2023 0 3
rlabel polysilicon 1227 -2017 1227 -2017 0 1
rlabel polysilicon 1227 -2023 1227 -2023 0 3
rlabel polysilicon 1234 -2017 1234 -2017 0 1
rlabel polysilicon 1234 -2023 1234 -2023 0 3
rlabel polysilicon 1241 -2017 1241 -2017 0 1
rlabel polysilicon 1241 -2023 1241 -2023 0 3
rlabel polysilicon 1248 -2017 1248 -2017 0 1
rlabel polysilicon 1248 -2023 1248 -2023 0 3
rlabel polysilicon 1255 -2017 1255 -2017 0 1
rlabel polysilicon 1255 -2023 1255 -2023 0 3
rlabel polysilicon 1262 -2017 1262 -2017 0 1
rlabel polysilicon 1262 -2023 1262 -2023 0 3
rlabel polysilicon 1269 -2017 1269 -2017 0 1
rlabel polysilicon 1269 -2023 1269 -2023 0 3
rlabel polysilicon 1276 -2017 1276 -2017 0 1
rlabel polysilicon 1276 -2023 1276 -2023 0 3
rlabel polysilicon 1283 -2017 1283 -2017 0 1
rlabel polysilicon 1283 -2023 1283 -2023 0 3
rlabel polysilicon 1293 -2017 1293 -2017 0 2
rlabel polysilicon 1290 -2023 1290 -2023 0 3
rlabel polysilicon 1293 -2023 1293 -2023 0 4
rlabel polysilicon 1297 -2017 1297 -2017 0 1
rlabel polysilicon 1297 -2023 1297 -2023 0 3
rlabel polysilicon 1304 -2017 1304 -2017 0 1
rlabel polysilicon 1304 -2023 1304 -2023 0 3
rlabel polysilicon 1311 -2017 1311 -2017 0 1
rlabel polysilicon 1311 -2023 1311 -2023 0 3
rlabel polysilicon 1318 -2017 1318 -2017 0 1
rlabel polysilicon 1318 -2023 1318 -2023 0 3
rlabel polysilicon 1325 -2017 1325 -2017 0 1
rlabel polysilicon 1325 -2023 1325 -2023 0 3
rlabel polysilicon 1332 -2017 1332 -2017 0 1
rlabel polysilicon 1332 -2023 1332 -2023 0 3
rlabel polysilicon 1339 -2017 1339 -2017 0 1
rlabel polysilicon 1339 -2023 1339 -2023 0 3
rlabel polysilicon 1346 -2017 1346 -2017 0 1
rlabel polysilicon 1346 -2023 1346 -2023 0 3
rlabel polysilicon 1353 -2017 1353 -2017 0 1
rlabel polysilicon 1353 -2023 1353 -2023 0 3
rlabel polysilicon 1360 -2017 1360 -2017 0 1
rlabel polysilicon 1360 -2023 1360 -2023 0 3
rlabel polysilicon 1367 -2017 1367 -2017 0 1
rlabel polysilicon 1367 -2023 1367 -2023 0 3
rlabel polysilicon 1374 -2017 1374 -2017 0 1
rlabel polysilicon 1374 -2023 1374 -2023 0 3
rlabel polysilicon 1381 -2017 1381 -2017 0 1
rlabel polysilicon 1384 -2017 1384 -2017 0 2
rlabel polysilicon 1381 -2023 1381 -2023 0 3
rlabel polysilicon 1388 -2017 1388 -2017 0 1
rlabel polysilicon 1388 -2023 1388 -2023 0 3
rlabel polysilicon 1395 -2017 1395 -2017 0 1
rlabel polysilicon 1395 -2023 1395 -2023 0 3
rlabel polysilicon 1402 -2017 1402 -2017 0 1
rlabel polysilicon 1402 -2023 1402 -2023 0 3
rlabel polysilicon 1409 -2017 1409 -2017 0 1
rlabel polysilicon 1409 -2023 1409 -2023 0 3
rlabel polysilicon 1416 -2017 1416 -2017 0 1
rlabel polysilicon 1416 -2023 1416 -2023 0 3
rlabel polysilicon 1423 -2017 1423 -2017 0 1
rlabel polysilicon 1423 -2023 1423 -2023 0 3
rlabel polysilicon 1430 -2017 1430 -2017 0 1
rlabel polysilicon 1430 -2023 1430 -2023 0 3
rlabel polysilicon 1437 -2017 1437 -2017 0 1
rlabel polysilicon 1437 -2023 1437 -2023 0 3
rlabel polysilicon 1444 -2017 1444 -2017 0 1
rlabel polysilicon 1444 -2023 1444 -2023 0 3
rlabel polysilicon 1451 -2017 1451 -2017 0 1
rlabel polysilicon 1451 -2023 1451 -2023 0 3
rlabel polysilicon 1458 -2017 1458 -2017 0 1
rlabel polysilicon 1458 -2023 1458 -2023 0 3
rlabel polysilicon 1465 -2017 1465 -2017 0 1
rlabel polysilicon 1465 -2023 1465 -2023 0 3
rlabel polysilicon 1472 -2017 1472 -2017 0 1
rlabel polysilicon 1472 -2023 1472 -2023 0 3
rlabel polysilicon 1479 -2017 1479 -2017 0 1
rlabel polysilicon 1479 -2023 1479 -2023 0 3
rlabel polysilicon 1486 -2017 1486 -2017 0 1
rlabel polysilicon 1486 -2023 1486 -2023 0 3
rlabel polysilicon 1493 -2017 1493 -2017 0 1
rlabel polysilicon 1493 -2023 1493 -2023 0 3
rlabel polysilicon 1500 -2017 1500 -2017 0 1
rlabel polysilicon 1500 -2023 1500 -2023 0 3
rlabel polysilicon 1507 -2017 1507 -2017 0 1
rlabel polysilicon 1507 -2023 1507 -2023 0 3
rlabel polysilicon 1514 -2017 1514 -2017 0 1
rlabel polysilicon 1514 -2023 1514 -2023 0 3
rlabel polysilicon 1521 -2017 1521 -2017 0 1
rlabel polysilicon 1521 -2023 1521 -2023 0 3
rlabel polysilicon 1528 -2017 1528 -2017 0 1
rlabel polysilicon 1528 -2023 1528 -2023 0 3
rlabel polysilicon 1535 -2017 1535 -2017 0 1
rlabel polysilicon 1535 -2023 1535 -2023 0 3
rlabel polysilicon 1542 -2017 1542 -2017 0 1
rlabel polysilicon 1542 -2023 1542 -2023 0 3
rlabel polysilicon 1549 -2017 1549 -2017 0 1
rlabel polysilicon 1549 -2023 1549 -2023 0 3
rlabel polysilicon 1556 -2017 1556 -2017 0 1
rlabel polysilicon 1556 -2023 1556 -2023 0 3
rlabel polysilicon 1563 -2017 1563 -2017 0 1
rlabel polysilicon 1563 -2023 1563 -2023 0 3
rlabel polysilicon 1570 -2017 1570 -2017 0 1
rlabel polysilicon 1570 -2023 1570 -2023 0 3
rlabel polysilicon 1577 -2017 1577 -2017 0 1
rlabel polysilicon 1577 -2023 1577 -2023 0 3
rlabel polysilicon 1584 -2017 1584 -2017 0 1
rlabel polysilicon 1584 -2023 1584 -2023 0 3
rlabel polysilicon 1591 -2017 1591 -2017 0 1
rlabel polysilicon 1591 -2023 1591 -2023 0 3
rlabel polysilicon 1594 -2023 1594 -2023 0 4
rlabel polysilicon 1598 -2017 1598 -2017 0 1
rlabel polysilicon 1598 -2023 1598 -2023 0 3
rlabel polysilicon 1605 -2017 1605 -2017 0 1
rlabel polysilicon 1605 -2023 1605 -2023 0 3
rlabel polysilicon 1612 -2017 1612 -2017 0 1
rlabel polysilicon 1612 -2023 1612 -2023 0 3
rlabel polysilicon 1619 -2017 1619 -2017 0 1
rlabel polysilicon 1619 -2023 1619 -2023 0 3
rlabel polysilicon 1626 -2017 1626 -2017 0 1
rlabel polysilicon 1626 -2023 1626 -2023 0 3
rlabel polysilicon 1633 -2017 1633 -2017 0 1
rlabel polysilicon 1633 -2023 1633 -2023 0 3
rlabel polysilicon 1640 -2017 1640 -2017 0 1
rlabel polysilicon 1640 -2023 1640 -2023 0 3
rlabel polysilicon 1647 -2017 1647 -2017 0 1
rlabel polysilicon 1647 -2023 1647 -2023 0 3
rlabel polysilicon 1654 -2017 1654 -2017 0 1
rlabel polysilicon 1654 -2023 1654 -2023 0 3
rlabel polysilicon 1661 -2017 1661 -2017 0 1
rlabel polysilicon 1661 -2023 1661 -2023 0 3
rlabel polysilicon 1668 -2017 1668 -2017 0 1
rlabel polysilicon 1668 -2023 1668 -2023 0 3
rlabel polysilicon 1675 -2017 1675 -2017 0 1
rlabel polysilicon 1675 -2023 1675 -2023 0 3
rlabel polysilicon 1682 -2017 1682 -2017 0 1
rlabel polysilicon 1682 -2023 1682 -2023 0 3
rlabel polysilicon 1689 -2017 1689 -2017 0 1
rlabel polysilicon 1689 -2023 1689 -2023 0 3
rlabel polysilicon 1696 -2017 1696 -2017 0 1
rlabel polysilicon 1696 -2023 1696 -2023 0 3
rlabel polysilicon 1703 -2017 1703 -2017 0 1
rlabel polysilicon 1703 -2023 1703 -2023 0 3
rlabel polysilicon 1710 -2017 1710 -2017 0 1
rlabel polysilicon 1710 -2023 1710 -2023 0 3
rlabel polysilicon 1717 -2017 1717 -2017 0 1
rlabel polysilicon 1717 -2023 1717 -2023 0 3
rlabel polysilicon 1724 -2017 1724 -2017 0 1
rlabel polysilicon 1724 -2023 1724 -2023 0 3
rlabel polysilicon 1731 -2017 1731 -2017 0 1
rlabel polysilicon 1731 -2023 1731 -2023 0 3
rlabel polysilicon 1738 -2017 1738 -2017 0 1
rlabel polysilicon 1738 -2023 1738 -2023 0 3
rlabel polysilicon 1745 -2023 1745 -2023 0 3
rlabel polysilicon 1748 -2023 1748 -2023 0 4
rlabel polysilicon 1752 -2017 1752 -2017 0 1
rlabel polysilicon 1752 -2023 1752 -2023 0 3
rlabel polysilicon 1759 -2017 1759 -2017 0 1
rlabel polysilicon 1759 -2023 1759 -2023 0 3
rlabel polysilicon 1766 -2017 1766 -2017 0 1
rlabel polysilicon 1766 -2023 1766 -2023 0 3
rlabel polysilicon 1773 -2017 1773 -2017 0 1
rlabel polysilicon 1773 -2023 1773 -2023 0 3
rlabel polysilicon 1780 -2017 1780 -2017 0 1
rlabel polysilicon 1780 -2023 1780 -2023 0 3
rlabel polysilicon 1787 -2017 1787 -2017 0 1
rlabel polysilicon 1787 -2023 1787 -2023 0 3
rlabel polysilicon 1794 -2017 1794 -2017 0 1
rlabel polysilicon 1794 -2023 1794 -2023 0 3
rlabel polysilicon 1801 -2017 1801 -2017 0 1
rlabel polysilicon 1801 -2023 1801 -2023 0 3
rlabel polysilicon 1808 -2017 1808 -2017 0 1
rlabel polysilicon 1808 -2023 1808 -2023 0 3
rlabel polysilicon 30 -2172 30 -2172 0 1
rlabel polysilicon 30 -2178 30 -2178 0 3
rlabel polysilicon 37 -2172 37 -2172 0 1
rlabel polysilicon 37 -2178 37 -2178 0 3
rlabel polysilicon 44 -2172 44 -2172 0 1
rlabel polysilicon 44 -2178 44 -2178 0 3
rlabel polysilicon 51 -2172 51 -2172 0 1
rlabel polysilicon 51 -2178 51 -2178 0 3
rlabel polysilicon 61 -2172 61 -2172 0 2
rlabel polysilicon 61 -2178 61 -2178 0 4
rlabel polysilicon 65 -2172 65 -2172 0 1
rlabel polysilicon 65 -2178 65 -2178 0 3
rlabel polysilicon 72 -2172 72 -2172 0 1
rlabel polysilicon 72 -2178 72 -2178 0 3
rlabel polysilicon 79 -2172 79 -2172 0 1
rlabel polysilicon 79 -2178 79 -2178 0 3
rlabel polysilicon 86 -2172 86 -2172 0 1
rlabel polysilicon 86 -2178 86 -2178 0 3
rlabel polysilicon 93 -2172 93 -2172 0 1
rlabel polysilicon 96 -2172 96 -2172 0 2
rlabel polysilicon 93 -2178 93 -2178 0 3
rlabel polysilicon 96 -2178 96 -2178 0 4
rlabel polysilicon 103 -2172 103 -2172 0 2
rlabel polysilicon 100 -2178 100 -2178 0 3
rlabel polysilicon 103 -2178 103 -2178 0 4
rlabel polysilicon 107 -2172 107 -2172 0 1
rlabel polysilicon 110 -2172 110 -2172 0 2
rlabel polysilicon 110 -2178 110 -2178 0 4
rlabel polysilicon 114 -2172 114 -2172 0 1
rlabel polysilicon 114 -2178 114 -2178 0 3
rlabel polysilicon 121 -2172 121 -2172 0 1
rlabel polysilicon 124 -2172 124 -2172 0 2
rlabel polysilicon 124 -2178 124 -2178 0 4
rlabel polysilicon 128 -2172 128 -2172 0 1
rlabel polysilicon 131 -2172 131 -2172 0 2
rlabel polysilicon 128 -2178 128 -2178 0 3
rlabel polysilicon 131 -2178 131 -2178 0 4
rlabel polysilicon 135 -2172 135 -2172 0 1
rlabel polysilicon 135 -2178 135 -2178 0 3
rlabel polysilicon 142 -2172 142 -2172 0 1
rlabel polysilicon 142 -2178 142 -2178 0 3
rlabel polysilicon 149 -2172 149 -2172 0 1
rlabel polysilicon 149 -2178 149 -2178 0 3
rlabel polysilicon 156 -2172 156 -2172 0 1
rlabel polysilicon 156 -2178 156 -2178 0 3
rlabel polysilicon 163 -2172 163 -2172 0 1
rlabel polysilicon 163 -2178 163 -2178 0 3
rlabel polysilicon 170 -2172 170 -2172 0 1
rlabel polysilicon 170 -2178 170 -2178 0 3
rlabel polysilicon 177 -2172 177 -2172 0 1
rlabel polysilicon 177 -2178 177 -2178 0 3
rlabel polysilicon 184 -2172 184 -2172 0 1
rlabel polysilicon 184 -2178 184 -2178 0 3
rlabel polysilicon 191 -2172 191 -2172 0 1
rlabel polysilicon 191 -2178 191 -2178 0 3
rlabel polysilicon 198 -2172 198 -2172 0 1
rlabel polysilicon 201 -2172 201 -2172 0 2
rlabel polysilicon 201 -2178 201 -2178 0 4
rlabel polysilicon 205 -2172 205 -2172 0 1
rlabel polysilicon 205 -2178 205 -2178 0 3
rlabel polysilicon 212 -2172 212 -2172 0 1
rlabel polysilicon 212 -2178 212 -2178 0 3
rlabel polysilicon 219 -2172 219 -2172 0 1
rlabel polysilicon 219 -2178 219 -2178 0 3
rlabel polysilicon 226 -2172 226 -2172 0 1
rlabel polysilicon 229 -2172 229 -2172 0 2
rlabel polysilicon 226 -2178 226 -2178 0 3
rlabel polysilicon 229 -2178 229 -2178 0 4
rlabel polysilicon 233 -2172 233 -2172 0 1
rlabel polysilicon 233 -2178 233 -2178 0 3
rlabel polysilicon 240 -2172 240 -2172 0 1
rlabel polysilicon 240 -2178 240 -2178 0 3
rlabel polysilicon 247 -2172 247 -2172 0 1
rlabel polysilicon 250 -2172 250 -2172 0 2
rlabel polysilicon 250 -2178 250 -2178 0 4
rlabel polysilicon 254 -2172 254 -2172 0 1
rlabel polysilicon 257 -2178 257 -2178 0 4
rlabel polysilicon 261 -2172 261 -2172 0 1
rlabel polysilicon 261 -2178 261 -2178 0 3
rlabel polysilicon 268 -2172 268 -2172 0 1
rlabel polysilicon 268 -2178 268 -2178 0 3
rlabel polysilicon 275 -2172 275 -2172 0 1
rlabel polysilicon 278 -2172 278 -2172 0 2
rlabel polysilicon 282 -2172 282 -2172 0 1
rlabel polysilicon 282 -2178 282 -2178 0 3
rlabel polysilicon 289 -2172 289 -2172 0 1
rlabel polysilicon 292 -2172 292 -2172 0 2
rlabel polysilicon 296 -2172 296 -2172 0 1
rlabel polysilicon 296 -2178 296 -2178 0 3
rlabel polysilicon 303 -2172 303 -2172 0 1
rlabel polysilicon 303 -2178 303 -2178 0 3
rlabel polysilicon 310 -2172 310 -2172 0 1
rlabel polysilicon 310 -2178 310 -2178 0 3
rlabel polysilicon 317 -2172 317 -2172 0 1
rlabel polysilicon 317 -2178 317 -2178 0 3
rlabel polysilicon 324 -2172 324 -2172 0 1
rlabel polysilicon 324 -2178 324 -2178 0 3
rlabel polysilicon 331 -2172 331 -2172 0 1
rlabel polysilicon 331 -2178 331 -2178 0 3
rlabel polysilicon 338 -2172 338 -2172 0 1
rlabel polysilicon 338 -2178 338 -2178 0 3
rlabel polysilicon 345 -2172 345 -2172 0 1
rlabel polysilicon 345 -2178 345 -2178 0 3
rlabel polysilicon 352 -2172 352 -2172 0 1
rlabel polysilicon 352 -2178 352 -2178 0 3
rlabel polysilicon 359 -2172 359 -2172 0 1
rlabel polysilicon 359 -2178 359 -2178 0 3
rlabel polysilicon 366 -2172 366 -2172 0 1
rlabel polysilicon 366 -2178 366 -2178 0 3
rlabel polysilicon 373 -2172 373 -2172 0 1
rlabel polysilicon 376 -2178 376 -2178 0 4
rlabel polysilicon 380 -2172 380 -2172 0 1
rlabel polysilicon 380 -2178 380 -2178 0 3
rlabel polysilicon 387 -2172 387 -2172 0 1
rlabel polysilicon 387 -2178 387 -2178 0 3
rlabel polysilicon 394 -2172 394 -2172 0 1
rlabel polysilicon 394 -2178 394 -2178 0 3
rlabel polysilicon 401 -2172 401 -2172 0 1
rlabel polysilicon 401 -2178 401 -2178 0 3
rlabel polysilicon 408 -2172 408 -2172 0 1
rlabel polysilicon 408 -2178 408 -2178 0 3
rlabel polysilicon 418 -2172 418 -2172 0 2
rlabel polysilicon 415 -2178 415 -2178 0 3
rlabel polysilicon 418 -2178 418 -2178 0 4
rlabel polysilicon 422 -2172 422 -2172 0 1
rlabel polysilicon 422 -2178 422 -2178 0 3
rlabel polysilicon 429 -2172 429 -2172 0 1
rlabel polysilicon 436 -2172 436 -2172 0 1
rlabel polysilicon 436 -2178 436 -2178 0 3
rlabel polysilicon 443 -2172 443 -2172 0 1
rlabel polysilicon 443 -2178 443 -2178 0 3
rlabel polysilicon 450 -2172 450 -2172 0 1
rlabel polysilicon 450 -2178 450 -2178 0 3
rlabel polysilicon 457 -2172 457 -2172 0 1
rlabel polysilicon 457 -2178 457 -2178 0 3
rlabel polysilicon 464 -2172 464 -2172 0 1
rlabel polysilicon 464 -2178 464 -2178 0 3
rlabel polysilicon 471 -2172 471 -2172 0 1
rlabel polysilicon 471 -2178 471 -2178 0 3
rlabel polysilicon 478 -2172 478 -2172 0 1
rlabel polysilicon 478 -2178 478 -2178 0 3
rlabel polysilicon 485 -2172 485 -2172 0 1
rlabel polysilicon 485 -2178 485 -2178 0 3
rlabel polysilicon 492 -2172 492 -2172 0 1
rlabel polysilicon 492 -2178 492 -2178 0 3
rlabel polysilicon 499 -2172 499 -2172 0 1
rlabel polysilicon 499 -2178 499 -2178 0 3
rlabel polysilicon 506 -2172 506 -2172 0 1
rlabel polysilicon 506 -2178 506 -2178 0 3
rlabel polysilicon 513 -2172 513 -2172 0 1
rlabel polysilicon 516 -2172 516 -2172 0 2
rlabel polysilicon 513 -2178 513 -2178 0 3
rlabel polysilicon 516 -2178 516 -2178 0 4
rlabel polysilicon 520 -2172 520 -2172 0 1
rlabel polysilicon 520 -2178 520 -2178 0 3
rlabel polysilicon 527 -2172 527 -2172 0 1
rlabel polysilicon 527 -2178 527 -2178 0 3
rlabel polysilicon 534 -2178 534 -2178 0 3
rlabel polysilicon 541 -2172 541 -2172 0 1
rlabel polysilicon 541 -2178 541 -2178 0 3
rlabel polysilicon 548 -2172 548 -2172 0 1
rlabel polysilicon 548 -2178 548 -2178 0 3
rlabel polysilicon 555 -2172 555 -2172 0 1
rlabel polysilicon 558 -2172 558 -2172 0 2
rlabel polysilicon 555 -2178 555 -2178 0 3
rlabel polysilicon 558 -2178 558 -2178 0 4
rlabel polysilicon 562 -2172 562 -2172 0 1
rlabel polysilicon 562 -2178 562 -2178 0 3
rlabel polysilicon 569 -2172 569 -2172 0 1
rlabel polysilicon 569 -2178 569 -2178 0 3
rlabel polysilicon 576 -2172 576 -2172 0 1
rlabel polysilicon 576 -2178 576 -2178 0 3
rlabel polysilicon 583 -2172 583 -2172 0 1
rlabel polysilicon 586 -2172 586 -2172 0 2
rlabel polysilicon 583 -2178 583 -2178 0 3
rlabel polysilicon 586 -2178 586 -2178 0 4
rlabel polysilicon 590 -2172 590 -2172 0 1
rlabel polysilicon 590 -2178 590 -2178 0 3
rlabel polysilicon 597 -2172 597 -2172 0 1
rlabel polysilicon 597 -2178 597 -2178 0 3
rlabel polysilicon 604 -2172 604 -2172 0 1
rlabel polysilicon 604 -2178 604 -2178 0 3
rlabel polysilicon 611 -2172 611 -2172 0 1
rlabel polysilicon 614 -2172 614 -2172 0 2
rlabel polysilicon 614 -2178 614 -2178 0 4
rlabel polysilicon 618 -2172 618 -2172 0 1
rlabel polysilicon 618 -2178 618 -2178 0 3
rlabel polysilicon 625 -2172 625 -2172 0 1
rlabel polysilicon 628 -2172 628 -2172 0 2
rlabel polysilicon 625 -2178 625 -2178 0 3
rlabel polysilicon 628 -2178 628 -2178 0 4
rlabel polysilicon 632 -2172 632 -2172 0 1
rlabel polysilicon 632 -2178 632 -2178 0 3
rlabel polysilicon 639 -2172 639 -2172 0 1
rlabel polysilicon 639 -2178 639 -2178 0 3
rlabel polysilicon 646 -2172 646 -2172 0 1
rlabel polysilicon 646 -2178 646 -2178 0 3
rlabel polysilicon 653 -2172 653 -2172 0 1
rlabel polysilicon 653 -2178 653 -2178 0 3
rlabel polysilicon 660 -2172 660 -2172 0 1
rlabel polysilicon 660 -2178 660 -2178 0 3
rlabel polysilicon 667 -2172 667 -2172 0 1
rlabel polysilicon 667 -2178 667 -2178 0 3
rlabel polysilicon 674 -2172 674 -2172 0 1
rlabel polysilicon 674 -2178 674 -2178 0 3
rlabel polysilicon 681 -2172 681 -2172 0 1
rlabel polysilicon 681 -2178 681 -2178 0 3
rlabel polysilicon 688 -2172 688 -2172 0 1
rlabel polysilicon 688 -2178 688 -2178 0 3
rlabel polysilicon 695 -2172 695 -2172 0 1
rlabel polysilicon 695 -2178 695 -2178 0 3
rlabel polysilicon 702 -2172 702 -2172 0 1
rlabel polysilicon 705 -2172 705 -2172 0 2
rlabel polysilicon 702 -2178 702 -2178 0 3
rlabel polysilicon 712 -2172 712 -2172 0 2
rlabel polysilicon 709 -2178 709 -2178 0 3
rlabel polysilicon 716 -2172 716 -2172 0 1
rlabel polysilicon 716 -2178 716 -2178 0 3
rlabel polysilicon 723 -2172 723 -2172 0 1
rlabel polysilicon 723 -2178 723 -2178 0 3
rlabel polysilicon 730 -2172 730 -2172 0 1
rlabel polysilicon 730 -2178 730 -2178 0 3
rlabel polysilicon 737 -2172 737 -2172 0 1
rlabel polysilicon 737 -2178 737 -2178 0 3
rlabel polysilicon 744 -2172 744 -2172 0 1
rlabel polysilicon 744 -2178 744 -2178 0 3
rlabel polysilicon 751 -2172 751 -2172 0 1
rlabel polysilicon 751 -2178 751 -2178 0 3
rlabel polysilicon 758 -2172 758 -2172 0 1
rlabel polysilicon 758 -2178 758 -2178 0 3
rlabel polysilicon 765 -2172 765 -2172 0 1
rlabel polysilicon 765 -2178 765 -2178 0 3
rlabel polysilicon 772 -2172 772 -2172 0 1
rlabel polysilicon 772 -2178 772 -2178 0 3
rlabel polysilicon 779 -2172 779 -2172 0 1
rlabel polysilicon 779 -2178 779 -2178 0 3
rlabel polysilicon 786 -2172 786 -2172 0 1
rlabel polysilicon 786 -2178 786 -2178 0 3
rlabel polysilicon 793 -2172 793 -2172 0 1
rlabel polysilicon 793 -2178 793 -2178 0 3
rlabel polysilicon 803 -2172 803 -2172 0 2
rlabel polysilicon 803 -2178 803 -2178 0 4
rlabel polysilicon 807 -2172 807 -2172 0 1
rlabel polysilicon 807 -2178 807 -2178 0 3
rlabel polysilicon 814 -2172 814 -2172 0 1
rlabel polysilicon 817 -2172 817 -2172 0 2
rlabel polysilicon 814 -2178 814 -2178 0 3
rlabel polysilicon 817 -2178 817 -2178 0 4
rlabel polysilicon 821 -2172 821 -2172 0 1
rlabel polysilicon 821 -2178 821 -2178 0 3
rlabel polysilicon 824 -2178 824 -2178 0 4
rlabel polysilicon 831 -2172 831 -2172 0 2
rlabel polysilicon 831 -2178 831 -2178 0 4
rlabel polysilicon 835 -2172 835 -2172 0 1
rlabel polysilicon 835 -2178 835 -2178 0 3
rlabel polysilicon 842 -2172 842 -2172 0 1
rlabel polysilicon 842 -2178 842 -2178 0 3
rlabel polysilicon 849 -2172 849 -2172 0 1
rlabel polysilicon 849 -2178 849 -2178 0 3
rlabel polysilicon 856 -2172 856 -2172 0 1
rlabel polysilicon 856 -2178 856 -2178 0 3
rlabel polysilicon 863 -2172 863 -2172 0 1
rlabel polysilicon 863 -2178 863 -2178 0 3
rlabel polysilicon 873 -2172 873 -2172 0 2
rlabel polysilicon 873 -2178 873 -2178 0 4
rlabel polysilicon 877 -2172 877 -2172 0 1
rlabel polysilicon 877 -2178 877 -2178 0 3
rlabel polysilicon 884 -2172 884 -2172 0 1
rlabel polysilicon 884 -2178 884 -2178 0 3
rlabel polysilicon 891 -2172 891 -2172 0 1
rlabel polysilicon 891 -2178 891 -2178 0 3
rlabel polysilicon 898 -2172 898 -2172 0 1
rlabel polysilicon 898 -2178 898 -2178 0 3
rlabel polysilicon 905 -2172 905 -2172 0 1
rlabel polysilicon 905 -2178 905 -2178 0 3
rlabel polysilicon 912 -2172 912 -2172 0 1
rlabel polysilicon 912 -2178 912 -2178 0 3
rlabel polysilicon 919 -2172 919 -2172 0 1
rlabel polysilicon 919 -2178 919 -2178 0 3
rlabel polysilicon 929 -2172 929 -2172 0 2
rlabel polysilicon 926 -2178 926 -2178 0 3
rlabel polysilicon 929 -2178 929 -2178 0 4
rlabel polysilicon 933 -2172 933 -2172 0 1
rlabel polysilicon 933 -2178 933 -2178 0 3
rlabel polysilicon 940 -2172 940 -2172 0 1
rlabel polysilicon 940 -2178 940 -2178 0 3
rlabel polysilicon 947 -2172 947 -2172 0 1
rlabel polysilicon 947 -2178 947 -2178 0 3
rlabel polysilicon 954 -2172 954 -2172 0 1
rlabel polysilicon 954 -2178 954 -2178 0 3
rlabel polysilicon 961 -2172 961 -2172 0 1
rlabel polysilicon 961 -2178 961 -2178 0 3
rlabel polysilicon 968 -2172 968 -2172 0 1
rlabel polysilicon 968 -2178 968 -2178 0 3
rlabel polysilicon 975 -2172 975 -2172 0 1
rlabel polysilicon 978 -2172 978 -2172 0 2
rlabel polysilicon 975 -2178 975 -2178 0 3
rlabel polysilicon 978 -2178 978 -2178 0 4
rlabel polysilicon 982 -2172 982 -2172 0 1
rlabel polysilicon 982 -2178 982 -2178 0 3
rlabel polysilicon 989 -2172 989 -2172 0 1
rlabel polysilicon 989 -2178 989 -2178 0 3
rlabel polysilicon 996 -2172 996 -2172 0 1
rlabel polysilicon 999 -2172 999 -2172 0 2
rlabel polysilicon 996 -2178 996 -2178 0 3
rlabel polysilicon 999 -2178 999 -2178 0 4
rlabel polysilicon 1003 -2172 1003 -2172 0 1
rlabel polysilicon 1003 -2178 1003 -2178 0 3
rlabel polysilicon 1010 -2172 1010 -2172 0 1
rlabel polysilicon 1010 -2178 1010 -2178 0 3
rlabel polysilicon 1017 -2172 1017 -2172 0 1
rlabel polysilicon 1017 -2178 1017 -2178 0 3
rlabel polysilicon 1024 -2172 1024 -2172 0 1
rlabel polysilicon 1027 -2172 1027 -2172 0 2
rlabel polysilicon 1024 -2178 1024 -2178 0 3
rlabel polysilicon 1027 -2178 1027 -2178 0 4
rlabel polysilicon 1031 -2172 1031 -2172 0 1
rlabel polysilicon 1031 -2178 1031 -2178 0 3
rlabel polysilicon 1038 -2172 1038 -2172 0 1
rlabel polysilicon 1038 -2178 1038 -2178 0 3
rlabel polysilicon 1045 -2172 1045 -2172 0 1
rlabel polysilicon 1045 -2178 1045 -2178 0 3
rlabel polysilicon 1052 -2172 1052 -2172 0 1
rlabel polysilicon 1052 -2178 1052 -2178 0 3
rlabel polysilicon 1059 -2172 1059 -2172 0 1
rlabel polysilicon 1062 -2172 1062 -2172 0 2
rlabel polysilicon 1059 -2178 1059 -2178 0 3
rlabel polysilicon 1062 -2178 1062 -2178 0 4
rlabel polysilicon 1066 -2172 1066 -2172 0 1
rlabel polysilicon 1066 -2178 1066 -2178 0 3
rlabel polysilicon 1073 -2172 1073 -2172 0 1
rlabel polysilicon 1073 -2178 1073 -2178 0 3
rlabel polysilicon 1080 -2172 1080 -2172 0 1
rlabel polysilicon 1080 -2178 1080 -2178 0 3
rlabel polysilicon 1087 -2172 1087 -2172 0 1
rlabel polysilicon 1087 -2178 1087 -2178 0 3
rlabel polysilicon 1094 -2172 1094 -2172 0 1
rlabel polysilicon 1094 -2178 1094 -2178 0 3
rlabel polysilicon 1101 -2172 1101 -2172 0 1
rlabel polysilicon 1101 -2178 1101 -2178 0 3
rlabel polysilicon 1108 -2172 1108 -2172 0 1
rlabel polysilicon 1108 -2178 1108 -2178 0 3
rlabel polysilicon 1115 -2172 1115 -2172 0 1
rlabel polysilicon 1115 -2178 1115 -2178 0 3
rlabel polysilicon 1125 -2172 1125 -2172 0 2
rlabel polysilicon 1122 -2178 1122 -2178 0 3
rlabel polysilicon 1125 -2178 1125 -2178 0 4
rlabel polysilicon 1129 -2172 1129 -2172 0 1
rlabel polysilicon 1132 -2172 1132 -2172 0 2
rlabel polysilicon 1129 -2178 1129 -2178 0 3
rlabel polysilicon 1132 -2178 1132 -2178 0 4
rlabel polysilicon 1136 -2172 1136 -2172 0 1
rlabel polysilicon 1136 -2178 1136 -2178 0 3
rlabel polysilicon 1143 -2172 1143 -2172 0 1
rlabel polysilicon 1143 -2178 1143 -2178 0 3
rlabel polysilicon 1150 -2172 1150 -2172 0 1
rlabel polysilicon 1150 -2178 1150 -2178 0 3
rlabel polysilicon 1157 -2172 1157 -2172 0 1
rlabel polysilicon 1157 -2178 1157 -2178 0 3
rlabel polysilicon 1164 -2172 1164 -2172 0 1
rlabel polysilicon 1164 -2178 1164 -2178 0 3
rlabel polysilicon 1171 -2172 1171 -2172 0 1
rlabel polysilicon 1171 -2178 1171 -2178 0 3
rlabel polysilicon 1178 -2172 1178 -2172 0 1
rlabel polysilicon 1178 -2178 1178 -2178 0 3
rlabel polysilicon 1185 -2172 1185 -2172 0 1
rlabel polysilicon 1185 -2178 1185 -2178 0 3
rlabel polysilicon 1192 -2172 1192 -2172 0 1
rlabel polysilicon 1195 -2172 1195 -2172 0 2
rlabel polysilicon 1192 -2178 1192 -2178 0 3
rlabel polysilicon 1195 -2178 1195 -2178 0 4
rlabel polysilicon 1199 -2172 1199 -2172 0 1
rlabel polysilicon 1199 -2178 1199 -2178 0 3
rlabel polysilicon 1206 -2172 1206 -2172 0 1
rlabel polysilicon 1206 -2178 1206 -2178 0 3
rlabel polysilicon 1213 -2172 1213 -2172 0 1
rlabel polysilicon 1213 -2178 1213 -2178 0 3
rlabel polysilicon 1220 -2172 1220 -2172 0 1
rlabel polysilicon 1220 -2178 1220 -2178 0 3
rlabel polysilicon 1227 -2172 1227 -2172 0 1
rlabel polysilicon 1227 -2178 1227 -2178 0 3
rlabel polysilicon 1234 -2172 1234 -2172 0 1
rlabel polysilicon 1234 -2178 1234 -2178 0 3
rlabel polysilicon 1241 -2172 1241 -2172 0 1
rlabel polysilicon 1241 -2178 1241 -2178 0 3
rlabel polysilicon 1248 -2172 1248 -2172 0 1
rlabel polysilicon 1248 -2178 1248 -2178 0 3
rlabel polysilicon 1255 -2172 1255 -2172 0 1
rlabel polysilicon 1255 -2178 1255 -2178 0 3
rlabel polysilicon 1262 -2172 1262 -2172 0 1
rlabel polysilicon 1262 -2178 1262 -2178 0 3
rlabel polysilicon 1269 -2172 1269 -2172 0 1
rlabel polysilicon 1269 -2178 1269 -2178 0 3
rlabel polysilicon 1276 -2172 1276 -2172 0 1
rlabel polysilicon 1276 -2178 1276 -2178 0 3
rlabel polysilicon 1283 -2172 1283 -2172 0 1
rlabel polysilicon 1283 -2178 1283 -2178 0 3
rlabel polysilicon 1290 -2172 1290 -2172 0 1
rlabel polysilicon 1290 -2178 1290 -2178 0 3
rlabel polysilicon 1297 -2172 1297 -2172 0 1
rlabel polysilicon 1297 -2178 1297 -2178 0 3
rlabel polysilicon 1304 -2172 1304 -2172 0 1
rlabel polysilicon 1304 -2178 1304 -2178 0 3
rlabel polysilicon 1311 -2172 1311 -2172 0 1
rlabel polysilicon 1314 -2172 1314 -2172 0 2
rlabel polysilicon 1311 -2178 1311 -2178 0 3
rlabel polysilicon 1314 -2178 1314 -2178 0 4
rlabel polysilicon 1318 -2172 1318 -2172 0 1
rlabel polysilicon 1318 -2178 1318 -2178 0 3
rlabel polysilicon 1325 -2172 1325 -2172 0 1
rlabel polysilicon 1325 -2178 1325 -2178 0 3
rlabel polysilicon 1332 -2172 1332 -2172 0 1
rlabel polysilicon 1332 -2178 1332 -2178 0 3
rlabel polysilicon 1339 -2172 1339 -2172 0 1
rlabel polysilicon 1339 -2178 1339 -2178 0 3
rlabel polysilicon 1346 -2172 1346 -2172 0 1
rlabel polysilicon 1346 -2178 1346 -2178 0 3
rlabel polysilicon 1353 -2172 1353 -2172 0 1
rlabel polysilicon 1353 -2178 1353 -2178 0 3
rlabel polysilicon 1360 -2172 1360 -2172 0 1
rlabel polysilicon 1360 -2178 1360 -2178 0 3
rlabel polysilicon 1367 -2172 1367 -2172 0 1
rlabel polysilicon 1367 -2178 1367 -2178 0 3
rlabel polysilicon 1374 -2172 1374 -2172 0 1
rlabel polysilicon 1374 -2178 1374 -2178 0 3
rlabel polysilicon 1381 -2172 1381 -2172 0 1
rlabel polysilicon 1381 -2178 1381 -2178 0 3
rlabel polysilicon 1388 -2172 1388 -2172 0 1
rlabel polysilicon 1388 -2178 1388 -2178 0 3
rlabel polysilicon 1395 -2172 1395 -2172 0 1
rlabel polysilicon 1395 -2178 1395 -2178 0 3
rlabel polysilicon 1402 -2172 1402 -2172 0 1
rlabel polysilicon 1402 -2178 1402 -2178 0 3
rlabel polysilicon 1409 -2172 1409 -2172 0 1
rlabel polysilicon 1409 -2178 1409 -2178 0 3
rlabel polysilicon 1412 -2178 1412 -2178 0 4
rlabel polysilicon 1416 -2172 1416 -2172 0 1
rlabel polysilicon 1416 -2178 1416 -2178 0 3
rlabel polysilicon 1423 -2172 1423 -2172 0 1
rlabel polysilicon 1423 -2178 1423 -2178 0 3
rlabel polysilicon 1430 -2172 1430 -2172 0 1
rlabel polysilicon 1430 -2178 1430 -2178 0 3
rlabel polysilicon 1437 -2172 1437 -2172 0 1
rlabel polysilicon 1437 -2178 1437 -2178 0 3
rlabel polysilicon 1444 -2172 1444 -2172 0 1
rlabel polysilicon 1444 -2178 1444 -2178 0 3
rlabel polysilicon 1451 -2172 1451 -2172 0 1
rlabel polysilicon 1451 -2178 1451 -2178 0 3
rlabel polysilicon 1458 -2172 1458 -2172 0 1
rlabel polysilicon 1458 -2178 1458 -2178 0 3
rlabel polysilicon 1465 -2172 1465 -2172 0 1
rlabel polysilicon 1465 -2178 1465 -2178 0 3
rlabel polysilicon 1472 -2172 1472 -2172 0 1
rlabel polysilicon 1472 -2178 1472 -2178 0 3
rlabel polysilicon 1479 -2172 1479 -2172 0 1
rlabel polysilicon 1479 -2178 1479 -2178 0 3
rlabel polysilicon 1486 -2172 1486 -2172 0 1
rlabel polysilicon 1486 -2178 1486 -2178 0 3
rlabel polysilicon 1493 -2172 1493 -2172 0 1
rlabel polysilicon 1493 -2178 1493 -2178 0 3
rlabel polysilicon 1500 -2172 1500 -2172 0 1
rlabel polysilicon 1500 -2178 1500 -2178 0 3
rlabel polysilicon 1507 -2172 1507 -2172 0 1
rlabel polysilicon 1507 -2178 1507 -2178 0 3
rlabel polysilicon 1514 -2172 1514 -2172 0 1
rlabel polysilicon 1514 -2178 1514 -2178 0 3
rlabel polysilicon 1521 -2172 1521 -2172 0 1
rlabel polysilicon 1521 -2178 1521 -2178 0 3
rlabel polysilicon 1528 -2172 1528 -2172 0 1
rlabel polysilicon 1528 -2178 1528 -2178 0 3
rlabel polysilicon 1535 -2172 1535 -2172 0 1
rlabel polysilicon 1535 -2178 1535 -2178 0 3
rlabel polysilicon 1542 -2172 1542 -2172 0 1
rlabel polysilicon 1542 -2178 1542 -2178 0 3
rlabel polysilicon 1549 -2172 1549 -2172 0 1
rlabel polysilicon 1549 -2178 1549 -2178 0 3
rlabel polysilicon 1556 -2172 1556 -2172 0 1
rlabel polysilicon 1556 -2178 1556 -2178 0 3
rlabel polysilicon 1563 -2172 1563 -2172 0 1
rlabel polysilicon 1563 -2178 1563 -2178 0 3
rlabel polysilicon 1570 -2172 1570 -2172 0 1
rlabel polysilicon 1570 -2178 1570 -2178 0 3
rlabel polysilicon 1577 -2172 1577 -2172 0 1
rlabel polysilicon 1577 -2178 1577 -2178 0 3
rlabel polysilicon 1584 -2172 1584 -2172 0 1
rlabel polysilicon 1584 -2178 1584 -2178 0 3
rlabel polysilicon 1591 -2172 1591 -2172 0 1
rlabel polysilicon 1594 -2172 1594 -2172 0 2
rlabel polysilicon 1591 -2178 1591 -2178 0 3
rlabel polysilicon 1598 -2172 1598 -2172 0 1
rlabel polysilicon 1598 -2178 1598 -2178 0 3
rlabel polysilicon 1605 -2172 1605 -2172 0 1
rlabel polysilicon 1605 -2178 1605 -2178 0 3
rlabel polysilicon 1612 -2172 1612 -2172 0 1
rlabel polysilicon 1612 -2178 1612 -2178 0 3
rlabel polysilicon 1619 -2172 1619 -2172 0 1
rlabel polysilicon 1619 -2178 1619 -2178 0 3
rlabel polysilicon 1626 -2172 1626 -2172 0 1
rlabel polysilicon 1626 -2178 1626 -2178 0 3
rlabel polysilicon 1633 -2172 1633 -2172 0 1
rlabel polysilicon 1633 -2178 1633 -2178 0 3
rlabel polysilicon 1640 -2172 1640 -2172 0 1
rlabel polysilicon 1640 -2178 1640 -2178 0 3
rlabel polysilicon 1647 -2172 1647 -2172 0 1
rlabel polysilicon 1647 -2178 1647 -2178 0 3
rlabel polysilicon 1654 -2172 1654 -2172 0 1
rlabel polysilicon 1654 -2178 1654 -2178 0 3
rlabel polysilicon 1661 -2172 1661 -2172 0 1
rlabel polysilicon 1661 -2178 1661 -2178 0 3
rlabel polysilicon 1668 -2172 1668 -2172 0 1
rlabel polysilicon 1668 -2178 1668 -2178 0 3
rlabel polysilicon 1675 -2172 1675 -2172 0 1
rlabel polysilicon 1675 -2178 1675 -2178 0 3
rlabel polysilicon 1682 -2172 1682 -2172 0 1
rlabel polysilicon 1682 -2178 1682 -2178 0 3
rlabel polysilicon 1689 -2172 1689 -2172 0 1
rlabel polysilicon 1689 -2178 1689 -2178 0 3
rlabel polysilicon 1696 -2172 1696 -2172 0 1
rlabel polysilicon 1696 -2178 1696 -2178 0 3
rlabel polysilicon 1703 -2172 1703 -2172 0 1
rlabel polysilicon 1703 -2178 1703 -2178 0 3
rlabel polysilicon 1710 -2172 1710 -2172 0 1
rlabel polysilicon 1713 -2172 1713 -2172 0 2
rlabel polysilicon 1710 -2178 1710 -2178 0 3
rlabel polysilicon 1713 -2178 1713 -2178 0 4
rlabel polysilicon 1717 -2178 1717 -2178 0 3
rlabel polysilicon 1720 -2178 1720 -2178 0 4
rlabel polysilicon 1724 -2172 1724 -2172 0 1
rlabel polysilicon 1724 -2178 1724 -2178 0 3
rlabel polysilicon 1731 -2172 1731 -2172 0 1
rlabel polysilicon 1731 -2178 1731 -2178 0 3
rlabel polysilicon 1738 -2172 1738 -2172 0 1
rlabel polysilicon 1738 -2178 1738 -2178 0 3
rlabel polysilicon 30 -2301 30 -2301 0 1
rlabel polysilicon 30 -2307 30 -2307 0 3
rlabel polysilicon 44 -2301 44 -2301 0 1
rlabel polysilicon 44 -2307 44 -2307 0 3
rlabel polysilicon 58 -2301 58 -2301 0 1
rlabel polysilicon 58 -2307 58 -2307 0 3
rlabel polysilicon 65 -2301 65 -2301 0 1
rlabel polysilicon 65 -2307 65 -2307 0 3
rlabel polysilicon 72 -2301 72 -2301 0 1
rlabel polysilicon 72 -2307 72 -2307 0 3
rlabel polysilicon 79 -2301 79 -2301 0 1
rlabel polysilicon 79 -2307 79 -2307 0 3
rlabel polysilicon 86 -2301 86 -2301 0 1
rlabel polysilicon 86 -2307 86 -2307 0 3
rlabel polysilicon 93 -2301 93 -2301 0 1
rlabel polysilicon 93 -2307 93 -2307 0 3
rlabel polysilicon 100 -2301 100 -2301 0 1
rlabel polysilicon 100 -2307 100 -2307 0 3
rlabel polysilicon 107 -2301 107 -2301 0 1
rlabel polysilicon 107 -2307 107 -2307 0 3
rlabel polysilicon 114 -2301 114 -2301 0 1
rlabel polysilicon 114 -2307 114 -2307 0 3
rlabel polysilicon 121 -2301 121 -2301 0 1
rlabel polysilicon 121 -2307 121 -2307 0 3
rlabel polysilicon 128 -2301 128 -2301 0 1
rlabel polysilicon 128 -2307 128 -2307 0 3
rlabel polysilicon 135 -2301 135 -2301 0 1
rlabel polysilicon 138 -2301 138 -2301 0 2
rlabel polysilicon 138 -2307 138 -2307 0 4
rlabel polysilicon 142 -2301 142 -2301 0 1
rlabel polysilicon 145 -2301 145 -2301 0 2
rlabel polysilicon 142 -2307 142 -2307 0 3
rlabel polysilicon 149 -2301 149 -2301 0 1
rlabel polysilicon 152 -2301 152 -2301 0 2
rlabel polysilicon 149 -2307 149 -2307 0 3
rlabel polysilicon 152 -2307 152 -2307 0 4
rlabel polysilicon 156 -2301 156 -2301 0 1
rlabel polysilicon 156 -2307 156 -2307 0 3
rlabel polysilicon 163 -2301 163 -2301 0 1
rlabel polysilicon 163 -2307 163 -2307 0 3
rlabel polysilicon 170 -2301 170 -2301 0 1
rlabel polysilicon 170 -2307 170 -2307 0 3
rlabel polysilicon 177 -2301 177 -2301 0 1
rlabel polysilicon 177 -2307 177 -2307 0 3
rlabel polysilicon 184 -2301 184 -2301 0 1
rlabel polysilicon 184 -2307 184 -2307 0 3
rlabel polysilicon 191 -2301 191 -2301 0 1
rlabel polysilicon 191 -2307 191 -2307 0 3
rlabel polysilicon 198 -2301 198 -2301 0 1
rlabel polysilicon 198 -2307 198 -2307 0 3
rlabel polysilicon 205 -2301 205 -2301 0 1
rlabel polysilicon 208 -2301 208 -2301 0 2
rlabel polysilicon 208 -2307 208 -2307 0 4
rlabel polysilicon 215 -2301 215 -2301 0 2
rlabel polysilicon 212 -2307 212 -2307 0 3
rlabel polysilicon 215 -2307 215 -2307 0 4
rlabel polysilicon 219 -2301 219 -2301 0 1
rlabel polysilicon 219 -2307 219 -2307 0 3
rlabel polysilicon 226 -2301 226 -2301 0 1
rlabel polysilicon 226 -2307 226 -2307 0 3
rlabel polysilicon 233 -2301 233 -2301 0 1
rlabel polysilicon 233 -2307 233 -2307 0 3
rlabel polysilicon 240 -2301 240 -2301 0 1
rlabel polysilicon 240 -2307 240 -2307 0 3
rlabel polysilicon 247 -2301 247 -2301 0 1
rlabel polysilicon 247 -2307 247 -2307 0 3
rlabel polysilicon 254 -2301 254 -2301 0 1
rlabel polysilicon 254 -2307 254 -2307 0 3
rlabel polysilicon 261 -2301 261 -2301 0 1
rlabel polysilicon 261 -2307 261 -2307 0 3
rlabel polysilicon 268 -2301 268 -2301 0 1
rlabel polysilicon 268 -2307 268 -2307 0 3
rlabel polysilicon 275 -2301 275 -2301 0 1
rlabel polysilicon 275 -2307 275 -2307 0 3
rlabel polysilicon 282 -2301 282 -2301 0 1
rlabel polysilicon 285 -2301 285 -2301 0 2
rlabel polysilicon 282 -2307 282 -2307 0 3
rlabel polysilicon 289 -2301 289 -2301 0 1
rlabel polysilicon 289 -2307 289 -2307 0 3
rlabel polysilicon 296 -2301 296 -2301 0 1
rlabel polysilicon 296 -2307 296 -2307 0 3
rlabel polysilicon 303 -2301 303 -2301 0 1
rlabel polysilicon 303 -2307 303 -2307 0 3
rlabel polysilicon 310 -2301 310 -2301 0 1
rlabel polysilicon 310 -2307 310 -2307 0 3
rlabel polysilicon 317 -2301 317 -2301 0 1
rlabel polysilicon 317 -2307 317 -2307 0 3
rlabel polysilicon 324 -2301 324 -2301 0 1
rlabel polysilicon 324 -2307 324 -2307 0 3
rlabel polysilicon 331 -2301 331 -2301 0 1
rlabel polysilicon 331 -2307 331 -2307 0 3
rlabel polysilicon 338 -2301 338 -2301 0 1
rlabel polysilicon 338 -2307 338 -2307 0 3
rlabel polysilicon 345 -2301 345 -2301 0 1
rlabel polysilicon 345 -2307 345 -2307 0 3
rlabel polysilicon 352 -2301 352 -2301 0 1
rlabel polysilicon 352 -2307 352 -2307 0 3
rlabel polysilicon 359 -2301 359 -2301 0 1
rlabel polysilicon 359 -2307 359 -2307 0 3
rlabel polysilicon 366 -2301 366 -2301 0 1
rlabel polysilicon 366 -2307 366 -2307 0 3
rlabel polysilicon 373 -2301 373 -2301 0 1
rlabel polysilicon 373 -2307 373 -2307 0 3
rlabel polysilicon 380 -2301 380 -2301 0 1
rlabel polysilicon 380 -2307 380 -2307 0 3
rlabel polysilicon 387 -2301 387 -2301 0 1
rlabel polysilicon 387 -2307 387 -2307 0 3
rlabel polysilicon 394 -2301 394 -2301 0 1
rlabel polysilicon 394 -2307 394 -2307 0 3
rlabel polysilicon 401 -2301 401 -2301 0 1
rlabel polysilicon 401 -2307 401 -2307 0 3
rlabel polysilicon 408 -2301 408 -2301 0 1
rlabel polysilicon 408 -2307 408 -2307 0 3
rlabel polysilicon 415 -2301 415 -2301 0 1
rlabel polysilicon 415 -2307 415 -2307 0 3
rlabel polysilicon 422 -2301 422 -2301 0 1
rlabel polysilicon 422 -2307 422 -2307 0 3
rlabel polysilicon 429 -2307 429 -2307 0 3
rlabel polysilicon 436 -2301 436 -2301 0 1
rlabel polysilicon 436 -2307 436 -2307 0 3
rlabel polysilicon 443 -2301 443 -2301 0 1
rlabel polysilicon 443 -2307 443 -2307 0 3
rlabel polysilicon 450 -2301 450 -2301 0 1
rlabel polysilicon 450 -2307 450 -2307 0 3
rlabel polysilicon 453 -2307 453 -2307 0 4
rlabel polysilicon 457 -2301 457 -2301 0 1
rlabel polysilicon 457 -2307 457 -2307 0 3
rlabel polysilicon 464 -2301 464 -2301 0 1
rlabel polysilicon 464 -2307 464 -2307 0 3
rlabel polysilicon 471 -2301 471 -2301 0 1
rlabel polysilicon 471 -2307 471 -2307 0 3
rlabel polysilicon 478 -2301 478 -2301 0 1
rlabel polysilicon 478 -2307 478 -2307 0 3
rlabel polysilicon 485 -2301 485 -2301 0 1
rlabel polysilicon 495 -2301 495 -2301 0 2
rlabel polysilicon 492 -2307 492 -2307 0 3
rlabel polysilicon 495 -2307 495 -2307 0 4
rlabel polysilicon 499 -2301 499 -2301 0 1
rlabel polysilicon 499 -2307 499 -2307 0 3
rlabel polysilicon 506 -2301 506 -2301 0 1
rlabel polysilicon 509 -2301 509 -2301 0 2
rlabel polysilicon 506 -2307 506 -2307 0 3
rlabel polysilicon 509 -2307 509 -2307 0 4
rlabel polysilicon 513 -2301 513 -2301 0 1
rlabel polysilicon 513 -2307 513 -2307 0 3
rlabel polysilicon 520 -2301 520 -2301 0 1
rlabel polysilicon 520 -2307 520 -2307 0 3
rlabel polysilicon 527 -2301 527 -2301 0 1
rlabel polysilicon 527 -2307 527 -2307 0 3
rlabel polysilicon 534 -2301 534 -2301 0 1
rlabel polysilicon 534 -2307 534 -2307 0 3
rlabel polysilicon 541 -2301 541 -2301 0 1
rlabel polysilicon 541 -2307 541 -2307 0 3
rlabel polysilicon 548 -2301 548 -2301 0 1
rlabel polysilicon 548 -2307 548 -2307 0 3
rlabel polysilicon 555 -2301 555 -2301 0 1
rlabel polysilicon 555 -2307 555 -2307 0 3
rlabel polysilicon 562 -2301 562 -2301 0 1
rlabel polysilicon 562 -2307 562 -2307 0 3
rlabel polysilicon 569 -2301 569 -2301 0 1
rlabel polysilicon 569 -2307 569 -2307 0 3
rlabel polysilicon 579 -2301 579 -2301 0 2
rlabel polysilicon 576 -2307 576 -2307 0 3
rlabel polysilicon 579 -2307 579 -2307 0 4
rlabel polysilicon 583 -2301 583 -2301 0 1
rlabel polysilicon 583 -2307 583 -2307 0 3
rlabel polysilicon 590 -2301 590 -2301 0 1
rlabel polysilicon 590 -2307 590 -2307 0 3
rlabel polysilicon 597 -2301 597 -2301 0 1
rlabel polysilicon 600 -2301 600 -2301 0 2
rlabel polysilicon 600 -2307 600 -2307 0 4
rlabel polysilicon 604 -2301 604 -2301 0 1
rlabel polysilicon 604 -2307 604 -2307 0 3
rlabel polysilicon 611 -2301 611 -2301 0 1
rlabel polysilicon 611 -2307 611 -2307 0 3
rlabel polysilicon 618 -2301 618 -2301 0 1
rlabel polysilicon 618 -2307 618 -2307 0 3
rlabel polysilicon 628 -2301 628 -2301 0 2
rlabel polysilicon 625 -2307 625 -2307 0 3
rlabel polysilicon 632 -2301 632 -2301 0 1
rlabel polysilicon 632 -2307 632 -2307 0 3
rlabel polysilicon 642 -2301 642 -2301 0 2
rlabel polysilicon 639 -2307 639 -2307 0 3
rlabel polysilicon 642 -2307 642 -2307 0 4
rlabel polysilicon 646 -2301 646 -2301 0 1
rlabel polysilicon 646 -2307 646 -2307 0 3
rlabel polysilicon 653 -2301 653 -2301 0 1
rlabel polysilicon 653 -2307 653 -2307 0 3
rlabel polysilicon 660 -2301 660 -2301 0 1
rlabel polysilicon 660 -2307 660 -2307 0 3
rlabel polysilicon 667 -2301 667 -2301 0 1
rlabel polysilicon 670 -2301 670 -2301 0 2
rlabel polysilicon 670 -2307 670 -2307 0 4
rlabel polysilicon 677 -2301 677 -2301 0 2
rlabel polysilicon 677 -2307 677 -2307 0 4
rlabel polysilicon 681 -2301 681 -2301 0 1
rlabel polysilicon 681 -2307 681 -2307 0 3
rlabel polysilicon 688 -2301 688 -2301 0 1
rlabel polysilicon 691 -2301 691 -2301 0 2
rlabel polysilicon 688 -2307 688 -2307 0 3
rlabel polysilicon 691 -2307 691 -2307 0 4
rlabel polysilicon 698 -2301 698 -2301 0 2
rlabel polysilicon 695 -2307 695 -2307 0 3
rlabel polysilicon 702 -2301 702 -2301 0 1
rlabel polysilicon 705 -2301 705 -2301 0 2
rlabel polysilicon 702 -2307 702 -2307 0 3
rlabel polysilicon 705 -2307 705 -2307 0 4
rlabel polysilicon 709 -2301 709 -2301 0 1
rlabel polysilicon 709 -2307 709 -2307 0 3
rlabel polysilicon 716 -2301 716 -2301 0 1
rlabel polysilicon 716 -2307 716 -2307 0 3
rlabel polysilicon 723 -2301 723 -2301 0 1
rlabel polysilicon 723 -2307 723 -2307 0 3
rlabel polysilicon 730 -2301 730 -2301 0 1
rlabel polysilicon 730 -2307 730 -2307 0 3
rlabel polysilicon 737 -2301 737 -2301 0 1
rlabel polysilicon 737 -2307 737 -2307 0 3
rlabel polysilicon 744 -2301 744 -2301 0 1
rlabel polysilicon 744 -2307 744 -2307 0 3
rlabel polysilicon 751 -2301 751 -2301 0 1
rlabel polysilicon 751 -2307 751 -2307 0 3
rlabel polysilicon 758 -2301 758 -2301 0 1
rlabel polysilicon 761 -2301 761 -2301 0 2
rlabel polysilicon 758 -2307 758 -2307 0 3
rlabel polysilicon 761 -2307 761 -2307 0 4
rlabel polysilicon 765 -2301 765 -2301 0 1
rlabel polysilicon 765 -2307 765 -2307 0 3
rlabel polysilicon 772 -2301 772 -2301 0 1
rlabel polysilicon 772 -2307 772 -2307 0 3
rlabel polysilicon 779 -2301 779 -2301 0 1
rlabel polysilicon 779 -2307 779 -2307 0 3
rlabel polysilicon 782 -2307 782 -2307 0 4
rlabel polysilicon 786 -2301 786 -2301 0 1
rlabel polysilicon 786 -2307 786 -2307 0 3
rlabel polysilicon 793 -2301 793 -2301 0 1
rlabel polysilicon 793 -2307 793 -2307 0 3
rlabel polysilicon 800 -2301 800 -2301 0 1
rlabel polysilicon 800 -2307 800 -2307 0 3
rlabel polysilicon 807 -2301 807 -2301 0 1
rlabel polysilicon 807 -2307 807 -2307 0 3
rlabel polysilicon 814 -2301 814 -2301 0 1
rlabel polysilicon 814 -2307 814 -2307 0 3
rlabel polysilicon 821 -2301 821 -2301 0 1
rlabel polysilicon 821 -2307 821 -2307 0 3
rlabel polysilicon 828 -2301 828 -2301 0 1
rlabel polysilicon 828 -2307 828 -2307 0 3
rlabel polysilicon 835 -2301 835 -2301 0 1
rlabel polysilicon 838 -2301 838 -2301 0 2
rlabel polysilicon 835 -2307 835 -2307 0 3
rlabel polysilicon 838 -2307 838 -2307 0 4
rlabel polysilicon 842 -2301 842 -2301 0 1
rlabel polysilicon 842 -2307 842 -2307 0 3
rlabel polysilicon 849 -2301 849 -2301 0 1
rlabel polysilicon 849 -2307 849 -2307 0 3
rlabel polysilicon 856 -2301 856 -2301 0 1
rlabel polysilicon 856 -2307 856 -2307 0 3
rlabel polysilicon 863 -2301 863 -2301 0 1
rlabel polysilicon 866 -2301 866 -2301 0 2
rlabel polysilicon 863 -2307 863 -2307 0 3
rlabel polysilicon 866 -2307 866 -2307 0 4
rlabel polysilicon 870 -2301 870 -2301 0 1
rlabel polysilicon 873 -2301 873 -2301 0 2
rlabel polysilicon 870 -2307 870 -2307 0 3
rlabel polysilicon 873 -2307 873 -2307 0 4
rlabel polysilicon 877 -2301 877 -2301 0 1
rlabel polysilicon 877 -2307 877 -2307 0 3
rlabel polysilicon 884 -2301 884 -2301 0 1
rlabel polysilicon 884 -2307 884 -2307 0 3
rlabel polysilicon 891 -2301 891 -2301 0 1
rlabel polysilicon 891 -2307 891 -2307 0 3
rlabel polysilicon 898 -2301 898 -2301 0 1
rlabel polysilicon 898 -2307 898 -2307 0 3
rlabel polysilicon 905 -2301 905 -2301 0 1
rlabel polysilicon 905 -2307 905 -2307 0 3
rlabel polysilicon 912 -2301 912 -2301 0 1
rlabel polysilicon 912 -2307 912 -2307 0 3
rlabel polysilicon 915 -2307 915 -2307 0 4
rlabel polysilicon 919 -2301 919 -2301 0 1
rlabel polysilicon 919 -2307 919 -2307 0 3
rlabel polysilicon 926 -2301 926 -2301 0 1
rlabel polysilicon 926 -2307 926 -2307 0 3
rlabel polysilicon 933 -2301 933 -2301 0 1
rlabel polysilicon 933 -2307 933 -2307 0 3
rlabel polysilicon 943 -2301 943 -2301 0 2
rlabel polysilicon 940 -2307 940 -2307 0 3
rlabel polysilicon 943 -2307 943 -2307 0 4
rlabel polysilicon 947 -2301 947 -2301 0 1
rlabel polysilicon 947 -2307 947 -2307 0 3
rlabel polysilicon 954 -2301 954 -2301 0 1
rlabel polysilicon 954 -2307 954 -2307 0 3
rlabel polysilicon 961 -2301 961 -2301 0 1
rlabel polysilicon 961 -2307 961 -2307 0 3
rlabel polysilicon 968 -2301 968 -2301 0 1
rlabel polysilicon 968 -2307 968 -2307 0 3
rlabel polysilicon 975 -2301 975 -2301 0 1
rlabel polysilicon 975 -2307 975 -2307 0 3
rlabel polysilicon 982 -2301 982 -2301 0 1
rlabel polysilicon 982 -2307 982 -2307 0 3
rlabel polysilicon 989 -2301 989 -2301 0 1
rlabel polysilicon 989 -2307 989 -2307 0 3
rlabel polysilicon 992 -2307 992 -2307 0 4
rlabel polysilicon 996 -2301 996 -2301 0 1
rlabel polysilicon 996 -2307 996 -2307 0 3
rlabel polysilicon 1003 -2301 1003 -2301 0 1
rlabel polysilicon 1003 -2307 1003 -2307 0 3
rlabel polysilicon 1010 -2301 1010 -2301 0 1
rlabel polysilicon 1010 -2307 1010 -2307 0 3
rlabel polysilicon 1017 -2301 1017 -2301 0 1
rlabel polysilicon 1020 -2301 1020 -2301 0 2
rlabel polysilicon 1017 -2307 1017 -2307 0 3
rlabel polysilicon 1020 -2307 1020 -2307 0 4
rlabel polysilicon 1024 -2301 1024 -2301 0 1
rlabel polysilicon 1027 -2301 1027 -2301 0 2
rlabel polysilicon 1024 -2307 1024 -2307 0 3
rlabel polysilicon 1031 -2301 1031 -2301 0 1
rlabel polysilicon 1031 -2307 1031 -2307 0 3
rlabel polysilicon 1038 -2301 1038 -2301 0 1
rlabel polysilicon 1041 -2301 1041 -2301 0 2
rlabel polysilicon 1038 -2307 1038 -2307 0 3
rlabel polysilicon 1041 -2307 1041 -2307 0 4
rlabel polysilicon 1045 -2301 1045 -2301 0 1
rlabel polysilicon 1045 -2307 1045 -2307 0 3
rlabel polysilicon 1052 -2301 1052 -2301 0 1
rlabel polysilicon 1052 -2307 1052 -2307 0 3
rlabel polysilicon 1059 -2301 1059 -2301 0 1
rlabel polysilicon 1059 -2307 1059 -2307 0 3
rlabel polysilicon 1066 -2301 1066 -2301 0 1
rlabel polysilicon 1066 -2307 1066 -2307 0 3
rlabel polysilicon 1073 -2301 1073 -2301 0 1
rlabel polysilicon 1073 -2307 1073 -2307 0 3
rlabel polysilicon 1080 -2301 1080 -2301 0 1
rlabel polysilicon 1080 -2307 1080 -2307 0 3
rlabel polysilicon 1087 -2301 1087 -2301 0 1
rlabel polysilicon 1087 -2307 1087 -2307 0 3
rlabel polysilicon 1094 -2301 1094 -2301 0 1
rlabel polysilicon 1094 -2307 1094 -2307 0 3
rlabel polysilicon 1101 -2301 1101 -2301 0 1
rlabel polysilicon 1101 -2307 1101 -2307 0 3
rlabel polysilicon 1108 -2301 1108 -2301 0 1
rlabel polysilicon 1108 -2307 1108 -2307 0 3
rlabel polysilicon 1115 -2301 1115 -2301 0 1
rlabel polysilicon 1115 -2307 1115 -2307 0 3
rlabel polysilicon 1122 -2301 1122 -2301 0 1
rlabel polysilicon 1122 -2307 1122 -2307 0 3
rlabel polysilicon 1129 -2301 1129 -2301 0 1
rlabel polysilicon 1129 -2307 1129 -2307 0 3
rlabel polysilicon 1136 -2301 1136 -2301 0 1
rlabel polysilicon 1136 -2307 1136 -2307 0 3
rlabel polysilicon 1143 -2301 1143 -2301 0 1
rlabel polysilicon 1143 -2307 1143 -2307 0 3
rlabel polysilicon 1150 -2301 1150 -2301 0 1
rlabel polysilicon 1150 -2307 1150 -2307 0 3
rlabel polysilicon 1157 -2301 1157 -2301 0 1
rlabel polysilicon 1157 -2307 1157 -2307 0 3
rlabel polysilicon 1164 -2301 1164 -2301 0 1
rlabel polysilicon 1164 -2307 1164 -2307 0 3
rlabel polysilicon 1174 -2301 1174 -2301 0 2
rlabel polysilicon 1171 -2307 1171 -2307 0 3
rlabel polysilicon 1174 -2307 1174 -2307 0 4
rlabel polysilicon 1178 -2301 1178 -2301 0 1
rlabel polysilicon 1178 -2307 1178 -2307 0 3
rlabel polysilicon 1185 -2301 1185 -2301 0 1
rlabel polysilicon 1185 -2307 1185 -2307 0 3
rlabel polysilicon 1192 -2301 1192 -2301 0 1
rlabel polysilicon 1192 -2307 1192 -2307 0 3
rlabel polysilicon 1202 -2301 1202 -2301 0 2
rlabel polysilicon 1202 -2307 1202 -2307 0 4
rlabel polysilicon 1206 -2301 1206 -2301 0 1
rlabel polysilicon 1206 -2307 1206 -2307 0 3
rlabel polysilicon 1213 -2301 1213 -2301 0 1
rlabel polysilicon 1213 -2307 1213 -2307 0 3
rlabel polysilicon 1220 -2301 1220 -2301 0 1
rlabel polysilicon 1220 -2307 1220 -2307 0 3
rlabel polysilicon 1227 -2301 1227 -2301 0 1
rlabel polysilicon 1227 -2307 1227 -2307 0 3
rlabel polysilicon 1234 -2301 1234 -2301 0 1
rlabel polysilicon 1234 -2307 1234 -2307 0 3
rlabel polysilicon 1241 -2301 1241 -2301 0 1
rlabel polysilicon 1241 -2307 1241 -2307 0 3
rlabel polysilicon 1244 -2307 1244 -2307 0 4
rlabel polysilicon 1248 -2301 1248 -2301 0 1
rlabel polysilicon 1248 -2307 1248 -2307 0 3
rlabel polysilicon 1255 -2301 1255 -2301 0 1
rlabel polysilicon 1255 -2307 1255 -2307 0 3
rlabel polysilicon 1262 -2301 1262 -2301 0 1
rlabel polysilicon 1262 -2307 1262 -2307 0 3
rlabel polysilicon 1269 -2301 1269 -2301 0 1
rlabel polysilicon 1269 -2307 1269 -2307 0 3
rlabel polysilicon 1276 -2301 1276 -2301 0 1
rlabel polysilicon 1276 -2307 1276 -2307 0 3
rlabel polysilicon 1283 -2301 1283 -2301 0 1
rlabel polysilicon 1283 -2307 1283 -2307 0 3
rlabel polysilicon 1290 -2301 1290 -2301 0 1
rlabel polysilicon 1290 -2307 1290 -2307 0 3
rlabel polysilicon 1297 -2301 1297 -2301 0 1
rlabel polysilicon 1297 -2307 1297 -2307 0 3
rlabel polysilicon 1304 -2301 1304 -2301 0 1
rlabel polysilicon 1304 -2307 1304 -2307 0 3
rlabel polysilicon 1311 -2301 1311 -2301 0 1
rlabel polysilicon 1311 -2307 1311 -2307 0 3
rlabel polysilicon 1318 -2301 1318 -2301 0 1
rlabel polysilicon 1318 -2307 1318 -2307 0 3
rlabel polysilicon 1325 -2301 1325 -2301 0 1
rlabel polysilicon 1325 -2307 1325 -2307 0 3
rlabel polysilicon 1332 -2301 1332 -2301 0 1
rlabel polysilicon 1332 -2307 1332 -2307 0 3
rlabel polysilicon 1339 -2301 1339 -2301 0 1
rlabel polysilicon 1339 -2307 1339 -2307 0 3
rlabel polysilicon 1346 -2301 1346 -2301 0 1
rlabel polysilicon 1346 -2307 1346 -2307 0 3
rlabel polysilicon 1353 -2301 1353 -2301 0 1
rlabel polysilicon 1353 -2307 1353 -2307 0 3
rlabel polysilicon 1360 -2301 1360 -2301 0 1
rlabel polysilicon 1360 -2307 1360 -2307 0 3
rlabel polysilicon 1367 -2301 1367 -2301 0 1
rlabel polysilicon 1367 -2307 1367 -2307 0 3
rlabel polysilicon 1374 -2301 1374 -2301 0 1
rlabel polysilicon 1374 -2307 1374 -2307 0 3
rlabel polysilicon 1381 -2301 1381 -2301 0 1
rlabel polysilicon 1381 -2307 1381 -2307 0 3
rlabel polysilicon 1388 -2301 1388 -2301 0 1
rlabel polysilicon 1388 -2307 1388 -2307 0 3
rlabel polysilicon 1395 -2301 1395 -2301 0 1
rlabel polysilicon 1395 -2307 1395 -2307 0 3
rlabel polysilicon 1402 -2301 1402 -2301 0 1
rlabel polysilicon 1402 -2307 1402 -2307 0 3
rlabel polysilicon 1409 -2301 1409 -2301 0 1
rlabel polysilicon 1412 -2301 1412 -2301 0 2
rlabel polysilicon 1409 -2307 1409 -2307 0 3
rlabel polysilicon 1416 -2301 1416 -2301 0 1
rlabel polysilicon 1416 -2307 1416 -2307 0 3
rlabel polysilicon 1423 -2301 1423 -2301 0 1
rlabel polysilicon 1423 -2307 1423 -2307 0 3
rlabel polysilicon 1430 -2301 1430 -2301 0 1
rlabel polysilicon 1430 -2307 1430 -2307 0 3
rlabel polysilicon 1437 -2301 1437 -2301 0 1
rlabel polysilicon 1437 -2307 1437 -2307 0 3
rlabel polysilicon 1444 -2301 1444 -2301 0 1
rlabel polysilicon 1444 -2307 1444 -2307 0 3
rlabel polysilicon 1451 -2301 1451 -2301 0 1
rlabel polysilicon 1451 -2307 1451 -2307 0 3
rlabel polysilicon 1458 -2301 1458 -2301 0 1
rlabel polysilicon 1458 -2307 1458 -2307 0 3
rlabel polysilicon 1465 -2301 1465 -2301 0 1
rlabel polysilicon 1465 -2307 1465 -2307 0 3
rlabel polysilicon 1472 -2301 1472 -2301 0 1
rlabel polysilicon 1472 -2307 1472 -2307 0 3
rlabel polysilicon 1479 -2301 1479 -2301 0 1
rlabel polysilicon 1479 -2307 1479 -2307 0 3
rlabel polysilicon 1486 -2301 1486 -2301 0 1
rlabel polysilicon 1486 -2307 1486 -2307 0 3
rlabel polysilicon 1493 -2301 1493 -2301 0 1
rlabel polysilicon 1493 -2307 1493 -2307 0 3
rlabel polysilicon 1500 -2301 1500 -2301 0 1
rlabel polysilicon 1500 -2307 1500 -2307 0 3
rlabel polysilicon 1507 -2301 1507 -2301 0 1
rlabel polysilicon 1507 -2307 1507 -2307 0 3
rlabel polysilicon 1514 -2301 1514 -2301 0 1
rlabel polysilicon 1514 -2307 1514 -2307 0 3
rlabel polysilicon 1521 -2301 1521 -2301 0 1
rlabel polysilicon 1521 -2307 1521 -2307 0 3
rlabel polysilicon 1528 -2301 1528 -2301 0 1
rlabel polysilicon 1528 -2307 1528 -2307 0 3
rlabel polysilicon 1535 -2301 1535 -2301 0 1
rlabel polysilicon 1535 -2307 1535 -2307 0 3
rlabel polysilicon 1542 -2301 1542 -2301 0 1
rlabel polysilicon 1542 -2307 1542 -2307 0 3
rlabel polysilicon 1549 -2301 1549 -2301 0 1
rlabel polysilicon 1549 -2307 1549 -2307 0 3
rlabel polysilicon 1556 -2301 1556 -2301 0 1
rlabel polysilicon 1556 -2307 1556 -2307 0 3
rlabel polysilicon 1563 -2301 1563 -2301 0 1
rlabel polysilicon 1563 -2307 1563 -2307 0 3
rlabel polysilicon 1570 -2301 1570 -2301 0 1
rlabel polysilicon 1570 -2307 1570 -2307 0 3
rlabel polysilicon 1577 -2301 1577 -2301 0 1
rlabel polysilicon 1577 -2307 1577 -2307 0 3
rlabel polysilicon 1584 -2301 1584 -2301 0 1
rlabel polysilicon 1584 -2307 1584 -2307 0 3
rlabel polysilicon 1591 -2301 1591 -2301 0 1
rlabel polysilicon 1591 -2307 1591 -2307 0 3
rlabel polysilicon 1598 -2301 1598 -2301 0 1
rlabel polysilicon 1598 -2307 1598 -2307 0 3
rlabel polysilicon 1605 -2301 1605 -2301 0 1
rlabel polysilicon 1605 -2307 1605 -2307 0 3
rlabel polysilicon 1612 -2301 1612 -2301 0 1
rlabel polysilicon 1612 -2307 1612 -2307 0 3
rlabel polysilicon 1619 -2301 1619 -2301 0 1
rlabel polysilicon 1619 -2307 1619 -2307 0 3
rlabel polysilicon 1626 -2301 1626 -2301 0 1
rlabel polysilicon 1626 -2307 1626 -2307 0 3
rlabel polysilicon 1633 -2301 1633 -2301 0 1
rlabel polysilicon 1633 -2307 1633 -2307 0 3
rlabel polysilicon 1640 -2301 1640 -2301 0 1
rlabel polysilicon 1640 -2307 1640 -2307 0 3
rlabel polysilicon 1647 -2301 1647 -2301 0 1
rlabel polysilicon 1650 -2301 1650 -2301 0 2
rlabel polysilicon 1647 -2307 1647 -2307 0 3
rlabel polysilicon 1650 -2307 1650 -2307 0 4
rlabel polysilicon 1654 -2307 1654 -2307 0 3
rlabel polysilicon 1661 -2301 1661 -2301 0 1
rlabel polysilicon 1661 -2307 1661 -2307 0 3
rlabel polysilicon 1668 -2301 1668 -2301 0 1
rlabel polysilicon 1671 -2301 1671 -2301 0 2
rlabel polysilicon 1668 -2307 1668 -2307 0 3
rlabel polysilicon 1671 -2307 1671 -2307 0 4
rlabel polysilicon 1675 -2301 1675 -2301 0 1
rlabel polysilicon 1675 -2307 1675 -2307 0 3
rlabel polysilicon 1682 -2301 1682 -2301 0 1
rlabel polysilicon 1682 -2307 1682 -2307 0 3
rlabel polysilicon 1689 -2301 1689 -2301 0 1
rlabel polysilicon 1689 -2307 1689 -2307 0 3
rlabel polysilicon 1696 -2301 1696 -2301 0 1
rlabel polysilicon 1696 -2307 1696 -2307 0 3
rlabel polysilicon 44 -2422 44 -2422 0 1
rlabel polysilicon 44 -2428 44 -2428 0 3
rlabel polysilicon 51 -2422 51 -2422 0 1
rlabel polysilicon 51 -2428 51 -2428 0 3
rlabel polysilicon 58 -2422 58 -2422 0 1
rlabel polysilicon 58 -2428 58 -2428 0 3
rlabel polysilicon 65 -2422 65 -2422 0 1
rlabel polysilicon 65 -2428 65 -2428 0 3
rlabel polysilicon 72 -2422 72 -2422 0 1
rlabel polysilicon 72 -2428 72 -2428 0 3
rlabel polysilicon 79 -2422 79 -2422 0 1
rlabel polysilicon 79 -2428 79 -2428 0 3
rlabel polysilicon 86 -2422 86 -2422 0 1
rlabel polysilicon 86 -2428 86 -2428 0 3
rlabel polysilicon 93 -2422 93 -2422 0 1
rlabel polysilicon 93 -2428 93 -2428 0 3
rlabel polysilicon 100 -2422 100 -2422 0 1
rlabel polysilicon 100 -2428 100 -2428 0 3
rlabel polysilicon 107 -2428 107 -2428 0 3
rlabel polysilicon 110 -2428 110 -2428 0 4
rlabel polysilicon 114 -2422 114 -2422 0 1
rlabel polysilicon 117 -2422 117 -2422 0 2
rlabel polysilicon 114 -2428 114 -2428 0 3
rlabel polysilicon 117 -2428 117 -2428 0 4
rlabel polysilicon 121 -2422 121 -2422 0 1
rlabel polysilicon 121 -2428 121 -2428 0 3
rlabel polysilicon 128 -2422 128 -2422 0 1
rlabel polysilicon 128 -2428 128 -2428 0 3
rlabel polysilicon 135 -2422 135 -2422 0 1
rlabel polysilicon 135 -2428 135 -2428 0 3
rlabel polysilicon 142 -2422 142 -2422 0 1
rlabel polysilicon 142 -2428 142 -2428 0 3
rlabel polysilicon 149 -2422 149 -2422 0 1
rlabel polysilicon 149 -2428 149 -2428 0 3
rlabel polysilicon 156 -2422 156 -2422 0 1
rlabel polysilicon 156 -2428 156 -2428 0 3
rlabel polysilicon 163 -2422 163 -2422 0 1
rlabel polysilicon 163 -2428 163 -2428 0 3
rlabel polysilicon 170 -2422 170 -2422 0 1
rlabel polysilicon 170 -2428 170 -2428 0 3
rlabel polysilicon 177 -2422 177 -2422 0 1
rlabel polysilicon 177 -2428 177 -2428 0 3
rlabel polysilicon 184 -2422 184 -2422 0 1
rlabel polysilicon 184 -2428 184 -2428 0 3
rlabel polysilicon 191 -2422 191 -2422 0 1
rlabel polysilicon 191 -2428 191 -2428 0 3
rlabel polysilicon 198 -2422 198 -2422 0 1
rlabel polysilicon 198 -2428 198 -2428 0 3
rlabel polysilicon 205 -2422 205 -2422 0 1
rlabel polysilicon 205 -2428 205 -2428 0 3
rlabel polysilicon 212 -2422 212 -2422 0 1
rlabel polysilicon 212 -2428 212 -2428 0 3
rlabel polysilicon 219 -2422 219 -2422 0 1
rlabel polysilicon 219 -2428 219 -2428 0 3
rlabel polysilicon 226 -2422 226 -2422 0 1
rlabel polysilicon 229 -2422 229 -2422 0 2
rlabel polysilicon 229 -2428 229 -2428 0 4
rlabel polysilicon 233 -2422 233 -2422 0 1
rlabel polysilicon 233 -2428 233 -2428 0 3
rlabel polysilicon 240 -2422 240 -2422 0 1
rlabel polysilicon 240 -2428 240 -2428 0 3
rlabel polysilicon 247 -2422 247 -2422 0 1
rlabel polysilicon 247 -2428 247 -2428 0 3
rlabel polysilicon 254 -2422 254 -2422 0 1
rlabel polysilicon 254 -2428 254 -2428 0 3
rlabel polysilicon 261 -2422 261 -2422 0 1
rlabel polysilicon 261 -2428 261 -2428 0 3
rlabel polysilicon 268 -2422 268 -2422 0 1
rlabel polysilicon 268 -2428 268 -2428 0 3
rlabel polysilicon 275 -2422 275 -2422 0 1
rlabel polysilicon 275 -2428 275 -2428 0 3
rlabel polysilicon 282 -2422 282 -2422 0 1
rlabel polysilicon 285 -2422 285 -2422 0 2
rlabel polysilicon 282 -2428 282 -2428 0 3
rlabel polysilicon 289 -2422 289 -2422 0 1
rlabel polysilicon 289 -2428 289 -2428 0 3
rlabel polysilicon 296 -2422 296 -2422 0 1
rlabel polysilicon 296 -2428 296 -2428 0 3
rlabel polysilicon 303 -2422 303 -2422 0 1
rlabel polysilicon 303 -2428 303 -2428 0 3
rlabel polysilicon 310 -2422 310 -2422 0 1
rlabel polysilicon 310 -2428 310 -2428 0 3
rlabel polysilicon 317 -2422 317 -2422 0 1
rlabel polysilicon 317 -2428 317 -2428 0 3
rlabel polysilicon 324 -2422 324 -2422 0 1
rlabel polysilicon 324 -2428 324 -2428 0 3
rlabel polysilicon 331 -2422 331 -2422 0 1
rlabel polysilicon 331 -2428 331 -2428 0 3
rlabel polysilicon 338 -2422 338 -2422 0 1
rlabel polysilicon 338 -2428 338 -2428 0 3
rlabel polysilicon 345 -2422 345 -2422 0 1
rlabel polysilicon 345 -2428 345 -2428 0 3
rlabel polysilicon 352 -2422 352 -2422 0 1
rlabel polysilicon 352 -2428 352 -2428 0 3
rlabel polysilicon 359 -2422 359 -2422 0 1
rlabel polysilicon 359 -2428 359 -2428 0 3
rlabel polysilicon 366 -2422 366 -2422 0 1
rlabel polysilicon 366 -2428 366 -2428 0 3
rlabel polysilicon 373 -2422 373 -2422 0 1
rlabel polysilicon 373 -2428 373 -2428 0 3
rlabel polysilicon 380 -2422 380 -2422 0 1
rlabel polysilicon 380 -2428 380 -2428 0 3
rlabel polysilicon 387 -2422 387 -2422 0 1
rlabel polysilicon 387 -2428 387 -2428 0 3
rlabel polysilicon 394 -2422 394 -2422 0 1
rlabel polysilicon 394 -2428 394 -2428 0 3
rlabel polysilicon 401 -2422 401 -2422 0 1
rlabel polysilicon 404 -2422 404 -2422 0 2
rlabel polysilicon 401 -2428 401 -2428 0 3
rlabel polysilicon 404 -2428 404 -2428 0 4
rlabel polysilicon 408 -2422 408 -2422 0 1
rlabel polysilicon 408 -2428 408 -2428 0 3
rlabel polysilicon 415 -2422 415 -2422 0 1
rlabel polysilicon 415 -2428 415 -2428 0 3
rlabel polysilicon 422 -2422 422 -2422 0 1
rlabel polysilicon 422 -2428 422 -2428 0 3
rlabel polysilicon 429 -2422 429 -2422 0 1
rlabel polysilicon 429 -2428 429 -2428 0 3
rlabel polysilicon 436 -2422 436 -2422 0 1
rlabel polysilicon 436 -2428 436 -2428 0 3
rlabel polysilicon 443 -2422 443 -2422 0 1
rlabel polysilicon 443 -2428 443 -2428 0 3
rlabel polysilicon 450 -2422 450 -2422 0 1
rlabel polysilicon 450 -2428 450 -2428 0 3
rlabel polysilicon 457 -2422 457 -2422 0 1
rlabel polysilicon 457 -2428 457 -2428 0 3
rlabel polysilicon 464 -2422 464 -2422 0 1
rlabel polysilicon 464 -2428 464 -2428 0 3
rlabel polysilicon 471 -2422 471 -2422 0 1
rlabel polysilicon 471 -2428 471 -2428 0 3
rlabel polysilicon 478 -2422 478 -2422 0 1
rlabel polysilicon 478 -2428 478 -2428 0 3
rlabel polysilicon 485 -2428 485 -2428 0 3
rlabel polysilicon 492 -2422 492 -2422 0 1
rlabel polysilicon 492 -2428 492 -2428 0 3
rlabel polysilicon 499 -2422 499 -2422 0 1
rlabel polysilicon 499 -2428 499 -2428 0 3
rlabel polysilicon 506 -2422 506 -2422 0 1
rlabel polysilicon 506 -2428 506 -2428 0 3
rlabel polysilicon 513 -2422 513 -2422 0 1
rlabel polysilicon 513 -2428 513 -2428 0 3
rlabel polysilicon 520 -2422 520 -2422 0 1
rlabel polysilicon 523 -2422 523 -2422 0 2
rlabel polysilicon 520 -2428 520 -2428 0 3
rlabel polysilicon 523 -2428 523 -2428 0 4
rlabel polysilicon 527 -2422 527 -2422 0 1
rlabel polysilicon 527 -2428 527 -2428 0 3
rlabel polysilicon 534 -2422 534 -2422 0 1
rlabel polysilicon 534 -2428 534 -2428 0 3
rlabel polysilicon 541 -2422 541 -2422 0 1
rlabel polysilicon 541 -2428 541 -2428 0 3
rlabel polysilicon 548 -2422 548 -2422 0 1
rlabel polysilicon 548 -2428 548 -2428 0 3
rlabel polysilicon 555 -2422 555 -2422 0 1
rlabel polysilicon 555 -2428 555 -2428 0 3
rlabel polysilicon 562 -2422 562 -2422 0 1
rlabel polysilicon 562 -2428 562 -2428 0 3
rlabel polysilicon 565 -2428 565 -2428 0 4
rlabel polysilicon 569 -2422 569 -2422 0 1
rlabel polysilicon 569 -2428 569 -2428 0 3
rlabel polysilicon 576 -2422 576 -2422 0 1
rlabel polysilicon 576 -2428 576 -2428 0 3
rlabel polysilicon 583 -2422 583 -2422 0 1
rlabel polysilicon 586 -2422 586 -2422 0 2
rlabel polysilicon 583 -2428 583 -2428 0 3
rlabel polysilicon 586 -2428 586 -2428 0 4
rlabel polysilicon 590 -2422 590 -2422 0 1
rlabel polysilicon 590 -2428 590 -2428 0 3
rlabel polysilicon 597 -2422 597 -2422 0 1
rlabel polysilicon 597 -2428 597 -2428 0 3
rlabel polysilicon 604 -2422 604 -2422 0 1
rlabel polysilicon 604 -2428 604 -2428 0 3
rlabel polysilicon 611 -2422 611 -2422 0 1
rlabel polysilicon 611 -2428 611 -2428 0 3
rlabel polysilicon 614 -2428 614 -2428 0 4
rlabel polysilicon 618 -2422 618 -2422 0 1
rlabel polysilicon 621 -2422 621 -2422 0 2
rlabel polysilicon 618 -2428 618 -2428 0 3
rlabel polysilicon 621 -2428 621 -2428 0 4
rlabel polysilicon 625 -2422 625 -2422 0 1
rlabel polysilicon 625 -2428 625 -2428 0 3
rlabel polysilicon 632 -2422 632 -2422 0 1
rlabel polysilicon 635 -2422 635 -2422 0 2
rlabel polysilicon 632 -2428 632 -2428 0 3
rlabel polysilicon 639 -2422 639 -2422 0 1
rlabel polysilicon 639 -2428 639 -2428 0 3
rlabel polysilicon 646 -2422 646 -2422 0 1
rlabel polysilicon 649 -2422 649 -2422 0 2
rlabel polysilicon 646 -2428 646 -2428 0 3
rlabel polysilicon 649 -2428 649 -2428 0 4
rlabel polysilicon 653 -2422 653 -2422 0 1
rlabel polysilicon 653 -2428 653 -2428 0 3
rlabel polysilicon 660 -2422 660 -2422 0 1
rlabel polysilicon 660 -2428 660 -2428 0 3
rlabel polysilicon 667 -2422 667 -2422 0 1
rlabel polysilicon 667 -2428 667 -2428 0 3
rlabel polysilicon 674 -2422 674 -2422 0 1
rlabel polysilicon 674 -2428 674 -2428 0 3
rlabel polysilicon 681 -2422 681 -2422 0 1
rlabel polysilicon 684 -2422 684 -2422 0 2
rlabel polysilicon 681 -2428 681 -2428 0 3
rlabel polysilicon 684 -2428 684 -2428 0 4
rlabel polysilicon 688 -2422 688 -2422 0 1
rlabel polysilicon 688 -2428 688 -2428 0 3
rlabel polysilicon 695 -2422 695 -2422 0 1
rlabel polysilicon 695 -2428 695 -2428 0 3
rlabel polysilicon 702 -2422 702 -2422 0 1
rlabel polysilicon 702 -2428 702 -2428 0 3
rlabel polysilicon 709 -2422 709 -2422 0 1
rlabel polysilicon 709 -2428 709 -2428 0 3
rlabel polysilicon 716 -2422 716 -2422 0 1
rlabel polysilicon 716 -2428 716 -2428 0 3
rlabel polysilicon 723 -2422 723 -2422 0 1
rlabel polysilicon 723 -2428 723 -2428 0 3
rlabel polysilicon 730 -2422 730 -2422 0 1
rlabel polysilicon 733 -2422 733 -2422 0 2
rlabel polysilicon 730 -2428 730 -2428 0 3
rlabel polysilicon 733 -2428 733 -2428 0 4
rlabel polysilicon 737 -2422 737 -2422 0 1
rlabel polysilicon 740 -2422 740 -2422 0 2
rlabel polysilicon 737 -2428 737 -2428 0 3
rlabel polysilicon 740 -2428 740 -2428 0 4
rlabel polysilicon 744 -2422 744 -2422 0 1
rlabel polysilicon 747 -2422 747 -2422 0 2
rlabel polysilicon 744 -2428 744 -2428 0 3
rlabel polysilicon 747 -2428 747 -2428 0 4
rlabel polysilicon 751 -2422 751 -2422 0 1
rlabel polysilicon 751 -2428 751 -2428 0 3
rlabel polysilicon 758 -2422 758 -2422 0 1
rlabel polysilicon 758 -2428 758 -2428 0 3
rlabel polysilicon 765 -2422 765 -2422 0 1
rlabel polysilicon 765 -2428 765 -2428 0 3
rlabel polysilicon 772 -2422 772 -2422 0 1
rlabel polysilicon 775 -2422 775 -2422 0 2
rlabel polysilicon 772 -2428 772 -2428 0 3
rlabel polysilicon 775 -2428 775 -2428 0 4
rlabel polysilicon 779 -2422 779 -2422 0 1
rlabel polysilicon 779 -2428 779 -2428 0 3
rlabel polysilicon 786 -2422 786 -2422 0 1
rlabel polysilicon 786 -2428 786 -2428 0 3
rlabel polysilicon 793 -2422 793 -2422 0 1
rlabel polysilicon 793 -2428 793 -2428 0 3
rlabel polysilicon 800 -2422 800 -2422 0 1
rlabel polysilicon 800 -2428 800 -2428 0 3
rlabel polysilicon 807 -2422 807 -2422 0 1
rlabel polysilicon 807 -2428 807 -2428 0 3
rlabel polysilicon 814 -2422 814 -2422 0 1
rlabel polysilicon 814 -2428 814 -2428 0 3
rlabel polysilicon 821 -2422 821 -2422 0 1
rlabel polysilicon 821 -2428 821 -2428 0 3
rlabel polysilicon 828 -2422 828 -2422 0 1
rlabel polysilicon 828 -2428 828 -2428 0 3
rlabel polysilicon 835 -2422 835 -2422 0 1
rlabel polysilicon 835 -2428 835 -2428 0 3
rlabel polysilicon 838 -2428 838 -2428 0 4
rlabel polysilicon 842 -2422 842 -2422 0 1
rlabel polysilicon 842 -2428 842 -2428 0 3
rlabel polysilicon 849 -2428 849 -2428 0 3
rlabel polysilicon 852 -2428 852 -2428 0 4
rlabel polysilicon 859 -2422 859 -2422 0 2
rlabel polysilicon 856 -2428 856 -2428 0 3
rlabel polysilicon 859 -2428 859 -2428 0 4
rlabel polysilicon 863 -2422 863 -2422 0 1
rlabel polysilicon 863 -2428 863 -2428 0 3
rlabel polysilicon 870 -2422 870 -2422 0 1
rlabel polysilicon 870 -2428 870 -2428 0 3
rlabel polysilicon 877 -2422 877 -2422 0 1
rlabel polysilicon 877 -2428 877 -2428 0 3
rlabel polysilicon 884 -2422 884 -2422 0 1
rlabel polysilicon 884 -2428 884 -2428 0 3
rlabel polysilicon 891 -2422 891 -2422 0 1
rlabel polysilicon 891 -2428 891 -2428 0 3
rlabel polysilicon 898 -2422 898 -2422 0 1
rlabel polysilicon 898 -2428 898 -2428 0 3
rlabel polysilicon 905 -2422 905 -2422 0 1
rlabel polysilicon 905 -2428 905 -2428 0 3
rlabel polysilicon 912 -2422 912 -2422 0 1
rlabel polysilicon 912 -2428 912 -2428 0 3
rlabel polysilicon 919 -2422 919 -2422 0 1
rlabel polysilicon 919 -2428 919 -2428 0 3
rlabel polysilicon 926 -2422 926 -2422 0 1
rlabel polysilicon 929 -2422 929 -2422 0 2
rlabel polysilicon 926 -2428 926 -2428 0 3
rlabel polysilicon 929 -2428 929 -2428 0 4
rlabel polysilicon 933 -2422 933 -2422 0 1
rlabel polysilicon 933 -2428 933 -2428 0 3
rlabel polysilicon 940 -2422 940 -2422 0 1
rlabel polysilicon 940 -2428 940 -2428 0 3
rlabel polysilicon 947 -2422 947 -2422 0 1
rlabel polysilicon 947 -2428 947 -2428 0 3
rlabel polysilicon 954 -2422 954 -2422 0 1
rlabel polysilicon 954 -2428 954 -2428 0 3
rlabel polysilicon 961 -2422 961 -2422 0 1
rlabel polysilicon 961 -2428 961 -2428 0 3
rlabel polysilicon 971 -2422 971 -2422 0 2
rlabel polysilicon 968 -2428 968 -2428 0 3
rlabel polysilicon 971 -2428 971 -2428 0 4
rlabel polysilicon 975 -2422 975 -2422 0 1
rlabel polysilicon 975 -2428 975 -2428 0 3
rlabel polysilicon 982 -2422 982 -2422 0 1
rlabel polysilicon 982 -2428 982 -2428 0 3
rlabel polysilicon 989 -2422 989 -2422 0 1
rlabel polysilicon 992 -2422 992 -2422 0 2
rlabel polysilicon 989 -2428 989 -2428 0 3
rlabel polysilicon 996 -2422 996 -2422 0 1
rlabel polysilicon 996 -2428 996 -2428 0 3
rlabel polysilicon 1003 -2422 1003 -2422 0 1
rlabel polysilicon 1003 -2428 1003 -2428 0 3
rlabel polysilicon 1010 -2422 1010 -2422 0 1
rlabel polysilicon 1010 -2428 1010 -2428 0 3
rlabel polysilicon 1017 -2422 1017 -2422 0 1
rlabel polysilicon 1017 -2428 1017 -2428 0 3
rlabel polysilicon 1024 -2422 1024 -2422 0 1
rlabel polysilicon 1024 -2428 1024 -2428 0 3
rlabel polysilicon 1031 -2422 1031 -2422 0 1
rlabel polysilicon 1031 -2428 1031 -2428 0 3
rlabel polysilicon 1038 -2422 1038 -2422 0 1
rlabel polysilicon 1038 -2428 1038 -2428 0 3
rlabel polysilicon 1045 -2422 1045 -2422 0 1
rlabel polysilicon 1045 -2428 1045 -2428 0 3
rlabel polysilicon 1052 -2422 1052 -2422 0 1
rlabel polysilicon 1052 -2428 1052 -2428 0 3
rlabel polysilicon 1059 -2422 1059 -2422 0 1
rlabel polysilicon 1059 -2428 1059 -2428 0 3
rlabel polysilicon 1066 -2422 1066 -2422 0 1
rlabel polysilicon 1066 -2428 1066 -2428 0 3
rlabel polysilicon 1073 -2422 1073 -2422 0 1
rlabel polysilicon 1073 -2428 1073 -2428 0 3
rlabel polysilicon 1080 -2422 1080 -2422 0 1
rlabel polysilicon 1080 -2428 1080 -2428 0 3
rlabel polysilicon 1087 -2422 1087 -2422 0 1
rlabel polysilicon 1087 -2428 1087 -2428 0 3
rlabel polysilicon 1094 -2422 1094 -2422 0 1
rlabel polysilicon 1094 -2428 1094 -2428 0 3
rlabel polysilicon 1104 -2422 1104 -2422 0 2
rlabel polysilicon 1104 -2428 1104 -2428 0 4
rlabel polysilicon 1108 -2422 1108 -2422 0 1
rlabel polysilicon 1108 -2428 1108 -2428 0 3
rlabel polysilicon 1115 -2422 1115 -2422 0 1
rlabel polysilicon 1115 -2428 1115 -2428 0 3
rlabel polysilicon 1122 -2422 1122 -2422 0 1
rlabel polysilicon 1125 -2428 1125 -2428 0 4
rlabel polysilicon 1129 -2422 1129 -2422 0 1
rlabel polysilicon 1129 -2428 1129 -2428 0 3
rlabel polysilicon 1136 -2422 1136 -2422 0 1
rlabel polysilicon 1136 -2428 1136 -2428 0 3
rlabel polysilicon 1143 -2422 1143 -2422 0 1
rlabel polysilicon 1143 -2428 1143 -2428 0 3
rlabel polysilicon 1150 -2422 1150 -2422 0 1
rlabel polysilicon 1150 -2428 1150 -2428 0 3
rlabel polysilicon 1157 -2422 1157 -2422 0 1
rlabel polysilicon 1157 -2428 1157 -2428 0 3
rlabel polysilicon 1164 -2422 1164 -2422 0 1
rlabel polysilicon 1164 -2428 1164 -2428 0 3
rlabel polysilicon 1171 -2422 1171 -2422 0 1
rlabel polysilicon 1171 -2428 1171 -2428 0 3
rlabel polysilicon 1178 -2422 1178 -2422 0 1
rlabel polysilicon 1178 -2428 1178 -2428 0 3
rlabel polysilicon 1185 -2422 1185 -2422 0 1
rlabel polysilicon 1185 -2428 1185 -2428 0 3
rlabel polysilicon 1188 -2428 1188 -2428 0 4
rlabel polysilicon 1192 -2422 1192 -2422 0 1
rlabel polysilicon 1192 -2428 1192 -2428 0 3
rlabel polysilicon 1199 -2422 1199 -2422 0 1
rlabel polysilicon 1202 -2422 1202 -2422 0 2
rlabel polysilicon 1199 -2428 1199 -2428 0 3
rlabel polysilicon 1202 -2428 1202 -2428 0 4
rlabel polysilicon 1206 -2422 1206 -2422 0 1
rlabel polysilicon 1206 -2428 1206 -2428 0 3
rlabel polysilicon 1213 -2422 1213 -2422 0 1
rlabel polysilicon 1213 -2428 1213 -2428 0 3
rlabel polysilicon 1220 -2422 1220 -2422 0 1
rlabel polysilicon 1220 -2428 1220 -2428 0 3
rlabel polysilicon 1227 -2422 1227 -2422 0 1
rlabel polysilicon 1227 -2428 1227 -2428 0 3
rlabel polysilicon 1234 -2422 1234 -2422 0 1
rlabel polysilicon 1237 -2422 1237 -2422 0 2
rlabel polysilicon 1237 -2428 1237 -2428 0 4
rlabel polysilicon 1241 -2422 1241 -2422 0 1
rlabel polysilicon 1241 -2428 1241 -2428 0 3
rlabel polysilicon 1248 -2422 1248 -2422 0 1
rlabel polysilicon 1251 -2422 1251 -2422 0 2
rlabel polysilicon 1251 -2428 1251 -2428 0 4
rlabel polysilicon 1255 -2422 1255 -2422 0 1
rlabel polysilicon 1255 -2428 1255 -2428 0 3
rlabel polysilicon 1262 -2422 1262 -2422 0 1
rlabel polysilicon 1262 -2428 1262 -2428 0 3
rlabel polysilicon 1269 -2422 1269 -2422 0 1
rlabel polysilicon 1269 -2428 1269 -2428 0 3
rlabel polysilicon 1276 -2422 1276 -2422 0 1
rlabel polysilicon 1276 -2428 1276 -2428 0 3
rlabel polysilicon 1283 -2422 1283 -2422 0 1
rlabel polysilicon 1283 -2428 1283 -2428 0 3
rlabel polysilicon 1290 -2422 1290 -2422 0 1
rlabel polysilicon 1293 -2422 1293 -2422 0 2
rlabel polysilicon 1290 -2428 1290 -2428 0 3
rlabel polysilicon 1297 -2422 1297 -2422 0 1
rlabel polysilicon 1297 -2428 1297 -2428 0 3
rlabel polysilicon 1304 -2422 1304 -2422 0 1
rlabel polysilicon 1304 -2428 1304 -2428 0 3
rlabel polysilicon 1311 -2422 1311 -2422 0 1
rlabel polysilicon 1311 -2428 1311 -2428 0 3
rlabel polysilicon 1318 -2422 1318 -2422 0 1
rlabel polysilicon 1318 -2428 1318 -2428 0 3
rlabel polysilicon 1325 -2422 1325 -2422 0 1
rlabel polysilicon 1325 -2428 1325 -2428 0 3
rlabel polysilicon 1332 -2422 1332 -2422 0 1
rlabel polysilicon 1332 -2428 1332 -2428 0 3
rlabel polysilicon 1339 -2422 1339 -2422 0 1
rlabel polysilicon 1339 -2428 1339 -2428 0 3
rlabel polysilicon 1346 -2422 1346 -2422 0 1
rlabel polysilicon 1346 -2428 1346 -2428 0 3
rlabel polysilicon 1353 -2422 1353 -2422 0 1
rlabel polysilicon 1353 -2428 1353 -2428 0 3
rlabel polysilicon 1363 -2422 1363 -2422 0 2
rlabel polysilicon 1360 -2428 1360 -2428 0 3
rlabel polysilicon 1363 -2428 1363 -2428 0 4
rlabel polysilicon 1367 -2422 1367 -2422 0 1
rlabel polysilicon 1367 -2428 1367 -2428 0 3
rlabel polysilicon 1374 -2422 1374 -2422 0 1
rlabel polysilicon 1374 -2428 1374 -2428 0 3
rlabel polysilicon 1381 -2422 1381 -2422 0 1
rlabel polysilicon 1381 -2428 1381 -2428 0 3
rlabel polysilicon 1384 -2428 1384 -2428 0 4
rlabel polysilicon 1388 -2422 1388 -2422 0 1
rlabel polysilicon 1388 -2428 1388 -2428 0 3
rlabel polysilicon 1395 -2422 1395 -2422 0 1
rlabel polysilicon 1395 -2428 1395 -2428 0 3
rlabel polysilicon 1402 -2422 1402 -2422 0 1
rlabel polysilicon 1402 -2428 1402 -2428 0 3
rlabel polysilicon 1409 -2422 1409 -2422 0 1
rlabel polysilicon 1409 -2428 1409 -2428 0 3
rlabel polysilicon 1416 -2422 1416 -2422 0 1
rlabel polysilicon 1416 -2428 1416 -2428 0 3
rlabel polysilicon 1423 -2422 1423 -2422 0 1
rlabel polysilicon 1423 -2428 1423 -2428 0 3
rlabel polysilicon 1430 -2422 1430 -2422 0 1
rlabel polysilicon 1430 -2428 1430 -2428 0 3
rlabel polysilicon 1437 -2422 1437 -2422 0 1
rlabel polysilicon 1437 -2428 1437 -2428 0 3
rlabel polysilicon 1444 -2422 1444 -2422 0 1
rlabel polysilicon 1444 -2428 1444 -2428 0 3
rlabel polysilicon 1451 -2422 1451 -2422 0 1
rlabel polysilicon 1451 -2428 1451 -2428 0 3
rlabel polysilicon 1458 -2422 1458 -2422 0 1
rlabel polysilicon 1458 -2428 1458 -2428 0 3
rlabel polysilicon 1465 -2422 1465 -2422 0 1
rlabel polysilicon 1465 -2428 1465 -2428 0 3
rlabel polysilicon 1472 -2422 1472 -2422 0 1
rlabel polysilicon 1472 -2428 1472 -2428 0 3
rlabel polysilicon 1479 -2422 1479 -2422 0 1
rlabel polysilicon 1479 -2428 1479 -2428 0 3
rlabel polysilicon 1486 -2422 1486 -2422 0 1
rlabel polysilicon 1486 -2428 1486 -2428 0 3
rlabel polysilicon 1493 -2422 1493 -2422 0 1
rlabel polysilicon 1493 -2428 1493 -2428 0 3
rlabel polysilicon 1500 -2422 1500 -2422 0 1
rlabel polysilicon 1500 -2428 1500 -2428 0 3
rlabel polysilicon 1507 -2422 1507 -2422 0 1
rlabel polysilicon 1507 -2428 1507 -2428 0 3
rlabel polysilicon 1514 -2422 1514 -2422 0 1
rlabel polysilicon 1514 -2428 1514 -2428 0 3
rlabel polysilicon 1521 -2422 1521 -2422 0 1
rlabel polysilicon 1521 -2428 1521 -2428 0 3
rlabel polysilicon 1528 -2422 1528 -2422 0 1
rlabel polysilicon 1528 -2428 1528 -2428 0 3
rlabel polysilicon 1535 -2422 1535 -2422 0 1
rlabel polysilicon 1535 -2428 1535 -2428 0 3
rlabel polysilicon 1542 -2422 1542 -2422 0 1
rlabel polysilicon 1542 -2428 1542 -2428 0 3
rlabel polysilicon 1549 -2422 1549 -2422 0 1
rlabel polysilicon 1549 -2428 1549 -2428 0 3
rlabel polysilicon 1556 -2422 1556 -2422 0 1
rlabel polysilicon 1556 -2428 1556 -2428 0 3
rlabel polysilicon 1563 -2422 1563 -2422 0 1
rlabel polysilicon 1563 -2428 1563 -2428 0 3
rlabel polysilicon 1570 -2422 1570 -2422 0 1
rlabel polysilicon 1570 -2428 1570 -2428 0 3
rlabel polysilicon 1577 -2422 1577 -2422 0 1
rlabel polysilicon 1577 -2428 1577 -2428 0 3
rlabel polysilicon 1584 -2422 1584 -2422 0 1
rlabel polysilicon 1584 -2428 1584 -2428 0 3
rlabel polysilicon 1591 -2422 1591 -2422 0 1
rlabel polysilicon 1591 -2428 1591 -2428 0 3
rlabel polysilicon 1598 -2422 1598 -2422 0 1
rlabel polysilicon 1598 -2428 1598 -2428 0 3
rlabel polysilicon 1605 -2422 1605 -2422 0 1
rlabel polysilicon 1605 -2428 1605 -2428 0 3
rlabel polysilicon 1612 -2422 1612 -2422 0 1
rlabel polysilicon 1612 -2428 1612 -2428 0 3
rlabel polysilicon 1619 -2422 1619 -2422 0 1
rlabel polysilicon 1622 -2422 1622 -2422 0 2
rlabel polysilicon 1619 -2428 1619 -2428 0 3
rlabel polysilicon 1622 -2428 1622 -2428 0 4
rlabel polysilicon 1626 -2422 1626 -2422 0 1
rlabel polysilicon 1626 -2428 1626 -2428 0 3
rlabel polysilicon 1633 -2422 1633 -2422 0 1
rlabel polysilicon 1633 -2428 1633 -2428 0 3
rlabel polysilicon 1640 -2428 1640 -2428 0 3
rlabel polysilicon 1643 -2428 1643 -2428 0 4
rlabel polysilicon 1650 -2422 1650 -2422 0 2
rlabel polysilicon 1647 -2428 1647 -2428 0 3
rlabel polysilicon 1650 -2428 1650 -2428 0 4
rlabel polysilicon 1654 -2422 1654 -2422 0 1
rlabel polysilicon 1654 -2428 1654 -2428 0 3
rlabel polysilicon 1661 -2422 1661 -2422 0 1
rlabel polysilicon 1661 -2428 1661 -2428 0 3
rlabel polysilicon 51 -2541 51 -2541 0 1
rlabel polysilicon 51 -2547 51 -2547 0 3
rlabel polysilicon 58 -2541 58 -2541 0 1
rlabel polysilicon 58 -2547 58 -2547 0 3
rlabel polysilicon 65 -2541 65 -2541 0 1
rlabel polysilicon 65 -2547 65 -2547 0 3
rlabel polysilicon 72 -2541 72 -2541 0 1
rlabel polysilicon 72 -2547 72 -2547 0 3
rlabel polysilicon 79 -2541 79 -2541 0 1
rlabel polysilicon 79 -2547 79 -2547 0 3
rlabel polysilicon 86 -2541 86 -2541 0 1
rlabel polysilicon 89 -2541 89 -2541 0 2
rlabel polysilicon 86 -2547 86 -2547 0 3
rlabel polysilicon 89 -2547 89 -2547 0 4
rlabel polysilicon 93 -2541 93 -2541 0 1
rlabel polysilicon 93 -2547 93 -2547 0 3
rlabel polysilicon 100 -2541 100 -2541 0 1
rlabel polysilicon 100 -2547 100 -2547 0 3
rlabel polysilicon 107 -2541 107 -2541 0 1
rlabel polysilicon 107 -2547 107 -2547 0 3
rlabel polysilicon 114 -2541 114 -2541 0 1
rlabel polysilicon 114 -2547 114 -2547 0 3
rlabel polysilicon 121 -2541 121 -2541 0 1
rlabel polysilicon 121 -2547 121 -2547 0 3
rlabel polysilicon 128 -2541 128 -2541 0 1
rlabel polysilicon 128 -2547 128 -2547 0 3
rlabel polysilicon 135 -2541 135 -2541 0 1
rlabel polysilicon 135 -2547 135 -2547 0 3
rlabel polysilicon 142 -2541 142 -2541 0 1
rlabel polysilicon 142 -2547 142 -2547 0 3
rlabel polysilicon 149 -2541 149 -2541 0 1
rlabel polysilicon 149 -2547 149 -2547 0 3
rlabel polysilicon 156 -2541 156 -2541 0 1
rlabel polysilicon 156 -2547 156 -2547 0 3
rlabel polysilicon 163 -2541 163 -2541 0 1
rlabel polysilicon 163 -2547 163 -2547 0 3
rlabel polysilicon 170 -2541 170 -2541 0 1
rlabel polysilicon 173 -2541 173 -2541 0 2
rlabel polysilicon 170 -2547 170 -2547 0 3
rlabel polysilicon 177 -2541 177 -2541 0 1
rlabel polysilicon 177 -2547 177 -2547 0 3
rlabel polysilicon 184 -2541 184 -2541 0 1
rlabel polysilicon 184 -2547 184 -2547 0 3
rlabel polysilicon 191 -2541 191 -2541 0 1
rlabel polysilicon 191 -2547 191 -2547 0 3
rlabel polysilicon 198 -2541 198 -2541 0 1
rlabel polysilicon 198 -2547 198 -2547 0 3
rlabel polysilicon 205 -2541 205 -2541 0 1
rlabel polysilicon 205 -2547 205 -2547 0 3
rlabel polysilicon 212 -2541 212 -2541 0 1
rlabel polysilicon 215 -2541 215 -2541 0 2
rlabel polysilicon 212 -2547 212 -2547 0 3
rlabel polysilicon 215 -2547 215 -2547 0 4
rlabel polysilicon 219 -2541 219 -2541 0 1
rlabel polysilicon 219 -2547 219 -2547 0 3
rlabel polysilicon 226 -2541 226 -2541 0 1
rlabel polysilicon 226 -2547 226 -2547 0 3
rlabel polysilicon 233 -2541 233 -2541 0 1
rlabel polysilicon 233 -2547 233 -2547 0 3
rlabel polysilicon 240 -2541 240 -2541 0 1
rlabel polysilicon 240 -2547 240 -2547 0 3
rlabel polysilicon 247 -2541 247 -2541 0 1
rlabel polysilicon 247 -2547 247 -2547 0 3
rlabel polysilicon 254 -2541 254 -2541 0 1
rlabel polysilicon 257 -2541 257 -2541 0 2
rlabel polysilicon 254 -2547 254 -2547 0 3
rlabel polysilicon 257 -2547 257 -2547 0 4
rlabel polysilicon 261 -2541 261 -2541 0 1
rlabel polysilicon 261 -2547 261 -2547 0 3
rlabel polysilicon 268 -2541 268 -2541 0 1
rlabel polysilicon 268 -2547 268 -2547 0 3
rlabel polysilicon 275 -2541 275 -2541 0 1
rlabel polysilicon 278 -2541 278 -2541 0 2
rlabel polysilicon 275 -2547 275 -2547 0 3
rlabel polysilicon 278 -2547 278 -2547 0 4
rlabel polysilicon 282 -2541 282 -2541 0 1
rlabel polysilicon 285 -2541 285 -2541 0 2
rlabel polysilicon 282 -2547 282 -2547 0 3
rlabel polysilicon 289 -2541 289 -2541 0 1
rlabel polysilicon 289 -2547 289 -2547 0 3
rlabel polysilicon 292 -2547 292 -2547 0 4
rlabel polysilicon 296 -2541 296 -2541 0 1
rlabel polysilicon 303 -2541 303 -2541 0 1
rlabel polysilicon 303 -2547 303 -2547 0 3
rlabel polysilicon 310 -2541 310 -2541 0 1
rlabel polysilicon 310 -2547 310 -2547 0 3
rlabel polysilicon 317 -2541 317 -2541 0 1
rlabel polysilicon 317 -2547 317 -2547 0 3
rlabel polysilicon 324 -2541 324 -2541 0 1
rlabel polysilicon 324 -2547 324 -2547 0 3
rlabel polysilicon 331 -2541 331 -2541 0 1
rlabel polysilicon 331 -2547 331 -2547 0 3
rlabel polysilicon 338 -2541 338 -2541 0 1
rlabel polysilicon 338 -2547 338 -2547 0 3
rlabel polysilicon 345 -2541 345 -2541 0 1
rlabel polysilicon 345 -2547 345 -2547 0 3
rlabel polysilicon 352 -2541 352 -2541 0 1
rlabel polysilicon 352 -2547 352 -2547 0 3
rlabel polysilicon 359 -2541 359 -2541 0 1
rlabel polysilicon 359 -2547 359 -2547 0 3
rlabel polysilicon 366 -2541 366 -2541 0 1
rlabel polysilicon 366 -2547 366 -2547 0 3
rlabel polysilicon 373 -2541 373 -2541 0 1
rlabel polysilicon 373 -2547 373 -2547 0 3
rlabel polysilicon 380 -2541 380 -2541 0 1
rlabel polysilicon 380 -2547 380 -2547 0 3
rlabel polysilicon 387 -2541 387 -2541 0 1
rlabel polysilicon 390 -2541 390 -2541 0 2
rlabel polysilicon 390 -2547 390 -2547 0 4
rlabel polysilicon 394 -2541 394 -2541 0 1
rlabel polysilicon 394 -2547 394 -2547 0 3
rlabel polysilicon 401 -2541 401 -2541 0 1
rlabel polysilicon 401 -2547 401 -2547 0 3
rlabel polysilicon 408 -2541 408 -2541 0 1
rlabel polysilicon 408 -2547 408 -2547 0 3
rlabel polysilicon 415 -2547 415 -2547 0 3
rlabel polysilicon 418 -2547 418 -2547 0 4
rlabel polysilicon 422 -2541 422 -2541 0 1
rlabel polysilicon 422 -2547 422 -2547 0 3
rlabel polysilicon 429 -2541 429 -2541 0 1
rlabel polysilicon 429 -2547 429 -2547 0 3
rlabel polysilicon 436 -2541 436 -2541 0 1
rlabel polysilicon 436 -2547 436 -2547 0 3
rlabel polysilicon 443 -2541 443 -2541 0 1
rlabel polysilicon 443 -2547 443 -2547 0 3
rlabel polysilicon 450 -2541 450 -2541 0 1
rlabel polysilicon 450 -2547 450 -2547 0 3
rlabel polysilicon 457 -2541 457 -2541 0 1
rlabel polysilicon 457 -2547 457 -2547 0 3
rlabel polysilicon 464 -2541 464 -2541 0 1
rlabel polysilicon 464 -2547 464 -2547 0 3
rlabel polysilicon 471 -2541 471 -2541 0 1
rlabel polysilicon 471 -2547 471 -2547 0 3
rlabel polysilicon 478 -2541 478 -2541 0 1
rlabel polysilicon 481 -2541 481 -2541 0 2
rlabel polysilicon 481 -2547 481 -2547 0 4
rlabel polysilicon 485 -2541 485 -2541 0 1
rlabel polysilicon 485 -2547 485 -2547 0 3
rlabel polysilicon 492 -2541 492 -2541 0 1
rlabel polysilicon 492 -2547 492 -2547 0 3
rlabel polysilicon 499 -2541 499 -2541 0 1
rlabel polysilicon 499 -2547 499 -2547 0 3
rlabel polysilicon 506 -2541 506 -2541 0 1
rlabel polysilicon 506 -2547 506 -2547 0 3
rlabel polysilicon 513 -2541 513 -2541 0 1
rlabel polysilicon 513 -2547 513 -2547 0 3
rlabel polysilicon 520 -2541 520 -2541 0 1
rlabel polysilicon 520 -2547 520 -2547 0 3
rlabel polysilicon 527 -2541 527 -2541 0 1
rlabel polysilicon 530 -2541 530 -2541 0 2
rlabel polysilicon 530 -2547 530 -2547 0 4
rlabel polysilicon 534 -2541 534 -2541 0 1
rlabel polysilicon 534 -2547 534 -2547 0 3
rlabel polysilicon 541 -2541 541 -2541 0 1
rlabel polysilicon 541 -2547 541 -2547 0 3
rlabel polysilicon 544 -2547 544 -2547 0 4
rlabel polysilicon 548 -2541 548 -2541 0 1
rlabel polysilicon 548 -2547 548 -2547 0 3
rlabel polysilicon 555 -2541 555 -2541 0 1
rlabel polysilicon 555 -2547 555 -2547 0 3
rlabel polysilicon 562 -2541 562 -2541 0 1
rlabel polysilicon 565 -2541 565 -2541 0 2
rlabel polysilicon 562 -2547 562 -2547 0 3
rlabel polysilicon 565 -2547 565 -2547 0 4
rlabel polysilicon 569 -2541 569 -2541 0 1
rlabel polysilicon 572 -2541 572 -2541 0 2
rlabel polysilicon 569 -2547 569 -2547 0 3
rlabel polysilicon 572 -2547 572 -2547 0 4
rlabel polysilicon 576 -2541 576 -2541 0 1
rlabel polysilicon 576 -2547 576 -2547 0 3
rlabel polysilicon 583 -2541 583 -2541 0 1
rlabel polysilicon 583 -2547 583 -2547 0 3
rlabel polysilicon 590 -2541 590 -2541 0 1
rlabel polysilicon 590 -2547 590 -2547 0 3
rlabel polysilicon 597 -2541 597 -2541 0 1
rlabel polysilicon 600 -2541 600 -2541 0 2
rlabel polysilicon 597 -2547 597 -2547 0 3
rlabel polysilicon 600 -2547 600 -2547 0 4
rlabel polysilicon 604 -2541 604 -2541 0 1
rlabel polysilicon 604 -2547 604 -2547 0 3
rlabel polysilicon 611 -2541 611 -2541 0 1
rlabel polysilicon 611 -2547 611 -2547 0 3
rlabel polysilicon 618 -2541 618 -2541 0 1
rlabel polysilicon 618 -2547 618 -2547 0 3
rlabel polysilicon 625 -2541 625 -2541 0 1
rlabel polysilicon 625 -2547 625 -2547 0 3
rlabel polysilicon 632 -2541 632 -2541 0 1
rlabel polysilicon 632 -2547 632 -2547 0 3
rlabel polysilicon 639 -2541 639 -2541 0 1
rlabel polysilicon 639 -2547 639 -2547 0 3
rlabel polysilicon 646 -2541 646 -2541 0 1
rlabel polysilicon 646 -2547 646 -2547 0 3
rlabel polysilicon 653 -2541 653 -2541 0 1
rlabel polysilicon 653 -2547 653 -2547 0 3
rlabel polysilicon 660 -2541 660 -2541 0 1
rlabel polysilicon 660 -2547 660 -2547 0 3
rlabel polysilicon 667 -2547 667 -2547 0 3
rlabel polysilicon 670 -2547 670 -2547 0 4
rlabel polysilicon 674 -2541 674 -2541 0 1
rlabel polysilicon 674 -2547 674 -2547 0 3
rlabel polysilicon 681 -2541 681 -2541 0 1
rlabel polysilicon 681 -2547 681 -2547 0 3
rlabel polysilicon 688 -2541 688 -2541 0 1
rlabel polysilicon 688 -2547 688 -2547 0 3
rlabel polysilicon 695 -2541 695 -2541 0 1
rlabel polysilicon 695 -2547 695 -2547 0 3
rlabel polysilicon 702 -2541 702 -2541 0 1
rlabel polysilicon 702 -2547 702 -2547 0 3
rlabel polysilicon 709 -2541 709 -2541 0 1
rlabel polysilicon 709 -2547 709 -2547 0 3
rlabel polysilicon 716 -2541 716 -2541 0 1
rlabel polysilicon 716 -2547 716 -2547 0 3
rlabel polysilicon 723 -2541 723 -2541 0 1
rlabel polysilicon 723 -2547 723 -2547 0 3
rlabel polysilicon 730 -2541 730 -2541 0 1
rlabel polysilicon 730 -2547 730 -2547 0 3
rlabel polysilicon 733 -2547 733 -2547 0 4
rlabel polysilicon 737 -2541 737 -2541 0 1
rlabel polysilicon 740 -2541 740 -2541 0 2
rlabel polysilicon 737 -2547 737 -2547 0 3
rlabel polysilicon 740 -2547 740 -2547 0 4
rlabel polysilicon 744 -2541 744 -2541 0 1
rlabel polysilicon 744 -2547 744 -2547 0 3
rlabel polysilicon 747 -2547 747 -2547 0 4
rlabel polysilicon 751 -2547 751 -2547 0 3
rlabel polysilicon 754 -2547 754 -2547 0 4
rlabel polysilicon 758 -2541 758 -2541 0 1
rlabel polysilicon 758 -2547 758 -2547 0 3
rlabel polysilicon 765 -2541 765 -2541 0 1
rlabel polysilicon 765 -2547 765 -2547 0 3
rlabel polysilicon 772 -2541 772 -2541 0 1
rlabel polysilicon 772 -2547 772 -2547 0 3
rlabel polysilicon 779 -2541 779 -2541 0 1
rlabel polysilicon 779 -2547 779 -2547 0 3
rlabel polysilicon 786 -2541 786 -2541 0 1
rlabel polysilicon 786 -2547 786 -2547 0 3
rlabel polysilicon 789 -2547 789 -2547 0 4
rlabel polysilicon 793 -2541 793 -2541 0 1
rlabel polysilicon 793 -2547 793 -2547 0 3
rlabel polysilicon 800 -2541 800 -2541 0 1
rlabel polysilicon 803 -2541 803 -2541 0 2
rlabel polysilicon 800 -2547 800 -2547 0 3
rlabel polysilicon 803 -2547 803 -2547 0 4
rlabel polysilicon 807 -2541 807 -2541 0 1
rlabel polysilicon 810 -2541 810 -2541 0 2
rlabel polysilicon 810 -2547 810 -2547 0 4
rlabel polysilicon 814 -2541 814 -2541 0 1
rlabel polysilicon 814 -2547 814 -2547 0 3
rlabel polysilicon 821 -2541 821 -2541 0 1
rlabel polysilicon 821 -2547 821 -2547 0 3
rlabel polysilicon 828 -2541 828 -2541 0 1
rlabel polysilicon 831 -2541 831 -2541 0 2
rlabel polysilicon 828 -2547 828 -2547 0 3
rlabel polysilicon 831 -2547 831 -2547 0 4
rlabel polysilicon 835 -2541 835 -2541 0 1
rlabel polysilicon 835 -2547 835 -2547 0 3
rlabel polysilicon 842 -2541 842 -2541 0 1
rlabel polysilicon 842 -2547 842 -2547 0 3
rlabel polysilicon 849 -2541 849 -2541 0 1
rlabel polysilicon 849 -2547 849 -2547 0 3
rlabel polysilicon 856 -2541 856 -2541 0 1
rlabel polysilicon 856 -2547 856 -2547 0 3
rlabel polysilicon 863 -2541 863 -2541 0 1
rlabel polysilicon 863 -2547 863 -2547 0 3
rlabel polysilicon 870 -2541 870 -2541 0 1
rlabel polysilicon 870 -2547 870 -2547 0 3
rlabel polysilicon 877 -2541 877 -2541 0 1
rlabel polysilicon 877 -2547 877 -2547 0 3
rlabel polysilicon 884 -2541 884 -2541 0 1
rlabel polysilicon 884 -2547 884 -2547 0 3
rlabel polysilicon 891 -2541 891 -2541 0 1
rlabel polysilicon 891 -2547 891 -2547 0 3
rlabel polysilicon 901 -2541 901 -2541 0 2
rlabel polysilicon 898 -2547 898 -2547 0 3
rlabel polysilicon 901 -2547 901 -2547 0 4
rlabel polysilicon 905 -2541 905 -2541 0 1
rlabel polysilicon 905 -2547 905 -2547 0 3
rlabel polysilicon 912 -2541 912 -2541 0 1
rlabel polysilicon 912 -2547 912 -2547 0 3
rlabel polysilicon 919 -2541 919 -2541 0 1
rlabel polysilicon 919 -2547 919 -2547 0 3
rlabel polysilicon 926 -2541 926 -2541 0 1
rlabel polysilicon 926 -2547 926 -2547 0 3
rlabel polysilicon 933 -2541 933 -2541 0 1
rlabel polysilicon 933 -2547 933 -2547 0 3
rlabel polysilicon 940 -2541 940 -2541 0 1
rlabel polysilicon 940 -2547 940 -2547 0 3
rlabel polysilicon 947 -2541 947 -2541 0 1
rlabel polysilicon 947 -2547 947 -2547 0 3
rlabel polysilicon 954 -2541 954 -2541 0 1
rlabel polysilicon 954 -2547 954 -2547 0 3
rlabel polysilicon 961 -2541 961 -2541 0 1
rlabel polysilicon 961 -2547 961 -2547 0 3
rlabel polysilicon 968 -2541 968 -2541 0 1
rlabel polysilicon 968 -2547 968 -2547 0 3
rlabel polysilicon 975 -2541 975 -2541 0 1
rlabel polysilicon 975 -2547 975 -2547 0 3
rlabel polysilicon 982 -2541 982 -2541 0 1
rlabel polysilicon 982 -2547 982 -2547 0 3
rlabel polysilicon 989 -2541 989 -2541 0 1
rlabel polysilicon 989 -2547 989 -2547 0 3
rlabel polysilicon 996 -2541 996 -2541 0 1
rlabel polysilicon 996 -2547 996 -2547 0 3
rlabel polysilicon 1003 -2541 1003 -2541 0 1
rlabel polysilicon 1003 -2547 1003 -2547 0 3
rlabel polysilicon 1010 -2541 1010 -2541 0 1
rlabel polysilicon 1013 -2541 1013 -2541 0 2
rlabel polysilicon 1010 -2547 1010 -2547 0 3
rlabel polysilicon 1017 -2541 1017 -2541 0 1
rlabel polysilicon 1017 -2547 1017 -2547 0 3
rlabel polysilicon 1024 -2541 1024 -2541 0 1
rlabel polysilicon 1027 -2541 1027 -2541 0 2
rlabel polysilicon 1031 -2541 1031 -2541 0 1
rlabel polysilicon 1031 -2547 1031 -2547 0 3
rlabel polysilicon 1038 -2541 1038 -2541 0 1
rlabel polysilicon 1038 -2547 1038 -2547 0 3
rlabel polysilicon 1045 -2541 1045 -2541 0 1
rlabel polysilicon 1045 -2547 1045 -2547 0 3
rlabel polysilicon 1052 -2541 1052 -2541 0 1
rlabel polysilicon 1052 -2547 1052 -2547 0 3
rlabel polysilicon 1059 -2541 1059 -2541 0 1
rlabel polysilicon 1059 -2547 1059 -2547 0 3
rlabel polysilicon 1066 -2541 1066 -2541 0 1
rlabel polysilicon 1066 -2547 1066 -2547 0 3
rlabel polysilicon 1073 -2541 1073 -2541 0 1
rlabel polysilicon 1073 -2547 1073 -2547 0 3
rlabel polysilicon 1080 -2541 1080 -2541 0 1
rlabel polysilicon 1080 -2547 1080 -2547 0 3
rlabel polysilicon 1087 -2541 1087 -2541 0 1
rlabel polysilicon 1087 -2547 1087 -2547 0 3
rlabel polysilicon 1094 -2541 1094 -2541 0 1
rlabel polysilicon 1094 -2547 1094 -2547 0 3
rlabel polysilicon 1101 -2541 1101 -2541 0 1
rlabel polysilicon 1101 -2547 1101 -2547 0 3
rlabel polysilicon 1108 -2541 1108 -2541 0 1
rlabel polysilicon 1108 -2547 1108 -2547 0 3
rlabel polysilicon 1115 -2541 1115 -2541 0 1
rlabel polysilicon 1115 -2547 1115 -2547 0 3
rlabel polysilicon 1122 -2541 1122 -2541 0 1
rlabel polysilicon 1122 -2547 1122 -2547 0 3
rlabel polysilicon 1129 -2541 1129 -2541 0 1
rlabel polysilicon 1129 -2547 1129 -2547 0 3
rlabel polysilicon 1136 -2541 1136 -2541 0 1
rlabel polysilicon 1136 -2547 1136 -2547 0 3
rlabel polysilicon 1146 -2541 1146 -2541 0 2
rlabel polysilicon 1143 -2547 1143 -2547 0 3
rlabel polysilicon 1146 -2547 1146 -2547 0 4
rlabel polysilicon 1150 -2541 1150 -2541 0 1
rlabel polysilicon 1150 -2547 1150 -2547 0 3
rlabel polysilicon 1157 -2541 1157 -2541 0 1
rlabel polysilicon 1157 -2547 1157 -2547 0 3
rlabel polysilicon 1164 -2541 1164 -2541 0 1
rlabel polysilicon 1164 -2547 1164 -2547 0 3
rlabel polysilicon 1171 -2541 1171 -2541 0 1
rlabel polysilicon 1171 -2547 1171 -2547 0 3
rlabel polysilicon 1178 -2541 1178 -2541 0 1
rlabel polysilicon 1178 -2547 1178 -2547 0 3
rlabel polysilicon 1185 -2541 1185 -2541 0 1
rlabel polysilicon 1185 -2547 1185 -2547 0 3
rlabel polysilicon 1192 -2541 1192 -2541 0 1
rlabel polysilicon 1192 -2547 1192 -2547 0 3
rlabel polysilicon 1199 -2541 1199 -2541 0 1
rlabel polysilicon 1199 -2547 1199 -2547 0 3
rlabel polysilicon 1206 -2541 1206 -2541 0 1
rlabel polysilicon 1206 -2547 1206 -2547 0 3
rlabel polysilicon 1213 -2541 1213 -2541 0 1
rlabel polysilicon 1213 -2547 1213 -2547 0 3
rlabel polysilicon 1220 -2541 1220 -2541 0 1
rlabel polysilicon 1220 -2547 1220 -2547 0 3
rlabel polysilicon 1227 -2541 1227 -2541 0 1
rlabel polysilicon 1227 -2547 1227 -2547 0 3
rlabel polysilicon 1234 -2541 1234 -2541 0 1
rlabel polysilicon 1234 -2547 1234 -2547 0 3
rlabel polysilicon 1241 -2541 1241 -2541 0 1
rlabel polysilicon 1241 -2547 1241 -2547 0 3
rlabel polysilicon 1248 -2541 1248 -2541 0 1
rlabel polysilicon 1251 -2541 1251 -2541 0 2
rlabel polysilicon 1248 -2547 1248 -2547 0 3
rlabel polysilicon 1251 -2547 1251 -2547 0 4
rlabel polysilicon 1255 -2541 1255 -2541 0 1
rlabel polysilicon 1255 -2547 1255 -2547 0 3
rlabel polysilicon 1262 -2541 1262 -2541 0 1
rlabel polysilicon 1262 -2547 1262 -2547 0 3
rlabel polysilicon 1269 -2541 1269 -2541 0 1
rlabel polysilicon 1269 -2547 1269 -2547 0 3
rlabel polysilicon 1276 -2541 1276 -2541 0 1
rlabel polysilicon 1276 -2547 1276 -2547 0 3
rlabel polysilicon 1283 -2541 1283 -2541 0 1
rlabel polysilicon 1283 -2547 1283 -2547 0 3
rlabel polysilicon 1290 -2541 1290 -2541 0 1
rlabel polysilicon 1290 -2547 1290 -2547 0 3
rlabel polysilicon 1297 -2541 1297 -2541 0 1
rlabel polysilicon 1297 -2547 1297 -2547 0 3
rlabel polysilicon 1304 -2541 1304 -2541 0 1
rlabel polysilicon 1304 -2547 1304 -2547 0 3
rlabel polysilicon 1311 -2541 1311 -2541 0 1
rlabel polysilicon 1311 -2547 1311 -2547 0 3
rlabel polysilicon 1318 -2541 1318 -2541 0 1
rlabel polysilicon 1318 -2547 1318 -2547 0 3
rlabel polysilicon 1325 -2541 1325 -2541 0 1
rlabel polysilicon 1325 -2547 1325 -2547 0 3
rlabel polysilicon 1332 -2541 1332 -2541 0 1
rlabel polysilicon 1332 -2547 1332 -2547 0 3
rlabel polysilicon 1339 -2541 1339 -2541 0 1
rlabel polysilicon 1339 -2547 1339 -2547 0 3
rlabel polysilicon 1346 -2541 1346 -2541 0 1
rlabel polysilicon 1346 -2547 1346 -2547 0 3
rlabel polysilicon 1353 -2541 1353 -2541 0 1
rlabel polysilicon 1353 -2547 1353 -2547 0 3
rlabel polysilicon 1360 -2541 1360 -2541 0 1
rlabel polysilicon 1360 -2547 1360 -2547 0 3
rlabel polysilicon 1367 -2541 1367 -2541 0 1
rlabel polysilicon 1367 -2547 1367 -2547 0 3
rlabel polysilicon 1374 -2541 1374 -2541 0 1
rlabel polysilicon 1374 -2547 1374 -2547 0 3
rlabel polysilicon 1381 -2541 1381 -2541 0 1
rlabel polysilicon 1381 -2547 1381 -2547 0 3
rlabel polysilicon 1388 -2541 1388 -2541 0 1
rlabel polysilicon 1388 -2547 1388 -2547 0 3
rlabel polysilicon 1395 -2541 1395 -2541 0 1
rlabel polysilicon 1395 -2547 1395 -2547 0 3
rlabel polysilicon 1405 -2541 1405 -2541 0 2
rlabel polysilicon 1405 -2547 1405 -2547 0 4
rlabel polysilicon 1409 -2541 1409 -2541 0 1
rlabel polysilicon 1409 -2547 1409 -2547 0 3
rlabel polysilicon 1416 -2541 1416 -2541 0 1
rlabel polysilicon 1416 -2547 1416 -2547 0 3
rlabel polysilicon 1423 -2541 1423 -2541 0 1
rlabel polysilicon 1423 -2547 1423 -2547 0 3
rlabel polysilicon 1430 -2541 1430 -2541 0 1
rlabel polysilicon 1430 -2547 1430 -2547 0 3
rlabel polysilicon 1437 -2541 1437 -2541 0 1
rlabel polysilicon 1437 -2547 1437 -2547 0 3
rlabel polysilicon 1444 -2541 1444 -2541 0 1
rlabel polysilicon 1444 -2547 1444 -2547 0 3
rlabel polysilicon 1451 -2541 1451 -2541 0 1
rlabel polysilicon 1451 -2547 1451 -2547 0 3
rlabel polysilicon 1458 -2541 1458 -2541 0 1
rlabel polysilicon 1458 -2547 1458 -2547 0 3
rlabel polysilicon 1465 -2541 1465 -2541 0 1
rlabel polysilicon 1465 -2547 1465 -2547 0 3
rlabel polysilicon 1472 -2541 1472 -2541 0 1
rlabel polysilicon 1472 -2547 1472 -2547 0 3
rlabel polysilicon 1479 -2541 1479 -2541 0 1
rlabel polysilicon 1479 -2547 1479 -2547 0 3
rlabel polysilicon 1486 -2541 1486 -2541 0 1
rlabel polysilicon 1486 -2547 1486 -2547 0 3
rlabel polysilicon 1493 -2541 1493 -2541 0 1
rlabel polysilicon 1493 -2547 1493 -2547 0 3
rlabel polysilicon 1500 -2541 1500 -2541 0 1
rlabel polysilicon 1500 -2547 1500 -2547 0 3
rlabel polysilicon 1507 -2541 1507 -2541 0 1
rlabel polysilicon 1507 -2547 1507 -2547 0 3
rlabel polysilicon 1514 -2541 1514 -2541 0 1
rlabel polysilicon 1514 -2547 1514 -2547 0 3
rlabel polysilicon 1521 -2541 1521 -2541 0 1
rlabel polysilicon 1521 -2547 1521 -2547 0 3
rlabel polysilicon 1528 -2541 1528 -2541 0 1
rlabel polysilicon 1528 -2547 1528 -2547 0 3
rlabel polysilicon 1535 -2541 1535 -2541 0 1
rlabel polysilicon 1535 -2547 1535 -2547 0 3
rlabel polysilicon 1542 -2541 1542 -2541 0 1
rlabel polysilicon 1542 -2547 1542 -2547 0 3
rlabel polysilicon 1549 -2541 1549 -2541 0 1
rlabel polysilicon 1549 -2547 1549 -2547 0 3
rlabel polysilicon 1556 -2541 1556 -2541 0 1
rlabel polysilicon 1556 -2547 1556 -2547 0 3
rlabel polysilicon 1563 -2541 1563 -2541 0 1
rlabel polysilicon 1563 -2547 1563 -2547 0 3
rlabel polysilicon 1570 -2541 1570 -2541 0 1
rlabel polysilicon 1570 -2547 1570 -2547 0 3
rlabel polysilicon 1577 -2541 1577 -2541 0 1
rlabel polysilicon 1577 -2547 1577 -2547 0 3
rlabel polysilicon 1587 -2541 1587 -2541 0 2
rlabel polysilicon 1584 -2547 1584 -2547 0 3
rlabel polysilicon 1587 -2547 1587 -2547 0 4
rlabel polysilicon 1591 -2541 1591 -2541 0 1
rlabel polysilicon 1591 -2547 1591 -2547 0 3
rlabel polysilicon 1598 -2541 1598 -2541 0 1
rlabel polysilicon 1598 -2547 1598 -2547 0 3
rlabel polysilicon 1605 -2541 1605 -2541 0 1
rlabel polysilicon 1605 -2547 1605 -2547 0 3
rlabel polysilicon 1612 -2541 1612 -2541 0 1
rlabel polysilicon 1615 -2541 1615 -2541 0 2
rlabel polysilicon 1612 -2547 1612 -2547 0 3
rlabel polysilicon 1615 -2547 1615 -2547 0 4
rlabel polysilicon 1640 -2541 1640 -2541 0 1
rlabel polysilicon 1640 -2547 1640 -2547 0 3
rlabel polysilicon 44 -2670 44 -2670 0 1
rlabel polysilicon 44 -2676 44 -2676 0 3
rlabel polysilicon 51 -2670 51 -2670 0 1
rlabel polysilicon 51 -2676 51 -2676 0 3
rlabel polysilicon 58 -2670 58 -2670 0 1
rlabel polysilicon 58 -2676 58 -2676 0 3
rlabel polysilicon 65 -2670 65 -2670 0 1
rlabel polysilicon 65 -2676 65 -2676 0 3
rlabel polysilicon 72 -2670 72 -2670 0 1
rlabel polysilicon 72 -2676 72 -2676 0 3
rlabel polysilicon 79 -2670 79 -2670 0 1
rlabel polysilicon 79 -2676 79 -2676 0 3
rlabel polysilicon 86 -2670 86 -2670 0 1
rlabel polysilicon 86 -2676 86 -2676 0 3
rlabel polysilicon 93 -2670 93 -2670 0 1
rlabel polysilicon 93 -2676 93 -2676 0 3
rlabel polysilicon 100 -2670 100 -2670 0 1
rlabel polysilicon 100 -2676 100 -2676 0 3
rlabel polysilicon 107 -2670 107 -2670 0 1
rlabel polysilicon 107 -2676 107 -2676 0 3
rlabel polysilicon 114 -2670 114 -2670 0 1
rlabel polysilicon 114 -2676 114 -2676 0 3
rlabel polysilicon 121 -2670 121 -2670 0 1
rlabel polysilicon 121 -2676 121 -2676 0 3
rlabel polysilicon 131 -2670 131 -2670 0 2
rlabel polysilicon 128 -2676 128 -2676 0 3
rlabel polysilicon 131 -2676 131 -2676 0 4
rlabel polysilicon 135 -2670 135 -2670 0 1
rlabel polysilicon 135 -2676 135 -2676 0 3
rlabel polysilicon 142 -2670 142 -2670 0 1
rlabel polysilicon 142 -2676 142 -2676 0 3
rlabel polysilicon 149 -2670 149 -2670 0 1
rlabel polysilicon 152 -2670 152 -2670 0 2
rlabel polysilicon 149 -2676 149 -2676 0 3
rlabel polysilicon 152 -2676 152 -2676 0 4
rlabel polysilicon 156 -2670 156 -2670 0 1
rlabel polysilicon 156 -2676 156 -2676 0 3
rlabel polysilicon 163 -2670 163 -2670 0 1
rlabel polysilicon 163 -2676 163 -2676 0 3
rlabel polysilicon 170 -2670 170 -2670 0 1
rlabel polysilicon 170 -2676 170 -2676 0 3
rlabel polysilicon 180 -2670 180 -2670 0 2
rlabel polysilicon 177 -2676 177 -2676 0 3
rlabel polysilicon 184 -2670 184 -2670 0 1
rlabel polysilicon 184 -2676 184 -2676 0 3
rlabel polysilicon 191 -2670 191 -2670 0 1
rlabel polysilicon 191 -2676 191 -2676 0 3
rlabel polysilicon 201 -2670 201 -2670 0 2
rlabel polysilicon 198 -2676 198 -2676 0 3
rlabel polysilicon 201 -2676 201 -2676 0 4
rlabel polysilicon 205 -2670 205 -2670 0 1
rlabel polysilicon 208 -2670 208 -2670 0 2
rlabel polysilicon 205 -2676 205 -2676 0 3
rlabel polysilicon 208 -2676 208 -2676 0 4
rlabel polysilicon 212 -2670 212 -2670 0 1
rlabel polysilicon 212 -2676 212 -2676 0 3
rlabel polysilicon 219 -2670 219 -2670 0 1
rlabel polysilicon 219 -2676 219 -2676 0 3
rlabel polysilicon 226 -2670 226 -2670 0 1
rlabel polysilicon 226 -2676 226 -2676 0 3
rlabel polysilicon 233 -2670 233 -2670 0 1
rlabel polysilicon 236 -2670 236 -2670 0 2
rlabel polysilicon 233 -2676 233 -2676 0 3
rlabel polysilicon 236 -2676 236 -2676 0 4
rlabel polysilicon 240 -2670 240 -2670 0 1
rlabel polysilicon 240 -2676 240 -2676 0 3
rlabel polysilicon 247 -2670 247 -2670 0 1
rlabel polysilicon 247 -2676 247 -2676 0 3
rlabel polysilicon 254 -2670 254 -2670 0 1
rlabel polysilicon 254 -2676 254 -2676 0 3
rlabel polysilicon 261 -2670 261 -2670 0 1
rlabel polysilicon 264 -2670 264 -2670 0 2
rlabel polysilicon 264 -2676 264 -2676 0 4
rlabel polysilicon 268 -2670 268 -2670 0 1
rlabel polysilicon 268 -2676 268 -2676 0 3
rlabel polysilicon 275 -2670 275 -2670 0 1
rlabel polysilicon 275 -2676 275 -2676 0 3
rlabel polysilicon 282 -2670 282 -2670 0 1
rlabel polysilicon 282 -2676 282 -2676 0 3
rlabel polysilicon 289 -2670 289 -2670 0 1
rlabel polysilicon 289 -2676 289 -2676 0 3
rlabel polysilicon 296 -2670 296 -2670 0 1
rlabel polysilicon 296 -2676 296 -2676 0 3
rlabel polysilicon 303 -2670 303 -2670 0 1
rlabel polysilicon 303 -2676 303 -2676 0 3
rlabel polysilicon 310 -2670 310 -2670 0 1
rlabel polysilicon 310 -2676 310 -2676 0 3
rlabel polysilicon 317 -2670 317 -2670 0 1
rlabel polysilicon 317 -2676 317 -2676 0 3
rlabel polysilicon 324 -2670 324 -2670 0 1
rlabel polysilicon 324 -2676 324 -2676 0 3
rlabel polysilicon 331 -2670 331 -2670 0 1
rlabel polysilicon 331 -2676 331 -2676 0 3
rlabel polysilicon 338 -2670 338 -2670 0 1
rlabel polysilicon 338 -2676 338 -2676 0 3
rlabel polysilicon 345 -2670 345 -2670 0 1
rlabel polysilicon 345 -2676 345 -2676 0 3
rlabel polysilicon 352 -2670 352 -2670 0 1
rlabel polysilicon 352 -2676 352 -2676 0 3
rlabel polysilicon 359 -2670 359 -2670 0 1
rlabel polysilicon 359 -2676 359 -2676 0 3
rlabel polysilicon 366 -2670 366 -2670 0 1
rlabel polysilicon 366 -2676 366 -2676 0 3
rlabel polysilicon 376 -2670 376 -2670 0 2
rlabel polysilicon 373 -2676 373 -2676 0 3
rlabel polysilicon 380 -2670 380 -2670 0 1
rlabel polysilicon 380 -2676 380 -2676 0 3
rlabel polysilicon 387 -2670 387 -2670 0 1
rlabel polysilicon 387 -2676 387 -2676 0 3
rlabel polysilicon 394 -2676 394 -2676 0 3
rlabel polysilicon 397 -2676 397 -2676 0 4
rlabel polysilicon 401 -2670 401 -2670 0 1
rlabel polysilicon 401 -2676 401 -2676 0 3
rlabel polysilicon 408 -2670 408 -2670 0 1
rlabel polysilicon 408 -2676 408 -2676 0 3
rlabel polysilicon 415 -2670 415 -2670 0 1
rlabel polysilicon 415 -2676 415 -2676 0 3
rlabel polysilicon 422 -2670 422 -2670 0 1
rlabel polysilicon 425 -2670 425 -2670 0 2
rlabel polysilicon 422 -2676 422 -2676 0 3
rlabel polysilicon 425 -2676 425 -2676 0 4
rlabel polysilicon 429 -2670 429 -2670 0 1
rlabel polysilicon 429 -2676 429 -2676 0 3
rlabel polysilicon 436 -2670 436 -2670 0 1
rlabel polysilicon 436 -2676 436 -2676 0 3
rlabel polysilicon 443 -2670 443 -2670 0 1
rlabel polysilicon 443 -2676 443 -2676 0 3
rlabel polysilicon 450 -2670 450 -2670 0 1
rlabel polysilicon 450 -2676 450 -2676 0 3
rlabel polysilicon 457 -2670 457 -2670 0 1
rlabel polysilicon 457 -2676 457 -2676 0 3
rlabel polysilicon 464 -2670 464 -2670 0 1
rlabel polysilicon 464 -2676 464 -2676 0 3
rlabel polysilicon 471 -2670 471 -2670 0 1
rlabel polysilicon 471 -2676 471 -2676 0 3
rlabel polysilicon 478 -2670 478 -2670 0 1
rlabel polysilicon 478 -2676 478 -2676 0 3
rlabel polysilicon 485 -2670 485 -2670 0 1
rlabel polysilicon 485 -2676 485 -2676 0 3
rlabel polysilicon 492 -2670 492 -2670 0 1
rlabel polysilicon 492 -2676 492 -2676 0 3
rlabel polysilicon 499 -2670 499 -2670 0 1
rlabel polysilicon 502 -2670 502 -2670 0 2
rlabel polysilicon 499 -2676 499 -2676 0 3
rlabel polysilicon 506 -2670 506 -2670 0 1
rlabel polysilicon 506 -2676 506 -2676 0 3
rlabel polysilicon 513 -2670 513 -2670 0 1
rlabel polysilicon 513 -2676 513 -2676 0 3
rlabel polysilicon 520 -2670 520 -2670 0 1
rlabel polysilicon 520 -2676 520 -2676 0 3
rlabel polysilicon 527 -2670 527 -2670 0 1
rlabel polysilicon 527 -2676 527 -2676 0 3
rlabel polysilicon 534 -2670 534 -2670 0 1
rlabel polysilicon 534 -2676 534 -2676 0 3
rlabel polysilicon 541 -2670 541 -2670 0 1
rlabel polysilicon 541 -2676 541 -2676 0 3
rlabel polysilicon 548 -2670 548 -2670 0 1
rlabel polysilicon 548 -2676 548 -2676 0 3
rlabel polysilicon 555 -2670 555 -2670 0 1
rlabel polysilicon 555 -2676 555 -2676 0 3
rlabel polysilicon 562 -2670 562 -2670 0 1
rlabel polysilicon 562 -2676 562 -2676 0 3
rlabel polysilicon 569 -2670 569 -2670 0 1
rlabel polysilicon 569 -2676 569 -2676 0 3
rlabel polysilicon 576 -2670 576 -2670 0 1
rlabel polysilicon 576 -2676 576 -2676 0 3
rlabel polysilicon 583 -2670 583 -2670 0 1
rlabel polysilicon 583 -2676 583 -2676 0 3
rlabel polysilicon 590 -2670 590 -2670 0 1
rlabel polysilicon 590 -2676 590 -2676 0 3
rlabel polysilicon 597 -2670 597 -2670 0 1
rlabel polysilicon 597 -2676 597 -2676 0 3
rlabel polysilicon 604 -2670 604 -2670 0 1
rlabel polysilicon 604 -2676 604 -2676 0 3
rlabel polysilicon 611 -2670 611 -2670 0 1
rlabel polysilicon 614 -2670 614 -2670 0 2
rlabel polysilicon 611 -2676 611 -2676 0 3
rlabel polysilicon 614 -2676 614 -2676 0 4
rlabel polysilicon 618 -2670 618 -2670 0 1
rlabel polysilicon 618 -2676 618 -2676 0 3
rlabel polysilicon 625 -2670 625 -2670 0 1
rlabel polysilicon 625 -2676 625 -2676 0 3
rlabel polysilicon 632 -2670 632 -2670 0 1
rlabel polysilicon 632 -2676 632 -2676 0 3
rlabel polysilicon 639 -2670 639 -2670 0 1
rlabel polysilicon 639 -2676 639 -2676 0 3
rlabel polysilicon 646 -2670 646 -2670 0 1
rlabel polysilicon 649 -2676 649 -2676 0 4
rlabel polysilicon 653 -2670 653 -2670 0 1
rlabel polysilicon 656 -2670 656 -2670 0 2
rlabel polysilicon 653 -2676 653 -2676 0 3
rlabel polysilicon 656 -2676 656 -2676 0 4
rlabel polysilicon 660 -2670 660 -2670 0 1
rlabel polysilicon 660 -2676 660 -2676 0 3
rlabel polysilicon 667 -2670 667 -2670 0 1
rlabel polysilicon 667 -2676 667 -2676 0 3
rlabel polysilicon 674 -2670 674 -2670 0 1
rlabel polysilicon 674 -2676 674 -2676 0 3
rlabel polysilicon 681 -2670 681 -2670 0 1
rlabel polysilicon 681 -2676 681 -2676 0 3
rlabel polysilicon 688 -2670 688 -2670 0 1
rlabel polysilicon 688 -2676 688 -2676 0 3
rlabel polysilicon 695 -2670 695 -2670 0 1
rlabel polysilicon 695 -2676 695 -2676 0 3
rlabel polysilicon 702 -2670 702 -2670 0 1
rlabel polysilicon 702 -2676 702 -2676 0 3
rlabel polysilicon 709 -2670 709 -2670 0 1
rlabel polysilicon 709 -2676 709 -2676 0 3
rlabel polysilicon 719 -2670 719 -2670 0 2
rlabel polysilicon 723 -2670 723 -2670 0 1
rlabel polysilicon 723 -2676 723 -2676 0 3
rlabel polysilicon 730 -2670 730 -2670 0 1
rlabel polysilicon 733 -2670 733 -2670 0 2
rlabel polysilicon 733 -2676 733 -2676 0 4
rlabel polysilicon 737 -2670 737 -2670 0 1
rlabel polysilicon 737 -2676 737 -2676 0 3
rlabel polysilicon 744 -2670 744 -2670 0 1
rlabel polysilicon 744 -2676 744 -2676 0 3
rlabel polysilicon 751 -2670 751 -2670 0 1
rlabel polysilicon 751 -2676 751 -2676 0 3
rlabel polysilicon 758 -2670 758 -2670 0 1
rlabel polysilicon 758 -2676 758 -2676 0 3
rlabel polysilicon 765 -2670 765 -2670 0 1
rlabel polysilicon 765 -2676 765 -2676 0 3
rlabel polysilicon 772 -2670 772 -2670 0 1
rlabel polysilicon 772 -2676 772 -2676 0 3
rlabel polysilicon 779 -2670 779 -2670 0 1
rlabel polysilicon 779 -2676 779 -2676 0 3
rlabel polysilicon 786 -2670 786 -2670 0 1
rlabel polysilicon 786 -2676 786 -2676 0 3
rlabel polysilicon 793 -2670 793 -2670 0 1
rlabel polysilicon 793 -2676 793 -2676 0 3
rlabel polysilicon 803 -2670 803 -2670 0 2
rlabel polysilicon 800 -2676 800 -2676 0 3
rlabel polysilicon 803 -2676 803 -2676 0 4
rlabel polysilicon 807 -2670 807 -2670 0 1
rlabel polysilicon 807 -2676 807 -2676 0 3
rlabel polysilicon 814 -2670 814 -2670 0 1
rlabel polysilicon 814 -2676 814 -2676 0 3
rlabel polysilicon 821 -2670 821 -2670 0 1
rlabel polysilicon 821 -2676 821 -2676 0 3
rlabel polysilicon 828 -2670 828 -2670 0 1
rlabel polysilicon 828 -2676 828 -2676 0 3
rlabel polysilicon 835 -2670 835 -2670 0 1
rlabel polysilicon 835 -2676 835 -2676 0 3
rlabel polysilicon 842 -2670 842 -2670 0 1
rlabel polysilicon 842 -2676 842 -2676 0 3
rlabel polysilicon 849 -2670 849 -2670 0 1
rlabel polysilicon 849 -2676 849 -2676 0 3
rlabel polysilicon 859 -2670 859 -2670 0 2
rlabel polysilicon 856 -2676 856 -2676 0 3
rlabel polysilicon 859 -2676 859 -2676 0 4
rlabel polysilicon 863 -2670 863 -2670 0 1
rlabel polysilicon 863 -2676 863 -2676 0 3
rlabel polysilicon 870 -2670 870 -2670 0 1
rlabel polysilicon 870 -2676 870 -2676 0 3
rlabel polysilicon 877 -2670 877 -2670 0 1
rlabel polysilicon 880 -2670 880 -2670 0 2
rlabel polysilicon 877 -2676 877 -2676 0 3
rlabel polysilicon 880 -2676 880 -2676 0 4
rlabel polysilicon 884 -2670 884 -2670 0 1
rlabel polysilicon 887 -2670 887 -2670 0 2
rlabel polysilicon 884 -2676 884 -2676 0 3
rlabel polysilicon 887 -2676 887 -2676 0 4
rlabel polysilicon 891 -2670 891 -2670 0 1
rlabel polysilicon 891 -2676 891 -2676 0 3
rlabel polysilicon 898 -2670 898 -2670 0 1
rlabel polysilicon 901 -2670 901 -2670 0 2
rlabel polysilicon 898 -2676 898 -2676 0 3
rlabel polysilicon 901 -2676 901 -2676 0 4
rlabel polysilicon 905 -2670 905 -2670 0 1
rlabel polysilicon 905 -2676 905 -2676 0 3
rlabel polysilicon 912 -2670 912 -2670 0 1
rlabel polysilicon 912 -2676 912 -2676 0 3
rlabel polysilicon 919 -2670 919 -2670 0 1
rlabel polysilicon 919 -2676 919 -2676 0 3
rlabel polysilicon 926 -2670 926 -2670 0 1
rlabel polysilicon 926 -2676 926 -2676 0 3
rlabel polysilicon 933 -2670 933 -2670 0 1
rlabel polysilicon 933 -2676 933 -2676 0 3
rlabel polysilicon 940 -2670 940 -2670 0 1
rlabel polysilicon 940 -2676 940 -2676 0 3
rlabel polysilicon 947 -2670 947 -2670 0 1
rlabel polysilicon 950 -2670 950 -2670 0 2
rlabel polysilicon 947 -2676 947 -2676 0 3
rlabel polysilicon 950 -2676 950 -2676 0 4
rlabel polysilicon 954 -2670 954 -2670 0 1
rlabel polysilicon 957 -2670 957 -2670 0 2
rlabel polysilicon 954 -2676 954 -2676 0 3
rlabel polysilicon 957 -2676 957 -2676 0 4
rlabel polysilicon 961 -2670 961 -2670 0 1
rlabel polysilicon 961 -2676 961 -2676 0 3
rlabel polysilicon 968 -2670 968 -2670 0 1
rlabel polysilicon 971 -2670 971 -2670 0 2
rlabel polysilicon 971 -2676 971 -2676 0 4
rlabel polysilicon 975 -2670 975 -2670 0 1
rlabel polysilicon 978 -2670 978 -2670 0 2
rlabel polysilicon 975 -2676 975 -2676 0 3
rlabel polysilicon 978 -2676 978 -2676 0 4
rlabel polysilicon 982 -2670 982 -2670 0 1
rlabel polysilicon 982 -2676 982 -2676 0 3
rlabel polysilicon 989 -2670 989 -2670 0 1
rlabel polysilicon 989 -2676 989 -2676 0 3
rlabel polysilicon 996 -2670 996 -2670 0 1
rlabel polysilicon 996 -2676 996 -2676 0 3
rlabel polysilicon 1003 -2670 1003 -2670 0 1
rlabel polysilicon 1003 -2676 1003 -2676 0 3
rlabel polysilicon 1010 -2670 1010 -2670 0 1
rlabel polysilicon 1010 -2676 1010 -2676 0 3
rlabel polysilicon 1017 -2670 1017 -2670 0 1
rlabel polysilicon 1017 -2676 1017 -2676 0 3
rlabel polysilicon 1024 -2670 1024 -2670 0 1
rlabel polysilicon 1027 -2670 1027 -2670 0 2
rlabel polysilicon 1024 -2676 1024 -2676 0 3
rlabel polysilicon 1031 -2670 1031 -2670 0 1
rlabel polysilicon 1031 -2676 1031 -2676 0 3
rlabel polysilicon 1038 -2670 1038 -2670 0 1
rlabel polysilicon 1038 -2676 1038 -2676 0 3
rlabel polysilicon 1045 -2670 1045 -2670 0 1
rlabel polysilicon 1045 -2676 1045 -2676 0 3
rlabel polysilicon 1052 -2670 1052 -2670 0 1
rlabel polysilicon 1052 -2676 1052 -2676 0 3
rlabel polysilicon 1059 -2670 1059 -2670 0 1
rlabel polysilicon 1059 -2676 1059 -2676 0 3
rlabel polysilicon 1066 -2670 1066 -2670 0 1
rlabel polysilicon 1066 -2676 1066 -2676 0 3
rlabel polysilicon 1073 -2670 1073 -2670 0 1
rlabel polysilicon 1073 -2676 1073 -2676 0 3
rlabel polysilicon 1080 -2670 1080 -2670 0 1
rlabel polysilicon 1080 -2676 1080 -2676 0 3
rlabel polysilicon 1087 -2670 1087 -2670 0 1
rlabel polysilicon 1090 -2670 1090 -2670 0 2
rlabel polysilicon 1090 -2676 1090 -2676 0 4
rlabel polysilicon 1094 -2670 1094 -2670 0 1
rlabel polysilicon 1094 -2676 1094 -2676 0 3
rlabel polysilicon 1101 -2670 1101 -2670 0 1
rlabel polysilicon 1101 -2676 1101 -2676 0 3
rlabel polysilicon 1108 -2670 1108 -2670 0 1
rlabel polysilicon 1108 -2676 1108 -2676 0 3
rlabel polysilicon 1115 -2670 1115 -2670 0 1
rlabel polysilicon 1115 -2676 1115 -2676 0 3
rlabel polysilicon 1122 -2670 1122 -2670 0 1
rlabel polysilicon 1122 -2676 1122 -2676 0 3
rlabel polysilicon 1129 -2670 1129 -2670 0 1
rlabel polysilicon 1129 -2676 1129 -2676 0 3
rlabel polysilicon 1136 -2670 1136 -2670 0 1
rlabel polysilicon 1136 -2676 1136 -2676 0 3
rlabel polysilicon 1143 -2670 1143 -2670 0 1
rlabel polysilicon 1143 -2676 1143 -2676 0 3
rlabel polysilicon 1150 -2670 1150 -2670 0 1
rlabel polysilicon 1153 -2670 1153 -2670 0 2
rlabel polysilicon 1150 -2676 1150 -2676 0 3
rlabel polysilicon 1153 -2676 1153 -2676 0 4
rlabel polysilicon 1157 -2670 1157 -2670 0 1
rlabel polysilicon 1157 -2676 1157 -2676 0 3
rlabel polysilicon 1164 -2670 1164 -2670 0 1
rlabel polysilicon 1164 -2676 1164 -2676 0 3
rlabel polysilicon 1171 -2670 1171 -2670 0 1
rlabel polysilicon 1171 -2676 1171 -2676 0 3
rlabel polysilicon 1178 -2670 1178 -2670 0 1
rlabel polysilicon 1178 -2676 1178 -2676 0 3
rlabel polysilicon 1185 -2670 1185 -2670 0 1
rlabel polysilicon 1188 -2670 1188 -2670 0 2
rlabel polysilicon 1185 -2676 1185 -2676 0 3
rlabel polysilicon 1188 -2676 1188 -2676 0 4
rlabel polysilicon 1192 -2670 1192 -2670 0 1
rlabel polysilicon 1192 -2676 1192 -2676 0 3
rlabel polysilicon 1199 -2670 1199 -2670 0 1
rlabel polysilicon 1199 -2676 1199 -2676 0 3
rlabel polysilicon 1206 -2670 1206 -2670 0 1
rlabel polysilicon 1206 -2676 1206 -2676 0 3
rlabel polysilicon 1213 -2670 1213 -2670 0 1
rlabel polysilicon 1213 -2676 1213 -2676 0 3
rlabel polysilicon 1220 -2670 1220 -2670 0 1
rlabel polysilicon 1220 -2676 1220 -2676 0 3
rlabel polysilicon 1227 -2670 1227 -2670 0 1
rlabel polysilicon 1227 -2676 1227 -2676 0 3
rlabel polysilicon 1234 -2670 1234 -2670 0 1
rlabel polysilicon 1234 -2676 1234 -2676 0 3
rlabel polysilicon 1241 -2670 1241 -2670 0 1
rlabel polysilicon 1241 -2676 1241 -2676 0 3
rlabel polysilicon 1248 -2670 1248 -2670 0 1
rlabel polysilicon 1248 -2676 1248 -2676 0 3
rlabel polysilicon 1255 -2670 1255 -2670 0 1
rlabel polysilicon 1255 -2676 1255 -2676 0 3
rlabel polysilicon 1262 -2670 1262 -2670 0 1
rlabel polysilicon 1262 -2676 1262 -2676 0 3
rlabel polysilicon 1269 -2670 1269 -2670 0 1
rlabel polysilicon 1269 -2676 1269 -2676 0 3
rlabel polysilicon 1276 -2670 1276 -2670 0 1
rlabel polysilicon 1276 -2676 1276 -2676 0 3
rlabel polysilicon 1283 -2670 1283 -2670 0 1
rlabel polysilicon 1283 -2676 1283 -2676 0 3
rlabel polysilicon 1290 -2670 1290 -2670 0 1
rlabel polysilicon 1290 -2676 1290 -2676 0 3
rlabel polysilicon 1297 -2670 1297 -2670 0 1
rlabel polysilicon 1297 -2676 1297 -2676 0 3
rlabel polysilicon 1304 -2670 1304 -2670 0 1
rlabel polysilicon 1304 -2676 1304 -2676 0 3
rlabel polysilicon 1311 -2670 1311 -2670 0 1
rlabel polysilicon 1311 -2676 1311 -2676 0 3
rlabel polysilicon 1318 -2670 1318 -2670 0 1
rlabel polysilicon 1318 -2676 1318 -2676 0 3
rlabel polysilicon 1325 -2670 1325 -2670 0 1
rlabel polysilicon 1325 -2676 1325 -2676 0 3
rlabel polysilicon 1332 -2670 1332 -2670 0 1
rlabel polysilicon 1332 -2676 1332 -2676 0 3
rlabel polysilicon 1339 -2670 1339 -2670 0 1
rlabel polysilicon 1339 -2676 1339 -2676 0 3
rlabel polysilicon 1346 -2670 1346 -2670 0 1
rlabel polysilicon 1346 -2676 1346 -2676 0 3
rlabel polysilicon 1353 -2670 1353 -2670 0 1
rlabel polysilicon 1353 -2676 1353 -2676 0 3
rlabel polysilicon 1360 -2670 1360 -2670 0 1
rlabel polysilicon 1360 -2676 1360 -2676 0 3
rlabel polysilicon 1367 -2670 1367 -2670 0 1
rlabel polysilicon 1367 -2676 1367 -2676 0 3
rlabel polysilicon 1374 -2670 1374 -2670 0 1
rlabel polysilicon 1374 -2676 1374 -2676 0 3
rlabel polysilicon 1381 -2670 1381 -2670 0 1
rlabel polysilicon 1381 -2676 1381 -2676 0 3
rlabel polysilicon 1388 -2670 1388 -2670 0 1
rlabel polysilicon 1388 -2676 1388 -2676 0 3
rlabel polysilicon 1395 -2670 1395 -2670 0 1
rlabel polysilicon 1395 -2676 1395 -2676 0 3
rlabel polysilicon 1402 -2670 1402 -2670 0 1
rlabel polysilicon 1402 -2676 1402 -2676 0 3
rlabel polysilicon 1409 -2670 1409 -2670 0 1
rlabel polysilicon 1409 -2676 1409 -2676 0 3
rlabel polysilicon 1416 -2670 1416 -2670 0 1
rlabel polysilicon 1416 -2676 1416 -2676 0 3
rlabel polysilicon 1423 -2670 1423 -2670 0 1
rlabel polysilicon 1423 -2676 1423 -2676 0 3
rlabel polysilicon 1430 -2670 1430 -2670 0 1
rlabel polysilicon 1430 -2676 1430 -2676 0 3
rlabel polysilicon 1437 -2670 1437 -2670 0 1
rlabel polysilicon 1437 -2676 1437 -2676 0 3
rlabel polysilicon 1444 -2670 1444 -2670 0 1
rlabel polysilicon 1444 -2676 1444 -2676 0 3
rlabel polysilicon 1451 -2670 1451 -2670 0 1
rlabel polysilicon 1451 -2676 1451 -2676 0 3
rlabel polysilicon 1458 -2670 1458 -2670 0 1
rlabel polysilicon 1458 -2676 1458 -2676 0 3
rlabel polysilicon 1465 -2670 1465 -2670 0 1
rlabel polysilicon 1465 -2676 1465 -2676 0 3
rlabel polysilicon 1472 -2670 1472 -2670 0 1
rlabel polysilicon 1472 -2676 1472 -2676 0 3
rlabel polysilicon 1479 -2670 1479 -2670 0 1
rlabel polysilicon 1479 -2676 1479 -2676 0 3
rlabel polysilicon 1486 -2670 1486 -2670 0 1
rlabel polysilicon 1486 -2676 1486 -2676 0 3
rlabel polysilicon 1493 -2670 1493 -2670 0 1
rlabel polysilicon 1493 -2676 1493 -2676 0 3
rlabel polysilicon 1500 -2670 1500 -2670 0 1
rlabel polysilicon 1500 -2676 1500 -2676 0 3
rlabel polysilicon 1507 -2670 1507 -2670 0 1
rlabel polysilicon 1507 -2676 1507 -2676 0 3
rlabel polysilicon 1514 -2670 1514 -2670 0 1
rlabel polysilicon 1514 -2676 1514 -2676 0 3
rlabel polysilicon 1521 -2670 1521 -2670 0 1
rlabel polysilicon 1521 -2676 1521 -2676 0 3
rlabel polysilicon 1528 -2670 1528 -2670 0 1
rlabel polysilicon 1528 -2676 1528 -2676 0 3
rlabel polysilicon 1535 -2670 1535 -2670 0 1
rlabel polysilicon 1535 -2676 1535 -2676 0 3
rlabel polysilicon 1542 -2670 1542 -2670 0 1
rlabel polysilicon 1542 -2676 1542 -2676 0 3
rlabel polysilicon 1549 -2670 1549 -2670 0 1
rlabel polysilicon 1549 -2676 1549 -2676 0 3
rlabel polysilicon 1556 -2670 1556 -2670 0 1
rlabel polysilicon 1556 -2676 1556 -2676 0 3
rlabel polysilicon 1563 -2670 1563 -2670 0 1
rlabel polysilicon 1563 -2676 1563 -2676 0 3
rlabel polysilicon 1570 -2670 1570 -2670 0 1
rlabel polysilicon 1570 -2676 1570 -2676 0 3
rlabel polysilicon 1577 -2670 1577 -2670 0 1
rlabel polysilicon 1577 -2676 1577 -2676 0 3
rlabel polysilicon 1584 -2670 1584 -2670 0 1
rlabel polysilicon 1584 -2676 1584 -2676 0 3
rlabel polysilicon 1591 -2670 1591 -2670 0 1
rlabel polysilicon 1591 -2676 1591 -2676 0 3
rlabel polysilicon 1598 -2670 1598 -2670 0 1
rlabel polysilicon 1598 -2676 1598 -2676 0 3
rlabel polysilicon 1605 -2670 1605 -2670 0 1
rlabel polysilicon 1605 -2676 1605 -2676 0 3
rlabel polysilicon 1612 -2670 1612 -2670 0 1
rlabel polysilicon 1612 -2676 1612 -2676 0 3
rlabel polysilicon 1619 -2670 1619 -2670 0 1
rlabel polysilicon 1619 -2676 1619 -2676 0 3
rlabel polysilicon 1626 -2670 1626 -2670 0 1
rlabel polysilicon 1629 -2670 1629 -2670 0 2
rlabel polysilicon 1626 -2676 1626 -2676 0 3
rlabel polysilicon 1629 -2676 1629 -2676 0 4
rlabel polysilicon 1636 -2670 1636 -2670 0 2
rlabel polysilicon 1633 -2676 1633 -2676 0 3
rlabel polysilicon 1636 -2676 1636 -2676 0 4
rlabel polysilicon 44 -2783 44 -2783 0 1
rlabel polysilicon 44 -2789 44 -2789 0 3
rlabel polysilicon 58 -2783 58 -2783 0 1
rlabel polysilicon 58 -2789 58 -2789 0 3
rlabel polysilicon 65 -2783 65 -2783 0 1
rlabel polysilicon 65 -2789 65 -2789 0 3
rlabel polysilicon 72 -2783 72 -2783 0 1
rlabel polysilicon 72 -2789 72 -2789 0 3
rlabel polysilicon 79 -2783 79 -2783 0 1
rlabel polysilicon 79 -2789 79 -2789 0 3
rlabel polysilicon 86 -2783 86 -2783 0 1
rlabel polysilicon 86 -2789 86 -2789 0 3
rlabel polysilicon 93 -2783 93 -2783 0 1
rlabel polysilicon 93 -2789 93 -2789 0 3
rlabel polysilicon 100 -2783 100 -2783 0 1
rlabel polysilicon 100 -2789 100 -2789 0 3
rlabel polysilicon 107 -2783 107 -2783 0 1
rlabel polysilicon 107 -2789 107 -2789 0 3
rlabel polysilicon 110 -2789 110 -2789 0 4
rlabel polysilicon 114 -2783 114 -2783 0 1
rlabel polysilicon 114 -2789 114 -2789 0 3
rlabel polysilicon 121 -2783 121 -2783 0 1
rlabel polysilicon 124 -2783 124 -2783 0 2
rlabel polysilicon 121 -2789 121 -2789 0 3
rlabel polysilicon 124 -2789 124 -2789 0 4
rlabel polysilicon 128 -2783 128 -2783 0 1
rlabel polysilicon 131 -2783 131 -2783 0 2
rlabel polysilicon 128 -2789 128 -2789 0 3
rlabel polysilicon 135 -2783 135 -2783 0 1
rlabel polysilicon 138 -2783 138 -2783 0 2
rlabel polysilicon 135 -2789 135 -2789 0 3
rlabel polysilicon 138 -2789 138 -2789 0 4
rlabel polysilicon 142 -2783 142 -2783 0 1
rlabel polysilicon 142 -2789 142 -2789 0 3
rlabel polysilicon 149 -2783 149 -2783 0 1
rlabel polysilicon 149 -2789 149 -2789 0 3
rlabel polysilicon 156 -2783 156 -2783 0 1
rlabel polysilicon 159 -2783 159 -2783 0 2
rlabel polysilicon 159 -2789 159 -2789 0 4
rlabel polysilicon 163 -2783 163 -2783 0 1
rlabel polysilicon 163 -2789 163 -2789 0 3
rlabel polysilicon 170 -2783 170 -2783 0 1
rlabel polysilicon 170 -2789 170 -2789 0 3
rlabel polysilicon 177 -2783 177 -2783 0 1
rlabel polysilicon 177 -2789 177 -2789 0 3
rlabel polysilicon 184 -2783 184 -2783 0 1
rlabel polysilicon 184 -2789 184 -2789 0 3
rlabel polysilicon 191 -2783 191 -2783 0 1
rlabel polysilicon 191 -2789 191 -2789 0 3
rlabel polysilicon 198 -2783 198 -2783 0 1
rlabel polysilicon 198 -2789 198 -2789 0 3
rlabel polysilicon 205 -2783 205 -2783 0 1
rlabel polysilicon 205 -2789 205 -2789 0 3
rlabel polysilicon 212 -2783 212 -2783 0 1
rlabel polysilicon 215 -2783 215 -2783 0 2
rlabel polysilicon 212 -2789 212 -2789 0 3
rlabel polysilicon 215 -2789 215 -2789 0 4
rlabel polysilicon 219 -2783 219 -2783 0 1
rlabel polysilicon 219 -2789 219 -2789 0 3
rlabel polysilicon 226 -2783 226 -2783 0 1
rlabel polysilicon 226 -2789 226 -2789 0 3
rlabel polysilicon 233 -2789 233 -2789 0 3
rlabel polysilicon 236 -2789 236 -2789 0 4
rlabel polysilicon 240 -2783 240 -2783 0 1
rlabel polysilicon 240 -2789 240 -2789 0 3
rlabel polysilicon 247 -2783 247 -2783 0 1
rlabel polysilicon 247 -2789 247 -2789 0 3
rlabel polysilicon 254 -2783 254 -2783 0 1
rlabel polysilicon 254 -2789 254 -2789 0 3
rlabel polysilicon 261 -2783 261 -2783 0 1
rlabel polysilicon 264 -2783 264 -2783 0 2
rlabel polysilicon 264 -2789 264 -2789 0 4
rlabel polysilicon 268 -2783 268 -2783 0 1
rlabel polysilicon 268 -2789 268 -2789 0 3
rlabel polysilicon 275 -2783 275 -2783 0 1
rlabel polysilicon 275 -2789 275 -2789 0 3
rlabel polysilicon 282 -2789 282 -2789 0 3
rlabel polysilicon 289 -2783 289 -2783 0 1
rlabel polysilicon 292 -2783 292 -2783 0 2
rlabel polysilicon 292 -2789 292 -2789 0 4
rlabel polysilicon 296 -2783 296 -2783 0 1
rlabel polysilicon 296 -2789 296 -2789 0 3
rlabel polysilicon 303 -2783 303 -2783 0 1
rlabel polysilicon 303 -2789 303 -2789 0 3
rlabel polysilicon 310 -2783 310 -2783 0 1
rlabel polysilicon 310 -2789 310 -2789 0 3
rlabel polysilicon 317 -2783 317 -2783 0 1
rlabel polysilicon 317 -2789 317 -2789 0 3
rlabel polysilicon 324 -2783 324 -2783 0 1
rlabel polysilicon 324 -2789 324 -2789 0 3
rlabel polysilicon 331 -2783 331 -2783 0 1
rlabel polysilicon 331 -2789 331 -2789 0 3
rlabel polysilicon 338 -2783 338 -2783 0 1
rlabel polysilicon 338 -2789 338 -2789 0 3
rlabel polysilicon 345 -2783 345 -2783 0 1
rlabel polysilicon 345 -2789 345 -2789 0 3
rlabel polysilicon 352 -2783 352 -2783 0 1
rlabel polysilicon 352 -2789 352 -2789 0 3
rlabel polysilicon 359 -2783 359 -2783 0 1
rlabel polysilicon 359 -2789 359 -2789 0 3
rlabel polysilicon 366 -2783 366 -2783 0 1
rlabel polysilicon 366 -2789 366 -2789 0 3
rlabel polysilicon 373 -2783 373 -2783 0 1
rlabel polysilicon 373 -2789 373 -2789 0 3
rlabel polysilicon 380 -2783 380 -2783 0 1
rlabel polysilicon 380 -2789 380 -2789 0 3
rlabel polysilicon 387 -2783 387 -2783 0 1
rlabel polysilicon 387 -2789 387 -2789 0 3
rlabel polysilicon 394 -2783 394 -2783 0 1
rlabel polysilicon 394 -2789 394 -2789 0 3
rlabel polysilicon 401 -2783 401 -2783 0 1
rlabel polysilicon 401 -2789 401 -2789 0 3
rlabel polysilicon 408 -2783 408 -2783 0 1
rlabel polysilicon 408 -2789 408 -2789 0 3
rlabel polysilicon 415 -2783 415 -2783 0 1
rlabel polysilicon 415 -2789 415 -2789 0 3
rlabel polysilicon 422 -2783 422 -2783 0 1
rlabel polysilicon 422 -2789 422 -2789 0 3
rlabel polysilicon 429 -2783 429 -2783 0 1
rlabel polysilicon 429 -2789 429 -2789 0 3
rlabel polysilicon 436 -2783 436 -2783 0 1
rlabel polysilicon 436 -2789 436 -2789 0 3
rlabel polysilicon 446 -2783 446 -2783 0 2
rlabel polysilicon 443 -2789 443 -2789 0 3
rlabel polysilicon 446 -2789 446 -2789 0 4
rlabel polysilicon 450 -2783 450 -2783 0 1
rlabel polysilicon 450 -2789 450 -2789 0 3
rlabel polysilicon 457 -2783 457 -2783 0 1
rlabel polysilicon 457 -2789 457 -2789 0 3
rlabel polysilicon 464 -2783 464 -2783 0 1
rlabel polysilicon 464 -2789 464 -2789 0 3
rlabel polysilicon 471 -2783 471 -2783 0 1
rlabel polysilicon 471 -2789 471 -2789 0 3
rlabel polysilicon 478 -2783 478 -2783 0 1
rlabel polysilicon 485 -2783 485 -2783 0 1
rlabel polysilicon 485 -2789 485 -2789 0 3
rlabel polysilicon 492 -2783 492 -2783 0 1
rlabel polysilicon 492 -2789 492 -2789 0 3
rlabel polysilicon 499 -2783 499 -2783 0 1
rlabel polysilicon 499 -2789 499 -2789 0 3
rlabel polysilicon 506 -2783 506 -2783 0 1
rlabel polysilicon 506 -2789 506 -2789 0 3
rlabel polysilicon 513 -2783 513 -2783 0 1
rlabel polysilicon 513 -2789 513 -2789 0 3
rlabel polysilicon 520 -2783 520 -2783 0 1
rlabel polysilicon 520 -2789 520 -2789 0 3
rlabel polysilicon 527 -2783 527 -2783 0 1
rlabel polysilicon 527 -2789 527 -2789 0 3
rlabel polysilicon 534 -2783 534 -2783 0 1
rlabel polysilicon 534 -2789 534 -2789 0 3
rlabel polysilicon 541 -2783 541 -2783 0 1
rlabel polysilicon 541 -2789 541 -2789 0 3
rlabel polysilicon 548 -2783 548 -2783 0 1
rlabel polysilicon 548 -2789 548 -2789 0 3
rlabel polysilicon 555 -2783 555 -2783 0 1
rlabel polysilicon 555 -2789 555 -2789 0 3
rlabel polysilicon 562 -2783 562 -2783 0 1
rlabel polysilicon 565 -2783 565 -2783 0 2
rlabel polysilicon 562 -2789 562 -2789 0 3
rlabel polysilicon 565 -2789 565 -2789 0 4
rlabel polysilicon 569 -2783 569 -2783 0 1
rlabel polysilicon 569 -2789 569 -2789 0 3
rlabel polysilicon 576 -2783 576 -2783 0 1
rlabel polysilicon 576 -2789 576 -2789 0 3
rlabel polysilicon 583 -2783 583 -2783 0 1
rlabel polysilicon 583 -2789 583 -2789 0 3
rlabel polysilicon 590 -2789 590 -2789 0 3
rlabel polysilicon 593 -2789 593 -2789 0 4
rlabel polysilicon 597 -2783 597 -2783 0 1
rlabel polysilicon 597 -2789 597 -2789 0 3
rlabel polysilicon 604 -2783 604 -2783 0 1
rlabel polysilicon 604 -2789 604 -2789 0 3
rlabel polysilicon 611 -2783 611 -2783 0 1
rlabel polysilicon 611 -2789 611 -2789 0 3
rlabel polysilicon 618 -2783 618 -2783 0 1
rlabel polysilicon 618 -2789 618 -2789 0 3
rlabel polysilicon 625 -2783 625 -2783 0 1
rlabel polysilicon 625 -2789 625 -2789 0 3
rlabel polysilicon 632 -2783 632 -2783 0 1
rlabel polysilicon 632 -2789 632 -2789 0 3
rlabel polysilicon 639 -2783 639 -2783 0 1
rlabel polysilicon 639 -2789 639 -2789 0 3
rlabel polysilicon 646 -2783 646 -2783 0 1
rlabel polysilicon 646 -2789 646 -2789 0 3
rlabel polysilicon 653 -2783 653 -2783 0 1
rlabel polysilicon 653 -2789 653 -2789 0 3
rlabel polysilicon 660 -2783 660 -2783 0 1
rlabel polysilicon 663 -2783 663 -2783 0 2
rlabel polysilicon 660 -2789 660 -2789 0 3
rlabel polysilicon 663 -2789 663 -2789 0 4
rlabel polysilicon 667 -2783 667 -2783 0 1
rlabel polysilicon 667 -2789 667 -2789 0 3
rlabel polysilicon 670 -2789 670 -2789 0 4
rlabel polysilicon 674 -2783 674 -2783 0 1
rlabel polysilicon 677 -2783 677 -2783 0 2
rlabel polysilicon 677 -2789 677 -2789 0 4
rlabel polysilicon 681 -2783 681 -2783 0 1
rlabel polysilicon 681 -2789 681 -2789 0 3
rlabel polysilicon 691 -2783 691 -2783 0 2
rlabel polysilicon 688 -2789 688 -2789 0 3
rlabel polysilicon 695 -2783 695 -2783 0 1
rlabel polysilicon 695 -2789 695 -2789 0 3
rlabel polysilicon 702 -2783 702 -2783 0 1
rlabel polysilicon 702 -2789 702 -2789 0 3
rlabel polysilicon 709 -2783 709 -2783 0 1
rlabel polysilicon 709 -2789 709 -2789 0 3
rlabel polysilicon 716 -2783 716 -2783 0 1
rlabel polysilicon 716 -2789 716 -2789 0 3
rlabel polysilicon 723 -2783 723 -2783 0 1
rlabel polysilicon 723 -2789 723 -2789 0 3
rlabel polysilicon 730 -2783 730 -2783 0 1
rlabel polysilicon 730 -2789 730 -2789 0 3
rlabel polysilicon 737 -2783 737 -2783 0 1
rlabel polysilicon 737 -2789 737 -2789 0 3
rlabel polysilicon 744 -2783 744 -2783 0 1
rlabel polysilicon 747 -2783 747 -2783 0 2
rlabel polysilicon 744 -2789 744 -2789 0 3
rlabel polysilicon 747 -2789 747 -2789 0 4
rlabel polysilicon 751 -2783 751 -2783 0 1
rlabel polysilicon 751 -2789 751 -2789 0 3
rlabel polysilicon 758 -2783 758 -2783 0 1
rlabel polysilicon 761 -2783 761 -2783 0 2
rlabel polysilicon 761 -2789 761 -2789 0 4
rlabel polysilicon 765 -2783 765 -2783 0 1
rlabel polysilicon 765 -2789 765 -2789 0 3
rlabel polysilicon 772 -2783 772 -2783 0 1
rlabel polysilicon 772 -2789 772 -2789 0 3
rlabel polysilicon 779 -2783 779 -2783 0 1
rlabel polysilicon 782 -2783 782 -2783 0 2
rlabel polysilicon 779 -2789 779 -2789 0 3
rlabel polysilicon 786 -2783 786 -2783 0 1
rlabel polysilicon 786 -2789 786 -2789 0 3
rlabel polysilicon 789 -2789 789 -2789 0 4
rlabel polysilicon 793 -2783 793 -2783 0 1
rlabel polysilicon 793 -2789 793 -2789 0 3
rlabel polysilicon 800 -2783 800 -2783 0 1
rlabel polysilicon 800 -2789 800 -2789 0 3
rlabel polysilicon 807 -2789 807 -2789 0 3
rlabel polysilicon 810 -2789 810 -2789 0 4
rlabel polysilicon 814 -2783 814 -2783 0 1
rlabel polysilicon 817 -2783 817 -2783 0 2
rlabel polysilicon 814 -2789 814 -2789 0 3
rlabel polysilicon 817 -2789 817 -2789 0 4
rlabel polysilicon 821 -2783 821 -2783 0 1
rlabel polysilicon 821 -2789 821 -2789 0 3
rlabel polysilicon 828 -2783 828 -2783 0 1
rlabel polysilicon 828 -2789 828 -2789 0 3
rlabel polysilicon 835 -2783 835 -2783 0 1
rlabel polysilicon 835 -2789 835 -2789 0 3
rlabel polysilicon 842 -2783 842 -2783 0 1
rlabel polysilicon 845 -2783 845 -2783 0 2
rlabel polysilicon 842 -2789 842 -2789 0 3
rlabel polysilicon 845 -2789 845 -2789 0 4
rlabel polysilicon 849 -2783 849 -2783 0 1
rlabel polysilicon 849 -2789 849 -2789 0 3
rlabel polysilicon 856 -2783 856 -2783 0 1
rlabel polysilicon 856 -2789 856 -2789 0 3
rlabel polysilicon 863 -2783 863 -2783 0 1
rlabel polysilicon 863 -2789 863 -2789 0 3
rlabel polysilicon 870 -2783 870 -2783 0 1
rlabel polysilicon 870 -2789 870 -2789 0 3
rlabel polysilicon 877 -2783 877 -2783 0 1
rlabel polysilicon 880 -2783 880 -2783 0 2
rlabel polysilicon 877 -2789 877 -2789 0 3
rlabel polysilicon 880 -2789 880 -2789 0 4
rlabel polysilicon 884 -2783 884 -2783 0 1
rlabel polysilicon 884 -2789 884 -2789 0 3
rlabel polysilicon 891 -2783 891 -2783 0 1
rlabel polysilicon 891 -2789 891 -2789 0 3
rlabel polysilicon 898 -2783 898 -2783 0 1
rlabel polysilicon 898 -2789 898 -2789 0 3
rlabel polysilicon 905 -2783 905 -2783 0 1
rlabel polysilicon 908 -2783 908 -2783 0 2
rlabel polysilicon 905 -2789 905 -2789 0 3
rlabel polysilicon 908 -2789 908 -2789 0 4
rlabel polysilicon 912 -2783 912 -2783 0 1
rlabel polysilicon 912 -2789 912 -2789 0 3
rlabel polysilicon 919 -2783 919 -2783 0 1
rlabel polysilicon 919 -2789 919 -2789 0 3
rlabel polysilicon 926 -2783 926 -2783 0 1
rlabel polysilicon 926 -2789 926 -2789 0 3
rlabel polysilicon 933 -2783 933 -2783 0 1
rlabel polysilicon 933 -2789 933 -2789 0 3
rlabel polysilicon 940 -2783 940 -2783 0 1
rlabel polysilicon 940 -2789 940 -2789 0 3
rlabel polysilicon 947 -2783 947 -2783 0 1
rlabel polysilicon 947 -2789 947 -2789 0 3
rlabel polysilicon 954 -2783 954 -2783 0 1
rlabel polysilicon 954 -2789 954 -2789 0 3
rlabel polysilicon 961 -2783 961 -2783 0 1
rlabel polysilicon 961 -2789 961 -2789 0 3
rlabel polysilicon 968 -2783 968 -2783 0 1
rlabel polysilicon 968 -2789 968 -2789 0 3
rlabel polysilicon 975 -2783 975 -2783 0 1
rlabel polysilicon 975 -2789 975 -2789 0 3
rlabel polysilicon 982 -2783 982 -2783 0 1
rlabel polysilicon 982 -2789 982 -2789 0 3
rlabel polysilicon 989 -2783 989 -2783 0 1
rlabel polysilicon 989 -2789 989 -2789 0 3
rlabel polysilicon 996 -2783 996 -2783 0 1
rlabel polysilicon 996 -2789 996 -2789 0 3
rlabel polysilicon 1003 -2789 1003 -2789 0 3
rlabel polysilicon 1006 -2789 1006 -2789 0 4
rlabel polysilicon 1010 -2783 1010 -2783 0 1
rlabel polysilicon 1010 -2789 1010 -2789 0 3
rlabel polysilicon 1017 -2783 1017 -2783 0 1
rlabel polysilicon 1017 -2789 1017 -2789 0 3
rlabel polysilicon 1024 -2783 1024 -2783 0 1
rlabel polysilicon 1024 -2789 1024 -2789 0 3
rlabel polysilicon 1031 -2783 1031 -2783 0 1
rlabel polysilicon 1031 -2789 1031 -2789 0 3
rlabel polysilicon 1038 -2783 1038 -2783 0 1
rlabel polysilicon 1038 -2789 1038 -2789 0 3
rlabel polysilicon 1045 -2783 1045 -2783 0 1
rlabel polysilicon 1045 -2789 1045 -2789 0 3
rlabel polysilicon 1052 -2783 1052 -2783 0 1
rlabel polysilicon 1052 -2789 1052 -2789 0 3
rlabel polysilicon 1059 -2783 1059 -2783 0 1
rlabel polysilicon 1059 -2789 1059 -2789 0 3
rlabel polysilicon 1066 -2783 1066 -2783 0 1
rlabel polysilicon 1066 -2789 1066 -2789 0 3
rlabel polysilicon 1073 -2783 1073 -2783 0 1
rlabel polysilicon 1073 -2789 1073 -2789 0 3
rlabel polysilicon 1080 -2783 1080 -2783 0 1
rlabel polysilicon 1080 -2789 1080 -2789 0 3
rlabel polysilicon 1087 -2783 1087 -2783 0 1
rlabel polysilicon 1087 -2789 1087 -2789 0 3
rlabel polysilicon 1094 -2783 1094 -2783 0 1
rlabel polysilicon 1094 -2789 1094 -2789 0 3
rlabel polysilicon 1101 -2783 1101 -2783 0 1
rlabel polysilicon 1101 -2789 1101 -2789 0 3
rlabel polysilicon 1108 -2783 1108 -2783 0 1
rlabel polysilicon 1108 -2789 1108 -2789 0 3
rlabel polysilicon 1115 -2783 1115 -2783 0 1
rlabel polysilicon 1115 -2789 1115 -2789 0 3
rlabel polysilicon 1122 -2783 1122 -2783 0 1
rlabel polysilicon 1122 -2789 1122 -2789 0 3
rlabel polysilicon 1129 -2783 1129 -2783 0 1
rlabel polysilicon 1129 -2789 1129 -2789 0 3
rlabel polysilicon 1136 -2783 1136 -2783 0 1
rlabel polysilicon 1136 -2789 1136 -2789 0 3
rlabel polysilicon 1143 -2783 1143 -2783 0 1
rlabel polysilicon 1143 -2789 1143 -2789 0 3
rlabel polysilicon 1150 -2783 1150 -2783 0 1
rlabel polysilicon 1150 -2789 1150 -2789 0 3
rlabel polysilicon 1157 -2783 1157 -2783 0 1
rlabel polysilicon 1160 -2783 1160 -2783 0 2
rlabel polysilicon 1157 -2789 1157 -2789 0 3
rlabel polysilicon 1160 -2789 1160 -2789 0 4
rlabel polysilicon 1164 -2783 1164 -2783 0 1
rlabel polysilicon 1164 -2789 1164 -2789 0 3
rlabel polysilicon 1171 -2783 1171 -2783 0 1
rlabel polysilicon 1171 -2789 1171 -2789 0 3
rlabel polysilicon 1178 -2783 1178 -2783 0 1
rlabel polysilicon 1178 -2789 1178 -2789 0 3
rlabel polysilicon 1185 -2783 1185 -2783 0 1
rlabel polysilicon 1188 -2783 1188 -2783 0 2
rlabel polysilicon 1185 -2789 1185 -2789 0 3
rlabel polysilicon 1192 -2783 1192 -2783 0 1
rlabel polysilicon 1192 -2789 1192 -2789 0 3
rlabel polysilicon 1199 -2783 1199 -2783 0 1
rlabel polysilicon 1199 -2789 1199 -2789 0 3
rlabel polysilicon 1206 -2783 1206 -2783 0 1
rlabel polysilicon 1206 -2789 1206 -2789 0 3
rlabel polysilicon 1213 -2783 1213 -2783 0 1
rlabel polysilicon 1213 -2789 1213 -2789 0 3
rlabel polysilicon 1220 -2783 1220 -2783 0 1
rlabel polysilicon 1220 -2789 1220 -2789 0 3
rlabel polysilicon 1227 -2783 1227 -2783 0 1
rlabel polysilicon 1227 -2789 1227 -2789 0 3
rlabel polysilicon 1234 -2783 1234 -2783 0 1
rlabel polysilicon 1234 -2789 1234 -2789 0 3
rlabel polysilicon 1241 -2783 1241 -2783 0 1
rlabel polysilicon 1241 -2789 1241 -2789 0 3
rlabel polysilicon 1248 -2783 1248 -2783 0 1
rlabel polysilicon 1248 -2789 1248 -2789 0 3
rlabel polysilicon 1255 -2783 1255 -2783 0 1
rlabel polysilicon 1255 -2789 1255 -2789 0 3
rlabel polysilicon 1262 -2783 1262 -2783 0 1
rlabel polysilicon 1262 -2789 1262 -2789 0 3
rlabel polysilicon 1269 -2783 1269 -2783 0 1
rlabel polysilicon 1269 -2789 1269 -2789 0 3
rlabel polysilicon 1276 -2783 1276 -2783 0 1
rlabel polysilicon 1276 -2789 1276 -2789 0 3
rlabel polysilicon 1283 -2783 1283 -2783 0 1
rlabel polysilicon 1283 -2789 1283 -2789 0 3
rlabel polysilicon 1290 -2783 1290 -2783 0 1
rlabel polysilicon 1290 -2789 1290 -2789 0 3
rlabel polysilicon 1300 -2783 1300 -2783 0 2
rlabel polysilicon 1297 -2789 1297 -2789 0 3
rlabel polysilicon 1300 -2789 1300 -2789 0 4
rlabel polysilicon 1304 -2783 1304 -2783 0 1
rlabel polysilicon 1304 -2789 1304 -2789 0 3
rlabel polysilicon 1311 -2783 1311 -2783 0 1
rlabel polysilicon 1311 -2789 1311 -2789 0 3
rlabel polysilicon 1318 -2783 1318 -2783 0 1
rlabel polysilicon 1318 -2789 1318 -2789 0 3
rlabel polysilicon 1325 -2783 1325 -2783 0 1
rlabel polysilicon 1325 -2789 1325 -2789 0 3
rlabel polysilicon 1332 -2783 1332 -2783 0 1
rlabel polysilicon 1332 -2789 1332 -2789 0 3
rlabel polysilicon 1339 -2783 1339 -2783 0 1
rlabel polysilicon 1339 -2789 1339 -2789 0 3
rlabel polysilicon 1346 -2783 1346 -2783 0 1
rlabel polysilicon 1346 -2789 1346 -2789 0 3
rlabel polysilicon 1353 -2783 1353 -2783 0 1
rlabel polysilicon 1353 -2789 1353 -2789 0 3
rlabel polysilicon 1360 -2783 1360 -2783 0 1
rlabel polysilicon 1360 -2789 1360 -2789 0 3
rlabel polysilicon 1367 -2783 1367 -2783 0 1
rlabel polysilicon 1367 -2789 1367 -2789 0 3
rlabel polysilicon 1374 -2783 1374 -2783 0 1
rlabel polysilicon 1374 -2789 1374 -2789 0 3
rlabel polysilicon 1381 -2783 1381 -2783 0 1
rlabel polysilicon 1381 -2789 1381 -2789 0 3
rlabel polysilicon 1388 -2783 1388 -2783 0 1
rlabel polysilicon 1388 -2789 1388 -2789 0 3
rlabel polysilicon 1395 -2783 1395 -2783 0 1
rlabel polysilicon 1395 -2789 1395 -2789 0 3
rlabel polysilicon 1402 -2783 1402 -2783 0 1
rlabel polysilicon 1402 -2789 1402 -2789 0 3
rlabel polysilicon 1409 -2783 1409 -2783 0 1
rlabel polysilicon 1409 -2789 1409 -2789 0 3
rlabel polysilicon 1416 -2783 1416 -2783 0 1
rlabel polysilicon 1416 -2789 1416 -2789 0 3
rlabel polysilicon 1423 -2783 1423 -2783 0 1
rlabel polysilicon 1423 -2789 1423 -2789 0 3
rlabel polysilicon 1430 -2783 1430 -2783 0 1
rlabel polysilicon 1430 -2789 1430 -2789 0 3
rlabel polysilicon 1437 -2783 1437 -2783 0 1
rlabel polysilicon 1437 -2789 1437 -2789 0 3
rlabel polysilicon 1444 -2783 1444 -2783 0 1
rlabel polysilicon 1444 -2789 1444 -2789 0 3
rlabel polysilicon 1451 -2783 1451 -2783 0 1
rlabel polysilicon 1451 -2789 1451 -2789 0 3
rlabel polysilicon 1458 -2783 1458 -2783 0 1
rlabel polysilicon 1458 -2789 1458 -2789 0 3
rlabel polysilicon 1465 -2783 1465 -2783 0 1
rlabel polysilicon 1465 -2789 1465 -2789 0 3
rlabel polysilicon 1472 -2783 1472 -2783 0 1
rlabel polysilicon 1472 -2789 1472 -2789 0 3
rlabel polysilicon 1479 -2783 1479 -2783 0 1
rlabel polysilicon 1479 -2789 1479 -2789 0 3
rlabel polysilicon 1486 -2783 1486 -2783 0 1
rlabel polysilicon 1486 -2789 1486 -2789 0 3
rlabel polysilicon 1493 -2783 1493 -2783 0 1
rlabel polysilicon 1493 -2789 1493 -2789 0 3
rlabel polysilicon 1500 -2783 1500 -2783 0 1
rlabel polysilicon 1500 -2789 1500 -2789 0 3
rlabel polysilicon 1507 -2783 1507 -2783 0 1
rlabel polysilicon 1507 -2789 1507 -2789 0 3
rlabel polysilicon 1514 -2783 1514 -2783 0 1
rlabel polysilicon 1514 -2789 1514 -2789 0 3
rlabel polysilicon 1521 -2783 1521 -2783 0 1
rlabel polysilicon 1524 -2783 1524 -2783 0 2
rlabel polysilicon 1521 -2789 1521 -2789 0 3
rlabel polysilicon 72 -2908 72 -2908 0 1
rlabel polysilicon 72 -2914 72 -2914 0 3
rlabel polysilicon 79 -2908 79 -2908 0 1
rlabel polysilicon 79 -2914 79 -2914 0 3
rlabel polysilicon 86 -2908 86 -2908 0 1
rlabel polysilicon 86 -2914 86 -2914 0 3
rlabel polysilicon 93 -2908 93 -2908 0 1
rlabel polysilicon 93 -2914 93 -2914 0 3
rlabel polysilicon 103 -2908 103 -2908 0 2
rlabel polysilicon 103 -2914 103 -2914 0 4
rlabel polysilicon 107 -2908 107 -2908 0 1
rlabel polysilicon 107 -2914 107 -2914 0 3
rlabel polysilicon 114 -2908 114 -2908 0 1
rlabel polysilicon 114 -2914 114 -2914 0 3
rlabel polysilicon 121 -2908 121 -2908 0 1
rlabel polysilicon 124 -2908 124 -2908 0 2
rlabel polysilicon 121 -2914 121 -2914 0 3
rlabel polysilicon 124 -2914 124 -2914 0 4
rlabel polysilicon 128 -2908 128 -2908 0 1
rlabel polysilicon 128 -2914 128 -2914 0 3
rlabel polysilicon 135 -2908 135 -2908 0 1
rlabel polysilicon 135 -2914 135 -2914 0 3
rlabel polysilicon 142 -2908 142 -2908 0 1
rlabel polysilicon 145 -2908 145 -2908 0 2
rlabel polysilicon 142 -2914 142 -2914 0 3
rlabel polysilicon 145 -2914 145 -2914 0 4
rlabel polysilicon 149 -2908 149 -2908 0 1
rlabel polysilicon 149 -2914 149 -2914 0 3
rlabel polysilicon 156 -2908 156 -2908 0 1
rlabel polysilicon 156 -2914 156 -2914 0 3
rlabel polysilicon 163 -2908 163 -2908 0 1
rlabel polysilicon 163 -2914 163 -2914 0 3
rlabel polysilicon 170 -2908 170 -2908 0 1
rlabel polysilicon 170 -2914 170 -2914 0 3
rlabel polysilicon 177 -2908 177 -2908 0 1
rlabel polysilicon 177 -2914 177 -2914 0 3
rlabel polysilicon 184 -2908 184 -2908 0 1
rlabel polysilicon 184 -2914 184 -2914 0 3
rlabel polysilicon 191 -2908 191 -2908 0 1
rlabel polysilicon 191 -2914 191 -2914 0 3
rlabel polysilicon 198 -2908 198 -2908 0 1
rlabel polysilicon 198 -2914 198 -2914 0 3
rlabel polysilicon 205 -2908 205 -2908 0 1
rlabel polysilicon 208 -2908 208 -2908 0 2
rlabel polysilicon 205 -2914 205 -2914 0 3
rlabel polysilicon 208 -2914 208 -2914 0 4
rlabel polysilicon 212 -2908 212 -2908 0 1
rlabel polysilicon 212 -2914 212 -2914 0 3
rlabel polysilicon 219 -2908 219 -2908 0 1
rlabel polysilicon 219 -2914 219 -2914 0 3
rlabel polysilicon 226 -2908 226 -2908 0 1
rlabel polysilicon 229 -2908 229 -2908 0 2
rlabel polysilicon 229 -2914 229 -2914 0 4
rlabel polysilicon 233 -2908 233 -2908 0 1
rlabel polysilicon 233 -2914 233 -2914 0 3
rlabel polysilicon 240 -2908 240 -2908 0 1
rlabel polysilicon 240 -2914 240 -2914 0 3
rlabel polysilicon 247 -2908 247 -2908 0 1
rlabel polysilicon 250 -2908 250 -2908 0 2
rlabel polysilicon 247 -2914 247 -2914 0 3
rlabel polysilicon 250 -2914 250 -2914 0 4
rlabel polysilicon 254 -2908 254 -2908 0 1
rlabel polysilicon 254 -2914 254 -2914 0 3
rlabel polysilicon 261 -2908 261 -2908 0 1
rlabel polysilicon 261 -2914 261 -2914 0 3
rlabel polysilicon 268 -2908 268 -2908 0 1
rlabel polysilicon 268 -2914 268 -2914 0 3
rlabel polysilicon 275 -2908 275 -2908 0 1
rlabel polysilicon 278 -2908 278 -2908 0 2
rlabel polysilicon 275 -2914 275 -2914 0 3
rlabel polysilicon 278 -2914 278 -2914 0 4
rlabel polysilicon 282 -2908 282 -2908 0 1
rlabel polysilicon 285 -2908 285 -2908 0 2
rlabel polysilicon 282 -2914 282 -2914 0 3
rlabel polysilicon 285 -2914 285 -2914 0 4
rlabel polysilicon 292 -2908 292 -2908 0 2
rlabel polysilicon 289 -2914 289 -2914 0 3
rlabel polysilicon 292 -2914 292 -2914 0 4
rlabel polysilicon 296 -2908 296 -2908 0 1
rlabel polysilicon 296 -2914 296 -2914 0 3
rlabel polysilicon 303 -2908 303 -2908 0 1
rlabel polysilicon 303 -2914 303 -2914 0 3
rlabel polysilicon 310 -2908 310 -2908 0 1
rlabel polysilicon 310 -2914 310 -2914 0 3
rlabel polysilicon 317 -2908 317 -2908 0 1
rlabel polysilicon 317 -2914 317 -2914 0 3
rlabel polysilicon 324 -2908 324 -2908 0 1
rlabel polysilicon 324 -2914 324 -2914 0 3
rlabel polysilicon 331 -2908 331 -2908 0 1
rlabel polysilicon 331 -2914 331 -2914 0 3
rlabel polysilicon 338 -2908 338 -2908 0 1
rlabel polysilicon 338 -2914 338 -2914 0 3
rlabel polysilicon 345 -2908 345 -2908 0 1
rlabel polysilicon 345 -2914 345 -2914 0 3
rlabel polysilicon 352 -2908 352 -2908 0 1
rlabel polysilicon 352 -2914 352 -2914 0 3
rlabel polysilicon 359 -2908 359 -2908 0 1
rlabel polysilicon 359 -2914 359 -2914 0 3
rlabel polysilicon 366 -2908 366 -2908 0 1
rlabel polysilicon 366 -2914 366 -2914 0 3
rlabel polysilicon 373 -2908 373 -2908 0 1
rlabel polysilicon 373 -2914 373 -2914 0 3
rlabel polysilicon 380 -2908 380 -2908 0 1
rlabel polysilicon 380 -2914 380 -2914 0 3
rlabel polysilicon 387 -2908 387 -2908 0 1
rlabel polysilicon 387 -2914 387 -2914 0 3
rlabel polysilicon 394 -2908 394 -2908 0 1
rlabel polysilicon 394 -2914 394 -2914 0 3
rlabel polysilicon 401 -2908 401 -2908 0 1
rlabel polysilicon 401 -2914 401 -2914 0 3
rlabel polysilicon 408 -2908 408 -2908 0 1
rlabel polysilicon 408 -2914 408 -2914 0 3
rlabel polysilicon 415 -2908 415 -2908 0 1
rlabel polysilicon 415 -2914 415 -2914 0 3
rlabel polysilicon 422 -2908 422 -2908 0 1
rlabel polysilicon 422 -2914 422 -2914 0 3
rlabel polysilicon 429 -2908 429 -2908 0 1
rlabel polysilicon 429 -2914 429 -2914 0 3
rlabel polysilicon 436 -2908 436 -2908 0 1
rlabel polysilicon 436 -2914 436 -2914 0 3
rlabel polysilicon 443 -2908 443 -2908 0 1
rlabel polysilicon 443 -2914 443 -2914 0 3
rlabel polysilicon 450 -2908 450 -2908 0 1
rlabel polysilicon 450 -2914 450 -2914 0 3
rlabel polysilicon 457 -2908 457 -2908 0 1
rlabel polysilicon 457 -2914 457 -2914 0 3
rlabel polysilicon 464 -2908 464 -2908 0 1
rlabel polysilicon 464 -2914 464 -2914 0 3
rlabel polysilicon 471 -2908 471 -2908 0 1
rlabel polysilicon 471 -2914 471 -2914 0 3
rlabel polysilicon 478 -2908 478 -2908 0 1
rlabel polysilicon 478 -2914 478 -2914 0 3
rlabel polysilicon 485 -2908 485 -2908 0 1
rlabel polysilicon 485 -2914 485 -2914 0 3
rlabel polysilicon 495 -2908 495 -2908 0 2
rlabel polysilicon 492 -2914 492 -2914 0 3
rlabel polysilicon 495 -2914 495 -2914 0 4
rlabel polysilicon 499 -2908 499 -2908 0 1
rlabel polysilicon 499 -2914 499 -2914 0 3
rlabel polysilicon 506 -2908 506 -2908 0 1
rlabel polysilicon 506 -2914 506 -2914 0 3
rlabel polysilicon 513 -2908 513 -2908 0 1
rlabel polysilicon 513 -2914 513 -2914 0 3
rlabel polysilicon 520 -2908 520 -2908 0 1
rlabel polysilicon 520 -2914 520 -2914 0 3
rlabel polysilicon 527 -2908 527 -2908 0 1
rlabel polysilicon 527 -2914 527 -2914 0 3
rlabel polysilicon 534 -2908 534 -2908 0 1
rlabel polysilicon 534 -2914 534 -2914 0 3
rlabel polysilicon 541 -2908 541 -2908 0 1
rlabel polysilicon 541 -2914 541 -2914 0 3
rlabel polysilicon 548 -2908 548 -2908 0 1
rlabel polysilicon 548 -2914 548 -2914 0 3
rlabel polysilicon 555 -2908 555 -2908 0 1
rlabel polysilicon 558 -2908 558 -2908 0 2
rlabel polysilicon 562 -2908 562 -2908 0 1
rlabel polysilicon 562 -2914 562 -2914 0 3
rlabel polysilicon 569 -2908 569 -2908 0 1
rlabel polysilicon 569 -2914 569 -2914 0 3
rlabel polysilicon 576 -2908 576 -2908 0 1
rlabel polysilicon 576 -2914 576 -2914 0 3
rlabel polysilicon 583 -2914 583 -2914 0 3
rlabel polysilicon 586 -2914 586 -2914 0 4
rlabel polysilicon 590 -2908 590 -2908 0 1
rlabel polysilicon 590 -2914 590 -2914 0 3
rlabel polysilicon 597 -2908 597 -2908 0 1
rlabel polysilicon 597 -2914 597 -2914 0 3
rlabel polysilicon 604 -2908 604 -2908 0 1
rlabel polysilicon 604 -2914 604 -2914 0 3
rlabel polysilicon 611 -2908 611 -2908 0 1
rlabel polysilicon 611 -2914 611 -2914 0 3
rlabel polysilicon 618 -2908 618 -2908 0 1
rlabel polysilicon 618 -2914 618 -2914 0 3
rlabel polysilicon 625 -2908 625 -2908 0 1
rlabel polysilicon 625 -2914 625 -2914 0 3
rlabel polysilicon 632 -2908 632 -2908 0 1
rlabel polysilicon 632 -2914 632 -2914 0 3
rlabel polysilicon 639 -2908 639 -2908 0 1
rlabel polysilicon 642 -2908 642 -2908 0 2
rlabel polysilicon 639 -2914 639 -2914 0 3
rlabel polysilicon 642 -2914 642 -2914 0 4
rlabel polysilicon 646 -2908 646 -2908 0 1
rlabel polysilicon 646 -2914 646 -2914 0 3
rlabel polysilicon 653 -2908 653 -2908 0 1
rlabel polysilicon 653 -2914 653 -2914 0 3
rlabel polysilicon 660 -2908 660 -2908 0 1
rlabel polysilicon 663 -2908 663 -2908 0 2
rlabel polysilicon 660 -2914 660 -2914 0 3
rlabel polysilicon 663 -2914 663 -2914 0 4
rlabel polysilicon 667 -2908 667 -2908 0 1
rlabel polysilicon 667 -2914 667 -2914 0 3
rlabel polysilicon 674 -2908 674 -2908 0 1
rlabel polysilicon 674 -2914 674 -2914 0 3
rlabel polysilicon 681 -2908 681 -2908 0 1
rlabel polysilicon 681 -2914 681 -2914 0 3
rlabel polysilicon 688 -2908 688 -2908 0 1
rlabel polysilicon 688 -2914 688 -2914 0 3
rlabel polysilicon 695 -2908 695 -2908 0 1
rlabel polysilicon 695 -2914 695 -2914 0 3
rlabel polysilicon 702 -2908 702 -2908 0 1
rlabel polysilicon 705 -2908 705 -2908 0 2
rlabel polysilicon 702 -2914 702 -2914 0 3
rlabel polysilicon 705 -2914 705 -2914 0 4
rlabel polysilicon 709 -2908 709 -2908 0 1
rlabel polysilicon 709 -2914 709 -2914 0 3
rlabel polysilicon 716 -2908 716 -2908 0 1
rlabel polysilicon 716 -2914 716 -2914 0 3
rlabel polysilicon 723 -2908 723 -2908 0 1
rlabel polysilicon 723 -2914 723 -2914 0 3
rlabel polysilicon 730 -2908 730 -2908 0 1
rlabel polysilicon 730 -2914 730 -2914 0 3
rlabel polysilicon 737 -2908 737 -2908 0 1
rlabel polysilicon 737 -2914 737 -2914 0 3
rlabel polysilicon 744 -2908 744 -2908 0 1
rlabel polysilicon 744 -2914 744 -2914 0 3
rlabel polysilicon 747 -2914 747 -2914 0 4
rlabel polysilicon 751 -2908 751 -2908 0 1
rlabel polysilicon 751 -2914 751 -2914 0 3
rlabel polysilicon 758 -2908 758 -2908 0 1
rlabel polysilicon 761 -2908 761 -2908 0 2
rlabel polysilicon 758 -2914 758 -2914 0 3
rlabel polysilicon 761 -2914 761 -2914 0 4
rlabel polysilicon 765 -2908 765 -2908 0 1
rlabel polysilicon 765 -2914 765 -2914 0 3
rlabel polysilicon 772 -2908 772 -2908 0 1
rlabel polysilicon 772 -2914 772 -2914 0 3
rlabel polysilicon 779 -2908 779 -2908 0 1
rlabel polysilicon 779 -2914 779 -2914 0 3
rlabel polysilicon 786 -2908 786 -2908 0 1
rlabel polysilicon 786 -2914 786 -2914 0 3
rlabel polysilicon 793 -2908 793 -2908 0 1
rlabel polysilicon 793 -2914 793 -2914 0 3
rlabel polysilicon 800 -2908 800 -2908 0 1
rlabel polysilicon 800 -2914 800 -2914 0 3
rlabel polysilicon 807 -2908 807 -2908 0 1
rlabel polysilicon 807 -2914 807 -2914 0 3
rlabel polysilicon 814 -2908 814 -2908 0 1
rlabel polysilicon 814 -2914 814 -2914 0 3
rlabel polysilicon 821 -2908 821 -2908 0 1
rlabel polysilicon 824 -2908 824 -2908 0 2
rlabel polysilicon 821 -2914 821 -2914 0 3
rlabel polysilicon 824 -2914 824 -2914 0 4
rlabel polysilicon 828 -2908 828 -2908 0 1
rlabel polysilicon 828 -2914 828 -2914 0 3
rlabel polysilicon 835 -2908 835 -2908 0 1
rlabel polysilicon 838 -2908 838 -2908 0 2
rlabel polysilicon 835 -2914 835 -2914 0 3
rlabel polysilicon 838 -2914 838 -2914 0 4
rlabel polysilicon 842 -2908 842 -2908 0 1
rlabel polysilicon 845 -2908 845 -2908 0 2
rlabel polysilicon 842 -2914 842 -2914 0 3
rlabel polysilicon 849 -2908 849 -2908 0 1
rlabel polysilicon 849 -2914 849 -2914 0 3
rlabel polysilicon 856 -2908 856 -2908 0 1
rlabel polysilicon 856 -2914 856 -2914 0 3
rlabel polysilicon 866 -2908 866 -2908 0 2
rlabel polysilicon 863 -2914 863 -2914 0 3
rlabel polysilicon 866 -2914 866 -2914 0 4
rlabel polysilicon 870 -2908 870 -2908 0 1
rlabel polysilicon 870 -2914 870 -2914 0 3
rlabel polysilicon 877 -2908 877 -2908 0 1
rlabel polysilicon 877 -2914 877 -2914 0 3
rlabel polysilicon 884 -2908 884 -2908 0 1
rlabel polysilicon 884 -2914 884 -2914 0 3
rlabel polysilicon 891 -2908 891 -2908 0 1
rlabel polysilicon 891 -2914 891 -2914 0 3
rlabel polysilicon 898 -2908 898 -2908 0 1
rlabel polysilicon 898 -2914 898 -2914 0 3
rlabel polysilicon 905 -2908 905 -2908 0 1
rlabel polysilicon 912 -2908 912 -2908 0 1
rlabel polysilicon 915 -2908 915 -2908 0 2
rlabel polysilicon 912 -2914 912 -2914 0 3
rlabel polysilicon 915 -2914 915 -2914 0 4
rlabel polysilicon 919 -2908 919 -2908 0 1
rlabel polysilicon 922 -2908 922 -2908 0 2
rlabel polysilicon 919 -2914 919 -2914 0 3
rlabel polysilicon 922 -2914 922 -2914 0 4
rlabel polysilicon 926 -2908 926 -2908 0 1
rlabel polysilicon 926 -2914 926 -2914 0 3
rlabel polysilicon 933 -2908 933 -2908 0 1
rlabel polysilicon 933 -2914 933 -2914 0 3
rlabel polysilicon 940 -2908 940 -2908 0 1
rlabel polysilicon 940 -2914 940 -2914 0 3
rlabel polysilicon 947 -2908 947 -2908 0 1
rlabel polysilicon 947 -2914 947 -2914 0 3
rlabel polysilicon 950 -2914 950 -2914 0 4
rlabel polysilicon 954 -2908 954 -2908 0 1
rlabel polysilicon 957 -2908 957 -2908 0 2
rlabel polysilicon 954 -2914 954 -2914 0 3
rlabel polysilicon 957 -2914 957 -2914 0 4
rlabel polysilicon 961 -2908 961 -2908 0 1
rlabel polysilicon 961 -2914 961 -2914 0 3
rlabel polysilicon 968 -2908 968 -2908 0 1
rlabel polysilicon 968 -2914 968 -2914 0 3
rlabel polysilicon 975 -2908 975 -2908 0 1
rlabel polysilicon 975 -2914 975 -2914 0 3
rlabel polysilicon 982 -2908 982 -2908 0 1
rlabel polysilicon 982 -2914 982 -2914 0 3
rlabel polysilicon 989 -2908 989 -2908 0 1
rlabel polysilicon 989 -2914 989 -2914 0 3
rlabel polysilicon 996 -2908 996 -2908 0 1
rlabel polysilicon 996 -2914 996 -2914 0 3
rlabel polysilicon 1003 -2908 1003 -2908 0 1
rlabel polysilicon 1003 -2914 1003 -2914 0 3
rlabel polysilicon 1010 -2908 1010 -2908 0 1
rlabel polysilicon 1010 -2914 1010 -2914 0 3
rlabel polysilicon 1017 -2908 1017 -2908 0 1
rlabel polysilicon 1020 -2908 1020 -2908 0 2
rlabel polysilicon 1017 -2914 1017 -2914 0 3
rlabel polysilicon 1020 -2914 1020 -2914 0 4
rlabel polysilicon 1024 -2908 1024 -2908 0 1
rlabel polysilicon 1024 -2914 1024 -2914 0 3
rlabel polysilicon 1031 -2908 1031 -2908 0 1
rlabel polysilicon 1031 -2914 1031 -2914 0 3
rlabel polysilicon 1038 -2908 1038 -2908 0 1
rlabel polysilicon 1038 -2914 1038 -2914 0 3
rlabel polysilicon 1045 -2908 1045 -2908 0 1
rlabel polysilicon 1045 -2914 1045 -2914 0 3
rlabel polysilicon 1052 -2908 1052 -2908 0 1
rlabel polysilicon 1052 -2914 1052 -2914 0 3
rlabel polysilicon 1059 -2908 1059 -2908 0 1
rlabel polysilicon 1059 -2914 1059 -2914 0 3
rlabel polysilicon 1066 -2908 1066 -2908 0 1
rlabel polysilicon 1066 -2914 1066 -2914 0 3
rlabel polysilicon 1073 -2908 1073 -2908 0 1
rlabel polysilicon 1073 -2914 1073 -2914 0 3
rlabel polysilicon 1080 -2908 1080 -2908 0 1
rlabel polysilicon 1080 -2914 1080 -2914 0 3
rlabel polysilicon 1087 -2908 1087 -2908 0 1
rlabel polysilicon 1087 -2914 1087 -2914 0 3
rlabel polysilicon 1094 -2908 1094 -2908 0 1
rlabel polysilicon 1097 -2908 1097 -2908 0 2
rlabel polysilicon 1094 -2914 1094 -2914 0 3
rlabel polysilicon 1097 -2914 1097 -2914 0 4
rlabel polysilicon 1101 -2908 1101 -2908 0 1
rlabel polysilicon 1101 -2914 1101 -2914 0 3
rlabel polysilicon 1108 -2908 1108 -2908 0 1
rlabel polysilicon 1108 -2914 1108 -2914 0 3
rlabel polysilicon 1115 -2908 1115 -2908 0 1
rlabel polysilicon 1115 -2914 1115 -2914 0 3
rlabel polysilicon 1122 -2908 1122 -2908 0 1
rlabel polysilicon 1122 -2914 1122 -2914 0 3
rlabel polysilicon 1129 -2908 1129 -2908 0 1
rlabel polysilicon 1129 -2914 1129 -2914 0 3
rlabel polysilicon 1136 -2908 1136 -2908 0 1
rlabel polysilicon 1136 -2914 1136 -2914 0 3
rlabel polysilicon 1143 -2908 1143 -2908 0 1
rlabel polysilicon 1143 -2914 1143 -2914 0 3
rlabel polysilicon 1150 -2908 1150 -2908 0 1
rlabel polysilicon 1150 -2914 1150 -2914 0 3
rlabel polysilicon 1157 -2908 1157 -2908 0 1
rlabel polysilicon 1157 -2914 1157 -2914 0 3
rlabel polysilicon 1164 -2908 1164 -2908 0 1
rlabel polysilicon 1164 -2914 1164 -2914 0 3
rlabel polysilicon 1171 -2908 1171 -2908 0 1
rlabel polysilicon 1171 -2914 1171 -2914 0 3
rlabel polysilicon 1178 -2908 1178 -2908 0 1
rlabel polysilicon 1178 -2914 1178 -2914 0 3
rlabel polysilicon 1185 -2908 1185 -2908 0 1
rlabel polysilicon 1185 -2914 1185 -2914 0 3
rlabel polysilicon 1192 -2908 1192 -2908 0 1
rlabel polysilicon 1192 -2914 1192 -2914 0 3
rlabel polysilicon 1199 -2908 1199 -2908 0 1
rlabel polysilicon 1199 -2914 1199 -2914 0 3
rlabel polysilicon 1206 -2908 1206 -2908 0 1
rlabel polysilicon 1206 -2914 1206 -2914 0 3
rlabel polysilicon 1213 -2908 1213 -2908 0 1
rlabel polysilicon 1213 -2914 1213 -2914 0 3
rlabel polysilicon 1220 -2908 1220 -2908 0 1
rlabel polysilicon 1220 -2914 1220 -2914 0 3
rlabel polysilicon 1227 -2908 1227 -2908 0 1
rlabel polysilicon 1227 -2914 1227 -2914 0 3
rlabel polysilicon 1230 -2914 1230 -2914 0 4
rlabel polysilicon 1234 -2908 1234 -2908 0 1
rlabel polysilicon 1234 -2914 1234 -2914 0 3
rlabel polysilicon 1241 -2908 1241 -2908 0 1
rlabel polysilicon 1241 -2914 1241 -2914 0 3
rlabel polysilicon 1248 -2908 1248 -2908 0 1
rlabel polysilicon 1248 -2914 1248 -2914 0 3
rlabel polysilicon 1255 -2908 1255 -2908 0 1
rlabel polysilicon 1255 -2914 1255 -2914 0 3
rlabel polysilicon 1262 -2908 1262 -2908 0 1
rlabel polysilicon 1262 -2914 1262 -2914 0 3
rlabel polysilicon 1269 -2908 1269 -2908 0 1
rlabel polysilicon 1269 -2914 1269 -2914 0 3
rlabel polysilicon 1276 -2908 1276 -2908 0 1
rlabel polysilicon 1276 -2914 1276 -2914 0 3
rlabel polysilicon 1283 -2908 1283 -2908 0 1
rlabel polysilicon 1283 -2914 1283 -2914 0 3
rlabel polysilicon 1290 -2908 1290 -2908 0 1
rlabel polysilicon 1290 -2914 1290 -2914 0 3
rlabel polysilicon 1297 -2908 1297 -2908 0 1
rlabel polysilicon 1297 -2914 1297 -2914 0 3
rlabel polysilicon 1304 -2908 1304 -2908 0 1
rlabel polysilicon 1304 -2914 1304 -2914 0 3
rlabel polysilicon 1311 -2908 1311 -2908 0 1
rlabel polysilicon 1311 -2914 1311 -2914 0 3
rlabel polysilicon 1318 -2908 1318 -2908 0 1
rlabel polysilicon 1318 -2914 1318 -2914 0 3
rlabel polysilicon 1325 -2908 1325 -2908 0 1
rlabel polysilicon 1325 -2914 1325 -2914 0 3
rlabel polysilicon 1332 -2908 1332 -2908 0 1
rlabel polysilicon 1332 -2914 1332 -2914 0 3
rlabel polysilicon 1339 -2908 1339 -2908 0 1
rlabel polysilicon 1339 -2914 1339 -2914 0 3
rlabel polysilicon 1346 -2908 1346 -2908 0 1
rlabel polysilicon 1346 -2914 1346 -2914 0 3
rlabel polysilicon 1353 -2908 1353 -2908 0 1
rlabel polysilicon 1353 -2914 1353 -2914 0 3
rlabel polysilicon 1363 -2908 1363 -2908 0 2
rlabel polysilicon 1360 -2914 1360 -2914 0 3
rlabel polysilicon 1367 -2908 1367 -2908 0 1
rlabel polysilicon 1367 -2914 1367 -2914 0 3
rlabel polysilicon 1374 -2908 1374 -2908 0 1
rlabel polysilicon 1374 -2914 1374 -2914 0 3
rlabel polysilicon 1381 -2908 1381 -2908 0 1
rlabel polysilicon 1381 -2914 1381 -2914 0 3
rlabel polysilicon 1388 -2908 1388 -2908 0 1
rlabel polysilicon 1388 -2914 1388 -2914 0 3
rlabel polysilicon 1395 -2908 1395 -2908 0 1
rlabel polysilicon 1395 -2914 1395 -2914 0 3
rlabel polysilicon 1402 -2908 1402 -2908 0 1
rlabel polysilicon 1402 -2914 1402 -2914 0 3
rlabel polysilicon 1409 -2908 1409 -2908 0 1
rlabel polysilicon 1409 -2914 1409 -2914 0 3
rlabel polysilicon 1416 -2908 1416 -2908 0 1
rlabel polysilicon 1416 -2914 1416 -2914 0 3
rlabel polysilicon 1423 -2908 1423 -2908 0 1
rlabel polysilicon 1423 -2914 1423 -2914 0 3
rlabel polysilicon 1430 -2908 1430 -2908 0 1
rlabel polysilicon 1430 -2914 1430 -2914 0 3
rlabel polysilicon 86 -3027 86 -3027 0 1
rlabel polysilicon 86 -3033 86 -3033 0 3
rlabel polysilicon 93 -3027 93 -3027 0 1
rlabel polysilicon 93 -3033 93 -3033 0 3
rlabel polysilicon 100 -3027 100 -3027 0 1
rlabel polysilicon 100 -3033 100 -3033 0 3
rlabel polysilicon 107 -3027 107 -3027 0 1
rlabel polysilicon 107 -3033 107 -3033 0 3
rlabel polysilicon 114 -3027 114 -3027 0 1
rlabel polysilicon 114 -3033 114 -3033 0 3
rlabel polysilicon 121 -3027 121 -3027 0 1
rlabel polysilicon 121 -3033 121 -3033 0 3
rlabel polysilicon 128 -3027 128 -3027 0 1
rlabel polysilicon 128 -3033 128 -3033 0 3
rlabel polysilicon 135 -3027 135 -3027 0 1
rlabel polysilicon 135 -3033 135 -3033 0 3
rlabel polysilicon 142 -3027 142 -3027 0 1
rlabel polysilicon 142 -3033 142 -3033 0 3
rlabel polysilicon 149 -3027 149 -3027 0 1
rlabel polysilicon 149 -3033 149 -3033 0 3
rlabel polysilicon 152 -3033 152 -3033 0 4
rlabel polysilicon 156 -3027 156 -3027 0 1
rlabel polysilicon 156 -3033 156 -3033 0 3
rlabel polysilicon 163 -3027 163 -3027 0 1
rlabel polysilicon 166 -3027 166 -3027 0 2
rlabel polysilicon 163 -3033 163 -3033 0 3
rlabel polysilicon 166 -3033 166 -3033 0 4
rlabel polysilicon 170 -3027 170 -3027 0 1
rlabel polysilicon 170 -3033 170 -3033 0 3
rlabel polysilicon 177 -3027 177 -3027 0 1
rlabel polysilicon 177 -3033 177 -3033 0 3
rlabel polysilicon 184 -3027 184 -3027 0 1
rlabel polysilicon 184 -3033 184 -3033 0 3
rlabel polysilicon 191 -3027 191 -3027 0 1
rlabel polysilicon 191 -3033 191 -3033 0 3
rlabel polysilicon 198 -3027 198 -3027 0 1
rlabel polysilicon 198 -3033 198 -3033 0 3
rlabel polysilicon 208 -3027 208 -3027 0 2
rlabel polysilicon 208 -3033 208 -3033 0 4
rlabel polysilicon 212 -3027 212 -3027 0 1
rlabel polysilicon 212 -3033 212 -3033 0 3
rlabel polysilicon 219 -3027 219 -3027 0 1
rlabel polysilicon 222 -3027 222 -3027 0 2
rlabel polysilicon 219 -3033 219 -3033 0 3
rlabel polysilicon 226 -3027 226 -3027 0 1
rlabel polysilicon 226 -3033 226 -3033 0 3
rlabel polysilicon 233 -3027 233 -3027 0 1
rlabel polysilicon 233 -3033 233 -3033 0 3
rlabel polysilicon 240 -3027 240 -3027 0 1
rlabel polysilicon 240 -3033 240 -3033 0 3
rlabel polysilicon 247 -3027 247 -3027 0 1
rlabel polysilicon 254 -3027 254 -3027 0 1
rlabel polysilicon 254 -3033 254 -3033 0 3
rlabel polysilicon 261 -3027 261 -3027 0 1
rlabel polysilicon 264 -3027 264 -3027 0 2
rlabel polysilicon 261 -3033 261 -3033 0 3
rlabel polysilicon 268 -3027 268 -3027 0 1
rlabel polysilicon 268 -3033 268 -3033 0 3
rlabel polysilicon 275 -3027 275 -3027 0 1
rlabel polysilicon 275 -3033 275 -3033 0 3
rlabel polysilicon 282 -3027 282 -3027 0 1
rlabel polysilicon 289 -3027 289 -3027 0 1
rlabel polysilicon 289 -3033 289 -3033 0 3
rlabel polysilicon 296 -3027 296 -3027 0 1
rlabel polysilicon 296 -3033 296 -3033 0 3
rlabel polysilicon 303 -3027 303 -3027 0 1
rlabel polysilicon 303 -3033 303 -3033 0 3
rlabel polysilicon 310 -3027 310 -3027 0 1
rlabel polysilicon 310 -3033 310 -3033 0 3
rlabel polysilicon 317 -3027 317 -3027 0 1
rlabel polysilicon 317 -3033 317 -3033 0 3
rlabel polysilicon 324 -3027 324 -3027 0 1
rlabel polysilicon 324 -3033 324 -3033 0 3
rlabel polysilicon 331 -3027 331 -3027 0 1
rlabel polysilicon 331 -3033 331 -3033 0 3
rlabel polysilicon 338 -3027 338 -3027 0 1
rlabel polysilicon 338 -3033 338 -3033 0 3
rlabel polysilicon 345 -3027 345 -3027 0 1
rlabel polysilicon 345 -3033 345 -3033 0 3
rlabel polysilicon 352 -3027 352 -3027 0 1
rlabel polysilicon 352 -3033 352 -3033 0 3
rlabel polysilicon 359 -3027 359 -3027 0 1
rlabel polysilicon 359 -3033 359 -3033 0 3
rlabel polysilicon 366 -3027 366 -3027 0 1
rlabel polysilicon 366 -3033 366 -3033 0 3
rlabel polysilicon 373 -3027 373 -3027 0 1
rlabel polysilicon 373 -3033 373 -3033 0 3
rlabel polysilicon 380 -3027 380 -3027 0 1
rlabel polysilicon 380 -3033 380 -3033 0 3
rlabel polysilicon 387 -3027 387 -3027 0 1
rlabel polysilicon 387 -3033 387 -3033 0 3
rlabel polysilicon 394 -3027 394 -3027 0 1
rlabel polysilicon 394 -3033 394 -3033 0 3
rlabel polysilicon 401 -3027 401 -3027 0 1
rlabel polysilicon 401 -3033 401 -3033 0 3
rlabel polysilicon 408 -3027 408 -3027 0 1
rlabel polysilicon 411 -3027 411 -3027 0 2
rlabel polysilicon 408 -3033 408 -3033 0 3
rlabel polysilicon 411 -3033 411 -3033 0 4
rlabel polysilicon 415 -3027 415 -3027 0 1
rlabel polysilicon 415 -3033 415 -3033 0 3
rlabel polysilicon 422 -3027 422 -3027 0 1
rlabel polysilicon 422 -3033 422 -3033 0 3
rlabel polysilicon 429 -3027 429 -3027 0 1
rlabel polysilicon 429 -3033 429 -3033 0 3
rlabel polysilicon 436 -3027 436 -3027 0 1
rlabel polysilicon 436 -3033 436 -3033 0 3
rlabel polysilicon 443 -3027 443 -3027 0 1
rlabel polysilicon 443 -3033 443 -3033 0 3
rlabel polysilicon 450 -3027 450 -3027 0 1
rlabel polysilicon 450 -3033 450 -3033 0 3
rlabel polysilicon 457 -3027 457 -3027 0 1
rlabel polysilicon 457 -3033 457 -3033 0 3
rlabel polysilicon 464 -3027 464 -3027 0 1
rlabel polysilicon 464 -3033 464 -3033 0 3
rlabel polysilicon 471 -3027 471 -3027 0 1
rlabel polysilicon 471 -3033 471 -3033 0 3
rlabel polysilicon 478 -3027 478 -3027 0 1
rlabel polysilicon 478 -3033 478 -3033 0 3
rlabel polysilicon 485 -3027 485 -3027 0 1
rlabel polysilicon 485 -3033 485 -3033 0 3
rlabel polysilicon 492 -3027 492 -3027 0 1
rlabel polysilicon 492 -3033 492 -3033 0 3
rlabel polysilicon 499 -3027 499 -3027 0 1
rlabel polysilicon 499 -3033 499 -3033 0 3
rlabel polysilicon 509 -3033 509 -3033 0 4
rlabel polysilicon 513 -3027 513 -3027 0 1
rlabel polysilicon 513 -3033 513 -3033 0 3
rlabel polysilicon 520 -3027 520 -3027 0 1
rlabel polysilicon 520 -3033 520 -3033 0 3
rlabel polysilicon 527 -3027 527 -3027 0 1
rlabel polysilicon 527 -3033 527 -3033 0 3
rlabel polysilicon 534 -3027 534 -3027 0 1
rlabel polysilicon 534 -3033 534 -3033 0 3
rlabel polysilicon 541 -3027 541 -3027 0 1
rlabel polysilicon 541 -3033 541 -3033 0 3
rlabel polysilicon 548 -3027 548 -3027 0 1
rlabel polysilicon 548 -3033 548 -3033 0 3
rlabel polysilicon 555 -3027 555 -3027 0 1
rlabel polysilicon 555 -3033 555 -3033 0 3
rlabel polysilicon 562 -3027 562 -3027 0 1
rlabel polysilicon 562 -3033 562 -3033 0 3
rlabel polysilicon 569 -3027 569 -3027 0 1
rlabel polysilicon 569 -3033 569 -3033 0 3
rlabel polysilicon 576 -3027 576 -3027 0 1
rlabel polysilicon 576 -3033 576 -3033 0 3
rlabel polysilicon 583 -3027 583 -3027 0 1
rlabel polysilicon 583 -3033 583 -3033 0 3
rlabel polysilicon 590 -3027 590 -3027 0 1
rlabel polysilicon 590 -3033 590 -3033 0 3
rlabel polysilicon 597 -3027 597 -3027 0 1
rlabel polysilicon 597 -3033 597 -3033 0 3
rlabel polysilicon 604 -3027 604 -3027 0 1
rlabel polysilicon 604 -3033 604 -3033 0 3
rlabel polysilicon 611 -3027 611 -3027 0 1
rlabel polysilicon 611 -3033 611 -3033 0 3
rlabel polysilicon 618 -3027 618 -3027 0 1
rlabel polysilicon 618 -3033 618 -3033 0 3
rlabel polysilicon 625 -3027 625 -3027 0 1
rlabel polysilicon 625 -3033 625 -3033 0 3
rlabel polysilicon 632 -3027 632 -3027 0 1
rlabel polysilicon 635 -3027 635 -3027 0 2
rlabel polysilicon 635 -3033 635 -3033 0 4
rlabel polysilicon 639 -3027 639 -3027 0 1
rlabel polysilicon 639 -3033 639 -3033 0 3
rlabel polysilicon 646 -3027 646 -3027 0 1
rlabel polysilicon 649 -3027 649 -3027 0 2
rlabel polysilicon 649 -3033 649 -3033 0 4
rlabel polysilicon 653 -3027 653 -3027 0 1
rlabel polysilicon 653 -3033 653 -3033 0 3
rlabel polysilicon 660 -3027 660 -3027 0 1
rlabel polysilicon 663 -3027 663 -3027 0 2
rlabel polysilicon 660 -3033 660 -3033 0 3
rlabel polysilicon 667 -3027 667 -3027 0 1
rlabel polysilicon 667 -3033 667 -3033 0 3
rlabel polysilicon 674 -3027 674 -3027 0 1
rlabel polysilicon 674 -3033 674 -3033 0 3
rlabel polysilicon 681 -3027 681 -3027 0 1
rlabel polysilicon 681 -3033 681 -3033 0 3
rlabel polysilicon 688 -3027 688 -3027 0 1
rlabel polysilicon 691 -3027 691 -3027 0 2
rlabel polysilicon 688 -3033 688 -3033 0 3
rlabel polysilicon 691 -3033 691 -3033 0 4
rlabel polysilicon 695 -3027 695 -3027 0 1
rlabel polysilicon 698 -3027 698 -3027 0 2
rlabel polysilicon 695 -3033 695 -3033 0 3
rlabel polysilicon 698 -3033 698 -3033 0 4
rlabel polysilicon 702 -3027 702 -3027 0 1
rlabel polysilicon 702 -3033 702 -3033 0 3
rlabel polysilicon 709 -3027 709 -3027 0 1
rlabel polysilicon 709 -3033 709 -3033 0 3
rlabel polysilicon 716 -3027 716 -3027 0 1
rlabel polysilicon 716 -3033 716 -3033 0 3
rlabel polysilicon 723 -3027 723 -3027 0 1
rlabel polysilicon 723 -3033 723 -3033 0 3
rlabel polysilicon 730 -3027 730 -3027 0 1
rlabel polysilicon 730 -3033 730 -3033 0 3
rlabel polysilicon 733 -3033 733 -3033 0 4
rlabel polysilicon 737 -3027 737 -3027 0 1
rlabel polysilicon 737 -3033 737 -3033 0 3
rlabel polysilicon 744 -3027 744 -3027 0 1
rlabel polysilicon 744 -3033 744 -3033 0 3
rlabel polysilicon 751 -3027 751 -3027 0 1
rlabel polysilicon 754 -3027 754 -3027 0 2
rlabel polysilicon 754 -3033 754 -3033 0 4
rlabel polysilicon 758 -3027 758 -3027 0 1
rlabel polysilicon 758 -3033 758 -3033 0 3
rlabel polysilicon 768 -3027 768 -3027 0 2
rlabel polysilicon 765 -3033 765 -3033 0 3
rlabel polysilicon 772 -3027 772 -3027 0 1
rlabel polysilicon 772 -3033 772 -3033 0 3
rlabel polysilicon 779 -3027 779 -3027 0 1
rlabel polysilicon 779 -3033 779 -3033 0 3
rlabel polysilicon 786 -3027 786 -3027 0 1
rlabel polysilicon 789 -3027 789 -3027 0 2
rlabel polysilicon 786 -3033 786 -3033 0 3
rlabel polysilicon 789 -3033 789 -3033 0 4
rlabel polysilicon 793 -3027 793 -3027 0 1
rlabel polysilicon 793 -3033 793 -3033 0 3
rlabel polysilicon 800 -3027 800 -3027 0 1
rlabel polysilicon 800 -3033 800 -3033 0 3
rlabel polysilicon 807 -3027 807 -3027 0 1
rlabel polysilicon 807 -3033 807 -3033 0 3
rlabel polysilicon 814 -3027 814 -3027 0 1
rlabel polysilicon 814 -3033 814 -3033 0 3
rlabel polysilicon 821 -3027 821 -3027 0 1
rlabel polysilicon 821 -3033 821 -3033 0 3
rlabel polysilicon 828 -3027 828 -3027 0 1
rlabel polysilicon 828 -3033 828 -3033 0 3
rlabel polysilicon 835 -3027 835 -3027 0 1
rlabel polysilicon 838 -3027 838 -3027 0 2
rlabel polysilicon 835 -3033 835 -3033 0 3
rlabel polysilicon 838 -3033 838 -3033 0 4
rlabel polysilicon 842 -3027 842 -3027 0 1
rlabel polysilicon 842 -3033 842 -3033 0 3
rlabel polysilicon 849 -3027 849 -3027 0 1
rlabel polysilicon 849 -3033 849 -3033 0 3
rlabel polysilicon 856 -3027 856 -3027 0 1
rlabel polysilicon 856 -3033 856 -3033 0 3
rlabel polysilicon 863 -3027 863 -3027 0 1
rlabel polysilicon 866 -3027 866 -3027 0 2
rlabel polysilicon 863 -3033 863 -3033 0 3
rlabel polysilicon 866 -3033 866 -3033 0 4
rlabel polysilicon 870 -3027 870 -3027 0 1
rlabel polysilicon 873 -3027 873 -3027 0 2
rlabel polysilicon 873 -3033 873 -3033 0 4
rlabel polysilicon 877 -3027 877 -3027 0 1
rlabel polysilicon 877 -3033 877 -3033 0 3
rlabel polysilicon 884 -3027 884 -3027 0 1
rlabel polysilicon 884 -3033 884 -3033 0 3
rlabel polysilicon 887 -3033 887 -3033 0 4
rlabel polysilicon 891 -3027 891 -3027 0 1
rlabel polysilicon 891 -3033 891 -3033 0 3
rlabel polysilicon 898 -3027 898 -3027 0 1
rlabel polysilicon 898 -3033 898 -3033 0 3
rlabel polysilicon 905 -3033 905 -3033 0 3
rlabel polysilicon 912 -3027 912 -3027 0 1
rlabel polysilicon 915 -3027 915 -3027 0 2
rlabel polysilicon 912 -3033 912 -3033 0 3
rlabel polysilicon 919 -3027 919 -3027 0 1
rlabel polysilicon 922 -3027 922 -3027 0 2
rlabel polysilicon 919 -3033 919 -3033 0 3
rlabel polysilicon 922 -3033 922 -3033 0 4
rlabel polysilicon 926 -3027 926 -3027 0 1
rlabel polysilicon 926 -3033 926 -3033 0 3
rlabel polysilicon 933 -3027 933 -3027 0 1
rlabel polysilicon 933 -3033 933 -3033 0 3
rlabel polysilicon 940 -3027 940 -3027 0 1
rlabel polysilicon 940 -3033 940 -3033 0 3
rlabel polysilicon 947 -3027 947 -3027 0 1
rlabel polysilicon 947 -3033 947 -3033 0 3
rlabel polysilicon 954 -3027 954 -3027 0 1
rlabel polysilicon 954 -3033 954 -3033 0 3
rlabel polysilicon 961 -3027 961 -3027 0 1
rlabel polysilicon 961 -3033 961 -3033 0 3
rlabel polysilicon 968 -3027 968 -3027 0 1
rlabel polysilicon 968 -3033 968 -3033 0 3
rlabel polysilicon 975 -3027 975 -3027 0 1
rlabel polysilicon 975 -3033 975 -3033 0 3
rlabel polysilicon 982 -3027 982 -3027 0 1
rlabel polysilicon 982 -3033 982 -3033 0 3
rlabel polysilicon 989 -3027 989 -3027 0 1
rlabel polysilicon 989 -3033 989 -3033 0 3
rlabel polysilicon 996 -3027 996 -3027 0 1
rlabel polysilicon 996 -3033 996 -3033 0 3
rlabel polysilicon 1003 -3027 1003 -3027 0 1
rlabel polysilicon 1003 -3033 1003 -3033 0 3
rlabel polysilicon 1010 -3027 1010 -3027 0 1
rlabel polysilicon 1010 -3033 1010 -3033 0 3
rlabel polysilicon 1017 -3027 1017 -3027 0 1
rlabel polysilicon 1020 -3033 1020 -3033 0 4
rlabel polysilicon 1024 -3027 1024 -3027 0 1
rlabel polysilicon 1024 -3033 1024 -3033 0 3
rlabel polysilicon 1031 -3027 1031 -3027 0 1
rlabel polysilicon 1031 -3033 1031 -3033 0 3
rlabel polysilicon 1038 -3027 1038 -3027 0 1
rlabel polysilicon 1038 -3033 1038 -3033 0 3
rlabel polysilicon 1045 -3027 1045 -3027 0 1
rlabel polysilicon 1045 -3033 1045 -3033 0 3
rlabel polysilicon 1052 -3027 1052 -3027 0 1
rlabel polysilicon 1052 -3033 1052 -3033 0 3
rlabel polysilicon 1059 -3027 1059 -3027 0 1
rlabel polysilicon 1059 -3033 1059 -3033 0 3
rlabel polysilicon 1066 -3027 1066 -3027 0 1
rlabel polysilicon 1066 -3033 1066 -3033 0 3
rlabel polysilicon 1073 -3027 1073 -3027 0 1
rlabel polysilicon 1076 -3027 1076 -3027 0 2
rlabel polysilicon 1073 -3033 1073 -3033 0 3
rlabel polysilicon 1080 -3027 1080 -3027 0 1
rlabel polysilicon 1080 -3033 1080 -3033 0 3
rlabel polysilicon 1087 -3027 1087 -3027 0 1
rlabel polysilicon 1087 -3033 1087 -3033 0 3
rlabel polysilicon 1094 -3027 1094 -3027 0 1
rlabel polysilicon 1094 -3033 1094 -3033 0 3
rlabel polysilicon 1101 -3027 1101 -3027 0 1
rlabel polysilicon 1101 -3033 1101 -3033 0 3
rlabel polysilicon 1108 -3027 1108 -3027 0 1
rlabel polysilicon 1108 -3033 1108 -3033 0 3
rlabel polysilicon 1115 -3027 1115 -3027 0 1
rlabel polysilicon 1115 -3033 1115 -3033 0 3
rlabel polysilicon 1122 -3027 1122 -3027 0 1
rlabel polysilicon 1122 -3033 1122 -3033 0 3
rlabel polysilicon 1129 -3027 1129 -3027 0 1
rlabel polysilicon 1129 -3033 1129 -3033 0 3
rlabel polysilicon 1136 -3027 1136 -3027 0 1
rlabel polysilicon 1136 -3033 1136 -3033 0 3
rlabel polysilicon 1143 -3027 1143 -3027 0 1
rlabel polysilicon 1143 -3033 1143 -3033 0 3
rlabel polysilicon 1150 -3033 1150 -3033 0 3
rlabel polysilicon 1153 -3033 1153 -3033 0 4
rlabel polysilicon 1157 -3027 1157 -3027 0 1
rlabel polysilicon 1157 -3033 1157 -3033 0 3
rlabel polysilicon 1164 -3027 1164 -3027 0 1
rlabel polysilicon 1164 -3033 1164 -3033 0 3
rlabel polysilicon 1171 -3027 1171 -3027 0 1
rlabel polysilicon 1171 -3033 1171 -3033 0 3
rlabel polysilicon 1178 -3027 1178 -3027 0 1
rlabel polysilicon 1178 -3033 1178 -3033 0 3
rlabel polysilicon 1185 -3027 1185 -3027 0 1
rlabel polysilicon 1185 -3033 1185 -3033 0 3
rlabel polysilicon 1192 -3027 1192 -3027 0 1
rlabel polysilicon 1192 -3033 1192 -3033 0 3
rlabel polysilicon 1199 -3027 1199 -3027 0 1
rlabel polysilicon 1199 -3033 1199 -3033 0 3
rlabel polysilicon 1206 -3027 1206 -3027 0 1
rlabel polysilicon 1206 -3033 1206 -3033 0 3
rlabel polysilicon 1213 -3027 1213 -3027 0 1
rlabel polysilicon 1213 -3033 1213 -3033 0 3
rlabel polysilicon 1220 -3027 1220 -3027 0 1
rlabel polysilicon 1220 -3033 1220 -3033 0 3
rlabel polysilicon 1227 -3027 1227 -3027 0 1
rlabel polysilicon 1230 -3027 1230 -3027 0 2
rlabel polysilicon 1227 -3033 1227 -3033 0 3
rlabel polysilicon 1234 -3027 1234 -3027 0 1
rlabel polysilicon 1234 -3033 1234 -3033 0 3
rlabel polysilicon 1241 -3027 1241 -3027 0 1
rlabel polysilicon 1241 -3033 1241 -3033 0 3
rlabel polysilicon 1248 -3027 1248 -3027 0 1
rlabel polysilicon 1248 -3033 1248 -3033 0 3
rlabel polysilicon 1255 -3027 1255 -3027 0 1
rlabel polysilicon 1255 -3033 1255 -3033 0 3
rlabel polysilicon 1262 -3027 1262 -3027 0 1
rlabel polysilicon 1262 -3033 1262 -3033 0 3
rlabel polysilicon 1269 -3027 1269 -3027 0 1
rlabel polysilicon 1269 -3033 1269 -3033 0 3
rlabel polysilicon 1276 -3027 1276 -3027 0 1
rlabel polysilicon 1276 -3033 1276 -3033 0 3
rlabel polysilicon 1283 -3027 1283 -3027 0 1
rlabel polysilicon 1283 -3033 1283 -3033 0 3
rlabel polysilicon 1290 -3027 1290 -3027 0 1
rlabel polysilicon 1290 -3033 1290 -3033 0 3
rlabel polysilicon 1297 -3027 1297 -3027 0 1
rlabel polysilicon 1297 -3033 1297 -3033 0 3
rlabel polysilicon 1304 -3027 1304 -3027 0 1
rlabel polysilicon 1304 -3033 1304 -3033 0 3
rlabel polysilicon 1311 -3027 1311 -3027 0 1
rlabel polysilicon 1311 -3033 1311 -3033 0 3
rlabel polysilicon 1318 -3027 1318 -3027 0 1
rlabel polysilicon 1318 -3033 1318 -3033 0 3
rlabel polysilicon 1325 -3027 1325 -3027 0 1
rlabel polysilicon 1325 -3033 1325 -3033 0 3
rlabel polysilicon 1332 -3027 1332 -3027 0 1
rlabel polysilicon 1332 -3033 1332 -3033 0 3
rlabel polysilicon 1339 -3027 1339 -3027 0 1
rlabel polysilicon 1339 -3033 1339 -3033 0 3
rlabel polysilicon 1346 -3027 1346 -3027 0 1
rlabel polysilicon 1346 -3033 1346 -3033 0 3
rlabel polysilicon 1353 -3027 1353 -3027 0 1
rlabel polysilicon 1353 -3033 1353 -3033 0 3
rlabel polysilicon 1360 -3027 1360 -3027 0 1
rlabel polysilicon 1360 -3033 1360 -3033 0 3
rlabel polysilicon 1367 -3027 1367 -3027 0 1
rlabel polysilicon 1367 -3033 1367 -3033 0 3
rlabel polysilicon 1374 -3027 1374 -3027 0 1
rlabel polysilicon 1374 -3033 1374 -3033 0 3
rlabel polysilicon 1381 -3027 1381 -3027 0 1
rlabel polysilicon 1381 -3033 1381 -3033 0 3
rlabel polysilicon 1388 -3027 1388 -3027 0 1
rlabel polysilicon 1388 -3033 1388 -3033 0 3
rlabel polysilicon 1395 -3027 1395 -3027 0 1
rlabel polysilicon 1395 -3033 1395 -3033 0 3
rlabel polysilicon 1402 -3027 1402 -3027 0 1
rlabel polysilicon 1402 -3033 1402 -3033 0 3
rlabel polysilicon 1409 -3027 1409 -3027 0 1
rlabel polysilicon 1409 -3033 1409 -3033 0 3
rlabel polysilicon 100 -3138 100 -3138 0 1
rlabel polysilicon 100 -3144 100 -3144 0 3
rlabel polysilicon 107 -3138 107 -3138 0 1
rlabel polysilicon 107 -3144 107 -3144 0 3
rlabel polysilicon 114 -3138 114 -3138 0 1
rlabel polysilicon 114 -3144 114 -3144 0 3
rlabel polysilicon 121 -3138 121 -3138 0 1
rlabel polysilicon 121 -3144 121 -3144 0 3
rlabel polysilicon 128 -3138 128 -3138 0 1
rlabel polysilicon 128 -3144 128 -3144 0 3
rlabel polysilicon 135 -3138 135 -3138 0 1
rlabel polysilicon 135 -3144 135 -3144 0 3
rlabel polysilicon 142 -3138 142 -3138 0 1
rlabel polysilicon 142 -3144 142 -3144 0 3
rlabel polysilicon 149 -3138 149 -3138 0 1
rlabel polysilicon 149 -3144 149 -3144 0 3
rlabel polysilicon 156 -3138 156 -3138 0 1
rlabel polysilicon 156 -3144 156 -3144 0 3
rlabel polysilicon 159 -3144 159 -3144 0 4
rlabel polysilicon 163 -3138 163 -3138 0 1
rlabel polysilicon 163 -3144 163 -3144 0 3
rlabel polysilicon 170 -3138 170 -3138 0 1
rlabel polysilicon 170 -3144 170 -3144 0 3
rlabel polysilicon 177 -3138 177 -3138 0 1
rlabel polysilicon 177 -3144 177 -3144 0 3
rlabel polysilicon 184 -3138 184 -3138 0 1
rlabel polysilicon 184 -3144 184 -3144 0 3
rlabel polysilicon 191 -3138 191 -3138 0 1
rlabel polysilicon 191 -3144 191 -3144 0 3
rlabel polysilicon 198 -3138 198 -3138 0 1
rlabel polysilicon 198 -3144 198 -3144 0 3
rlabel polysilicon 205 -3138 205 -3138 0 1
rlabel polysilicon 205 -3144 205 -3144 0 3
rlabel polysilicon 212 -3138 212 -3138 0 1
rlabel polysilicon 212 -3144 212 -3144 0 3
rlabel polysilicon 222 -3138 222 -3138 0 2
rlabel polysilicon 222 -3144 222 -3144 0 4
rlabel polysilicon 226 -3138 226 -3138 0 1
rlabel polysilicon 229 -3138 229 -3138 0 2
rlabel polysilicon 229 -3144 229 -3144 0 4
rlabel polysilicon 233 -3138 233 -3138 0 1
rlabel polysilicon 233 -3144 233 -3144 0 3
rlabel polysilicon 240 -3138 240 -3138 0 1
rlabel polysilicon 240 -3144 240 -3144 0 3
rlabel polysilicon 247 -3138 247 -3138 0 1
rlabel polysilicon 247 -3144 247 -3144 0 3
rlabel polysilicon 250 -3144 250 -3144 0 4
rlabel polysilicon 254 -3138 254 -3138 0 1
rlabel polysilicon 257 -3138 257 -3138 0 2
rlabel polysilicon 261 -3138 261 -3138 0 1
rlabel polysilicon 261 -3144 261 -3144 0 3
rlabel polysilicon 268 -3138 268 -3138 0 1
rlabel polysilicon 268 -3144 268 -3144 0 3
rlabel polysilicon 275 -3138 275 -3138 0 1
rlabel polysilicon 275 -3144 275 -3144 0 3
rlabel polysilicon 282 -3144 282 -3144 0 3
rlabel polysilicon 289 -3138 289 -3138 0 1
rlabel polysilicon 289 -3144 289 -3144 0 3
rlabel polysilicon 296 -3138 296 -3138 0 1
rlabel polysilicon 296 -3144 296 -3144 0 3
rlabel polysilicon 303 -3138 303 -3138 0 1
rlabel polysilicon 303 -3144 303 -3144 0 3
rlabel polysilicon 310 -3138 310 -3138 0 1
rlabel polysilicon 310 -3144 310 -3144 0 3
rlabel polysilicon 317 -3138 317 -3138 0 1
rlabel polysilicon 317 -3144 317 -3144 0 3
rlabel polysilicon 324 -3138 324 -3138 0 1
rlabel polysilicon 327 -3138 327 -3138 0 2
rlabel polysilicon 324 -3144 324 -3144 0 3
rlabel polysilicon 327 -3144 327 -3144 0 4
rlabel polysilicon 331 -3138 331 -3138 0 1
rlabel polysilicon 331 -3144 331 -3144 0 3
rlabel polysilicon 338 -3138 338 -3138 0 1
rlabel polysilicon 338 -3144 338 -3144 0 3
rlabel polysilicon 345 -3138 345 -3138 0 1
rlabel polysilicon 345 -3144 345 -3144 0 3
rlabel polysilicon 352 -3138 352 -3138 0 1
rlabel polysilicon 352 -3144 352 -3144 0 3
rlabel polysilicon 359 -3138 359 -3138 0 1
rlabel polysilicon 359 -3144 359 -3144 0 3
rlabel polysilicon 366 -3138 366 -3138 0 1
rlabel polysilicon 366 -3144 366 -3144 0 3
rlabel polysilicon 373 -3138 373 -3138 0 1
rlabel polysilicon 373 -3144 373 -3144 0 3
rlabel polysilicon 380 -3138 380 -3138 0 1
rlabel polysilicon 380 -3144 380 -3144 0 3
rlabel polysilicon 387 -3144 387 -3144 0 3
rlabel polysilicon 390 -3144 390 -3144 0 4
rlabel polysilicon 394 -3138 394 -3138 0 1
rlabel polysilicon 394 -3144 394 -3144 0 3
rlabel polysilicon 401 -3138 401 -3138 0 1
rlabel polysilicon 401 -3144 401 -3144 0 3
rlabel polysilicon 411 -3138 411 -3138 0 2
rlabel polysilicon 408 -3144 408 -3144 0 3
rlabel polysilicon 411 -3144 411 -3144 0 4
rlabel polysilicon 415 -3138 415 -3138 0 1
rlabel polysilicon 415 -3144 415 -3144 0 3
rlabel polysilicon 422 -3138 422 -3138 0 1
rlabel polysilicon 422 -3144 422 -3144 0 3
rlabel polysilicon 429 -3138 429 -3138 0 1
rlabel polysilicon 429 -3144 429 -3144 0 3
rlabel polysilicon 436 -3138 436 -3138 0 1
rlabel polysilicon 436 -3144 436 -3144 0 3
rlabel polysilicon 443 -3138 443 -3138 0 1
rlabel polysilicon 443 -3144 443 -3144 0 3
rlabel polysilicon 450 -3138 450 -3138 0 1
rlabel polysilicon 450 -3144 450 -3144 0 3
rlabel polysilicon 457 -3138 457 -3138 0 1
rlabel polysilicon 457 -3144 457 -3144 0 3
rlabel polysilicon 464 -3138 464 -3138 0 1
rlabel polysilicon 464 -3144 464 -3144 0 3
rlabel polysilicon 471 -3138 471 -3138 0 1
rlabel polysilicon 471 -3144 471 -3144 0 3
rlabel polysilicon 478 -3138 478 -3138 0 1
rlabel polysilicon 478 -3144 478 -3144 0 3
rlabel polysilicon 485 -3138 485 -3138 0 1
rlabel polysilicon 485 -3144 485 -3144 0 3
rlabel polysilicon 492 -3138 492 -3138 0 1
rlabel polysilicon 492 -3144 492 -3144 0 3
rlabel polysilicon 499 -3138 499 -3138 0 1
rlabel polysilicon 499 -3144 499 -3144 0 3
rlabel polysilicon 506 -3138 506 -3138 0 1
rlabel polysilicon 506 -3144 506 -3144 0 3
rlabel polysilicon 513 -3138 513 -3138 0 1
rlabel polysilicon 516 -3138 516 -3138 0 2
rlabel polysilicon 513 -3144 513 -3144 0 3
rlabel polysilicon 516 -3144 516 -3144 0 4
rlabel polysilicon 520 -3138 520 -3138 0 1
rlabel polysilicon 520 -3144 520 -3144 0 3
rlabel polysilicon 527 -3138 527 -3138 0 1
rlabel polysilicon 527 -3144 527 -3144 0 3
rlabel polysilicon 534 -3138 534 -3138 0 1
rlabel polysilicon 534 -3144 534 -3144 0 3
rlabel polysilicon 541 -3138 541 -3138 0 1
rlabel polysilicon 541 -3144 541 -3144 0 3
rlabel polysilicon 548 -3138 548 -3138 0 1
rlabel polysilicon 548 -3144 548 -3144 0 3
rlabel polysilicon 555 -3138 555 -3138 0 1
rlabel polysilicon 555 -3144 555 -3144 0 3
rlabel polysilicon 562 -3138 562 -3138 0 1
rlabel polysilicon 562 -3144 562 -3144 0 3
rlabel polysilicon 569 -3138 569 -3138 0 1
rlabel polysilicon 569 -3144 569 -3144 0 3
rlabel polysilicon 576 -3138 576 -3138 0 1
rlabel polysilicon 576 -3144 576 -3144 0 3
rlabel polysilicon 583 -3138 583 -3138 0 1
rlabel polysilicon 583 -3144 583 -3144 0 3
rlabel polysilicon 590 -3138 590 -3138 0 1
rlabel polysilicon 590 -3144 590 -3144 0 3
rlabel polysilicon 593 -3144 593 -3144 0 4
rlabel polysilicon 597 -3138 597 -3138 0 1
rlabel polysilicon 597 -3144 597 -3144 0 3
rlabel polysilicon 607 -3138 607 -3138 0 2
rlabel polysilicon 604 -3144 604 -3144 0 3
rlabel polysilicon 607 -3144 607 -3144 0 4
rlabel polysilicon 611 -3138 611 -3138 0 1
rlabel polysilicon 611 -3144 611 -3144 0 3
rlabel polysilicon 618 -3138 618 -3138 0 1
rlabel polysilicon 618 -3144 618 -3144 0 3
rlabel polysilicon 625 -3138 625 -3138 0 1
rlabel polysilicon 625 -3144 625 -3144 0 3
rlabel polysilicon 632 -3138 632 -3138 0 1
rlabel polysilicon 632 -3144 632 -3144 0 3
rlabel polysilicon 639 -3138 639 -3138 0 1
rlabel polysilicon 639 -3144 639 -3144 0 3
rlabel polysilicon 646 -3138 646 -3138 0 1
rlabel polysilicon 649 -3138 649 -3138 0 2
rlabel polysilicon 646 -3144 646 -3144 0 3
rlabel polysilicon 653 -3138 653 -3138 0 1
rlabel polysilicon 653 -3144 653 -3144 0 3
rlabel polysilicon 660 -3138 660 -3138 0 1
rlabel polysilicon 660 -3144 660 -3144 0 3
rlabel polysilicon 667 -3138 667 -3138 0 1
rlabel polysilicon 667 -3144 667 -3144 0 3
rlabel polysilicon 674 -3138 674 -3138 0 1
rlabel polysilicon 674 -3144 674 -3144 0 3
rlabel polysilicon 681 -3138 681 -3138 0 1
rlabel polysilicon 681 -3144 681 -3144 0 3
rlabel polysilicon 688 -3138 688 -3138 0 1
rlabel polysilicon 688 -3144 688 -3144 0 3
rlabel polysilicon 695 -3138 695 -3138 0 1
rlabel polysilicon 698 -3138 698 -3138 0 2
rlabel polysilicon 695 -3144 695 -3144 0 3
rlabel polysilicon 698 -3144 698 -3144 0 4
rlabel polysilicon 702 -3138 702 -3138 0 1
rlabel polysilicon 702 -3144 702 -3144 0 3
rlabel polysilicon 709 -3138 709 -3138 0 1
rlabel polysilicon 709 -3144 709 -3144 0 3
rlabel polysilicon 716 -3138 716 -3138 0 1
rlabel polysilicon 716 -3144 716 -3144 0 3
rlabel polysilicon 723 -3138 723 -3138 0 1
rlabel polysilicon 723 -3144 723 -3144 0 3
rlabel polysilicon 730 -3138 730 -3138 0 1
rlabel polysilicon 733 -3138 733 -3138 0 2
rlabel polysilicon 730 -3144 730 -3144 0 3
rlabel polysilicon 737 -3138 737 -3138 0 1
rlabel polysilicon 740 -3138 740 -3138 0 2
rlabel polysilicon 737 -3144 737 -3144 0 3
rlabel polysilicon 740 -3144 740 -3144 0 4
rlabel polysilicon 744 -3138 744 -3138 0 1
rlabel polysilicon 747 -3138 747 -3138 0 2
rlabel polysilicon 744 -3144 744 -3144 0 3
rlabel polysilicon 747 -3144 747 -3144 0 4
rlabel polysilicon 751 -3138 751 -3138 0 1
rlabel polysilicon 751 -3144 751 -3144 0 3
rlabel polysilicon 761 -3138 761 -3138 0 2
rlabel polysilicon 758 -3144 758 -3144 0 3
rlabel polysilicon 761 -3144 761 -3144 0 4
rlabel polysilicon 765 -3138 765 -3138 0 1
rlabel polysilicon 765 -3144 765 -3144 0 3
rlabel polysilicon 772 -3138 772 -3138 0 1
rlabel polysilicon 772 -3144 772 -3144 0 3
rlabel polysilicon 779 -3138 779 -3138 0 1
rlabel polysilicon 779 -3144 779 -3144 0 3
rlabel polysilicon 786 -3138 786 -3138 0 1
rlabel polysilicon 786 -3144 786 -3144 0 3
rlabel polysilicon 793 -3138 793 -3138 0 1
rlabel polysilicon 796 -3138 796 -3138 0 2
rlabel polysilicon 793 -3144 793 -3144 0 3
rlabel polysilicon 796 -3144 796 -3144 0 4
rlabel polysilicon 800 -3138 800 -3138 0 1
rlabel polysilicon 800 -3144 800 -3144 0 3
rlabel polysilicon 807 -3138 807 -3138 0 1
rlabel polysilicon 810 -3138 810 -3138 0 2
rlabel polysilicon 807 -3144 807 -3144 0 3
rlabel polysilicon 810 -3144 810 -3144 0 4
rlabel polysilicon 814 -3138 814 -3138 0 1
rlabel polysilicon 814 -3144 814 -3144 0 3
rlabel polysilicon 821 -3138 821 -3138 0 1
rlabel polysilicon 821 -3144 821 -3144 0 3
rlabel polysilicon 828 -3138 828 -3138 0 1
rlabel polysilicon 828 -3144 828 -3144 0 3
rlabel polysilicon 835 -3138 835 -3138 0 1
rlabel polysilicon 835 -3144 835 -3144 0 3
rlabel polysilicon 842 -3138 842 -3138 0 1
rlabel polysilicon 842 -3144 842 -3144 0 3
rlabel polysilicon 849 -3138 849 -3138 0 1
rlabel polysilicon 849 -3144 849 -3144 0 3
rlabel polysilicon 856 -3138 856 -3138 0 1
rlabel polysilicon 856 -3144 856 -3144 0 3
rlabel polysilicon 863 -3138 863 -3138 0 1
rlabel polysilicon 863 -3144 863 -3144 0 3
rlabel polysilicon 870 -3138 870 -3138 0 1
rlabel polysilicon 870 -3144 870 -3144 0 3
rlabel polysilicon 877 -3138 877 -3138 0 1
rlabel polysilicon 877 -3144 877 -3144 0 3
rlabel polysilicon 884 -3138 884 -3138 0 1
rlabel polysilicon 884 -3144 884 -3144 0 3
rlabel polysilicon 891 -3138 891 -3138 0 1
rlabel polysilicon 891 -3144 891 -3144 0 3
rlabel polysilicon 898 -3138 898 -3138 0 1
rlabel polysilicon 901 -3138 901 -3138 0 2
rlabel polysilicon 898 -3144 898 -3144 0 3
rlabel polysilicon 901 -3144 901 -3144 0 4
rlabel polysilicon 905 -3138 905 -3138 0 1
rlabel polysilicon 905 -3144 905 -3144 0 3
rlabel polysilicon 912 -3138 912 -3138 0 1
rlabel polysilicon 915 -3138 915 -3138 0 2
rlabel polysilicon 915 -3144 915 -3144 0 4
rlabel polysilicon 919 -3138 919 -3138 0 1
rlabel polysilicon 919 -3144 919 -3144 0 3
rlabel polysilicon 926 -3138 926 -3138 0 1
rlabel polysilicon 926 -3144 926 -3144 0 3
rlabel polysilicon 933 -3138 933 -3138 0 1
rlabel polysilicon 933 -3144 933 -3144 0 3
rlabel polysilicon 940 -3138 940 -3138 0 1
rlabel polysilicon 940 -3144 940 -3144 0 3
rlabel polysilicon 947 -3138 947 -3138 0 1
rlabel polysilicon 947 -3144 947 -3144 0 3
rlabel polysilicon 954 -3138 954 -3138 0 1
rlabel polysilicon 954 -3144 954 -3144 0 3
rlabel polysilicon 961 -3138 961 -3138 0 1
rlabel polysilicon 961 -3144 961 -3144 0 3
rlabel polysilicon 968 -3138 968 -3138 0 1
rlabel polysilicon 968 -3144 968 -3144 0 3
rlabel polysilicon 975 -3138 975 -3138 0 1
rlabel polysilicon 975 -3144 975 -3144 0 3
rlabel polysilicon 982 -3138 982 -3138 0 1
rlabel polysilicon 982 -3144 982 -3144 0 3
rlabel polysilicon 989 -3138 989 -3138 0 1
rlabel polysilicon 989 -3144 989 -3144 0 3
rlabel polysilicon 996 -3138 996 -3138 0 1
rlabel polysilicon 996 -3144 996 -3144 0 3
rlabel polysilicon 1003 -3138 1003 -3138 0 1
rlabel polysilicon 1003 -3144 1003 -3144 0 3
rlabel polysilicon 1010 -3138 1010 -3138 0 1
rlabel polysilicon 1010 -3144 1010 -3144 0 3
rlabel polysilicon 1017 -3138 1017 -3138 0 1
rlabel polysilicon 1017 -3144 1017 -3144 0 3
rlabel polysilicon 1024 -3138 1024 -3138 0 1
rlabel polysilicon 1024 -3144 1024 -3144 0 3
rlabel polysilicon 1031 -3138 1031 -3138 0 1
rlabel polysilicon 1031 -3144 1031 -3144 0 3
rlabel polysilicon 1038 -3138 1038 -3138 0 1
rlabel polysilicon 1038 -3144 1038 -3144 0 3
rlabel polysilicon 1045 -3138 1045 -3138 0 1
rlabel polysilicon 1045 -3144 1045 -3144 0 3
rlabel polysilicon 1052 -3138 1052 -3138 0 1
rlabel polysilicon 1052 -3144 1052 -3144 0 3
rlabel polysilicon 1059 -3138 1059 -3138 0 1
rlabel polysilicon 1059 -3144 1059 -3144 0 3
rlabel polysilicon 1066 -3138 1066 -3138 0 1
rlabel polysilicon 1066 -3144 1066 -3144 0 3
rlabel polysilicon 1073 -3138 1073 -3138 0 1
rlabel polysilicon 1073 -3144 1073 -3144 0 3
rlabel polysilicon 1080 -3138 1080 -3138 0 1
rlabel polysilicon 1080 -3144 1080 -3144 0 3
rlabel polysilicon 1087 -3138 1087 -3138 0 1
rlabel polysilicon 1087 -3144 1087 -3144 0 3
rlabel polysilicon 1094 -3138 1094 -3138 0 1
rlabel polysilicon 1094 -3144 1094 -3144 0 3
rlabel polysilicon 1101 -3138 1101 -3138 0 1
rlabel polysilicon 1101 -3144 1101 -3144 0 3
rlabel polysilicon 1108 -3138 1108 -3138 0 1
rlabel polysilicon 1108 -3144 1108 -3144 0 3
rlabel polysilicon 1115 -3138 1115 -3138 0 1
rlabel polysilicon 1115 -3144 1115 -3144 0 3
rlabel polysilicon 1122 -3138 1122 -3138 0 1
rlabel polysilicon 1122 -3144 1122 -3144 0 3
rlabel polysilicon 1129 -3138 1129 -3138 0 1
rlabel polysilicon 1129 -3144 1129 -3144 0 3
rlabel polysilicon 1136 -3138 1136 -3138 0 1
rlabel polysilicon 1136 -3144 1136 -3144 0 3
rlabel polysilicon 1143 -3138 1143 -3138 0 1
rlabel polysilicon 1143 -3144 1143 -3144 0 3
rlabel polysilicon 1150 -3138 1150 -3138 0 1
rlabel polysilicon 1150 -3144 1150 -3144 0 3
rlabel polysilicon 1157 -3138 1157 -3138 0 1
rlabel polysilicon 1157 -3144 1157 -3144 0 3
rlabel polysilicon 1164 -3138 1164 -3138 0 1
rlabel polysilicon 1164 -3144 1164 -3144 0 3
rlabel polysilicon 1171 -3138 1171 -3138 0 1
rlabel polysilicon 1171 -3144 1171 -3144 0 3
rlabel polysilicon 1178 -3138 1178 -3138 0 1
rlabel polysilicon 1178 -3144 1178 -3144 0 3
rlabel polysilicon 1185 -3138 1185 -3138 0 1
rlabel polysilicon 1185 -3144 1185 -3144 0 3
rlabel polysilicon 1192 -3138 1192 -3138 0 1
rlabel polysilicon 1192 -3144 1192 -3144 0 3
rlabel polysilicon 1202 -3138 1202 -3138 0 2
rlabel polysilicon 1199 -3144 1199 -3144 0 3
rlabel polysilicon 1202 -3144 1202 -3144 0 4
rlabel polysilicon 1209 -3138 1209 -3138 0 2
rlabel polysilicon 1206 -3144 1206 -3144 0 3
rlabel polysilicon 1209 -3144 1209 -3144 0 4
rlabel polysilicon 1213 -3138 1213 -3138 0 1
rlabel polysilicon 1213 -3144 1213 -3144 0 3
rlabel polysilicon 1220 -3138 1220 -3138 0 1
rlabel polysilicon 1220 -3144 1220 -3144 0 3
rlabel polysilicon 1227 -3138 1227 -3138 0 1
rlabel polysilicon 1227 -3144 1227 -3144 0 3
rlabel polysilicon 1234 -3138 1234 -3138 0 1
rlabel polysilicon 1234 -3144 1234 -3144 0 3
rlabel polysilicon 1241 -3138 1241 -3138 0 1
rlabel polysilicon 1241 -3144 1241 -3144 0 3
rlabel polysilicon 1248 -3138 1248 -3138 0 1
rlabel polysilicon 1248 -3144 1248 -3144 0 3
rlabel polysilicon 1255 -3138 1255 -3138 0 1
rlabel polysilicon 1255 -3144 1255 -3144 0 3
rlabel polysilicon 1262 -3138 1262 -3138 0 1
rlabel polysilicon 1262 -3144 1262 -3144 0 3
rlabel polysilicon 1269 -3138 1269 -3138 0 1
rlabel polysilicon 1269 -3144 1269 -3144 0 3
rlabel polysilicon 1276 -3138 1276 -3138 0 1
rlabel polysilicon 1276 -3144 1276 -3144 0 3
rlabel polysilicon 1283 -3138 1283 -3138 0 1
rlabel polysilicon 1283 -3144 1283 -3144 0 3
rlabel polysilicon 1290 -3138 1290 -3138 0 1
rlabel polysilicon 1290 -3144 1290 -3144 0 3
rlabel polysilicon 1297 -3138 1297 -3138 0 1
rlabel polysilicon 1297 -3144 1297 -3144 0 3
rlabel polysilicon 1304 -3138 1304 -3138 0 1
rlabel polysilicon 1304 -3144 1304 -3144 0 3
rlabel polysilicon 1311 -3138 1311 -3138 0 1
rlabel polysilicon 1311 -3144 1311 -3144 0 3
rlabel polysilicon 1318 -3138 1318 -3138 0 1
rlabel polysilicon 1318 -3144 1318 -3144 0 3
rlabel polysilicon 1325 -3138 1325 -3138 0 1
rlabel polysilicon 1325 -3144 1325 -3144 0 3
rlabel polysilicon 1332 -3138 1332 -3138 0 1
rlabel polysilicon 1335 -3138 1335 -3138 0 2
rlabel polysilicon 1332 -3144 1332 -3144 0 3
rlabel polysilicon 1335 -3144 1335 -3144 0 4
rlabel polysilicon 1339 -3138 1339 -3138 0 1
rlabel polysilicon 1339 -3144 1339 -3144 0 3
rlabel polysilicon 1353 -3138 1353 -3138 0 1
rlabel polysilicon 1353 -3144 1353 -3144 0 3
rlabel polysilicon 1360 -3138 1360 -3138 0 1
rlabel polysilicon 1360 -3144 1360 -3144 0 3
rlabel polysilicon 1367 -3138 1367 -3138 0 1
rlabel polysilicon 1367 -3144 1367 -3144 0 3
rlabel polysilicon 1374 -3138 1374 -3138 0 1
rlabel polysilicon 1374 -3144 1374 -3144 0 3
rlabel polysilicon 163 -3231 163 -3231 0 1
rlabel polysilicon 163 -3237 163 -3237 0 3
rlabel polysilicon 170 -3231 170 -3231 0 1
rlabel polysilicon 170 -3237 170 -3237 0 3
rlabel polysilicon 177 -3231 177 -3231 0 1
rlabel polysilicon 177 -3237 177 -3237 0 3
rlabel polysilicon 184 -3231 184 -3231 0 1
rlabel polysilicon 187 -3231 187 -3231 0 2
rlabel polysilicon 184 -3237 184 -3237 0 3
rlabel polysilicon 187 -3237 187 -3237 0 4
rlabel polysilicon 191 -3231 191 -3231 0 1
rlabel polysilicon 191 -3237 191 -3237 0 3
rlabel polysilicon 198 -3231 198 -3231 0 1
rlabel polysilicon 198 -3237 198 -3237 0 3
rlabel polysilicon 205 -3231 205 -3231 0 1
rlabel polysilicon 205 -3237 205 -3237 0 3
rlabel polysilicon 212 -3231 212 -3231 0 1
rlabel polysilicon 212 -3237 212 -3237 0 3
rlabel polysilicon 219 -3231 219 -3231 0 1
rlabel polysilicon 219 -3237 219 -3237 0 3
rlabel polysilicon 226 -3231 226 -3231 0 1
rlabel polysilicon 226 -3237 226 -3237 0 3
rlabel polysilicon 233 -3231 233 -3231 0 1
rlabel polysilicon 233 -3237 233 -3237 0 3
rlabel polysilicon 240 -3231 240 -3231 0 1
rlabel polysilicon 240 -3237 240 -3237 0 3
rlabel polysilicon 247 -3231 247 -3231 0 1
rlabel polysilicon 247 -3237 247 -3237 0 3
rlabel polysilicon 254 -3231 254 -3231 0 1
rlabel polysilicon 254 -3237 254 -3237 0 3
rlabel polysilicon 261 -3231 261 -3231 0 1
rlabel polysilicon 261 -3237 261 -3237 0 3
rlabel polysilicon 268 -3231 268 -3231 0 1
rlabel polysilicon 268 -3237 268 -3237 0 3
rlabel polysilicon 275 -3231 275 -3231 0 1
rlabel polysilicon 275 -3237 275 -3237 0 3
rlabel polysilicon 282 -3231 282 -3231 0 1
rlabel polysilicon 285 -3231 285 -3231 0 2
rlabel polysilicon 282 -3237 282 -3237 0 3
rlabel polysilicon 289 -3231 289 -3231 0 1
rlabel polysilicon 289 -3237 289 -3237 0 3
rlabel polysilicon 296 -3231 296 -3231 0 1
rlabel polysilicon 296 -3237 296 -3237 0 3
rlabel polysilicon 303 -3231 303 -3231 0 1
rlabel polysilicon 303 -3237 303 -3237 0 3
rlabel polysilicon 310 -3231 310 -3231 0 1
rlabel polysilicon 310 -3237 310 -3237 0 3
rlabel polysilicon 317 -3231 317 -3231 0 1
rlabel polysilicon 317 -3237 317 -3237 0 3
rlabel polysilicon 324 -3231 324 -3231 0 1
rlabel polysilicon 324 -3237 324 -3237 0 3
rlabel polysilicon 331 -3231 331 -3231 0 1
rlabel polysilicon 331 -3237 331 -3237 0 3
rlabel polysilicon 338 -3231 338 -3231 0 1
rlabel polysilicon 338 -3237 338 -3237 0 3
rlabel polysilicon 345 -3231 345 -3231 0 1
rlabel polysilicon 345 -3237 345 -3237 0 3
rlabel polysilicon 352 -3231 352 -3231 0 1
rlabel polysilicon 352 -3237 352 -3237 0 3
rlabel polysilicon 359 -3231 359 -3231 0 1
rlabel polysilicon 359 -3237 359 -3237 0 3
rlabel polysilicon 366 -3231 366 -3231 0 1
rlabel polysilicon 366 -3237 366 -3237 0 3
rlabel polysilicon 373 -3231 373 -3231 0 1
rlabel polysilicon 373 -3237 373 -3237 0 3
rlabel polysilicon 380 -3231 380 -3231 0 1
rlabel polysilicon 380 -3237 380 -3237 0 3
rlabel polysilicon 387 -3231 387 -3231 0 1
rlabel polysilicon 387 -3237 387 -3237 0 3
rlabel polysilicon 394 -3231 394 -3231 0 1
rlabel polysilicon 394 -3237 394 -3237 0 3
rlabel polysilicon 401 -3231 401 -3231 0 1
rlabel polysilicon 401 -3237 401 -3237 0 3
rlabel polysilicon 408 -3231 408 -3231 0 1
rlabel polysilicon 408 -3237 408 -3237 0 3
rlabel polysilicon 415 -3231 415 -3231 0 1
rlabel polysilicon 415 -3237 415 -3237 0 3
rlabel polysilicon 422 -3231 422 -3231 0 1
rlabel polysilicon 422 -3237 422 -3237 0 3
rlabel polysilicon 429 -3231 429 -3231 0 1
rlabel polysilicon 429 -3237 429 -3237 0 3
rlabel polysilicon 436 -3231 436 -3231 0 1
rlabel polysilicon 436 -3237 436 -3237 0 3
rlabel polysilicon 443 -3231 443 -3231 0 1
rlabel polysilicon 443 -3237 443 -3237 0 3
rlabel polysilicon 450 -3231 450 -3231 0 1
rlabel polysilicon 450 -3237 450 -3237 0 3
rlabel polysilicon 457 -3231 457 -3231 0 1
rlabel polysilicon 460 -3231 460 -3231 0 2
rlabel polysilicon 457 -3237 457 -3237 0 3
rlabel polysilicon 460 -3237 460 -3237 0 4
rlabel polysilicon 464 -3231 464 -3231 0 1
rlabel polysilicon 464 -3237 464 -3237 0 3
rlabel polysilicon 471 -3231 471 -3231 0 1
rlabel polysilicon 471 -3237 471 -3237 0 3
rlabel polysilicon 478 -3231 478 -3231 0 1
rlabel polysilicon 478 -3237 478 -3237 0 3
rlabel polysilicon 481 -3237 481 -3237 0 4
rlabel polysilicon 485 -3231 485 -3231 0 1
rlabel polysilicon 485 -3237 485 -3237 0 3
rlabel polysilicon 492 -3231 492 -3231 0 1
rlabel polysilicon 492 -3237 492 -3237 0 3
rlabel polysilicon 499 -3231 499 -3231 0 1
rlabel polysilicon 499 -3237 499 -3237 0 3
rlabel polysilicon 506 -3231 506 -3231 0 1
rlabel polysilicon 506 -3237 506 -3237 0 3
rlabel polysilicon 513 -3231 513 -3231 0 1
rlabel polysilicon 513 -3237 513 -3237 0 3
rlabel polysilicon 520 -3231 520 -3231 0 1
rlabel polysilicon 520 -3237 520 -3237 0 3
rlabel polysilicon 527 -3231 527 -3231 0 1
rlabel polysilicon 527 -3237 527 -3237 0 3
rlabel polysilicon 534 -3231 534 -3231 0 1
rlabel polysilicon 534 -3237 534 -3237 0 3
rlabel polysilicon 544 -3231 544 -3231 0 2
rlabel polysilicon 541 -3237 541 -3237 0 3
rlabel polysilicon 544 -3237 544 -3237 0 4
rlabel polysilicon 548 -3231 548 -3231 0 1
rlabel polysilicon 548 -3237 548 -3237 0 3
rlabel polysilicon 555 -3231 555 -3231 0 1
rlabel polysilicon 555 -3237 555 -3237 0 3
rlabel polysilicon 562 -3231 562 -3231 0 1
rlabel polysilicon 562 -3237 562 -3237 0 3
rlabel polysilicon 569 -3231 569 -3231 0 1
rlabel polysilicon 569 -3237 569 -3237 0 3
rlabel polysilicon 576 -3231 576 -3231 0 1
rlabel polysilicon 579 -3237 579 -3237 0 4
rlabel polysilicon 583 -3231 583 -3231 0 1
rlabel polysilicon 583 -3237 583 -3237 0 3
rlabel polysilicon 590 -3231 590 -3231 0 1
rlabel polysilicon 590 -3237 590 -3237 0 3
rlabel polysilicon 597 -3231 597 -3231 0 1
rlabel polysilicon 597 -3237 597 -3237 0 3
rlabel polysilicon 604 -3231 604 -3231 0 1
rlabel polysilicon 604 -3237 604 -3237 0 3
rlabel polysilicon 611 -3231 611 -3231 0 1
rlabel polysilicon 611 -3237 611 -3237 0 3
rlabel polysilicon 618 -3231 618 -3231 0 1
rlabel polysilicon 618 -3237 618 -3237 0 3
rlabel polysilicon 625 -3231 625 -3231 0 1
rlabel polysilicon 625 -3237 625 -3237 0 3
rlabel polysilicon 632 -3231 632 -3231 0 1
rlabel polysilicon 635 -3231 635 -3231 0 2
rlabel polysilicon 639 -3231 639 -3231 0 1
rlabel polysilicon 639 -3237 639 -3237 0 3
rlabel polysilicon 646 -3231 646 -3231 0 1
rlabel polysilicon 646 -3237 646 -3237 0 3
rlabel polysilicon 653 -3231 653 -3231 0 1
rlabel polysilicon 653 -3237 653 -3237 0 3
rlabel polysilicon 660 -3231 660 -3231 0 1
rlabel polysilicon 660 -3237 660 -3237 0 3
rlabel polysilicon 667 -3231 667 -3231 0 1
rlabel polysilicon 667 -3237 667 -3237 0 3
rlabel polysilicon 674 -3231 674 -3231 0 1
rlabel polysilicon 674 -3237 674 -3237 0 3
rlabel polysilicon 681 -3231 681 -3231 0 1
rlabel polysilicon 681 -3237 681 -3237 0 3
rlabel polysilicon 688 -3231 688 -3231 0 1
rlabel polysilicon 688 -3237 688 -3237 0 3
rlabel polysilicon 695 -3231 695 -3231 0 1
rlabel polysilicon 695 -3237 695 -3237 0 3
rlabel polysilicon 702 -3231 702 -3231 0 1
rlabel polysilicon 702 -3237 702 -3237 0 3
rlabel polysilicon 709 -3231 709 -3231 0 1
rlabel polysilicon 709 -3237 709 -3237 0 3
rlabel polysilicon 712 -3237 712 -3237 0 4
rlabel polysilicon 716 -3231 716 -3231 0 1
rlabel polysilicon 716 -3237 716 -3237 0 3
rlabel polysilicon 723 -3231 723 -3231 0 1
rlabel polysilicon 723 -3237 723 -3237 0 3
rlabel polysilicon 730 -3231 730 -3231 0 1
rlabel polysilicon 730 -3237 730 -3237 0 3
rlabel polysilicon 737 -3231 737 -3231 0 1
rlabel polysilicon 737 -3237 737 -3237 0 3
rlabel polysilicon 744 -3231 744 -3231 0 1
rlabel polysilicon 747 -3231 747 -3231 0 2
rlabel polysilicon 744 -3237 744 -3237 0 3
rlabel polysilicon 747 -3237 747 -3237 0 4
rlabel polysilicon 751 -3231 751 -3231 0 1
rlabel polysilicon 754 -3231 754 -3231 0 2
rlabel polysilicon 751 -3237 751 -3237 0 3
rlabel polysilicon 754 -3237 754 -3237 0 4
rlabel polysilicon 758 -3231 758 -3231 0 1
rlabel polysilicon 758 -3237 758 -3237 0 3
rlabel polysilicon 765 -3231 765 -3231 0 1
rlabel polysilicon 768 -3231 768 -3231 0 2
rlabel polysilicon 768 -3237 768 -3237 0 4
rlabel polysilicon 772 -3231 772 -3231 0 1
rlabel polysilicon 772 -3237 772 -3237 0 3
rlabel polysilicon 779 -3231 779 -3231 0 1
rlabel polysilicon 779 -3237 779 -3237 0 3
rlabel polysilicon 786 -3231 786 -3231 0 1
rlabel polysilicon 786 -3237 786 -3237 0 3
rlabel polysilicon 793 -3231 793 -3231 0 1
rlabel polysilicon 793 -3237 793 -3237 0 3
rlabel polysilicon 800 -3231 800 -3231 0 1
rlabel polysilicon 800 -3237 800 -3237 0 3
rlabel polysilicon 807 -3231 807 -3231 0 1
rlabel polysilicon 810 -3231 810 -3231 0 2
rlabel polysilicon 807 -3237 807 -3237 0 3
rlabel polysilicon 810 -3237 810 -3237 0 4
rlabel polysilicon 814 -3231 814 -3231 0 1
rlabel polysilicon 814 -3237 814 -3237 0 3
rlabel polysilicon 821 -3231 821 -3231 0 1
rlabel polysilicon 821 -3237 821 -3237 0 3
rlabel polysilicon 828 -3231 828 -3231 0 1
rlabel polysilicon 828 -3237 828 -3237 0 3
rlabel polysilicon 835 -3231 835 -3231 0 1
rlabel polysilicon 835 -3237 835 -3237 0 3
rlabel polysilicon 842 -3231 842 -3231 0 1
rlabel polysilicon 842 -3237 842 -3237 0 3
rlabel polysilicon 849 -3231 849 -3231 0 1
rlabel polysilicon 849 -3237 849 -3237 0 3
rlabel polysilicon 856 -3231 856 -3231 0 1
rlabel polysilicon 856 -3237 856 -3237 0 3
rlabel polysilicon 863 -3231 863 -3231 0 1
rlabel polysilicon 863 -3237 863 -3237 0 3
rlabel polysilicon 870 -3231 870 -3231 0 1
rlabel polysilicon 870 -3237 870 -3237 0 3
rlabel polysilicon 877 -3231 877 -3231 0 1
rlabel polysilicon 877 -3237 877 -3237 0 3
rlabel polysilicon 884 -3231 884 -3231 0 1
rlabel polysilicon 884 -3237 884 -3237 0 3
rlabel polysilicon 891 -3231 891 -3231 0 1
rlabel polysilicon 894 -3231 894 -3231 0 2
rlabel polysilicon 891 -3237 891 -3237 0 3
rlabel polysilicon 898 -3231 898 -3231 0 1
rlabel polysilicon 898 -3237 898 -3237 0 3
rlabel polysilicon 905 -3231 905 -3231 0 1
rlabel polysilicon 905 -3237 905 -3237 0 3
rlabel polysilicon 912 -3231 912 -3231 0 1
rlabel polysilicon 912 -3237 912 -3237 0 3
rlabel polysilicon 919 -3231 919 -3231 0 1
rlabel polysilicon 919 -3237 919 -3237 0 3
rlabel polysilicon 926 -3231 926 -3231 0 1
rlabel polysilicon 926 -3237 926 -3237 0 3
rlabel polysilicon 933 -3231 933 -3231 0 1
rlabel polysilicon 933 -3237 933 -3237 0 3
rlabel polysilicon 940 -3231 940 -3231 0 1
rlabel polysilicon 943 -3231 943 -3231 0 2
rlabel polysilicon 940 -3237 940 -3237 0 3
rlabel polysilicon 947 -3231 947 -3231 0 1
rlabel polysilicon 947 -3237 947 -3237 0 3
rlabel polysilicon 954 -3231 954 -3231 0 1
rlabel polysilicon 954 -3237 954 -3237 0 3
rlabel polysilicon 961 -3231 961 -3231 0 1
rlabel polysilicon 961 -3237 961 -3237 0 3
rlabel polysilicon 964 -3237 964 -3237 0 4
rlabel polysilicon 968 -3231 968 -3231 0 1
rlabel polysilicon 968 -3237 968 -3237 0 3
rlabel polysilicon 975 -3231 975 -3231 0 1
rlabel polysilicon 975 -3237 975 -3237 0 3
rlabel polysilicon 982 -3231 982 -3231 0 1
rlabel polysilicon 982 -3237 982 -3237 0 3
rlabel polysilicon 989 -3231 989 -3231 0 1
rlabel polysilicon 989 -3237 989 -3237 0 3
rlabel polysilicon 996 -3231 996 -3231 0 1
rlabel polysilicon 996 -3237 996 -3237 0 3
rlabel polysilicon 1003 -3231 1003 -3231 0 1
rlabel polysilicon 1003 -3237 1003 -3237 0 3
rlabel polysilicon 1010 -3231 1010 -3231 0 1
rlabel polysilicon 1010 -3237 1010 -3237 0 3
rlabel polysilicon 1017 -3231 1017 -3231 0 1
rlabel polysilicon 1017 -3237 1017 -3237 0 3
rlabel polysilicon 1024 -3231 1024 -3231 0 1
rlabel polysilicon 1024 -3237 1024 -3237 0 3
rlabel polysilicon 1031 -3231 1031 -3231 0 1
rlabel polysilicon 1031 -3237 1031 -3237 0 3
rlabel polysilicon 1038 -3231 1038 -3231 0 1
rlabel polysilicon 1038 -3237 1038 -3237 0 3
rlabel polysilicon 1045 -3231 1045 -3231 0 1
rlabel polysilicon 1045 -3237 1045 -3237 0 3
rlabel polysilicon 1052 -3231 1052 -3231 0 1
rlabel polysilicon 1052 -3237 1052 -3237 0 3
rlabel polysilicon 1059 -3231 1059 -3231 0 1
rlabel polysilicon 1059 -3237 1059 -3237 0 3
rlabel polysilicon 1066 -3231 1066 -3231 0 1
rlabel polysilicon 1066 -3237 1066 -3237 0 3
rlabel polysilicon 1073 -3231 1073 -3231 0 1
rlabel polysilicon 1073 -3237 1073 -3237 0 3
rlabel polysilicon 1080 -3231 1080 -3231 0 1
rlabel polysilicon 1080 -3237 1080 -3237 0 3
rlabel polysilicon 1087 -3231 1087 -3231 0 1
rlabel polysilicon 1087 -3237 1087 -3237 0 3
rlabel polysilicon 1094 -3231 1094 -3231 0 1
rlabel polysilicon 1094 -3237 1094 -3237 0 3
rlabel polysilicon 1101 -3231 1101 -3231 0 1
rlabel polysilicon 1101 -3237 1101 -3237 0 3
rlabel polysilicon 1108 -3231 1108 -3231 0 1
rlabel polysilicon 1108 -3237 1108 -3237 0 3
rlabel polysilicon 1115 -3231 1115 -3231 0 1
rlabel polysilicon 1115 -3237 1115 -3237 0 3
rlabel polysilicon 1122 -3231 1122 -3231 0 1
rlabel polysilicon 1122 -3237 1122 -3237 0 3
rlabel polysilicon 1129 -3231 1129 -3231 0 1
rlabel polysilicon 1129 -3237 1129 -3237 0 3
rlabel polysilicon 1136 -3231 1136 -3231 0 1
rlabel polysilicon 1136 -3237 1136 -3237 0 3
rlabel polysilicon 1143 -3231 1143 -3231 0 1
rlabel polysilicon 1143 -3237 1143 -3237 0 3
rlabel polysilicon 1150 -3231 1150 -3231 0 1
rlabel polysilicon 1150 -3237 1150 -3237 0 3
rlabel polysilicon 1157 -3231 1157 -3231 0 1
rlabel polysilicon 1157 -3237 1157 -3237 0 3
rlabel polysilicon 1164 -3231 1164 -3231 0 1
rlabel polysilicon 1167 -3231 1167 -3231 0 2
rlabel polysilicon 1164 -3237 1164 -3237 0 3
rlabel polysilicon 1171 -3231 1171 -3231 0 1
rlabel polysilicon 1171 -3237 1171 -3237 0 3
rlabel polysilicon 1178 -3231 1178 -3231 0 1
rlabel polysilicon 1178 -3237 1178 -3237 0 3
rlabel polysilicon 1185 -3231 1185 -3231 0 1
rlabel polysilicon 1185 -3237 1185 -3237 0 3
rlabel polysilicon 1192 -3231 1192 -3231 0 1
rlabel polysilicon 1192 -3237 1192 -3237 0 3
rlabel polysilicon 1199 -3231 1199 -3231 0 1
rlabel polysilicon 1202 -3231 1202 -3231 0 2
rlabel polysilicon 1202 -3237 1202 -3237 0 4
rlabel polysilicon 1206 -3231 1206 -3231 0 1
rlabel polysilicon 1206 -3237 1206 -3237 0 3
rlabel polysilicon 1213 -3231 1213 -3231 0 1
rlabel polysilicon 1213 -3237 1213 -3237 0 3
rlabel polysilicon 1220 -3231 1220 -3231 0 1
rlabel polysilicon 1220 -3237 1220 -3237 0 3
rlabel polysilicon 1230 -3231 1230 -3231 0 2
rlabel polysilicon 1227 -3237 1227 -3237 0 3
rlabel polysilicon 1234 -3231 1234 -3231 0 1
rlabel polysilicon 1234 -3237 1234 -3237 0 3
rlabel polysilicon 1241 -3231 1241 -3231 0 1
rlabel polysilicon 1241 -3237 1241 -3237 0 3
rlabel polysilicon 1248 -3231 1248 -3231 0 1
rlabel polysilicon 1248 -3237 1248 -3237 0 3
rlabel polysilicon 1255 -3231 1255 -3231 0 1
rlabel polysilicon 1255 -3237 1255 -3237 0 3
rlabel polysilicon 1258 -3237 1258 -3237 0 4
rlabel polysilicon 1262 -3231 1262 -3231 0 1
rlabel polysilicon 1262 -3237 1262 -3237 0 3
rlabel polysilicon 1269 -3231 1269 -3231 0 1
rlabel polysilicon 1269 -3237 1269 -3237 0 3
rlabel polysilicon 1276 -3231 1276 -3231 0 1
rlabel polysilicon 1276 -3237 1276 -3237 0 3
rlabel polysilicon 1283 -3231 1283 -3231 0 1
rlabel polysilicon 1286 -3231 1286 -3231 0 2
rlabel polysilicon 1283 -3237 1283 -3237 0 3
rlabel polysilicon 1290 -3231 1290 -3231 0 1
rlabel polysilicon 1293 -3231 1293 -3231 0 2
rlabel polysilicon 1293 -3237 1293 -3237 0 4
rlabel polysilicon 1297 -3231 1297 -3231 0 1
rlabel polysilicon 1297 -3237 1297 -3237 0 3
rlabel polysilicon 1304 -3231 1304 -3231 0 1
rlabel polysilicon 1304 -3237 1304 -3237 0 3
rlabel polysilicon 1346 -3231 1346 -3231 0 1
rlabel polysilicon 1346 -3237 1346 -3237 0 3
rlabel polysilicon 1353 -3231 1353 -3231 0 1
rlabel polysilicon 1353 -3237 1353 -3237 0 3
rlabel polysilicon 1360 -3231 1360 -3231 0 1
rlabel polysilicon 1360 -3237 1360 -3237 0 3
rlabel polysilicon 156 -3308 156 -3308 0 1
rlabel polysilicon 156 -3314 156 -3314 0 3
rlabel polysilicon 163 -3308 163 -3308 0 1
rlabel polysilicon 163 -3314 163 -3314 0 3
rlabel polysilicon 170 -3308 170 -3308 0 1
rlabel polysilicon 170 -3314 170 -3314 0 3
rlabel polysilicon 177 -3308 177 -3308 0 1
rlabel polysilicon 177 -3314 177 -3314 0 3
rlabel polysilicon 184 -3308 184 -3308 0 1
rlabel polysilicon 184 -3314 184 -3314 0 3
rlabel polysilicon 191 -3308 191 -3308 0 1
rlabel polysilicon 191 -3314 191 -3314 0 3
rlabel polysilicon 198 -3308 198 -3308 0 1
rlabel polysilicon 201 -3308 201 -3308 0 2
rlabel polysilicon 205 -3308 205 -3308 0 1
rlabel polysilicon 205 -3314 205 -3314 0 3
rlabel polysilicon 212 -3308 212 -3308 0 1
rlabel polysilicon 212 -3314 212 -3314 0 3
rlabel polysilicon 219 -3308 219 -3308 0 1
rlabel polysilicon 219 -3314 219 -3314 0 3
rlabel polysilicon 226 -3308 226 -3308 0 1
rlabel polysilicon 226 -3314 226 -3314 0 3
rlabel polysilicon 233 -3308 233 -3308 0 1
rlabel polysilicon 233 -3314 233 -3314 0 3
rlabel polysilicon 243 -3308 243 -3308 0 2
rlabel polysilicon 243 -3314 243 -3314 0 4
rlabel polysilicon 247 -3308 247 -3308 0 1
rlabel polysilicon 247 -3314 247 -3314 0 3
rlabel polysilicon 254 -3308 254 -3308 0 1
rlabel polysilicon 254 -3314 254 -3314 0 3
rlabel polysilicon 261 -3308 261 -3308 0 1
rlabel polysilicon 261 -3314 261 -3314 0 3
rlabel polysilicon 268 -3308 268 -3308 0 1
rlabel polysilicon 268 -3314 268 -3314 0 3
rlabel polysilicon 275 -3308 275 -3308 0 1
rlabel polysilicon 275 -3314 275 -3314 0 3
rlabel polysilicon 282 -3308 282 -3308 0 1
rlabel polysilicon 282 -3314 282 -3314 0 3
rlabel polysilicon 289 -3308 289 -3308 0 1
rlabel polysilicon 289 -3314 289 -3314 0 3
rlabel polysilicon 296 -3308 296 -3308 0 1
rlabel polysilicon 296 -3314 296 -3314 0 3
rlabel polysilicon 303 -3308 303 -3308 0 1
rlabel polysilicon 303 -3314 303 -3314 0 3
rlabel polysilicon 310 -3308 310 -3308 0 1
rlabel polysilicon 310 -3314 310 -3314 0 3
rlabel polysilicon 317 -3308 317 -3308 0 1
rlabel polysilicon 317 -3314 317 -3314 0 3
rlabel polysilicon 324 -3308 324 -3308 0 1
rlabel polysilicon 324 -3314 324 -3314 0 3
rlabel polysilicon 331 -3308 331 -3308 0 1
rlabel polysilicon 331 -3314 331 -3314 0 3
rlabel polysilicon 338 -3308 338 -3308 0 1
rlabel polysilicon 338 -3314 338 -3314 0 3
rlabel polysilicon 345 -3308 345 -3308 0 1
rlabel polysilicon 345 -3314 345 -3314 0 3
rlabel polysilicon 352 -3308 352 -3308 0 1
rlabel polysilicon 352 -3314 352 -3314 0 3
rlabel polysilicon 359 -3308 359 -3308 0 1
rlabel polysilicon 359 -3314 359 -3314 0 3
rlabel polysilicon 366 -3308 366 -3308 0 1
rlabel polysilicon 366 -3314 366 -3314 0 3
rlabel polysilicon 373 -3308 373 -3308 0 1
rlabel polysilicon 373 -3314 373 -3314 0 3
rlabel polysilicon 380 -3308 380 -3308 0 1
rlabel polysilicon 380 -3314 380 -3314 0 3
rlabel polysilicon 387 -3308 387 -3308 0 1
rlabel polysilicon 387 -3314 387 -3314 0 3
rlabel polysilicon 394 -3308 394 -3308 0 1
rlabel polysilicon 394 -3314 394 -3314 0 3
rlabel polysilicon 401 -3308 401 -3308 0 1
rlabel polysilicon 401 -3314 401 -3314 0 3
rlabel polysilicon 408 -3308 408 -3308 0 1
rlabel polysilicon 408 -3314 408 -3314 0 3
rlabel polysilicon 415 -3308 415 -3308 0 1
rlabel polysilicon 415 -3314 415 -3314 0 3
rlabel polysilicon 422 -3308 422 -3308 0 1
rlabel polysilicon 422 -3314 422 -3314 0 3
rlabel polysilicon 429 -3308 429 -3308 0 1
rlabel polysilicon 429 -3314 429 -3314 0 3
rlabel polysilicon 436 -3308 436 -3308 0 1
rlabel polysilicon 436 -3314 436 -3314 0 3
rlabel polysilicon 443 -3308 443 -3308 0 1
rlabel polysilicon 443 -3314 443 -3314 0 3
rlabel polysilicon 450 -3308 450 -3308 0 1
rlabel polysilicon 450 -3314 450 -3314 0 3
rlabel polysilicon 457 -3308 457 -3308 0 1
rlabel polysilicon 457 -3314 457 -3314 0 3
rlabel polysilicon 464 -3308 464 -3308 0 1
rlabel polysilicon 464 -3314 464 -3314 0 3
rlabel polysilicon 471 -3308 471 -3308 0 1
rlabel polysilicon 471 -3314 471 -3314 0 3
rlabel polysilicon 478 -3308 478 -3308 0 1
rlabel polysilicon 478 -3314 478 -3314 0 3
rlabel polysilicon 485 -3308 485 -3308 0 1
rlabel polysilicon 488 -3308 488 -3308 0 2
rlabel polysilicon 485 -3314 485 -3314 0 3
rlabel polysilicon 492 -3308 492 -3308 0 1
rlabel polysilicon 492 -3314 492 -3314 0 3
rlabel polysilicon 499 -3308 499 -3308 0 1
rlabel polysilicon 499 -3314 499 -3314 0 3
rlabel polysilicon 506 -3308 506 -3308 0 1
rlabel polysilicon 506 -3314 506 -3314 0 3
rlabel polysilicon 513 -3308 513 -3308 0 1
rlabel polysilicon 513 -3314 513 -3314 0 3
rlabel polysilicon 520 -3308 520 -3308 0 1
rlabel polysilicon 520 -3314 520 -3314 0 3
rlabel polysilicon 527 -3308 527 -3308 0 1
rlabel polysilicon 527 -3314 527 -3314 0 3
rlabel polysilicon 537 -3308 537 -3308 0 2
rlabel polysilicon 534 -3314 534 -3314 0 3
rlabel polysilicon 537 -3314 537 -3314 0 4
rlabel polysilicon 541 -3308 541 -3308 0 1
rlabel polysilicon 541 -3314 541 -3314 0 3
rlabel polysilicon 548 -3308 548 -3308 0 1
rlabel polysilicon 548 -3314 548 -3314 0 3
rlabel polysilicon 555 -3308 555 -3308 0 1
rlabel polysilicon 555 -3314 555 -3314 0 3
rlabel polysilicon 562 -3308 562 -3308 0 1
rlabel polysilicon 562 -3314 562 -3314 0 3
rlabel polysilicon 569 -3308 569 -3308 0 1
rlabel polysilicon 569 -3314 569 -3314 0 3
rlabel polysilicon 576 -3308 576 -3308 0 1
rlabel polysilicon 576 -3314 576 -3314 0 3
rlabel polysilicon 583 -3308 583 -3308 0 1
rlabel polysilicon 583 -3314 583 -3314 0 3
rlabel polysilicon 590 -3308 590 -3308 0 1
rlabel polysilicon 590 -3314 590 -3314 0 3
rlabel polysilicon 597 -3308 597 -3308 0 1
rlabel polysilicon 597 -3314 597 -3314 0 3
rlabel polysilicon 604 -3308 604 -3308 0 1
rlabel polysilicon 604 -3314 604 -3314 0 3
rlabel polysilicon 611 -3308 611 -3308 0 1
rlabel polysilicon 614 -3308 614 -3308 0 2
rlabel polysilicon 614 -3314 614 -3314 0 4
rlabel polysilicon 618 -3308 618 -3308 0 1
rlabel polysilicon 618 -3314 618 -3314 0 3
rlabel polysilicon 625 -3308 625 -3308 0 1
rlabel polysilicon 625 -3314 625 -3314 0 3
rlabel polysilicon 632 -3308 632 -3308 0 1
rlabel polysilicon 632 -3314 632 -3314 0 3
rlabel polysilicon 639 -3308 639 -3308 0 1
rlabel polysilicon 639 -3314 639 -3314 0 3
rlabel polysilicon 646 -3308 646 -3308 0 1
rlabel polysilicon 646 -3314 646 -3314 0 3
rlabel polysilicon 653 -3308 653 -3308 0 1
rlabel polysilicon 656 -3308 656 -3308 0 2
rlabel polysilicon 653 -3314 653 -3314 0 3
rlabel polysilicon 656 -3314 656 -3314 0 4
rlabel polysilicon 660 -3308 660 -3308 0 1
rlabel polysilicon 663 -3308 663 -3308 0 2
rlabel polysilicon 660 -3314 660 -3314 0 3
rlabel polysilicon 663 -3314 663 -3314 0 4
rlabel polysilicon 667 -3308 667 -3308 0 1
rlabel polysilicon 670 -3308 670 -3308 0 2
rlabel polysilicon 667 -3314 667 -3314 0 3
rlabel polysilicon 670 -3314 670 -3314 0 4
rlabel polysilicon 674 -3308 674 -3308 0 1
rlabel polysilicon 674 -3314 674 -3314 0 3
rlabel polysilicon 681 -3308 681 -3308 0 1
rlabel polysilicon 681 -3314 681 -3314 0 3
rlabel polysilicon 688 -3308 688 -3308 0 1
rlabel polysilicon 691 -3308 691 -3308 0 2
rlabel polysilicon 688 -3314 688 -3314 0 3
rlabel polysilicon 691 -3314 691 -3314 0 4
rlabel polysilicon 695 -3308 695 -3308 0 1
rlabel polysilicon 695 -3314 695 -3314 0 3
rlabel polysilicon 702 -3308 702 -3308 0 1
rlabel polysilicon 702 -3314 702 -3314 0 3
rlabel polysilicon 709 -3308 709 -3308 0 1
rlabel polysilicon 709 -3314 709 -3314 0 3
rlabel polysilicon 716 -3308 716 -3308 0 1
rlabel polysilicon 716 -3314 716 -3314 0 3
rlabel polysilicon 723 -3308 723 -3308 0 1
rlabel polysilicon 723 -3314 723 -3314 0 3
rlabel polysilicon 733 -3308 733 -3308 0 2
rlabel polysilicon 730 -3314 730 -3314 0 3
rlabel polysilicon 737 -3308 737 -3308 0 1
rlabel polysilicon 737 -3314 737 -3314 0 3
rlabel polysilicon 744 -3308 744 -3308 0 1
rlabel polysilicon 744 -3314 744 -3314 0 3
rlabel polysilicon 751 -3308 751 -3308 0 1
rlabel polysilicon 751 -3314 751 -3314 0 3
rlabel polysilicon 758 -3308 758 -3308 0 1
rlabel polysilicon 758 -3314 758 -3314 0 3
rlabel polysilicon 761 -3314 761 -3314 0 4
rlabel polysilicon 765 -3308 765 -3308 0 1
rlabel polysilicon 765 -3314 765 -3314 0 3
rlabel polysilicon 772 -3308 772 -3308 0 1
rlabel polysilicon 772 -3314 772 -3314 0 3
rlabel polysilicon 779 -3308 779 -3308 0 1
rlabel polysilicon 779 -3314 779 -3314 0 3
rlabel polysilicon 786 -3308 786 -3308 0 1
rlabel polysilicon 786 -3314 786 -3314 0 3
rlabel polysilicon 793 -3308 793 -3308 0 1
rlabel polysilicon 793 -3314 793 -3314 0 3
rlabel polysilicon 800 -3308 800 -3308 0 1
rlabel polysilicon 800 -3314 800 -3314 0 3
rlabel polysilicon 807 -3308 807 -3308 0 1
rlabel polysilicon 807 -3314 807 -3314 0 3
rlabel polysilicon 814 -3308 814 -3308 0 1
rlabel polysilicon 814 -3314 814 -3314 0 3
rlabel polysilicon 821 -3308 821 -3308 0 1
rlabel polysilicon 824 -3308 824 -3308 0 2
rlabel polysilicon 824 -3314 824 -3314 0 4
rlabel polysilicon 828 -3308 828 -3308 0 1
rlabel polysilicon 828 -3314 828 -3314 0 3
rlabel polysilicon 838 -3308 838 -3308 0 2
rlabel polysilicon 835 -3314 835 -3314 0 3
rlabel polysilicon 838 -3314 838 -3314 0 4
rlabel polysilicon 842 -3308 842 -3308 0 1
rlabel polysilicon 842 -3314 842 -3314 0 3
rlabel polysilicon 849 -3308 849 -3308 0 1
rlabel polysilicon 849 -3314 849 -3314 0 3
rlabel polysilicon 859 -3308 859 -3308 0 2
rlabel polysilicon 856 -3314 856 -3314 0 3
rlabel polysilicon 859 -3314 859 -3314 0 4
rlabel polysilicon 863 -3308 863 -3308 0 1
rlabel polysilicon 863 -3314 863 -3314 0 3
rlabel polysilicon 873 -3308 873 -3308 0 2
rlabel polysilicon 870 -3314 870 -3314 0 3
rlabel polysilicon 873 -3314 873 -3314 0 4
rlabel polysilicon 877 -3308 877 -3308 0 1
rlabel polysilicon 877 -3314 877 -3314 0 3
rlabel polysilicon 884 -3308 884 -3308 0 1
rlabel polysilicon 884 -3314 884 -3314 0 3
rlabel polysilicon 891 -3308 891 -3308 0 1
rlabel polysilicon 894 -3308 894 -3308 0 2
rlabel polysilicon 891 -3314 891 -3314 0 3
rlabel polysilicon 894 -3314 894 -3314 0 4
rlabel polysilicon 898 -3308 898 -3308 0 1
rlabel polysilicon 898 -3314 898 -3314 0 3
rlabel polysilicon 905 -3308 905 -3308 0 1
rlabel polysilicon 905 -3314 905 -3314 0 3
rlabel polysilicon 912 -3308 912 -3308 0 1
rlabel polysilicon 912 -3314 912 -3314 0 3
rlabel polysilicon 919 -3308 919 -3308 0 1
rlabel polysilicon 919 -3314 919 -3314 0 3
rlabel polysilicon 926 -3308 926 -3308 0 1
rlabel polysilicon 926 -3314 926 -3314 0 3
rlabel polysilicon 933 -3308 933 -3308 0 1
rlabel polysilicon 933 -3314 933 -3314 0 3
rlabel polysilicon 940 -3308 940 -3308 0 1
rlabel polysilicon 940 -3314 940 -3314 0 3
rlabel polysilicon 947 -3308 947 -3308 0 1
rlabel polysilicon 947 -3314 947 -3314 0 3
rlabel polysilicon 954 -3308 954 -3308 0 1
rlabel polysilicon 954 -3314 954 -3314 0 3
rlabel polysilicon 961 -3308 961 -3308 0 1
rlabel polysilicon 961 -3314 961 -3314 0 3
rlabel polysilicon 968 -3308 968 -3308 0 1
rlabel polysilicon 968 -3314 968 -3314 0 3
rlabel polysilicon 975 -3308 975 -3308 0 1
rlabel polysilicon 975 -3314 975 -3314 0 3
rlabel polysilicon 982 -3308 982 -3308 0 1
rlabel polysilicon 982 -3314 982 -3314 0 3
rlabel polysilicon 989 -3308 989 -3308 0 1
rlabel polysilicon 989 -3314 989 -3314 0 3
rlabel polysilicon 996 -3308 996 -3308 0 1
rlabel polysilicon 996 -3314 996 -3314 0 3
rlabel polysilicon 1003 -3308 1003 -3308 0 1
rlabel polysilicon 1006 -3308 1006 -3308 0 2
rlabel polysilicon 1003 -3314 1003 -3314 0 3
rlabel polysilicon 1010 -3308 1010 -3308 0 1
rlabel polysilicon 1010 -3314 1010 -3314 0 3
rlabel polysilicon 1017 -3308 1017 -3308 0 1
rlabel polysilicon 1017 -3314 1017 -3314 0 3
rlabel polysilicon 1024 -3308 1024 -3308 0 1
rlabel polysilicon 1027 -3308 1027 -3308 0 2
rlabel polysilicon 1027 -3314 1027 -3314 0 4
rlabel polysilicon 1031 -3308 1031 -3308 0 1
rlabel polysilicon 1031 -3314 1031 -3314 0 3
rlabel polysilicon 1038 -3308 1038 -3308 0 1
rlabel polysilicon 1038 -3314 1038 -3314 0 3
rlabel polysilicon 1045 -3308 1045 -3308 0 1
rlabel polysilicon 1045 -3314 1045 -3314 0 3
rlabel polysilicon 1052 -3308 1052 -3308 0 1
rlabel polysilicon 1052 -3314 1052 -3314 0 3
rlabel polysilicon 1059 -3308 1059 -3308 0 1
rlabel polysilicon 1059 -3314 1059 -3314 0 3
rlabel polysilicon 1066 -3308 1066 -3308 0 1
rlabel polysilicon 1066 -3314 1066 -3314 0 3
rlabel polysilicon 1073 -3308 1073 -3308 0 1
rlabel polysilicon 1073 -3314 1073 -3314 0 3
rlabel polysilicon 1080 -3308 1080 -3308 0 1
rlabel polysilicon 1080 -3314 1080 -3314 0 3
rlabel polysilicon 1087 -3308 1087 -3308 0 1
rlabel polysilicon 1087 -3314 1087 -3314 0 3
rlabel polysilicon 1094 -3308 1094 -3308 0 1
rlabel polysilicon 1094 -3314 1094 -3314 0 3
rlabel polysilicon 1101 -3308 1101 -3308 0 1
rlabel polysilicon 1101 -3314 1101 -3314 0 3
rlabel polysilicon 1108 -3308 1108 -3308 0 1
rlabel polysilicon 1108 -3314 1108 -3314 0 3
rlabel polysilicon 1115 -3308 1115 -3308 0 1
rlabel polysilicon 1115 -3314 1115 -3314 0 3
rlabel polysilicon 1122 -3308 1122 -3308 0 1
rlabel polysilicon 1122 -3314 1122 -3314 0 3
rlabel polysilicon 1129 -3308 1129 -3308 0 1
rlabel polysilicon 1129 -3314 1129 -3314 0 3
rlabel polysilicon 1136 -3308 1136 -3308 0 1
rlabel polysilicon 1136 -3314 1136 -3314 0 3
rlabel polysilicon 1139 -3314 1139 -3314 0 4
rlabel polysilicon 1143 -3308 1143 -3308 0 1
rlabel polysilicon 1143 -3314 1143 -3314 0 3
rlabel polysilicon 1150 -3308 1150 -3308 0 1
rlabel polysilicon 1150 -3314 1150 -3314 0 3
rlabel polysilicon 1157 -3308 1157 -3308 0 1
rlabel polysilicon 1157 -3314 1157 -3314 0 3
rlabel polysilicon 1164 -3308 1164 -3308 0 1
rlabel polysilicon 1164 -3314 1164 -3314 0 3
rlabel polysilicon 1171 -3308 1171 -3308 0 1
rlabel polysilicon 1171 -3314 1171 -3314 0 3
rlabel polysilicon 1178 -3308 1178 -3308 0 1
rlabel polysilicon 1178 -3314 1178 -3314 0 3
rlabel polysilicon 1185 -3308 1185 -3308 0 1
rlabel polysilicon 1185 -3314 1185 -3314 0 3
rlabel polysilicon 1192 -3308 1192 -3308 0 1
rlabel polysilicon 1192 -3314 1192 -3314 0 3
rlabel polysilicon 1199 -3308 1199 -3308 0 1
rlabel polysilicon 1199 -3314 1199 -3314 0 3
rlabel polysilicon 1206 -3308 1206 -3308 0 1
rlabel polysilicon 1206 -3314 1206 -3314 0 3
rlabel polysilicon 1213 -3308 1213 -3308 0 1
rlabel polysilicon 1213 -3314 1213 -3314 0 3
rlabel polysilicon 1220 -3308 1220 -3308 0 1
rlabel polysilicon 1220 -3314 1220 -3314 0 3
rlabel polysilicon 1227 -3308 1227 -3308 0 1
rlabel polysilicon 1227 -3314 1227 -3314 0 3
rlabel polysilicon 1234 -3308 1234 -3308 0 1
rlabel polysilicon 1234 -3314 1234 -3314 0 3
rlabel polysilicon 1241 -3308 1241 -3308 0 1
rlabel polysilicon 1241 -3314 1241 -3314 0 3
rlabel polysilicon 1248 -3308 1248 -3308 0 1
rlabel polysilicon 1248 -3314 1248 -3314 0 3
rlabel polysilicon 1255 -3308 1255 -3308 0 1
rlabel polysilicon 1255 -3314 1255 -3314 0 3
rlabel polysilicon 1262 -3308 1262 -3308 0 1
rlabel polysilicon 1262 -3314 1262 -3314 0 3
rlabel polysilicon 1272 -3308 1272 -3308 0 2
rlabel polysilicon 1269 -3314 1269 -3314 0 3
rlabel polysilicon 1272 -3314 1272 -3314 0 4
rlabel polysilicon 1276 -3308 1276 -3308 0 1
rlabel polysilicon 1276 -3314 1276 -3314 0 3
rlabel polysilicon 1290 -3308 1290 -3308 0 1
rlabel polysilicon 1290 -3314 1290 -3314 0 3
rlabel polysilicon 1339 -3308 1339 -3308 0 1
rlabel polysilicon 1339 -3314 1339 -3314 0 3
rlabel polysilicon 1346 -3308 1346 -3308 0 1
rlabel polysilicon 1346 -3314 1346 -3314 0 3
rlabel polysilicon 1353 -3308 1353 -3308 0 1
rlabel polysilicon 1353 -3314 1353 -3314 0 3
rlabel polysilicon 198 -3381 198 -3381 0 1
rlabel polysilicon 198 -3387 198 -3387 0 3
rlabel polysilicon 205 -3381 205 -3381 0 1
rlabel polysilicon 205 -3387 205 -3387 0 3
rlabel polysilicon 212 -3381 212 -3381 0 1
rlabel polysilicon 212 -3387 212 -3387 0 3
rlabel polysilicon 219 -3381 219 -3381 0 1
rlabel polysilicon 219 -3387 219 -3387 0 3
rlabel polysilicon 226 -3381 226 -3381 0 1
rlabel polysilicon 226 -3387 226 -3387 0 3
rlabel polysilicon 233 -3381 233 -3381 0 1
rlabel polysilicon 233 -3387 233 -3387 0 3
rlabel polysilicon 240 -3381 240 -3381 0 1
rlabel polysilicon 240 -3387 240 -3387 0 3
rlabel polysilicon 247 -3381 247 -3381 0 1
rlabel polysilicon 247 -3387 247 -3387 0 3
rlabel polysilicon 254 -3381 254 -3381 0 1
rlabel polysilicon 254 -3387 254 -3387 0 3
rlabel polysilicon 261 -3387 261 -3387 0 3
rlabel polysilicon 271 -3381 271 -3381 0 2
rlabel polysilicon 268 -3387 268 -3387 0 3
rlabel polysilicon 271 -3387 271 -3387 0 4
rlabel polysilicon 275 -3381 275 -3381 0 1
rlabel polysilicon 278 -3387 278 -3387 0 4
rlabel polysilicon 282 -3381 282 -3381 0 1
rlabel polysilicon 282 -3387 282 -3387 0 3
rlabel polysilicon 289 -3381 289 -3381 0 1
rlabel polysilicon 289 -3387 289 -3387 0 3
rlabel polysilicon 296 -3381 296 -3381 0 1
rlabel polysilicon 296 -3387 296 -3387 0 3
rlabel polysilicon 303 -3381 303 -3381 0 1
rlabel polysilicon 303 -3387 303 -3387 0 3
rlabel polysilicon 310 -3381 310 -3381 0 1
rlabel polysilicon 310 -3387 310 -3387 0 3
rlabel polysilicon 317 -3381 317 -3381 0 1
rlabel polysilicon 317 -3387 317 -3387 0 3
rlabel polysilicon 324 -3381 324 -3381 0 1
rlabel polysilicon 324 -3387 324 -3387 0 3
rlabel polysilicon 331 -3381 331 -3381 0 1
rlabel polysilicon 331 -3387 331 -3387 0 3
rlabel polysilicon 338 -3381 338 -3381 0 1
rlabel polysilicon 338 -3387 338 -3387 0 3
rlabel polysilicon 345 -3381 345 -3381 0 1
rlabel polysilicon 345 -3387 345 -3387 0 3
rlabel polysilicon 352 -3381 352 -3381 0 1
rlabel polysilicon 352 -3387 352 -3387 0 3
rlabel polysilicon 359 -3381 359 -3381 0 1
rlabel polysilicon 359 -3387 359 -3387 0 3
rlabel polysilicon 366 -3381 366 -3381 0 1
rlabel polysilicon 366 -3387 366 -3387 0 3
rlabel polysilicon 373 -3381 373 -3381 0 1
rlabel polysilicon 373 -3387 373 -3387 0 3
rlabel polysilicon 380 -3381 380 -3381 0 1
rlabel polysilicon 380 -3387 380 -3387 0 3
rlabel polysilicon 387 -3381 387 -3381 0 1
rlabel polysilicon 387 -3387 387 -3387 0 3
rlabel polysilicon 394 -3381 394 -3381 0 1
rlabel polysilicon 394 -3387 394 -3387 0 3
rlabel polysilicon 401 -3381 401 -3381 0 1
rlabel polysilicon 404 -3381 404 -3381 0 2
rlabel polysilicon 404 -3387 404 -3387 0 4
rlabel polysilicon 408 -3381 408 -3381 0 1
rlabel polysilicon 411 -3381 411 -3381 0 2
rlabel polysilicon 408 -3387 408 -3387 0 3
rlabel polysilicon 411 -3387 411 -3387 0 4
rlabel polysilicon 415 -3381 415 -3381 0 1
rlabel polysilicon 415 -3387 415 -3387 0 3
rlabel polysilicon 422 -3381 422 -3381 0 1
rlabel polysilicon 425 -3381 425 -3381 0 2
rlabel polysilicon 422 -3387 422 -3387 0 3
rlabel polysilicon 429 -3381 429 -3381 0 1
rlabel polysilicon 429 -3387 429 -3387 0 3
rlabel polysilicon 436 -3381 436 -3381 0 1
rlabel polysilicon 436 -3387 436 -3387 0 3
rlabel polysilicon 443 -3381 443 -3381 0 1
rlabel polysilicon 443 -3387 443 -3387 0 3
rlabel polysilicon 450 -3381 450 -3381 0 1
rlabel polysilicon 450 -3387 450 -3387 0 3
rlabel polysilicon 457 -3381 457 -3381 0 1
rlabel polysilicon 457 -3387 457 -3387 0 3
rlabel polysilicon 464 -3381 464 -3381 0 1
rlabel polysilicon 464 -3387 464 -3387 0 3
rlabel polysilicon 471 -3381 471 -3381 0 1
rlabel polysilicon 471 -3387 471 -3387 0 3
rlabel polysilicon 474 -3387 474 -3387 0 4
rlabel polysilicon 478 -3381 478 -3381 0 1
rlabel polysilicon 478 -3387 478 -3387 0 3
rlabel polysilicon 485 -3381 485 -3381 0 1
rlabel polysilicon 485 -3387 485 -3387 0 3
rlabel polysilicon 492 -3381 492 -3381 0 1
rlabel polysilicon 492 -3387 492 -3387 0 3
rlabel polysilicon 499 -3381 499 -3381 0 1
rlabel polysilicon 499 -3387 499 -3387 0 3
rlabel polysilicon 506 -3381 506 -3381 0 1
rlabel polysilicon 506 -3387 506 -3387 0 3
rlabel polysilicon 513 -3381 513 -3381 0 1
rlabel polysilicon 513 -3387 513 -3387 0 3
rlabel polysilicon 520 -3381 520 -3381 0 1
rlabel polysilicon 520 -3387 520 -3387 0 3
rlabel polysilicon 527 -3381 527 -3381 0 1
rlabel polysilicon 534 -3381 534 -3381 0 1
rlabel polysilicon 534 -3387 534 -3387 0 3
rlabel polysilicon 541 -3381 541 -3381 0 1
rlabel polysilicon 544 -3381 544 -3381 0 2
rlabel polysilicon 541 -3387 541 -3387 0 3
rlabel polysilicon 548 -3381 548 -3381 0 1
rlabel polysilicon 548 -3387 548 -3387 0 3
rlabel polysilicon 555 -3381 555 -3381 0 1
rlabel polysilicon 558 -3381 558 -3381 0 2
rlabel polysilicon 558 -3387 558 -3387 0 4
rlabel polysilicon 562 -3381 562 -3381 0 1
rlabel polysilicon 562 -3387 562 -3387 0 3
rlabel polysilicon 569 -3381 569 -3381 0 1
rlabel polysilicon 572 -3381 572 -3381 0 2
rlabel polysilicon 569 -3387 569 -3387 0 3
rlabel polysilicon 572 -3387 572 -3387 0 4
rlabel polysilicon 576 -3381 576 -3381 0 1
rlabel polysilicon 579 -3381 579 -3381 0 2
rlabel polysilicon 576 -3387 576 -3387 0 3
rlabel polysilicon 579 -3387 579 -3387 0 4
rlabel polysilicon 583 -3381 583 -3381 0 1
rlabel polysilicon 583 -3387 583 -3387 0 3
rlabel polysilicon 590 -3381 590 -3381 0 1
rlabel polysilicon 590 -3387 590 -3387 0 3
rlabel polysilicon 597 -3381 597 -3381 0 1
rlabel polysilicon 597 -3387 597 -3387 0 3
rlabel polysilicon 604 -3381 604 -3381 0 1
rlabel polysilicon 604 -3387 604 -3387 0 3
rlabel polysilicon 611 -3381 611 -3381 0 1
rlabel polysilicon 611 -3387 611 -3387 0 3
rlabel polysilicon 618 -3381 618 -3381 0 1
rlabel polysilicon 618 -3387 618 -3387 0 3
rlabel polysilicon 625 -3381 625 -3381 0 1
rlabel polysilicon 625 -3387 625 -3387 0 3
rlabel polysilicon 632 -3381 632 -3381 0 1
rlabel polysilicon 632 -3387 632 -3387 0 3
rlabel polysilicon 639 -3381 639 -3381 0 1
rlabel polysilicon 639 -3387 639 -3387 0 3
rlabel polysilicon 646 -3381 646 -3381 0 1
rlabel polysilicon 646 -3387 646 -3387 0 3
rlabel polysilicon 653 -3381 653 -3381 0 1
rlabel polysilicon 656 -3381 656 -3381 0 2
rlabel polysilicon 656 -3387 656 -3387 0 4
rlabel polysilicon 660 -3381 660 -3381 0 1
rlabel polysilicon 660 -3387 660 -3387 0 3
rlabel polysilicon 667 -3381 667 -3381 0 1
rlabel polysilicon 667 -3387 667 -3387 0 3
rlabel polysilicon 674 -3381 674 -3381 0 1
rlabel polysilicon 674 -3387 674 -3387 0 3
rlabel polysilicon 681 -3381 681 -3381 0 1
rlabel polysilicon 681 -3387 681 -3387 0 3
rlabel polysilicon 688 -3381 688 -3381 0 1
rlabel polysilicon 688 -3387 688 -3387 0 3
rlabel polysilicon 695 -3381 695 -3381 0 1
rlabel polysilicon 695 -3387 695 -3387 0 3
rlabel polysilicon 702 -3381 702 -3381 0 1
rlabel polysilicon 702 -3387 702 -3387 0 3
rlabel polysilicon 709 -3381 709 -3381 0 1
rlabel polysilicon 709 -3387 709 -3387 0 3
rlabel polysilicon 716 -3381 716 -3381 0 1
rlabel polysilicon 716 -3387 716 -3387 0 3
rlabel polysilicon 723 -3381 723 -3381 0 1
rlabel polysilicon 723 -3387 723 -3387 0 3
rlabel polysilicon 730 -3381 730 -3381 0 1
rlabel polysilicon 730 -3387 730 -3387 0 3
rlabel polysilicon 737 -3381 737 -3381 0 1
rlabel polysilicon 737 -3387 737 -3387 0 3
rlabel polysilicon 744 -3381 744 -3381 0 1
rlabel polysilicon 744 -3387 744 -3387 0 3
rlabel polysilicon 751 -3381 751 -3381 0 1
rlabel polysilicon 751 -3387 751 -3387 0 3
rlabel polysilicon 761 -3381 761 -3381 0 2
rlabel polysilicon 758 -3387 758 -3387 0 3
rlabel polysilicon 765 -3381 765 -3381 0 1
rlabel polysilicon 765 -3387 765 -3387 0 3
rlabel polysilicon 772 -3381 772 -3381 0 1
rlabel polysilicon 772 -3387 772 -3387 0 3
rlabel polysilicon 779 -3381 779 -3381 0 1
rlabel polysilicon 779 -3387 779 -3387 0 3
rlabel polysilicon 786 -3381 786 -3381 0 1
rlabel polysilicon 786 -3387 786 -3387 0 3
rlabel polysilicon 793 -3381 793 -3381 0 1
rlabel polysilicon 793 -3387 793 -3387 0 3
rlabel polysilicon 796 -3387 796 -3387 0 4
rlabel polysilicon 800 -3381 800 -3381 0 1
rlabel polysilicon 800 -3387 800 -3387 0 3
rlabel polysilicon 807 -3381 807 -3381 0 1
rlabel polysilicon 807 -3387 807 -3387 0 3
rlabel polysilicon 814 -3381 814 -3381 0 1
rlabel polysilicon 814 -3387 814 -3387 0 3
rlabel polysilicon 821 -3381 821 -3381 0 1
rlabel polysilicon 821 -3387 821 -3387 0 3
rlabel polysilicon 828 -3381 828 -3381 0 1
rlabel polysilicon 828 -3387 828 -3387 0 3
rlabel polysilicon 835 -3381 835 -3381 0 1
rlabel polysilicon 835 -3387 835 -3387 0 3
rlabel polysilicon 842 -3381 842 -3381 0 1
rlabel polysilicon 842 -3387 842 -3387 0 3
rlabel polysilicon 849 -3381 849 -3381 0 1
rlabel polysilicon 849 -3387 849 -3387 0 3
rlabel polysilicon 856 -3381 856 -3381 0 1
rlabel polysilicon 856 -3387 856 -3387 0 3
rlabel polysilicon 863 -3381 863 -3381 0 1
rlabel polysilicon 863 -3387 863 -3387 0 3
rlabel polysilicon 870 -3381 870 -3381 0 1
rlabel polysilicon 870 -3387 870 -3387 0 3
rlabel polysilicon 877 -3381 877 -3381 0 1
rlabel polysilicon 877 -3387 877 -3387 0 3
rlabel polysilicon 884 -3381 884 -3381 0 1
rlabel polysilicon 884 -3387 884 -3387 0 3
rlabel polysilicon 891 -3381 891 -3381 0 1
rlabel polysilicon 891 -3387 891 -3387 0 3
rlabel polysilicon 898 -3381 898 -3381 0 1
rlabel polysilicon 898 -3387 898 -3387 0 3
rlabel polysilicon 905 -3381 905 -3381 0 1
rlabel polysilicon 905 -3387 905 -3387 0 3
rlabel polysilicon 912 -3381 912 -3381 0 1
rlabel polysilicon 912 -3387 912 -3387 0 3
rlabel polysilicon 919 -3381 919 -3381 0 1
rlabel polysilicon 919 -3387 919 -3387 0 3
rlabel polysilicon 926 -3381 926 -3381 0 1
rlabel polysilicon 926 -3387 926 -3387 0 3
rlabel polysilicon 933 -3381 933 -3381 0 1
rlabel polysilicon 933 -3387 933 -3387 0 3
rlabel polysilicon 940 -3381 940 -3381 0 1
rlabel polysilicon 940 -3387 940 -3387 0 3
rlabel polysilicon 947 -3381 947 -3381 0 1
rlabel polysilicon 947 -3387 947 -3387 0 3
rlabel polysilicon 954 -3381 954 -3381 0 1
rlabel polysilicon 957 -3387 957 -3387 0 4
rlabel polysilicon 961 -3381 961 -3381 0 1
rlabel polysilicon 961 -3387 961 -3387 0 3
rlabel polysilicon 968 -3381 968 -3381 0 1
rlabel polysilicon 968 -3387 968 -3387 0 3
rlabel polysilicon 975 -3381 975 -3381 0 1
rlabel polysilicon 975 -3387 975 -3387 0 3
rlabel polysilicon 982 -3381 982 -3381 0 1
rlabel polysilicon 982 -3387 982 -3387 0 3
rlabel polysilicon 989 -3381 989 -3381 0 1
rlabel polysilicon 989 -3387 989 -3387 0 3
rlabel polysilicon 996 -3381 996 -3381 0 1
rlabel polysilicon 996 -3387 996 -3387 0 3
rlabel polysilicon 1003 -3381 1003 -3381 0 1
rlabel polysilicon 1003 -3387 1003 -3387 0 3
rlabel polysilicon 1010 -3381 1010 -3381 0 1
rlabel polysilicon 1013 -3381 1013 -3381 0 2
rlabel polysilicon 1010 -3387 1010 -3387 0 3
rlabel polysilicon 1013 -3387 1013 -3387 0 4
rlabel polysilicon 1017 -3381 1017 -3381 0 1
rlabel polysilicon 1017 -3387 1017 -3387 0 3
rlabel polysilicon 1024 -3381 1024 -3381 0 1
rlabel polysilicon 1024 -3387 1024 -3387 0 3
rlabel polysilicon 1031 -3381 1031 -3381 0 1
rlabel polysilicon 1031 -3387 1031 -3387 0 3
rlabel polysilicon 1041 -3381 1041 -3381 0 2
rlabel polysilicon 1038 -3387 1038 -3387 0 3
rlabel polysilicon 1045 -3381 1045 -3381 0 1
rlabel polysilicon 1045 -3387 1045 -3387 0 3
rlabel polysilicon 1052 -3381 1052 -3381 0 1
rlabel polysilicon 1055 -3381 1055 -3381 0 2
rlabel polysilicon 1059 -3381 1059 -3381 0 1
rlabel polysilicon 1059 -3387 1059 -3387 0 3
rlabel polysilicon 1066 -3381 1066 -3381 0 1
rlabel polysilicon 1069 -3381 1069 -3381 0 2
rlabel polysilicon 1066 -3387 1066 -3387 0 3
rlabel polysilicon 1073 -3381 1073 -3381 0 1
rlabel polysilicon 1073 -3387 1073 -3387 0 3
rlabel polysilicon 1080 -3381 1080 -3381 0 1
rlabel polysilicon 1080 -3387 1080 -3387 0 3
rlabel polysilicon 1087 -3381 1087 -3381 0 1
rlabel polysilicon 1087 -3387 1087 -3387 0 3
rlabel polysilicon 1094 -3381 1094 -3381 0 1
rlabel polysilicon 1094 -3387 1094 -3387 0 3
rlabel polysilicon 1101 -3381 1101 -3381 0 1
rlabel polysilicon 1101 -3387 1101 -3387 0 3
rlabel polysilicon 1122 -3381 1122 -3381 0 1
rlabel polysilicon 1122 -3387 1122 -3387 0 3
rlabel polysilicon 1129 -3381 1129 -3381 0 1
rlabel polysilicon 1129 -3387 1129 -3387 0 3
rlabel polysilicon 1181 -3381 1181 -3381 0 2
rlabel polysilicon 1181 -3387 1181 -3387 0 4
rlabel polysilicon 1185 -3381 1185 -3381 0 1
rlabel polysilicon 1185 -3387 1185 -3387 0 3
rlabel polysilicon 1192 -3381 1192 -3381 0 1
rlabel polysilicon 1192 -3387 1192 -3387 0 3
rlabel polysilicon 1339 -3381 1339 -3381 0 1
rlabel polysilicon 1339 -3387 1339 -3387 0 3
rlabel polysilicon 1346 -3381 1346 -3381 0 1
rlabel polysilicon 1346 -3387 1346 -3387 0 3
rlabel polysilicon 1349 -3387 1349 -3387 0 4
rlabel polysilicon 1353 -3381 1353 -3381 0 1
rlabel polysilicon 1353 -3387 1353 -3387 0 3
rlabel polysilicon 247 -3444 247 -3444 0 1
rlabel polysilicon 247 -3450 247 -3450 0 3
rlabel polysilicon 261 -3444 261 -3444 0 1
rlabel polysilicon 261 -3450 261 -3450 0 3
rlabel polysilicon 292 -3444 292 -3444 0 2
rlabel polysilicon 289 -3450 289 -3450 0 3
rlabel polysilicon 292 -3450 292 -3450 0 4
rlabel polysilicon 310 -3444 310 -3444 0 1
rlabel polysilicon 310 -3450 310 -3450 0 3
rlabel polysilicon 317 -3444 317 -3444 0 1
rlabel polysilicon 317 -3450 317 -3450 0 3
rlabel polysilicon 324 -3444 324 -3444 0 1
rlabel polysilicon 324 -3450 324 -3450 0 3
rlabel polysilicon 331 -3444 331 -3444 0 1
rlabel polysilicon 331 -3450 331 -3450 0 3
rlabel polysilicon 338 -3444 338 -3444 0 1
rlabel polysilicon 338 -3450 338 -3450 0 3
rlabel polysilicon 345 -3444 345 -3444 0 1
rlabel polysilicon 348 -3444 348 -3444 0 2
rlabel polysilicon 352 -3444 352 -3444 0 1
rlabel polysilicon 352 -3450 352 -3450 0 3
rlabel polysilicon 359 -3444 359 -3444 0 1
rlabel polysilicon 359 -3450 359 -3450 0 3
rlabel polysilicon 366 -3444 366 -3444 0 1
rlabel polysilicon 373 -3444 373 -3444 0 1
rlabel polysilicon 373 -3450 373 -3450 0 3
rlabel polysilicon 380 -3444 380 -3444 0 1
rlabel polysilicon 380 -3450 380 -3450 0 3
rlabel polysilicon 387 -3444 387 -3444 0 1
rlabel polysilicon 394 -3444 394 -3444 0 1
rlabel polysilicon 394 -3450 394 -3450 0 3
rlabel polysilicon 401 -3444 401 -3444 0 1
rlabel polysilicon 408 -3444 408 -3444 0 1
rlabel polysilicon 408 -3450 408 -3450 0 3
rlabel polysilicon 415 -3444 415 -3444 0 1
rlabel polysilicon 415 -3450 415 -3450 0 3
rlabel polysilicon 422 -3444 422 -3444 0 1
rlabel polysilicon 422 -3450 422 -3450 0 3
rlabel polysilicon 429 -3444 429 -3444 0 1
rlabel polysilicon 429 -3450 429 -3450 0 3
rlabel polysilicon 436 -3444 436 -3444 0 1
rlabel polysilicon 436 -3450 436 -3450 0 3
rlabel polysilicon 446 -3444 446 -3444 0 2
rlabel polysilicon 443 -3450 443 -3450 0 3
rlabel polysilicon 446 -3450 446 -3450 0 4
rlabel polysilicon 450 -3444 450 -3444 0 1
rlabel polysilicon 450 -3450 450 -3450 0 3
rlabel polysilicon 457 -3444 457 -3444 0 1
rlabel polysilicon 457 -3450 457 -3450 0 3
rlabel polysilicon 464 -3444 464 -3444 0 1
rlabel polysilicon 464 -3450 464 -3450 0 3
rlabel polysilicon 471 -3444 471 -3444 0 1
rlabel polysilicon 471 -3450 471 -3450 0 3
rlabel polysilicon 478 -3444 478 -3444 0 1
rlabel polysilicon 478 -3450 478 -3450 0 3
rlabel polysilicon 485 -3444 485 -3444 0 1
rlabel polysilicon 485 -3450 485 -3450 0 3
rlabel polysilicon 492 -3444 492 -3444 0 1
rlabel polysilicon 492 -3450 492 -3450 0 3
rlabel polysilicon 499 -3444 499 -3444 0 1
rlabel polysilicon 502 -3444 502 -3444 0 2
rlabel polysilicon 499 -3450 499 -3450 0 3
rlabel polysilicon 506 -3444 506 -3444 0 1
rlabel polysilicon 506 -3450 506 -3450 0 3
rlabel polysilicon 513 -3444 513 -3444 0 1
rlabel polysilicon 513 -3450 513 -3450 0 3
rlabel polysilicon 520 -3444 520 -3444 0 1
rlabel polysilicon 520 -3450 520 -3450 0 3
rlabel polysilicon 530 -3444 530 -3444 0 2
rlabel polysilicon 527 -3450 527 -3450 0 3
rlabel polysilicon 530 -3450 530 -3450 0 4
rlabel polysilicon 534 -3444 534 -3444 0 1
rlabel polysilicon 534 -3450 534 -3450 0 3
rlabel polysilicon 541 -3444 541 -3444 0 1
rlabel polysilicon 541 -3450 541 -3450 0 3
rlabel polysilicon 548 -3444 548 -3444 0 1
rlabel polysilicon 548 -3450 548 -3450 0 3
rlabel polysilicon 555 -3444 555 -3444 0 1
rlabel polysilicon 555 -3450 555 -3450 0 3
rlabel polysilicon 562 -3444 562 -3444 0 1
rlabel polysilicon 562 -3450 562 -3450 0 3
rlabel polysilicon 569 -3444 569 -3444 0 1
rlabel polysilicon 569 -3450 569 -3450 0 3
rlabel polysilicon 576 -3444 576 -3444 0 1
rlabel polysilicon 576 -3450 576 -3450 0 3
rlabel polysilicon 583 -3444 583 -3444 0 1
rlabel polysilicon 583 -3450 583 -3450 0 3
rlabel polysilicon 590 -3444 590 -3444 0 1
rlabel polysilicon 590 -3450 590 -3450 0 3
rlabel polysilicon 597 -3444 597 -3444 0 1
rlabel polysilicon 597 -3450 597 -3450 0 3
rlabel polysilicon 604 -3444 604 -3444 0 1
rlabel polysilicon 604 -3450 604 -3450 0 3
rlabel polysilicon 611 -3444 611 -3444 0 1
rlabel polysilicon 611 -3450 611 -3450 0 3
rlabel polysilicon 618 -3444 618 -3444 0 1
rlabel polysilicon 618 -3450 618 -3450 0 3
rlabel polysilicon 625 -3444 625 -3444 0 1
rlabel polysilicon 625 -3450 625 -3450 0 3
rlabel polysilicon 632 -3444 632 -3444 0 1
rlabel polysilicon 632 -3450 632 -3450 0 3
rlabel polysilicon 639 -3444 639 -3444 0 1
rlabel polysilicon 639 -3450 639 -3450 0 3
rlabel polysilicon 646 -3444 646 -3444 0 1
rlabel polysilicon 649 -3444 649 -3444 0 2
rlabel polysilicon 649 -3450 649 -3450 0 4
rlabel polysilicon 653 -3444 653 -3444 0 1
rlabel polysilicon 653 -3450 653 -3450 0 3
rlabel polysilicon 660 -3444 660 -3444 0 1
rlabel polysilicon 660 -3450 660 -3450 0 3
rlabel polysilicon 667 -3444 667 -3444 0 1
rlabel polysilicon 667 -3450 667 -3450 0 3
rlabel polysilicon 674 -3444 674 -3444 0 1
rlabel polysilicon 674 -3450 674 -3450 0 3
rlabel polysilicon 681 -3444 681 -3444 0 1
rlabel polysilicon 681 -3450 681 -3450 0 3
rlabel polysilicon 691 -3444 691 -3444 0 2
rlabel polysilicon 688 -3450 688 -3450 0 3
rlabel polysilicon 691 -3450 691 -3450 0 4
rlabel polysilicon 695 -3444 695 -3444 0 1
rlabel polysilicon 695 -3450 695 -3450 0 3
rlabel polysilicon 702 -3444 702 -3444 0 1
rlabel polysilicon 702 -3450 702 -3450 0 3
rlabel polysilicon 709 -3444 709 -3444 0 1
rlabel polysilicon 709 -3450 709 -3450 0 3
rlabel polysilicon 716 -3444 716 -3444 0 1
rlabel polysilicon 716 -3450 716 -3450 0 3
rlabel polysilicon 723 -3444 723 -3444 0 1
rlabel polysilicon 723 -3450 723 -3450 0 3
rlabel polysilicon 730 -3444 730 -3444 0 1
rlabel polysilicon 730 -3450 730 -3450 0 3
rlabel polysilicon 737 -3444 737 -3444 0 1
rlabel polysilicon 740 -3444 740 -3444 0 2
rlabel polysilicon 737 -3450 737 -3450 0 3
rlabel polysilicon 740 -3450 740 -3450 0 4
rlabel polysilicon 744 -3444 744 -3444 0 1
rlabel polysilicon 744 -3450 744 -3450 0 3
rlabel polysilicon 751 -3444 751 -3444 0 1
rlabel polysilicon 751 -3450 751 -3450 0 3
rlabel polysilicon 758 -3444 758 -3444 0 1
rlabel polysilicon 765 -3444 765 -3444 0 1
rlabel polysilicon 765 -3450 765 -3450 0 3
rlabel polysilicon 772 -3444 772 -3444 0 1
rlabel polysilicon 772 -3450 772 -3450 0 3
rlabel polysilicon 779 -3444 779 -3444 0 1
rlabel polysilicon 779 -3450 779 -3450 0 3
rlabel polysilicon 786 -3444 786 -3444 0 1
rlabel polysilicon 786 -3450 786 -3450 0 3
rlabel polysilicon 793 -3444 793 -3444 0 1
rlabel polysilicon 793 -3450 793 -3450 0 3
rlabel polysilicon 800 -3444 800 -3444 0 1
rlabel polysilicon 800 -3450 800 -3450 0 3
rlabel polysilicon 807 -3444 807 -3444 0 1
rlabel polysilicon 807 -3450 807 -3450 0 3
rlabel polysilicon 814 -3444 814 -3444 0 1
rlabel polysilicon 814 -3450 814 -3450 0 3
rlabel polysilicon 824 -3444 824 -3444 0 2
rlabel polysilicon 821 -3450 821 -3450 0 3
rlabel polysilicon 824 -3450 824 -3450 0 4
rlabel polysilicon 828 -3444 828 -3444 0 1
rlabel polysilicon 828 -3450 828 -3450 0 3
rlabel polysilicon 835 -3444 835 -3444 0 1
rlabel polysilicon 835 -3450 835 -3450 0 3
rlabel polysilicon 842 -3444 842 -3444 0 1
rlabel polysilicon 842 -3450 842 -3450 0 3
rlabel polysilicon 849 -3444 849 -3444 0 1
rlabel polysilicon 849 -3450 849 -3450 0 3
rlabel polysilicon 859 -3444 859 -3444 0 2
rlabel polysilicon 856 -3450 856 -3450 0 3
rlabel polysilicon 859 -3450 859 -3450 0 4
rlabel polysilicon 863 -3444 863 -3444 0 1
rlabel polysilicon 863 -3450 863 -3450 0 3
rlabel polysilicon 873 -3444 873 -3444 0 2
rlabel polysilicon 870 -3450 870 -3450 0 3
rlabel polysilicon 877 -3444 877 -3444 0 1
rlabel polysilicon 877 -3450 877 -3450 0 3
rlabel polysilicon 884 -3444 884 -3444 0 1
rlabel polysilicon 887 -3444 887 -3444 0 2
rlabel polysilicon 884 -3450 884 -3450 0 3
rlabel polysilicon 887 -3450 887 -3450 0 4
rlabel polysilicon 891 -3444 891 -3444 0 1
rlabel polysilicon 891 -3450 891 -3450 0 3
rlabel polysilicon 898 -3450 898 -3450 0 3
rlabel polysilicon 901 -3450 901 -3450 0 4
rlabel polysilicon 905 -3444 905 -3444 0 1
rlabel polysilicon 905 -3450 905 -3450 0 3
rlabel polysilicon 912 -3444 912 -3444 0 1
rlabel polysilicon 912 -3450 912 -3450 0 3
rlabel polysilicon 919 -3444 919 -3444 0 1
rlabel polysilicon 919 -3450 919 -3450 0 3
rlabel polysilicon 926 -3444 926 -3444 0 1
rlabel polysilicon 926 -3450 926 -3450 0 3
rlabel polysilicon 933 -3444 933 -3444 0 1
rlabel polysilicon 933 -3450 933 -3450 0 3
rlabel polysilicon 936 -3450 936 -3450 0 4
rlabel polysilicon 940 -3444 940 -3444 0 1
rlabel polysilicon 940 -3450 940 -3450 0 3
rlabel polysilicon 943 -3450 943 -3450 0 4
rlabel polysilicon 947 -3444 947 -3444 0 1
rlabel polysilicon 947 -3450 947 -3450 0 3
rlabel polysilicon 954 -3444 954 -3444 0 1
rlabel polysilicon 954 -3450 954 -3450 0 3
rlabel polysilicon 961 -3444 961 -3444 0 1
rlabel polysilicon 961 -3450 961 -3450 0 3
rlabel polysilicon 968 -3444 968 -3444 0 1
rlabel polysilicon 968 -3450 968 -3450 0 3
rlabel polysilicon 975 -3444 975 -3444 0 1
rlabel polysilicon 975 -3450 975 -3450 0 3
rlabel polysilicon 982 -3444 982 -3444 0 1
rlabel polysilicon 982 -3450 982 -3450 0 3
rlabel polysilicon 1003 -3444 1003 -3444 0 1
rlabel polysilicon 1003 -3450 1003 -3450 0 3
rlabel polysilicon 1010 -3444 1010 -3444 0 1
rlabel polysilicon 1010 -3450 1010 -3450 0 3
rlabel polysilicon 1024 -3444 1024 -3444 0 1
rlabel polysilicon 1027 -3444 1027 -3444 0 2
rlabel polysilicon 1027 -3450 1027 -3450 0 4
rlabel polysilicon 1031 -3444 1031 -3444 0 1
rlabel polysilicon 1031 -3450 1031 -3450 0 3
rlabel polysilicon 1038 -3444 1038 -3444 0 1
rlabel polysilicon 1038 -3450 1038 -3450 0 3
rlabel polysilicon 1045 -3444 1045 -3444 0 1
rlabel polysilicon 1045 -3450 1045 -3450 0 3
rlabel polysilicon 1087 -3444 1087 -3444 0 1
rlabel polysilicon 1087 -3450 1087 -3450 0 3
rlabel polysilicon 1094 -3444 1094 -3444 0 1
rlabel polysilicon 1094 -3450 1094 -3450 0 3
rlabel polysilicon 1115 -3444 1115 -3444 0 1
rlabel polysilicon 1115 -3450 1115 -3450 0 3
rlabel polysilicon 1136 -3444 1136 -3444 0 1
rlabel polysilicon 1136 -3450 1136 -3450 0 3
rlabel polysilicon 1178 -3444 1178 -3444 0 1
rlabel polysilicon 1178 -3450 1178 -3450 0 3
rlabel polysilicon 1339 -3444 1339 -3444 0 1
rlabel polysilicon 1339 -3450 1339 -3450 0 3
rlabel polysilicon 1342 -3450 1342 -3450 0 4
rlabel polysilicon 1346 -3444 1346 -3444 0 1
rlabel polysilicon 1349 -3444 1349 -3444 0 2
rlabel polysilicon 1346 -3450 1346 -3450 0 3
rlabel polysilicon 1353 -3444 1353 -3444 0 1
rlabel polysilicon 1353 -3450 1353 -3450 0 3
rlabel polysilicon 247 -3501 247 -3501 0 1
rlabel polysilicon 247 -3507 247 -3507 0 3
rlabel polysilicon 261 -3501 261 -3501 0 1
rlabel polysilicon 261 -3507 261 -3507 0 3
rlabel polysilicon 275 -3501 275 -3501 0 1
rlabel polysilicon 275 -3507 275 -3507 0 3
rlabel polysilicon 331 -3501 331 -3501 0 1
rlabel polysilicon 331 -3507 331 -3507 0 3
rlabel polysilicon 338 -3501 338 -3501 0 1
rlabel polysilicon 338 -3507 338 -3507 0 3
rlabel polysilicon 345 -3501 345 -3501 0 1
rlabel polysilicon 345 -3507 345 -3507 0 3
rlabel polysilicon 352 -3501 352 -3501 0 1
rlabel polysilicon 352 -3507 352 -3507 0 3
rlabel polysilicon 359 -3501 359 -3501 0 1
rlabel polysilicon 359 -3507 359 -3507 0 3
rlabel polysilicon 366 -3501 366 -3501 0 1
rlabel polysilicon 366 -3507 366 -3507 0 3
rlabel polysilicon 373 -3501 373 -3501 0 1
rlabel polysilicon 373 -3507 373 -3507 0 3
rlabel polysilicon 380 -3501 380 -3501 0 1
rlabel polysilicon 380 -3507 380 -3507 0 3
rlabel polysilicon 387 -3507 387 -3507 0 3
rlabel polysilicon 394 -3501 394 -3501 0 1
rlabel polysilicon 394 -3507 394 -3507 0 3
rlabel polysilicon 401 -3507 401 -3507 0 3
rlabel polysilicon 408 -3501 408 -3501 0 1
rlabel polysilicon 408 -3507 408 -3507 0 3
rlabel polysilicon 415 -3501 415 -3501 0 1
rlabel polysilicon 415 -3507 415 -3507 0 3
rlabel polysilicon 422 -3501 422 -3501 0 1
rlabel polysilicon 425 -3501 425 -3501 0 2
rlabel polysilicon 422 -3507 422 -3507 0 3
rlabel polysilicon 425 -3507 425 -3507 0 4
rlabel polysilicon 429 -3501 429 -3501 0 1
rlabel polysilicon 429 -3507 429 -3507 0 3
rlabel polysilicon 436 -3501 436 -3501 0 1
rlabel polysilicon 436 -3507 436 -3507 0 3
rlabel polysilicon 443 -3501 443 -3501 0 1
rlabel polysilicon 443 -3507 443 -3507 0 3
rlabel polysilicon 450 -3501 450 -3501 0 1
rlabel polysilicon 450 -3507 450 -3507 0 3
rlabel polysilicon 457 -3501 457 -3501 0 1
rlabel polysilicon 457 -3507 457 -3507 0 3
rlabel polysilicon 464 -3501 464 -3501 0 1
rlabel polysilicon 467 -3501 467 -3501 0 2
rlabel polysilicon 464 -3507 464 -3507 0 3
rlabel polysilicon 467 -3507 467 -3507 0 4
rlabel polysilicon 471 -3501 471 -3501 0 1
rlabel polysilicon 471 -3507 471 -3507 0 3
rlabel polysilicon 478 -3501 478 -3501 0 1
rlabel polysilicon 478 -3507 478 -3507 0 3
rlabel polysilicon 485 -3501 485 -3501 0 1
rlabel polysilicon 485 -3507 485 -3507 0 3
rlabel polysilicon 492 -3501 492 -3501 0 1
rlabel polysilicon 492 -3507 492 -3507 0 3
rlabel polysilicon 495 -3507 495 -3507 0 4
rlabel polysilicon 499 -3501 499 -3501 0 1
rlabel polysilicon 499 -3507 499 -3507 0 3
rlabel polysilicon 506 -3501 506 -3501 0 1
rlabel polysilicon 506 -3507 506 -3507 0 3
rlabel polysilicon 513 -3501 513 -3501 0 1
rlabel polysilicon 513 -3507 513 -3507 0 3
rlabel polysilicon 520 -3501 520 -3501 0 1
rlabel polysilicon 520 -3507 520 -3507 0 3
rlabel polysilicon 527 -3501 527 -3501 0 1
rlabel polysilicon 527 -3507 527 -3507 0 3
rlabel polysilicon 534 -3501 534 -3501 0 1
rlabel polysilicon 537 -3501 537 -3501 0 2
rlabel polysilicon 534 -3507 534 -3507 0 3
rlabel polysilicon 541 -3501 541 -3501 0 1
rlabel polysilicon 541 -3507 541 -3507 0 3
rlabel polysilicon 548 -3501 548 -3501 0 1
rlabel polysilicon 548 -3507 548 -3507 0 3
rlabel polysilicon 555 -3501 555 -3501 0 1
rlabel polysilicon 555 -3507 555 -3507 0 3
rlabel polysilicon 562 -3501 562 -3501 0 1
rlabel polysilicon 562 -3507 562 -3507 0 3
rlabel polysilicon 565 -3507 565 -3507 0 4
rlabel polysilicon 569 -3501 569 -3501 0 1
rlabel polysilicon 569 -3507 569 -3507 0 3
rlabel polysilicon 579 -3501 579 -3501 0 2
rlabel polysilicon 576 -3507 576 -3507 0 3
rlabel polysilicon 579 -3507 579 -3507 0 4
rlabel polysilicon 583 -3501 583 -3501 0 1
rlabel polysilicon 583 -3507 583 -3507 0 3
rlabel polysilicon 590 -3501 590 -3501 0 1
rlabel polysilicon 590 -3507 590 -3507 0 3
rlabel polysilicon 597 -3501 597 -3501 0 1
rlabel polysilicon 597 -3507 597 -3507 0 3
rlabel polysilicon 604 -3501 604 -3501 0 1
rlabel polysilicon 604 -3507 604 -3507 0 3
rlabel polysilicon 611 -3501 611 -3501 0 1
rlabel polysilicon 611 -3507 611 -3507 0 3
rlabel polysilicon 618 -3501 618 -3501 0 1
rlabel polysilicon 618 -3507 618 -3507 0 3
rlabel polysilicon 625 -3501 625 -3501 0 1
rlabel polysilicon 628 -3501 628 -3501 0 2
rlabel polysilicon 625 -3507 625 -3507 0 3
rlabel polysilicon 632 -3501 632 -3501 0 1
rlabel polysilicon 632 -3507 632 -3507 0 3
rlabel polysilicon 639 -3501 639 -3501 0 1
rlabel polysilicon 639 -3507 639 -3507 0 3
rlabel polysilicon 642 -3507 642 -3507 0 4
rlabel polysilicon 646 -3501 646 -3501 0 1
rlabel polysilicon 646 -3507 646 -3507 0 3
rlabel polysilicon 653 -3501 653 -3501 0 1
rlabel polysilicon 653 -3507 653 -3507 0 3
rlabel polysilicon 660 -3501 660 -3501 0 1
rlabel polysilicon 660 -3507 660 -3507 0 3
rlabel polysilicon 667 -3501 667 -3501 0 1
rlabel polysilicon 667 -3507 667 -3507 0 3
rlabel polysilicon 677 -3501 677 -3501 0 2
rlabel polysilicon 674 -3507 674 -3507 0 3
rlabel polysilicon 677 -3507 677 -3507 0 4
rlabel polysilicon 681 -3501 681 -3501 0 1
rlabel polysilicon 681 -3507 681 -3507 0 3
rlabel polysilicon 688 -3501 688 -3501 0 1
rlabel polysilicon 688 -3507 688 -3507 0 3
rlabel polysilicon 695 -3501 695 -3501 0 1
rlabel polysilicon 695 -3507 695 -3507 0 3
rlabel polysilicon 702 -3501 702 -3501 0 1
rlabel polysilicon 702 -3507 702 -3507 0 3
rlabel polysilicon 709 -3501 709 -3501 0 1
rlabel polysilicon 709 -3507 709 -3507 0 3
rlabel polysilicon 716 -3501 716 -3501 0 1
rlabel polysilicon 716 -3507 716 -3507 0 3
rlabel polysilicon 726 -3501 726 -3501 0 2
rlabel polysilicon 726 -3507 726 -3507 0 4
rlabel polysilicon 730 -3501 730 -3501 0 1
rlabel polysilicon 730 -3507 730 -3507 0 3
rlabel polysilicon 737 -3501 737 -3501 0 1
rlabel polysilicon 737 -3507 737 -3507 0 3
rlabel polysilicon 744 -3501 744 -3501 0 1
rlabel polysilicon 744 -3507 744 -3507 0 3
rlabel polysilicon 751 -3501 751 -3501 0 1
rlabel polysilicon 751 -3507 751 -3507 0 3
rlabel polysilicon 758 -3507 758 -3507 0 3
rlabel polysilicon 765 -3501 765 -3501 0 1
rlabel polysilicon 765 -3507 765 -3507 0 3
rlabel polysilicon 772 -3501 772 -3501 0 1
rlabel polysilicon 772 -3507 772 -3507 0 3
rlabel polysilicon 779 -3501 779 -3501 0 1
rlabel polysilicon 779 -3507 779 -3507 0 3
rlabel polysilicon 800 -3501 800 -3501 0 1
rlabel polysilicon 800 -3507 800 -3507 0 3
rlabel polysilicon 807 -3501 807 -3501 0 1
rlabel polysilicon 807 -3507 807 -3507 0 3
rlabel polysilicon 814 -3501 814 -3501 0 1
rlabel polysilicon 817 -3501 817 -3501 0 2
rlabel polysilicon 821 -3501 821 -3501 0 1
rlabel polysilicon 821 -3507 821 -3507 0 3
rlabel polysilicon 835 -3501 835 -3501 0 1
rlabel polysilicon 835 -3507 835 -3507 0 3
rlabel polysilicon 842 -3501 842 -3501 0 1
rlabel polysilicon 842 -3507 842 -3507 0 3
rlabel polysilicon 849 -3501 849 -3501 0 1
rlabel polysilicon 849 -3507 849 -3507 0 3
rlabel polysilicon 856 -3501 856 -3501 0 1
rlabel polysilicon 856 -3507 856 -3507 0 3
rlabel polysilicon 863 -3501 863 -3501 0 1
rlabel polysilicon 863 -3507 863 -3507 0 3
rlabel polysilicon 870 -3501 870 -3501 0 1
rlabel polysilicon 870 -3507 870 -3507 0 3
rlabel polysilicon 877 -3501 877 -3501 0 1
rlabel polysilicon 877 -3507 877 -3507 0 3
rlabel polysilicon 905 -3501 905 -3501 0 1
rlabel polysilicon 905 -3507 905 -3507 0 3
rlabel polysilicon 912 -3501 912 -3501 0 1
rlabel polysilicon 912 -3507 912 -3507 0 3
rlabel polysilicon 919 -3501 919 -3501 0 1
rlabel polysilicon 919 -3507 919 -3507 0 3
rlabel polysilicon 926 -3501 926 -3501 0 1
rlabel polysilicon 926 -3507 926 -3507 0 3
rlabel polysilicon 933 -3501 933 -3501 0 1
rlabel polysilicon 936 -3501 936 -3501 0 2
rlabel polysilicon 933 -3507 933 -3507 0 3
rlabel polysilicon 940 -3501 940 -3501 0 1
rlabel polysilicon 943 -3501 943 -3501 0 2
rlabel polysilicon 940 -3507 940 -3507 0 3
rlabel polysilicon 947 -3501 947 -3501 0 1
rlabel polysilicon 947 -3507 947 -3507 0 3
rlabel polysilicon 954 -3501 954 -3501 0 1
rlabel polysilicon 957 -3501 957 -3501 0 2
rlabel polysilicon 954 -3507 954 -3507 0 3
rlabel polysilicon 961 -3501 961 -3501 0 1
rlabel polysilicon 961 -3507 961 -3507 0 3
rlabel polysilicon 968 -3501 968 -3501 0 1
rlabel polysilicon 968 -3507 968 -3507 0 3
rlabel polysilicon 982 -3501 982 -3501 0 1
rlabel polysilicon 982 -3507 982 -3507 0 3
rlabel polysilicon 989 -3501 989 -3501 0 1
rlabel polysilicon 989 -3507 989 -3507 0 3
rlabel polysilicon 996 -3501 996 -3501 0 1
rlabel polysilicon 999 -3501 999 -3501 0 2
rlabel polysilicon 996 -3507 996 -3507 0 3
rlabel polysilicon 1003 -3501 1003 -3501 0 1
rlabel polysilicon 1003 -3507 1003 -3507 0 3
rlabel polysilicon 1010 -3501 1010 -3501 0 1
rlabel polysilicon 1010 -3507 1010 -3507 0 3
rlabel polysilicon 1052 -3501 1052 -3501 0 1
rlabel polysilicon 1052 -3507 1052 -3507 0 3
rlabel polysilicon 1080 -3501 1080 -3501 0 1
rlabel polysilicon 1080 -3507 1080 -3507 0 3
rlabel polysilicon 1087 -3501 1087 -3501 0 1
rlabel polysilicon 1087 -3507 1087 -3507 0 3
rlabel polysilicon 1108 -3501 1108 -3501 0 1
rlabel polysilicon 1108 -3507 1108 -3507 0 3
rlabel polysilicon 1122 -3501 1122 -3501 0 1
rlabel polysilicon 1122 -3507 1122 -3507 0 3
rlabel polysilicon 1150 -3501 1150 -3501 0 1
rlabel polysilicon 1150 -3507 1150 -3507 0 3
rlabel polysilicon 1171 -3501 1171 -3501 0 1
rlabel polysilicon 1174 -3501 1174 -3501 0 2
rlabel polysilicon 1171 -3507 1171 -3507 0 3
rlabel polysilicon 1178 -3501 1178 -3501 0 1
rlabel polysilicon 1178 -3507 1178 -3507 0 3
rlabel polysilicon 1339 -3501 1339 -3501 0 1
rlabel polysilicon 1342 -3501 1342 -3501 0 2
rlabel polysilicon 1339 -3507 1339 -3507 0 3
rlabel polysilicon 1346 -3501 1346 -3501 0 1
rlabel polysilicon 1346 -3507 1346 -3507 0 3
rlabel polysilicon 1349 -3507 1349 -3507 0 4
rlabel polysilicon 1353 -3501 1353 -3501 0 1
rlabel polysilicon 1353 -3507 1353 -3507 0 3
rlabel polysilicon 247 -3542 247 -3542 0 1
rlabel polysilicon 247 -3548 247 -3548 0 3
rlabel polysilicon 254 -3542 254 -3542 0 1
rlabel polysilicon 257 -3548 257 -3548 0 4
rlabel polysilicon 261 -3542 261 -3542 0 1
rlabel polysilicon 261 -3548 261 -3548 0 3
rlabel polysilicon 268 -3542 268 -3542 0 1
rlabel polysilicon 268 -3548 268 -3548 0 3
rlabel polysilicon 296 -3542 296 -3542 0 1
rlabel polysilicon 296 -3548 296 -3548 0 3
rlabel polysilicon 345 -3542 345 -3542 0 1
rlabel polysilicon 345 -3548 345 -3548 0 3
rlabel polysilicon 359 -3542 359 -3542 0 1
rlabel polysilicon 359 -3548 359 -3548 0 3
rlabel polysilicon 380 -3542 380 -3542 0 1
rlabel polysilicon 380 -3548 380 -3548 0 3
rlabel polysilicon 394 -3542 394 -3542 0 1
rlabel polysilicon 394 -3548 394 -3548 0 3
rlabel polysilicon 401 -3542 401 -3542 0 1
rlabel polysilicon 401 -3548 401 -3548 0 3
rlabel polysilicon 408 -3542 408 -3542 0 1
rlabel polysilicon 408 -3548 408 -3548 0 3
rlabel polysilicon 415 -3542 415 -3542 0 1
rlabel polysilicon 415 -3548 415 -3548 0 3
rlabel polysilicon 422 -3542 422 -3542 0 1
rlabel polysilicon 422 -3548 422 -3548 0 3
rlabel polysilicon 429 -3542 429 -3542 0 1
rlabel polysilicon 432 -3548 432 -3548 0 4
rlabel polysilicon 436 -3542 436 -3542 0 1
rlabel polysilicon 436 -3548 436 -3548 0 3
rlabel polysilicon 443 -3542 443 -3542 0 1
rlabel polysilicon 450 -3542 450 -3542 0 1
rlabel polysilicon 453 -3542 453 -3542 0 2
rlabel polysilicon 450 -3548 450 -3548 0 3
rlabel polysilicon 453 -3548 453 -3548 0 4
rlabel polysilicon 457 -3542 457 -3542 0 1
rlabel polysilicon 457 -3548 457 -3548 0 3
rlabel polysilicon 464 -3542 464 -3542 0 1
rlabel polysilicon 464 -3548 464 -3548 0 3
rlabel polysilicon 471 -3542 471 -3542 0 1
rlabel polysilicon 471 -3548 471 -3548 0 3
rlabel polysilicon 478 -3542 478 -3542 0 1
rlabel polysilicon 478 -3548 478 -3548 0 3
rlabel polysilicon 488 -3548 488 -3548 0 4
rlabel polysilicon 492 -3542 492 -3542 0 1
rlabel polysilicon 492 -3548 492 -3548 0 3
rlabel polysilicon 499 -3542 499 -3542 0 1
rlabel polysilicon 499 -3548 499 -3548 0 3
rlabel polysilicon 506 -3542 506 -3542 0 1
rlabel polysilicon 506 -3548 506 -3548 0 3
rlabel polysilicon 513 -3542 513 -3542 0 1
rlabel polysilicon 513 -3548 513 -3548 0 3
rlabel polysilicon 520 -3542 520 -3542 0 1
rlabel polysilicon 520 -3548 520 -3548 0 3
rlabel polysilicon 527 -3542 527 -3542 0 1
rlabel polysilicon 527 -3548 527 -3548 0 3
rlabel polysilicon 534 -3542 534 -3542 0 1
rlabel polysilicon 534 -3548 534 -3548 0 3
rlabel polysilicon 541 -3542 541 -3542 0 1
rlabel polysilicon 544 -3542 544 -3542 0 2
rlabel polysilicon 541 -3548 541 -3548 0 3
rlabel polysilicon 544 -3548 544 -3548 0 4
rlabel polysilicon 548 -3542 548 -3542 0 1
rlabel polysilicon 548 -3548 548 -3548 0 3
rlabel polysilicon 555 -3542 555 -3542 0 1
rlabel polysilicon 555 -3548 555 -3548 0 3
rlabel polysilicon 562 -3542 562 -3542 0 1
rlabel polysilicon 562 -3548 562 -3548 0 3
rlabel polysilicon 569 -3542 569 -3542 0 1
rlabel polysilicon 569 -3548 569 -3548 0 3
rlabel polysilicon 576 -3542 576 -3542 0 1
rlabel polysilicon 576 -3548 576 -3548 0 3
rlabel polysilicon 583 -3542 583 -3542 0 1
rlabel polysilicon 583 -3548 583 -3548 0 3
rlabel polysilicon 590 -3542 590 -3542 0 1
rlabel polysilicon 590 -3548 590 -3548 0 3
rlabel polysilicon 600 -3542 600 -3542 0 2
rlabel polysilicon 600 -3548 600 -3548 0 4
rlabel polysilicon 604 -3542 604 -3542 0 1
rlabel polysilicon 604 -3548 604 -3548 0 3
rlabel polysilicon 611 -3542 611 -3542 0 1
rlabel polysilicon 611 -3548 611 -3548 0 3
rlabel polysilicon 625 -3542 625 -3542 0 1
rlabel polysilicon 628 -3542 628 -3542 0 2
rlabel polysilicon 628 -3548 628 -3548 0 4
rlabel polysilicon 639 -3542 639 -3542 0 1
rlabel polysilicon 639 -3548 639 -3548 0 3
rlabel polysilicon 667 -3542 667 -3542 0 1
rlabel polysilicon 667 -3548 667 -3548 0 3
rlabel polysilicon 681 -3542 681 -3542 0 1
rlabel polysilicon 681 -3548 681 -3548 0 3
rlabel polysilicon 688 -3542 688 -3542 0 1
rlabel polysilicon 691 -3542 691 -3542 0 2
rlabel polysilicon 695 -3542 695 -3542 0 1
rlabel polysilicon 695 -3548 695 -3548 0 3
rlabel polysilicon 702 -3542 702 -3542 0 1
rlabel polysilicon 702 -3548 702 -3548 0 3
rlabel polysilicon 709 -3542 709 -3542 0 1
rlabel polysilicon 716 -3542 716 -3542 0 1
rlabel polysilicon 716 -3548 716 -3548 0 3
rlabel polysilicon 723 -3542 723 -3542 0 1
rlabel polysilicon 723 -3548 723 -3548 0 3
rlabel polysilicon 726 -3548 726 -3548 0 4
rlabel polysilicon 730 -3542 730 -3542 0 1
rlabel polysilicon 730 -3548 730 -3548 0 3
rlabel polysilicon 737 -3542 737 -3542 0 1
rlabel polysilicon 737 -3548 737 -3548 0 3
rlabel polysilicon 744 -3542 744 -3542 0 1
rlabel polysilicon 744 -3548 744 -3548 0 3
rlabel polysilicon 751 -3542 751 -3542 0 1
rlabel polysilicon 751 -3548 751 -3548 0 3
rlabel polysilicon 758 -3542 758 -3542 0 1
rlabel polysilicon 758 -3548 758 -3548 0 3
rlabel polysilicon 765 -3542 765 -3542 0 1
rlabel polysilicon 765 -3548 765 -3548 0 3
rlabel polysilicon 835 -3542 835 -3542 0 1
rlabel polysilicon 835 -3548 835 -3548 0 3
rlabel polysilicon 849 -3542 849 -3542 0 1
rlabel polysilicon 849 -3548 849 -3548 0 3
rlabel polysilicon 863 -3542 863 -3542 0 1
rlabel polysilicon 863 -3548 863 -3548 0 3
rlabel polysilicon 870 -3542 870 -3542 0 1
rlabel polysilicon 870 -3548 870 -3548 0 3
rlabel polysilicon 877 -3542 877 -3542 0 1
rlabel polysilicon 877 -3548 877 -3548 0 3
rlabel polysilicon 884 -3542 884 -3542 0 1
rlabel polysilicon 884 -3548 884 -3548 0 3
rlabel polysilicon 891 -3542 891 -3542 0 1
rlabel polysilicon 891 -3548 891 -3548 0 3
rlabel polysilicon 898 -3542 898 -3542 0 1
rlabel polysilicon 898 -3548 898 -3548 0 3
rlabel polysilicon 905 -3542 905 -3542 0 1
rlabel polysilicon 905 -3548 905 -3548 0 3
rlabel polysilicon 912 -3542 912 -3542 0 1
rlabel polysilicon 912 -3548 912 -3548 0 3
rlabel polysilicon 922 -3542 922 -3542 0 2
rlabel polysilicon 919 -3548 919 -3548 0 3
rlabel polysilicon 926 -3542 926 -3542 0 1
rlabel polysilicon 926 -3548 926 -3548 0 3
rlabel polysilicon 933 -3542 933 -3542 0 1
rlabel polysilicon 933 -3548 933 -3548 0 3
rlabel polysilicon 940 -3542 940 -3542 0 1
rlabel polysilicon 943 -3542 943 -3542 0 2
rlabel polysilicon 947 -3542 947 -3542 0 1
rlabel polysilicon 947 -3548 947 -3548 0 3
rlabel polysilicon 968 -3542 968 -3542 0 1
rlabel polysilicon 968 -3548 968 -3548 0 3
rlabel polysilicon 975 -3542 975 -3542 0 1
rlabel polysilicon 975 -3548 975 -3548 0 3
rlabel polysilicon 989 -3542 989 -3542 0 1
rlabel polysilicon 989 -3548 989 -3548 0 3
rlabel polysilicon 1006 -3542 1006 -3542 0 2
rlabel polysilicon 1006 -3548 1006 -3548 0 4
rlabel polysilicon 1010 -3542 1010 -3542 0 1
rlabel polysilicon 1010 -3548 1010 -3548 0 3
rlabel polysilicon 1052 -3542 1052 -3542 0 1
rlabel polysilicon 1052 -3548 1052 -3548 0 3
rlabel polysilicon 1059 -3542 1059 -3542 0 1
rlabel polysilicon 1059 -3548 1059 -3548 0 3
rlabel polysilicon 1080 -3542 1080 -3542 0 1
rlabel polysilicon 1080 -3548 1080 -3548 0 3
rlabel polysilicon 1108 -3542 1108 -3542 0 1
rlabel polysilicon 1108 -3548 1108 -3548 0 3
rlabel polysilicon 1150 -3542 1150 -3542 0 1
rlabel polysilicon 1150 -3548 1150 -3548 0 3
rlabel polysilicon 1160 -3542 1160 -3542 0 2
rlabel polysilicon 1157 -3548 1157 -3548 0 3
rlabel polysilicon 261 -3579 261 -3579 0 1
rlabel polysilicon 264 -3585 264 -3585 0 4
rlabel polysilicon 268 -3579 268 -3579 0 1
rlabel polysilicon 268 -3585 268 -3585 0 3
rlabel polysilicon 310 -3579 310 -3579 0 1
rlabel polysilicon 310 -3585 310 -3585 0 3
rlabel polysilicon 327 -3579 327 -3579 0 2
rlabel polysilicon 324 -3585 324 -3585 0 3
rlabel polysilicon 327 -3585 327 -3585 0 4
rlabel polysilicon 352 -3579 352 -3579 0 1
rlabel polysilicon 352 -3585 352 -3585 0 3
rlabel polysilicon 359 -3579 359 -3579 0 1
rlabel polysilicon 359 -3585 359 -3585 0 3
rlabel polysilicon 366 -3579 366 -3579 0 1
rlabel polysilicon 366 -3585 366 -3585 0 3
rlabel polysilicon 376 -3579 376 -3579 0 2
rlabel polysilicon 376 -3585 376 -3585 0 4
rlabel polysilicon 394 -3579 394 -3579 0 1
rlabel polysilicon 394 -3585 394 -3585 0 3
rlabel polysilicon 401 -3579 401 -3579 0 1
rlabel polysilicon 404 -3585 404 -3585 0 4
rlabel polysilicon 408 -3579 408 -3579 0 1
rlabel polysilicon 408 -3585 408 -3585 0 3
rlabel polysilicon 415 -3579 415 -3579 0 1
rlabel polysilicon 415 -3585 415 -3585 0 3
rlabel polysilicon 436 -3579 436 -3579 0 1
rlabel polysilicon 436 -3585 436 -3585 0 3
rlabel polysilicon 443 -3579 443 -3579 0 1
rlabel polysilicon 443 -3585 443 -3585 0 3
rlabel polysilicon 446 -3585 446 -3585 0 4
rlabel polysilicon 450 -3579 450 -3579 0 1
rlabel polysilicon 450 -3585 450 -3585 0 3
rlabel polysilicon 457 -3579 457 -3579 0 1
rlabel polysilicon 457 -3585 457 -3585 0 3
rlabel polysilicon 464 -3579 464 -3579 0 1
rlabel polysilicon 464 -3585 464 -3585 0 3
rlabel polysilicon 471 -3579 471 -3579 0 1
rlabel polysilicon 471 -3585 471 -3585 0 3
rlabel polysilicon 478 -3579 478 -3579 0 1
rlabel polysilicon 478 -3585 478 -3585 0 3
rlabel polysilicon 485 -3579 485 -3579 0 1
rlabel polysilicon 488 -3579 488 -3579 0 2
rlabel polysilicon 492 -3579 492 -3579 0 1
rlabel polysilicon 492 -3585 492 -3585 0 3
rlabel polysilicon 499 -3579 499 -3579 0 1
rlabel polysilicon 499 -3585 499 -3585 0 3
rlabel polysilicon 506 -3579 506 -3579 0 1
rlabel polysilicon 506 -3585 506 -3585 0 3
rlabel polysilicon 513 -3579 513 -3579 0 1
rlabel polysilicon 516 -3585 516 -3585 0 4
rlabel polysilicon 520 -3579 520 -3579 0 1
rlabel polysilicon 520 -3585 520 -3585 0 3
rlabel polysilicon 527 -3579 527 -3579 0 1
rlabel polysilicon 527 -3585 527 -3585 0 3
rlabel polysilicon 534 -3579 534 -3579 0 1
rlabel polysilicon 534 -3585 534 -3585 0 3
rlabel polysilicon 541 -3579 541 -3579 0 1
rlabel polysilicon 541 -3585 541 -3585 0 3
rlabel polysilicon 548 -3579 548 -3579 0 1
rlabel polysilicon 548 -3585 548 -3585 0 3
rlabel polysilicon 555 -3579 555 -3579 0 1
rlabel polysilicon 555 -3585 555 -3585 0 3
rlabel polysilicon 562 -3579 562 -3579 0 1
rlabel polysilicon 562 -3585 562 -3585 0 3
rlabel polysilicon 569 -3579 569 -3579 0 1
rlabel polysilicon 569 -3585 569 -3585 0 3
rlabel polysilicon 597 -3579 597 -3579 0 1
rlabel polysilicon 597 -3585 597 -3585 0 3
rlabel polysilicon 611 -3579 611 -3579 0 1
rlabel polysilicon 611 -3585 611 -3585 0 3
rlabel polysilicon 618 -3579 618 -3579 0 1
rlabel polysilicon 618 -3585 618 -3585 0 3
rlabel polysilicon 646 -3579 646 -3579 0 1
rlabel polysilicon 646 -3585 646 -3585 0 3
rlabel polysilicon 660 -3579 660 -3579 0 1
rlabel polysilicon 660 -3585 660 -3585 0 3
rlabel polysilicon 677 -3579 677 -3579 0 2
rlabel polysilicon 674 -3585 674 -3585 0 3
rlabel polysilicon 677 -3585 677 -3585 0 4
rlabel polysilicon 688 -3579 688 -3579 0 1
rlabel polysilicon 688 -3585 688 -3585 0 3
rlabel polysilicon 695 -3579 695 -3579 0 1
rlabel polysilicon 695 -3585 695 -3585 0 3
rlabel polysilicon 702 -3579 702 -3579 0 1
rlabel polysilicon 702 -3585 702 -3585 0 3
rlabel polysilicon 709 -3585 709 -3585 0 3
rlabel polysilicon 716 -3579 716 -3579 0 1
rlabel polysilicon 716 -3585 716 -3585 0 3
rlabel polysilicon 723 -3579 723 -3579 0 1
rlabel polysilicon 726 -3579 726 -3579 0 2
rlabel polysilicon 723 -3585 723 -3585 0 3
rlabel polysilicon 730 -3579 730 -3579 0 1
rlabel polysilicon 730 -3585 730 -3585 0 3
rlabel polysilicon 737 -3579 737 -3579 0 1
rlabel polysilicon 737 -3585 737 -3585 0 3
rlabel polysilicon 744 -3579 744 -3579 0 1
rlabel polysilicon 744 -3585 744 -3585 0 3
rlabel polysilicon 751 -3579 751 -3579 0 1
rlabel polysilicon 751 -3585 751 -3585 0 3
rlabel polysilicon 758 -3579 758 -3579 0 1
rlabel polysilicon 758 -3585 758 -3585 0 3
rlabel polysilicon 765 -3579 765 -3579 0 1
rlabel polysilicon 765 -3585 765 -3585 0 3
rlabel polysilicon 849 -3579 849 -3579 0 1
rlabel polysilicon 849 -3585 849 -3585 0 3
rlabel polysilicon 856 -3579 856 -3579 0 1
rlabel polysilicon 856 -3585 856 -3585 0 3
rlabel polysilicon 891 -3579 891 -3579 0 1
rlabel polysilicon 891 -3585 891 -3585 0 3
rlabel polysilicon 901 -3579 901 -3579 0 2
rlabel polysilicon 901 -3585 901 -3585 0 4
rlabel polysilicon 905 -3579 905 -3579 0 1
rlabel polysilicon 905 -3585 905 -3585 0 3
rlabel polysilicon 912 -3579 912 -3579 0 1
rlabel polysilicon 912 -3585 912 -3585 0 3
rlabel polysilicon 919 -3579 919 -3579 0 1
rlabel polysilicon 922 -3579 922 -3579 0 2
rlabel polysilicon 926 -3579 926 -3579 0 1
rlabel polysilicon 926 -3585 926 -3585 0 3
rlabel polysilicon 940 -3579 940 -3579 0 1
rlabel polysilicon 940 -3585 940 -3585 0 3
rlabel polysilicon 968 -3579 968 -3579 0 1
rlabel polysilicon 968 -3585 968 -3585 0 3
rlabel polysilicon 975 -3579 975 -3579 0 1
rlabel polysilicon 975 -3585 975 -3585 0 3
rlabel polysilicon 982 -3579 982 -3579 0 1
rlabel polysilicon 982 -3585 982 -3585 0 3
rlabel polysilicon 985 -3585 985 -3585 0 4
rlabel polysilicon 989 -3579 989 -3579 0 1
rlabel polysilicon 989 -3585 989 -3585 0 3
rlabel polysilicon 1038 -3579 1038 -3579 0 1
rlabel polysilicon 1038 -3585 1038 -3585 0 3
rlabel polysilicon 1052 -3579 1052 -3579 0 1
rlabel polysilicon 1052 -3585 1052 -3585 0 3
rlabel polysilicon 1083 -3585 1083 -3585 0 4
rlabel polysilicon 1087 -3579 1087 -3579 0 1
rlabel polysilicon 1087 -3585 1087 -3585 0 3
rlabel polysilicon 1108 -3579 1108 -3579 0 1
rlabel polysilicon 1108 -3585 1108 -3585 0 3
rlabel polysilicon 327 -3602 327 -3602 0 2
rlabel polysilicon 352 -3602 352 -3602 0 1
rlabel polysilicon 401 -3602 401 -3602 0 1
rlabel polysilicon 401 -3608 401 -3608 0 3
rlabel polysilicon 408 -3602 408 -3602 0 1
rlabel polysilicon 457 -3602 457 -3602 0 1
rlabel polysilicon 457 -3608 457 -3608 0 3
rlabel polysilicon 471 -3602 471 -3602 0 1
rlabel polysilicon 471 -3608 471 -3608 0 3
rlabel polysilicon 492 -3602 492 -3602 0 1
rlabel polysilicon 492 -3608 492 -3608 0 3
rlabel polysilicon 506 -3602 506 -3602 0 1
rlabel polysilicon 506 -3608 506 -3608 0 3
rlabel polysilicon 516 -3602 516 -3602 0 2
rlabel polysilicon 513 -3608 513 -3608 0 3
rlabel polysilicon 516 -3608 516 -3608 0 4
rlabel polysilicon 520 -3602 520 -3602 0 1
rlabel polysilicon 520 -3608 520 -3608 0 3
rlabel polysilicon 544 -3602 544 -3602 0 2
rlabel polysilicon 541 -3608 541 -3608 0 3
rlabel polysilicon 548 -3602 548 -3602 0 1
rlabel polysilicon 548 -3608 548 -3608 0 3
rlabel polysilicon 555 -3602 555 -3602 0 1
rlabel polysilicon 555 -3608 555 -3608 0 3
rlabel polysilicon 562 -3602 562 -3602 0 1
rlabel polysilicon 562 -3608 562 -3608 0 3
rlabel polysilicon 569 -3602 569 -3602 0 1
rlabel polysilicon 569 -3608 569 -3608 0 3
rlabel polysilicon 576 -3602 576 -3602 0 1
rlabel polysilicon 576 -3608 576 -3608 0 3
rlabel polysilicon 597 -3602 597 -3602 0 1
rlabel polysilicon 597 -3608 597 -3608 0 3
rlabel polysilicon 604 -3602 604 -3602 0 1
rlabel polysilicon 604 -3608 604 -3608 0 3
rlabel polysilicon 614 -3602 614 -3602 0 2
rlabel polysilicon 611 -3608 611 -3608 0 3
rlabel polysilicon 681 -3602 681 -3602 0 1
rlabel polysilicon 684 -3608 684 -3608 0 4
rlabel polysilicon 695 -3602 695 -3602 0 1
rlabel polysilicon 695 -3608 695 -3608 0 3
rlabel polysilicon 702 -3602 702 -3602 0 1
rlabel polysilicon 702 -3608 702 -3608 0 3
rlabel polysilicon 709 -3602 709 -3602 0 1
rlabel polysilicon 709 -3608 709 -3608 0 3
rlabel polysilicon 712 -3608 712 -3608 0 4
rlabel polysilicon 716 -3602 716 -3602 0 1
rlabel polysilicon 716 -3608 716 -3608 0 3
rlabel polysilicon 723 -3602 723 -3602 0 1
rlabel polysilicon 723 -3608 723 -3608 0 3
rlabel polysilicon 730 -3602 730 -3602 0 1
rlabel polysilicon 730 -3608 730 -3608 0 3
rlabel polysilicon 737 -3602 737 -3602 0 1
rlabel polysilicon 737 -3608 737 -3608 0 3
rlabel polysilicon 744 -3602 744 -3602 0 1
rlabel polysilicon 744 -3608 744 -3608 0 3
rlabel polysilicon 751 -3602 751 -3602 0 1
rlabel polysilicon 751 -3608 751 -3608 0 3
rlabel polysilicon 758 -3602 758 -3602 0 1
rlabel polysilicon 758 -3608 758 -3608 0 3
rlabel polysilicon 761 -3608 761 -3608 0 4
rlabel polysilicon 765 -3602 765 -3602 0 1
rlabel polysilicon 765 -3608 765 -3608 0 3
rlabel polysilicon 772 -3602 772 -3602 0 1
rlabel polysilicon 772 -3608 772 -3608 0 3
rlabel polysilicon 856 -3602 856 -3602 0 1
rlabel polysilicon 856 -3608 856 -3608 0 3
rlabel polysilicon 863 -3602 863 -3602 0 1
rlabel polysilicon 863 -3608 863 -3608 0 3
rlabel polysilicon 905 -3602 905 -3602 0 1
rlabel polysilicon 908 -3602 908 -3602 0 2
rlabel polysilicon 919 -3602 919 -3602 0 1
rlabel polysilicon 919 -3608 919 -3608 0 3
rlabel polysilicon 926 -3602 926 -3602 0 1
rlabel polysilicon 926 -3608 926 -3608 0 3
rlabel polysilicon 975 -3602 975 -3602 0 1
rlabel polysilicon 975 -3608 975 -3608 0 3
rlabel polysilicon 982 -3602 982 -3602 0 1
rlabel polysilicon 982 -3608 982 -3608 0 3
rlabel polysilicon 1031 -3602 1031 -3602 0 1
rlabel polysilicon 1031 -3608 1031 -3608 0 3
rlabel polysilicon 1045 -3602 1045 -3602 0 1
rlabel polysilicon 1045 -3608 1045 -3608 0 3
rlabel polysilicon 1052 -3602 1052 -3602 0 1
rlabel polysilicon 1052 -3608 1052 -3608 0 3
rlabel polysilicon 1108 -3602 1108 -3602 0 1
rlabel polysilicon 1108 -3608 1108 -3608 0 3
rlabel polysilicon 401 -3627 401 -3627 0 1
rlabel polysilicon 401 -3633 401 -3633 0 3
rlabel polysilicon 408 -3633 408 -3633 0 3
rlabel polysilicon 464 -3627 464 -3627 0 1
rlabel polysilicon 464 -3633 464 -3633 0 3
rlabel polysilicon 471 -3627 471 -3627 0 1
rlabel polysilicon 471 -3633 471 -3633 0 3
rlabel polysilicon 527 -3627 527 -3627 0 1
rlabel polysilicon 527 -3633 527 -3633 0 3
rlabel polysilicon 562 -3627 562 -3627 0 1
rlabel polysilicon 562 -3633 562 -3633 0 3
rlabel polysilicon 569 -3627 569 -3627 0 1
rlabel polysilicon 569 -3633 569 -3633 0 3
rlabel polysilicon 576 -3627 576 -3627 0 1
rlabel polysilicon 576 -3633 576 -3633 0 3
rlabel polysilicon 583 -3627 583 -3627 0 1
rlabel polysilicon 583 -3633 583 -3633 0 3
rlabel polysilicon 590 -3627 590 -3627 0 1
rlabel polysilicon 590 -3633 590 -3633 0 3
rlabel polysilicon 702 -3627 702 -3627 0 1
rlabel polysilicon 702 -3633 702 -3633 0 3
rlabel polysilicon 709 -3627 709 -3627 0 1
rlabel polysilicon 712 -3627 712 -3627 0 2
rlabel polysilicon 709 -3633 709 -3633 0 3
rlabel polysilicon 716 -3627 716 -3627 0 1
rlabel polysilicon 716 -3633 716 -3633 0 3
rlabel polysilicon 723 -3627 723 -3627 0 1
rlabel polysilicon 723 -3633 723 -3633 0 3
rlabel polysilicon 744 -3627 744 -3627 0 1
rlabel polysilicon 744 -3633 744 -3633 0 3
rlabel polysilicon 751 -3627 751 -3627 0 1
rlabel polysilicon 751 -3633 751 -3633 0 3
rlabel polysilicon 758 -3627 758 -3627 0 1
rlabel polysilicon 758 -3633 758 -3633 0 3
rlabel polysilicon 765 -3627 765 -3627 0 1
rlabel polysilicon 765 -3633 765 -3633 0 3
rlabel polysilicon 775 -3627 775 -3627 0 2
rlabel polysilicon 772 -3633 772 -3633 0 3
rlabel polysilicon 800 -3627 800 -3627 0 1
rlabel polysilicon 800 -3633 800 -3633 0 3
rlabel polysilicon 856 -3627 856 -3627 0 1
rlabel polysilicon 856 -3633 856 -3633 0 3
rlabel polysilicon 863 -3627 863 -3627 0 1
rlabel polysilicon 863 -3633 863 -3633 0 3
rlabel polysilicon 926 -3627 926 -3627 0 1
rlabel polysilicon 926 -3633 926 -3633 0 3
rlabel polysilicon 933 -3627 933 -3627 0 1
rlabel polysilicon 933 -3633 933 -3633 0 3
rlabel polysilicon 982 -3627 982 -3627 0 1
rlabel polysilicon 982 -3633 982 -3633 0 3
rlabel polysilicon 1003 -3627 1003 -3627 0 1
rlabel polysilicon 1003 -3633 1003 -3633 0 3
rlabel polysilicon 1031 -3627 1031 -3627 0 1
rlabel polysilicon 1031 -3633 1031 -3633 0 3
rlabel polysilicon 1052 -3633 1052 -3633 0 3
rlabel polysilicon 1055 -3633 1055 -3633 0 4
rlabel polysilicon 1059 -3627 1059 -3627 0 1
rlabel polysilicon 1059 -3633 1059 -3633 0 3
rlabel polysilicon 1080 -3627 1080 -3627 0 1
rlabel polysilicon 1080 -3633 1080 -3633 0 3
rlabel polysilicon 1108 -3627 1108 -3627 0 1
rlabel polysilicon 1108 -3633 1108 -3633 0 3
rlabel polysilicon 401 -3642 401 -3642 0 1
rlabel polysilicon 401 -3648 401 -3648 0 3
rlabel polysilicon 408 -3642 408 -3642 0 1
rlabel polysilicon 408 -3648 408 -3648 0 3
rlabel polysilicon 464 -3642 464 -3642 0 1
rlabel polysilicon 464 -3648 464 -3648 0 3
rlabel polysilicon 474 -3642 474 -3642 0 2
rlabel polysilicon 474 -3648 474 -3648 0 4
rlabel polysilicon 527 -3642 527 -3642 0 1
rlabel polysilicon 527 -3648 527 -3648 0 3
rlabel polysilicon 572 -3642 572 -3642 0 2
rlabel polysilicon 569 -3648 569 -3648 0 3
rlabel polysilicon 576 -3642 576 -3642 0 1
rlabel polysilicon 576 -3648 576 -3648 0 3
rlabel polysilicon 583 -3642 583 -3642 0 1
rlabel polysilicon 583 -3648 583 -3648 0 3
rlabel polysilicon 586 -3648 586 -3648 0 4
rlabel polysilicon 590 -3642 590 -3642 0 1
rlabel polysilicon 590 -3648 590 -3648 0 3
rlabel polysilicon 597 -3642 597 -3642 0 1
rlabel polysilicon 597 -3648 597 -3648 0 3
rlabel polysilicon 709 -3642 709 -3642 0 1
rlabel polysilicon 709 -3648 709 -3648 0 3
rlabel polysilicon 716 -3642 716 -3642 0 1
rlabel polysilicon 719 -3642 719 -3642 0 2
rlabel polysilicon 716 -3648 716 -3648 0 3
rlabel polysilicon 719 -3648 719 -3648 0 4
rlabel polysilicon 723 -3642 723 -3642 0 1
rlabel polysilicon 723 -3648 723 -3648 0 3
rlabel polysilicon 751 -3642 751 -3642 0 1
rlabel polysilicon 751 -3648 751 -3648 0 3
rlabel polysilicon 758 -3642 758 -3642 0 1
rlabel polysilicon 758 -3648 758 -3648 0 3
rlabel polysilicon 765 -3642 765 -3642 0 1
rlabel polysilicon 765 -3648 765 -3648 0 3
rlabel polysilicon 859 -3642 859 -3642 0 2
rlabel polysilicon 856 -3648 856 -3648 0 3
rlabel polysilicon 863 -3642 863 -3642 0 1
rlabel polysilicon 863 -3648 863 -3648 0 3
rlabel polysilicon 926 -3642 926 -3642 0 1
rlabel polysilicon 929 -3642 929 -3642 0 2
rlabel polysilicon 929 -3648 929 -3648 0 4
rlabel polysilicon 933 -3642 933 -3642 0 1
rlabel polysilicon 933 -3648 933 -3648 0 3
rlabel polysilicon 985 -3642 985 -3642 0 2
rlabel polysilicon 985 -3648 985 -3648 0 4
rlabel polysilicon 989 -3642 989 -3642 0 1
rlabel polysilicon 989 -3648 989 -3648 0 3
rlabel polysilicon 1031 -3642 1031 -3642 0 1
rlabel polysilicon 1034 -3642 1034 -3642 0 2
rlabel polysilicon 1094 -3642 1094 -3642 0 1
rlabel polysilicon 1094 -3648 1094 -3648 0 3
rlabel polysilicon 1111 -3642 1111 -3642 0 2
rlabel polysilicon 1108 -3648 1108 -3648 0 3
rlabel polysilicon 401 -3657 401 -3657 0 1
rlabel polysilicon 404 -3663 404 -3663 0 4
rlabel polysilicon 408 -3657 408 -3657 0 1
rlabel polysilicon 408 -3663 408 -3663 0 3
rlabel polysilicon 527 -3663 527 -3663 0 3
rlabel polysilicon 534 -3657 534 -3657 0 1
rlabel polysilicon 534 -3663 534 -3663 0 3
rlabel polysilicon 758 -3657 758 -3657 0 1
rlabel polysilicon 758 -3663 758 -3663 0 3
rlabel polysilicon 765 -3657 765 -3657 0 1
rlabel polysilicon 765 -3663 765 -3663 0 3
rlabel polysilicon 768 -3663 768 -3663 0 4
rlabel polysilicon 772 -3657 772 -3657 0 1
rlabel polysilicon 772 -3663 772 -3663 0 3
rlabel metal2 226 1 226 1 0 net=6047
rlabel metal2 366 1 366 1 0 net=2763
rlabel metal2 415 1 415 1 0 net=1753
rlabel metal2 590 1 590 1 0 net=7649
rlabel metal2 667 1 667 1 0 net=11501
rlabel metal2 705 1 705 1 0 net=11123
rlabel metal2 254 -1 254 -1 0 net=11889
rlabel metal2 401 -1 401 -1 0 net=10253
rlabel metal2 457 -1 457 -1 0 net=4171
rlabel metal2 492 -1 492 -1 0 net=6711
rlabel metal2 765 -1 765 -1 0 net=11437
rlabel metal2 803 -1 803 -1 0 net=10049
rlabel metal2 275 -3 275 -3 0 net=3753
rlabel metal2 506 -3 506 -3 0 net=7403
rlabel metal2 516 -3 516 -3 0 net=7095
rlabel metal2 534 -3 534 -3 0 net=3591
rlabel metal2 317 -5 317 -5 0 net=4443
rlabel metal2 429 -5 429 -5 0 net=6013
rlabel metal2 135 -16 135 -16 0 net=1879
rlabel metal2 303 -16 303 -16 0 net=4445
rlabel metal2 327 -16 327 -16 0 net=3861
rlabel metal2 383 -16 383 -16 0 net=7225
rlabel metal2 541 -16 541 -16 0 net=7551
rlabel metal2 565 -16 565 -16 0 net=4155
rlabel metal2 765 -16 765 -16 0 net=11439
rlabel metal2 765 -16 765 -16 0 net=11439
rlabel metal2 775 -16 775 -16 0 net=11393
rlabel metal2 821 -16 821 -16 0 net=11363
rlabel metal2 191 -18 191 -18 0 net=6049
rlabel metal2 310 -18 310 -18 0 net=6423
rlabel metal2 345 -18 345 -18 0 net=2765
rlabel metal2 373 -18 373 -18 0 net=3139
rlabel metal2 450 -18 450 -18 0 net=10255
rlabel metal2 527 -18 527 -18 0 net=7097
rlabel metal2 569 -18 569 -18 0 net=3593
rlabel metal2 632 -18 632 -18 0 net=12081
rlabel metal2 674 -18 674 -18 0 net=11503
rlabel metal2 782 -18 782 -18 0 net=10485
rlabel metal2 828 -18 828 -18 0 net=11125
rlabel metal2 205 -20 205 -20 0 net=11891
rlabel metal2 331 -20 331 -20 0 net=7517
rlabel metal2 488 -20 488 -20 0 net=11647
rlabel metal2 569 -20 569 -20 0 net=7999
rlabel metal2 842 -20 842 -20 0 net=10051
rlabel metal2 212 -22 212 -22 0 net=3755
rlabel metal2 331 -22 331 -22 0 net=5899
rlabel metal2 408 -22 408 -22 0 net=9099
rlabel metal2 471 -22 471 -22 0 net=4173
rlabel metal2 471 -22 471 -22 0 net=4173
rlabel metal2 492 -22 492 -22 0 net=6713
rlabel metal2 492 -22 492 -22 0 net=6713
rlabel metal2 506 -22 506 -22 0 net=7405
rlabel metal2 576 -22 576 -22 0 net=7651
rlabel metal2 635 -22 635 -22 0 net=4993
rlabel metal2 660 -22 660 -22 0 net=7533
rlabel metal2 226 -24 226 -24 0 net=10909
rlabel metal2 352 -24 352 -24 0 net=1755
rlabel metal2 436 -24 436 -24 0 net=6014
rlabel metal2 450 -24 450 -24 0 net=6553
rlabel metal2 639 -24 639 -24 0 net=10367
rlabel metal2 254 -26 254 -26 0 net=5035
rlabel metal2 376 -26 376 -26 0 net=7639
rlabel metal2 443 -26 443 -26 0 net=298
rlabel metal2 299 -28 299 -28 0 net=4463
rlabel metal2 457 -28 457 -28 0 net=5527
rlabel metal2 317 -30 317 -30 0 net=3343
rlabel metal2 618 -30 618 -30 0 net=9841
rlabel metal2 387 -32 387 -32 0 net=3585
rlabel metal2 401 -32 401 -32 0 net=3415
rlabel metal2 618 -32 618 -32 0 net=11751
rlabel metal2 359 -34 359 -34 0 net=2561
rlabel metal2 79 -45 79 -45 0 net=9061
rlabel metal2 268 -45 268 -45 0 net=5901
rlabel metal2 345 -45 345 -45 0 net=2767
rlabel metal2 345 -45 345 -45 0 net=2767
rlabel metal2 380 -45 380 -45 0 net=3862
rlabel metal2 450 -45 450 -45 0 net=6393
rlabel metal2 618 -45 618 -45 0 net=6769
rlabel metal2 856 -45 856 -45 0 net=10053
rlabel metal2 877 -45 877 -45 0 net=11127
rlabel metal2 919 -45 919 -45 0 net=11365
rlabel metal2 100 -47 100 -47 0 net=1881
rlabel metal2 142 -47 142 -47 0 net=1468
rlabel metal2 380 -47 380 -47 0 net=3911
rlabel metal2 576 -47 576 -47 0 net=7653
rlabel metal2 632 -47 632 -47 0 net=4995
rlabel metal2 667 -47 667 -47 0 net=12083
rlabel metal2 758 -47 758 -47 0 net=12111
rlabel metal2 128 -49 128 -49 0 net=6565
rlabel metal2 278 -49 278 -49 0 net=4446
rlabel metal2 310 -49 310 -49 0 net=3351
rlabel metal2 310 -49 310 -49 0 net=3351
rlabel metal2 324 -49 324 -49 0 net=6477
rlabel metal2 478 -49 478 -49 0 net=7519
rlabel metal2 639 -49 639 -49 0 net=9843
rlabel metal2 695 -49 695 -49 0 net=11505
rlabel metal2 761 -49 761 -49 0 net=11149
rlabel metal2 149 -51 149 -51 0 net=3345
rlabel metal2 397 -51 397 -51 0 net=4059
rlabel metal2 408 -51 408 -51 0 net=9101
rlabel metal2 541 -51 541 -51 0 net=7099
rlabel metal2 576 -51 576 -51 0 net=3595
rlabel metal2 590 -51 590 -51 0 net=6729
rlabel metal2 660 -51 660 -51 0 net=7535
rlabel metal2 702 -51 702 -51 0 net=10369
rlabel metal2 765 -51 765 -51 0 net=11441
rlabel metal2 786 -51 786 -51 0 net=11753
rlabel metal2 156 -53 156 -53 0 net=5037
rlabel metal2 289 -53 289 -53 0 net=10249
rlabel metal2 422 -53 422 -53 0 net=7640
rlabel metal2 485 -53 485 -53 0 net=6091
rlabel metal2 702 -53 702 -53 0 net=7521
rlabel metal2 163 -55 163 -55 0 net=1709
rlabel metal2 184 -55 184 -55 0 net=6051
rlabel metal2 219 -55 219 -55 0 net=3527
rlabel metal2 464 -55 464 -55 0 net=12121
rlabel metal2 709 -55 709 -55 0 net=4157
rlabel metal2 793 -55 793 -55 0 net=10487
rlabel metal2 170 -57 170 -57 0 net=7379
rlabel metal2 303 -57 303 -57 0 net=2563
rlabel metal2 366 -57 366 -57 0 net=8977
rlabel metal2 499 -57 499 -57 0 net=8001
rlabel metal2 625 -57 625 -57 0 net=8039
rlabel metal2 800 -57 800 -57 0 net=11395
rlabel metal2 177 -59 177 -59 0 net=7781
rlabel metal2 222 -59 222 -59 0 net=5141
rlabel metal2 415 -59 415 -59 0 net=4465
rlabel metal2 436 -59 436 -59 0 net=4175
rlabel metal2 520 -59 520 -59 0 net=10257
rlabel metal2 177 -61 177 -61 0 net=6491
rlabel metal2 527 -61 527 -61 0 net=6555
rlabel metal2 555 -61 555 -61 0 net=11649
rlabel metal2 180 -63 180 -63 0 net=11892
rlabel metal2 226 -63 226 -63 0 net=10911
rlabel metal2 261 -63 261 -63 0 net=6369
rlabel metal2 317 -63 317 -63 0 net=1757
rlabel metal2 369 -63 369 -63 0 net=8127
rlabel metal2 527 -63 527 -63 0 net=5671
rlabel metal2 191 -65 191 -65 0 net=3757
rlabel metal2 226 -65 226 -65 0 net=11179
rlabel metal2 646 -65 646 -65 0 net=5529
rlabel metal2 205 -67 205 -67 0 net=3141
rlabel metal2 415 -67 415 -67 0 net=3417
rlabel metal2 534 -67 534 -67 0 net=7227
rlabel metal2 681 -67 681 -67 0 net=11813
rlabel metal2 229 -69 229 -69 0 net=6357
rlabel metal2 450 -69 450 -69 0 net=1376
rlabel metal2 513 -69 513 -69 0 net=7407
rlabel metal2 548 -69 548 -69 0 net=7553
rlabel metal2 569 -69 569 -69 0 net=11955
rlabel metal2 646 -69 646 -69 0 net=9771
rlabel metal2 243 -71 243 -71 0 net=2733
rlabel metal2 369 -71 369 -71 0 net=1389
rlabel metal2 331 -73 331 -73 0 net=8661
rlabel metal2 338 -75 338 -75 0 net=6425
rlabel metal2 457 -75 457 -75 0 net=5943
rlabel metal2 338 -77 338 -77 0 net=6907
rlabel metal2 373 -79 373 -79 0 net=3587
rlabel metal2 492 -79 492 -79 0 net=6715
rlabel metal2 548 -79 548 -79 0 net=8223
rlabel metal2 492 -81 492 -81 0 net=6687
rlabel metal2 593 -83 593 -83 0 net=8783
rlabel metal2 79 -94 79 -94 0 net=9062
rlabel metal2 418 -94 418 -94 0 net=8219
rlabel metal2 814 -94 814 -94 0 net=10489
rlabel metal2 856 -94 856 -94 0 net=11755
rlabel metal2 940 -94 940 -94 0 net=3449
rlabel metal2 114 -96 114 -96 0 net=6908
rlabel metal2 352 -96 352 -96 0 net=2735
rlabel metal2 432 -96 432 -96 0 net=10258
rlabel metal2 730 -96 730 -96 0 net=11442
rlabel metal2 842 -96 842 -96 0 net=10425
rlabel metal2 968 -96 968 -96 0 net=11367
rlabel metal2 100 -98 100 -98 0 net=1883
rlabel metal2 128 -98 128 -98 0 net=6566
rlabel metal2 250 -98 250 -98 0 net=8163
rlabel metal2 744 -98 744 -98 0 net=10371
rlabel metal2 870 -98 870 -98 0 net=12113
rlabel metal2 100 -100 100 -100 0 net=961
rlabel metal2 149 -100 149 -100 0 net=3346
rlabel metal2 352 -100 352 -100 0 net=3419
rlabel metal2 443 -100 443 -100 0 net=7689
rlabel metal2 744 -100 744 -100 0 net=4159
rlabel metal2 863 -100 863 -100 0 net=10055
rlabel metal2 891 -100 891 -100 0 net=11151
rlabel metal2 156 -102 156 -102 0 net=5038
rlabel metal2 240 -102 240 -102 0 net=4093
rlabel metal2 446 -102 446 -102 0 net=8224
rlabel metal2 558 -102 558 -102 0 net=6345
rlabel metal2 163 -104 163 -104 0 net=1711
rlabel metal2 163 -104 163 -104 0 net=1711
rlabel metal2 205 -104 205 -104 0 net=3143
rlabel metal2 453 -104 453 -104 0 net=11650
rlabel metal2 723 -104 723 -104 0 net=12085
rlabel metal2 905 -104 905 -104 0 net=11129
rlabel metal2 205 -106 205 -106 0 net=4837
rlabel metal2 282 -106 282 -106 0 net=3352
rlabel metal2 324 -106 324 -106 0 net=6479
rlabel metal2 506 -106 506 -106 0 net=9103
rlabel metal2 793 -106 793 -106 0 net=11815
rlabel metal2 149 -108 149 -108 0 net=5717
rlabel metal2 292 -108 292 -108 0 net=6426
rlabel metal2 499 -108 499 -108 0 net=8002
rlabel metal2 513 -108 513 -108 0 net=6717
rlabel metal2 642 -108 642 -108 0 net=10795
rlabel metal2 145 -110 145 -110 0 net=4291
rlabel metal2 513 -110 513 -110 0 net=1623
rlabel metal2 688 -110 688 -110 0 net=9845
rlabel metal2 821 -110 821 -110 0 net=11397
rlabel metal2 170 -112 170 -112 0 net=7380
rlabel metal2 296 -112 296 -112 0 net=925
rlabel metal2 562 -112 562 -112 0 net=7101
rlabel metal2 646 -112 646 -112 0 net=9773
rlabel metal2 660 -112 660 -112 0 net=7229
rlabel metal2 170 -114 170 -114 0 net=11419
rlabel metal2 485 -114 485 -114 0 net=6093
rlabel metal2 569 -114 569 -114 0 net=12135
rlabel metal2 215 -116 215 -116 0 net=4091
rlabel metal2 268 -116 268 -116 0 net=5902
rlabel metal2 303 -116 303 -116 0 net=2564
rlabel metal2 569 -116 569 -116 0 net=4997
rlabel metal2 646 -116 646 -116 0 net=6731
rlabel metal2 660 -116 660 -116 0 net=6809
rlabel metal2 751 -116 751 -116 0 net=11507
rlabel metal2 177 -118 177 -118 0 net=1144
rlabel metal2 310 -118 310 -118 0 net=1759
rlabel metal2 324 -118 324 -118 0 net=3913
rlabel metal2 471 -118 471 -118 0 net=6725
rlabel metal2 653 -118 653 -118 0 net=6771
rlabel metal2 177 -120 177 -120 0 net=6371
rlabel metal2 268 -120 268 -120 0 net=4229
rlabel metal2 359 -120 359 -120 0 net=5143
rlabel metal2 548 -120 548 -120 0 net=5965
rlabel metal2 754 -120 754 -120 0 net=9571
rlabel metal2 191 -122 191 -122 0 net=3759
rlabel metal2 278 -122 278 -122 0 net=1070
rlabel metal2 345 -122 345 -122 0 net=2769
rlabel metal2 471 -122 471 -122 0 net=7520
rlabel metal2 618 -122 618 -122 0 net=11957
rlabel metal2 142 -124 142 -124 0 net=7583
rlabel metal2 450 -124 450 -124 0 net=251
rlabel metal2 649 -124 649 -124 0 net=1
rlabel metal2 184 -126 184 -126 0 net=6053
rlabel metal2 212 -126 212 -126 0 net=3203
rlabel metal2 436 -126 436 -126 0 net=4177
rlabel metal2 534 -126 534 -126 0 net=7409
rlabel metal2 667 -126 667 -126 0 net=7537
rlabel metal2 184 -128 184 -128 0 net=12053
rlabel metal2 555 -128 555 -128 0 net=7555
rlabel metal2 674 -128 674 -128 0 net=8785
rlabel metal2 198 -130 198 -130 0 net=7783
rlabel metal2 254 -130 254 -130 0 net=10913
rlabel metal2 457 -130 457 -130 0 net=5945
rlabel metal2 583 -130 583 -130 0 net=11181
rlabel metal2 198 -132 198 -132 0 net=3529
rlabel metal2 240 -132 240 -132 0 net=3231
rlabel metal2 285 -132 285 -132 0 net=5955
rlabel metal2 457 -132 457 -132 0 net=5957
rlabel metal2 583 -132 583 -132 0 net=6395
rlabel metal2 674 -132 674 -132 0 net=3073
rlabel metal2 765 -132 765 -132 0 net=8041
rlabel metal2 219 -134 219 -134 0 net=2311
rlabel metal2 285 -134 285 -134 0 net=3211
rlabel metal2 492 -134 492 -134 0 net=6689
rlabel metal2 688 -134 688 -134 0 net=7523
rlabel metal2 716 -134 716 -134 0 net=5531
rlabel metal2 422 -136 422 -136 0 net=4467
rlabel metal2 520 -136 520 -136 0 net=8129
rlabel metal2 401 -138 401 -138 0 net=4061
rlabel metal2 520 -138 520 -138 0 net=5673
rlabel metal2 590 -138 590 -138 0 net=8662
rlabel metal2 695 -138 695 -138 0 net=12123
rlabel metal2 373 -140 373 -140 0 net=3589
rlabel metal2 429 -140 429 -140 0 net=6359
rlabel metal2 597 -140 597 -140 0 net=7655
rlabel metal2 289 -142 289 -142 0 net=10251
rlabel metal2 429 -142 429 -142 0 net=9451
rlabel metal2 233 -144 233 -144 0 net=7119
rlabel metal2 478 -144 478 -144 0 net=8979
rlabel metal2 681 -144 681 -144 0 net=9341
rlabel metal2 478 -146 478 -146 0 net=3597
rlabel metal2 702 -146 702 -146 0 net=7617
rlabel metal2 464 -148 464 -148 0 net=6493
rlabel metal2 464 -150 464 -150 0 net=11073
rlabel metal2 541 -152 541 -152 0 net=6557
rlabel metal2 488 -154 488 -154 0 net=5389
rlabel metal2 72 -165 72 -165 0 net=8211
rlabel metal2 450 -165 450 -165 0 net=4178
rlabel metal2 495 -165 495 -165 0 net=8980
rlabel metal2 618 -165 618 -165 0 net=12086
rlabel metal2 870 -165 870 -165 0 net=10057
rlabel metal2 954 -165 954 -165 0 net=12115
rlabel metal2 100 -167 100 -167 0 net=2569
rlabel metal2 135 -167 135 -167 0 net=3421
rlabel metal2 390 -167 390 -167 0 net=5956
rlabel metal2 453 -167 453 -167 0 net=6360
rlabel metal2 541 -167 541 -167 0 net=5391
rlabel metal2 618 -167 618 -167 0 net=5533
rlabel metal2 730 -167 730 -167 0 net=8165
rlabel metal2 100 -169 100 -169 0 net=1885
rlabel metal2 124 -169 124 -169 0 net=11857
rlabel metal2 107 -171 107 -171 0 net=9145
rlabel metal2 877 -171 877 -171 0 net=11183
rlabel metal2 110 -173 110 -173 0 net=994
rlabel metal2 457 -173 457 -173 0 net=5959
rlabel metal2 621 -173 621 -173 0 net=8225
rlabel metal2 114 -175 114 -175 0 net=4469
rlabel metal2 509 -175 509 -175 0 net=12071
rlabel metal2 149 -177 149 -177 0 net=5718
rlabel metal2 254 -177 254 -177 0 net=4005
rlabel metal2 467 -177 467 -177 0 net=3074
rlabel metal2 695 -177 695 -177 0 net=7749
rlabel metal2 730 -177 730 -177 0 net=7231
rlabel metal2 1003 -177 1003 -177 0 net=11369
rlabel metal2 156 -179 156 -179 0 net=1397
rlabel metal2 506 -179 506 -179 0 net=6961
rlabel metal2 695 -179 695 -179 0 net=7539
rlabel metal2 996 -179 996 -179 0 net=11245
rlabel metal2 170 -181 170 -181 0 net=11420
rlabel metal2 310 -181 310 -181 0 net=1760
rlabel metal2 352 -181 352 -181 0 net=2649
rlabel metal2 506 -181 506 -181 0 net=5675
rlabel metal2 625 -181 625 -181 0 net=6719
rlabel metal2 625 -181 625 -181 0 net=6719
rlabel metal2 632 -181 632 -181 0 net=6727
rlabel metal2 786 -181 786 -181 0 net=8043
rlabel metal2 884 -181 884 -181 0 net=11959
rlabel metal2 166 -183 166 -183 0 net=7427
rlabel metal2 562 -183 562 -183 0 net=6095
rlabel metal2 667 -183 667 -183 0 net=7557
rlabel metal2 828 -183 828 -183 0 net=10797
rlabel metal2 173 -185 173 -185 0 net=493
rlabel metal2 310 -185 310 -185 0 net=1955
rlabel metal2 488 -185 488 -185 0 net=409
rlabel metal2 835 -185 835 -185 0 net=10373
rlabel metal2 891 -185 891 -185 0 net=11399
rlabel metal2 184 -187 184 -187 0 net=12054
rlabel metal2 471 -187 471 -187 0 net=3229
rlabel metal2 562 -187 562 -187 0 net=5509
rlabel metal2 814 -187 814 -187 0 net=9847
rlabel metal2 898 -187 898 -187 0 net=11509
rlabel metal2 163 -189 163 -189 0 net=1713
rlabel metal2 198 -189 198 -189 0 net=3531
rlabel metal2 198 -189 198 -189 0 net=3531
rlabel metal2 208 -189 208 -189 0 net=7784
rlabel metal2 219 -189 219 -189 0 net=2313
rlabel metal2 261 -189 261 -189 0 net=3761
rlabel metal2 639 -189 639 -189 0 net=7103
rlabel metal2 814 -189 814 -189 0 net=7699
rlabel metal2 856 -189 856 -189 0 net=11075
rlabel metal2 163 -191 163 -191 0 net=9017
rlabel metal2 905 -191 905 -191 0 net=11817
rlabel metal2 177 -193 177 -193 0 net=6373
rlabel metal2 667 -193 667 -193 0 net=4161
rlabel metal2 758 -193 758 -193 0 net=8221
rlabel metal2 912 -193 912 -193 0 net=12125
rlabel metal2 177 -195 177 -195 0 net=4231
rlabel metal2 324 -195 324 -195 0 net=3915
rlabel metal2 653 -195 653 -195 0 net=6773
rlabel metal2 779 -195 779 -195 0 net=9105
rlabel metal2 919 -195 919 -195 0 net=11757
rlabel metal2 121 -197 121 -197 0 net=1703
rlabel metal2 380 -197 380 -197 0 net=6481
rlabel metal2 597 -197 597 -197 0 net=6559
rlabel metal2 793 -197 793 -197 0 net=9453
rlabel metal2 926 -197 926 -197 0 net=11131
rlabel metal2 212 -199 212 -199 0 net=3205
rlabel metal2 380 -199 380 -199 0 net=4063
rlabel metal2 432 -199 432 -199 0 net=6103
rlabel metal2 712 -199 712 -199 0 net=1
rlabel metal2 821 -199 821 -199 0 net=9573
rlabel metal2 933 -199 933 -199 0 net=12137
rlabel metal2 219 -201 219 -201 0 net=1983
rlabel metal2 282 -201 282 -201 0 net=10252
rlabel metal2 394 -201 394 -201 0 net=2736
rlabel metal2 737 -201 737 -201 0 net=7619
rlabel metal2 842 -201 842 -201 0 net=10427
rlabel metal2 943 -201 943 -201 0 net=10689
rlabel metal2 961 -201 961 -201 0 net=11153
rlabel metal2 222 -203 222 -203 0 net=2593
rlabel metal2 331 -203 331 -203 0 net=3213
rlabel metal2 464 -203 464 -203 0 net=3599
rlabel metal2 611 -203 611 -203 0 net=7411
rlabel metal2 754 -203 754 -203 0 net=10507
rlabel metal2 947 -203 947 -203 0 net=11185
rlabel metal2 226 -205 226 -205 0 net=4092
rlabel metal2 285 -205 285 -205 0 net=1207
rlabel metal2 681 -205 681 -205 0 net=10733
rlabel metal2 968 -205 968 -205 0 net=6347
rlabel metal2 226 -207 226 -207 0 net=5967
rlabel metal2 681 -207 681 -207 0 net=10579
rlabel metal2 975 -207 975 -207 0 net=3450
rlabel metal2 240 -209 240 -209 0 net=3233
rlabel metal2 289 -209 289 -209 0 net=1943
rlabel metal2 705 -209 705 -209 0 net=10853
rlabel metal2 250 -211 250 -211 0 net=1155
rlabel metal2 317 -211 317 -211 0 net=10915
rlabel metal2 261 -213 261 -213 0 net=2267
rlabel metal2 478 -213 478 -213 0 net=9483
rlabel metal2 271 -215 271 -215 0 net=1813
rlabel metal2 359 -215 359 -215 0 net=2771
rlabel metal2 394 -215 394 -215 0 net=4293
rlabel metal2 415 -215 415 -215 0 net=1625
rlabel metal2 548 -215 548 -215 0 net=6397
rlabel metal2 772 -215 772 -215 0 net=8787
rlabel metal2 849 -215 849 -215 0 net=10491
rlabel metal2 205 -217 205 -217 0 net=4839
rlabel metal2 366 -217 366 -217 0 net=2949
rlabel metal2 723 -217 723 -217 0 net=7657
rlabel metal2 205 -219 205 -219 0 net=1388
rlabel metal2 513 -219 513 -219 0 net=6810
rlabel metal2 765 -219 765 -219 0 net=9343
rlabel metal2 257 -221 257 -221 0 net=6059
rlabel metal2 604 -221 604 -221 0 net=6691
rlabel metal2 765 -221 765 -221 0 net=7695
rlabel metal2 345 -223 345 -223 0 net=7584
rlabel metal2 646 -223 646 -223 0 net=6733
rlabel metal2 278 -225 278 -225 0 net=2989
rlabel metal2 401 -225 401 -225 0 net=3590
rlabel metal2 569 -225 569 -225 0 net=4999
rlabel metal2 401 -227 401 -227 0 net=7645
rlabel metal2 534 -229 534 -229 0 net=5947
rlabel metal2 576 -229 576 -229 0 net=6495
rlabel metal2 233 -231 233 -231 0 net=7121
rlabel metal2 191 -233 191 -233 0 net=6055
rlabel metal2 534 -233 534 -233 0 net=9774
rlabel metal2 191 -235 191 -235 0 net=1845
rlabel metal2 800 -235 800 -235 0 net=8131
rlabel metal2 709 -237 709 -237 0 net=7691
rlabel metal2 387 -239 387 -239 0 net=7491
rlabel metal2 387 -241 387 -241 0 net=5145
rlabel metal2 443 -243 443 -243 0 net=4095
rlabel metal2 296 -245 296 -245 0 net=101
rlabel metal2 296 -247 296 -247 0 net=3145
rlabel metal2 338 -249 338 -249 0 net=11975
rlabel metal2 54 -260 54 -260 0 net=531
rlabel metal2 296 -260 296 -260 0 net=3147
rlabel metal2 481 -260 481 -260 0 net=7122
rlabel metal2 614 -260 614 -260 0 net=11184
rlabel metal2 1038 -260 1038 -260 0 net=11155
rlabel metal2 72 -262 72 -262 0 net=8212
rlabel metal2 124 -262 124 -262 0 net=379
rlabel metal2 219 -262 219 -262 0 net=9106
rlabel metal2 947 -262 947 -262 0 net=10581
rlabel metal2 1052 -262 1052 -262 0 net=11859
rlabel metal2 79 -264 79 -264 0 net=11029
rlabel metal2 86 -266 86 -266 0 net=1887
rlabel metal2 110 -266 110 -266 0 net=1181
rlabel metal2 345 -266 345 -266 0 net=2991
rlabel metal2 481 -266 481 -266 0 net=8222
rlabel metal2 898 -266 898 -266 0 net=9575
rlabel metal2 954 -266 954 -266 0 net=10691
rlabel metal2 93 -268 93 -268 0 net=3371
rlabel metal2 635 -268 635 -268 0 net=10929
rlabel metal2 100 -270 100 -270 0 net=2773
rlabel metal2 401 -270 401 -270 0 net=3230
rlabel metal2 485 -270 485 -270 0 net=5676
rlabel metal2 516 -270 516 -270 0 net=6728
rlabel metal2 726 -270 726 -270 0 net=10921
rlabel metal2 124 -272 124 -272 0 net=9241
rlabel metal2 1059 -272 1059 -272 0 net=11371
rlabel metal2 128 -274 128 -274 0 net=2571
rlabel metal2 142 -274 142 -274 0 net=1847
rlabel metal2 219 -274 219 -274 0 net=5001
rlabel metal2 663 -274 663 -274 0 net=11510
rlabel metal2 1073 -274 1073 -274 0 net=11961
rlabel metal2 128 -276 128 -276 0 net=4703
rlabel metal2 240 -276 240 -276 0 net=2269
rlabel metal2 289 -276 289 -276 0 net=1945
rlabel metal2 359 -276 359 -276 0 net=4841
rlabel metal2 457 -276 457 -276 0 net=3917
rlabel metal2 530 -276 530 -276 0 net=158
rlabel metal2 849 -276 849 -276 0 net=9345
rlabel metal2 954 -276 954 -276 0 net=8227
rlabel metal2 149 -278 149 -278 0 net=6057
rlabel metal2 254 -278 254 -278 0 net=4006
rlabel metal2 604 -278 604 -278 0 net=10798
rlabel metal2 1080 -278 1080 -278 0 net=12073
rlabel metal2 156 -280 156 -280 0 net=5677
rlabel metal2 488 -280 488 -280 0 net=9041
rlabel metal2 1087 -280 1087 -280 0 net=12117
rlabel metal2 163 -282 163 -282 0 net=3762
rlabel metal2 467 -282 467 -282 0 net=8463
rlabel metal2 1094 -282 1094 -282 0 net=12139
rlabel metal2 82 -284 82 -284 0 net=3025
rlabel metal2 492 -284 492 -284 0 net=7412
rlabel metal2 744 -284 744 -284 0 net=7527
rlabel metal2 877 -284 877 -284 0 net=9485
rlabel metal2 163 -286 163 -286 0 net=1627
rlabel metal2 541 -286 541 -286 0 net=7232
rlabel metal2 765 -286 765 -286 0 net=11963
rlabel metal2 184 -288 184 -288 0 net=1715
rlabel metal2 198 -288 198 -288 0 net=3533
rlabel metal2 212 -288 212 -288 0 net=3207
rlabel metal2 513 -288 513 -288 0 net=5661
rlabel metal2 544 -288 544 -288 0 net=10781
rlabel metal2 58 -290 58 -290 0 net=4913
rlabel metal2 254 -290 254 -290 0 net=5147
rlabel metal2 408 -290 408 -290 0 net=6061
rlabel metal2 768 -290 768 -290 0 net=9454
rlabel metal2 933 -290 933 -290 0 net=10509
rlabel metal2 107 -292 107 -292 0 net=5167
rlabel metal2 268 -292 268 -292 0 net=1985
rlabel metal2 296 -292 296 -292 0 net=1553
rlabel metal2 320 -292 320 -292 0 net=6374
rlabel metal2 646 -292 646 -292 0 net=6497
rlabel metal2 779 -292 779 -292 0 net=7621
rlabel metal2 884 -292 884 -292 0 net=10375
rlabel metal2 107 -294 107 -294 0 net=3235
rlabel metal2 303 -294 303 -294 0 net=2595
rlabel metal2 387 -294 387 -294 0 net=6945
rlabel metal2 548 -294 548 -294 0 net=6398
rlabel metal2 597 -294 597 -294 0 net=6105
rlabel metal2 751 -294 751 -294 0 net=7647
rlabel metal2 891 -294 891 -294 0 net=9849
rlabel metal2 114 -296 114 -296 0 net=4471
rlabel metal2 562 -296 562 -296 0 net=5511
rlabel metal2 625 -296 625 -296 0 net=6721
rlabel metal2 702 -296 702 -296 0 net=7105
rlabel metal2 831 -296 831 -296 0 net=11186
rlabel metal2 1003 -296 1003 -296 0 net=11247
rlabel metal2 135 -298 135 -298 0 net=3423
rlabel metal2 247 -298 247 -298 0 net=2315
rlabel metal2 275 -298 275 -298 0 net=3215
rlabel metal2 471 -298 471 -298 0 net=6633
rlabel metal2 786 -298 786 -298 0 net=7697
rlabel metal2 177 -300 177 -300 0 net=4233
rlabel metal2 415 -300 415 -300 0 net=2891
rlabel metal2 569 -300 569 -300 0 net=5949
rlabel metal2 632 -300 632 -300 0 net=6097
rlabel metal2 772 -300 772 -300 0 net=7659
rlabel metal2 940 -300 940 -300 0 net=10059
rlabel metal2 1010 -300 1010 -300 0 net=11133
rlabel metal2 177 -302 177 -302 0 net=4529
rlabel metal2 499 -302 499 -302 0 net=4097
rlabel metal2 569 -302 569 -302 0 net=7692
rlabel metal2 807 -302 807 -302 0 net=8133
rlabel metal2 236 -304 236 -304 0 net=8069
rlabel metal2 968 -304 968 -304 0 net=10855
rlabel metal2 303 -306 303 -306 0 net=4037
rlabel metal2 513 -306 513 -306 0 net=8655
rlabel metal2 1017 -306 1017 -306 0 net=11401
rlabel metal2 114 -308 114 -308 0 net=5193
rlabel metal2 520 -308 520 -308 0 net=7429
rlabel metal2 793 -308 793 -308 0 net=7751
rlabel metal2 968 -308 968 -308 0 net=8167
rlabel metal2 317 -310 317 -310 0 net=2651
rlabel metal2 366 -310 366 -310 0 net=2951
rlabel metal2 464 -310 464 -310 0 net=3601
rlabel metal2 520 -310 520 -310 0 net=6483
rlabel metal2 576 -310 576 -310 0 net=5285
rlabel metal2 814 -310 814 -310 0 net=7701
rlabel metal2 961 -310 961 -310 0 net=10735
rlabel metal2 310 -312 310 -312 0 net=1957
rlabel metal2 404 -312 404 -312 0 net=8649
rlabel metal2 975 -312 975 -312 0 net=10917
rlabel metal2 310 -314 310 -314 0 net=1705
rlabel metal2 485 -314 485 -314 0 net=2575
rlabel metal2 821 -314 821 -314 0 net=8789
rlabel metal2 863 -314 863 -314 0 net=8045
rlabel metal2 982 -314 982 -314 0 net=11077
rlabel metal2 324 -316 324 -316 0 net=1815
rlabel metal2 527 -316 527 -316 0 net=11573
rlabel metal2 583 -318 583 -318 0 net=11976
rlabel metal2 632 -320 632 -320 0 net=12126
rlabel metal2 586 -322 586 -322 0 net=10465
rlabel metal2 586 -324 586 -324 0 net=8135
rlabel metal2 989 -324 989 -324 0 net=11819
rlabel metal2 639 -326 639 -326 0 net=4163
rlabel metal2 674 -326 674 -326 0 net=6963
rlabel metal2 835 -326 835 -326 0 net=9019
rlabel metal2 607 -328 607 -328 0 net=7257
rlabel metal2 842 -328 842 -328 0 net=6349
rlabel metal2 611 -330 611 -330 0 net=5561
rlabel metal2 684 -330 684 -330 0 net=8445
rlabel metal2 870 -330 870 -330 0 net=9147
rlabel metal2 1024 -330 1024 -330 0 net=11759
rlabel metal2 72 -332 72 -332 0 net=4919
rlabel metal2 618 -332 618 -332 0 net=5535
rlabel metal2 688 -332 688 -332 0 net=7559
rlabel metal2 919 -332 919 -332 0 net=10493
rlabel metal2 450 -334 450 -334 0 net=5741
rlabel metal2 653 -334 653 -334 0 net=6561
rlabel metal2 695 -334 695 -334 0 net=7541
rlabel metal2 926 -334 926 -334 0 net=10429
rlabel metal2 226 -336 226 -336 0 net=5969
rlabel metal2 709 -336 709 -336 0 net=7493
rlabel metal2 226 -338 226 -338 0 net=4353
rlabel metal2 446 -338 446 -338 0 net=4219
rlabel metal2 488 -338 488 -338 0 net=7795
rlabel metal2 555 -340 555 -340 0 net=5393
rlabel metal2 660 -340 660 -340 0 net=6693
rlabel metal2 719 -340 719 -340 0 net=8283
rlabel metal2 394 -342 394 -342 0 net=4295
rlabel metal2 590 -342 590 -342 0 net=5961
rlabel metal2 723 -342 723 -342 0 net=6735
rlabel metal2 845 -342 845 -342 0 net=8987
rlabel metal2 173 -344 173 -344 0 net=4357
rlabel metal2 590 -344 590 -344 0 net=11187
rlabel metal2 758 -346 758 -346 0 net=6775
rlabel metal2 380 -348 380 -348 0 net=4065
rlabel metal2 786 -348 786 -348 0 net=8025
rlabel metal2 170 -350 170 -350 0 net=3173
rlabel metal2 51 -352 51 -352 0 net=8137
rlabel metal2 58 -363 58 -363 0 net=7698
rlabel metal2 1227 -363 1227 -363 0 net=11373
rlabel metal2 1332 -363 1332 -363 0 net=11633
rlabel metal2 65 -365 65 -365 0 net=5679
rlabel metal2 366 -365 366 -365 0 net=5663
rlabel metal2 548 -365 548 -365 0 net=4473
rlabel metal2 548 -365 548 -365 0 net=4473
rlabel metal2 558 -365 558 -365 0 net=7660
rlabel metal2 919 -365 919 -365 0 net=7797
rlabel metal2 79 -367 79 -367 0 net=6375
rlabel metal2 96 -367 96 -367 0 net=8136
rlabel metal2 1038 -367 1038 -367 0 net=9043
rlabel metal2 1300 -367 1300 -367 0 net=11289
rlabel metal2 114 -369 114 -369 0 net=5194
rlabel metal2 485 -369 485 -369 0 net=4066
rlabel metal2 786 -369 786 -369 0 net=11248
rlabel metal2 1234 -369 1234 -369 0 net=11403
rlabel metal2 124 -371 124 -371 0 net=4704
rlabel metal2 149 -371 149 -371 0 net=6058
rlabel metal2 163 -371 163 -371 0 net=1629
rlabel metal2 296 -371 296 -371 0 net=1554
rlabel metal2 530 -371 530 -371 0 net=7542
rlabel metal2 891 -371 891 -371 0 net=8229
rlabel metal2 996 -371 996 -371 0 net=10061
rlabel metal2 1248 -371 1248 -371 0 net=11761
rlabel metal2 128 -373 128 -373 0 net=4038
rlabel metal2 310 -373 310 -373 0 net=1706
rlabel metal2 565 -373 565 -373 0 net=10922
rlabel metal2 1157 -373 1157 -373 0 net=10857
rlabel metal2 1255 -373 1255 -373 0 net=11821
rlabel metal2 152 -375 152 -375 0 net=1332
rlabel metal2 184 -375 184 -375 0 net=5169
rlabel metal2 380 -375 380 -375 0 net=3175
rlabel metal2 488 -375 488 -375 0 net=8464
rlabel metal2 1136 -375 1136 -375 0 net=10693
rlabel metal2 1262 -375 1262 -375 0 net=11861
rlabel metal2 163 -377 163 -377 0 net=5951
rlabel metal2 677 -377 677 -377 0 net=8134
rlabel metal2 1087 -377 1087 -377 0 net=11189
rlabel metal2 1276 -377 1276 -377 0 net=11965
rlabel metal2 170 -379 170 -379 0 net=11962
rlabel metal2 1290 -379 1290 -379 0 net=12119
rlabel metal2 170 -381 170 -381 0 net=1717
rlabel metal2 198 -381 198 -381 0 net=3425
rlabel metal2 513 -381 513 -381 0 net=5286
rlabel metal2 800 -381 800 -381 0 net=6737
rlabel metal2 831 -381 831 -381 0 net=9148
rlabel metal2 1024 -381 1024 -381 0 net=8989
rlabel metal2 1115 -381 1115 -381 0 net=10495
rlabel metal2 184 -383 184 -383 0 net=4355
rlabel metal2 240 -383 240 -383 0 net=2271
rlabel metal2 240 -383 240 -383 0 net=2271
rlabel metal2 247 -383 247 -383 0 net=3989
rlabel metal2 516 -383 516 -383 0 net=10625
rlabel metal2 191 -385 191 -385 0 net=5261
rlabel metal2 579 -385 579 -385 0 net=12140
rlabel metal2 198 -387 198 -387 0 net=3535
rlabel metal2 219 -387 219 -387 0 net=5003
rlabel metal2 534 -387 534 -387 0 net=4099
rlabel metal2 562 -387 562 -387 0 net=5513
rlabel metal2 604 -387 604 -387 0 net=492
rlabel metal2 726 -387 726 -387 0 net=10736
rlabel metal2 1150 -387 1150 -387 0 net=10783
rlabel metal2 124 -389 124 -389 0 net=7961
rlabel metal2 607 -389 607 -389 0 net=8627
rlabel metal2 1066 -389 1066 -389 0 net=9487
rlabel metal2 1164 -389 1164 -389 0 net=10919
rlabel metal2 135 -391 135 -391 0 net=2573
rlabel metal2 219 -391 219 -391 0 net=2935
rlabel metal2 684 -391 684 -391 0 net=10510
rlabel metal2 1122 -391 1122 -391 0 net=10931
rlabel metal2 1185 -391 1185 -391 0 net=11031
rlabel metal2 135 -393 135 -393 0 net=6063
rlabel metal2 754 -393 754 -393 0 net=11574
rlabel metal2 226 -395 226 -395 0 net=4235
rlabel metal2 457 -395 457 -395 0 net=3208
rlabel metal2 632 -395 632 -395 0 net=8467
rlabel metal2 800 -395 800 -395 0 net=6351
rlabel metal2 849 -395 849 -395 0 net=8791
rlabel metal2 1094 -395 1094 -395 0 net=10377
rlabel metal2 1192 -395 1192 -395 0 net=11079
rlabel metal2 296 -397 296 -397 0 net=5515
rlabel metal2 576 -397 576 -397 0 net=9975
rlabel metal2 1206 -397 1206 -397 0 net=11157
rlabel metal2 303 -399 303 -399 0 net=1947
rlabel metal2 373 -399 373 -399 0 net=2597
rlabel metal2 481 -399 481 -399 0 net=9045
rlabel metal2 1101 -399 1101 -399 0 net=10431
rlabel metal2 310 -401 310 -401 0 net=1693
rlabel metal2 716 -401 716 -401 0 net=6847
rlabel metal2 898 -401 898 -401 0 net=9347
rlabel metal2 324 -403 324 -403 0 net=1816
rlabel metal2 576 -403 576 -403 0 net=2576
rlabel metal2 828 -403 828 -403 0 net=7107
rlabel metal2 905 -403 905 -403 0 net=7703
rlabel metal2 107 -405 107 -405 0 net=3237
rlabel metal2 579 -405 579 -405 0 net=10571
rlabel metal2 107 -407 107 -407 0 net=2605
rlabel metal2 289 -407 289 -407 0 net=1987
rlabel metal2 331 -407 331 -407 0 net=5129
rlabel metal2 583 -407 583 -407 0 net=628
rlabel metal2 849 -407 849 -407 0 net=6777
rlabel metal2 1031 -407 1031 -407 0 net=10583
rlabel metal2 1052 -407 1052 -407 0 net=9243
rlabel metal2 1101 -407 1101 -407 0 net=11135
rlabel metal2 177 -409 177 -409 0 net=4531
rlabel metal2 583 -409 583 -409 0 net=4547
rlabel metal2 719 -409 719 -409 0 net=9809
rlabel metal2 968 -409 968 -409 0 net=8169
rlabel metal2 1010 -409 1010 -409 0 net=8657
rlabel metal2 1108 -409 1108 -409 0 net=10467
rlabel metal2 156 -411 156 -411 0 net=9265
rlabel metal2 131 -413 131 -413 0 net=1575
rlabel metal2 177 -413 177 -413 0 net=4739
rlabel metal2 586 -413 586 -413 0 net=7648
rlabel metal2 912 -413 912 -413 0 net=7753
rlabel metal2 233 -415 233 -415 0 net=5963
rlabel metal2 723 -415 723 -415 0 net=6033
rlabel metal2 926 -415 926 -415 0 net=8027
rlabel metal2 338 -417 338 -417 0 net=2491
rlabel metal2 520 -417 520 -417 0 net=6485
rlabel metal2 940 -417 940 -417 0 net=8071
rlabel metal2 345 -419 345 -419 0 net=3149
rlabel metal2 506 -419 506 -419 0 net=3919
rlabel metal2 597 -419 597 -419 0 net=9850
rlabel metal2 149 -421 149 -421 0 net=6271
rlabel metal2 373 -423 373 -423 0 net=3779
rlabel metal2 702 -423 702 -423 0 net=6695
rlabel metal2 835 -423 835 -423 0 net=7259
rlabel metal2 982 -423 982 -423 0 net=8285
rlabel metal2 380 -425 380 -425 0 net=3027
rlabel metal2 611 -425 611 -425 0 net=4921
rlabel metal2 632 -425 632 -425 0 net=7494
rlabel metal2 387 -427 387 -427 0 net=6947
rlabel metal2 635 -427 635 -427 0 net=12074
rlabel metal2 352 -429 352 -429 0 net=1959
rlabel metal2 394 -429 394 -429 0 net=4358
rlabel metal2 642 -429 642 -429 0 net=8197
rlabel metal2 72 -431 72 -431 0 net=3667
rlabel metal2 401 -431 401 -431 0 net=4843
rlabel metal2 72 -433 72 -433 0 net=1889
rlabel metal2 100 -433 100 -433 0 net=2774
rlabel metal2 401 -433 401 -433 0 net=3603
rlabel metal2 660 -433 660 -433 0 net=10341
rlabel metal2 86 -435 86 -435 0 net=4915
rlabel metal2 422 -435 422 -435 0 net=2953
rlabel metal2 499 -435 499 -435 0 net=4296
rlabel metal2 660 -435 660 -435 0 net=5563
rlabel metal2 684 -435 684 -435 0 net=9143
rlabel metal2 100 -437 100 -437 0 net=3217
rlabel metal2 415 -437 415 -437 0 net=2893
rlabel metal2 429 -437 429 -437 0 net=2993
rlabel metal2 555 -437 555 -437 0 net=9431
rlabel metal2 212 -439 212 -439 0 net=8650
rlabel metal2 254 -441 254 -441 0 net=5149
rlabel metal2 667 -441 667 -441 0 net=5537
rlabel metal2 730 -441 730 -441 0 net=6499
rlabel metal2 772 -441 772 -441 0 net=7641
rlabel metal2 947 -441 947 -441 0 net=9577
rlabel metal2 254 -443 254 -443 0 net=2199
rlabel metal2 534 -443 534 -443 0 net=7853
rlabel metal2 317 -445 317 -445 0 net=2653
rlabel metal2 667 -445 667 -445 0 net=6965
rlabel metal2 870 -445 870 -445 0 net=7561
rlabel metal2 933 -445 933 -445 0 net=8047
rlabel metal2 268 -447 268 -447 0 net=2317
rlabel metal2 355 -447 355 -447 0 net=4341
rlabel metal2 590 -447 590 -447 0 net=5039
rlabel metal2 877 -447 877 -447 0 net=7623
rlabel metal2 93 -449 93 -449 0 net=3372
rlabel metal2 590 -449 590 -449 0 net=5395
rlabel metal2 688 -449 688 -449 0 net=6563
rlabel metal2 887 -449 887 -449 0 net=5219
rlabel metal2 51 -451 51 -451 0 net=8138
rlabel metal2 702 -451 702 -451 0 net=6099
rlabel metal2 744 -451 744 -451 0 net=6107
rlabel metal2 789 -451 789 -451 0 net=7179
rlabel metal2 569 -453 569 -453 0 net=5929
rlabel metal2 674 -453 674 -453 0 net=5353
rlabel metal2 751 -453 751 -453 0 net=7431
rlabel metal2 142 -455 142 -455 0 net=1849
rlabel metal2 695 -455 695 -455 0 net=5971
rlabel metal2 758 -455 758 -455 0 net=11511
rlabel metal2 142 -457 142 -457 0 net=4871
rlabel metal2 695 -457 695 -457 0 net=9961
rlabel metal2 789 -459 789 -459 0 net=8497
rlabel metal2 807 -461 807 -461 0 net=8447
rlabel metal2 779 -463 779 -463 0 net=6635
rlabel metal2 821 -463 821 -463 0 net=7529
rlabel metal2 639 -465 639 -465 0 net=4165
rlabel metal2 639 -467 639 -467 0 net=9020
rlabel metal2 611 -469 611 -469 0 net=9457
rlabel metal2 646 -471 646 -471 0 net=6723
rlabel metal2 618 -473 618 -473 0 net=5743
rlabel metal2 450 -475 450 -475 0 net=4221
rlabel metal2 450 -477 450 -477 0 net=2457
rlabel metal2 58 -488 58 -488 0 net=5397
rlabel metal2 611 -488 611 -488 0 net=9044
rlabel metal2 1346 -488 1346 -488 0 net=11823
rlabel metal2 1346 -488 1346 -488 0 net=11823
rlabel metal2 1377 -488 1377 -488 0 net=11405
rlabel metal2 65 -490 65 -490 0 net=5681
rlabel metal2 310 -490 310 -490 0 net=1694
rlabel metal2 373 -490 373 -490 0 net=3780
rlabel metal2 625 -490 625 -490 0 net=4922
rlabel metal2 698 -490 698 -490 0 net=7798
rlabel metal2 51 -492 51 -492 0 net=2067
rlabel metal2 68 -492 68 -492 0 net=2574
rlabel metal2 212 -492 212 -492 0 net=2937
rlabel metal2 233 -492 233 -492 0 net=5964
rlabel metal2 768 -492 768 -492 0 net=11404
rlabel metal2 72 -494 72 -494 0 net=1890
rlabel metal2 114 -494 114 -494 0 net=1026
rlabel metal2 131 -494 131 -494 0 net=1869
rlabel metal2 338 -494 338 -494 0 net=2492
rlabel metal2 831 -494 831 -494 0 net=11080
rlabel metal2 1325 -494 1325 -494 0 net=11863
rlabel metal2 72 -496 72 -496 0 net=6377
rlabel metal2 124 -496 124 -496 0 net=6948
rlabel metal2 513 -496 513 -496 0 net=4844
rlabel metal2 978 -496 978 -496 0 net=11087
rlabel metal2 128 -498 128 -498 0 net=3991
rlabel metal2 254 -498 254 -498 0 net=2200
rlabel metal2 569 -498 569 -498 0 net=1850
rlabel metal2 849 -498 849 -498 0 net=6779
rlabel metal2 849 -498 849 -498 0 net=6779
rlabel metal2 863 -498 863 -498 0 net=6849
rlabel metal2 863 -498 863 -498 0 net=6849
rlabel metal2 884 -498 884 -498 0 net=12120
rlabel metal2 152 -500 152 -500 0 net=1718
rlabel metal2 177 -500 177 -500 0 net=4741
rlabel metal2 373 -500 373 -500 0 net=5201
rlabel metal2 782 -500 782 -500 0 net=7754
rlabel metal2 1206 -500 1206 -500 0 net=10573
rlabel metal2 1206 -500 1206 -500 0 net=10573
rlabel metal2 152 -502 152 -502 0 net=4356
rlabel metal2 198 -502 198 -502 0 net=3537
rlabel metal2 215 -502 215 -502 0 net=6486
rlabel metal2 933 -502 933 -502 0 net=7625
rlabel metal2 933 -502 933 -502 0 net=7625
rlabel metal2 954 -502 954 -502 0 net=9811
rlabel metal2 156 -504 156 -504 0 net=1576
rlabel metal2 586 -504 586 -504 0 net=6564
rlabel metal2 887 -504 887 -504 0 net=10511
rlabel metal2 163 -506 163 -506 0 net=5953
rlabel metal2 646 -506 646 -506 0 net=5744
rlabel metal2 688 -506 688 -506 0 net=7211
rlabel metal2 891 -506 891 -506 0 net=8231
rlabel metal2 163 -508 163 -508 0 net=2599
rlabel metal2 460 -508 460 -508 0 net=6724
rlabel metal2 870 -508 870 -508 0 net=5041
rlabel metal2 156 -510 156 -510 0 net=7017
rlabel metal2 912 -510 912 -510 0 net=7563
rlabel metal2 968 -510 968 -510 0 net=11513
rlabel metal2 177 -512 177 -512 0 net=4115
rlabel metal2 688 -512 688 -512 0 net=4167
rlabel metal2 786 -512 786 -512 0 net=10496
rlabel metal2 184 -514 184 -514 0 net=5931
rlabel metal2 705 -514 705 -514 0 net=7432
rlabel metal2 1045 -514 1045 -514 0 net=6273
rlabel metal2 219 -516 219 -516 0 net=3238
rlabel metal2 499 -516 499 -516 0 net=8028
rlabel metal2 1045 -516 1045 -516 0 net=7369
rlabel metal2 222 -518 222 -518 0 net=8139
rlabel metal2 982 -518 982 -518 0 net=8049
rlabel metal2 982 -518 982 -518 0 net=8049
rlabel metal2 989 -518 989 -518 0 net=8171
rlabel metal2 1087 -518 1087 -518 0 net=11191
rlabel metal2 240 -520 240 -520 0 net=2273
rlabel metal2 296 -520 296 -520 0 net=5517
rlabel metal2 653 -520 653 -520 0 net=5355
rlabel metal2 754 -520 754 -520 0 net=8628
rlabel metal2 1178 -520 1178 -520 0 net=10343
rlabel metal2 243 -522 243 -522 0 net=7547
rlabel metal2 614 -522 614 -522 0 net=9365
rlabel metal2 1178 -522 1178 -522 0 net=10695
rlabel metal2 268 -524 268 -524 0 net=5651
rlabel metal2 380 -524 380 -524 0 net=3029
rlabel metal2 513 -524 513 -524 0 net=6966
rlabel metal2 709 -524 709 -524 0 net=5539
rlabel metal2 709 -524 709 -524 0 net=5539
rlabel metal2 716 -524 716 -524 0 net=9348
rlabel metal2 268 -526 268 -526 0 net=5131
rlabel metal2 359 -526 359 -526 0 net=5170
rlabel metal2 719 -526 719 -526 0 net=7704
rlabel metal2 1248 -526 1248 -526 0 net=10859
rlabel metal2 107 -528 107 -528 0 net=2607
rlabel metal2 397 -528 397 -528 0 net=477
rlabel metal2 737 -528 737 -528 0 net=5973
rlabel metal2 751 -528 751 -528 0 net=6619
rlabel metal2 1241 -528 1241 -528 0 net=10785
rlabel metal2 107 -530 107 -530 0 net=9813
rlabel metal2 835 -530 835 -530 0 net=7181
rlabel metal2 901 -530 901 -530 0 net=8651
rlabel metal2 1150 -530 1150 -530 0 net=9977
rlabel metal2 159 -532 159 -532 0 net=10747
rlabel metal2 296 -534 296 -534 0 net=3605
rlabel metal2 408 -534 408 -534 0 net=2655
rlabel metal2 499 -534 499 -534 0 net=7579
rlabel metal2 926 -534 926 -534 0 net=9047
rlabel metal2 1164 -534 1164 -534 0 net=10063
rlabel metal2 317 -536 317 -536 0 net=2319
rlabel metal2 401 -536 401 -536 0 net=3797
rlabel metal2 733 -536 733 -536 0 net=6647
rlabel metal2 772 -536 772 -536 0 net=5220
rlabel metal2 1073 -536 1073 -536 0 net=8991
rlabel metal2 1171 -536 1171 -536 0 net=10379
rlabel metal2 303 -538 303 -538 0 net=1949
rlabel metal2 324 -538 324 -538 0 net=1989
rlabel metal2 366 -538 366 -538 0 net=5665
rlabel metal2 786 -538 786 -538 0 net=6353
rlabel metal2 814 -538 814 -538 0 net=6697
rlabel metal2 835 -538 835 -538 0 net=6739
rlabel metal2 856 -538 856 -538 0 net=8659
rlabel metal2 1073 -538 1073 -538 0 net=9267
rlabel metal2 1185 -538 1185 -538 0 net=10469
rlabel metal2 261 -540 261 -540 0 net=1631
rlabel metal2 324 -540 324 -540 0 net=1961
rlabel metal2 415 -540 415 -540 0 net=2995
rlabel metal2 502 -540 502 -540 0 net=8468
rlabel metal2 821 -540 821 -540 0 net=7531
rlabel metal2 919 -540 919 -540 0 net=8499
rlabel metal2 1108 -540 1108 -540 0 net=10433
rlabel metal2 387 -542 387 -542 0 net=3369
rlabel metal2 502 -542 502 -542 0 net=11032
rlabel metal2 443 -544 443 -544 0 net=4223
rlabel metal2 674 -544 674 -544 0 net=9089
rlabel metal2 1101 -544 1101 -544 0 net=11137
rlabel metal2 1276 -544 1276 -544 0 net=11291
rlabel metal2 450 -546 450 -546 0 net=2459
rlabel metal2 492 -546 492 -546 0 net=5005
rlabel metal2 660 -546 660 -546 0 net=5565
rlabel metal2 730 -546 730 -546 0 net=6501
rlabel metal2 807 -546 807 -546 0 net=6637
rlabel metal2 919 -546 919 -546 0 net=8073
rlabel metal2 1003 -546 1003 -546 0 net=8287
rlabel metal2 1094 -546 1094 -546 0 net=9245
rlabel metal2 1115 -546 1115 -546 0 net=9433
rlabel metal2 1304 -546 1304 -546 0 net=11375
rlabel metal2 121 -548 121 -548 0 net=9723
rlabel metal2 1311 -548 1311 -548 0 net=11763
rlabel metal2 121 -550 121 -550 0 net=5445
rlabel metal2 534 -550 534 -550 0 net=5514
rlabel metal2 590 -550 590 -550 0 net=2103
rlabel metal2 604 -550 604 -550 0 net=7963
rlabel metal2 975 -550 975 -550 0 net=9531
rlabel metal2 1094 -550 1094 -550 0 net=9459
rlabel metal2 1332 -550 1332 -550 0 net=11635
rlabel metal2 93 -552 93 -552 0 net=11927
rlabel metal2 142 -554 142 -554 0 net=4873
rlabel metal2 635 -554 635 -554 0 net=9919
rlabel metal2 135 -556 135 -556 0 net=6065
rlabel metal2 394 -556 394 -556 0 net=3669
rlabel metal2 537 -556 537 -556 0 net=7108
rlabel metal2 940 -556 940 -556 0 net=7643
rlabel metal2 135 -558 135 -558 0 net=10920
rlabel metal2 149 -560 149 -560 0 net=7679
rlabel metal2 149 -562 149 -562 0 net=1344
rlabel metal2 779 -562 779 -562 0 net=10799
rlabel metal2 191 -564 191 -564 0 net=5262
rlabel metal2 429 -564 429 -564 0 net=5151
rlabel metal2 639 -564 639 -564 0 net=5263
rlabel metal2 793 -564 793 -564 0 net=9144
rlabel metal2 191 -566 191 -566 0 net=3427
rlabel metal2 492 -566 492 -566 0 net=4549
rlabel metal2 660 -566 660 -566 0 net=5895
rlabel metal2 1269 -566 1269 -566 0 net=11159
rlabel metal2 345 -568 345 -568 0 net=3151
rlabel metal2 436 -568 436 -568 0 net=2955
rlabel metal2 471 -568 471 -568 0 net=4343
rlabel metal2 583 -568 583 -568 0 net=5367
rlabel metal2 1290 -568 1290 -568 0 net=11967
rlabel metal2 198 -570 198 -570 0 net=12141
rlabel metal2 250 -572 250 -572 0 net=4683
rlabel metal2 352 -572 352 -572 0 net=2219
rlabel metal2 422 -574 422 -574 0 net=2895
rlabel metal2 464 -574 464 -574 0 net=3177
rlabel metal2 485 -574 485 -574 0 net=6101
rlabel metal2 100 -576 100 -576 0 net=3219
rlabel metal2 478 -576 478 -576 0 net=2281
rlabel metal2 86 -578 86 -578 0 net=4917
rlabel metal2 422 -578 422 -578 0 net=3921
rlabel metal2 527 -578 527 -578 0 net=4533
rlabel metal2 79 -580 79 -580 0 net=1533
rlabel metal2 520 -580 520 -580 0 net=6035
rlabel metal2 527 -582 527 -582 0 net=6545
rlabel metal2 548 -584 548 -584 0 net=4475
rlabel metal2 723 -584 723 -584 0 net=7261
rlabel metal2 226 -586 226 -586 0 net=4237
rlabel metal2 555 -586 555 -586 0 net=996
rlabel metal2 905 -586 905 -586 0 net=7855
rlabel metal2 40 -588 40 -588 0 net=2235
rlabel metal2 541 -588 541 -588 0 net=4101
rlabel metal2 947 -588 947 -588 0 net=8199
rlabel metal2 40 -590 40 -590 0 net=5359
rlabel metal2 541 -590 541 -590 0 net=8448
rlabel metal2 1010 -592 1010 -592 0 net=10933
rlabel metal2 1220 -592 1220 -592 0 net=10627
rlabel metal2 807 -594 807 -594 0 net=10655
rlabel metal2 961 -596 961 -596 0 net=9579
rlabel metal2 961 -598 961 -598 0 net=8793
rlabel metal2 1066 -600 1066 -600 0 net=9489
rlabel metal2 1136 -602 1136 -602 0 net=9963
rlabel metal2 1038 -604 1038 -604 0 net=10585
rlabel metal2 758 -606 758 -606 0 net=8825
rlabel metal2 758 -608 758 -608 0 net=6109
rlabel metal2 765 -610 765 -610 0 net=8643
rlabel metal2 44 -621 44 -621 0 net=11307
rlabel metal2 387 -621 387 -621 0 net=3370
rlabel metal2 649 -621 649 -621 0 net=9724
rlabel metal2 1185 -621 1185 -621 0 net=10471
rlabel metal2 1472 -621 1472 -621 0 net=6275
rlabel metal2 51 -623 51 -623 0 net=2068
rlabel metal2 527 -623 527 -623 0 net=7564
rlabel metal2 975 -623 975 -623 0 net=7371
rlabel metal2 1059 -623 1059 -623 0 net=9367
rlabel metal2 1234 -623 1234 -623 0 net=6621
rlabel metal2 51 -625 51 -625 0 net=5653
rlabel metal2 397 -625 397 -625 0 net=92
rlabel metal2 684 -625 684 -625 0 net=10860
rlabel metal2 1311 -625 1311 -625 0 net=11765
rlabel metal2 72 -627 72 -627 0 net=6378
rlabel metal2 107 -627 107 -627 0 net=9814
rlabel metal2 698 -627 698 -627 0 net=7532
rlabel metal2 887 -627 887 -627 0 net=9246
rlabel metal2 1136 -627 1136 -627 0 net=9965
rlabel metal2 1353 -627 1353 -627 0 net=11406
rlabel metal2 1388 -627 1388 -627 0 net=10513
rlabel metal2 65 -629 65 -629 0 net=8403
rlabel metal2 1157 -629 1157 -629 0 net=10587
rlabel metal2 1332 -629 1332 -629 0 net=11929
rlabel metal2 65 -631 65 -631 0 net=2237
rlabel metal2 233 -631 233 -631 0 net=6901
rlabel metal2 537 -631 537 -631 0 net=7262
rlabel metal2 730 -631 730 -631 0 net=10344
rlabel metal2 1227 -631 1227 -631 0 net=10657
rlabel metal2 1276 -631 1276 -631 0 net=11293
rlabel metal2 1356 -631 1356 -631 0 net=5042
rlabel metal2 72 -633 72 -633 0 net=5203
rlabel metal2 429 -633 429 -633 0 net=3152
rlabel metal2 541 -633 541 -633 0 net=5954
rlabel metal2 702 -633 702 -633 0 net=8232
rlabel metal2 82 -635 82 -635 0 net=4918
rlabel metal2 114 -635 114 -635 0 net=3003
rlabel metal2 128 -635 128 -635 0 net=3993
rlabel metal2 243 -635 243 -635 0 net=2195
rlabel metal2 432 -635 432 -635 0 net=6648
rlabel metal2 772 -635 772 -635 0 net=11636
rlabel metal2 1360 -635 1360 -635 0 net=12143
rlabel metal2 86 -637 86 -637 0 net=1535
rlabel metal2 128 -637 128 -637 0 net=4103
rlabel metal2 702 -637 702 -637 0 net=6111
rlabel metal2 768 -637 768 -637 0 net=10865
rlabel metal2 86 -639 86 -639 0 net=5567
rlabel metal2 705 -639 705 -639 0 net=6515
rlabel metal2 898 -639 898 -639 0 net=10934
rlabel metal2 1017 -639 1017 -639 0 net=8501
rlabel metal2 1129 -639 1129 -639 0 net=9921
rlabel metal2 1269 -639 1269 -639 0 net=11161
rlabel metal2 138 -641 138 -641 0 net=970
rlabel metal2 247 -641 247 -641 0 net=8660
rlabel metal2 863 -641 863 -641 0 net=6851
rlabel metal2 940 -641 940 -641 0 net=7681
rlabel metal2 1080 -641 1080 -641 0 net=8993
rlabel metal2 1157 -641 1157 -641 0 net=10065
rlabel metal2 1171 -641 1171 -641 0 net=10381
rlabel metal2 1290 -641 1290 -641 0 net=11969
rlabel metal2 107 -643 107 -643 0 net=8021
rlabel metal2 250 -643 250 -643 0 net=3741
rlabel metal2 555 -643 555 -643 0 net=28
rlabel metal2 772 -643 772 -643 0 net=5751
rlabel metal2 954 -643 954 -643 0 net=7965
rlabel metal2 1052 -643 1052 -643 0 net=9091
rlabel metal2 1192 -643 1192 -643 0 net=11139
rlabel metal2 142 -645 142 -645 0 net=6066
rlabel metal2 159 -645 159 -645 0 net=11443
rlabel metal2 149 -647 149 -647 0 net=2711
rlabel metal2 250 -647 250 -647 0 net=2282
rlabel metal2 485 -647 485 -647 0 net=6102
rlabel metal2 674 -647 674 -647 0 net=6639
rlabel metal2 831 -647 831 -647 0 net=10696
rlabel metal2 1206 -647 1206 -647 0 net=10575
rlabel metal2 1290 -647 1290 -647 0 net=11377
rlabel metal2 1325 -647 1325 -647 0 net=11865
rlabel metal2 152 -649 152 -649 0 net=9434
rlabel metal2 1241 -649 1241 -649 0 net=10749
rlabel metal2 156 -651 156 -651 0 net=2125
rlabel metal2 807 -651 807 -651 0 net=11824
rlabel metal2 163 -653 163 -653 0 net=2600
rlabel metal2 443 -653 443 -653 0 net=4225
rlabel metal2 586 -653 586 -653 0 net=9279
rlabel metal2 1248 -653 1248 -653 0 net=10787
rlabel metal2 163 -655 163 -655 0 net=2049
rlabel metal2 695 -655 695 -655 0 net=8675
rlabel metal2 1248 -655 1248 -655 0 net=10181
rlabel metal2 58 -657 58 -657 0 net=5399
rlabel metal2 709 -657 709 -657 0 net=5541
rlabel metal2 775 -657 775 -657 0 net=316
rlabel metal2 982 -657 982 -657 0 net=8051
rlabel metal2 1122 -657 1122 -657 0 net=9581
rlabel metal2 58 -659 58 -659 0 net=8529
rlabel metal2 170 -659 170 -659 0 net=2321
rlabel metal2 415 -659 415 -659 0 net=2997
rlabel metal2 450 -659 450 -659 0 net=2957
rlabel metal2 450 -659 450 -659 0 net=2957
rlabel metal2 457 -659 457 -659 0 net=2461
rlabel metal2 457 -659 457 -659 0 net=2461
rlabel metal2 471 -659 471 -659 0 net=3179
rlabel metal2 565 -659 565 -659 0 net=9535
rlabel metal2 187 -661 187 -661 0 net=3538
rlabel metal2 219 -661 219 -661 0 net=1963
rlabel metal2 345 -661 345 -661 0 net=4685
rlabel metal2 716 -661 716 -661 0 net=11035
rlabel metal2 124 -663 124 -663 0 net=4129
rlabel metal2 373 -663 373 -663 0 net=3221
rlabel metal2 471 -663 471 -663 0 net=2105
rlabel metal2 607 -663 607 -663 0 net=10083
rlabel metal2 149 -665 149 -665 0 net=3569
rlabel metal2 716 -665 716 -665 0 net=6699
rlabel metal2 856 -665 856 -665 0 net=11853
rlabel metal2 198 -667 198 -667 0 net=5221
rlabel metal2 198 -667 198 -667 0 net=5221
rlabel metal2 201 -667 201 -667 0 net=2938
rlabel metal2 268 -667 268 -667 0 net=5133
rlabel metal2 380 -667 380 -667 0 net=4551
rlabel metal2 719 -667 719 -667 0 net=9460
rlabel metal2 205 -669 205 -669 0 net=5369
rlabel metal2 723 -669 723 -669 0 net=11192
rlabel metal2 212 -671 212 -671 0 net=2221
rlabel metal2 401 -671 401 -671 0 net=3799
rlabel metal2 464 -671 464 -671 0 net=3731
rlabel metal2 726 -671 726 -671 0 net=7827
rlabel metal2 1024 -671 1024 -671 0 net=8645
rlabel metal2 268 -673 268 -673 0 net=3127
rlabel metal2 733 -673 733 -673 0 net=7203
rlabel metal2 961 -673 961 -673 0 net=8795
rlabel metal2 275 -675 275 -675 0 net=5683
rlabel metal2 779 -675 779 -675 0 net=7644
rlabel metal2 1003 -675 1003 -675 0 net=8289
rlabel metal2 254 -677 254 -677 0 net=1907
rlabel metal2 282 -677 282 -677 0 net=1870
rlabel metal2 611 -677 611 -677 0 net=7549
rlabel metal2 1006 -677 1006 -677 0 net=9812
rlabel metal2 282 -679 282 -679 0 net=1929
rlabel metal2 737 -679 737 -679 0 net=5975
rlabel metal2 786 -679 786 -679 0 net=6355
rlabel metal2 877 -679 877 -679 0 net=7183
rlabel metal2 968 -679 968 -679 0 net=8141
rlabel metal2 121 -681 121 -681 0 net=5447
rlabel metal2 744 -681 744 -681 0 net=5667
rlabel metal2 793 -681 793 -681 0 net=11841
rlabel metal2 121 -683 121 -683 0 net=9268
rlabel metal2 296 -685 296 -685 0 net=3607
rlabel metal2 646 -685 646 -685 0 net=5519
rlabel metal2 793 -685 793 -685 0 net=11514
rlabel metal2 289 -687 289 -687 0 net=2275
rlabel metal2 310 -687 310 -687 0 net=7581
rlabel metal2 905 -687 905 -687 0 net=7857
rlabel metal2 1031 -687 1031 -687 0 net=8653
rlabel metal2 1262 -687 1262 -687 0 net=10801
rlabel metal2 317 -689 317 -689 0 net=1951
rlabel metal2 352 -689 352 -689 0 net=5153
rlabel metal2 618 -689 618 -689 0 net=5006
rlabel metal2 733 -689 733 -689 0 net=8113
rlabel metal2 1108 -689 1108 -689 0 net=10435
rlabel metal2 317 -691 317 -691 0 net=3923
rlabel metal2 513 -691 513 -691 0 net=5477
rlabel metal2 800 -691 800 -691 0 net=6503
rlabel metal2 884 -691 884 -691 0 net=7213
rlabel metal2 989 -691 989 -691 0 net=8173
rlabel metal2 401 -693 401 -693 0 net=3017
rlabel metal2 660 -693 660 -693 0 net=5897
rlabel metal2 807 -693 807 -693 0 net=5825
rlabel metal2 933 -693 933 -693 0 net=7627
rlabel metal2 992 -693 992 -693 0 net=9978
rlabel metal2 408 -695 408 -695 0 net=2657
rlabel metal2 513 -695 513 -695 0 net=3671
rlabel metal2 576 -695 576 -695 0 net=4535
rlabel metal2 660 -695 660 -695 0 net=4169
rlabel metal2 814 -695 814 -695 0 net=6547
rlabel metal2 905 -695 905 -695 0 net=11088
rlabel metal2 68 -697 68 -697 0 net=5279
rlabel metal2 821 -697 821 -697 0 net=6741
rlabel metal2 884 -697 884 -697 0 net=9048
rlabel metal2 1031 -697 1031 -697 0 net=7889
rlabel metal2 1062 -697 1062 -697 0 net=10677
rlabel metal2 96 -699 96 -699 0 net=8809
rlabel metal2 828 -699 828 -699 0 net=7415
rlabel metal2 1038 -699 1038 -699 0 net=8827
rlabel metal2 1220 -699 1220 -699 0 net=10629
rlabel metal2 135 -701 135 -701 0 net=7901
rlabel metal2 1066 -701 1066 -701 0 net=9491
rlabel metal2 135 -703 135 -703 0 net=5361
rlabel metal2 359 -703 359 -703 0 net=2609
rlabel metal2 422 -703 422 -703 0 net=2897
rlabel metal2 520 -703 520 -703 0 net=6037
rlabel metal2 667 -703 667 -703 0 net=6791
rlabel metal2 1087 -703 1087 -703 0 net=9533
rlabel metal2 184 -705 184 -705 0 net=5933
rlabel metal2 359 -705 359 -705 0 net=5357
rlabel metal2 667 -705 667 -705 0 net=6079
rlabel metal2 870 -705 870 -705 0 net=7019
rlabel metal2 947 -705 947 -705 0 net=8201
rlabel metal2 436 -707 436 -707 0 net=6441
rlabel metal2 520 -709 520 -709 0 net=4875
rlabel metal2 653 -709 653 -709 0 net=5213
rlabel metal2 835 -709 835 -709 0 net=5195
rlabel metal2 919 -709 919 -709 0 net=8075
rlabel metal2 534 -711 534 -711 0 net=4476
rlabel metal2 849 -711 849 -711 0 net=6781
rlabel metal2 548 -713 548 -713 0 net=4239
rlabel metal2 709 -713 709 -713 0 net=6135
rlabel metal2 919 -713 919 -713 0 net=8855
rlabel metal2 548 -715 548 -715 0 net=5265
rlabel metal2 394 -717 394 -717 0 net=4745
rlabel metal2 177 -719 177 -719 0 net=4117
rlabel metal2 562 -719 562 -719 0 net=4345
rlabel metal2 177 -721 177 -721 0 net=3031
rlabel metal2 191 -723 191 -723 0 net=3429
rlabel metal2 191 -725 191 -725 0 net=4743
rlabel metal2 303 -727 303 -727 0 net=1632
rlabel metal2 303 -729 303 -729 0 net=1547
rlabel metal2 331 -731 331 -731 0 net=1991
rlabel metal2 184 -733 184 -733 0 net=4393
rlabel metal2 37 -744 37 -744 0 net=8531
rlabel metal2 79 -744 79 -744 0 net=633
rlabel metal2 922 -744 922 -744 0 net=11444
rlabel metal2 1416 -744 1416 -744 0 net=11842
rlabel metal2 1633 -744 1633 -744 0 net=6277
rlabel metal2 44 -746 44 -746 0 net=11309
rlabel metal2 1570 -746 1570 -746 0 net=10515
rlabel metal2 44 -748 44 -748 0 net=2959
rlabel metal2 467 -748 467 -748 0 net=10861
rlabel metal2 1500 -748 1500 -748 0 net=6623
rlabel metal2 58 -750 58 -750 0 net=3571
rlabel metal2 166 -750 166 -750 0 net=11225
rlabel metal2 1521 -750 1521 -750 0 net=12145
rlabel metal2 1605 -750 1605 -750 0 net=6001
rlabel metal2 82 -752 82 -752 0 net=4643
rlabel metal2 607 -752 607 -752 0 net=6504
rlabel metal2 884 -752 884 -752 0 net=11997
rlabel metal2 93 -754 93 -754 0 net=5898
rlabel metal2 807 -754 807 -754 0 net=5827
rlabel metal2 807 -754 807 -754 0 net=5827
rlabel metal2 821 -754 821 -754 0 net=6743
rlabel metal2 905 -754 905 -754 0 net=10788
rlabel metal2 1353 -754 1353 -754 0 net=11295
rlabel metal2 93 -756 93 -756 0 net=3743
rlabel metal2 537 -756 537 -756 0 net=691
rlabel metal2 730 -756 730 -756 0 net=5668
rlabel metal2 782 -756 782 -756 0 net=9534
rlabel metal2 1241 -756 1241 -756 0 net=10085
rlabel metal2 1430 -756 1430 -756 0 net=8857
rlabel metal2 33 -758 33 -758 0 net=4849
rlabel metal2 558 -758 558 -758 0 net=11877
rlabel metal2 103 -760 103 -760 0 net=5134
rlabel metal2 485 -760 485 -760 0 net=2903
rlabel metal2 565 -760 565 -760 0 net=8174
rlabel metal2 1122 -760 1122 -760 0 net=8647
rlabel metal2 124 -762 124 -762 0 net=11417
rlabel metal2 128 -764 128 -764 0 net=4105
rlabel metal2 138 -764 138 -764 0 net=10866
rlabel metal2 1367 -764 1367 -764 0 net=11855
rlabel metal2 128 -766 128 -766 0 net=4537
rlabel metal2 632 -766 632 -766 0 net=4747
rlabel metal2 649 -766 649 -766 0 net=10189
rlabel metal2 1374 -766 1374 -766 0 net=11867
rlabel metal2 142 -768 142 -768 0 net=5191
rlabel metal2 730 -768 730 -768 0 net=5543
rlabel metal2 765 -768 765 -768 0 net=5977
rlabel metal2 828 -768 828 -768 0 net=7184
rlabel metal2 1003 -768 1003 -768 0 net=484
rlabel metal2 149 -770 149 -770 0 net=4687
rlabel metal2 628 -770 628 -770 0 net=10307
rlabel metal2 1388 -770 1388 -770 0 net=11971
rlabel metal2 184 -772 184 -772 0 net=11835
rlabel metal2 184 -774 184 -774 0 net=5223
rlabel metal2 205 -774 205 -774 0 net=5371
rlabel metal2 488 -774 488 -774 0 net=811
rlabel metal2 576 -774 576 -774 0 net=6700
rlabel metal2 733 -774 733 -774 0 net=883
rlabel metal2 187 -776 187 -776 0 net=8290
rlabel metal2 1227 -776 1227 -776 0 net=9923
rlabel metal2 191 -778 191 -778 0 net=4744
rlabel metal2 240 -778 240 -778 0 net=2713
rlabel metal2 471 -778 471 -778 0 net=2107
rlabel metal2 576 -778 576 -778 0 net=6356
rlabel metal2 870 -778 870 -778 0 net=11777
rlabel metal2 191 -780 191 -780 0 net=6439
rlabel metal2 471 -780 471 -780 0 net=3181
rlabel metal2 499 -780 499 -780 0 net=4347
rlabel metal2 625 -780 625 -780 0 net=6112
rlabel metal2 709 -780 709 -780 0 net=10382
rlabel metal2 1283 -780 1283 -780 0 net=10631
rlabel metal2 198 -782 198 -782 0 net=4077
rlabel metal2 579 -782 579 -782 0 net=7550
rlabel metal2 1038 -782 1038 -782 0 net=7903
rlabel metal2 1136 -782 1136 -782 0 net=8995
rlabel metal2 1269 -782 1269 -782 0 net=10577
rlabel metal2 205 -784 205 -784 0 net=2253
rlabel metal2 247 -784 247 -784 0 net=9280
rlabel metal2 1206 -784 1206 -784 0 net=9583
rlabel metal2 1381 -784 1381 -784 0 net=11931
rlabel metal2 233 -786 233 -786 0 net=6903
rlabel metal2 1080 -786 1080 -786 0 net=8143
rlabel metal2 1157 -786 1157 -786 0 net=10067
rlabel metal2 23 -788 23 -788 0 net=5497
rlabel metal2 250 -788 250 -788 0 net=11469
rlabel metal2 79 -790 79 -790 0 net=3539
rlabel metal2 275 -790 275 -790 0 net=4552
rlabel metal2 429 -790 429 -790 0 net=2659
rlabel metal2 534 -790 534 -790 0 net=7875
rlabel metal2 1171 -790 1171 -790 0 net=8829
rlabel metal2 135 -792 135 -792 0 net=5363
rlabel metal2 583 -792 583 -792 0 net=4227
rlabel metal2 642 -792 642 -792 0 net=8803
rlabel metal2 1248 -792 1248 -792 0 net=10183
rlabel metal2 1290 -792 1290 -792 0 net=11379
rlabel metal2 65 -794 65 -794 0 net=2238
rlabel metal2 590 -794 590 -794 0 net=10143
rlabel metal2 65 -796 65 -796 0 net=4039
rlabel metal2 842 -796 842 -796 0 net=6517
rlabel metal2 877 -796 877 -796 0 net=8797
rlabel metal2 1262 -796 1262 -796 0 net=10437
rlabel metal2 170 -798 170 -798 0 net=2323
rlabel metal2 408 -798 408 -798 0 net=2611
rlabel metal2 569 -798 569 -798 0 net=4241
rlabel metal2 593 -798 593 -798 0 net=8233
rlabel metal2 1185 -798 1185 -798 0 net=9369
rlabel metal2 1304 -798 1304 -798 0 net=10751
rlabel metal2 275 -800 275 -800 0 net=1577
rlabel metal2 814 -800 814 -800 0 net=8811
rlabel metal2 1318 -800 1318 -800 0 net=10803
rlabel metal2 289 -802 289 -802 0 net=5154
rlabel metal2 359 -802 359 -802 0 net=5358
rlabel metal2 908 -802 908 -802 0 net=9469
rlabel metal2 1325 -802 1325 -802 0 net=11037
rlabel metal2 163 -804 163 -804 0 net=2051
rlabel metal2 303 -804 303 -804 0 net=1549
rlabel metal2 303 -804 303 -804 0 net=1549
rlabel metal2 310 -804 310 -804 0 net=7582
rlabel metal2 765 -804 765 -804 0 net=5197
rlabel metal2 842 -804 842 -804 0 net=6137
rlabel metal2 856 -804 856 -804 0 net=9377
rlabel metal2 1332 -804 1332 -804 0 net=11141
rlabel metal2 261 -806 261 -806 0 net=5935
rlabel metal2 1339 -806 1339 -806 0 net=11163
rlabel metal2 261 -808 261 -808 0 net=1931
rlabel metal2 310 -808 310 -808 0 net=2197
rlabel metal2 408 -808 408 -808 0 net=2463
rlabel metal2 541 -808 541 -808 0 net=3609
rlabel metal2 586 -808 586 -808 0 net=9925
rlabel metal2 268 -810 268 -810 0 net=3129
rlabel metal2 387 -810 387 -810 0 net=2899
rlabel metal2 432 -810 432 -810 0 net=6399
rlabel metal2 859 -810 859 -810 0 net=11766
rlabel metal2 177 -812 177 -812 0 net=3033
rlabel metal2 457 -812 457 -812 0 net=4941
rlabel metal2 646 -812 646 -812 0 net=7271
rlabel metal2 716 -812 716 -812 0 net=5187
rlabel metal2 912 -812 912 -812 0 net=10472
rlabel metal2 177 -814 177 -814 0 net=2223
rlabel metal2 254 -814 254 -814 0 net=1909
rlabel metal2 282 -814 282 -814 0 net=4441
rlabel metal2 513 -814 513 -814 0 net=3673
rlabel metal2 565 -814 565 -814 0 net=8759
rlabel metal2 1192 -814 1192 -814 0 net=9537
rlabel metal2 1297 -814 1297 -814 0 net=10679
rlabel metal2 110 -816 110 -816 0 net=9715
rlabel metal2 156 -818 156 -818 0 net=2127
rlabel metal2 317 -818 317 -818 0 net=3924
rlabel metal2 653 -818 653 -818 0 net=8781
rlabel metal2 1255 -818 1255 -818 0 net=10659
rlabel metal2 156 -820 156 -820 0 net=3925
rlabel metal2 338 -820 338 -820 0 net=1993
rlabel metal2 338 -820 338 -820 0 net=1993
rlabel metal2 345 -820 345 -820 0 net=4131
rlabel metal2 656 -820 656 -820 0 net=8796
rlabel metal2 1234 -820 1234 -820 0 net=9967
rlabel metal2 135 -822 135 -822 0 net=9307
rlabel metal2 212 -824 212 -824 0 net=1965
rlabel metal2 226 -824 226 -824 0 net=3995
rlabel metal2 660 -824 660 -824 0 net=4170
rlabel metal2 887 -824 887 -824 0 net=8711
rlabel metal2 121 -826 121 -826 0 net=7283
rlabel metal2 345 -826 345 -826 0 net=5267
rlabel metal2 667 -826 667 -826 0 net=6081
rlabel metal2 912 -826 912 -826 0 net=9093
rlabel metal2 114 -828 114 -828 0 net=3005
rlabel metal2 667 -828 667 -828 0 net=5155
rlabel metal2 695 -828 695 -828 0 net=5400
rlabel metal2 740 -828 740 -828 0 net=9713
rlabel metal2 51 -830 51 -830 0 net=5655
rlabel metal2 751 -830 751 -830 0 net=5685
rlabel metal2 919 -830 919 -830 0 net=6443
rlabel metal2 100 -832 100 -832 0 net=1537
rlabel metal2 170 -832 170 -832 0 net=2709
rlabel metal2 681 -832 681 -832 0 net=5215
rlabel metal2 772 -832 772 -832 0 net=5753
rlabel metal2 929 -832 929 -832 0 net=10588
rlabel metal2 51 -834 51 -834 0 net=9815
rlabel metal2 100 -836 100 -836 0 net=9311
rlabel metal2 352 -838 352 -838 0 net=3733
rlabel metal2 681 -838 681 -838 0 net=5449
rlabel metal2 744 -838 744 -838 0 net=5479
rlabel metal2 786 -838 786 -838 0 net=5521
rlabel metal2 947 -838 947 -838 0 net=6783
rlabel metal2 947 -838 947 -838 0 net=6783
rlabel metal2 954 -838 954 -838 0 net=7205
rlabel metal2 1006 -838 1006 -838 0 net=9789
rlabel metal2 72 -840 72 -840 0 net=5205
rlabel metal2 786 -840 786 -840 0 net=11515
rlabel metal2 72 -842 72 -842 0 net=4395
rlabel metal2 415 -842 415 -842 0 net=3801
rlabel metal2 688 -842 688 -842 0 net=5281
rlabel metal2 933 -842 933 -842 0 net=6793
rlabel metal2 982 -842 982 -842 0 net=7629
rlabel metal2 1052 -842 1052 -842 0 net=8053
rlabel metal2 296 -844 296 -844 0 net=2277
rlabel metal2 401 -844 401 -844 0 net=3019
rlabel metal2 688 -844 688 -844 0 net=2559
rlabel metal2 831 -844 831 -844 0 net=7791
rlabel metal2 1066 -844 1066 -844 0 net=8077
rlabel metal2 324 -846 324 -846 0 net=1952
rlabel metal2 831 -846 831 -846 0 net=10743
rlabel metal2 324 -848 324 -848 0 net=4877
rlabel metal2 891 -848 891 -848 0 net=6549
rlabel metal2 1017 -848 1017 -848 0 net=7829
rlabel metal2 1101 -848 1101 -848 0 net=8405
rlabel metal2 401 -850 401 -850 0 net=2999
rlabel metal2 506 -850 506 -850 0 net=3431
rlabel metal2 611 -850 611 -850 0 net=6039
rlabel metal2 926 -850 926 -850 0 net=7021
rlabel metal2 989 -850 989 -850 0 net=7935
rlabel metal2 1108 -850 1108 -850 0 net=9493
rlabel metal2 86 -852 86 -852 0 net=5569
rlabel metal2 611 -852 611 -852 0 net=8654
rlabel metal2 107 -854 107 -854 0 net=8023
rlabel metal2 107 -856 107 -856 0 net=9641
rlabel metal2 989 -856 989 -856 0 net=7029
rlabel metal2 1017 -856 1017 -856 0 net=7301
rlabel metal2 1115 -856 1115 -856 0 net=8503
rlabel metal2 373 -858 373 -858 0 net=3223
rlabel metal2 1045 -858 1045 -858 0 net=7967
rlabel metal2 1129 -858 1129 -858 0 net=8677
rlabel metal2 373 -860 373 -860 0 net=4119
rlabel metal2 1010 -860 1010 -860 0 net=7683
rlabel metal2 1073 -860 1073 -860 0 net=8115
rlabel metal2 229 -862 229 -862 0 net=2287
rlabel metal2 968 -862 968 -862 0 net=7215
rlabel metal2 1024 -862 1024 -862 0 net=7859
rlabel metal2 1087 -862 1087 -862 0 net=8203
rlabel metal2 478 -864 478 -864 0 net=7341
rlabel metal2 1031 -864 1031 -864 0 net=7891
rlabel metal2 940 -866 940 -866 0 net=7417
rlabel metal2 975 -866 975 -866 0 net=7373
rlabel metal2 674 -868 674 -868 0 net=6641
rlabel metal2 674 -870 674 -870 0 net=4681
rlabel metal2 898 -870 898 -870 0 net=6853
rlabel metal2 898 -872 898 -872 0 net=5693
rlabel metal2 30 -883 30 -883 0 net=4397
rlabel metal2 89 -883 89 -883 0 net=1538
rlabel metal2 135 -883 135 -883 0 net=4442
rlabel metal2 292 -883 292 -883 0 net=1994
rlabel metal2 450 -883 450 -883 0 net=5372
rlabel metal2 618 -883 618 -883 0 net=4132
rlabel metal2 740 -883 740 -883 0 net=10752
rlabel metal2 1521 -883 1521 -883 0 net=11999
rlabel metal2 1696 -883 1696 -883 0 net=6279
rlabel metal2 65 -885 65 -885 0 net=4041
rlabel metal2 663 -885 663 -885 0 net=11856
rlabel metal2 1591 -885 1591 -885 0 net=12146
rlabel metal2 1619 -885 1619 -885 0 net=6625
rlabel metal2 65 -887 65 -887 0 net=3001
rlabel metal2 422 -887 422 -887 0 net=3035
rlabel metal2 457 -887 457 -887 0 net=4942
rlabel metal2 957 -887 957 -887 0 net=11164
rlabel metal2 1598 -887 1598 -887 0 net=10517
rlabel metal2 1633 -887 1633 -887 0 net=8859
rlabel metal2 72 -889 72 -889 0 net=4243
rlabel metal2 597 -889 597 -889 0 net=4228
rlabel metal2 635 -889 635 -889 0 net=11296
rlabel metal2 86 -891 86 -891 0 net=11221
rlabel metal2 103 -893 103 -893 0 net=5192
rlabel metal2 149 -893 149 -893 0 net=4689
rlabel metal2 761 -893 761 -893 0 net=6040
rlabel metal2 905 -893 905 -893 0 net=11142
rlabel metal2 107 -895 107 -895 0 net=3006
rlabel metal2 135 -895 135 -895 0 net=2901
rlabel metal2 422 -895 422 -895 0 net=5291
rlabel metal2 761 -895 761 -895 0 net=5669
rlabel metal2 898 -895 898 -895 0 net=5695
rlabel metal2 908 -895 908 -895 0 net=9494
rlabel metal2 1374 -895 1374 -895 0 net=10309
rlabel metal2 110 -897 110 -897 0 net=5373
rlabel metal2 387 -897 387 -897 0 net=5687
rlabel metal2 873 -897 873 -897 0 net=11711
rlabel metal2 114 -899 114 -899 0 net=3021
rlabel metal2 457 -899 457 -899 0 net=5157
rlabel metal2 691 -899 691 -899 0 net=8078
rlabel metal2 1206 -899 1206 -899 0 net=8805
rlabel metal2 1514 -899 1514 -899 0 net=11973
rlabel metal2 142 -901 142 -901 0 net=4409
rlabel metal2 499 -901 499 -901 0 net=4349
rlabel metal2 705 -901 705 -901 0 net=8406
rlabel metal2 1220 -901 1220 -901 0 net=8813
rlabel metal2 149 -903 149 -903 0 net=2225
rlabel metal2 184 -903 184 -903 0 net=5224
rlabel metal2 226 -903 226 -903 0 net=1910
rlabel metal2 275 -903 275 -903 0 net=1579
rlabel metal2 275 -903 275 -903 0 net=1579
rlabel metal2 296 -903 296 -903 0 net=1523
rlabel metal2 877 -903 877 -903 0 net=8054
rlabel metal2 1234 -903 1234 -903 0 net=9309
rlabel metal2 128 -905 128 -905 0 net=4539
rlabel metal2 184 -905 184 -905 0 net=1829
rlabel metal2 254 -905 254 -905 0 net=2129
rlabel metal2 254 -905 254 -905 0 net=2129
rlabel metal2 261 -905 261 -905 0 net=1933
rlabel metal2 303 -905 303 -905 0 net=1550
rlabel metal2 611 -905 611 -905 0 net=1695
rlabel metal2 964 -905 964 -905 0 net=11691
rlabel metal2 128 -907 128 -907 0 net=2585
rlabel metal2 796 -907 796 -907 0 net=9584
rlabel metal2 1395 -907 1395 -907 0 net=10661
rlabel metal2 138 -909 138 -909 0 net=2117
rlabel metal2 303 -909 303 -909 0 net=1551
rlabel metal2 586 -909 586 -909 0 net=8648
rlabel metal2 163 -911 163 -911 0 net=6904
rlabel metal2 1038 -911 1038 -911 0 net=7631
rlabel metal2 1248 -911 1248 -911 0 net=9313
rlabel metal2 1430 -911 1430 -911 0 net=10805
rlabel metal2 163 -913 163 -913 0 net=4879
rlabel metal2 331 -913 331 -913 0 net=2279
rlabel metal2 415 -913 415 -913 0 net=5189
rlabel metal2 768 -913 768 -913 0 net=11301
rlabel metal2 93 -915 93 -915 0 net=3745
rlabel metal2 373 -915 373 -915 0 net=4121
rlabel metal2 506 -915 506 -915 0 net=3225
rlabel metal2 506 -915 506 -915 0 net=3225
rlabel metal2 548 -915 548 -915 0 net=4107
rlabel metal2 786 -915 786 -915 0 net=11868
rlabel metal2 86 -917 86 -917 0 net=3681
rlabel metal2 166 -917 166 -917 0 net=3802
rlabel metal2 548 -917 548 -917 0 net=12059
rlabel metal2 170 -919 170 -919 0 net=2710
rlabel metal2 513 -919 513 -919 0 net=3075
rlabel metal2 912 -919 912 -919 0 net=9094
rlabel metal2 933 -919 933 -919 0 net=6551
rlabel metal2 1059 -919 1059 -919 0 net=10578
rlabel metal2 1486 -919 1486 -919 0 net=11471
rlabel metal2 170 -921 170 -921 0 net=2255
rlabel metal2 247 -921 247 -921 0 net=2053
rlabel metal2 310 -921 310 -921 0 net=2198
rlabel metal2 646 -921 646 -921 0 net=7273
rlabel metal2 733 -921 733 -921 0 net=7983
rlabel metal2 1493 -921 1493 -921 0 net=11837
rlabel metal2 191 -923 191 -923 0 net=6440
rlabel metal2 765 -923 765 -923 0 net=5199
rlabel metal2 810 -923 810 -923 0 net=12075
rlabel metal2 79 -925 79 -925 0 net=3541
rlabel metal2 198 -925 198 -925 0 net=4079
rlabel metal2 765 -925 765 -925 0 net=5936
rlabel metal2 1339 -925 1339 -925 0 net=9969
rlabel metal2 79 -927 79 -927 0 net=2539
rlabel metal2 569 -927 569 -927 0 net=3611
rlabel metal2 569 -927 569 -927 0 net=3611
rlabel metal2 576 -927 576 -927 0 net=4373
rlabel metal2 856 -927 856 -927 0 net=6401
rlabel metal2 919 -927 919 -927 0 net=6445
rlabel metal2 968 -927 968 -927 0 net=7419
rlabel metal2 975 -927 975 -927 0 net=6855
rlabel metal2 1062 -927 1062 -927 0 net=9924
rlabel metal2 1437 -927 1437 -927 0 net=10863
rlabel metal2 124 -929 124 -929 0 net=494
rlabel metal2 205 -929 205 -929 0 net=3331
rlabel metal2 646 -929 646 -929 0 net=7905
rlabel metal2 1101 -929 1101 -929 0 net=7937
rlabel metal2 1262 -929 1262 -929 0 net=9371
rlabel metal2 1444 -929 1444 -929 0 net=11779
rlabel metal2 226 -931 226 -931 0 net=2171
rlabel metal2 583 -931 583 -931 0 net=5657
rlabel metal2 772 -931 772 -931 0 net=5481
rlabel metal2 1458 -931 1458 -931 0 net=11227
rlabel metal2 229 -933 229 -933 0 net=8024
rlabel metal2 1150 -933 1150 -933 0 net=10439
rlabel metal2 1458 -933 1458 -933 0 net=11879
rlabel metal2 121 -935 121 -935 0 net=10589
rlabel metal2 233 -937 233 -937 0 net=11418
rlabel metal2 89 -939 89 -939 0 net=3781
rlabel metal2 236 -939 236 -939 0 net=11667
rlabel metal2 240 -941 240 -941 0 net=3735
rlabel metal2 373 -941 373 -941 0 net=2465
rlabel metal2 436 -941 436 -941 0 net=3997
rlabel metal2 1255 -941 1255 -941 0 net=10745
rlabel metal2 261 -943 261 -943 0 net=2661
rlabel metal2 436 -943 436 -943 0 net=5217
rlabel metal2 730 -943 730 -943 0 net=5545
rlabel metal2 856 -943 856 -943 0 net=10975
rlabel metal2 289 -945 289 -945 0 net=8005
rlabel metal2 1255 -945 1255 -945 0 net=10185
rlabel metal2 1276 -945 1276 -945 0 net=9379
rlabel metal2 1276 -945 1276 -945 0 net=9379
rlabel metal2 1297 -945 1297 -945 0 net=9717
rlabel metal2 37 -947 37 -947 0 net=8533
rlabel metal2 1304 -947 1304 -947 0 net=9791
rlabel metal2 313 -949 313 -949 0 net=2369
rlabel metal2 345 -949 345 -949 0 net=5269
rlabel metal2 576 -949 576 -949 0 net=4749
rlabel metal2 709 -949 709 -949 0 net=2560
rlabel metal2 863 -949 863 -949 0 net=6519
rlabel metal2 940 -949 940 -949 0 net=6643
rlabel metal2 1178 -949 1178 -949 0 net=8713
rlabel metal2 1346 -949 1346 -949 0 net=10191
rlabel metal2 1381 -949 1381 -949 0 net=6003
rlabel metal2 317 -951 317 -951 0 net=1607
rlabel metal2 474 -951 474 -951 0 net=4682
rlabel metal2 800 -951 800 -951 0 net=6083
rlabel metal2 968 -951 968 -951 0 net=7303
rlabel metal2 1031 -951 1031 -951 0 net=7375
rlabel metal2 1353 -951 1353 -951 0 net=10069
rlabel metal2 345 -953 345 -953 0 net=2715
rlabel metal2 394 -953 394 -953 0 net=2289
rlabel metal2 429 -953 429 -953 0 net=6179
rlabel metal2 632 -953 632 -953 0 net=6859
rlabel metal2 849 -953 849 -953 0 net=5523
rlabel metal2 870 -953 870 -953 0 net=9643
rlabel metal2 107 -955 107 -955 0 net=9135
rlabel metal2 870 -955 870 -955 0 net=7745
rlabel metal2 1199 -955 1199 -955 0 net=8799
rlabel metal2 1353 -955 1353 -955 0 net=10681
rlabel metal2 352 -957 352 -957 0 net=2325
rlabel metal2 394 -957 394 -957 0 net=3795
rlabel metal2 800 -957 800 -957 0 net=5979
rlabel metal2 877 -957 877 -957 0 net=10086
rlabel metal2 366 -959 366 -959 0 net=3183
rlabel metal2 478 -959 478 -959 0 net=2109
rlabel metal2 604 -959 604 -959 0 net=4645
rlabel metal2 751 -959 751 -959 0 net=5283
rlabel metal2 884 -959 884 -959 0 net=6745
rlabel metal2 898 -959 898 -959 0 net=8782
rlabel metal2 1283 -959 1283 -959 0 net=9471
rlabel metal2 37 -961 37 -961 0 net=3507
rlabel metal2 520 -961 520 -961 0 net=3433
rlabel metal2 604 -961 604 -961 0 net=11175
rlabel metal2 380 -963 380 -963 0 net=2905
rlabel metal2 492 -963 492 -963 0 net=2613
rlabel metal2 527 -963 527 -963 0 net=4851
rlabel metal2 884 -963 884 -963 0 net=7023
rlabel metal2 1003 -963 1003 -963 0 net=7207
rlabel metal2 1115 -963 1115 -963 0 net=8117
rlabel metal2 1290 -963 1290 -963 0 net=9539
rlabel metal2 44 -965 44 -965 0 net=2961
rlabel metal2 534 -965 534 -965 0 net=5365
rlabel metal2 947 -965 947 -965 0 net=6785
rlabel metal2 1052 -965 1052 -965 0 net=7793
rlabel metal2 1213 -965 1213 -965 0 net=11517
rlabel metal2 44 -967 44 -967 0 net=295
rlabel metal2 58 -967 58 -967 0 net=3573
rlabel metal2 537 -967 537 -967 0 net=9063
rlabel metal2 975 -967 975 -967 0 net=9623
rlabel metal2 54 -969 54 -969 0 net=11310
rlabel metal2 58 -971 58 -971 0 net=8235
rlabel metal2 1164 -971 1164 -971 0 net=8505
rlabel metal2 100 -973 100 -973 0 net=8819
rlabel metal2 23 -975 23 -975 0 net=5499
rlabel metal2 219 -975 219 -975 0 net=7285
rlabel metal2 978 -975 978 -975 0 net=174
rlabel metal2 359 -977 359 -977 0 net=3131
rlabel metal2 551 -977 551 -977 0 net=5206
rlabel metal2 880 -977 880 -977 0 net=10671
rlabel metal2 1129 -977 1129 -977 0 net=8205
rlabel metal2 212 -979 212 -979 0 net=1967
rlabel metal2 443 -979 443 -979 0 net=5571
rlabel metal2 744 -979 744 -979 0 net=5159
rlabel metal2 1003 -979 1003 -979 0 net=7969
rlabel metal2 1122 -979 1122 -979 0 net=8145
rlabel metal2 1164 -979 1164 -979 0 net=8679
rlabel metal2 156 -981 156 -981 0 net=3927
rlabel metal2 467 -981 467 -981 0 net=7247
rlabel metal2 156 -983 156 -983 0 net=4407
rlabel metal2 835 -983 835 -983 0 net=5755
rlabel metal2 212 -985 212 -985 0 net=3675
rlabel metal2 614 -985 614 -985 0 net=5225
rlabel metal2 835 -985 835 -985 0 net=6139
rlabel metal2 1024 -985 1024 -985 0 net=7343
rlabel metal2 541 -987 541 -987 0 net=3101
rlabel metal2 618 -987 618 -987 0 net=4359
rlabel metal2 796 -987 796 -987 0 net=6755
rlabel metal2 1045 -987 1045 -987 0 net=7685
rlabel metal2 625 -989 625 -989 0 net=5450
rlabel metal2 842 -989 842 -989 0 net=9001
rlabel metal2 639 -991 639 -991 0 net=7743
rlabel metal2 639 -993 639 -993 0 net=3973
rlabel metal2 954 -993 954 -993 0 net=6795
rlabel metal2 1062 -993 1062 -993 0 net=10632
rlabel metal2 681 -995 681 -995 0 net=8421
rlabel metal2 789 -997 789 -997 0 net=10225
rlabel metal2 954 -999 954 -999 0 net=10144
rlabel metal2 989 -1001 989 -1001 0 net=7031
rlabel metal2 1066 -1001 1066 -1001 0 net=7831
rlabel metal2 1451 -1001 1451 -1001 0 net=11039
rlabel metal2 989 -1003 989 -1003 0 net=10951
rlabel metal2 1010 -1005 1010 -1005 0 net=7217
rlabel metal2 1311 -1005 1311 -1005 0 net=9817
rlabel metal2 534 -1007 534 -1007 0 net=7443
rlabel metal2 1066 -1009 1066 -1009 0 net=8830
rlabel metal2 1073 -1011 1073 -1011 0 net=7861
rlabel metal2 1402 -1011 1402 -1011 0 net=11933
rlabel metal2 628 -1013 628 -1013 0 net=7053
rlabel metal2 1080 -1013 1080 -1013 0 net=7877
rlabel metal2 779 -1015 779 -1015 0 net=7059
rlabel metal2 779 -1017 779 -1017 0 net=5829
rlabel metal2 828 -1017 828 -1017 0 net=6411
rlabel metal2 807 -1019 807 -1019 0 net=6627
rlabel metal2 828 -1021 828 -1021 0 net=9714
rlabel metal2 1360 -1023 1360 -1023 0 net=11381
rlabel metal2 1318 -1025 1318 -1025 0 net=9927
rlabel metal2 1185 -1027 1185 -1027 0 net=8761
rlabel metal2 1185 -1029 1185 -1029 0 net=8997
rlabel metal2 1087 -1031 1087 -1031 0 net=7893
rlabel metal2 201 -1033 201 -1033 0 net=7123
rlabel metal2 44 -1044 44 -1044 0 net=3737
rlabel metal2 261 -1044 261 -1044 0 net=2662
rlabel metal2 653 -1044 653 -1044 0 net=4043
rlabel metal2 653 -1044 653 -1044 0 net=4043
rlabel metal2 681 -1044 681 -1044 0 net=6644
rlabel metal2 1710 -1044 1710 -1044 0 net=8861
rlabel metal2 65 -1046 65 -1046 0 net=3002
rlabel metal2 499 -1046 499 -1046 0 net=4123
rlabel metal2 681 -1046 681 -1046 0 net=4361
rlabel metal2 719 -1046 719 -1046 0 net=10310
rlabel metal2 1724 -1046 1724 -1046 0 net=6281
rlabel metal2 1724 -1046 1724 -1046 0 net=6281
rlabel metal2 65 -1048 65 -1048 0 net=3965
rlabel metal2 579 -1048 579 -1048 0 net=7744
rlabel metal2 86 -1050 86 -1050 0 net=6084
rlabel metal2 957 -1050 957 -1050 0 net=9310
rlabel metal2 89 -1052 89 -1052 0 net=10976
rlabel metal2 1626 -1052 1626 -1052 0 net=11839
rlabel metal2 93 -1054 93 -1054 0 net=3682
rlabel metal2 198 -1054 198 -1054 0 net=2280
rlabel metal2 408 -1054 408 -1054 0 net=2290
rlabel metal2 590 -1054 590 -1054 0 net=8806
rlabel metal2 51 -1056 51 -1056 0 net=4247
rlabel metal2 597 -1056 597 -1056 0 net=5572
rlabel metal2 723 -1056 723 -1056 0 net=8814
rlabel metal2 51 -1058 51 -1058 0 net=3435
rlabel metal2 600 -1058 600 -1058 0 net=6628
rlabel metal2 1062 -1058 1062 -1058 0 net=10737
rlabel metal2 93 -1060 93 -1060 0 net=3929
rlabel metal2 450 -1060 450 -1060 0 net=3037
rlabel metal2 513 -1060 513 -1060 0 net=3077
rlabel metal2 569 -1060 569 -1060 0 net=3612
rlabel metal2 614 -1060 614 -1060 0 net=5366
rlabel metal2 940 -1060 940 -1060 0 net=6857
rlabel metal2 1069 -1060 1069 -1060 0 net=11974
rlabel metal2 54 -1062 54 -1062 0 net=2823
rlabel metal2 450 -1062 450 -1062 0 net=2615
rlabel metal2 527 -1062 527 -1062 0 net=3132
rlabel metal2 726 -1062 726 -1062 0 net=1239
rlabel metal2 751 -1062 751 -1062 0 net=4852
rlabel metal2 810 -1062 810 -1062 0 net=6796
rlabel metal2 1129 -1062 1129 -1062 0 net=8147
rlabel metal2 1129 -1062 1129 -1062 0 net=8147
rlabel metal2 1143 -1062 1143 -1062 0 net=7939
rlabel metal2 1360 -1062 1360 -1062 0 net=11383
rlabel metal2 100 -1064 100 -1064 0 net=5500
rlabel metal2 292 -1064 292 -1064 0 net=139
rlabel metal2 702 -1064 702 -1064 0 net=4375
rlabel metal2 751 -1064 751 -1064 0 net=6004
rlabel metal2 1500 -1064 1500 -1064 0 net=11519
rlabel metal2 103 -1066 103 -1066 0 net=5482
rlabel metal2 1612 -1066 1612 -1066 0 net=11713
rlabel metal2 107 -1068 107 -1068 0 net=5190
rlabel metal2 464 -1068 464 -1068 0 net=7286
rlabel metal2 971 -1068 971 -1068 0 net=1068
rlabel metal2 1234 -1068 1234 -1068 0 net=6701
rlabel metal2 107 -1070 107 -1070 0 net=4195
rlabel metal2 758 -1070 758 -1070 0 net=7894
rlabel metal2 1276 -1070 1276 -1070 0 net=9381
rlabel metal2 1367 -1070 1367 -1070 0 net=9971
rlabel metal2 89 -1072 89 -1072 0 net=11767
rlabel metal2 110 -1074 110 -1074 0 net=9928
rlabel metal2 121 -1076 121 -1076 0 net=3998
rlabel metal2 1227 -1076 1227 -1076 0 net=8507
rlabel metal2 1381 -1076 1381 -1076 0 net=10807
rlabel metal2 121 -1078 121 -1078 0 net=5218
rlabel metal2 478 -1078 478 -1078 0 net=2111
rlabel metal2 621 -1078 621 -1078 0 net=8747
rlabel metal2 1290 -1078 1290 -1078 0 net=9473
rlabel metal2 1479 -1078 1479 -1078 0 net=11669
rlabel metal2 128 -1080 128 -1080 0 net=2587
rlabel metal2 506 -1080 506 -1080 0 net=3227
rlabel metal2 621 -1080 621 -1080 0 net=5756
rlabel metal2 1388 -1080 1388 -1080 0 net=9625
rlabel metal2 1640 -1080 1640 -1080 0 net=12001
rlabel metal2 128 -1082 128 -1082 0 net=5161
rlabel metal2 768 -1082 768 -1082 0 net=7376
rlabel metal2 1402 -1082 1402 -1082 0 net=11935
rlabel metal2 135 -1084 135 -1084 0 net=2902
rlabel metal2 506 -1084 506 -1084 0 net=7248
rlabel metal2 1255 -1084 1255 -1084 0 net=10187
rlabel metal2 1619 -1084 1619 -1084 0 net=11229
rlabel metal2 135 -1086 135 -1086 0 net=3333
rlabel metal2 208 -1086 208 -1086 0 net=7444
rlabel metal2 1339 -1086 1339 -1086 0 net=9315
rlabel metal2 1409 -1086 1409 -1086 0 net=9819
rlabel metal2 142 -1088 142 -1088 0 net=4411
rlabel metal2 628 -1088 628 -1088 0 net=10213
rlabel metal2 142 -1090 142 -1090 0 net=2227
rlabel metal2 166 -1090 166 -1090 0 net=1093
rlabel metal2 219 -1090 219 -1090 0 net=2055
rlabel metal2 261 -1090 261 -1090 0 net=1543
rlabel metal2 845 -1090 845 -1090 0 net=10440
rlabel metal2 1241 -1090 1241 -1090 0 net=8535
rlabel metal2 1311 -1090 1311 -1090 0 net=9645
rlabel metal2 149 -1092 149 -1092 0 net=1552
rlabel metal2 310 -1092 310 -1092 0 net=2371
rlabel metal2 352 -1092 352 -1092 0 net=2327
rlabel metal2 352 -1092 352 -1092 0 net=2327
rlabel metal2 359 -1092 359 -1092 0 net=1969
rlabel metal2 513 -1092 513 -1092 0 net=4750
rlabel metal2 702 -1092 702 -1092 0 net=6413
rlabel metal2 1437 -1092 1437 -1092 0 net=11881
rlabel metal2 170 -1094 170 -1094 0 net=2257
rlabel metal2 516 -1094 516 -1094 0 net=4901
rlabel metal2 786 -1094 786 -1094 0 net=5200
rlabel metal2 859 -1094 859 -1094 0 net=10603
rlabel metal2 170 -1096 170 -1096 0 net=3543
rlabel metal2 212 -1096 212 -1096 0 net=3677
rlabel metal2 331 -1096 331 -1096 0 net=2717
rlabel metal2 359 -1096 359 -1096 0 net=2963
rlabel metal2 520 -1096 520 -1096 0 net=3103
rlabel metal2 733 -1096 733 -1096 0 net=8367
rlabel metal2 1297 -1096 1297 -1096 0 net=9541
rlabel metal2 1458 -1096 1458 -1096 0 net=10227
rlabel metal2 47 -1098 47 -1098 0 net=710
rlabel metal2 744 -1098 744 -1098 0 net=6552
rlabel metal2 1010 -1098 1010 -1098 0 net=7209
rlabel metal2 1122 -1098 1122 -1098 0 net=7747
rlabel metal2 1346 -1098 1346 -1098 0 net=10193
rlabel metal2 1472 -1098 1472 -1098 0 net=10663
rlabel metal2 79 -1100 79 -1100 0 net=2541
rlabel metal2 212 -1100 212 -1100 0 net=2131
rlabel metal2 282 -1100 282 -1100 0 net=1935
rlabel metal2 366 -1100 366 -1100 0 net=3184
rlabel metal2 485 -1100 485 -1100 0 net=11171
rlabel metal2 79 -1102 79 -1102 0 net=8820
rlabel metal2 163 -1104 163 -1104 0 net=4880
rlabel metal2 275 -1104 275 -1104 0 net=1581
rlabel metal2 289 -1104 289 -1104 0 net=1609
rlabel metal2 366 -1104 366 -1104 0 net=6145
rlabel metal2 793 -1104 793 -1104 0 net=10864
rlabel metal2 114 -1106 114 -1106 0 net=3023
rlabel metal2 380 -1106 380 -1106 0 net=2907
rlabel metal2 807 -1106 807 -1106 0 net=7055
rlabel metal2 1115 -1106 1115 -1106 0 net=10673
rlabel metal2 114 -1108 114 -1108 0 net=5831
rlabel metal2 842 -1108 842 -1108 0 net=5325
rlabel metal2 1073 -1108 1073 -1108 0 net=7125
rlabel metal2 1115 -1108 1115 -1108 0 net=7687
rlabel metal2 1178 -1108 1178 -1108 0 net=7879
rlabel metal2 1332 -1108 1332 -1108 0 net=9003
rlabel metal2 1374 -1108 1374 -1108 0 net=11473
rlabel metal2 156 -1110 156 -1110 0 net=4408
rlabel metal2 296 -1110 296 -1110 0 net=1525
rlabel metal2 296 -1110 296 -1110 0 net=1525
rlabel metal2 380 -1110 380 -1110 0 net=4135
rlabel metal2 723 -1110 723 -1110 0 net=8299
rlabel metal2 1528 -1110 1528 -1110 0 net=10953
rlabel metal2 1556 -1110 1556 -1110 0 net=11177
rlabel metal2 156 -1112 156 -1112 0 net=7907
rlabel metal2 772 -1112 772 -1112 0 net=5547
rlabel metal2 849 -1112 849 -1112 0 net=9137
rlabel metal2 1542 -1112 1542 -1112 0 net=11781
rlabel metal2 75 -1114 75 -1114 0 net=6067
rlabel metal2 856 -1114 856 -1114 0 net=7495
rlabel metal2 1150 -1114 1150 -1114 0 net=8007
rlabel metal2 177 -1116 177 -1116 0 net=4540
rlabel metal2 646 -1116 646 -1116 0 net=4109
rlabel metal2 674 -1116 674 -1116 0 net=5227
rlabel metal2 835 -1116 835 -1116 0 net=6141
rlabel metal2 870 -1116 870 -1116 0 net=7327
rlabel metal2 1164 -1116 1164 -1116 0 net=8681
rlabel metal2 1248 -1116 1248 -1116 0 net=8801
rlabel metal2 177 -1118 177 -1118 0 net=1665
rlabel metal2 201 -1120 201 -1120 0 net=7463
rlabel metal2 1164 -1120 1164 -1120 0 net=8119
rlabel metal2 201 -1122 201 -1122 0 net=5158
rlabel metal2 537 -1122 537 -1122 0 net=4251
rlabel metal2 821 -1122 821 -1122 0 net=5284
rlabel metal2 873 -1122 873 -1122 0 net=10070
rlabel metal2 205 -1124 205 -1124 0 net=11707
rlabel metal2 236 -1126 236 -1126 0 net=8589
rlabel metal2 1353 -1126 1353 -1126 0 net=10683
rlabel metal2 240 -1128 240 -1128 0 net=3975
rlabel metal2 667 -1128 667 -1128 0 net=4351
rlabel metal2 821 -1128 821 -1128 0 net=7219
rlabel metal2 1185 -1128 1185 -1128 0 net=8999
rlabel metal2 1353 -1128 1353 -1128 0 net=9373
rlabel metal2 58 -1130 58 -1130 0 net=8237
rlabel metal2 835 -1130 835 -1130 0 net=7305
rlabel metal2 975 -1130 975 -1130 0 net=6787
rlabel metal2 1038 -1130 1038 -1130 0 net=7863
rlabel metal2 1395 -1130 1395 -1130 0 net=9793
rlabel metal2 58 -1132 58 -1132 0 net=6041
rlabel metal2 877 -1132 877 -1132 0 net=11899
rlabel metal2 247 -1134 247 -1134 0 net=2119
rlabel metal2 387 -1134 387 -1134 0 net=5689
rlabel metal2 625 -1134 625 -1134 0 net=4669
rlabel metal2 978 -1134 978 -1134 0 net=11361
rlabel metal2 163 -1136 163 -1136 0 net=5705
rlabel metal2 394 -1136 394 -1136 0 net=3796
rlabel metal2 894 -1136 894 -1136 0 net=9929
rlabel metal2 1444 -1136 1444 -1136 0 net=10591
rlabel metal2 226 -1138 226 -1138 0 net=2173
rlabel metal2 394 -1138 394 -1138 0 net=3891
rlabel metal2 877 -1138 877 -1138 0 net=7025
rlabel metal2 898 -1138 898 -1138 0 net=11302
rlabel metal2 30 -1140 30 -1140 0 net=4399
rlabel metal2 401 -1140 401 -1140 0 net=2239
rlabel metal2 639 -1140 639 -1140 0 net=4691
rlabel metal2 898 -1140 898 -1140 0 net=10703
rlabel metal2 1598 -1140 1598 -1140 0 net=10519
rlabel metal2 30 -1142 30 -1142 0 net=5659
rlabel metal2 709 -1142 709 -1142 0 net=4647
rlabel metal2 905 -1142 905 -1142 0 net=5697
rlabel metal2 905 -1142 905 -1142 0 net=5697
rlabel metal2 912 -1142 912 -1142 0 net=6402
rlabel metal2 989 -1142 989 -1142 0 net=9718
rlabel metal2 233 -1144 233 -1144 0 net=3783
rlabel metal2 709 -1144 709 -1144 0 net=4509
rlabel metal2 1101 -1144 1101 -1144 0 net=7633
rlabel metal2 1563 -1144 1563 -1144 0 net=11041
rlabel metal2 422 -1146 422 -1146 0 net=5293
rlabel metal2 912 -1146 912 -1146 0 net=6521
rlabel metal2 933 -1146 933 -1146 0 net=9065
rlabel metal2 1563 -1146 1563 -1146 0 net=11223
rlabel metal2 422 -1148 422 -1148 0 net=2747
rlabel metal2 726 -1148 726 -1148 0 net=5555
rlabel metal2 947 -1148 947 -1148 0 net=6747
rlabel metal2 989 -1148 989 -1148 0 net=9979
rlabel metal2 1591 -1148 1591 -1148 0 net=11693
rlabel metal2 324 -1150 324 -1150 0 net=3747
rlabel metal2 765 -1150 765 -1150 0 net=6571
rlabel metal2 954 -1150 954 -1150 0 net=10746
rlabel metal2 1647 -1150 1647 -1150 0 net=6626
rlabel metal2 100 -1152 100 -1152 0 net=2921
rlabel metal2 429 -1152 429 -1152 0 net=6181
rlabel metal2 814 -1152 814 -1152 0 net=6861
rlabel metal2 992 -1152 992 -1152 0 net=9615
rlabel metal2 1570 -1152 1570 -1152 0 net=12061
rlabel metal2 373 -1154 373 -1154 0 net=2467
rlabel metal2 457 -1154 457 -1154 0 net=1697
rlabel metal2 814 -1154 814 -1154 0 net=5525
rlabel metal2 919 -1154 919 -1154 0 net=6447
rlabel metal2 992 -1154 992 -1154 0 net=7984
rlabel metal2 373 -1156 373 -1156 0 net=4081
rlabel metal2 800 -1156 800 -1156 0 net=5981
rlabel metal2 996 -1156 996 -1156 0 net=6757
rlabel metal2 1031 -1156 1031 -1156 0 net=7275
rlabel metal2 1157 -1156 1157 -1156 0 net=8423
rlabel metal2 1486 -1156 1486 -1156 0 net=12077
rlabel metal2 338 -1158 338 -1158 0 net=5375
rlabel metal2 831 -1158 831 -1158 0 net=7083
rlabel metal2 1003 -1158 1003 -1158 0 net=7971
rlabel metal2 1283 -1158 1283 -1158 0 net=8763
rlabel metal2 184 -1160 184 -1160 0 net=1831
rlabel metal2 471 -1160 471 -1160 0 net=6403
rlabel metal2 957 -1160 957 -1160 0 net=9035
rlabel metal2 37 -1162 37 -1162 0 net=3509
rlabel metal2 562 -1162 562 -1162 0 net=5271
rlabel metal2 1003 -1162 1003 -1162 0 net=7033
rlabel metal2 37 -1164 37 -1164 0 net=4245
rlabel metal2 124 -1164 124 -1164 0 net=7445
rlabel metal2 184 -1166 184 -1166 0 net=4803
rlabel metal2 492 -1166 492 -1166 0 net=3575
rlabel metal2 611 -1166 611 -1166 0 net=5670
rlabel metal2 1017 -1166 1017 -1166 0 net=7421
rlabel metal2 492 -1168 492 -1168 0 net=4381
rlabel metal2 1017 -1168 1017 -1168 0 net=7061
rlabel metal2 635 -1170 635 -1170 0 net=7675
rlabel metal2 660 -1172 660 -1172 0 net=7794
rlabel metal2 901 -1174 901 -1174 0 net=8243
rlabel metal2 1024 -1176 1024 -1176 0 net=7345
rlabel metal2 1080 -1178 1080 -1178 0 net=8207
rlabel metal2 1136 -1180 1136 -1180 0 net=7833
rlabel metal2 1269 -1180 1269 -1180 0 net=8715
rlabel metal2 597 -1182 597 -1182 0 net=8523
rlabel metal2 607 -1184 607 -1184 0 net=9175
rlabel metal2 23 -1195 23 -1195 0 net=3967
rlabel metal2 79 -1195 79 -1195 0 net=1679
rlabel metal2 124 -1195 124 -1195 0 net=7688
rlabel metal2 1318 -1195 1318 -1195 0 net=9037
rlabel metal2 1318 -1195 1318 -1195 0 net=9037
rlabel metal2 1486 -1195 1486 -1195 0 net=12079
rlabel metal2 1717 -1195 1717 -1195 0 net=6283
rlabel metal2 1731 -1195 1731 -1195 0 net=8863
rlabel metal2 30 -1197 30 -1197 0 net=5660
rlabel metal2 93 -1197 93 -1197 0 net=3930
rlabel metal2 149 -1197 149 -1197 0 net=886
rlabel metal2 208 -1197 208 -1197 0 net=6182
rlabel metal2 810 -1197 810 -1197 0 net=7306
rlabel metal2 873 -1197 873 -1197 0 net=11042
rlabel metal2 1605 -1197 1605 -1197 0 net=11709
rlabel metal2 30 -1199 30 -1199 0 net=3817
rlabel metal2 506 -1199 506 -1199 0 net=2908
rlabel metal2 723 -1199 723 -1199 0 net=7972
rlabel metal2 1451 -1199 1451 -1199 0 net=10215
rlabel metal2 1500 -1199 1500 -1199 0 net=11521
rlabel metal2 1619 -1199 1619 -1199 0 net=11901
rlabel metal2 1675 -1199 1675 -1199 0 net=11230
rlabel metal2 58 -1201 58 -1201 0 net=6042
rlabel metal2 135 -1201 135 -1201 0 net=3334
rlabel metal2 541 -1201 541 -1201 0 net=4511
rlabel metal2 744 -1201 744 -1201 0 net=7834
rlabel metal2 1185 -1201 1185 -1201 0 net=9067
rlabel metal2 1465 -1201 1465 -1201 0 net=11769
rlabel metal2 1633 -1201 1633 -1201 0 net=10521
rlabel metal2 1633 -1201 1633 -1201 0 net=10521
rlabel metal2 1654 -1201 1654 -1201 0 net=11937
rlabel metal2 58 -1203 58 -1203 0 net=2121
rlabel metal2 250 -1203 250 -1203 0 net=2328
rlabel metal2 380 -1203 380 -1203 0 net=4137
rlabel metal2 744 -1203 744 -1203 0 net=5549
rlabel metal2 814 -1203 814 -1203 0 net=5526
rlabel metal2 901 -1203 901 -1203 0 net=10592
rlabel metal2 1591 -1203 1591 -1203 0 net=11695
rlabel metal2 1661 -1203 1661 -1203 0 net=10071
rlabel metal2 65 -1205 65 -1205 0 net=1539
rlabel metal2 205 -1205 205 -1205 0 net=1761
rlabel metal2 593 -1205 593 -1205 0 net=9980
rlabel metal2 1416 -1205 1416 -1205 0 net=9931
rlabel metal2 1542 -1205 1542 -1205 0 net=11783
rlabel metal2 96 -1207 96 -1207 0 net=10604
rlabel metal2 1528 -1207 1528 -1207 0 net=10955
rlabel metal2 121 -1209 121 -1209 0 net=10738
rlabel metal2 135 -1211 135 -1211 0 net=2965
rlabel metal2 380 -1211 380 -1211 0 net=2175
rlabel metal2 422 -1211 422 -1211 0 net=2748
rlabel metal2 530 -1211 530 -1211 0 net=7471
rlabel metal2 1206 -1211 1206 -1211 0 net=9617
rlabel metal2 1521 -1211 1521 -1211 0 net=12063
rlabel metal2 142 -1213 142 -1213 0 net=2229
rlabel metal2 163 -1213 163 -1213 0 net=9542
rlabel metal2 1325 -1213 1325 -1213 0 net=9795
rlabel metal2 1416 -1213 1416 -1213 0 net=11671
rlabel metal2 142 -1215 142 -1215 0 net=7748
rlabel metal2 1129 -1215 1129 -1215 0 net=8149
rlabel metal2 1241 -1215 1241 -1215 0 net=8537
rlabel metal2 1339 -1215 1339 -1215 0 net=9317
rlabel metal2 1409 -1215 1409 -1215 0 net=9821
rlabel metal2 124 -1217 124 -1217 0 net=9323
rlabel metal2 1437 -1217 1437 -1217 0 net=11883
rlabel metal2 163 -1219 163 -1219 0 net=8524
rlabel metal2 1213 -1219 1213 -1219 0 net=8301
rlabel metal2 1290 -1219 1290 -1219 0 net=9475
rlabel metal2 166 -1221 166 -1221 0 net=2455
rlabel metal2 492 -1221 492 -1221 0 net=4383
rlabel metal2 814 -1221 814 -1221 0 net=12002
rlabel metal2 166 -1223 166 -1223 0 net=8
rlabel metal2 492 -1223 492 -1223 0 net=4693
rlabel metal2 674 -1223 674 -1223 0 net=4253
rlabel metal2 768 -1223 768 -1223 0 net=12025
rlabel metal2 184 -1225 184 -1225 0 net=8238
rlabel metal2 695 -1225 695 -1225 0 net=3793
rlabel metal2 982 -1225 982 -1225 0 net=6863
rlabel metal2 1013 -1225 1013 -1225 0 net=9972
rlabel metal2 1374 -1225 1374 -1225 0 net=11475
rlabel metal2 82 -1227 82 -1227 0 net=7091
rlabel metal2 198 -1227 198 -1227 0 net=55
rlabel metal2 513 -1227 513 -1227 0 net=10311
rlabel metal2 198 -1229 198 -1229 0 net=4671
rlabel metal2 639 -1229 639 -1229 0 net=4045
rlabel metal2 709 -1229 709 -1229 0 net=4205
rlabel metal2 772 -1229 772 -1229 0 net=5229
rlabel metal2 894 -1229 894 -1229 0 net=6522
rlabel metal2 936 -1229 936 -1229 0 net=11840
rlabel metal2 156 -1231 156 -1231 0 net=7908
rlabel metal2 646 -1231 646 -1231 0 net=4111
rlabel metal2 828 -1231 828 -1231 0 net=10361
rlabel metal2 1535 -1231 1535 -1231 0 net=11173
rlabel metal2 156 -1233 156 -1233 0 net=1799
rlabel metal2 646 -1233 646 -1233 0 net=3979
rlabel metal2 831 -1233 831 -1233 0 net=6858
rlabel metal2 957 -1233 957 -1233 0 net=11362
rlabel metal2 233 -1235 233 -1235 0 net=2718
rlabel metal2 352 -1235 352 -1235 0 net=2617
rlabel metal2 478 -1235 478 -1235 0 net=4805
rlabel metal2 884 -1235 884 -1235 0 net=6405
rlabel metal2 971 -1235 971 -1235 0 net=10674
rlabel metal2 212 -1237 212 -1237 0 net=2133
rlabel metal2 387 -1237 387 -1237 0 net=3039
rlabel metal2 576 -1237 576 -1237 0 net=10441
rlabel metal2 191 -1239 191 -1239 0 net=2543
rlabel metal2 233 -1239 233 -1239 0 net=4721
rlabel metal2 597 -1239 597 -1239 0 net=10873
rlabel metal2 177 -1241 177 -1241 0 net=1667
rlabel metal2 236 -1241 236 -1241 0 net=9753
rlabel metal2 1472 -1241 1472 -1241 0 net=10665
rlabel metal2 177 -1243 177 -1243 0 net=2057
rlabel metal2 240 -1243 240 -1243 0 net=3977
rlabel metal2 653 -1243 653 -1243 0 net=2401
rlabel metal2 975 -1243 975 -1243 0 net=6789
rlabel metal2 1276 -1243 1276 -1243 0 net=8749
rlabel metal2 1356 -1243 1356 -1243 0 net=10977
rlabel metal2 219 -1245 219 -1245 0 net=4385
rlabel metal2 821 -1245 821 -1245 0 net=7221
rlabel metal2 898 -1245 898 -1245 0 net=5699
rlabel metal2 975 -1245 975 -1245 0 net=138
rlabel metal2 1045 -1245 1045 -1245 0 net=11178
rlabel metal2 152 -1247 152 -1247 0 net=5725
rlabel metal2 982 -1247 982 -1247 0 net=9000
rlabel metal2 1381 -1247 1381 -1247 0 net=10809
rlabel metal2 240 -1249 240 -1249 0 net=2069
rlabel metal2 821 -1249 821 -1249 0 net=7210
rlabel metal2 1031 -1249 1031 -1249 0 net=7277
rlabel metal2 1395 -1249 1395 -1249 0 net=8611
rlabel metal2 254 -1251 254 -1251 0 net=1937
rlabel metal2 394 -1251 394 -1251 0 net=3893
rlabel metal2 478 -1251 478 -1251 0 net=3228
rlabel metal2 544 -1251 544 -1251 0 net=9193
rlabel metal2 1423 -1251 1423 -1251 0 net=10195
rlabel metal2 1556 -1251 1556 -1251 0 net=11165
rlabel metal2 37 -1253 37 -1253 0 net=4246
rlabel metal2 562 -1253 562 -1253 0 net=3577
rlabel metal2 611 -1253 611 -1253 0 net=948
rlabel metal2 989 -1253 989 -1253 0 net=7328
rlabel metal2 1080 -1253 1080 -1253 0 net=8209
rlabel metal2 1388 -1253 1388 -1253 0 net=9627
rlabel metal2 1612 -1253 1612 -1253 0 net=11715
rlabel metal2 37 -1255 37 -1255 0 net=3749
rlabel metal2 614 -1255 614 -1255 0 net=11109
rlabel metal2 278 -1257 278 -1257 0 net=7056
rlabel metal2 989 -1257 989 -1257 0 net=7465
rlabel metal2 1108 -1257 1108 -1257 0 net=7677
rlabel metal2 1549 -1257 1549 -1257 0 net=11385
rlabel metal2 296 -1259 296 -1259 0 net=1527
rlabel metal2 296 -1259 296 -1259 0 net=1527
rlabel metal2 310 -1259 310 -1259 0 net=2372
rlabel metal2 548 -1259 548 -1259 0 net=3079
rlabel metal2 751 -1259 751 -1259 0 net=9287
rlabel metal2 1493 -1259 1493 -1259 0 net=10685
rlabel metal2 310 -1261 310 -1261 0 net=1805
rlabel metal2 471 -1261 471 -1261 0 net=3511
rlabel metal2 751 -1261 751 -1261 0 net=4903
rlabel metal2 807 -1261 807 -1261 0 net=7351
rlabel metal2 1129 -1261 1129 -1261 0 net=8509
rlabel metal2 1255 -1261 1255 -1261 0 net=8591
rlabel metal2 317 -1263 317 -1263 0 net=3024
rlabel metal2 1003 -1263 1003 -1263 0 net=7035
rlabel metal2 1108 -1263 1108 -1263 0 net=9375
rlabel metal2 282 -1265 282 -1265 0 net=1583
rlabel metal2 324 -1265 324 -1265 0 net=2923
rlabel metal2 394 -1265 394 -1265 0 net=6971
rlabel metal2 1003 -1265 1003 -1265 0 net=6703
rlabel metal2 1353 -1265 1353 -1265 0 net=9277
rlabel metal2 170 -1267 170 -1267 0 net=3545
rlabel metal2 345 -1267 345 -1267 0 net=2259
rlabel metal2 429 -1267 429 -1267 0 net=2468
rlabel metal2 555 -1267 555 -1267 0 net=3169
rlabel metal2 870 -1267 870 -1267 0 net=7063
rlabel metal2 1024 -1267 1024 -1267 0 net=7347
rlabel metal2 1143 -1267 1143 -1267 0 net=7941
rlabel metal2 1220 -1267 1220 -1267 0 net=8369
rlabel metal2 170 -1269 170 -1269 0 net=5691
rlabel metal2 877 -1269 877 -1269 0 net=7027
rlabel metal2 282 -1271 282 -1271 0 net=3899
rlabel metal2 996 -1271 996 -1271 0 net=6759
rlabel metal2 1045 -1271 1045 -1271 0 net=8121
rlabel metal2 1171 -1271 1171 -1271 0 net=8683
rlabel metal2 338 -1273 338 -1273 0 net=1833
rlabel metal2 443 -1273 443 -1273 0 net=2825
rlabel metal2 450 -1273 450 -1273 0 net=3785
rlabel metal2 590 -1273 590 -1273 0 net=4249
rlabel metal2 933 -1273 933 -1273 0 net=6573
rlabel metal2 1010 -1273 1010 -1273 0 net=8903
rlabel metal2 1094 -1273 1094 -1273 0 net=7497
rlabel metal2 1199 -1273 1199 -1273 0 net=8245
rlabel metal2 86 -1275 86 -1275 0 net=3823
rlabel metal2 933 -1275 933 -1275 0 net=7422
rlabel metal2 1094 -1275 1094 -1275 0 net=8425
rlabel metal2 1164 -1275 1164 -1275 0 net=7881
rlabel metal2 261 -1277 261 -1277 0 net=1545
rlabel metal2 408 -1277 408 -1277 0 net=1971
rlabel metal2 443 -1277 443 -1277 0 net=3105
rlabel metal2 534 -1277 534 -1277 0 net=2113
rlabel metal2 947 -1277 947 -1277 0 net=6749
rlabel metal2 1048 -1277 1048 -1277 0 net=10188
rlabel metal2 44 -1279 44 -1279 0 net=3739
rlabel metal2 569 -1279 569 -1279 0 net=4413
rlabel metal2 947 -1279 947 -1279 0 net=671
rlabel metal2 44 -1281 44 -1281 0 net=3705
rlabel metal2 226 -1281 226 -1281 0 net=4401
rlabel metal2 954 -1281 954 -1281 0 net=8291
rlabel metal2 1360 -1281 1360 -1281 0 net=9383
rlabel metal2 75 -1283 75 -1283 0 net=2249
rlabel metal2 226 -1283 226 -1283 0 net=1699
rlabel metal2 471 -1283 471 -1283 0 net=2143
rlabel metal2 863 -1283 863 -1283 0 net=5983
rlabel metal2 961 -1283 961 -1283 0 net=7085
rlabel metal2 1101 -1283 1101 -1283 0 net=7635
rlabel metal2 1150 -1283 1150 -1283 0 net=8009
rlabel metal2 1304 -1283 1304 -1283 0 net=9177
rlabel metal2 261 -1285 261 -1285 0 net=1775
rlabel metal2 425 -1285 425 -1285 0 net=8595
rlabel metal2 415 -1287 415 -1287 0 net=4363
rlabel metal2 702 -1287 702 -1287 0 net=6415
rlabel metal2 968 -1287 968 -1287 0 net=7953
rlabel metal2 366 -1289 366 -1289 0 net=6147
rlabel metal2 800 -1289 800 -1289 0 net=5377
rlabel metal2 919 -1289 919 -1289 0 net=6449
rlabel metal2 999 -1289 999 -1289 0 net=1
rlabel metal2 1038 -1289 1038 -1289 0 net=7865
rlabel metal2 1157 -1289 1157 -1289 0 net=8765
rlabel metal2 128 -1291 128 -1291 0 net=5163
rlabel metal2 842 -1291 842 -1291 0 net=5327
rlabel metal2 107 -1293 107 -1293 0 net=4197
rlabel metal2 303 -1293 303 -1293 0 net=3679
rlabel metal2 509 -1293 509 -1293 0 net=4352
rlabel metal2 842 -1293 842 -1293 0 net=6143
rlabel metal2 1052 -1293 1052 -1293 0 net=7447
rlabel metal2 107 -1295 107 -1295 0 net=5707
rlabel metal2 303 -1295 303 -1295 0 net=2241
rlabel metal2 628 -1295 628 -1295 0 net=6817
rlabel metal2 828 -1295 828 -1295 0 net=5321
rlabel metal2 1052 -1295 1052 -1295 0 net=11224
rlabel metal2 114 -1297 114 -1297 0 net=5833
rlabel metal2 632 -1297 632 -1297 0 net=4125
rlabel metal2 849 -1297 849 -1297 0 net=6069
rlabel metal2 1055 -1297 1055 -1297 0 net=9646
rlabel metal2 1507 -1297 1507 -1297 0 net=10705
rlabel metal2 114 -1299 114 -1299 0 net=2551
rlabel metal2 765 -1299 765 -1299 0 net=5273
rlabel metal2 1073 -1299 1073 -1299 0 net=7127
rlabel metal2 1311 -1299 1311 -1299 0 net=9005
rlabel metal2 1458 -1299 1458 -1299 0 net=10229
rlabel metal2 268 -1301 268 -1301 0 net=1611
rlabel metal2 373 -1301 373 -1301 0 net=4083
rlabel metal2 660 -1301 660 -1301 0 net=6881
rlabel metal2 1458 -1301 1458 -1301 0 net=9761
rlabel metal2 51 -1303 51 -1303 0 net=3437
rlabel metal2 373 -1303 373 -1303 0 net=2589
rlabel metal2 660 -1303 660 -1303 0 net=4648
rlabel metal2 765 -1303 765 -1303 0 net=7911
rlabel metal2 51 -1305 51 -1305 0 net=5855
rlabel metal2 730 -1305 730 -1305 0 net=4377
rlabel metal2 786 -1305 786 -1305 0 net=5295
rlabel metal2 257 -1307 257 -1307 0 net=3239
rlabel metal2 481 -1307 481 -1307 0 net=4273
rlabel metal2 786 -1307 786 -1307 0 net=8802
rlabel metal2 891 -1309 891 -1309 0 net=9269
rlabel metal2 891 -1311 891 -1311 0 net=5557
rlabel metal2 1248 -1311 1248 -1311 0 net=9139
rlabel metal2 82 -1313 82 -1313 0 net=6073
rlabel metal2 1269 -1313 1269 -1313 0 net=8717
rlabel metal2 93 -1315 93 -1315 0 net=9159
rlabel metal2 16 -1326 16 -1326 0 net=5857
rlabel metal2 58 -1326 58 -1326 0 net=2122
rlabel metal2 478 -1326 478 -1326 0 net=9278
rlabel metal2 1493 -1326 1493 -1326 0 net=8592
rlabel metal2 1738 -1326 1738 -1326 0 net=8865
rlabel metal2 37 -1328 37 -1328 0 net=3751
rlabel metal2 478 -1328 478 -1328 0 net=2827
rlabel metal2 579 -1328 579 -1328 0 net=8370
rlabel metal2 1346 -1328 1346 -1328 0 net=9270
rlabel metal2 1717 -1328 1717 -1328 0 net=6284
rlabel metal2 37 -1330 37 -1330 0 net=4833
rlabel metal2 233 -1330 233 -1330 0 net=3901
rlabel metal2 289 -1330 289 -1330 0 net=3438
rlabel metal2 597 -1330 597 -1330 0 net=3578
rlabel metal2 768 -1330 768 -1330 0 net=7498
rlabel metal2 1269 -1330 1269 -1330 0 net=9161
rlabel metal2 1269 -1330 1269 -1330 0 net=9161
rlabel metal2 1276 -1330 1276 -1330 0 net=9179
rlabel metal2 1493 -1330 1493 -1330 0 net=12065
rlabel metal2 1556 -1330 1556 -1330 0 net=11167
rlabel metal2 1556 -1330 1556 -1330 0 net=11167
rlabel metal2 1626 -1330 1626 -1330 0 net=11174
rlabel metal2 44 -1332 44 -1332 0 net=3706
rlabel metal2 82 -1332 82 -1332 0 net=8538
rlabel metal2 1521 -1332 1521 -1332 0 net=11111
rlabel metal2 1668 -1332 1668 -1332 0 net=11903
rlabel metal2 1668 -1332 1668 -1332 0 net=11903
rlabel metal2 1675 -1332 1675 -1332 0 net=11939
rlabel metal2 44 -1334 44 -1334 0 net=4673
rlabel metal2 212 -1334 212 -1334 0 net=2545
rlabel metal2 212 -1334 212 -1334 0 net=2545
rlabel metal2 240 -1334 240 -1334 0 net=2070
rlabel metal2 873 -1334 873 -1334 0 net=9628
rlabel metal2 1584 -1334 1584 -1334 0 net=10979
rlabel metal2 1682 -1334 1682 -1334 0 net=11710
rlabel metal2 51 -1336 51 -1336 0 net=3259
rlabel metal2 628 -1336 628 -1336 0 net=4384
rlabel metal2 786 -1336 786 -1336 0 net=6144
rlabel metal2 901 -1336 901 -1336 0 net=8426
rlabel metal2 1125 -1336 1125 -1336 0 net=11651
rlabel metal2 1696 -1336 1696 -1336 0 net=12027
rlabel metal2 75 -1338 75 -1338 0 net=1895
rlabel metal2 250 -1338 250 -1338 0 net=8596
rlabel metal2 1699 -1338 1699 -1338 0 net=10072
rlabel metal2 82 -1340 82 -1340 0 net=7678
rlabel metal2 86 -1342 86 -1342 0 net=2250
rlabel metal2 100 -1342 100 -1342 0 net=1681
rlabel metal2 100 -1342 100 -1342 0 net=1681
rlabel metal2 124 -1342 124 -1342 0 net=2230
rlabel metal2 170 -1342 170 -1342 0 net=5692
rlabel metal2 765 -1342 765 -1342 0 net=9553
rlabel metal2 93 -1344 93 -1344 0 net=7278
rlabel metal2 1283 -1344 1283 -1344 0 net=7129
rlabel metal2 96 -1346 96 -1346 0 net=3546
rlabel metal2 366 -1346 366 -1346 0 net=3680
rlabel metal2 590 -1346 590 -1346 0 net=2365
rlabel metal2 632 -1346 632 -1346 0 net=4085
rlabel metal2 796 -1346 796 -1346 0 net=9543
rlabel metal2 107 -1348 107 -1348 0 net=5709
rlabel metal2 177 -1348 177 -1348 0 net=2058
rlabel metal2 264 -1348 264 -1348 0 net=1584
rlabel metal2 324 -1348 324 -1348 0 net=4513
rlabel metal2 548 -1348 548 -1348 0 net=3081
rlabel metal2 597 -1348 597 -1348 0 net=5328
rlabel metal2 1136 -1348 1136 -1348 0 net=7473
rlabel metal2 107 -1350 107 -1350 0 net=10230
rlabel metal2 135 -1352 135 -1352 0 net=2966
rlabel metal2 460 -1352 460 -1352 0 net=9425
rlabel metal2 135 -1354 135 -1354 0 net=2071
rlabel metal2 506 -1354 506 -1354 0 net=1283
rlabel metal2 653 -1354 653 -1354 0 net=2402
rlabel metal2 821 -1354 821 -1354 0 net=6790
rlabel metal2 1262 -1354 1262 -1354 0 net=9039
rlabel metal2 1339 -1354 1339 -1354 0 net=10687
rlabel metal2 142 -1356 142 -1356 0 net=5303
rlabel metal2 828 -1356 828 -1356 0 net=11476
rlabel metal2 30 -1358 30 -1358 0 net=3819
rlabel metal2 149 -1358 149 -1358 0 net=3513
rlabel metal2 593 -1358 593 -1358 0 net=11721
rlabel metal2 26 -1360 26 -1360 0 net=4989
rlabel metal2 177 -1360 177 -1360 0 net=7093
rlabel metal2 191 -1360 191 -1360 0 net=1669
rlabel metal2 219 -1360 219 -1360 0 net=4387
rlabel metal2 520 -1360 520 -1360 0 net=5559
rlabel metal2 947 -1360 947 -1360 0 net=10956
rlabel metal2 117 -1362 117 -1362 0 net=10923
rlabel metal2 163 -1364 163 -1364 0 net=1501
rlabel metal2 219 -1364 219 -1364 0 net=1938
rlabel metal2 268 -1364 268 -1364 0 net=1613
rlabel metal2 268 -1364 268 -1364 0 net=1613
rlabel metal2 275 -1364 275 -1364 0 net=3786
rlabel metal2 457 -1364 457 -1364 0 net=4275
rlabel metal2 779 -1364 779 -1364 0 net=5231
rlabel metal2 891 -1364 891 -1364 0 net=7466
rlabel metal2 1010 -1364 1010 -1364 0 net=7942
rlabel metal2 1297 -1364 1297 -1364 0 net=9007
rlabel metal2 114 -1366 114 -1366 0 net=2553
rlabel metal2 275 -1366 275 -1366 0 net=2135
rlabel metal2 366 -1366 366 -1366 0 net=2027
rlabel metal2 695 -1366 695 -1366 0 net=3794
rlabel metal2 947 -1366 947 -1366 0 net=6451
rlabel metal2 978 -1366 978 -1366 0 net=11386
rlabel metal2 156 -1368 156 -1368 0 net=1801
rlabel metal2 247 -1368 247 -1368 0 net=9351
rlabel metal2 1612 -1368 1612 -1368 0 net=10523
rlabel metal2 156 -1370 156 -1370 0 net=3447
rlabel metal2 247 -1370 247 -1370 0 net=3999
rlabel metal2 282 -1370 282 -1370 0 net=2261
rlabel metal2 373 -1370 373 -1370 0 net=2591
rlabel metal2 1605 -1370 1605 -1370 0 net=11697
rlabel metal2 289 -1372 289 -1372 0 net=2529
rlabel metal2 436 -1372 436 -1372 0 net=3241
rlabel metal2 548 -1372 548 -1372 0 net=3171
rlabel metal2 562 -1372 562 -1372 0 net=2115
rlabel metal2 614 -1372 614 -1372 0 net=8091
rlabel metal2 828 -1372 828 -1372 0 net=5379
rlabel metal2 968 -1372 968 -1372 0 net=6761
rlabel metal2 1027 -1372 1027 -1372 0 net=11619
rlabel metal2 296 -1374 296 -1374 0 net=1528
rlabel metal2 618 -1374 618 -1374 0 net=3978
rlabel metal2 667 -1374 667 -1374 0 net=6819
rlabel metal2 1045 -1374 1045 -1374 0 net=8123
rlabel metal2 1055 -1374 1055 -1374 0 net=8718
rlabel metal2 1416 -1374 1416 -1374 0 net=11673
rlabel metal2 303 -1376 303 -1376 0 net=2243
rlabel metal2 352 -1376 352 -1376 0 net=2618
rlabel metal2 639 -1376 639 -1376 0 net=4047
rlabel metal2 688 -1376 688 -1376 0 net=9822
rlabel metal2 317 -1378 317 -1378 0 net=1595
rlabel metal2 835 -1378 835 -1378 0 net=5591
rlabel metal2 982 -1378 982 -1378 0 net=9825
rlabel metal2 1479 -1378 1479 -1378 0 net=10363
rlabel metal2 331 -1380 331 -1380 0 net=4723
rlabel metal2 590 -1380 590 -1380 0 net=10789
rlabel metal2 352 -1382 352 -1382 0 net=1973
rlabel metal2 415 -1382 415 -1382 0 net=4365
rlabel metal2 450 -1382 450 -1382 0 net=4807
rlabel metal2 863 -1382 863 -1382 0 net=9376
rlabel metal2 1129 -1382 1129 -1382 0 net=8511
rlabel metal2 1213 -1382 1213 -1382 0 net=8685
rlabel metal2 1304 -1382 1304 -1382 0 net=9325
rlabel metal2 338 -1384 338 -1384 0 net=1546
rlabel metal2 415 -1384 415 -1384 0 net=3740
rlabel metal2 604 -1384 604 -1384 0 net=4477
rlabel metal2 639 -1384 639 -1384 0 net=5296
rlabel metal2 1094 -1384 1094 -1384 0 net=8151
rlabel metal2 1255 -1384 1255 -1384 0 net=9319
rlabel metal2 261 -1386 261 -1386 0 net=1777
rlabel metal2 373 -1386 373 -1386 0 net=3825
rlabel metal2 611 -1386 611 -1386 0 net=9853
rlabel metal2 261 -1388 261 -1388 0 net=7923
rlabel metal2 1146 -1388 1146 -1388 0 net=11884
rlabel metal2 387 -1390 387 -1390 0 net=3041
rlabel metal2 534 -1390 534 -1390 0 net=5323
rlabel metal2 877 -1390 877 -1390 0 net=4250
rlabel metal2 940 -1390 940 -1390 0 net=6407
rlabel metal2 985 -1390 985 -1390 0 net=12080
rlabel metal2 303 -1392 303 -1392 0 net=1507
rlabel metal2 394 -1392 394 -1392 0 net=6973
rlabel metal2 1017 -1392 1017 -1392 0 net=6751
rlabel metal2 1171 -1392 1171 -1392 0 net=8303
rlabel metal2 1311 -1392 1311 -1392 0 net=9619
rlabel metal2 1654 -1392 1654 -1392 0 net=11785
rlabel metal2 205 -1394 205 -1394 0 net=1763
rlabel metal2 401 -1394 401 -1394 0 net=5835
rlabel metal2 877 -1394 877 -1394 0 net=5701
rlabel metal2 905 -1394 905 -1394 0 net=5727
rlabel metal2 1139 -1394 1139 -1394 0 net=8971
rlabel metal2 1325 -1394 1325 -1394 0 net=9797
rlabel metal2 79 -1396 79 -1396 0 net=301
rlabel metal2 940 -1396 940 -1396 0 net=6417
rlabel metal2 1017 -1396 1017 -1396 0 net=7087
rlabel metal2 1069 -1396 1069 -1396 0 net=11716
rlabel metal2 110 -1398 110 -1398 0 net=3701
rlabel metal2 401 -1398 401 -1398 0 net=3107
rlabel metal2 464 -1398 464 -1398 0 net=3895
rlabel metal2 653 -1398 653 -1398 0 net=4207
rlabel metal2 719 -1398 719 -1398 0 net=5984
rlabel metal2 1045 -1398 1045 -1398 0 net=7349
rlabel metal2 1185 -1398 1185 -1398 0 net=9069
rlabel metal2 1332 -1398 1332 -1398 0 net=9289
rlabel metal2 1402 -1398 1402 -1398 0 net=9763
rlabel metal2 1619 -1398 1619 -1398 0 net=11771
rlabel metal2 121 -1400 121 -1400 0 net=9651
rlabel metal2 1458 -1400 1458 -1400 0 net=10217
rlabel metal2 121 -1402 121 -1402 0 net=2177
rlabel metal2 464 -1402 464 -1402 0 net=3981
rlabel metal2 660 -1402 660 -1402 0 net=7028
rlabel metal2 1353 -1402 1353 -1402 0 net=11805
rlabel metal2 128 -1404 128 -1404 0 net=4199
rlabel metal2 660 -1404 660 -1404 0 net=4007
rlabel metal2 1087 -1404 1087 -1404 0 net=7867
rlabel metal2 1185 -1404 1185 -1404 0 net=9195
rlabel metal2 1486 -1404 1486 -1404 0 net=10443
rlabel metal2 128 -1406 128 -1406 0 net=2925
rlabel metal2 380 -1406 380 -1406 0 net=1835
rlabel metal2 485 -1406 485 -1406 0 net=2456
rlabel metal2 730 -1406 730 -1406 0 net=11557
rlabel metal2 23 -1408 23 -1408 0 net=3969
rlabel metal2 499 -1408 499 -1408 0 net=11683
rlabel metal2 65 -1410 65 -1410 0 net=1541
rlabel metal2 513 -1410 513 -1410 0 net=2859
rlabel metal2 1206 -1410 1206 -1410 0 net=8751
rlabel metal2 1353 -1410 1353 -1410 0 net=9477
rlabel metal2 1528 -1410 1528 -1410 0 net=10811
rlabel metal2 65 -1412 65 -1412 0 net=2001
rlabel metal2 226 -1412 226 -1412 0 net=1701
rlabel metal2 555 -1412 555 -1412 0 net=10211
rlabel metal2 310 -1414 310 -1414 0 net=1807
rlabel metal2 583 -1414 583 -1414 0 net=6177
rlabel metal2 1157 -1414 1157 -1414 0 net=8767
rlabel metal2 310 -1416 310 -1416 0 net=2145
rlabel metal2 677 -1416 677 -1416 0 net=8841
rlabel metal2 1248 -1416 1248 -1416 0 net=9141
rlabel metal2 58 -1418 58 -1418 0 net=3335
rlabel metal2 688 -1418 688 -1418 0 net=4127
rlabel metal2 709 -1418 709 -1418 0 net=4255
rlabel metal2 723 -1418 723 -1418 0 net=4138
rlabel metal2 800 -1418 800 -1418 0 net=5165
rlabel metal2 1248 -1418 1248 -1418 0 net=8613
rlabel metal2 695 -1420 695 -1420 0 net=4415
rlabel metal2 800 -1420 800 -1420 0 net=5275
rlabel metal2 866 -1420 866 -1420 0 net=11253
rlabel metal2 702 -1422 702 -1422 0 net=6865
rlabel metal2 1395 -1422 1395 -1422 0 net=9755
rlabel metal2 61 -1424 61 -1424 0 net=7249
rlabel metal2 1430 -1424 1430 -1424 0 net=9385
rlabel metal2 716 -1426 716 -1426 0 net=8239
rlabel metal2 1430 -1426 1430 -1426 0 net=9933
rlabel metal2 226 -1428 226 -1428 0 net=10293
rlabel metal2 723 -1430 723 -1430 0 net=8210
rlabel metal2 744 -1432 744 -1432 0 net=5551
rlabel metal2 814 -1432 814 -1432 0 net=6361
rlabel metal2 919 -1432 919 -1432 0 net=6071
rlabel metal2 975 -1432 975 -1432 0 net=6575
rlabel metal2 1367 -1432 1367 -1432 0 net=10197
rlabel metal2 737 -1434 737 -1434 0 net=4379
rlabel metal2 751 -1434 751 -1434 0 net=4905
rlabel metal2 814 -1434 814 -1434 0 net=7223
rlabel metal2 919 -1434 919 -1434 0 net=7037
rlabel metal2 1472 -1434 1472 -1434 0 net=10313
rlabel metal2 145 -1436 145 -1436 0 net=4591
rlabel metal2 758 -1436 758 -1436 0 net=7065
rlabel metal2 933 -1436 933 -1436 0 net=9981
rlabel metal2 1500 -1436 1500 -1436 0 net=10667
rlabel metal2 569 -1438 569 -1438 0 net=4403
rlabel metal2 824 -1438 824 -1438 0 net=9989
rlabel metal2 1535 -1438 1535 -1438 0 net=10875
rlabel metal2 509 -1440 509 -1440 0 net=3845
rlabel metal2 681 -1440 681 -1440 0 net=6149
rlabel metal2 933 -1440 933 -1440 0 net=11803
rlabel metal2 674 -1442 674 -1442 0 net=4113
rlabel metal2 849 -1442 849 -1442 0 net=6075
rlabel metal2 954 -1442 954 -1442 0 net=7637
rlabel metal2 1577 -1442 1577 -1442 0 net=11523
rlabel metal2 492 -1444 492 -1444 0 net=4694
rlabel metal2 856 -1444 856 -1444 0 net=6113
rlabel metal2 926 -1444 926 -1444 0 net=6705
rlabel metal2 1059 -1444 1059 -1444 0 net=7449
rlabel metal2 1143 -1444 1143 -1444 0 net=9387
rlabel metal2 1563 -1444 1563 -1444 0 net=10707
rlabel metal2 86 -1446 86 -1446 0 net=2719
rlabel metal2 1227 -1446 1227 -1446 0 net=8247
rlabel metal2 93 -1448 93 -1448 0 net=11205
rlabel metal2 530 -1448 530 -1448 0 net=10027
rlabel metal2 996 -1450 996 -1450 0 net=6883
rlabel metal2 1003 -1452 1003 -1452 0 net=8011
rlabel metal2 600 -1454 600 -1454 0 net=11343
rlabel metal2 1038 -1456 1038 -1456 0 net=7353
rlabel metal2 1115 -1458 1115 -1458 0 net=7883
rlabel metal2 1164 -1460 1164 -1460 0 net=8293
rlabel metal2 1080 -1462 1080 -1462 0 net=8905
rlabel metal2 1080 -1464 1080 -1464 0 net=7955
rlabel metal2 1052 -1466 1052 -1466 0 net=8469
rlabel metal2 912 -1468 912 -1468 0 net=7913
rlabel metal2 642 -1470 642 -1470 0 net=6019
rlabel metal2 16 -1481 16 -1481 0 net=5858
rlabel metal2 786 -1481 786 -1481 0 net=4086
rlabel metal2 870 -1481 870 -1481 0 net=7038
rlabel metal2 1024 -1481 1024 -1481 0 net=8152
rlabel metal2 1104 -1481 1104 -1481 0 net=10688
rlabel metal2 1745 -1481 1745 -1481 0 net=8867
rlabel metal2 23 -1483 23 -1483 0 net=4977
rlabel metal2 96 -1483 96 -1483 0 net=11722
rlabel metal2 30 -1485 30 -1485 0 net=4990
rlabel metal2 100 -1485 100 -1485 0 net=1683
rlabel metal2 100 -1485 100 -1485 0 net=1683
rlabel metal2 107 -1485 107 -1485 0 net=660
rlabel metal2 418 -1485 418 -1485 0 net=5317
rlabel metal2 786 -1485 786 -1485 0 net=6363
rlabel metal2 1024 -1485 1024 -1485 0 net=7869
rlabel metal2 1118 -1485 1118 -1485 0 net=12028
rlabel metal2 58 -1487 58 -1487 0 net=10212
rlabel metal2 61 -1489 61 -1489 0 net=668
rlabel metal2 142 -1489 142 -1489 0 net=3820
rlabel metal2 226 -1489 226 -1489 0 net=1808
rlabel metal2 373 -1489 373 -1489 0 net=3826
rlabel metal2 863 -1489 863 -1489 0 net=6419
rlabel metal2 1073 -1489 1073 -1489 0 net=5728
rlabel metal2 68 -1491 68 -1491 0 net=3172
rlabel metal2 555 -1491 555 -1491 0 net=1373
rlabel metal2 621 -1491 621 -1491 0 net=4256
rlabel metal2 719 -1491 719 -1491 0 net=8248
rlabel metal2 1640 -1491 1640 -1491 0 net=11905
rlabel metal2 72 -1493 72 -1493 0 net=2028
rlabel metal2 390 -1493 390 -1493 0 net=1542
rlabel metal2 443 -1493 443 -1493 0 net=1702
rlabel metal2 562 -1493 562 -1493 0 net=2116
rlabel metal2 733 -1493 733 -1493 0 net=6753
rlabel metal2 1073 -1493 1073 -1493 0 net=8253
rlabel metal2 1153 -1493 1153 -1493 0 net=9290
rlabel metal2 1339 -1493 1339 -1493 0 net=9827
rlabel metal2 1493 -1493 1493 -1493 0 net=12067
rlabel metal2 44 -1495 44 -1495 0 net=4675
rlabel metal2 107 -1495 107 -1495 0 net=2493
rlabel metal2 394 -1495 394 -1495 0 net=1764
rlabel metal2 866 -1495 866 -1495 0 net=8581
rlabel metal2 1122 -1495 1122 -1495 0 net=9040
rlabel metal2 1311 -1495 1311 -1495 0 net=9621
rlabel metal2 1416 -1495 1416 -1495 0 net=10445
rlabel metal2 1493 -1495 1493 -1495 0 net=10877
rlabel metal2 1563 -1495 1563 -1495 0 net=11653
rlabel metal2 1612 -1495 1612 -1495 0 net=10525
rlabel metal2 44 -1497 44 -1497 0 net=2557
rlabel metal2 394 -1497 394 -1497 0 net=3337
rlabel metal2 474 -1497 474 -1497 0 net=6072
rlabel metal2 989 -1497 989 -1497 0 net=6821
rlabel metal2 1125 -1497 1125 -1497 0 net=11940
rlabel metal2 30 -1499 30 -1499 0 net=4695
rlabel metal2 492 -1499 492 -1499 0 net=11206
rlabel metal2 905 -1499 905 -1499 0 net=6707
rlabel metal2 961 -1499 961 -1499 0 net=6763
rlabel metal2 975 -1499 975 -1499 0 net=6577
rlabel metal2 1087 -1499 1087 -1499 0 net=8305
rlabel metal2 1311 -1499 1311 -1499 0 net=9389
rlabel metal2 1486 -1499 1486 -1499 0 net=11675
rlabel metal2 114 -1501 114 -1501 0 net=4366
rlabel metal2 443 -1501 443 -1501 0 net=5759
rlabel metal2 114 -1503 114 -1503 0 net=4421
rlabel metal2 677 -1503 677 -1503 0 net=11558
rlabel metal2 1556 -1503 1556 -1503 0 net=11169
rlabel metal2 142 -1505 142 -1505 0 net=3109
rlabel metal2 408 -1505 408 -1505 0 net=4541
rlabel metal2 408 -1505 408 -1505 0 net=4541
rlabel metal2 422 -1505 422 -1505 0 net=3752
rlabel metal2 607 -1505 607 -1505 0 net=4048
rlabel metal2 730 -1505 730 -1505 0 net=9217
rlabel metal2 1325 -1505 1325 -1505 0 net=9765
rlabel metal2 1500 -1505 1500 -1505 0 net=10669
rlabel metal2 51 -1507 51 -1507 0 net=3261
rlabel metal2 436 -1507 436 -1507 0 net=2251
rlabel metal2 975 -1507 975 -1507 0 net=9427
rlabel metal2 1402 -1507 1402 -1507 0 net=10315
rlabel metal2 1535 -1507 1535 -1507 0 net=11525
rlabel metal2 1584 -1507 1584 -1507 0 net=11621
rlabel metal2 156 -1509 156 -1509 0 net=11147
rlabel metal2 1570 -1509 1570 -1509 0 net=11255
rlabel metal2 1584 -1509 1584 -1509 0 net=10709
rlabel metal2 156 -1511 156 -1511 0 net=2547
rlabel metal2 226 -1511 226 -1511 0 net=3931
rlabel metal2 261 -1511 261 -1511 0 net=2263
rlabel metal2 296 -1511 296 -1511 0 net=3897
rlabel metal2 632 -1511 632 -1511 0 net=7350
rlabel metal2 1048 -1511 1048 -1511 0 net=11595
rlabel metal2 1598 -1511 1598 -1511 0 net=11685
rlabel metal2 159 -1513 159 -1513 0 net=6178
rlabel metal2 635 -1513 635 -1513 0 net=2592
rlabel metal2 1549 -1513 1549 -1513 0 net=11543
rlabel metal2 149 -1515 149 -1515 0 net=3515
rlabel metal2 639 -1515 639 -1515 0 net=1002
rlabel metal2 149 -1517 149 -1517 0 net=1633
rlabel metal2 562 -1517 562 -1517 0 net=4114
rlabel metal2 712 -1517 712 -1517 0 net=11249
rlabel metal2 1619 -1517 1619 -1517 0 net=11699
rlabel metal2 191 -1519 191 -1519 0 net=3448
rlabel metal2 229 -1519 229 -1519 0 net=6408
rlabel metal2 1045 -1519 1045 -1519 0 net=5166
rlabel metal2 1139 -1519 1139 -1519 0 net=9386
rlabel metal2 1472 -1519 1472 -1519 0 net=11787
rlabel metal2 194 -1521 194 -1521 0 net=5324
rlabel metal2 541 -1521 541 -1521 0 net=3243
rlabel metal2 576 -1521 576 -1521 0 net=3082
rlabel metal2 604 -1521 604 -1521 0 net=4479
rlabel metal2 730 -1521 730 -1521 0 net=5233
rlabel metal2 796 -1521 796 -1521 0 net=10887
rlabel metal2 79 -1523 79 -1523 0 net=2383
rlabel metal2 604 -1523 604 -1523 0 net=11804
rlabel metal2 79 -1525 79 -1525 0 net=1803
rlabel metal2 198 -1525 198 -1525 0 net=1671
rlabel metal2 198 -1525 198 -1525 0 net=1671
rlabel metal2 212 -1525 212 -1525 0 net=1897
rlabel metal2 268 -1525 268 -1525 0 net=1615
rlabel metal2 310 -1525 310 -1525 0 net=2147
rlabel metal2 450 -1525 450 -1525 0 net=4808
rlabel metal2 499 -1525 499 -1525 0 net=4583
rlabel metal2 639 -1525 639 -1525 0 net=4009
rlabel metal2 747 -1525 747 -1525 0 net=7224
rlabel metal2 870 -1525 870 -1525 0 net=7089
rlabel metal2 1020 -1525 1020 -1525 0 net=11985
rlabel metal2 121 -1527 121 -1527 0 net=2179
rlabel metal2 299 -1527 299 -1527 0 net=1585
rlabel metal2 331 -1527 331 -1527 0 net=4725
rlabel metal2 450 -1527 450 -1527 0 net=2367
rlabel metal2 779 -1527 779 -1527 0 net=5277
rlabel metal2 891 -1527 891 -1527 0 net=8739
rlabel metal2 1143 -1527 1143 -1527 0 net=8753
rlabel metal2 1283 -1527 1283 -1527 0 net=9071
rlabel metal2 93 -1529 93 -1529 0 net=2941
rlabel metal2 163 -1529 163 -1529 0 net=1793
rlabel metal2 646 -1529 646 -1529 0 net=4201
rlabel metal2 646 -1529 646 -1529 0 net=4201
rlabel metal2 653 -1529 653 -1529 0 net=4209
rlabel metal2 653 -1529 653 -1529 0 net=4209
rlabel metal2 660 -1529 660 -1529 0 net=4417
rlabel metal2 719 -1529 719 -1529 0 net=9657
rlabel metal2 1346 -1529 1346 -1529 0 net=9855
rlabel metal2 1451 -1529 1451 -1529 0 net=10925
rlabel metal2 93 -1531 93 -1531 0 net=2366
rlabel metal2 674 -1531 674 -1531 0 net=4405
rlabel metal2 793 -1531 793 -1531 0 net=5553
rlabel metal2 891 -1531 891 -1531 0 net=6885
rlabel metal2 1017 -1531 1017 -1531 0 net=7130
rlabel metal2 51 -1533 51 -1533 0 net=8435
rlabel metal2 800 -1533 800 -1533 0 net=5837
rlabel metal2 898 -1533 898 -1533 0 net=6453
rlabel metal2 982 -1533 982 -1533 0 net=8241
rlabel metal2 1171 -1533 1171 -1533 0 net=8907
rlabel metal2 1258 -1533 1258 -1533 0 net=10649
rlabel metal2 1521 -1533 1521 -1533 0 net=11113
rlabel metal2 1626 -1533 1626 -1533 0 net=10981
rlabel metal2 205 -1535 205 -1535 0 net=3703
rlabel metal2 338 -1535 338 -1535 0 net=1779
rlabel metal2 464 -1535 464 -1535 0 net=3983
rlabel metal2 737 -1535 737 -1535 0 net=8111
rlabel metal2 996 -1535 996 -1535 0 net=7451
rlabel metal2 1062 -1535 1062 -1535 0 net=8769
rlabel metal2 1199 -1535 1199 -1535 0 net=11345
rlabel metal2 1521 -1535 1521 -1535 0 net=11807
rlabel metal2 191 -1537 191 -1537 0 net=9505
rlabel metal2 1206 -1537 1206 -1537 0 net=9545
rlabel metal2 1661 -1537 1661 -1537 0 net=11735
rlabel metal2 205 -1539 205 -1539 0 net=6020
rlabel metal2 926 -1539 926 -1539 0 net=8768
rlabel metal2 219 -1541 219 -1541 0 net=4001
rlabel metal2 303 -1541 303 -1541 0 net=1509
rlabel metal2 502 -1541 502 -1541 0 net=4128
rlabel metal2 758 -1541 758 -1541 0 net=7067
rlabel metal2 933 -1541 933 -1541 0 net=11825
rlabel metal2 184 -1543 184 -1543 0 net=1503
rlabel metal2 324 -1543 324 -1543 0 net=4515
rlabel metal2 758 -1543 758 -1543 0 net=9196
rlabel metal2 1227 -1543 1227 -1543 0 net=10029
rlabel metal2 135 -1545 135 -1545 0 net=2073
rlabel metal2 233 -1545 233 -1545 0 net=3903
rlabel metal2 338 -1545 338 -1545 0 net=6949
rlabel metal2 506 -1545 506 -1545 0 net=4388
rlabel metal2 842 -1545 842 -1545 0 net=5117
rlabel metal2 1129 -1545 1129 -1545 0 net=8687
rlabel metal2 1227 -1545 1227 -1545 0 net=7475
rlabel metal2 37 -1547 37 -1547 0 net=4835
rlabel metal2 233 -1547 233 -1547 0 net=7799
rlabel metal2 457 -1547 457 -1547 0 net=4277
rlabel metal2 513 -1547 513 -1547 0 net=2861
rlabel metal2 513 -1547 513 -1547 0 net=2861
rlabel metal2 520 -1547 520 -1547 0 net=5560
rlabel metal2 1185 -1547 1185 -1547 0 net=8973
rlabel metal2 1290 -1547 1290 -1547 0 net=9009
rlabel metal2 86 -1549 86 -1549 0 net=2721
rlabel metal2 457 -1549 457 -1549 0 net=3971
rlabel metal2 527 -1549 527 -1549 0 net=3043
rlabel metal2 569 -1549 569 -1549 0 net=3847
rlabel metal2 625 -1549 625 -1549 0 net=3381
rlabel metal2 933 -1549 933 -1549 0 net=8981
rlabel metal2 947 -1549 947 -1549 0 net=7251
rlabel metal2 1213 -1549 1213 -1549 0 net=9479
rlabel metal2 65 -1551 65 -1551 0 net=2003
rlabel metal2 590 -1551 590 -1551 0 net=5305
rlabel metal2 1031 -1551 1031 -1551 0 net=7885
rlabel metal2 1234 -1551 1234 -1551 0 net=9321
rlabel metal2 1297 -1551 1297 -1551 0 net=9757
rlabel metal2 65 -1553 65 -1553 0 net=7499
rlabel metal2 1241 -1553 1241 -1553 0 net=9353
rlabel metal2 1353 -1553 1353 -1553 0 net=9983
rlabel metal2 86 -1555 86 -1555 0 net=5593
rlabel metal2 873 -1555 873 -1555 0 net=1128
rlabel metal2 1318 -1555 1318 -1555 0 net=9555
rlabel metal2 1437 -1555 1437 -1555 0 net=10813
rlabel metal2 128 -1557 128 -1557 0 net=2927
rlabel metal2 527 -1557 527 -1557 0 net=513
rlabel metal2 128 -1559 128 -1559 0 net=2137
rlabel metal2 345 -1559 345 -1559 0 net=2245
rlabel metal2 485 -1559 485 -1559 0 net=4593
rlabel metal2 807 -1559 807 -1559 0 net=12069
rlabel metal2 170 -1561 170 -1561 0 net=5711
rlabel metal2 1115 -1561 1115 -1561 0 net=11485
rlabel metal2 170 -1563 170 -1563 0 net=1975
rlabel metal2 359 -1563 359 -1563 0 net=2829
rlabel metal2 667 -1563 667 -1563 0 net=10297
rlabel metal2 1367 -1563 1367 -1563 0 net=10199
rlabel metal2 254 -1565 254 -1565 0 net=2555
rlabel metal2 352 -1565 352 -1565 0 net=1837
rlabel metal2 478 -1565 478 -1565 0 net=5381
rlabel metal2 1367 -1565 1367 -1565 0 net=9991
rlabel metal2 275 -1567 275 -1567 0 net=1597
rlabel metal2 380 -1567 380 -1567 0 net=17
rlabel metal2 751 -1567 751 -1567 0 net=4907
rlabel metal2 821 -1567 821 -1567 0 net=8093
rlabel metal2 1430 -1567 1430 -1567 0 net=9935
rlabel metal2 289 -1569 289 -1569 0 net=2531
rlabel metal2 688 -1569 688 -1569 0 net=6975
rlabel metal2 1430 -1569 1430 -1569 0 net=10295
rlabel metal2 177 -1571 177 -1571 0 net=7094
rlabel metal2 614 -1571 614 -1571 0 net=11143
rlabel metal2 177 -1573 177 -1573 0 net=8815
rlabel metal2 716 -1573 716 -1573 0 net=6752
rlabel metal2 723 -1575 723 -1575 0 net=8629
rlabel metal2 723 -1577 723 -1577 0 net=4380
rlabel metal2 772 -1577 772 -1577 0 net=6115
rlabel metal2 1010 -1577 1010 -1577 0 net=7915
rlabel metal2 1108 -1577 1108 -1577 0 net=8513
rlabel metal2 548 -1579 548 -1579 0 net=3121
rlabel metal2 821 -1579 821 -1579 0 net=8295
rlabel metal2 1192 -1579 1192 -1579 0 net=9163
rlabel metal2 614 -1581 614 -1581 0 net=9461
rlabel metal2 726 -1583 726 -1583 0 net=7638
rlabel metal2 1052 -1583 1052 -1583 0 net=7957
rlabel metal2 1164 -1583 1164 -1583 0 net=8843
rlabel metal2 828 -1585 828 -1585 0 net=5703
rlabel metal2 954 -1585 954 -1585 0 net=7925
rlabel metal2 1220 -1585 1220 -1585 0 net=8615
rlabel metal2 849 -1587 849 -1587 0 net=6077
rlabel metal2 877 -1587 877 -1587 0 net=6151
rlabel metal2 1080 -1587 1080 -1587 0 net=8125
rlabel metal2 1248 -1587 1248 -1587 0 net=9327
rlabel metal2 702 -1589 702 -1589 0 net=6867
rlabel metal2 1101 -1589 1101 -1589 0 net=9142
rlabel metal2 292 -1591 292 -1591 0 net=5745
rlabel metal2 849 -1591 849 -1591 0 net=8013
rlabel metal2 1304 -1591 1304 -1591 0 net=9799
rlabel metal2 541 -1593 541 -1593 0 net=10345
rlabel metal2 1003 -1595 1003 -1595 0 net=7355
rlabel metal2 1381 -1595 1381 -1595 0 net=10219
rlabel metal2 1038 -1597 1038 -1597 0 net=8471
rlabel metal2 1458 -1597 1458 -1597 0 net=10365
rlabel metal2 1178 -1599 1178 -1599 0 net=9181
rlabel metal2 1479 -1599 1479 -1599 0 net=11773
rlabel metal2 264 -1601 264 -1601 0 net=11919
rlabel metal2 1276 -1603 1276 -1603 0 net=9653
rlabel metal2 1388 -1605 1388 -1605 0 net=10791
rlabel metal2 642 -1607 642 -1607 0 net=11431
rlabel metal2 16 -1618 16 -1618 0 net=4696
rlabel metal2 37 -1618 37 -1618 0 net=8807
rlabel metal2 296 -1618 296 -1618 0 net=3898
rlabel metal2 411 -1618 411 -1618 0 net=4567
rlabel metal2 758 -1618 758 -1618 0 net=1074
rlabel metal2 1115 -1618 1115 -1618 0 net=9556
rlabel metal2 1381 -1618 1381 -1618 0 net=10221
rlabel metal2 1479 -1618 1479 -1618 0 net=11775
rlabel metal2 1752 -1618 1752 -1618 0 net=8869
rlabel metal2 44 -1620 44 -1620 0 net=2558
rlabel metal2 268 -1620 268 -1620 0 net=1586
rlabel metal2 317 -1620 317 -1620 0 net=6185
rlabel metal2 929 -1620 929 -1620 0 net=9072
rlabel metal2 1717 -1620 1717 -1620 0 net=8631
rlabel metal2 44 -1622 44 -1622 0 net=2533
rlabel metal2 348 -1622 348 -1622 0 net=6754
rlabel metal2 933 -1622 933 -1622 0 net=8983
rlabel metal2 933 -1622 933 -1622 0 net=8983
rlabel metal2 961 -1622 961 -1622 0 net=6765
rlabel metal2 961 -1622 961 -1622 0 net=6765
rlabel metal2 996 -1622 996 -1622 0 net=7453
rlabel metal2 58 -1624 58 -1624 0 net=11114
rlabel metal2 1626 -1624 1626 -1624 0 net=11827
rlabel metal2 65 -1626 65 -1626 0 net=4991
rlabel metal2 513 -1626 513 -1626 0 net=2862
rlabel metal2 730 -1626 730 -1626 0 net=5235
rlabel metal2 761 -1626 761 -1626 0 net=11736
rlabel metal2 1668 -1626 1668 -1626 0 net=10526
rlabel metal2 72 -1628 72 -1628 0 net=4677
rlabel metal2 72 -1628 72 -1628 0 net=4677
rlabel metal2 79 -1628 79 -1628 0 net=1804
rlabel metal2 268 -1628 268 -1628 0 net=2041
rlabel metal2 324 -1628 324 -1628 0 net=2556
rlabel metal2 369 -1628 369 -1628 0 net=2148
rlabel metal2 432 -1628 432 -1628 0 net=3972
rlabel metal2 478 -1628 478 -1628 0 net=5382
rlabel metal2 632 -1628 632 -1628 0 net=3985
rlabel metal2 632 -1628 632 -1628 0 net=3985
rlabel metal2 639 -1628 639 -1628 0 net=4011
rlabel metal2 639 -1628 639 -1628 0 net=4011
rlabel metal2 667 -1628 667 -1628 0 net=5554
rlabel metal2 828 -1628 828 -1628 0 net=5704
rlabel metal2 919 -1628 919 -1628 0 net=342
rlabel metal2 975 -1628 975 -1628 0 net=9429
rlabel metal2 23 -1630 23 -1630 0 net=4979
rlabel metal2 373 -1630 373 -1630 0 net=1781
rlabel metal2 373 -1630 373 -1630 0 net=1781
rlabel metal2 387 -1630 387 -1630 0 net=2723
rlabel metal2 513 -1630 513 -1630 0 net=3353
rlabel metal2 667 -1630 667 -1630 0 net=4517
rlabel metal2 712 -1630 712 -1630 0 net=7870
rlabel metal2 1048 -1630 1048 -1630 0 net=10670
rlabel metal2 1640 -1630 1640 -1630 0 net=11907
rlabel metal2 61 -1632 61 -1632 0 net=6223
rlabel metal2 450 -1632 450 -1632 0 net=2368
rlabel metal2 793 -1632 793 -1632 0 net=8094
rlabel metal2 1486 -1632 1486 -1632 0 net=11677
rlabel metal2 79 -1634 79 -1634 0 net=3123
rlabel metal2 562 -1634 562 -1634 0 net=9271
rlabel metal2 1381 -1634 1381 -1634 0 net=10317
rlabel metal2 1500 -1634 1500 -1634 0 net=11251
rlabel metal2 1640 -1634 1640 -1634 0 net=10983
rlabel metal2 121 -1636 121 -1636 0 net=2942
rlabel metal2 548 -1636 548 -1636 0 net=3245
rlabel metal2 576 -1636 576 -1636 0 net=2384
rlabel metal2 975 -1636 975 -1636 0 net=10366
rlabel metal2 1514 -1636 1514 -1636 0 net=11433
rlabel metal2 121 -1638 121 -1638 0 net=4025
rlabel metal2 726 -1638 726 -1638 0 net=6454
rlabel metal2 996 -1638 996 -1638 0 net=8473
rlabel metal2 1059 -1638 1059 -1638 0 net=9936
rlabel metal2 1521 -1638 1521 -1638 0 net=11809
rlabel metal2 135 -1640 135 -1640 0 net=4836
rlabel metal2 674 -1640 674 -1640 0 net=4406
rlabel metal2 803 -1640 803 -1640 0 net=6379
rlabel metal2 863 -1640 863 -1640 0 net=6421
rlabel metal2 1115 -1640 1115 -1640 0 net=10073
rlabel metal2 1591 -1640 1591 -1640 0 net=11623
rlabel metal2 135 -1642 135 -1642 0 net=4481
rlabel metal2 702 -1642 702 -1642 0 net=5747
rlabel metal2 807 -1642 807 -1642 0 net=7543
rlabel metal2 1118 -1642 1118 -1642 0 net=9322
rlabel metal2 1241 -1642 1241 -1642 0 net=9355
rlabel metal2 1598 -1642 1598 -1642 0 net=11687
rlabel metal2 156 -1644 156 -1644 0 net=2549
rlabel metal2 450 -1644 450 -1644 0 net=2381
rlabel metal2 807 -1644 807 -1644 0 net=6811
rlabel metal2 992 -1644 992 -1644 0 net=11195
rlabel metal2 1647 -1644 1647 -1644 0 net=11921
rlabel metal2 156 -1646 156 -1646 0 net=8242
rlabel metal2 1003 -1646 1003 -1646 0 net=7357
rlabel metal2 1003 -1646 1003 -1646 0 net=7357
rlabel metal2 1052 -1646 1052 -1646 0 net=7959
rlabel metal2 1251 -1646 1251 -1646 0 net=12068
rlabel metal2 170 -1648 170 -1648 0 net=1977
rlabel metal2 338 -1648 338 -1648 0 net=6951
rlabel metal2 733 -1648 733 -1648 0 net=8112
rlabel metal2 982 -1648 982 -1648 0 net=6959
rlabel metal2 1101 -1648 1101 -1648 0 net=11387
rlabel metal2 1654 -1648 1654 -1648 0 net=11987
rlabel metal2 170 -1650 170 -1650 0 net=3704
rlabel metal2 338 -1650 338 -1650 0 net=4203
rlabel metal2 709 -1650 709 -1650 0 net=7719
rlabel metal2 1101 -1650 1101 -1650 0 net=8909
rlabel metal2 1213 -1650 1213 -1650 0 net=9481
rlabel metal2 1689 -1650 1689 -1650 0 net=10771
rlabel metal2 191 -1652 191 -1652 0 net=370
rlabel metal2 289 -1652 289 -1652 0 net=8015
rlabel metal2 863 -1652 863 -1652 0 net=6869
rlabel metal2 887 -1652 887 -1652 0 net=10296
rlabel metal2 1437 -1652 1437 -1652 0 net=10815
rlabel metal2 1619 -1652 1619 -1652 0 net=11701
rlabel metal2 191 -1654 191 -1654 0 net=7090
rlabel metal2 968 -1654 968 -1654 0 net=6579
rlabel metal2 1010 -1654 1010 -1654 0 net=7917
rlabel metal2 1153 -1654 1153 -1654 0 net=9622
rlabel metal2 1367 -1654 1367 -1654 0 net=9993
rlabel metal2 1465 -1654 1465 -1654 0 net=11145
rlabel metal2 194 -1656 194 -1656 0 net=11148
rlabel metal2 205 -1658 205 -1658 0 net=9073
rlabel metal2 1255 -1658 1255 -1658 0 net=11788
rlabel metal2 1493 -1658 1493 -1658 0 net=10879
rlabel metal2 51 -1660 51 -1660 0 net=8437
rlabel metal2 208 -1660 208 -1660 0 net=12070
rlabel metal2 51 -1662 51 -1662 0 net=4543
rlabel metal2 422 -1662 422 -1662 0 net=4727
rlabel metal2 737 -1662 737 -1662 0 net=11170
rlabel metal2 177 -1664 177 -1664 0 net=8817
rlabel metal2 1262 -1664 1262 -1664 0 net=9219
rlabel metal2 1507 -1664 1507 -1664 0 net=11347
rlabel metal2 212 -1666 212 -1666 0 net=1899
rlabel metal2 331 -1666 331 -1666 0 net=2669
rlabel metal2 1066 -1666 1066 -1666 0 net=10299
rlabel metal2 1563 -1666 1563 -1666 0 net=11655
rlabel metal2 86 -1668 86 -1668 0 net=5595
rlabel metal2 226 -1668 226 -1668 0 net=3933
rlabel metal2 597 -1668 597 -1668 0 net=3849
rlabel metal2 604 -1668 604 -1668 0 net=6822
rlabel metal2 1206 -1668 1206 -1668 0 net=9547
rlabel metal2 1367 -1668 1367 -1668 0 net=11545
rlabel metal2 1563 -1668 1563 -1668 0 net=11057
rlabel metal2 86 -1670 86 -1670 0 net=3111
rlabel metal2 184 -1670 184 -1670 0 net=2075
rlabel metal2 233 -1670 233 -1670 0 net=7801
rlabel metal2 1066 -1670 1066 -1670 0 net=10545
rlabel metal2 1535 -1670 1535 -1670 0 net=11527
rlabel metal2 1584 -1670 1584 -1670 0 net=10711
rlabel metal2 142 -1672 142 -1672 0 net=1795
rlabel metal2 184 -1672 184 -1672 0 net=1673
rlabel metal2 233 -1672 233 -1672 0 net=2265
rlabel metal2 278 -1672 278 -1672 0 net=7423
rlabel metal2 1073 -1672 1073 -1672 0 net=8255
rlabel metal2 1157 -1672 1157 -1672 0 net=8771
rlabel metal2 1220 -1672 1220 -1672 0 net=8617
rlabel metal2 1220 -1672 1220 -1672 0 net=8617
rlabel metal2 1269 -1672 1269 -1672 0 net=9463
rlabel metal2 107 -1674 107 -1674 0 net=2495
rlabel metal2 240 -1674 240 -1674 0 net=2181
rlabel metal2 436 -1674 436 -1674 0 net=2252
rlabel metal2 1073 -1674 1073 -1674 0 net=7477
rlabel metal2 1276 -1674 1276 -1674 0 net=9655
rlabel metal2 100 -1676 100 -1676 0 net=1685
rlabel metal2 149 -1676 149 -1676 0 net=1635
rlabel metal2 240 -1676 240 -1676 0 net=1617
rlabel metal2 296 -1676 296 -1676 0 net=2247
rlabel metal2 436 -1676 436 -1676 0 net=4419
rlabel metal2 772 -1676 772 -1676 0 net=6117
rlabel metal2 870 -1676 870 -1676 0 net=6152
rlabel metal2 905 -1676 905 -1676 0 net=6709
rlabel metal2 1304 -1676 1304 -1676 0 net=9801
rlabel metal2 1416 -1676 1416 -1676 0 net=10447
rlabel metal2 100 -1678 100 -1678 0 net=2029
rlabel metal2 478 -1678 478 -1678 0 net=5581
rlabel metal2 751 -1678 751 -1678 0 net=4909
rlabel metal2 782 -1678 782 -1678 0 net=11097
rlabel metal2 149 -1680 149 -1680 0 net=7755
rlabel metal2 751 -1680 751 -1680 0 net=5119
rlabel metal2 877 -1680 877 -1680 0 net=6887
rlabel metal2 905 -1680 905 -1680 0 net=7927
rlabel metal2 1020 -1680 1020 -1680 0 net=9111
rlabel metal2 1339 -1680 1339 -1680 0 net=9829
rlabel metal2 1423 -1680 1423 -1680 0 net=10651
rlabel metal2 282 -1682 282 -1682 0 net=1511
rlabel metal2 492 -1682 492 -1682 0 net=10779
rlabel metal2 359 -1684 359 -1684 0 net=2831
rlabel metal2 471 -1684 471 -1684 0 net=6667
rlabel metal2 499 -1684 499 -1684 0 net=4585
rlabel metal2 796 -1684 796 -1684 0 net=8003
rlabel metal2 1339 -1684 1339 -1684 0 net=9857
rlabel metal2 1353 -1684 1353 -1684 0 net=9985
rlabel metal2 352 -1686 352 -1686 0 net=1839
rlabel metal2 499 -1686 499 -1686 0 net=2929
rlabel metal2 527 -1686 527 -1686 0 net=10888
rlabel metal2 219 -1688 219 -1688 0 net=4003
rlabel metal2 359 -1688 359 -1688 0 net=1817
rlabel metal2 1118 -1688 1118 -1688 0 net=10611
rlabel metal2 1570 -1688 1570 -1688 0 net=11597
rlabel metal2 219 -1690 219 -1690 0 net=1599
rlabel metal2 380 -1690 380 -1690 0 net=592
rlabel metal2 534 -1690 534 -1690 0 net=3045
rlabel metal2 562 -1690 562 -1690 0 net=2753
rlabel metal2 884 -1690 884 -1690 0 net=6125
rlabel metal2 1150 -1690 1150 -1690 0 net=10263
rlabel metal2 1374 -1690 1374 -1690 0 net=10201
rlabel metal2 1528 -1690 1528 -1690 0 net=11487
rlabel metal2 173 -1692 173 -1692 0 net=738
rlabel metal2 380 -1692 380 -1692 0 net=3763
rlabel metal2 520 -1692 520 -1692 0 net=2967
rlabel metal2 912 -1692 912 -1692 0 net=7069
rlabel metal2 1164 -1692 1164 -1692 0 net=8845
rlabel metal2 1283 -1692 1283 -1692 0 net=9659
rlabel metal2 1374 -1692 1374 -1692 0 net=10347
rlabel metal2 177 -1694 177 -1694 0 net=11199
rlabel metal2 443 -1696 443 -1696 0 net=5761
rlabel metal2 873 -1696 873 -1696 0 net=9869
rlabel metal2 443 -1698 443 -1698 0 net=2283
rlabel metal2 534 -1698 534 -1698 0 net=3153
rlabel metal2 569 -1698 569 -1698 0 net=2005
rlabel metal2 723 -1698 723 -1698 0 net=6078
rlabel metal2 940 -1698 940 -1698 0 net=7501
rlabel metal2 1087 -1698 1087 -1698 0 net=8307
rlabel metal2 1178 -1698 1178 -1698 0 net=9183
rlabel metal2 1388 -1698 1388 -1698 0 net=10793
rlabel metal2 530 -1700 530 -1700 0 net=5712
rlabel metal2 929 -1700 929 -1700 0 net=8055
rlabel metal2 1108 -1700 1108 -1700 0 net=8515
rlabel metal2 1185 -1700 1185 -1700 0 net=8975
rlabel metal2 1297 -1700 1297 -1700 0 net=9759
rlabel metal2 128 -1702 128 -1702 0 net=2139
rlabel metal2 940 -1702 940 -1702 0 net=7253
rlabel metal2 1094 -1702 1094 -1702 0 net=8583
rlabel metal2 1199 -1702 1199 -1702 0 net=9507
rlabel metal2 1290 -1702 1290 -1702 0 net=9011
rlabel metal2 93 -1704 93 -1704 0 net=5859
rlabel metal2 541 -1704 541 -1704 0 net=11256
rlabel metal2 93 -1706 93 -1706 0 net=4429
rlabel metal2 765 -1706 765 -1706 0 net=5319
rlabel metal2 1108 -1706 1108 -1706 0 net=8755
rlabel metal2 1192 -1706 1192 -1706 0 net=9165
rlabel metal2 1451 -1706 1451 -1706 0 net=10927
rlabel metal2 96 -1708 96 -1708 0 net=7263
rlabel metal2 1129 -1708 1129 -1708 0 net=8689
rlabel metal2 1360 -1708 1360 -1708 0 net=10031
rlabel metal2 159 -1710 159 -1710 0 net=8317
rlabel metal2 1136 -1710 1136 -1710 0 net=8741
rlabel metal2 1325 -1710 1325 -1710 0 net=9767
rlabel metal2 247 -1712 247 -1712 0 net=1505
rlabel metal2 1311 -1712 1311 -1712 0 net=9391
rlabel metal2 247 -1714 247 -1714 0 net=4049
rlabel metal2 506 -1714 506 -1714 0 net=4279
rlabel metal2 821 -1714 821 -1714 0 net=8297
rlabel metal2 1248 -1714 1248 -1714 0 net=9329
rlabel metal2 394 -1716 394 -1716 0 net=3339
rlabel metal2 544 -1716 544 -1716 0 net=4435
rlabel metal2 621 -1716 621 -1716 0 net=8441
rlabel metal2 394 -1718 394 -1718 0 net=3263
rlabel metal2 569 -1718 569 -1718 0 net=3653
rlabel metal2 800 -1718 800 -1718 0 net=5839
rlabel metal2 828 -1718 828 -1718 0 net=8187
rlabel metal2 401 -1720 401 -1720 0 net=6673
rlabel metal2 583 -1720 583 -1720 0 net=3517
rlabel metal2 611 -1720 611 -1720 0 net=11331
rlabel metal2 114 -1722 114 -1722 0 net=4423
rlabel metal2 646 -1722 646 -1722 0 net=4211
rlabel metal2 670 -1722 670 -1722 0 net=8539
rlabel metal2 114 -1724 114 -1724 0 net=5307
rlabel metal2 597 -1724 597 -1724 0 net=3383
rlabel metal2 653 -1724 653 -1724 0 net=6365
rlabel metal2 800 -1724 800 -1724 0 net=8126
rlabel metal2 303 -1726 303 -1726 0 net=3905
rlabel metal2 590 -1726 590 -1726 0 net=6977
rlabel metal2 1031 -1726 1031 -1726 0 net=7887
rlabel metal2 1384 -1726 1384 -1726 0 net=1
rlabel metal2 303 -1728 303 -1728 0 net=4447
rlabel metal2 688 -1730 688 -1730 0 net=5278
rlabel metal2 926 -1730 926 -1730 0 net=6833
rlabel metal2 485 -1732 485 -1732 0 net=4594
rlabel metal2 345 -1734 345 -1734 0 net=2911
rlabel metal2 30 -1745 30 -1745 0 net=5861
rlabel metal2 159 -1745 159 -1745 0 net=639
rlabel metal2 534 -1745 534 -1745 0 net=3155
rlabel metal2 534 -1745 534 -1745 0 net=3155
rlabel metal2 541 -1745 541 -1745 0 net=4280
rlabel metal2 810 -1745 810 -1745 0 net=6888
rlabel metal2 884 -1745 884 -1745 0 net=7255
rlabel metal2 978 -1745 978 -1745 0 net=11146
rlabel metal2 1682 -1745 1682 -1745 0 net=11435
rlabel metal2 58 -1747 58 -1747 0 net=2931
rlabel metal2 502 -1747 502 -1747 0 net=5762
rlabel metal2 866 -1747 866 -1747 0 net=5937
rlabel metal2 61 -1749 61 -1749 0 net=4004
rlabel metal2 401 -1749 401 -1749 0 net=6675
rlabel metal2 989 -1749 989 -1749 0 net=11388
rlabel metal2 1748 -1749 1748 -1749 0 net=8870
rlabel metal2 1780 -1749 1780 -1749 0 net=8633
rlabel metal2 65 -1751 65 -1751 0 net=4992
rlabel metal2 264 -1751 264 -1751 0 net=1045
rlabel metal2 264 -1751 264 -1751 0 net=1045
rlabel metal2 275 -1751 275 -1751 0 net=2550
rlabel metal2 450 -1751 450 -1751 0 net=2382
rlabel metal2 1367 -1751 1367 -1751 0 net=11547
rlabel metal2 1752 -1751 1752 -1751 0 net=11923
rlabel metal2 65 -1753 65 -1753 0 net=8465
rlabel metal2 177 -1753 177 -1753 0 net=11252
rlabel metal2 1738 -1753 1738 -1753 0 net=11909
rlabel metal2 1759 -1753 1759 -1753 0 net=11989
rlabel metal2 1759 -1753 1759 -1753 0 net=11989
rlabel metal2 107 -1755 107 -1755 0 net=1687
rlabel metal2 159 -1755 159 -1755 0 net=2248
rlabel metal2 324 -1755 324 -1755 0 net=1978
rlabel metal2 604 -1755 604 -1755 0 net=3519
rlabel metal2 604 -1755 604 -1755 0 net=3519
rlabel metal2 618 -1755 618 -1755 0 net=4437
rlabel metal2 740 -1755 740 -1755 0 net=6422
rlabel metal2 1069 -1755 1069 -1755 0 net=10794
rlabel metal2 1612 -1755 1612 -1755 0 net=11333
rlabel metal2 1710 -1755 1710 -1755 0 net=11703
rlabel metal2 107 -1757 107 -1757 0 net=8298
rlabel metal2 1199 -1757 1199 -1757 0 net=8743
rlabel metal2 1332 -1757 1332 -1757 0 net=9549
rlabel metal2 1374 -1757 1374 -1757 0 net=10349
rlabel metal2 1605 -1757 1605 -1757 0 net=10713
rlabel metal2 1626 -1757 1626 -1757 0 net=10985
rlabel metal2 1696 -1757 1696 -1757 0 net=11657
rlabel metal2 110 -1759 110 -1759 0 net=2141
rlabel metal2 275 -1759 275 -1759 0 net=1851
rlabel metal2 814 -1759 814 -1759 0 net=6381
rlabel metal2 870 -1759 870 -1759 0 net=9591
rlabel metal2 1080 -1759 1080 -1759 0 net=7888
rlabel metal2 1160 -1759 1160 -1759 0 net=8004
rlabel metal2 1374 -1759 1374 -1759 0 net=10449
rlabel metal2 1528 -1759 1528 -1759 0 net=11201
rlabel metal2 114 -1761 114 -1761 0 net=5309
rlabel metal2 667 -1761 667 -1761 0 net=4519
rlabel metal2 793 -1761 793 -1761 0 net=5749
rlabel metal2 887 -1761 887 -1761 0 net=9272
rlabel metal2 1444 -1761 1444 -1761 0 net=9221
rlabel metal2 1528 -1761 1528 -1761 0 net=11349
rlabel metal2 1633 -1761 1633 -1761 0 net=11599
rlabel metal2 114 -1763 114 -1763 0 net=4981
rlabel metal2 408 -1763 408 -1763 0 net=2913
rlabel metal2 625 -1763 625 -1763 0 net=3851
rlabel metal2 677 -1763 677 -1763 0 net=4910
rlabel metal2 800 -1763 800 -1763 0 net=7502
rlabel metal2 1052 -1763 1052 -1763 0 net=7919
rlabel metal2 1052 -1763 1052 -1763 0 net=7919
rlabel metal2 1073 -1763 1073 -1763 0 net=7479
rlabel metal2 1108 -1763 1108 -1763 0 net=8757
rlabel metal2 1276 -1763 1276 -1763 0 net=9113
rlabel metal2 1430 -1763 1430 -1763 0 net=9995
rlabel metal2 1563 -1763 1563 -1763 0 net=11059
rlabel metal2 149 -1765 149 -1765 0 net=7757
rlabel metal2 1111 -1765 1111 -1765 0 net=11678
rlabel metal2 149 -1767 149 -1767 0 net=1675
rlabel metal2 191 -1767 191 -1767 0 net=4420
rlabel metal2 478 -1767 478 -1767 0 net=11941
rlabel metal2 170 -1769 170 -1769 0 net=2663
rlabel metal2 821 -1769 821 -1769 0 net=5841
rlabel metal2 891 -1769 891 -1769 0 net=9656
rlabel metal2 1549 -1769 1549 -1769 0 net=11529
rlabel metal2 180 -1771 180 -1771 0 net=2182
rlabel metal2 436 -1771 436 -1771 0 net=2285
rlabel metal2 625 -1771 625 -1771 0 net=5135
rlabel metal2 733 -1771 733 -1771 0 net=9275
rlabel metal2 1584 -1771 1584 -1771 0 net=11099
rlabel metal2 180 -1773 180 -1773 0 net=9430
rlabel metal2 184 -1775 184 -1775 0 net=3247
rlabel metal2 688 -1775 688 -1775 0 net=6960
rlabel metal2 989 -1775 989 -1775 0 net=6835
rlabel metal2 1041 -1775 1041 -1775 0 net=8976
rlabel metal2 1279 -1775 1279 -1775 0 net=10497
rlabel metal2 1570 -1775 1570 -1775 0 net=11489
rlabel metal2 191 -1777 191 -1777 0 net=10780
rlabel metal2 208 -1779 208 -1779 0 net=2839
rlabel metal2 548 -1779 548 -1779 0 net=7425
rlabel metal2 1017 -1779 1017 -1779 0 net=7803
rlabel metal2 1234 -1779 1234 -1779 0 net=9075
rlabel metal2 1521 -1779 1521 -1779 0 net=10817
rlabel metal2 1591 -1779 1591 -1779 0 net=11197
rlabel metal2 233 -1781 233 -1781 0 net=2266
rlabel metal2 348 -1781 348 -1781 0 net=2140
rlabel metal2 849 -1781 849 -1781 0 net=6119
rlabel metal2 915 -1781 915 -1781 0 net=9760
rlabel metal2 1507 -1781 1507 -1781 0 net=10613
rlabel metal2 233 -1783 233 -1783 0 net=3099
rlabel metal2 576 -1783 576 -1783 0 net=3935
rlabel metal2 695 -1783 695 -1783 0 net=4587
rlabel metal2 821 -1783 821 -1783 0 net=9508
rlabel metal2 1381 -1783 1381 -1783 0 net=10319
rlabel metal2 1556 -1783 1556 -1783 0 net=10881
rlabel metal2 240 -1785 240 -1785 0 net=1619
rlabel metal2 240 -1785 240 -1785 0 net=1619
rlabel metal2 268 -1785 268 -1785 0 net=2043
rlabel metal2 411 -1785 411 -1785 0 net=392
rlabel metal2 824 -1785 824 -1785 0 net=11477
rlabel metal2 268 -1787 268 -1787 0 net=3655
rlabel metal2 576 -1787 576 -1787 0 net=6165
rlabel metal2 919 -1787 919 -1787 0 net=11776
rlabel metal2 282 -1789 282 -1789 0 net=1513
rlabel metal2 317 -1789 317 -1789 0 net=6187
rlabel metal2 632 -1789 632 -1789 0 net=3987
rlabel metal2 702 -1789 702 -1789 0 net=8442
rlabel metal2 1220 -1789 1220 -1789 0 net=8619
rlabel metal2 1269 -1789 1269 -1789 0 net=9331
rlabel metal2 1465 -1789 1465 -1789 0 net=10203
rlabel metal2 1703 -1789 1703 -1789 0 net=11689
rlabel metal2 156 -1791 156 -1791 0 net=10023
rlabel metal2 1675 -1791 1675 -1791 0 net=11625
rlabel metal2 156 -1793 156 -1793 0 net=3563
rlabel metal2 639 -1793 639 -1793 0 net=4013
rlabel metal2 709 -1793 709 -1793 0 net=4729
rlabel metal2 828 -1793 828 -1793 0 net=7070
rlabel metal2 1171 -1793 1171 -1793 0 net=8407
rlabel metal2 198 -1795 198 -1795 0 net=1637
rlabel metal2 324 -1795 324 -1795 0 net=3265
rlabel metal2 415 -1795 415 -1795 0 net=1789
rlabel metal2 926 -1795 926 -1795 0 net=1506
rlabel metal2 1157 -1795 1157 -1795 0 net=9830
rlabel metal2 1675 -1795 1675 -1795 0 net=10773
rlabel metal2 198 -1797 198 -1797 0 net=3355
rlabel metal2 639 -1797 639 -1797 0 net=4213
rlabel metal2 709 -1797 709 -1797 0 net=4281
rlabel metal2 1115 -1797 1115 -1797 0 net=8517
rlabel metal2 1178 -1797 1178 -1797 0 net=8541
rlabel metal2 1276 -1797 1276 -1797 0 net=11587
rlabel metal2 247 -1799 247 -1799 0 net=4051
rlabel metal2 289 -1799 289 -1799 0 net=8017
rlabel metal2 1283 -1799 1283 -1799 0 net=9167
rlabel metal2 1416 -1799 1416 -1799 0 net=8349
rlabel metal2 121 -1801 121 -1801 0 net=4027
rlabel metal2 310 -1801 310 -1801 0 net=1901
rlabel metal2 422 -1801 422 -1801 0 net=1769
rlabel metal2 716 -1801 716 -1801 0 net=6953
rlabel metal2 1017 -1801 1017 -1801 0 net=9356
rlabel metal2 1731 -1801 1731 -1801 0 net=11829
rlabel metal2 93 -1803 93 -1803 0 net=4431
rlabel metal2 737 -1803 737 -1803 0 net=9585
rlabel metal2 1717 -1803 1717 -1803 0 net=11811
rlabel metal2 93 -1805 93 -1805 0 net=10153
rlabel metal2 303 -1805 303 -1805 0 net=4449
rlabel metal2 744 -1805 744 -1805 0 net=4568
rlabel metal2 919 -1805 919 -1805 0 net=6253
rlabel metal2 79 -1807 79 -1807 0 net=3125
rlabel metal2 331 -1807 331 -1807 0 net=2671
rlabel metal2 359 -1807 359 -1807 0 net=1819
rlabel metal2 674 -1807 674 -1807 0 net=3713
rlabel metal2 1153 -1807 1153 -1807 0 net=10145
rlabel metal2 79 -1809 79 -1809 0 net=3765
rlabel metal2 446 -1809 446 -1809 0 net=9495
rlabel metal2 121 -1811 121 -1811 0 net=3341
rlabel metal2 744 -1811 744 -1811 0 net=5121
rlabel metal2 758 -1811 758 -1811 0 net=5237
rlabel metal2 828 -1811 828 -1811 0 net=12029
rlabel metal2 135 -1813 135 -1813 0 net=4483
rlabel metal2 772 -1813 772 -1813 0 net=4569
rlabel metal2 100 -1815 100 -1815 0 net=2031
rlabel metal2 205 -1815 205 -1815 0 net=8439
rlabel metal2 331 -1815 331 -1815 0 net=4853
rlabel metal2 464 -1815 464 -1815 0 net=2833
rlabel metal2 611 -1815 611 -1815 0 net=4425
rlabel metal2 789 -1815 789 -1815 0 net=11679
rlabel metal2 100 -1817 100 -1817 0 net=2077
rlabel metal2 338 -1817 338 -1817 0 net=4204
rlabel metal2 506 -1817 506 -1817 0 net=3047
rlabel metal2 597 -1817 597 -1817 0 net=3385
rlabel metal2 849 -1817 849 -1817 0 net=8057
rlabel metal2 1101 -1817 1101 -1817 0 net=8911
rlabel metal2 1290 -1817 1290 -1817 0 net=7455
rlabel metal2 86 -1819 86 -1819 0 net=3113
rlabel metal2 597 -1819 597 -1819 0 net=4697
rlabel metal2 863 -1819 863 -1819 0 net=6871
rlabel metal2 1542 -1819 1542 -1819 0 net=9464
rlabel metal2 72 -1821 72 -1821 0 net=4679
rlabel metal2 205 -1821 205 -1821 0 net=8818
rlabel metal2 1458 -1821 1458 -1821 0 net=10075
rlabel metal2 44 -1823 44 -1823 0 net=2535
rlabel metal2 212 -1823 212 -1823 0 net=5597
rlabel metal2 863 -1823 863 -1823 0 net=6710
rlabel metal2 1423 -1823 1423 -1823 0 net=9987
rlabel metal2 44 -1825 44 -1825 0 net=2497
rlabel metal2 212 -1825 212 -1825 0 net=6669
rlabel metal2 912 -1825 912 -1825 0 net=6127
rlabel metal2 982 -1825 982 -1825 0 net=7960
rlabel metal2 1339 -1825 1339 -1825 0 net=9859
rlabel metal2 163 -1827 163 -1827 0 net=1707
rlabel metal2 926 -1827 926 -1827 0 net=10928
rlabel metal2 219 -1829 219 -1829 0 net=1601
rlabel metal2 338 -1829 338 -1829 0 net=433
rlabel metal2 471 -1829 471 -1829 0 net=1840
rlabel metal2 831 -1829 831 -1829 0 net=8095
rlabel metal2 1402 -1829 1402 -1829 0 net=10223
rlabel metal2 219 -1831 219 -1831 0 net=7233
rlabel metal2 929 -1831 929 -1831 0 net=9482
rlabel metal2 359 -1833 359 -1833 0 net=1783
rlabel metal2 380 -1833 380 -1833 0 net=2725
rlabel metal2 492 -1833 492 -1833 0 net=2503
rlabel metal2 936 -1833 936 -1833 0 net=8308
rlabel metal2 1206 -1833 1206 -1833 0 net=8773
rlabel metal2 1395 -1833 1395 -1833 0 net=9803
rlabel metal2 37 -1835 37 -1835 0 net=8808
rlabel metal2 947 -1835 947 -1835 0 net=7265
rlabel metal2 37 -1837 37 -1837 0 net=4545
rlabel metal2 247 -1837 247 -1837 0 net=3553
rlabel metal2 898 -1837 898 -1837 0 net=6813
rlabel metal2 975 -1837 975 -1837 0 net=9823
rlabel metal2 1206 -1837 1206 -1837 0 net=9185
rlabel metal2 1346 -1837 1346 -1837 0 net=9661
rlabel metal2 51 -1839 51 -1839 0 net=1797
rlabel metal2 373 -1839 373 -1839 0 net=2755
rlabel metal2 898 -1839 898 -1839 0 net=6529
rlabel metal2 933 -1839 933 -1839 0 net=8985
rlabel metal2 142 -1841 142 -1841 0 net=11421
rlabel metal2 401 -1841 401 -1841 0 net=2565
rlabel metal2 562 -1841 562 -1841 0 net=1565
rlabel metal2 856 -1841 856 -1841 0 net=5320
rlabel metal2 996 -1841 996 -1841 0 net=8475
rlabel metal2 1227 -1841 1227 -1841 0 net=8847
rlabel metal2 1297 -1841 1297 -1841 0 net=9013
rlabel metal2 429 -1843 429 -1843 0 net=3863
rlabel metal2 656 -1843 656 -1843 0 net=7909
rlabel metal2 1251 -1843 1251 -1843 0 net=10103
rlabel metal2 681 -1845 681 -1845 0 net=5583
rlabel metal2 961 -1845 961 -1845 0 net=6767
rlabel metal2 1003 -1845 1003 -1845 0 net=7359
rlabel metal2 1038 -1845 1038 -1845 0 net=7721
rlabel metal2 1143 -1845 1143 -1845 0 net=8691
rlabel metal2 1297 -1845 1297 -1845 0 net=10653
rlabel metal2 345 -1847 345 -1847 0 net=5171
rlabel metal2 1045 -1847 1045 -1847 0 net=10557
rlabel metal2 583 -1849 583 -1849 0 net=3907
rlabel metal2 835 -1849 835 -1849 0 net=6823
rlabel metal2 1024 -1849 1024 -1849 0 net=7545
rlabel metal2 1353 -1849 1353 -1849 0 net=10265
rlabel metal2 583 -1851 583 -1851 0 net=6979
rlabel metal2 653 -1851 653 -1851 0 net=6367
rlabel metal2 968 -1851 968 -1851 0 net=6580
rlabel metal2 1027 -1851 1027 -1851 0 net=11033
rlabel metal2 450 -1853 450 -1853 0 net=3133
rlabel metal2 968 -1853 968 -1853 0 net=2513
rlabel metal2 1048 -1853 1048 -1853 0 net=10157
rlabel metal2 590 -1855 590 -1855 0 net=2007
rlabel metal2 1066 -1855 1066 -1855 0 net=8319
rlabel metal2 1353 -1855 1353 -1855 0 net=10301
rlabel metal2 660 -1857 660 -1857 0 net=6333
rlabel metal2 905 -1857 905 -1857 0 net=7929
rlabel metal2 1451 -1857 1451 -1857 0 net=10033
rlabel metal2 807 -1859 807 -1859 0 net=9973
rlabel metal2 905 -1861 905 -1861 0 net=10546
rlabel metal2 1094 -1863 1094 -1863 0 net=8189
rlabel metal2 1409 -1863 1409 -1863 0 net=9871
rlabel metal2 194 -1865 194 -1865 0 net=9695
rlabel metal2 1094 -1867 1094 -1867 0 net=8257
rlabel metal2 1122 -1869 1122 -1869 0 net=8585
rlabel metal2 1185 -1871 1185 -1871 0 net=9769
rlabel metal2 1325 -1873 1325 -1873 0 net=9393
rlabel metal2 723 -1875 723 -1875 0 net=9199
rlabel metal2 387 -1877 387 -1877 0 net=6225
rlabel metal2 387 -1879 387 -1879 0 net=2969
rlabel metal2 250 -1881 250 -1881 0 net=3579
rlabel metal2 51 -1892 51 -1892 0 net=1798
rlabel metal2 233 -1892 233 -1892 0 net=3100
rlabel metal2 905 -1892 905 -1892 0 net=8758
rlabel metal2 1216 -1892 1216 -1892 0 net=7910
rlabel metal2 1234 -1892 1234 -1892 0 net=8621
rlabel metal2 1234 -1892 1234 -1892 0 net=8621
rlabel metal2 1276 -1892 1276 -1892 0 net=10224
rlabel metal2 1654 -1892 1654 -1892 0 net=11198
rlabel metal2 51 -1894 51 -1894 0 net=3657
rlabel metal2 296 -1894 296 -1894 0 net=1515
rlabel metal2 296 -1894 296 -1894 0 net=1515
rlabel metal2 303 -1894 303 -1894 0 net=3126
rlabel metal2 478 -1894 478 -1894 0 net=6189
rlabel metal2 912 -1894 912 -1894 0 net=6129
rlabel metal2 912 -1894 912 -1894 0 net=6129
rlabel metal2 919 -1894 919 -1894 0 net=6255
rlabel metal2 1017 -1894 1017 -1894 0 net=7546
rlabel metal2 1171 -1894 1171 -1894 0 net=8409
rlabel metal2 1171 -1894 1171 -1894 0 net=8409
rlabel metal2 1276 -1894 1276 -1894 0 net=8351
rlabel metal2 1668 -1894 1668 -1894 0 net=11531
rlabel metal2 1668 -1894 1668 -1894 0 net=11531
rlabel metal2 1773 -1894 1773 -1894 0 net=11436
rlabel metal2 65 -1896 65 -1896 0 net=8466
rlabel metal2 65 -1896 65 -1896 0 net=8466
rlabel metal2 68 -1896 68 -1896 0 net=7426
rlabel metal2 572 -1896 572 -1896 0 net=8986
rlabel metal2 1381 -1896 1381 -1896 0 net=9587
rlabel metal2 1409 -1896 1409 -1896 0 net=9696
rlabel metal2 1794 -1896 1794 -1896 0 net=5939
rlabel metal2 72 -1898 72 -1898 0 net=2536
rlabel metal2 135 -1898 135 -1898 0 net=2033
rlabel metal2 303 -1898 303 -1898 0 net=1567
rlabel metal2 593 -1898 593 -1898 0 net=9974
rlabel metal2 1493 -1898 1493 -1898 0 net=9223
rlabel metal2 72 -1900 72 -1900 0 net=1677
rlabel metal2 156 -1900 156 -1900 0 net=6797
rlabel metal2 240 -1900 240 -1900 0 net=1621
rlabel metal2 240 -1900 240 -1900 0 net=1621
rlabel metal2 250 -1900 250 -1900 0 net=372
rlabel metal2 562 -1900 562 -1900 0 net=6815
rlabel metal2 954 -1900 954 -1900 0 net=2514
rlabel metal2 1024 -1900 1024 -1900 0 net=11990
rlabel metal2 79 -1902 79 -1902 0 net=3767
rlabel metal2 345 -1902 345 -1902 0 net=5173
rlabel metal2 831 -1902 831 -1902 0 net=6872
rlabel metal2 1111 -1902 1111 -1902 0 net=11690
rlabel metal2 79 -1904 79 -1904 0 net=3387
rlabel metal2 646 -1904 646 -1904 0 net=5598
rlabel metal2 796 -1904 796 -1904 0 net=6382
rlabel metal2 849 -1904 849 -1904 0 net=8059
rlabel metal2 1279 -1904 1279 -1904 0 net=11885
rlabel metal2 86 -1906 86 -1906 0 net=4680
rlabel metal2 135 -1906 135 -1906 0 net=2567
rlabel metal2 436 -1906 436 -1906 0 net=2286
rlabel metal2 1024 -1906 1024 -1906 0 net=8191
rlabel metal2 1153 -1906 1153 -1906 0 net=11812
rlabel metal2 86 -1908 86 -1908 0 net=8440
rlabel metal2 324 -1908 324 -1908 0 net=3266
rlabel metal2 499 -1908 499 -1908 0 net=2431
rlabel metal2 922 -1908 922 -1908 0 net=794
rlabel metal2 1031 -1908 1031 -1908 0 net=7361
rlabel metal2 1115 -1908 1115 -1908 0 net=8519
rlabel metal2 1283 -1908 1283 -1908 0 net=9169
rlabel metal2 1283 -1908 1283 -1908 0 net=9169
rlabel metal2 1314 -1908 1314 -1908 0 net=11478
rlabel metal2 1731 -1908 1731 -1908 0 net=11911
rlabel metal2 89 -1910 89 -1910 0 net=7111
rlabel metal2 1353 -1910 1353 -1910 0 net=10303
rlabel metal2 1633 -1910 1633 -1910 0 net=11335
rlabel metal2 1752 -1910 1752 -1910 0 net=11943
rlabel metal2 100 -1912 100 -1912 0 net=2078
rlabel metal2 464 -1912 464 -1912 0 net=5750
rlabel metal2 926 -1912 926 -1912 0 net=6768
rlabel metal2 1003 -1912 1003 -1912 0 net=6825
rlabel metal2 1139 -1912 1139 -1912 0 net=3821
rlabel metal2 1780 -1912 1780 -1912 0 net=5077
rlabel metal2 100 -1914 100 -1914 0 net=11207
rlabel metal2 1801 -1914 1801 -1914 0 net=8635
rlabel metal2 110 -1916 110 -1916 0 net=4891
rlabel metal2 509 -1916 509 -1916 0 net=9197
rlabel metal2 1381 -1916 1381 -1916 0 net=10205
rlabel metal2 142 -1918 142 -1918 0 net=11423
rlabel metal2 142 -1920 142 -1920 0 net=9496
rlabel metal2 145 -1922 145 -1922 0 net=2987
rlabel metal2 324 -1922 324 -1922 0 net=1903
rlabel metal2 527 -1922 527 -1922 0 net=11588
rlabel metal2 149 -1924 149 -1924 0 net=407
rlabel metal2 212 -1924 212 -1924 0 net=6670
rlabel metal2 527 -1924 527 -1924 0 net=3715
rlabel metal2 723 -1924 723 -1924 0 net=6227
rlabel metal2 957 -1924 957 -1924 0 net=9114
rlabel metal2 1409 -1924 1409 -1924 0 net=10321
rlabel metal2 1626 -1924 1626 -1924 0 net=10987
rlabel metal2 156 -1926 156 -1926 0 net=3249
rlabel metal2 191 -1926 191 -1926 0 net=4459
rlabel metal2 334 -1926 334 -1926 0 net=1855
rlabel metal2 541 -1926 541 -1926 0 net=2841
rlabel metal2 618 -1926 618 -1926 0 net=5311
rlabel metal2 929 -1926 929 -1926 0 net=5941
rlabel metal2 1027 -1926 1027 -1926 0 net=11605
rlabel metal2 128 -1928 128 -1928 0 net=1689
rlabel metal2 191 -1928 191 -1928 0 net=1791
rlabel metal2 506 -1928 506 -1928 0 net=3049
rlabel metal2 597 -1928 597 -1928 0 net=4699
rlabel metal2 800 -1928 800 -1928 0 net=9824
rlabel metal2 1031 -1928 1031 -1928 0 net=7481
rlabel metal2 1143 -1928 1143 -1928 0 net=8745
rlabel metal2 1318 -1928 1318 -1928 0 net=9395
rlabel metal2 1374 -1928 1374 -1928 0 net=10451
rlabel metal2 1626 -1928 1626 -1928 0 net=10775
rlabel metal2 152 -1930 152 -1930 0 net=6537
rlabel metal2 457 -1930 457 -1930 0 net=3555
rlabel metal2 604 -1930 604 -1930 0 net=3521
rlabel metal2 604 -1930 604 -1930 0 net=3521
rlabel metal2 618 -1930 618 -1930 0 net=4215
rlabel metal2 653 -1930 653 -1930 0 net=7804
rlabel metal2 1248 -1930 1248 -1930 0 net=8849
rlabel metal2 1360 -1930 1360 -1930 0 net=9997
rlabel metal2 1675 -1930 1675 -1930 0 net=11659
rlabel metal2 37 -1932 37 -1932 0 net=4546
rlabel metal2 506 -1932 506 -1932 0 net=11991
rlabel metal2 159 -1934 159 -1934 0 net=4987
rlabel metal2 901 -1934 901 -1934 0 net=10867
rlabel metal2 1710 -1934 1710 -1934 0 net=11831
rlabel metal2 163 -1936 163 -1936 0 net=1708
rlabel metal2 254 -1936 254 -1936 0 net=2142
rlabel metal2 1059 -1936 1059 -1936 0 net=9593
rlabel metal2 1374 -1936 1374 -1936 0 net=9663
rlabel metal2 1423 -1936 1423 -1936 0 net=9861
rlabel metal2 163 -1938 163 -1938 0 net=5287
rlabel metal2 345 -1938 345 -1938 0 net=3865
rlabel metal2 632 -1938 632 -1938 0 net=3565
rlabel metal2 653 -1938 653 -1938 0 net=1995
rlabel metal2 1045 -1938 1045 -1938 0 net=10654
rlabel metal2 1395 -1938 1395 -1938 0 net=10159
rlabel metal2 93 -1940 93 -1940 0 net=10155
rlabel metal2 93 -1942 93 -1942 0 net=7819
rlabel metal2 198 -1942 198 -1942 0 net=3357
rlabel metal2 632 -1942 632 -1942 0 net=4015
rlabel metal2 737 -1942 737 -1942 0 net=4451
rlabel metal2 737 -1942 737 -1942 0 net=4451
rlabel metal2 751 -1942 751 -1942 0 net=4427
rlabel metal2 751 -1942 751 -1942 0 net=4427
rlabel metal2 772 -1942 772 -1942 0 net=4571
rlabel metal2 772 -1942 772 -1942 0 net=4571
rlabel metal2 793 -1942 793 -1942 0 net=4731
rlabel metal2 807 -1942 807 -1942 0 net=6368
rlabel metal2 968 -1942 968 -1942 0 net=8097
rlabel metal2 1423 -1942 1423 -1942 0 net=10267
rlabel metal2 103 -1944 103 -1944 0 net=9509
rlabel metal2 1437 -1944 1437 -1944 0 net=9873
rlabel metal2 1514 -1944 1514 -1944 0 net=10351
rlabel metal2 170 -1946 170 -1946 0 net=2665
rlabel metal2 460 -1946 460 -1946 0 net=3613
rlabel metal2 807 -1946 807 -1946 0 net=6121
rlabel metal2 933 -1946 933 -1946 0 net=6677
rlabel metal2 975 -1946 975 -1946 0 net=10105
rlabel metal2 1402 -1946 1402 -1946 0 net=9805
rlabel metal2 1535 -1946 1535 -1946 0 net=10559
rlabel metal2 110 -1948 110 -1948 0 net=10231
rlabel metal2 1563 -1948 1563 -1948 0 net=10883
rlabel metal2 170 -1950 170 -1950 0 net=1603
rlabel metal2 247 -1950 247 -1950 0 net=1853
rlabel metal2 373 -1950 373 -1950 0 net=2757
rlabel metal2 380 -1950 380 -1950 0 net=2727
rlabel metal2 639 -1950 639 -1950 0 net=2623
rlabel metal2 824 -1950 824 -1950 0 net=7256
rlabel metal2 891 -1950 891 -1950 0 net=9988
rlabel metal2 114 -1952 114 -1952 0 net=4983
rlabel metal2 835 -1952 835 -1952 0 net=2453
rlabel metal2 1010 -1952 1010 -1952 0 net=6955
rlabel metal2 1080 -1952 1080 -1952 0 net=4595
rlabel metal2 1157 -1952 1157 -1952 0 net=9770
rlabel metal2 1206 -1952 1206 -1952 0 net=9187
rlabel metal2 1430 -1952 1430 -1952 0 net=9077
rlabel metal2 114 -1954 114 -1954 0 net=4053
rlabel metal2 373 -1954 373 -1954 0 net=2505
rlabel metal2 667 -1954 667 -1954 0 net=3853
rlabel metal2 719 -1954 719 -1954 0 net=62
rlabel metal2 1122 -1954 1122 -1954 0 net=8587
rlabel metal2 131 -1956 131 -1956 0 net=3185
rlabel metal2 254 -1956 254 -1956 0 net=3157
rlabel metal2 667 -1956 667 -1956 0 net=4485
rlabel metal2 786 -1956 786 -1956 0 net=4589
rlabel metal2 989 -1956 989 -1956 0 net=6837
rlabel metal2 1020 -1956 1020 -1956 0 net=6991
rlabel metal2 1087 -1956 1087 -1956 0 net=7723
rlabel metal2 1129 -1956 1129 -1956 0 net=7931
rlabel metal2 1206 -1956 1206 -1956 0 net=8693
rlabel metal2 1262 -1956 1262 -1956 0 net=10147
rlabel metal2 177 -1958 177 -1958 0 net=406
rlabel metal2 989 -1958 989 -1958 0 net=10818
rlabel metal2 180 -1960 180 -1960 0 net=180
rlabel metal2 814 -1960 814 -1960 0 net=5239
rlabel metal2 877 -1960 877 -1960 0 net=6649
rlabel metal2 1052 -1960 1052 -1960 0 net=7921
rlabel metal2 1241 -1960 1241 -1960 0 net=8775
rlabel metal2 1297 -1960 1297 -1960 0 net=9201
rlabel metal2 1486 -1960 1486 -1960 0 net=11101
rlabel metal2 180 -1962 180 -1962 0 net=1770
rlabel metal2 534 -1962 534 -1962 0 net=3115
rlabel metal2 590 -1962 590 -1962 0 net=2009
rlabel metal2 810 -1962 810 -1962 0 net=9419
rlabel metal2 1528 -1962 1528 -1962 0 net=11351
rlabel metal2 1619 -1962 1619 -1962 0 net=11203
rlabel metal2 58 -1964 58 -1964 0 net=2933
rlabel metal2 758 -1964 758 -1964 0 net=8320
rlabel metal2 1073 -1964 1073 -1964 0 net=7759
rlabel metal2 1220 -1964 1220 -1964 0 net=8543
rlabel metal2 1311 -1964 1311 -1964 0 net=10935
rlabel metal2 1640 -1964 1640 -1964 0 net=11549
rlabel metal2 58 -1966 58 -1966 0 net=4283
rlabel metal2 814 -1966 814 -1966 0 net=5585
rlabel metal2 1052 -1966 1052 -1966 0 net=8019
rlabel metal2 1192 -1966 1192 -1966 0 net=8477
rlabel metal2 1269 -1966 1269 -1966 0 net=9333
rlabel metal2 1384 -1966 1384 -1966 0 net=1
rlabel metal2 1528 -1966 1528 -1966 0 net=10499
rlabel metal2 1682 -1966 1682 -1966 0 net=11681
rlabel metal2 198 -1968 198 -1968 0 net=2291
rlabel metal2 838 -1968 838 -1968 0 net=7266
rlabel metal2 1542 -1968 1542 -1968 0 net=10077
rlabel metal2 205 -1970 205 -1970 0 net=4029
rlabel metal2 387 -1970 387 -1970 0 net=2971
rlabel metal2 649 -1970 649 -1970 0 net=11843
rlabel metal2 212 -1972 212 -1972 0 net=11034
rlabel metal2 219 -1974 219 -1974 0 net=7235
rlabel metal2 1178 -1974 1178 -1974 0 net=8913
rlabel metal2 1388 -1974 1388 -1974 0 net=10035
rlabel metal2 1598 -1974 1598 -1974 0 net=10715
rlabel metal2 219 -1976 219 -1976 0 net=3295
rlabel metal2 394 -1976 394 -1976 0 net=4433
rlabel metal2 856 -1976 856 -1976 0 net=5843
rlabel metal2 1017 -1976 1017 -1976 0 net=7071
rlabel metal2 1178 -1976 1178 -1976 0 net=9551
rlabel metal2 1465 -1976 1465 -1976 0 net=10025
rlabel metal2 1612 -1976 1612 -1976 0 net=11491
rlabel metal2 264 -1978 264 -1978 0 net=5297
rlabel metal2 422 -1978 422 -1978 0 net=4439
rlabel metal2 870 -1978 870 -1978 0 net=9349
rlabel metal2 1038 -1978 1038 -1978 0 net=10605
rlabel metal2 1661 -1978 1661 -1978 0 net=11627
rlabel metal2 275 -1980 275 -1980 0 net=1785
rlabel metal2 709 -1980 709 -1980 0 net=6531
rlabel metal2 1038 -1980 1038 -1980 0 net=11600
rlabel metal2 1703 -1980 1703 -1980 0 net=11705
rlabel metal2 282 -1982 282 -1982 0 net=2813
rlabel metal2 716 -1982 716 -1982 0 net=5713
rlabel metal2 1066 -1982 1066 -1982 0 net=7457
rlabel metal2 1293 -1982 1293 -1982 0 net=11723
rlabel metal2 1738 -1982 1738 -1982 0 net=11925
rlabel metal2 359 -1984 359 -1984 0 net=3937
rlabel metal2 723 -1984 723 -1984 0 net=4307
rlabel metal2 1073 -1984 1073 -1984 0 net=8259
rlabel metal2 1192 -1984 1192 -1984 0 net=10243
rlabel metal2 1465 -1984 1465 -1984 0 net=11061
rlabel metal2 1766 -1984 1766 -1984 0 net=12031
rlabel metal2 366 -1986 366 -1986 0 net=2045
rlabel metal2 583 -1986 583 -1986 0 net=6981
rlabel metal2 1304 -1986 1304 -1986 0 net=9015
rlabel metal2 1591 -1986 1591 -1986 0 net=10615
rlabel metal2 317 -1988 317 -1988 0 net=1639
rlabel metal2 583 -1988 583 -1988 0 net=5137
rlabel metal2 628 -1988 628 -1988 0 net=9297
rlabel metal2 317 -1990 317 -1990 0 net=2915
rlabel metal2 625 -1990 625 -1990 0 net=3988
rlabel metal2 730 -1990 730 -1990 0 net=4367
rlabel metal2 1160 -1990 1160 -1990 0 net=11461
rlabel metal2 352 -1992 352 -1992 0 net=2673
rlabel metal2 576 -1992 576 -1992 0 net=6167
rlabel metal2 919 -1992 919 -1992 0 net=4599
rlabel metal2 30 -1994 30 -1994 0 net=5863
rlabel metal2 681 -1994 681 -1994 0 net=3909
rlabel metal2 961 -1994 961 -1994 0 net=7805
rlabel metal2 30 -1996 30 -1996 0 net=4855
rlabel metal2 681 -1996 681 -1996 0 net=4521
rlabel metal2 44 -1998 44 -1998 0 net=2498
rlabel metal2 744 -1998 744 -1998 0 net=5123
rlabel metal2 44 -2000 44 -2000 0 net=2123
rlabel metal2 660 -2000 660 -2000 0 net=6335
rlabel metal2 124 -2002 124 -2002 0 net=5849
rlabel metal2 520 -2002 520 -2002 0 net=3581
rlabel metal2 513 -2004 513 -2004 0 net=2835
rlabel metal2 450 -2006 450 -2006 0 net=3135
rlabel metal2 450 -2008 450 -2008 0 net=3625
rlabel metal2 121 -2010 121 -2010 0 net=3342
rlabel metal2 121 -2012 121 -2012 0 net=9276
rlabel metal2 656 -2014 656 -2014 0 net=5075
rlabel metal2 37 -2025 37 -2025 0 net=7079
rlabel metal2 632 -2025 632 -2025 0 net=4017
rlabel metal2 632 -2025 632 -2025 0 net=4017
rlabel metal2 667 -2025 667 -2025 0 net=4487
rlabel metal2 702 -2025 702 -2025 0 net=3614
rlabel metal2 964 -2025 964 -2025 0 net=8020
rlabel metal2 1062 -2025 1062 -2025 0 net=4596
rlabel metal2 1139 -2025 1139 -2025 0 net=9806
rlabel metal2 1479 -2025 1479 -2025 0 net=5076
rlabel metal2 44 -2027 44 -2027 0 net=2124
rlabel metal2 719 -2027 719 -2027 0 net=5312
rlabel metal2 929 -2027 929 -2027 0 net=8588
rlabel metal2 1591 -2027 1591 -2027 0 net=11463
rlabel metal2 1713 -2027 1713 -2027 0 net=5940
rlabel metal2 44 -2029 44 -2029 0 net=3951
rlabel metal2 222 -2029 222 -2029 0 net=1854
rlabel metal2 278 -2029 278 -2029 0 net=7112
rlabel metal2 1195 -2029 1195 -2029 0 net=9862
rlabel metal2 1591 -2029 1591 -2029 0 net=10617
rlabel metal2 1745 -2029 1745 -2029 0 net=5078
rlabel metal2 51 -2031 51 -2031 0 net=3658
rlabel metal2 229 -2031 229 -2031 0 net=8060
rlabel metal2 1213 -2031 1213 -2031 0 net=11682
rlabel metal2 51 -2033 51 -2033 0 net=1787
rlabel metal2 296 -2033 296 -2033 0 net=1517
rlabel metal2 296 -2033 296 -2033 0 net=1517
rlabel metal2 331 -2033 331 -2033 0 net=2046
rlabel metal2 516 -2033 516 -2033 0 net=4590
rlabel metal2 954 -2033 954 -2033 0 net=9188
rlabel metal2 1423 -2033 1423 -2033 0 net=10269
rlabel metal2 1444 -2033 1444 -2033 0 net=10453
rlabel metal2 1682 -2033 1682 -2033 0 net=11833
rlabel metal2 61 -2035 61 -2035 0 net=6982
rlabel metal2 1157 -2035 1157 -2035 0 net=7933
rlabel metal2 72 -2037 72 -2037 0 net=1678
rlabel metal2 240 -2037 240 -2037 0 net=1622
rlabel metal2 331 -2037 331 -2037 0 net=1809
rlabel metal2 464 -2037 464 -2037 0 net=2973
rlabel metal2 520 -2037 520 -2037 0 net=2837
rlabel metal2 555 -2037 555 -2037 0 net=2934
rlabel metal2 590 -2037 590 -2037 0 net=3557
rlabel metal2 614 -2037 614 -2037 0 net=10106
rlabel metal2 996 -2037 996 -2037 0 net=7337
rlabel metal2 1395 -2037 1395 -2037 0 net=10161
rlabel metal2 1430 -2037 1430 -2037 0 net=10353
rlabel metal2 72 -2039 72 -2039 0 net=2035
rlabel metal2 338 -2039 338 -2039 0 net=3768
rlabel metal2 667 -2039 667 -2039 0 net=4369
rlabel metal2 744 -2039 744 -2039 0 net=6337
rlabel metal2 744 -2039 744 -2039 0 net=6337
rlabel metal2 751 -2039 751 -2039 0 net=4428
rlabel metal2 898 -2039 898 -2039 0 net=9203
rlabel metal2 1314 -2039 1314 -2039 0 net=11706
rlabel metal2 100 -2041 100 -2041 0 net=4440
rlabel metal2 520 -2041 520 -2041 0 net=3117
rlabel metal2 558 -2041 558 -2041 0 net=10593
rlabel metal2 1703 -2041 1703 -2041 0 net=11887
rlabel metal2 103 -2043 103 -2043 0 net=4988
rlabel metal2 877 -2043 877 -2043 0 net=6651
rlabel metal2 996 -2043 996 -2043 0 net=9552
rlabel metal2 1195 -2043 1195 -2043 0 net=11532
rlabel metal2 1724 -2043 1724 -2043 0 net=4601
rlabel metal2 103 -2045 103 -2045 0 net=1792
rlabel metal2 205 -2045 205 -2045 0 net=4031
rlabel metal2 702 -2045 702 -2045 0 net=9874
rlabel metal2 1514 -2045 1514 -2045 0 net=10937
rlabel metal2 1594 -2045 1594 -2045 0 net=1
rlabel metal2 1626 -2045 1626 -2045 0 net=10777
rlabel metal2 110 -2047 110 -2047 0 net=2857
rlabel metal2 177 -2047 177 -2047 0 net=5139
rlabel metal2 751 -2047 751 -2047 0 net=4573
rlabel metal2 786 -2047 786 -2047 0 net=2010
rlabel metal2 999 -2047 999 -2047 0 net=11926
rlabel metal2 114 -2049 114 -2049 0 net=4055
rlabel metal2 761 -2049 761 -2049 0 net=2454
rlabel metal2 842 -2049 842 -2049 0 net=5241
rlabel metal2 842 -2049 842 -2049 0 net=5241
rlabel metal2 856 -2049 856 -2049 0 net=5845
rlabel metal2 887 -2049 887 -2049 0 net=11204
rlabel metal2 1626 -2049 1626 -2049 0 net=11629
rlabel metal2 1738 -2049 1738 -2049 0 net=9225
rlabel metal2 114 -2051 114 -2051 0 net=1997
rlabel metal2 786 -2051 786 -2051 0 net=2985
rlabel metal2 905 -2051 905 -2051 0 net=6191
rlabel metal2 999 -2051 999 -2051 0 net=6826
rlabel metal2 1157 -2051 1157 -2051 0 net=8411
rlabel metal2 1199 -2051 1199 -2051 0 net=9511
rlabel metal2 1395 -2051 1395 -2051 0 net=10323
rlabel metal2 1451 -2051 1451 -2051 0 net=9079
rlabel metal2 1570 -2051 1570 -2051 0 net=11209
rlabel metal2 1619 -2051 1619 -2051 0 net=11551
rlabel metal2 1661 -2051 1661 -2051 0 net=11993
rlabel metal2 121 -2053 121 -2053 0 net=10156
rlabel metal2 1507 -2053 1507 -2053 0 net=9589
rlabel metal2 121 -2055 121 -2055 0 net=894
rlabel metal2 572 -2055 572 -2055 0 net=4087
rlabel metal2 695 -2055 695 -2055 0 net=6169
rlabel metal2 912 -2055 912 -2055 0 net=6131
rlabel metal2 1017 -2055 1017 -2055 0 net=7073
rlabel metal2 1052 -2055 1052 -2055 0 net=7363
rlabel metal2 1164 -2055 1164 -2055 0 net=8851
rlabel metal2 1293 -2055 1293 -2055 0 net=9016
rlabel metal2 1409 -2055 1409 -2055 0 net=10245
rlabel metal2 1458 -2055 1458 -2055 0 net=10501
rlabel metal2 1577 -2055 1577 -2055 0 net=10717
rlabel metal2 124 -2057 124 -2057 0 net=3317
rlabel metal2 219 -2057 219 -2057 0 net=9149
rlabel metal2 1332 -2057 1332 -2057 0 net=10037
rlabel metal2 1500 -2057 1500 -2057 0 net=11725
rlabel metal2 124 -2059 124 -2059 0 net=2988
rlabel metal2 338 -2059 338 -2059 0 net=1841
rlabel metal2 1171 -2059 1171 -2059 0 net=8777
rlabel metal2 1283 -2059 1283 -2059 0 net=9171
rlabel metal2 1507 -2059 1507 -2059 0 net=10885
rlabel metal2 1584 -2059 1584 -2059 0 net=11353
rlabel metal2 1689 -2059 1689 -2059 0 net=10989
rlabel metal2 131 -2061 131 -2061 0 net=6816
rlabel metal2 569 -2061 569 -2061 0 net=8853
rlabel metal2 1283 -2061 1283 -2061 0 net=9397
rlabel metal2 1563 -2061 1563 -2061 0 net=11493
rlabel metal2 1689 -2061 1689 -2061 0 net=11845
rlabel metal2 131 -2063 131 -2063 0 net=11424
rlabel metal2 135 -2065 135 -2065 0 net=2568
rlabel metal2 359 -2065 359 -2065 0 net=3938
rlabel metal2 394 -2065 394 -2065 0 net=4434
rlabel metal2 817 -2065 817 -2065 0 net=9350
rlabel metal2 873 -2065 873 -2065 0 net=11645
rlabel metal2 1612 -2065 1612 -2065 0 net=11607
rlabel metal2 1654 -2065 1654 -2065 0 net=11945
rlabel metal2 30 -2067 30 -2067 0 net=4857
rlabel metal2 142 -2067 142 -2067 0 net=5729
rlabel metal2 912 -2067 912 -2067 0 net=6229
rlabel metal2 968 -2067 968 -2067 0 net=8099
rlabel metal2 1241 -2067 1241 -2067 0 net=8353
rlabel metal2 1318 -2067 1318 -2067 0 net=10207
rlabel metal2 1647 -2067 1647 -2067 0 net=11913
rlabel metal2 30 -2069 30 -2069 0 net=8897
rlabel metal2 142 -2069 142 -2069 0 net=4309
rlabel metal2 793 -2069 793 -2069 0 net=5175
rlabel metal2 831 -2069 831 -2069 0 net=8544
rlabel metal2 1381 -2069 1381 -2069 0 net=10607
rlabel metal2 1731 -2069 1731 -2069 0 net=8637
rlabel metal2 145 -2071 145 -2071 0 net=5942
rlabel metal2 1024 -2071 1024 -2071 0 net=8193
rlabel metal2 1255 -2071 1255 -2071 0 net=9335
rlabel metal2 184 -2073 184 -2073 0 net=1691
rlabel metal2 317 -2073 317 -2073 0 net=2917
rlabel metal2 366 -2073 366 -2073 0 net=1640
rlabel metal2 548 -2073 548 -2073 0 net=11337
rlabel metal2 184 -2075 184 -2075 0 net=3321
rlabel metal2 233 -2075 233 -2075 0 net=6799
rlabel metal2 922 -2075 922 -2075 0 net=7922
rlabel metal2 1290 -2075 1290 -2075 0 net=11089
rlabel metal2 65 -2077 65 -2077 0 net=2373
rlabel metal2 240 -2077 240 -2077 0 net=1743
rlabel metal2 317 -2077 317 -2077 0 net=1905
rlabel metal2 366 -2077 366 -2077 0 net=2759
rlabel metal2 541 -2077 541 -2077 0 net=3051
rlabel metal2 628 -2077 628 -2077 0 net=4325
rlabel metal2 796 -2077 796 -2077 0 net=8967
rlabel metal2 65 -2079 65 -2079 0 net=2515
rlabel metal2 709 -2079 709 -2079 0 net=6533
rlabel metal2 1024 -2079 1024 -2079 0 net=8746
rlabel metal2 1185 -2079 1185 -2079 0 net=8915
rlabel metal2 86 -2081 86 -2081 0 net=5721
rlabel metal2 247 -2081 247 -2081 0 net=6567
rlabel metal2 541 -2081 541 -2081 0 net=4985
rlabel metal2 835 -2081 835 -2081 0 net=5103
rlabel metal2 1066 -2081 1066 -2081 0 net=7459
rlabel metal2 1066 -2081 1066 -2081 0 net=7459
rlabel metal2 1073 -2081 1073 -2081 0 net=8261
rlabel metal2 1143 -2081 1143 -2081 0 net=9299
rlabel metal2 86 -2083 86 -2083 0 net=2517
rlabel metal2 695 -2083 695 -2083 0 net=4453
rlabel metal2 821 -2083 821 -2083 0 net=10026
rlabel metal2 191 -2085 191 -2085 0 net=3627
rlabel metal2 457 -2085 457 -2085 0 net=3523
rlabel metal2 681 -2085 681 -2085 0 net=4523
rlabel metal2 856 -2085 856 -2085 0 net=5247
rlabel metal2 919 -2085 919 -2085 0 net=9497
rlabel metal2 1304 -2085 1304 -2085 0 net=9999
rlabel metal2 1472 -2085 1472 -2085 0 net=10305
rlabel metal2 93 -2087 93 -2087 0 net=7821
rlabel metal2 933 -2087 933 -2087 0 net=6679
rlabel metal2 989 -2087 989 -2087 0 net=9049
rlabel metal2 1493 -2087 1493 -2087 0 net=10869
rlabel metal2 93 -2089 93 -2089 0 net=11336
rlabel metal2 163 -2091 163 -2091 0 net=5289
rlabel metal2 660 -2091 660 -2091 0 net=3583
rlabel metal2 807 -2091 807 -2091 0 net=6123
rlabel metal2 947 -2091 947 -2091 0 net=6257
rlabel metal2 1031 -2091 1031 -2091 0 net=7483
rlabel metal2 1080 -2091 1080 -2091 0 net=7761
rlabel metal2 1262 -2091 1262 -2091 0 net=10149
rlabel metal2 1486 -2091 1486 -2091 0 net=11103
rlabel metal2 1633 -2091 1633 -2091 0 net=11661
rlabel metal2 163 -2093 163 -2093 0 net=2683
rlabel metal2 978 -2093 978 -2093 0 net=9281
rlabel metal2 1269 -2093 1269 -2093 0 net=9421
rlabel metal2 1675 -2093 1675 -2093 0 net=12033
rlabel metal2 198 -2095 198 -2095 0 net=2293
rlabel metal2 394 -2095 394 -2095 0 net=3137
rlabel metal2 555 -2095 555 -2095 0 net=7763
rlabel metal2 1010 -2095 1010 -2095 0 net=6839
rlabel metal2 1087 -2095 1087 -2095 0 net=7237
rlabel metal2 198 -2097 198 -2097 0 net=2201
rlabel metal2 254 -2097 254 -2097 0 net=3159
rlabel metal2 583 -2097 583 -2097 0 net=10633
rlabel metal2 254 -2099 254 -2099 0 net=5864
rlabel metal2 807 -2099 807 -2099 0 net=5715
rlabel metal2 891 -2099 891 -2099 0 net=5179
rlabel metal2 1325 -2099 1325 -2099 0 net=9595
rlabel metal2 156 -2101 156 -2101 0 net=3251
rlabel metal2 716 -2101 716 -2101 0 net=9697
rlabel metal2 58 -2103 58 -2103 0 net=4285
rlabel metal2 268 -2103 268 -2103 0 net=4461
rlabel metal2 429 -2103 429 -2103 0 net=3359
rlabel metal2 716 -2103 716 -2103 0 net=6043
rlabel metal2 226 -2105 226 -2105 0 net=3187
rlabel metal2 282 -2105 282 -2105 0 net=2815
rlabel metal2 814 -2105 814 -2105 0 net=5587
rlabel metal2 982 -2105 982 -2105 0 net=6993
rlabel metal2 1087 -2105 1087 -2105 0 net=8521
rlabel metal2 226 -2107 226 -2107 0 net=8831
rlabel metal2 1227 -2107 1227 -2107 0 net=9107
rlabel metal2 282 -2109 282 -2109 0 net=3717
rlabel metal2 1010 -2109 1010 -2109 0 net=9665
rlabel metal2 289 -2111 289 -2111 0 net=5299
rlabel metal2 1059 -2111 1059 -2111 0 net=6671
rlabel metal2 170 -2113 170 -2113 0 net=1604
rlabel metal2 324 -2113 324 -2113 0 net=2507
rlabel metal2 380 -2113 380 -2113 0 net=3296
rlabel metal2 1094 -2113 1094 -2113 0 net=7725
rlabel metal2 1129 -2113 1129 -2113 0 net=3822
rlabel metal2 170 -2115 170 -2115 0 net=2729
rlabel metal2 527 -2115 527 -2115 0 net=4701
rlabel metal2 1101 -2115 1101 -2115 0 net=7807
rlabel metal2 1374 -2115 1374 -2115 0 net=11063
rlabel metal2 107 -2117 107 -2117 0 net=10533
rlabel metal2 107 -2119 107 -2119 0 net=3910
rlabel metal2 758 -2119 758 -2119 0 net=10527
rlabel metal2 345 -2121 345 -2121 0 net=3867
rlabel metal2 499 -2121 499 -2121 0 net=2433
rlabel metal2 765 -2121 765 -2121 0 net=5125
rlabel metal2 345 -2123 345 -2123 0 net=1857
rlabel metal2 499 -2123 499 -2123 0 net=2843
rlabel metal2 765 -2123 765 -2123 0 net=4733
rlabel metal2 303 -2125 303 -2125 0 net=1569
rlabel metal2 492 -2125 492 -2125 0 net=1822
rlabel metal2 303 -2127 303 -2127 0 net=3015
rlabel metal2 352 -2129 352 -2129 0 net=5851
rlabel metal2 352 -2131 352 -2131 0 net=1911
rlabel metal2 373 -2133 373 -2133 0 net=9198
rlabel metal2 128 -2135 128 -2135 0 net=9681
rlabel metal2 128 -2137 128 -2137 0 net=2775
rlabel metal2 380 -2137 380 -2137 0 net=3567
rlabel metal2 401 -2139 401 -2139 0 net=2667
rlabel metal2 646 -2139 646 -2139 0 net=3855
rlabel metal2 79 -2141 79 -2141 0 net=3389
rlabel metal2 408 -2141 408 -2141 0 net=2675
rlabel metal2 674 -2141 674 -2141 0 net=7003
rlabel metal2 79 -2143 79 -2143 0 net=6539
rlabel metal2 418 -2143 418 -2143 0 net=6873
rlabel metal2 408 -2145 408 -2145 0 net=4617
rlabel metal2 429 -2147 429 -2147 0 net=2577
rlabel metal2 436 -2149 436 -2149 0 net=4893
rlabel metal2 436 -2151 436 -2151 0 net=2625
rlabel metal2 618 -2153 618 -2153 0 net=4217
rlabel metal2 618 -2155 618 -2155 0 net=6957
rlabel metal2 1045 -2157 1045 -2157 0 net=8479
rlabel metal2 1206 -2159 1206 -2159 0 net=8695
rlabel metal2 1206 -2161 1206 -2161 0 net=8623
rlabel metal2 1234 -2163 1234 -2163 0 net=10233
rlabel metal2 1402 -2165 1402 -2165 0 net=10561
rlabel metal2 1535 -2167 1535 -2167 0 net=10079
rlabel metal2 152 -2169 152 -2169 0 net=11425
rlabel metal2 51 -2180 51 -2180 0 net=1788
rlabel metal2 418 -2180 418 -2180 0 net=6027
rlabel metal2 803 -2180 803 -2180 0 net=11846
rlabel metal2 1696 -2180 1696 -2180 0 net=10990
rlabel metal2 58 -2182 58 -2182 0 net=4859
rlabel metal2 145 -2182 145 -2182 0 net=5730
rlabel metal2 940 -2182 940 -2182 0 net=6132
rlabel metal2 1125 -2182 1125 -2182 0 net=10162
rlabel metal2 1549 -2182 1549 -2182 0 net=11427
rlabel metal2 1549 -2182 1549 -2182 0 net=11427
rlabel metal2 1563 -2182 1563 -2182 0 net=11495
rlabel metal2 1563 -2182 1563 -2182 0 net=11495
rlabel metal2 1640 -2182 1640 -2182 0 net=9590
rlabel metal2 72 -2184 72 -2184 0 net=2036
rlabel metal2 660 -2184 660 -2184 0 net=5301
rlabel metal2 866 -2184 866 -2184 0 net=7338
rlabel metal2 1409 -2184 1409 -2184 0 net=10247
rlabel metal2 1650 -2184 1650 -2184 0 net=10778
rlabel metal2 1671 -2184 1671 -2184 0 net=9226
rlabel metal2 93 -2186 93 -2186 0 net=1692
rlabel metal2 317 -2186 317 -2186 0 net=1906
rlabel metal2 380 -2186 380 -2186 0 net=3568
rlabel metal2 943 -2186 943 -2186 0 net=8522
rlabel metal2 1132 -2186 1132 -2186 0 net=11834
rlabel metal2 1689 -2186 1689 -2186 0 net=4603
rlabel metal2 93 -2188 93 -2188 0 net=2189
rlabel metal2 1262 -2188 1262 -2188 0 net=9283
rlabel metal2 1696 -2188 1696 -2188 0 net=8639
rlabel metal2 100 -2190 100 -2190 0 net=489
rlabel metal2 1059 -2190 1059 -2190 0 net=7461
rlabel metal2 1087 -2190 1087 -2190 0 net=8309
rlabel metal2 1150 -2190 1150 -2190 0 net=10529
rlabel metal2 1388 -2190 1388 -2190 0 net=6672
rlabel metal2 61 -2192 61 -2192 0 net=6935
rlabel metal2 107 -2192 107 -2192 0 net=4619
rlabel metal2 492 -2192 492 -2192 0 net=2668
rlabel metal2 586 -2192 586 -2192 0 net=6124
rlabel metal2 975 -2192 975 -2192 0 net=9172
rlabel metal2 1388 -2192 1388 -2192 0 net=10455
rlabel metal2 110 -2194 110 -2194 0 net=2059
rlabel metal2 201 -2194 201 -2194 0 net=4462
rlabel metal2 499 -2194 499 -2194 0 net=2844
rlabel metal2 873 -2194 873 -2194 0 net=9150
rlabel metal2 1311 -2194 1311 -2194 0 net=10886
rlabel metal2 72 -2196 72 -2196 0 net=3957
rlabel metal2 877 -2196 877 -2196 0 net=6801
rlabel metal2 933 -2196 933 -2196 0 net=6995
rlabel metal2 999 -2196 999 -2196 0 net=7762
rlabel metal2 1150 -2196 1150 -2196 0 net=9095
rlabel metal2 114 -2198 114 -2198 0 net=1999
rlabel metal2 499 -2198 499 -2198 0 net=2975
rlabel metal2 513 -2198 513 -2198 0 net=8489
rlabel metal2 1174 -2198 1174 -2198 0 net=8854
rlabel metal2 1262 -2198 1262 -2198 0 net=9699
rlabel metal2 1409 -2198 1409 -2198 0 net=10635
rlabel metal2 1507 -2198 1507 -2198 0 net=11091
rlabel metal2 114 -2200 114 -2200 0 net=5875
rlabel metal2 618 -2200 618 -2200 0 net=6958
rlabel metal2 688 -2200 688 -2200 0 net=2434
rlabel metal2 877 -2200 877 -2200 0 net=9109
rlabel metal2 1248 -2200 1248 -2200 0 net=9423
rlabel metal2 1311 -2200 1311 -2200 0 net=10039
rlabel metal2 1353 -2200 1353 -2200 0 net=10535
rlabel metal2 1542 -2200 1542 -2200 0 net=11355
rlabel metal2 121 -2202 121 -2202 0 net=3525
rlabel metal2 506 -2202 506 -2202 0 net=3252
rlabel metal2 583 -2202 583 -2202 0 net=3559
rlabel metal2 604 -2202 604 -2202 0 net=5290
rlabel metal2 905 -2202 905 -2202 0 net=6653
rlabel metal2 975 -2202 975 -2202 0 net=7075
rlabel metal2 1066 -2202 1066 -2202 0 net=8101
rlabel metal2 1227 -2202 1227 -2202 0 net=7239
rlabel metal2 1444 -2202 1444 -2202 0 net=9081
rlabel metal2 1598 -2202 1598 -2202 0 net=11663
rlabel metal2 44 -2204 44 -2204 0 net=3953
rlabel metal2 495 -2204 495 -2204 0 net=4327
rlabel metal2 611 -2204 611 -2204 0 net=4019
rlabel metal2 660 -2204 660 -2204 0 net=6231
rlabel metal2 961 -2204 961 -2204 0 net=6875
rlabel metal2 1020 -2204 1020 -2204 0 net=9887
rlabel metal2 1318 -2204 1318 -2204 0 net=10209
rlabel metal2 1374 -2204 1374 -2204 0 net=11065
rlabel metal2 44 -2206 44 -2206 0 net=7113
rlabel metal2 128 -2206 128 -2206 0 net=1475
rlabel metal2 156 -2206 156 -2206 0 net=4287
rlabel metal2 513 -2206 513 -2206 0 net=3119
rlabel metal2 534 -2206 534 -2206 0 net=2838
rlabel metal2 618 -2206 618 -2206 0 net=3857
rlabel metal2 688 -2206 688 -2206 0 net=5716
rlabel metal2 817 -2206 817 -2206 0 net=11979
rlabel metal2 128 -2208 128 -2208 0 net=4089
rlabel metal2 691 -2208 691 -2208 0 net=4326
rlabel metal2 761 -2208 761 -2208 0 net=6534
rlabel metal2 1027 -2208 1027 -2208 0 net=8696
rlabel metal2 1314 -2208 1314 -2208 0 net=10595
rlabel metal2 1381 -2208 1381 -2208 0 net=10609
rlabel metal2 131 -2210 131 -2210 0 net=2858
rlabel metal2 156 -2210 156 -2210 0 net=4033
rlabel metal2 520 -2210 520 -2210 0 net=3361
rlabel metal2 597 -2210 597 -2210 0 net=4057
rlabel metal2 698 -2210 698 -2210 0 net=2986
rlabel metal2 807 -2210 807 -2210 0 net=5847
rlabel metal2 978 -2210 978 -2210 0 net=11888
rlabel metal2 65 -2212 65 -2212 0 net=2516
rlabel metal2 982 -2212 982 -2212 0 net=7365
rlabel metal2 1062 -2212 1062 -2212 0 net=10135
rlabel metal2 1332 -2212 1332 -2212 0 net=10355
rlabel metal2 65 -2214 65 -2214 0 net=3719
rlabel metal2 285 -2214 285 -2214 0 net=11646
rlabel metal2 124 -2216 124 -2216 0 net=10623
rlabel metal2 1528 -2216 1528 -2216 0 net=11631
rlabel metal2 138 -2218 138 -2218 0 net=7785
rlabel metal2 709 -2218 709 -2218 0 net=10483
rlabel metal2 1626 -2218 1626 -2218 0 net=12035
rlabel metal2 163 -2220 163 -2220 0 net=2685
rlabel metal2 254 -2220 254 -2220 0 net=1843
rlabel metal2 359 -2220 359 -2220 0 net=2919
rlabel metal2 394 -2220 394 -2220 0 net=3138
rlabel metal2 600 -2220 600 -2220 0 net=7943
rlabel metal2 1080 -2220 1080 -2220 0 net=8263
rlabel metal2 1381 -2220 1381 -2220 0 net=10325
rlabel metal2 163 -2222 163 -2222 0 net=4525
rlabel metal2 786 -2222 786 -2222 0 net=5589
rlabel metal2 1003 -2222 1003 -2222 0 net=7485
rlabel metal2 1108 -2222 1108 -2222 0 net=4597
rlabel metal2 1395 -2222 1395 -2222 0 net=10271
rlabel metal2 170 -2224 170 -2224 0 net=2731
rlabel metal2 464 -2224 464 -2224 0 net=4371
rlabel metal2 674 -2224 674 -2224 0 net=7005
rlabel metal2 1017 -2224 1017 -2224 0 net=10306
rlabel metal2 30 -2226 30 -2226 0 net=8899
rlabel metal2 177 -2226 177 -2226 0 net=5140
rlabel metal2 667 -2226 667 -2226 0 net=7822
rlabel metal2 1024 -2226 1024 -2226 0 net=9557
rlabel metal2 1437 -2226 1437 -2226 0 net=11105
rlabel metal2 30 -2228 30 -2228 0 net=5443
rlabel metal2 212 -2228 212 -2228 0 net=2375
rlabel metal2 296 -2228 296 -2228 0 net=1519
rlabel metal2 303 -2228 303 -2228 0 net=3016
rlabel metal2 709 -2228 709 -2228 0 net=9205
rlabel metal2 1027 -2228 1027 -2228 0 net=8852
rlabel metal2 1556 -2228 1556 -2228 0 net=10719
rlabel metal2 177 -2230 177 -2230 0 net=4455
rlabel metal2 716 -2230 716 -2230 0 net=6045
rlabel metal2 1073 -2230 1073 -2230 0 net=8833
rlabel metal2 1577 -2230 1577 -2230 0 net=11995
rlabel metal2 184 -2232 184 -2232 0 net=3323
rlabel metal2 184 -2232 184 -2232 0 net=3323
rlabel metal2 215 -2232 215 -2232 0 net=9666
rlabel metal2 1115 -2232 1115 -2232 0 net=8195
rlabel metal2 219 -2234 219 -2234 0 net=2203
rlabel metal2 219 -2234 219 -2234 0 net=2203
rlabel metal2 226 -2234 226 -2234 0 net=4986
rlabel metal2 555 -2234 555 -2234 0 net=4218
rlabel metal2 681 -2234 681 -2234 0 net=3584
rlabel metal2 737 -2234 737 -2234 0 net=7143
rlabel metal2 1115 -2234 1115 -2234 0 net=8413
rlabel metal2 1178 -2234 1178 -2234 0 net=9499
rlabel metal2 1535 -2234 1535 -2234 0 net=10081
rlabel metal2 226 -2236 226 -2236 0 net=1745
rlabel metal2 261 -2236 261 -2236 0 net=2777
rlabel metal2 394 -2236 394 -2236 0 net=2677
rlabel metal2 509 -2236 509 -2236 0 net=4655
rlabel metal2 821 -2236 821 -2236 0 net=10753
rlabel metal2 229 -2238 229 -2238 0 net=10895
rlabel metal2 233 -2240 233 -2240 0 net=5723
rlabel metal2 1143 -2240 1143 -2240 0 net=9301
rlabel metal2 1199 -2240 1199 -2240 0 net=9513
rlabel metal2 233 -2242 233 -2242 0 net=3621
rlabel metal2 989 -2242 989 -2242 0 net=7765
rlabel metal2 1206 -2242 1206 -2242 0 net=8625
rlabel metal2 240 -2244 240 -2244 0 net=1979
rlabel metal2 625 -2244 625 -2244 0 net=7934
rlabel metal2 261 -2246 261 -2246 0 net=4067
rlabel metal2 1206 -2246 1206 -2246 0 net=8355
rlabel metal2 1479 -2246 1479 -2246 0 net=10871
rlabel metal2 268 -2248 268 -2248 0 net=3189
rlabel metal2 282 -2248 282 -2248 0 net=6192
rlabel metal2 989 -2248 989 -2248 0 net=7727
rlabel metal2 1143 -2248 1143 -2248 0 net=8917
rlabel metal2 1241 -2248 1241 -2248 0 net=9050
rlabel metal2 1493 -2248 1493 -2248 0 net=11211
rlabel metal2 268 -2250 268 -2250 0 net=1859
rlabel metal2 359 -2250 359 -2250 0 net=3011
rlabel metal2 898 -2250 898 -2250 0 net=6681
rlabel metal2 996 -2250 996 -2250 0 net=11297
rlabel metal2 1276 -2250 1276 -2250 0 net=10503
rlabel metal2 1570 -2250 1570 -2250 0 net=10619
rlabel metal2 79 -2252 79 -2252 0 net=6541
rlabel metal2 401 -2252 401 -2252 0 net=3391
rlabel metal2 628 -2252 628 -2252 0 net=9837
rlabel metal2 1591 -2252 1591 -2252 0 net=11609
rlabel metal2 79 -2254 79 -2254 0 net=10594
rlabel metal2 1605 -2254 1605 -2254 0 net=11465
rlabel metal2 103 -2256 103 -2256 0 net=10889
rlabel metal2 1521 -2256 1521 -2256 0 net=11339
rlabel metal2 1605 -2256 1605 -2256 0 net=11915
rlabel metal2 250 -2258 250 -2258 0 net=5425
rlabel metal2 471 -2258 471 -2258 0 net=6569
rlabel metal2 996 -2258 996 -2258 0 net=7809
rlabel metal2 1584 -2258 1584 -2258 0 net=11553
rlabel metal2 1647 -2258 1647 -2258 0 net=5207
rlabel metal2 296 -2260 296 -2260 0 net=2579
rlabel metal2 471 -2260 471 -2260 0 net=4895
rlabel metal2 821 -2260 821 -2260 0 net=5249
rlabel metal2 929 -2260 929 -2260 0 net=10765
rlabel metal2 1619 -2260 1619 -2260 0 net=11947
rlabel metal2 257 -2262 257 -2262 0 net=5615
rlabel metal2 856 -2262 856 -2262 0 net=6259
rlabel metal2 954 -2262 954 -2262 0 net=8969
rlabel metal2 1412 -2262 1412 -2262 0 net=1
rlabel metal2 303 -2264 303 -2264 0 net=1571
rlabel metal2 534 -2264 534 -2264 0 net=4489
rlabel metal2 814 -2264 814 -2264 0 net=7707
rlabel metal2 1010 -2264 1010 -2264 0 net=2435
rlabel metal2 191 -2266 191 -2266 0 net=3629
rlabel metal2 541 -2266 541 -2266 0 net=5243
rlabel metal2 1094 -2266 1094 -2266 0 net=8779
rlabel metal2 1213 -2266 1213 -2266 0 net=9337
rlabel metal2 149 -2268 149 -2268 0 net=1939
rlabel metal2 310 -2268 310 -2268 0 net=1811
rlabel metal2 338 -2268 338 -2268 0 net=1913
rlabel metal2 548 -2268 548 -2268 0 net=3053
rlabel metal2 632 -2268 632 -2268 0 net=5181
rlabel metal2 1255 -2268 1255 -2268 0 net=9683
rlabel metal2 86 -2270 86 -2270 0 net=2519
rlabel metal2 681 -2270 681 -2270 0 net=4575
rlabel metal2 758 -2270 758 -2270 0 net=5853
rlabel metal2 1234 -2270 1234 -2270 0 net=10235
rlabel metal2 86 -2272 86 -2272 0 net=4881
rlabel metal2 705 -2272 705 -2272 0 net=8321
rlabel metal2 1234 -2272 1234 -2272 0 net=9597
rlabel metal2 152 -2274 152 -2274 0 net=2405
rlabel metal2 730 -2274 730 -2274 0 net=5127
rlabel metal2 793 -2274 793 -2274 0 net=5177
rlabel metal2 1283 -2274 1283 -2274 0 net=9399
rlabel metal2 205 -2276 205 -2276 0 net=3319
rlabel metal2 814 -2276 814 -2276 0 net=6171
rlabel metal2 1283 -2276 1283 -2276 0 net=10001
rlabel metal2 317 -2278 317 -2278 0 net=2761
rlabel metal2 527 -2278 527 -2278 0 net=4702
rlabel metal2 884 -2278 884 -2278 0 net=8481
rlabel metal2 1304 -2278 1304 -2278 0 net=10151
rlabel metal2 142 -2280 142 -2280 0 net=4311
rlabel metal2 604 -2280 604 -2280 0 net=2183
rlabel metal2 1031 -2280 1031 -2280 0 net=6841
rlabel metal2 1360 -2280 1360 -2280 0 net=10563
rlabel metal2 142 -2282 142 -2282 0 net=7835
rlabel metal2 744 -2282 744 -2282 0 net=6339
rlabel metal2 1031 -2282 1031 -2282 0 net=6241
rlabel metal2 1402 -2282 1402 -2282 0 net=11727
rlabel metal2 205 -2284 205 -2284 0 net=11869
rlabel metal2 1500 -2284 1500 -2284 0 net=10939
rlabel metal2 324 -2286 324 -2286 0 net=2508
rlabel metal2 744 -2286 744 -2286 0 net=4735
rlabel metal2 324 -2288 324 -2288 0 net=2817
rlabel metal2 765 -2288 765 -2288 0 net=5105
rlabel metal2 331 -2290 331 -2290 0 net=2627
rlabel metal2 485 -2290 485 -2290 0 net=2863
rlabel metal2 366 -2292 366 -2292 0 net=2295
rlabel metal2 436 -2292 436 -2292 0 net=3161
rlabel metal2 835 -2292 835 -2292 0 net=11323
rlabel metal2 37 -2294 37 -2294 0 net=7081
rlabel metal2 387 -2296 387 -2296 0 net=3869
rlabel metal2 450 -2298 450 -2298 0 net=6827
rlabel metal2 30 -2309 30 -2309 0 net=5444
rlabel metal2 205 -2309 205 -2309 0 net=2205
rlabel metal2 254 -2309 254 -2309 0 net=1844
rlabel metal2 548 -2309 548 -2309 0 net=2406
rlabel metal2 971 -2309 971 -2309 0 net=8780
rlabel metal2 1115 -2309 1115 -2309 0 net=8415
rlabel metal2 1115 -2309 1115 -2309 0 net=8415
rlabel metal2 1143 -2309 1143 -2309 0 net=8919
rlabel metal2 1143 -2309 1143 -2309 0 net=8919
rlabel metal2 1174 -2309 1174 -2309 0 net=11212
rlabel metal2 1514 -2309 1514 -2309 0 net=11325
rlabel metal2 1514 -2309 1514 -2309 0 net=11325
rlabel metal2 1622 -2309 1622 -2309 0 net=8640
rlabel metal2 51 -2311 51 -2311 0 net=3013
rlabel metal2 387 -2311 387 -2311 0 net=3871
rlabel metal2 576 -2311 576 -2311 0 net=5302
rlabel metal2 835 -2311 835 -2311 0 net=10484
rlabel metal2 1465 -2311 1465 -2311 0 net=11067
rlabel metal2 1465 -2311 1465 -2311 0 net=11067
rlabel metal2 1493 -2311 1493 -2311 0 net=11357
rlabel metal2 1647 -2311 1647 -2311 0 net=4604
rlabel metal2 65 -2313 65 -2313 0 net=3721
rlabel metal2 79 -2313 79 -2313 0 net=7082
rlabel metal2 597 -2313 597 -2313 0 net=2797
rlabel metal2 779 -2313 779 -2313 0 net=10236
rlabel metal2 1437 -2313 1437 -2313 0 net=11107
rlabel metal2 1437 -2313 1437 -2313 0 net=11107
rlabel metal2 1451 -2313 1451 -2313 0 net=11193
rlabel metal2 65 -2315 65 -2315 0 net=4069
rlabel metal2 285 -2315 285 -2315 0 net=1812
rlabel metal2 317 -2315 317 -2315 0 net=2762
rlabel metal2 625 -2315 625 -2315 0 net=3320
rlabel metal2 821 -2315 821 -2315 0 net=5251
rlabel metal2 859 -2315 859 -2315 0 net=10624
rlabel metal2 1542 -2315 1542 -2315 0 net=11555
rlabel metal2 79 -2317 79 -2317 0 net=5427
rlabel metal2 415 -2317 415 -2317 0 net=2732
rlabel metal2 635 -2317 635 -2317 0 net=4565
rlabel metal2 677 -2317 677 -2317 0 net=5128
rlabel metal2 740 -2317 740 -2317 0 net=8196
rlabel metal2 128 -2319 128 -2319 0 net=4090
rlabel metal2 705 -2319 705 -2319 0 net=5848
rlabel metal2 866 -2319 866 -2319 0 net=9424
rlabel metal2 1251 -2319 1251 -2319 0 net=9400
rlabel metal2 1346 -2319 1346 -2319 0 net=10597
rlabel metal2 1430 -2319 1430 -2319 0 net=10891
rlabel metal2 1612 -2319 1612 -2319 0 net=11467
rlabel metal2 114 -2321 114 -2321 0 net=5877
rlabel metal2 873 -2321 873 -2321 0 net=10152
rlabel metal2 1311 -2321 1311 -2321 0 net=10041
rlabel metal2 1311 -2321 1311 -2321 0 net=10041
rlabel metal2 1374 -2321 1374 -2321 0 net=10273
rlabel metal2 1444 -2321 1444 -2321 0 net=9083
rlabel metal2 1612 -2321 1612 -2321 0 net=11981
rlabel metal2 114 -2323 114 -2323 0 net=4288
rlabel metal2 450 -2323 450 -2323 0 net=5724
rlabel metal2 1171 -2323 1171 -2323 0 net=6593
rlabel metal2 135 -2325 135 -2325 0 net=5245
rlabel metal2 562 -2325 562 -2325 0 net=5178
rlabel metal2 912 -2325 912 -2325 0 net=9514
rlabel metal2 1444 -2325 1444 -2325 0 net=10897
rlabel metal2 149 -2327 149 -2327 0 net=8103
rlabel metal2 1073 -2327 1073 -2327 0 net=8835
rlabel metal2 1164 -2327 1164 -2327 0 net=9303
rlabel metal2 1199 -2327 1199 -2327 0 net=8626
rlabel metal2 208 -2329 208 -2329 0 net=4372
rlabel metal2 492 -2329 492 -2329 0 net=1160
rlabel metal2 1052 -2329 1052 -2329 0 net=7945
rlabel metal2 1129 -2329 1129 -2329 0 net=11871
rlabel metal2 215 -2331 215 -2331 0 net=2818
rlabel metal2 359 -2331 359 -2331 0 net=4491
rlabel metal2 541 -2331 541 -2331 0 net=3393
rlabel metal2 579 -2331 579 -2331 0 net=8153
rlabel metal2 1073 -2331 1073 -2331 0 net=8265
rlabel metal2 1087 -2331 1087 -2331 0 net=8311
rlabel metal2 1087 -2331 1087 -2331 0 net=8311
rlabel metal2 1122 -2331 1122 -2331 0 net=8491
rlabel metal2 1157 -2331 1157 -2331 0 net=7767
rlabel metal2 1202 -2331 1202 -2331 0 net=10326
rlabel metal2 1472 -2331 1472 -2331 0 net=11093
rlabel metal2 1535 -2331 1535 -2331 0 net=11611
rlabel metal2 86 -2333 86 -2333 0 net=4883
rlabel metal2 590 -2333 590 -2333 0 net=4329
rlabel metal2 639 -2333 639 -2333 0 net=5854
rlabel metal2 891 -2333 891 -2333 0 net=6683
rlabel metal2 912 -2333 912 -2333 0 net=5407
rlabel metal2 1591 -2333 1591 -2333 0 net=11917
rlabel metal2 72 -2335 72 -2335 0 net=3959
rlabel metal2 639 -2335 639 -2335 0 net=4577
rlabel metal2 684 -2335 684 -2335 0 net=7039
rlabel metal2 842 -2335 842 -2335 0 net=6655
rlabel metal2 915 -2335 915 -2335 0 net=10610
rlabel metal2 1605 -2335 1605 -2335 0 net=11977
rlabel metal2 72 -2337 72 -2337 0 net=5183
rlabel metal2 667 -2337 667 -2337 0 net=6261
rlabel metal2 919 -2337 919 -2337 0 net=6046
rlabel metal2 919 -2337 919 -2337 0 net=6046
rlabel metal2 989 -2337 989 -2337 0 net=7729
rlabel metal2 1017 -2337 1017 -2337 0 net=4598
rlabel metal2 1122 -2337 1122 -2337 0 net=11996
rlabel metal2 86 -2339 86 -2339 0 net=5043
rlabel metal2 233 -2339 233 -2339 0 net=3623
rlabel metal2 261 -2339 261 -2339 0 net=3191
rlabel metal2 289 -2339 289 -2339 0 net=2377
rlabel metal2 436 -2339 436 -2339 0 net=3163
rlabel metal2 495 -2339 495 -2339 0 net=4058
rlabel metal2 681 -2339 681 -2339 0 net=10087
rlabel metal2 1185 -2339 1185 -2339 0 net=11299
rlabel metal2 117 -2341 117 -2341 0 net=2845
rlabel metal2 296 -2341 296 -2341 0 net=2581
rlabel metal2 632 -2341 632 -2341 0 net=8970
rlabel metal2 975 -2341 975 -2341 0 net=7077
rlabel metal2 1185 -2341 1185 -2341 0 net=10210
rlabel metal2 142 -2343 142 -2343 0 net=3547
rlabel metal2 247 -2343 247 -2343 0 net=2687
rlabel metal2 373 -2343 373 -2343 0 net=2779
rlabel metal2 478 -2343 478 -2343 0 net=6829
rlabel metal2 975 -2343 975 -2343 0 net=7367
rlabel metal2 989 -2343 989 -2343 0 net=7487
rlabel metal2 1020 -2343 1020 -2343 0 net=7462
rlabel metal2 1206 -2343 1206 -2343 0 net=8356
rlabel metal2 1248 -2343 1248 -2343 0 net=12036
rlabel metal2 142 -2345 142 -2345 0 net=1981
rlabel metal2 247 -2345 247 -2345 0 net=2629
rlabel metal2 373 -2345 373 -2345 0 net=2185
rlabel metal2 688 -2345 688 -2345 0 net=5590
rlabel metal2 849 -2345 849 -2345 0 net=7007
rlabel metal2 1003 -2345 1003 -2345 0 net=6243
rlabel metal2 1038 -2345 1038 -2345 0 net=10456
rlabel metal2 1570 -2345 1570 -2345 0 net=10621
rlabel metal2 170 -2347 170 -2347 0 net=8901
rlabel metal2 282 -2347 282 -2347 0 net=6983
rlabel metal2 996 -2347 996 -2347 0 net=7811
rlabel metal2 1045 -2347 1045 -2347 0 net=6843
rlabel metal2 1206 -2347 1206 -2347 0 net=8525
rlabel metal2 1367 -2347 1367 -2347 0 net=10941
rlabel metal2 170 -2349 170 -2349 0 net=1941
rlabel metal2 219 -2349 219 -2349 0 net=1747
rlabel metal2 240 -2349 240 -2349 0 net=2297
rlabel metal2 380 -2349 380 -2349 0 net=2920
rlabel metal2 422 -2349 422 -2349 0 net=2000
rlabel metal2 691 -2349 691 -2349 0 net=5807
rlabel metal2 786 -2349 786 -2349 0 net=3659
rlabel metal2 184 -2351 184 -2351 0 net=3325
rlabel metal2 226 -2351 226 -2351 0 net=6570
rlabel metal2 1059 -2351 1059 -2351 0 net=7241
rlabel metal2 1237 -2351 1237 -2351 0 net=10248
rlabel metal2 184 -2353 184 -2353 0 net=2865
rlabel metal2 499 -2353 499 -2353 0 net=2977
rlabel metal2 499 -2353 499 -2353 0 net=2977
rlabel metal2 506 -2353 506 -2353 0 net=4751
rlabel metal2 709 -2353 709 -2353 0 net=9207
rlabel metal2 1150 -2353 1150 -2353 0 net=9097
rlabel metal2 1241 -2353 1241 -2353 0 net=10872
rlabel metal2 1486 -2353 1486 -2353 0 net=11231
rlabel metal2 268 -2355 268 -2355 0 net=1861
rlabel metal2 422 -2355 422 -2355 0 net=3955
rlabel metal2 506 -2355 506 -2355 0 net=3055
rlabel metal2 604 -2355 604 -2355 0 net=4021
rlabel metal2 621 -2355 621 -2355 0 net=11445
rlabel metal2 1650 -2355 1650 -2355 0 net=10082
rlabel metal2 268 -2357 268 -2357 0 net=5865
rlabel metal2 838 -2357 838 -2357 0 net=11743
rlabel metal2 1661 -2357 1661 -2357 0 net=9285
rlabel metal2 282 -2359 282 -2359 0 net=11303
rlabel metal2 296 -2361 296 -2361 0 net=1915
rlabel metal2 345 -2361 345 -2361 0 net=6543
rlabel metal2 695 -2361 695 -2361 0 net=9110
rlabel metal2 947 -2361 947 -2361 0 net=7709
rlabel metal2 1150 -2361 1150 -2361 0 net=8371
rlabel metal2 1388 -2361 1388 -2361 0 net=10637
rlabel metal2 100 -2363 100 -2363 0 net=6937
rlabel metal2 709 -2363 709 -2363 0 net=6341
rlabel metal2 800 -2363 800 -2363 0 net=6029
rlabel metal2 947 -2363 947 -2363 0 net=6877
rlabel metal2 992 -2363 992 -2363 0 net=1
rlabel metal2 1220 -2363 1220 -2363 0 net=9559
rlabel metal2 1220 -2363 1220 -2363 0 net=9559
rlabel metal2 1241 -2363 1241 -2363 0 net=9889
rlabel metal2 1318 -2363 1318 -2363 0 net=10137
rlabel metal2 100 -2365 100 -2365 0 net=6173
rlabel metal2 870 -2365 870 -2365 0 net=9455
rlabel metal2 1318 -2365 1318 -2365 0 net=10357
rlabel metal2 1339 -2365 1339 -2365 0 net=10531
rlabel metal2 303 -2367 303 -2367 0 net=1573
rlabel metal2 303 -2367 303 -2367 0 net=1573
rlabel metal2 310 -2367 310 -2367 0 net=4897
rlabel metal2 509 -2367 509 -2367 0 net=3120
rlabel metal2 534 -2367 534 -2367 0 net=2939
rlabel metal2 1269 -2367 1269 -2367 0 net=9839
rlabel metal2 1332 -2367 1332 -2367 0 net=10537
rlabel metal2 58 -2369 58 -2369 0 net=4861
rlabel metal2 611 -2369 611 -2369 0 net=6889
rlabel metal2 870 -2369 870 -2369 0 net=6459
rlabel metal2 1255 -2369 1255 -2369 0 net=9685
rlabel metal2 1283 -2369 1283 -2369 0 net=10003
rlabel metal2 1339 -2369 1339 -2369 0 net=10565
rlabel metal2 44 -2371 44 -2371 0 net=7115
rlabel metal2 317 -2371 317 -2371 0 net=1645
rlabel metal2 716 -2371 716 -2371 0 net=4657
rlabel metal2 926 -2371 926 -2371 0 net=6803
rlabel metal2 1234 -2371 1234 -2371 0 net=9599
rlabel metal2 1262 -2371 1262 -2371 0 net=9701
rlabel metal2 1290 -2371 1290 -2371 0 net=11632
rlabel metal2 44 -2373 44 -2373 0 net=9059
rlabel metal2 898 -2373 898 -2373 0 net=6523
rlabel metal2 1017 -2373 1017 -2373 0 net=7307
rlabel metal2 1353 -2373 1353 -2373 0 net=10755
rlabel metal2 1528 -2373 1528 -2373 0 net=11429
rlabel metal2 331 -2375 331 -2375 0 net=4933
rlabel metal2 653 -2375 653 -2375 0 net=7787
rlabel metal2 1192 -2375 1192 -2375 0 net=10767
rlabel metal2 1549 -2375 1549 -2375 0 net=10721
rlabel metal2 107 -2377 107 -2377 0 net=4621
rlabel metal2 660 -2377 660 -2377 0 net=6233
rlabel metal2 1178 -2377 1178 -2377 0 net=9501
rlabel metal2 1213 -2377 1213 -2377 0 net=9339
rlabel metal2 1402 -2377 1402 -2377 0 net=11729
rlabel metal2 138 -2379 138 -2379 0 net=9401
rlabel metal2 1213 -2379 1213 -2379 0 net=11341
rlabel metal2 163 -2381 163 -2381 0 net=4527
rlabel metal2 723 -2381 723 -2381 0 net=7837
rlabel metal2 1276 -2381 1276 -2381 0 net=10505
rlabel metal2 1521 -2381 1521 -2381 0 net=11497
rlabel metal2 163 -2383 163 -2383 0 net=1521
rlabel metal2 436 -2383 436 -2383 0 net=3363
rlabel metal2 583 -2383 583 -2383 0 net=3561
rlabel metal2 723 -2383 723 -2383 0 net=5209
rlabel metal2 338 -2385 338 -2385 0 net=2521
rlabel metal2 366 -2385 366 -2385 0 net=4313
rlabel metal2 730 -2385 730 -2385 0 net=8482
rlabel metal2 1202 -2385 1202 -2385 0 net=12087
rlabel metal2 1563 -2385 1563 -2385 0 net=11665
rlabel metal2 156 -2387 156 -2387 0 net=4035
rlabel metal2 380 -2387 380 -2387 0 net=8697
rlabel metal2 1598 -2387 1598 -2387 0 net=11949
rlabel metal2 156 -2389 156 -2389 0 net=10097
rlabel metal2 747 -2389 747 -2389 0 net=10473
rlabel metal2 345 -2391 345 -2391 0 net=7377
rlabel metal2 751 -2391 751 -2391 0 net=9519
rlabel metal2 387 -2393 387 -2393 0 net=2679
rlabel metal2 404 -2393 404 -2393 0 net=2537
rlabel metal2 443 -2393 443 -2393 0 net=3631
rlabel metal2 520 -2393 520 -2393 0 net=10275
rlabel metal2 744 -2393 744 -2393 0 net=4737
rlabel metal2 128 -2395 128 -2395 0 net=6193
rlabel metal2 758 -2395 758 -2395 0 net=6487
rlabel metal2 443 -2397 443 -2397 0 net=1921
rlabel metal2 450 -2399 450 -2399 0 net=2303
rlabel metal2 453 -2401 453 -2401 0 net=7144
rlabel metal2 758 -2401 758 -2401 0 net=5107
rlabel metal2 775 -2401 775 -2401 0 net=11733
rlabel metal2 394 -2403 394 -2403 0 net=5007
rlabel metal2 765 -2403 765 -2403 0 net=5617
rlabel metal2 933 -2403 933 -2403 0 net=6997
rlabel metal2 457 -2405 457 -2405 0 net=2437
rlabel metal2 471 -2407 471 -2407 0 net=3859
rlabel metal2 642 -2407 642 -2407 0 net=7993
rlabel metal2 1010 -2407 1010 -2407 0 net=8323
rlabel metal2 121 -2409 121 -2409 0 net=3526
rlabel metal2 121 -2411 121 -2411 0 net=7693
rlabel metal2 527 -2411 527 -2411 0 net=9291
rlabel metal2 198 -2413 198 -2413 0 net=2061
rlabel metal2 93 -2415 93 -2415 0 net=2191
rlabel metal2 93 -2417 93 -2417 0 net=4457
rlabel metal2 152 -2419 152 -2419 0 net=1587
rlabel metal2 44 -2430 44 -2430 0 net=9060
rlabel metal2 562 -2430 562 -2430 0 net=10474
rlabel metal2 1444 -2430 1444 -2430 0 net=10899
rlabel metal2 1444 -2430 1444 -2430 0 net=10899
rlabel metal2 1500 -2430 1500 -2430 0 net=11447
rlabel metal2 1500 -2430 1500 -2430 0 net=11447
rlabel metal2 1615 -2430 1615 -2430 0 net=11468
rlabel metal2 93 -2432 93 -2432 0 net=4458
rlabel metal2 121 -2432 121 -2432 0 net=7694
rlabel metal2 831 -2432 831 -2432 0 net=11342
rlabel metal2 1234 -2432 1234 -2432 0 net=9775
rlabel metal2 1622 -2432 1622 -2432 0 net=9286
rlabel metal2 93 -2434 93 -2434 0 net=1923
rlabel metal2 471 -2434 471 -2434 0 net=3860
rlabel metal2 674 -2434 674 -2434 0 net=4566
rlabel metal2 747 -2434 747 -2434 0 net=11734
rlabel metal2 1626 -2434 1626 -2434 0 net=10622
rlabel metal2 107 -2436 107 -2436 0 net=11326
rlabel metal2 1577 -2436 1577 -2436 0 net=11873
rlabel metal2 107 -2438 107 -2438 0 net=1823
rlabel metal2 121 -2438 121 -2438 0 net=5211
rlabel metal2 737 -2438 737 -2438 0 net=9098
rlabel metal2 1248 -2438 1248 -2438 0 net=11978
rlabel metal2 135 -2440 135 -2440 0 net=5246
rlabel metal2 674 -2440 674 -2440 0 net=2737
rlabel metal2 1066 -2440 1066 -2440 0 net=7839
rlabel metal2 1185 -2440 1185 -2440 0 net=8935
rlabel metal2 1251 -2440 1251 -2440 0 net=10532
rlabel metal2 1549 -2440 1549 -2440 0 net=10723
rlabel metal2 135 -2442 135 -2442 0 net=2439
rlabel metal2 520 -2442 520 -2442 0 net=4528
rlabel metal2 681 -2442 681 -2442 0 net=4738
rlabel metal2 901 -2442 901 -2442 0 net=7368
rlabel metal2 989 -2442 989 -2442 0 net=7489
rlabel metal2 1104 -2442 1104 -2442 0 net=9340
rlabel metal2 1290 -2442 1290 -2442 0 net=10138
rlabel metal2 1549 -2442 1549 -2442 0 net=11745
rlabel metal2 142 -2444 142 -2444 0 net=1982
rlabel metal2 572 -2444 572 -2444 0 net=3562
rlabel metal2 723 -2444 723 -2444 0 net=5079
rlabel metal2 1199 -2444 1199 -2444 0 net=11108
rlabel metal2 142 -2446 142 -2446 0 net=2681
rlabel metal2 394 -2446 394 -2446 0 net=5009
rlabel metal2 569 -2446 569 -2446 0 net=4885
rlabel metal2 733 -2446 733 -2446 0 net=12037
rlabel metal2 163 -2448 163 -2448 0 net=1522
rlabel metal2 821 -2448 821 -2448 0 net=7041
rlabel metal2 1013 -2448 1013 -2448 0 net=11430
rlabel metal2 163 -2450 163 -2450 0 net=2047
rlabel metal2 394 -2450 394 -2450 0 net=2149
rlabel metal2 639 -2450 639 -2450 0 net=4579
rlabel metal2 681 -2450 681 -2450 0 net=2085
rlabel metal2 688 -2450 688 -2450 0 net=6544
rlabel metal2 821 -2450 821 -2450 0 net=3807
rlabel metal2 1493 -2450 1493 -2450 0 net=11359
rlabel metal2 170 -2452 170 -2452 0 net=1942
rlabel metal2 282 -2452 282 -2452 0 net=669
rlabel metal2 835 -2452 835 -2452 0 net=9208
rlabel metal2 1115 -2452 1115 -2452 0 net=8417
rlabel metal2 1115 -2452 1115 -2452 0 net=8417
rlabel metal2 1164 -2452 1164 -2452 0 net=7769
rlabel metal2 1220 -2452 1220 -2452 0 net=9561
rlabel metal2 1332 -2452 1332 -2452 0 net=10539
rlabel metal2 1486 -2452 1486 -2452 0 net=11233
rlabel metal2 51 -2454 51 -2454 0 net=3014
rlabel metal2 219 -2454 219 -2454 0 net=1749
rlabel metal2 229 -2454 229 -2454 0 net=227
rlabel metal2 51 -2456 51 -2456 0 net=8061
rlabel metal2 404 -2456 404 -2456 0 net=2538
rlabel metal2 583 -2456 583 -2456 0 net=11213
rlabel metal2 114 -2458 114 -2458 0 net=2095
rlabel metal2 240 -2458 240 -2458 0 net=2299
rlabel metal2 583 -2458 583 -2458 0 net=6343
rlabel metal2 740 -2458 740 -2458 0 net=6656
rlabel metal2 849 -2458 849 -2458 0 net=9456
rlabel metal2 1339 -2458 1339 -2458 0 net=10567
rlabel metal2 58 -2460 58 -2460 0 net=7117
rlabel metal2 128 -2460 128 -2460 0 net=6195
rlabel metal2 849 -2460 849 -2460 0 net=6031
rlabel metal2 919 -2460 919 -2460 0 net=9840
rlabel metal2 1346 -2460 1346 -2460 0 net=10599
rlabel metal2 58 -2462 58 -2462 0 net=7433
rlabel metal2 303 -2462 303 -2462 0 net=1574
rlabel metal2 758 -2462 758 -2462 0 net=5109
rlabel metal2 828 -2462 828 -2462 0 net=5253
rlabel metal2 852 -2462 852 -2462 0 net=7078
rlabel metal2 1192 -2462 1192 -2462 0 net=9503
rlabel metal2 1318 -2462 1318 -2462 0 net=10359
rlabel metal2 1353 -2462 1353 -2462 0 net=10757
rlabel metal2 79 -2464 79 -2464 0 net=5429
rlabel metal2 856 -2464 856 -2464 0 net=11747
rlabel metal2 79 -2466 79 -2466 0 net=2631
rlabel metal2 254 -2466 254 -2466 0 net=3624
rlabel metal2 303 -2466 303 -2466 0 net=3347
rlabel metal2 1143 -2466 1143 -2466 0 net=8921
rlabel metal2 1206 -2466 1206 -2466 0 net=8527
rlabel metal2 1360 -2466 1360 -2466 0 net=11666
rlabel metal2 247 -2468 247 -2468 0 net=3633
rlabel metal2 576 -2468 576 -2468 0 net=2582
rlabel metal2 793 -2468 793 -2468 0 net=6891
rlabel metal2 929 -2468 929 -2468 0 net=10506
rlabel metal2 1563 -2468 1563 -2468 0 net=11983
rlabel metal2 254 -2470 254 -2470 0 net=1203
rlabel metal2 933 -2470 933 -2470 0 net=7995
rlabel metal2 1171 -2470 1171 -2470 0 net=9305
rlabel metal2 1374 -2470 1374 -2470 0 net=10274
rlabel metal2 1384 -2470 1384 -2470 0 net=11918
rlabel metal2 338 -2472 338 -2472 0 net=2523
rlabel metal2 523 -2472 523 -2472 0 net=2943
rlabel metal2 586 -2472 586 -2472 0 net=9051
rlabel metal2 1241 -2472 1241 -2472 0 net=9891
rlabel metal2 324 -2474 324 -2474 0 net=2689
rlabel metal2 359 -2474 359 -2474 0 net=4492
rlabel metal2 590 -2474 590 -2474 0 net=3961
rlabel metal2 590 -2474 590 -2474 0 net=3961
rlabel metal2 600 -2474 600 -2474 0 net=6804
rlabel metal2 1024 -2474 1024 -2474 0 net=7789
rlabel metal2 1150 -2474 1150 -2474 0 net=8373
rlabel metal2 1202 -2474 1202 -2474 0 net=8641
rlabel metal2 1251 -2474 1251 -2474 0 net=9357
rlabel metal2 1269 -2474 1269 -2474 0 net=9687
rlabel metal2 233 -2476 233 -2476 0 net=3549
rlabel metal2 359 -2476 359 -2476 0 net=2781
rlabel metal2 604 -2476 604 -2476 0 net=4023
rlabel metal2 667 -2476 667 -2476 0 net=6263
rlabel metal2 905 -2476 905 -2476 0 net=6831
rlabel metal2 1024 -2476 1024 -2476 0 net=11300
rlabel metal2 233 -2478 233 -2478 0 net=2187
rlabel metal2 380 -2478 380 -2478 0 net=8699
rlabel metal2 898 -2478 898 -2478 0 net=6525
rlabel metal2 940 -2478 940 -2478 0 net=6999
rlabel metal2 940 -2478 940 -2478 0 net=6999
rlabel metal2 947 -2478 947 -2478 0 net=6879
rlabel metal2 1038 -2478 1038 -2478 0 net=7711
rlabel metal2 1206 -2478 1206 -2478 0 net=7735
rlabel metal2 296 -2480 296 -2480 0 net=1917
rlabel metal2 380 -2480 380 -2480 0 net=4753
rlabel metal2 709 -2480 709 -2480 0 net=5619
rlabel metal2 793 -2480 793 -2480 0 net=4659
rlabel metal2 828 -2480 828 -2480 0 net=10163
rlabel metal2 1507 -2480 1507 -2480 0 net=11613
rlabel metal2 1640 -2480 1640 -2480 0 net=6595
rlabel metal2 173 -2482 173 -2482 0 net=867
rlabel metal2 366 -2482 366 -2482 0 net=4314
rlabel metal2 618 -2482 618 -2482 0 net=6629
rlabel metal2 947 -2482 947 -2482 0 net=7947
rlabel metal2 1178 -2482 1178 -2482 0 net=9403
rlabel metal2 1276 -2482 1276 -2482 0 net=12089
rlabel metal2 366 -2484 366 -2484 0 net=2979
rlabel metal2 618 -2484 618 -2484 0 net=4331
rlabel metal2 639 -2484 639 -2484 0 net=4637
rlabel metal2 891 -2484 891 -2484 0 net=6685
rlabel metal2 1283 -2484 1283 -2484 0 net=9703
rlabel metal2 1535 -2484 1535 -2484 0 net=11731
rlabel metal2 401 -2486 401 -2486 0 net=3365
rlabel metal2 464 -2486 464 -2486 0 net=4623
rlabel metal2 695 -2486 695 -2486 0 net=6939
rlabel metal2 996 -2486 996 -2486 0 net=7731
rlabel metal2 1045 -2486 1045 -2486 0 net=8313
rlabel metal2 1129 -2486 1129 -2486 0 net=8493
rlabel metal2 1220 -2486 1220 -2486 0 net=7823
rlabel metal2 1304 -2486 1304 -2486 0 net=10005
rlabel metal2 1556 -2486 1556 -2486 0 net=11951
rlabel metal2 128 -2488 128 -2488 0 net=2037
rlabel metal2 1052 -2488 1052 -2488 0 net=8155
rlabel metal2 1304 -2488 1304 -2488 0 net=10043
rlabel metal2 1458 -2488 1458 -2488 0 net=9085
rlabel metal2 408 -2490 408 -2490 0 net=2379
rlabel metal2 485 -2490 485 -2490 0 net=3723
rlabel metal2 621 -2490 621 -2490 0 net=4663
rlabel metal2 702 -2490 702 -2490 0 net=5879
rlabel metal2 870 -2490 870 -2490 0 net=6461
rlabel metal2 926 -2490 926 -2490 0 net=6645
rlabel metal2 1146 -2490 1146 -2490 0 net=10997
rlabel metal2 65 -2492 65 -2492 0 net=4071
rlabel metal2 499 -2492 499 -2492 0 net=3395
rlabel metal2 569 -2492 569 -2492 0 net=8029
rlabel metal2 1255 -2492 1255 -2492 0 net=9601
rlabel metal2 65 -2494 65 -2494 0 net=6607
rlabel metal2 310 -2496 310 -2496 0 net=4899
rlabel metal2 436 -2496 436 -2496 0 net=2305
rlabel metal2 513 -2496 513 -2496 0 net=4863
rlabel metal2 737 -2496 737 -2496 0 net=1335
rlabel metal2 198 -2498 198 -2498 0 net=2193
rlabel metal2 352 -2498 352 -2498 0 net=4036
rlabel metal2 611 -2498 611 -2498 0 net=9189
rlabel metal2 89 -2500 89 -2500 0 net=5401
rlabel metal2 450 -2500 450 -2500 0 net=7985
rlabel metal2 625 -2500 625 -2500 0 net=5409
rlabel metal2 1052 -2500 1052 -2500 0 net=6845
rlabel metal2 198 -2502 198 -2502 0 net=2207
rlabel metal2 492 -2502 492 -2502 0 net=3165
rlabel metal2 527 -2502 527 -2502 0 net=9293
rlabel metal2 205 -2504 205 -2504 0 net=2063
rlabel metal2 345 -2504 345 -2504 0 net=7378
rlabel metal2 548 -2504 548 -2504 0 net=3873
rlabel metal2 649 -2504 649 -2504 0 net=10107
rlabel metal2 212 -2506 212 -2506 0 net=8902
rlabel metal2 289 -2506 289 -2506 0 net=2847
rlabel metal2 492 -2506 492 -2506 0 net=3661
rlabel metal2 800 -2506 800 -2506 0 net=11194
rlabel metal2 240 -2508 240 -2508 0 net=6085
rlabel metal2 548 -2508 548 -2508 0 net=2799
rlabel metal2 653 -2508 653 -2508 0 net=5809
rlabel metal2 807 -2508 807 -2508 0 net=11556
rlabel metal2 275 -2510 275 -2510 0 net=3956
rlabel metal2 506 -2510 506 -2510 0 net=3056
rlabel metal2 744 -2510 744 -2510 0 net=7841
rlabel metal2 1367 -2510 1367 -2510 0 net=10943
rlabel metal2 1521 -2510 1521 -2510 0 net=11499
rlabel metal2 86 -2512 86 -2512 0 net=5045
rlabel metal2 565 -2512 565 -2512 0 net=4709
rlabel metal2 765 -2512 765 -2512 0 net=5085
rlabel metal2 86 -2514 86 -2514 0 net=3007
rlabel metal2 779 -2514 779 -2514 0 net=4779
rlabel metal2 1479 -2514 1479 -2514 0 net=11305
rlabel metal2 156 -2516 156 -2516 0 net=10099
rlabel metal2 814 -2516 814 -2516 0 net=6235
rlabel metal2 884 -2516 884 -2516 0 net=6489
rlabel metal2 1010 -2516 1010 -2516 0 net=8325
rlabel metal2 1157 -2516 1157 -2516 0 net=10089
rlabel metal2 1472 -2516 1472 -2516 0 net=11095
rlabel metal2 100 -2518 100 -2518 0 net=6175
rlabel metal2 268 -2518 268 -2518 0 net=5867
rlabel metal2 884 -2518 884 -2518 0 net=6245
rlabel metal2 1073 -2518 1073 -2518 0 net=8267
rlabel metal2 1465 -2518 1465 -2518 0 net=11069
rlabel metal2 100 -2520 100 -2520 0 net=4935
rlabel metal2 534 -2520 534 -2520 0 net=2940
rlabel metal2 1073 -2520 1073 -2520 0 net=8837
rlabel metal2 1430 -2520 1430 -2520 0 net=10893
rlabel metal2 72 -2522 72 -2522 0 net=5185
rlabel metal2 786 -2522 786 -2522 0 net=8175
rlabel metal2 1423 -2522 1423 -2522 0 net=10769
rlabel metal2 72 -2524 72 -2524 0 net=3193
rlabel metal2 331 -2524 331 -2524 0 net=1863
rlabel metal2 912 -2524 912 -2524 0 net=6985
rlabel metal2 968 -2524 968 -2524 0 net=7145
rlabel metal2 1388 -2524 1388 -2524 0 net=10639
rlabel metal2 149 -2526 149 -2526 0 net=8105
rlabel metal2 149 -2528 149 -2528 0 net=3327
rlabel metal2 261 -2528 261 -2528 0 net=1647
rlabel metal2 555 -2528 555 -2528 0 net=10277
rlabel metal2 184 -2530 184 -2530 0 net=2867
rlabel metal2 278 -2530 278 -2530 0 net=4561
rlabel metal2 751 -2530 751 -2530 0 net=9521
rlabel metal2 968 -2530 968 -2530 0 net=7009
rlabel metal2 177 -2532 177 -2532 0 net=1589
rlabel metal2 191 -2532 191 -2532 0 net=2231
rlabel metal2 982 -2532 982 -2532 0 net=7309
rlabel metal2 177 -2534 177 -2534 0 net=1529
rlabel metal2 317 -2534 317 -2534 0 net=2079
rlabel metal2 1017 -2534 1017 -2534 0 net=7243
rlabel metal2 1031 -2536 1031 -2536 0 net=7813
rlabel metal2 971 -2538 971 -2538 0 net=7279
rlabel metal2 44 -2549 44 -2549 0 net=3349
rlabel metal2 387 -2549 387 -2549 0 net=4639
rlabel metal2 656 -2549 656 -2549 0 net=11746
rlabel metal2 1556 -2549 1556 -2549 0 net=11953
rlabel metal2 1584 -2549 1584 -2549 0 net=10724
rlabel metal2 1629 -2549 1629 -2549 0 net=6596
rlabel metal2 72 -2551 72 -2551 0 net=3194
rlabel metal2 303 -2551 303 -2551 0 net=2701
rlabel metal2 429 -2551 429 -2551 0 net=2301
rlabel metal2 429 -2551 429 -2551 0 net=2301
rlabel metal2 457 -2551 457 -2551 0 net=2525
rlabel metal2 527 -2551 527 -2551 0 net=2087
rlabel metal2 730 -2551 730 -2551 0 net=10894
rlabel metal2 1472 -2551 1472 -2551 0 net=11071
rlabel metal2 1556 -2551 1556 -2551 0 net=11847
rlabel metal2 72 -2553 72 -2553 0 net=4333
rlabel metal2 625 -2553 625 -2553 0 net=5411
rlabel metal2 849 -2553 849 -2553 0 net=6032
rlabel metal2 950 -2553 950 -2553 0 net=11096
rlabel metal2 1514 -2553 1514 -2553 0 net=11749
rlabel metal2 1591 -2553 1591 -2553 0 net=12091
rlabel metal2 86 -2555 86 -2555 0 net=695
rlabel metal2 212 -2555 212 -2555 0 net=4193
rlabel metal2 352 -2555 352 -2555 0 net=5403
rlabel metal2 737 -2555 737 -2555 0 net=11214
rlabel metal2 86 -2557 86 -2557 0 net=4581
rlabel metal2 737 -2557 737 -2557 0 net=4653
rlabel metal2 971 -2557 971 -2557 0 net=7840
rlabel metal2 1143 -2557 1143 -2557 0 net=10360
rlabel metal2 1405 -2557 1405 -2557 0 net=11500
rlabel metal2 1598 -2557 1598 -2557 0 net=9086
rlabel metal2 93 -2559 93 -2559 0 net=1925
rlabel metal2 233 -2559 233 -2559 0 net=2188
rlabel metal2 744 -2559 744 -2559 0 net=7790
rlabel metal2 1136 -2559 1136 -2559 0 net=8107
rlabel metal2 1188 -2559 1188 -2559 0 net=10770
rlabel metal2 1444 -2559 1444 -2559 0 net=10901
rlabel metal2 1507 -2559 1507 -2559 0 net=11615
rlabel metal2 1577 -2559 1577 -2559 0 net=11875
rlabel metal2 93 -2561 93 -2561 0 net=4133
rlabel metal2 534 -2561 534 -2561 0 net=5186
rlabel metal2 789 -2561 789 -2561 0 net=6686
rlabel metal2 1304 -2561 1304 -2561 0 net=10045
rlabel metal2 1409 -2561 1409 -2561 0 net=10569
rlabel metal2 121 -2563 121 -2563 0 net=5212
rlabel metal2 835 -2563 835 -2563 0 net=6197
rlabel metal2 887 -2563 887 -2563 0 net=9504
rlabel metal2 1304 -2563 1304 -2563 0 net=10759
rlabel metal2 1458 -2563 1458 -2563 0 net=10999
rlabel metal2 65 -2565 65 -2565 0 net=6609
rlabel metal2 135 -2565 135 -2565 0 net=2440
rlabel metal2 901 -2565 901 -2565 0 net=7490
rlabel metal2 1073 -2565 1073 -2565 0 net=8839
rlabel metal2 65 -2567 65 -2567 0 net=4937
rlabel metal2 135 -2567 135 -2567 0 net=1531
rlabel metal2 201 -2567 201 -2567 0 net=10327
rlabel metal2 100 -2569 100 -2569 0 net=1825
rlabel metal2 142 -2569 142 -2569 0 net=2682
rlabel metal2 422 -2569 422 -2569 0 net=10100
rlabel metal2 667 -2569 667 -2569 0 net=4887
rlabel metal2 730 -2569 730 -2569 0 net=1605
rlabel metal2 758 -2569 758 -2569 0 net=5431
rlabel metal2 954 -2569 954 -2569 0 net=9523
rlabel metal2 1388 -2569 1388 -2569 0 net=10279
rlabel metal2 107 -2571 107 -2571 0 net=3483
rlabel metal2 142 -2571 142 -2571 0 net=2065
rlabel metal2 215 -2571 215 -2571 0 net=989
rlabel metal2 450 -2571 450 -2571 0 net=7987
rlabel metal2 1129 -2571 1129 -2571 0 net=8031
rlabel metal2 1234 -2571 1234 -2571 0 net=9777
rlabel metal2 152 -2573 152 -2573 0 net=10739
rlabel metal2 163 -2575 163 -2575 0 net=2048
rlabel metal2 254 -2575 254 -2575 0 net=6832
rlabel metal2 978 -2575 978 -2575 0 net=9294
rlabel metal2 1346 -2575 1346 -2575 0 net=9893
rlabel metal2 1409 -2575 1409 -2575 0 net=12039
rlabel metal2 226 -2577 226 -2577 0 net=1751
rlabel metal2 275 -2577 275 -2577 0 net=5061
rlabel metal2 803 -2577 803 -2577 0 net=9306
rlabel metal2 1423 -2577 1423 -2577 0 net=10641
rlabel metal2 198 -2579 198 -2579 0 net=2209
rlabel metal2 268 -2579 268 -2579 0 net=2869
rlabel metal2 278 -2579 278 -2579 0 net=4664
rlabel metal2 828 -2579 828 -2579 0 net=6265
rlabel metal2 926 -2579 926 -2579 0 net=6490
rlabel metal2 961 -2579 961 -2579 0 net=7815
rlabel metal2 1066 -2579 1066 -2579 0 net=7843
rlabel metal2 1090 -2579 1090 -2579 0 net=11732
rlabel metal2 268 -2581 268 -2581 0 net=1771
rlabel metal2 380 -2581 380 -2581 0 net=4755
rlabel metal2 562 -2581 562 -2581 0 net=3962
rlabel metal2 597 -2581 597 -2581 0 net=12021
rlabel metal2 247 -2583 247 -2583 0 net=3635
rlabel metal2 600 -2583 600 -2583 0 net=10825
rlabel metal2 247 -2585 247 -2585 0 net=2194
rlabel metal2 317 -2585 317 -2585 0 net=2081
rlabel metal2 390 -2585 390 -2585 0 net=4900
rlabel metal2 450 -2585 450 -2585 0 net=2407
rlabel metal2 996 -2585 996 -2585 0 net=11984
rlabel metal2 89 -2587 89 -2587 0 net=11893
rlabel metal2 191 -2589 191 -2589 0 net=2233
rlabel metal2 345 -2589 345 -2589 0 net=2849
rlabel metal2 394 -2589 394 -2589 0 net=2151
rlabel metal2 457 -2589 457 -2589 0 net=4073
rlabel metal2 492 -2589 492 -2589 0 net=3663
rlabel metal2 625 -2589 625 -2589 0 net=5621
rlabel metal2 880 -2589 880 -2589 0 net=7287
rlabel metal2 1017 -2589 1017 -2589 0 net=7245
rlabel metal2 1318 -2589 1318 -2589 0 net=9689
rlabel metal2 1374 -2589 1374 -2589 0 net=10109
rlabel metal2 58 -2591 58 -2591 0 net=7435
rlabel metal2 282 -2591 282 -2591 0 net=2380
rlabel metal2 464 -2591 464 -2591 0 net=4625
rlabel metal2 565 -2591 565 -2591 0 net=11601
rlabel metal2 58 -2593 58 -2593 0 net=3551
rlabel metal2 345 -2593 345 -2593 0 net=1919
rlabel metal2 401 -2593 401 -2593 0 net=3367
rlabel metal2 464 -2593 464 -2593 0 net=3809
rlabel metal2 905 -2593 905 -2593 0 net=6527
rlabel metal2 1073 -2593 1073 -2593 0 net=9053
rlabel metal2 1251 -2593 1251 -2593 0 net=11360
rlabel metal2 233 -2595 233 -2595 0 net=3841
rlabel metal2 401 -2595 401 -2595 0 net=6429
rlabel metal2 555 -2595 555 -2595 0 net=4563
rlabel metal2 786 -2595 786 -2595 0 net=7661
rlabel metal2 1024 -2595 1024 -2595 0 net=11306
rlabel metal2 257 -2597 257 -2597 0 net=2385
rlabel metal2 481 -2597 481 -2597 0 net=3083
rlabel metal2 502 -2597 502 -2597 0 net=4139
rlabel metal2 611 -2597 611 -2597 0 net=3875
rlabel metal2 688 -2597 688 -2597 0 net=5869
rlabel metal2 821 -2597 821 -2597 0 net=6463
rlabel metal2 905 -2597 905 -2597 0 net=6880
rlabel metal2 1027 -2597 1027 -2597 0 net=8528
rlabel metal2 1493 -2597 1493 -2597 0 net=11235
rlabel metal2 156 -2599 156 -2599 0 net=6176
rlabel metal2 614 -2599 614 -2599 0 net=8593
rlabel metal2 1339 -2599 1339 -2599 0 net=9173
rlabel metal2 156 -2601 156 -2601 0 net=1299
rlabel metal2 261 -2601 261 -2601 0 net=1649
rlabel metal2 289 -2601 289 -2601 0 net=1641
rlabel metal2 485 -2601 485 -2601 0 net=2739
rlabel metal2 786 -2601 786 -2601 0 net=4661
rlabel metal2 814 -2601 814 -2601 0 net=5255
rlabel metal2 877 -2601 877 -2601 0 net=5019
rlabel metal2 912 -2601 912 -2601 0 net=6987
rlabel metal2 1038 -2601 1038 -2601 0 net=7733
rlabel metal2 1129 -2601 1129 -2601 0 net=9359
rlabel metal2 1269 -2601 1269 -2601 0 net=9405
rlabel metal2 1416 -2601 1416 -2601 0 net=10601
rlabel metal2 1500 -2601 1500 -2601 0 net=11449
rlabel metal2 163 -2603 163 -2603 0 net=2015
rlabel metal2 1038 -2603 1038 -2603 0 net=8419
rlabel metal2 1178 -2603 1178 -2603 0 net=8495
rlabel metal2 1451 -2603 1451 -2603 0 net=10945
rlabel metal2 240 -2605 240 -2605 0 net=6087
rlabel metal2 912 -2605 912 -2605 0 net=6941
rlabel metal2 1045 -2605 1045 -2605 0 net=8315
rlabel metal2 219 -2607 219 -2607 0 net=2097
rlabel metal2 261 -2607 261 -2607 0 net=3724
rlabel metal2 632 -2607 632 -2607 0 net=4711
rlabel metal2 632 -2607 632 -2607 0 net=4711
rlabel metal2 733 -2607 733 -2607 0 net=8213
rlabel metal2 1220 -2607 1220 -2607 0 net=7825
rlabel metal2 1269 -2607 1269 -2607 0 net=7339
rlabel metal2 219 -2609 219 -2609 0 net=4555
rlabel metal2 289 -2609 289 -2609 0 net=2691
rlabel metal2 520 -2609 520 -2609 0 net=3009
rlabel metal2 733 -2609 733 -2609 0 net=8642
rlabel metal2 1255 -2609 1255 -2609 0 net=9191
rlabel metal2 1367 -2609 1367 -2609 0 net=10091
rlabel metal2 338 -2611 338 -2611 0 net=3397
rlabel metal2 520 -2611 520 -2611 0 net=3949
rlabel metal2 555 -2611 555 -2611 0 net=3485
rlabel metal2 572 -2611 572 -2611 0 net=4024
rlabel metal2 793 -2611 793 -2611 0 net=5335
rlabel metal2 1052 -2611 1052 -2611 0 net=6846
rlabel metal2 1171 -2611 1171 -2611 0 net=8375
rlabel metal2 1227 -2611 1227 -2611 0 net=8449
rlabel metal2 1276 -2611 1276 -2611 0 net=9719
rlabel metal2 499 -2613 499 -2613 0 net=3279
rlabel metal2 569 -2613 569 -2613 0 net=5081
rlabel metal2 800 -2613 800 -2613 0 net=7267
rlabel metal2 1087 -2613 1087 -2613 0 net=8597
rlabel metal2 1241 -2613 1241 -2613 0 net=10165
rlabel metal2 1395 -2613 1395 -2613 0 net=10541
rlabel metal2 471 -2615 471 -2615 0 net=5011
rlabel metal2 863 -2615 863 -2615 0 net=8701
rlabel metal2 1332 -2615 1332 -2615 0 net=9705
rlabel metal2 359 -2617 359 -2617 0 net=2783
rlabel metal2 583 -2617 583 -2617 0 net=6344
rlabel metal2 863 -2617 863 -2617 0 net=6237
rlabel metal2 884 -2617 884 -2617 0 net=6247
rlabel metal2 940 -2617 940 -2617 0 net=7001
rlabel metal2 1031 -2617 1031 -2617 0 net=7281
rlabel metal2 1108 -2617 1108 -2617 0 net=7997
rlabel metal2 1213 -2617 1213 -2617 0 net=8937
rlabel metal2 1290 -2617 1290 -2617 0 net=9563
rlabel metal2 1353 -2617 1353 -2617 0 net=10007
rlabel metal2 208 -2619 208 -2619 0 net=7973
rlabel metal2 1115 -2619 1115 -2619 0 net=7771
rlabel metal2 1311 -2619 1311 -2619 0 net=9603
rlabel metal2 359 -2621 359 -2621 0 net=3877
rlabel metal2 583 -2621 583 -2621 0 net=5811
rlabel metal2 660 -2621 660 -2621 0 net=7949
rlabel metal2 1031 -2621 1031 -2621 0 net=7737
rlabel metal2 331 -2623 331 -2623 0 net=1864
rlabel metal2 670 -2623 670 -2623 0 net=9863
rlabel metal2 79 -2625 79 -2625 0 net=2633
rlabel metal2 604 -2625 604 -2625 0 net=5881
rlabel metal2 740 -2625 740 -2625 0 net=8275
rlabel metal2 79 -2627 79 -2627 0 net=2039
rlabel metal2 702 -2627 702 -2627 0 net=7043
rlabel metal2 1080 -2627 1080 -2627 0 net=8327
rlabel metal2 803 -2629 803 -2629 0 net=9151
rlabel metal2 810 -2631 810 -2631 0 net=1494
rlabel metal2 989 -2631 989 -2631 0 net=7147
rlabel metal2 1164 -2631 1164 -2631 0 net=8269
rlabel metal2 856 -2633 856 -2633 0 net=6893
rlabel metal2 884 -2633 884 -2633 0 net=6646
rlabel metal2 1157 -2633 1157 -2633 0 net=8177
rlabel metal2 1192 -2633 1192 -2633 0 net=8923
rlabel metal2 170 -2635 170 -2635 0 net=7871
rlabel metal2 1150 -2635 1150 -2635 0 net=8157
rlabel metal2 170 -2637 170 -2637 0 net=1591
rlabel metal2 751 -2637 751 -2637 0 net=8249
rlabel metal2 184 -2639 184 -2639 0 net=4389
rlabel metal2 859 -2639 859 -2639 0 net=7413
rlabel metal2 1150 -2639 1150 -2639 0 net=12055
rlabel metal2 506 -2641 506 -2641 0 net=5047
rlabel metal2 919 -2641 919 -2641 0 net=6631
rlabel metal2 982 -2641 982 -2641 0 net=7311
rlabel metal2 506 -2643 506 -2643 0 net=2801
rlabel metal2 919 -2643 919 -2643 0 net=6967
rlabel metal2 436 -2645 436 -2645 0 net=2307
rlabel metal2 968 -2645 968 -2645 0 net=7011
rlabel metal2 436 -2647 436 -2647 0 net=3167
rlabel metal2 968 -2647 968 -2647 0 net=7712
rlabel metal2 513 -2649 513 -2649 0 net=2945
rlabel metal2 1185 -2649 1185 -2649 0 net=12003
rlabel metal2 576 -2651 576 -2651 0 net=5087
rlabel metal2 765 -2653 765 -2653 0 net=5111
rlabel metal2 695 -2655 695 -2655 0 net=4865
rlabel metal2 695 -2657 695 -2657 0 net=4781
rlabel metal2 51 -2659 51 -2659 0 net=8063
rlabel metal2 51 -2661 51 -2661 0 net=3329
rlabel metal2 114 -2663 114 -2663 0 net=7118
rlabel metal2 114 -2665 114 -2665 0 net=2981
rlabel metal2 366 -2667 366 -2667 0 net=5903
rlabel metal2 44 -2678 44 -2678 0 net=3350
rlabel metal2 782 -2678 782 -2678 0 net=11750
rlabel metal2 44 -2680 44 -2680 0 net=4339
rlabel metal2 397 -2680 397 -2680 0 net=2302
rlabel metal2 436 -2680 436 -2680 0 net=3168
rlabel metal2 534 -2680 534 -2680 0 net=4757
rlabel metal2 649 -2680 649 -2680 0 net=4866
rlabel metal2 786 -2680 786 -2680 0 net=4662
rlabel metal2 908 -2680 908 -2680 0 net=7246
rlabel metal2 1524 -2680 1524 -2680 0 net=11876
rlabel metal2 51 -2682 51 -2682 0 net=3330
rlabel metal2 205 -2682 205 -2682 0 net=1920
rlabel metal2 394 -2682 394 -2682 0 net=2341
rlabel metal2 1262 -2682 1262 -2682 0 net=7826
rlabel metal2 58 -2684 58 -2684 0 net=3552
rlabel metal2 264 -2684 264 -2684 0 net=8594
rlabel metal2 58 -2686 58 -2686 0 net=6183
rlabel metal2 135 -2686 135 -2686 0 net=1532
rlabel metal2 198 -2686 198 -2686 0 net=2234
rlabel metal2 331 -2686 331 -2686 0 net=2635
rlabel metal2 446 -2686 446 -2686 0 net=10740
rlabel metal2 72 -2688 72 -2688 0 net=4334
rlabel metal2 681 -2688 681 -2688 0 net=5405
rlabel metal2 786 -2688 786 -2688 0 net=8840
rlabel metal2 1507 -2688 1507 -2688 0 net=12057
rlabel metal2 72 -2690 72 -2690 0 net=1593
rlabel metal2 177 -2690 177 -2690 0 net=2387
rlabel metal2 499 -2690 499 -2690 0 net=5337
rlabel metal2 800 -2690 800 -2690 0 net=7998
rlabel metal2 1185 -2690 1185 -2690 0 net=11072
rlabel metal2 79 -2692 79 -2692 0 net=2040
rlabel metal2 408 -2692 408 -2692 0 net=3368
rlabel metal2 534 -2692 534 -2692 0 net=5413
rlabel metal2 817 -2692 817 -2692 0 net=10570
rlabel metal2 79 -2694 79 -2694 0 net=5113
rlabel metal2 793 -2694 793 -2694 0 net=5257
rlabel metal2 877 -2694 877 -2694 0 net=7002
rlabel metal2 1024 -2694 1024 -2694 0 net=11637
rlabel metal2 1486 -2694 1486 -2694 0 net=12023
rlabel metal2 86 -2696 86 -2696 0 net=4582
rlabel metal2 576 -2696 576 -2696 0 net=5089
rlabel metal2 730 -2696 730 -2696 0 net=8281
rlabel metal2 1185 -2696 1185 -2696 0 net=9174
rlabel metal2 86 -2698 86 -2698 0 net=1827
rlabel metal2 114 -2698 114 -2698 0 net=2983
rlabel metal2 345 -2698 345 -2698 0 net=2083
rlabel metal2 373 -2698 373 -2698 0 net=2153
rlabel metal2 422 -2698 422 -2698 0 net=3281
rlabel metal2 576 -2698 576 -2698 0 net=4783
rlabel metal2 709 -2698 709 -2698 0 net=4564
rlabel metal2 737 -2698 737 -2698 0 net=4654
rlabel metal2 940 -2698 940 -2698 0 net=6632
rlabel metal2 957 -2698 957 -2698 0 net=8924
rlabel metal2 65 -2700 65 -2700 0 net=4939
rlabel metal2 124 -2700 124 -2700 0 net=4649
rlabel metal2 205 -2700 205 -2700 0 net=2099
rlabel metal2 264 -2700 264 -2700 0 net=4194
rlabel metal2 310 -2700 310 -2700 0 net=3707
rlabel metal2 653 -2700 653 -2700 0 net=8871
rlabel metal2 845 -2700 845 -2700 0 net=6427
rlabel metal2 933 -2700 933 -2700 0 net=6249
rlabel metal2 968 -2700 968 -2700 0 net=7289
rlabel metal2 1010 -2700 1010 -2700 0 net=7713
rlabel metal2 65 -2702 65 -2702 0 net=2791
rlabel metal2 156 -2702 156 -2702 0 net=3664
rlabel metal2 653 -2702 653 -2702 0 net=8109
rlabel metal2 1150 -2702 1150 -2702 0 net=11954
rlabel metal2 93 -2704 93 -2704 0 net=4134
rlabel metal2 170 -2704 170 -2704 0 net=2409
rlabel metal2 464 -2704 464 -2704 0 net=3811
rlabel metal2 569 -2704 569 -2704 0 net=5083
rlabel metal2 656 -2704 656 -2704 0 net=7282
rlabel metal2 1073 -2704 1073 -2704 0 net=9055
rlabel metal2 1241 -2704 1241 -2704 0 net=10167
rlabel metal2 93 -2706 93 -2706 0 net=3615
rlabel metal2 275 -2706 275 -2706 0 net=2871
rlabel metal2 275 -2706 275 -2706 0 net=2871
rlabel metal2 296 -2706 296 -2706 0 net=2785
rlabel metal2 520 -2706 520 -2706 0 net=3950
rlabel metal2 880 -2706 880 -2706 0 net=8496
rlabel metal2 100 -2708 100 -2708 0 net=2819
rlabel metal2 212 -2708 212 -2708 0 net=1927
rlabel metal2 352 -2708 352 -2708 0 net=6431
rlabel metal2 415 -2708 415 -2708 0 net=3487
rlabel metal2 569 -2708 569 -2708 0 net=3637
rlabel metal2 604 -2708 604 -2708 0 net=5883
rlabel metal2 744 -2708 744 -2708 0 net=1606
rlabel metal2 765 -2708 765 -2708 0 net=6465
rlabel metal2 880 -2708 880 -2708 0 net=7734
rlabel metal2 1150 -2708 1150 -2708 0 net=9865
rlabel metal2 128 -2710 128 -2710 0 net=4493
rlabel metal2 450 -2710 450 -2710 0 net=2803
rlabel metal2 555 -2710 555 -2710 0 net=5013
rlabel metal2 744 -2710 744 -2710 0 net=8316
rlabel metal2 135 -2712 135 -2712 0 net=3876
rlabel metal2 660 -2712 660 -2712 0 net=7950
rlabel metal2 1101 -2712 1101 -2712 0 net=8277
rlabel metal2 1241 -2712 1241 -2712 0 net=9605
rlabel metal2 1381 -2712 1381 -2712 0 net=11617
rlabel metal2 142 -2714 142 -2714 0 net=2066
rlabel metal2 401 -2714 401 -2714 0 net=3085
rlabel metal2 506 -2714 506 -2714 0 net=4889
rlabel metal2 674 -2714 674 -2714 0 net=3010
rlabel metal2 821 -2714 821 -2714 0 net=6199
rlabel metal2 884 -2714 884 -2714 0 net=6597
rlabel metal2 954 -2714 954 -2714 0 net=9851
rlabel metal2 1188 -2714 1188 -2714 0 net=10697
rlabel metal2 1430 -2714 1430 -2714 0 net=11001
rlabel metal2 142 -2716 142 -2716 0 net=2693
rlabel metal2 425 -2716 425 -2716 0 net=4943
rlabel metal2 611 -2716 611 -2716 0 net=6969
rlabel metal2 926 -2716 926 -2716 0 net=6989
rlabel metal2 1087 -2716 1087 -2716 0 net=8215
rlabel metal2 1262 -2716 1262 -2716 0 net=9707
rlabel metal2 1514 -2716 1514 -2716 0 net=12093
rlabel metal2 149 -2718 149 -2718 0 net=991
rlabel metal2 870 -2718 870 -2718 0 net=6895
rlabel metal2 933 -2718 933 -2718 0 net=7013
rlabel metal2 996 -2718 996 -2718 0 net=7313
rlabel metal2 1024 -2718 1024 -2718 0 net=7975
rlabel metal2 1129 -2718 1129 -2718 0 net=9361
rlabel metal2 1283 -2718 1283 -2718 0 net=10543
rlabel metal2 149 -2720 149 -2720 0 net=1773
rlabel metal2 464 -2720 464 -2720 0 net=4141
rlabel metal2 625 -2720 625 -2720 0 net=5623
rlabel metal2 779 -2720 779 -2720 0 net=8065
rlabel metal2 1108 -2720 1108 -2720 0 net=8251
rlabel metal2 1311 -2720 1311 -2720 0 net=10009
rlabel metal2 1451 -2720 1451 -2720 0 net=11451
rlabel metal2 156 -2722 156 -2722 0 net=7340
rlabel metal2 1353 -2722 1353 -2722 0 net=10329
rlabel metal2 163 -2724 163 -2724 0 net=2017
rlabel metal2 387 -2724 387 -2724 0 net=4641
rlabel metal2 660 -2724 660 -2724 0 net=9778
rlabel metal2 163 -2726 163 -2726 0 net=4557
rlabel metal2 226 -2726 226 -2726 0 net=2211
rlabel metal2 387 -2726 387 -2726 0 net=2309
rlabel metal2 562 -2726 562 -2726 0 net=4627
rlabel metal2 663 -2726 663 -2726 0 net=6383
rlabel metal2 901 -2726 901 -2726 0 net=9875
rlabel metal2 1367 -2726 1367 -2726 0 net=10643
rlabel metal2 138 -2728 138 -2728 0 net=11559
rlabel metal2 215 -2730 215 -2730 0 net=1752
rlabel metal2 408 -2730 408 -2730 0 net=2883
rlabel metal2 681 -2730 681 -2730 0 net=5049
rlabel metal2 849 -2730 849 -2730 0 net=7149
rlabel metal2 1115 -2730 1115 -2730 0 net=7773
rlabel metal2 1192 -2730 1192 -2730 0 net=10111
rlabel metal2 1444 -2730 1444 -2730 0 net=11271
rlabel metal2 219 -2732 219 -2732 0 net=2703
rlabel metal2 366 -2732 366 -2732 0 net=5905
rlabel metal2 856 -2732 856 -2732 0 net=6239
rlabel metal2 905 -2732 905 -2732 0 net=9131
rlabel metal2 1395 -2732 1395 -2732 0 net=10827
rlabel metal2 226 -2734 226 -2734 0 net=1765
rlabel metal2 254 -2734 254 -2734 0 net=1651
rlabel metal2 303 -2734 303 -2734 0 net=3399
rlabel metal2 471 -2734 471 -2734 0 net=2741
rlabel metal2 492 -2734 492 -2734 0 net=5329
rlabel metal2 691 -2734 691 -2734 0 net=7414
rlabel metal2 1115 -2734 1115 -2734 0 net=8451
rlabel metal2 1472 -2734 1472 -2734 0 net=11849
rlabel metal2 212 -2736 212 -2736 0 net=3401
rlabel metal2 527 -2736 527 -2736 0 net=2089
rlabel metal2 695 -2736 695 -2736 0 net=7873
rlabel metal2 1227 -2736 1227 -2736 0 net=9525
rlabel metal2 324 -2738 324 -2738 0 net=3843
rlabel metal2 478 -2738 478 -2738 0 net=2527
rlabel metal2 527 -2738 527 -2738 0 net=4713
rlabel metal2 702 -2738 702 -2738 0 net=7045
rlabel metal2 954 -2738 954 -2738 0 net=8033
rlabel metal2 1255 -2738 1255 -2738 0 net=8939
rlabel metal2 292 -2740 292 -2740 0 net=1095
rlabel metal2 548 -2740 548 -2740 0 net=6089
rlabel metal2 859 -2740 859 -2740 0 net=10991
rlabel metal2 324 -2742 324 -2742 0 net=2947
rlabel metal2 583 -2742 583 -2742 0 net=5813
rlabel metal2 702 -2742 702 -2742 0 net=5063
rlabel metal2 842 -2742 842 -2742 0 net=6528
rlabel metal2 1080 -2742 1080 -2742 0 net=8159
rlabel metal2 1255 -2742 1255 -2742 0 net=9691
rlabel metal2 338 -2744 338 -2744 0 net=3879
rlabel metal2 457 -2744 457 -2744 0 net=4075
rlabel metal2 583 -2744 583 -2744 0 net=5871
rlabel metal2 709 -2744 709 -2744 0 net=5433
rlabel metal2 863 -2744 863 -2744 0 net=6305
rlabel metal2 1160 -2744 1160 -2744 0 net=10383
rlabel metal2 184 -2746 184 -2746 0 net=4391
rlabel metal2 380 -2746 380 -2746 0 net=2851
rlabel metal2 758 -2746 758 -2746 0 net=9192
rlabel metal2 184 -2748 184 -2748 0 net=2499
rlabel metal2 828 -2748 828 -2748 0 net=6267
rlabel metal2 891 -2748 891 -2748 0 net=5020
rlabel metal2 961 -2748 961 -2748 0 net=7817
rlabel metal2 989 -2748 989 -2748 0 net=7663
rlabel metal2 1059 -2748 1059 -2748 0 net=8377
rlabel metal2 1346 -2748 1346 -2748 0 net=10281
rlabel metal2 121 -2750 121 -2750 0 net=6611
rlabel metal2 971 -2750 971 -2750 0 net=8420
rlabel metal2 1094 -2750 1094 -2750 0 net=8179
rlabel metal2 1220 -2750 1220 -2750 0 net=9435
rlabel metal2 121 -2752 121 -2752 0 net=240
rlabel metal2 317 -2752 317 -2752 0 net=1643
rlabel metal2 779 -2752 779 -2752 0 net=7131
rlabel metal2 975 -2752 975 -2752 0 net=7268
rlabel metal2 1136 -2752 1136 -2752 0 net=8599
rlabel metal2 1437 -2752 1437 -2752 0 net=11237
rlabel metal2 107 -2754 107 -2754 0 net=3484
rlabel metal2 191 -2754 191 -2754 0 net=7437
rlabel metal2 828 -2754 828 -2754 0 net=6943
rlabel metal2 947 -2754 947 -2754 0 net=4297
rlabel metal2 107 -2756 107 -2756 0 net=5785
rlabel metal2 289 -2756 289 -2756 0 net=7567
rlabel metal2 978 -2756 978 -2756 0 net=10602
rlabel metal2 667 -2758 667 -2758 0 net=6133
rlabel metal2 1017 -2758 1017 -2758 0 net=7739
rlabel metal2 1038 -2758 1038 -2758 0 net=7989
rlabel metal2 1164 -2758 1164 -2758 0 net=8703
rlabel metal2 1493 -2758 1493 -2758 0 net=12005
rlabel metal2 1031 -2760 1031 -2760 0 net=7845
rlabel metal2 1122 -2760 1122 -2760 0 net=9721
rlabel metal2 1045 -2762 1045 -2762 0 net=8329
rlabel metal2 1234 -2762 1234 -2762 0 net=9565
rlabel metal2 1066 -2764 1066 -2764 0 net=8271
rlabel metal2 1213 -2764 1213 -2764 0 net=9407
rlabel metal2 1332 -2764 1332 -2764 0 net=12041
rlabel metal2 1199 -2766 1199 -2766 0 net=9153
rlabel metal2 1318 -2766 1318 -2766 0 net=10093
rlabel metal2 887 -2768 887 -2768 0 net=10957
rlabel metal2 1248 -2770 1248 -2770 0 net=9647
rlabel metal2 1276 -2772 1276 -2772 0 net=9895
rlabel metal2 1409 -2772 1409 -2772 0 net=10947
rlabel metal2 1290 -2774 1290 -2774 0 net=11603
rlabel metal2 1304 -2776 1304 -2776 0 net=10761
rlabel metal2 1402 -2776 1402 -2776 0 net=10047
rlabel metal2 674 -2778 674 -2778 0 net=9955
rlabel metal2 1402 -2778 1402 -2778 0 net=10903
rlabel metal2 1479 -2780 1479 -2780 0 net=11895
rlabel metal2 58 -2791 58 -2791 0 net=6184
rlabel metal2 247 -2791 247 -2791 0 net=1928
rlabel metal2 296 -2791 296 -2791 0 net=2787
rlabel metal2 296 -2791 296 -2791 0 net=2787
rlabel metal2 303 -2791 303 -2791 0 net=3400
rlabel metal2 593 -2791 593 -2791 0 net=8282
rlabel metal2 747 -2791 747 -2791 0 net=9852
rlabel metal2 1160 -2791 1160 -2791 0 net=10048
rlabel metal2 65 -2793 65 -2793 0 net=2792
rlabel metal2 149 -2793 149 -2793 0 net=1774
rlabel metal2 285 -2793 285 -2793 0 net=3844
rlabel metal2 373 -2793 373 -2793 0 net=2155
rlabel metal2 373 -2793 373 -2793 0 net=2155
rlabel metal2 380 -2793 380 -2793 0 net=1644
rlabel metal2 499 -2793 499 -2793 0 net=5338
rlabel metal2 810 -2793 810 -2793 0 net=11896
rlabel metal2 86 -2795 86 -2795 0 net=1828
rlabel metal2 110 -2795 110 -2795 0 net=6944
rlabel metal2 845 -2795 845 -2795 0 net=7314
rlabel metal2 1006 -2795 1006 -2795 0 net=8940
rlabel metal2 86 -2797 86 -2797 0 net=7439
rlabel metal2 324 -2797 324 -2797 0 net=2948
rlabel metal2 730 -2797 730 -2797 0 net=5885
rlabel metal2 772 -2797 772 -2797 0 net=5406
rlabel metal2 996 -2797 996 -2797 0 net=8601
rlabel metal2 1297 -2797 1297 -2797 0 net=11618
rlabel metal2 93 -2799 93 -2799 0 net=3616
rlabel metal2 866 -2799 866 -2799 0 net=12024
rlabel metal2 93 -2801 93 -2801 0 net=2501
rlabel metal2 198 -2801 198 -2801 0 net=4650
rlabel metal2 310 -2801 310 -2801 0 net=3709
rlabel metal2 331 -2801 331 -2801 0 net=2984
rlabel metal2 499 -2801 499 -2801 0 net=4867
rlabel metal2 688 -2801 688 -2801 0 net=5624
rlabel metal2 737 -2801 737 -2801 0 net=5907
rlabel metal2 772 -2801 772 -2801 0 net=6599
rlabel metal2 898 -2801 898 -2801 0 net=6428
rlabel metal2 1297 -2801 1297 -2801 0 net=10829
rlabel metal2 107 -2803 107 -2803 0 net=6433
rlabel metal2 366 -2803 366 -2803 0 net=3283
rlabel metal2 429 -2803 429 -2803 0 net=2636
rlabel metal2 688 -2803 688 -2803 0 net=9867
rlabel metal2 1185 -2803 1185 -2803 0 net=9693
rlabel metal2 1325 -2803 1325 -2803 0 net=11239
rlabel metal2 100 -2805 100 -2805 0 net=2821
rlabel metal2 443 -2805 443 -2805 0 net=570
rlabel metal2 912 -2805 912 -2805 0 net=6134
rlabel metal2 1255 -2805 1255 -2805 0 net=10011
rlabel metal2 1363 -2805 1363 -2805 0 net=4553
rlabel metal2 114 -2807 114 -2807 0 net=4940
rlabel metal2 121 -2807 121 -2807 0 net=8110
rlabel metal2 723 -2807 723 -2807 0 net=7715
rlabel metal2 1020 -2807 1020 -2807 0 net=12058
rlabel metal2 114 -2809 114 -2809 0 net=2873
rlabel metal2 310 -2809 310 -2809 0 net=2885
rlabel metal2 443 -2809 443 -2809 0 net=5331
rlabel metal2 506 -2809 506 -2809 0 net=4890
rlabel metal2 828 -2809 828 -2809 0 net=7151
rlabel metal2 898 -2809 898 -2809 0 net=8035
rlabel metal2 1010 -2809 1010 -2809 0 net=8705
rlabel metal2 1311 -2809 1311 -2809 0 net=11003
rlabel metal2 338 -2811 338 -2811 0 net=3881
rlabel metal2 506 -2811 506 -2811 0 net=2091
rlabel metal2 653 -2811 653 -2811 0 net=7329
rlabel metal2 1097 -2811 1097 -2811 0 net=10544
rlabel metal2 1381 -2811 1381 -2811 0 net=2485
rlabel metal2 124 -2813 124 -2813 0 net=5451
rlabel metal2 345 -2813 345 -2813 0 net=2084
rlabel metal2 597 -2813 597 -2813 0 net=4642
rlabel metal2 842 -2813 842 -2813 0 net=7057
rlabel metal2 1003 -2813 1003 -2813 0 net=8279
rlabel metal2 1129 -2813 1129 -2813 0 net=7775
rlabel metal2 1150 -2813 1150 -2813 0 net=9877
rlabel metal2 1283 -2813 1283 -2813 0 net=10699
rlabel metal2 1430 -2813 1430 -2813 0 net=12007
rlabel metal2 44 -2815 44 -2815 0 net=4340
rlabel metal2 128 -2815 128 -2815 0 net=4076
rlabel metal2 520 -2815 520 -2815 0 net=2528
rlabel metal2 565 -2815 565 -2815 0 net=10457
rlabel metal2 1374 -2815 1374 -2815 0 net=11639
rlabel metal2 103 -2817 103 -2817 0 net=5383
rlabel metal2 135 -2817 135 -2817 0 net=1298
rlabel metal2 744 -2817 744 -2817 0 net=9937
rlabel metal2 1164 -2817 1164 -2817 0 net=9897
rlabel metal2 135 -2819 135 -2819 0 net=3639
rlabel metal2 590 -2819 590 -2819 0 net=4945
rlabel metal2 625 -2819 625 -2819 0 net=4299
rlabel metal2 1101 -2819 1101 -2819 0 net=9709
rlabel metal2 1276 -2819 1276 -2819 0 net=10645
rlabel metal2 142 -2821 142 -2821 0 net=2695
rlabel metal2 345 -2821 345 -2821 0 net=3087
rlabel metal2 408 -2821 408 -2821 0 net=3403
rlabel metal2 513 -2821 513 -2821 0 net=5435
rlabel metal2 744 -2821 744 -2821 0 net=8180
rlabel metal2 1129 -2821 1129 -2821 0 net=9409
rlabel metal2 1262 -2821 1262 -2821 0 net=10385
rlabel metal2 1367 -2821 1367 -2821 0 net=11561
rlabel metal2 142 -2823 142 -2823 0 net=5611
rlabel metal2 156 -2823 156 -2823 0 net=5015
rlabel metal2 597 -2823 597 -2823 0 net=5051
rlabel metal2 709 -2823 709 -2823 0 net=6909
rlabel metal2 1136 -2823 1136 -2823 0 net=9831
rlabel metal2 159 -2825 159 -2825 0 net=6240
rlabel metal2 1213 -2825 1213 -2825 0 net=10169
rlabel metal2 170 -2827 170 -2827 0 net=2411
rlabel metal2 317 -2827 317 -2827 0 net=4809
rlabel metal2 170 -2829 170 -2829 0 net=2329
rlabel metal2 261 -2829 261 -2829 0 net=3813
rlabel metal2 548 -2829 548 -2829 0 net=6090
rlabel metal2 681 -2829 681 -2829 0 net=7315
rlabel metal2 177 -2831 177 -2831 0 net=2389
rlabel metal2 520 -2831 520 -2831 0 net=6467
rlabel metal2 779 -2831 779 -2831 0 net=6613
rlabel metal2 177 -2833 177 -2833 0 net=2805
rlabel metal2 471 -2833 471 -2833 0 net=2743
rlabel metal2 527 -2833 527 -2833 0 net=4715
rlabel metal2 632 -2833 632 -2833 0 net=5815
rlabel metal2 765 -2833 765 -2833 0 net=6307
rlabel metal2 891 -2833 891 -2833 0 net=7665
rlabel metal2 184 -2835 184 -2835 0 net=2101
rlabel metal2 212 -2835 212 -2835 0 net=11604
rlabel metal2 72 -2837 72 -2837 0 net=1594
rlabel metal2 212 -2837 212 -2837 0 net=2509
rlabel metal2 352 -2837 352 -2837 0 net=2853
rlabel metal2 527 -2837 527 -2837 0 net=6153
rlabel metal2 989 -2837 989 -2837 0 net=8217
rlabel metal2 72 -2839 72 -2839 0 net=4559
rlabel metal2 191 -2839 191 -2839 0 net=5787
rlabel metal2 215 -2839 215 -2839 0 net=384
rlabel metal2 800 -2839 800 -2839 0 net=8873
rlabel metal2 842 -2839 842 -2839 0 net=7818
rlabel metal2 163 -2841 163 -2841 0 net=2019
rlabel metal2 380 -2841 380 -2841 0 net=3777
rlabel metal2 663 -2841 663 -2841 0 net=11311
rlabel metal2 191 -2843 191 -2843 0 net=4845
rlabel metal2 233 -2843 233 -2843 0 net=6021
rlabel metal2 800 -2843 800 -2843 0 net=6251
rlabel metal2 954 -2843 954 -2843 0 net=9667
rlabel metal2 226 -2845 226 -2845 0 net=1767
rlabel metal2 247 -2845 247 -2845 0 net=7874
rlabel metal2 845 -2845 845 -2845 0 net=9021
rlabel metal2 982 -2845 982 -2845 0 net=8273
rlabel metal2 226 -2847 226 -2847 0 net=5084
rlabel metal2 632 -2847 632 -2847 0 net=7977
rlabel metal2 1066 -2847 1066 -2847 0 net=9437
rlabel metal2 254 -2849 254 -2849 0 net=1653
rlabel metal2 387 -2849 387 -2849 0 net=2310
rlabel metal2 849 -2849 849 -2849 0 net=8067
rlabel metal2 219 -2851 219 -2851 0 net=2705
rlabel metal2 401 -2851 401 -2851 0 net=4143
rlabel metal2 534 -2851 534 -2851 0 net=5414
rlabel metal2 856 -2851 856 -2851 0 net=7133
rlabel metal2 1073 -2851 1073 -2851 0 net=9607
rlabel metal2 219 -2853 219 -2853 0 net=4955
rlabel metal2 912 -2853 912 -2853 0 net=10725
rlabel metal2 229 -2855 229 -2855 0 net=9747
rlabel metal2 534 -2855 534 -2855 0 net=5065
rlabel metal2 761 -2855 761 -2855 0 net=10101
rlabel metal2 1241 -2855 1241 -2855 0 net=10331
rlabel metal2 240 -2857 240 -2857 0 net=2213
rlabel metal2 264 -2857 264 -2857 0 net=4392
rlabel metal2 436 -2857 436 -2857 0 net=4495
rlabel metal2 541 -2857 541 -2857 0 net=4759
rlabel metal2 674 -2857 674 -2857 0 net=8079
rlabel metal2 761 -2857 761 -2857 0 net=6990
rlabel metal2 1353 -2857 1353 -2857 0 net=11851
rlabel metal2 79 -2859 79 -2859 0 net=5115
rlabel metal2 450 -2859 450 -2859 0 net=4785
rlabel metal2 618 -2859 618 -2859 0 net=4629
rlabel metal2 695 -2859 695 -2859 0 net=5259
rlabel metal2 814 -2859 814 -2859 0 net=6897
rlabel metal2 961 -2859 961 -2859 0 net=8331
rlabel metal2 1052 -2859 1052 -2859 0 net=9527
rlabel metal2 79 -2861 79 -2861 0 net=10461
rlabel metal2 359 -2861 359 -2861 0 net=3489
rlabel metal2 457 -2861 457 -2861 0 net=2909
rlabel metal2 919 -2861 919 -2861 0 net=9722
rlabel metal2 121 -2863 121 -2863 0 net=5637
rlabel metal2 793 -2863 793 -2863 0 net=6269
rlabel metal2 877 -2863 877 -2863 0 net=10259
rlabel metal2 240 -2865 240 -2865 0 net=6385
rlabel metal2 1045 -2865 1045 -2865 0 net=9155
rlabel metal2 394 -2867 394 -2867 0 net=2343
rlabel metal2 548 -2867 548 -2867 0 net=5091
rlabel metal2 786 -2867 786 -2867 0 net=4787
rlabel metal2 1122 -2867 1122 -2867 0 net=10095
rlabel metal2 145 -2869 145 -2869 0 net=3253
rlabel metal2 555 -2869 555 -2869 0 net=4665
rlabel metal2 611 -2869 611 -2869 0 net=6970
rlabel metal2 716 -2869 716 -2869 0 net=3725
rlabel metal2 786 -2869 786 -2869 0 net=6201
rlabel metal2 870 -2869 870 -2869 0 net=7047
rlabel metal2 1192 -2869 1192 -2869 0 net=10113
rlabel metal2 1318 -2869 1318 -2869 0 net=10763
rlabel metal2 569 -2871 569 -2871 0 net=7951
rlabel metal2 926 -2871 926 -2871 0 net=7015
rlabel metal2 1017 -2871 1017 -2871 0 net=7741
rlabel metal2 1332 -2871 1332 -2871 0 net=12043
rlabel metal2 576 -2873 576 -2873 0 net=7991
rlabel metal2 1332 -2873 1332 -2873 0 net=11273
rlabel metal2 583 -2875 583 -2875 0 net=5873
rlabel metal2 821 -2875 821 -2875 0 net=8252
rlabel metal2 933 -2877 933 -2877 0 net=7569
rlabel metal2 1017 -2877 1017 -2877 0 net=9247
rlabel metal2 1038 -2877 1038 -2877 0 net=9363
rlabel metal2 975 -2879 975 -2879 0 net=8379
rlabel metal2 1108 -2879 1108 -2879 0 net=9567
rlabel metal2 1059 -2881 1059 -2881 0 net=8161
rlabel metal2 1206 -2881 1206 -2881 0 net=10905
rlabel metal2 1080 -2883 1080 -2883 0 net=9057
rlabel metal2 1234 -2883 1234 -2883 0 net=10283
rlabel metal2 1402 -2883 1402 -2883 0 net=12095
rlabel metal2 1171 -2885 1171 -2885 0 net=9649
rlabel metal2 1346 -2885 1346 -2885 0 net=11453
rlabel metal2 1248 -2887 1248 -2887 0 net=10949
rlabel metal2 905 -2889 905 -2889 0 net=4179
rlabel metal2 905 -2891 905 -2891 0 net=7291
rlabel metal2 968 -2893 968 -2893 0 net=8453
rlabel metal2 1115 -2895 1115 -2895 0 net=9133
rlabel metal2 1178 -2897 1178 -2897 0 net=9957
rlabel metal2 1304 -2899 1304 -2899 0 net=10993
rlabel metal2 1416 -2901 1416 -2901 0 net=10959
rlabel metal2 1031 -2903 1031 -2903 0 net=7847
rlabel metal2 663 -2905 663 -2905 0 net=11407
rlabel metal2 72 -2916 72 -2916 0 net=4560
rlabel metal2 250 -2916 250 -2916 0 net=7952
rlabel metal2 583 -2916 583 -2916 0 net=34
rlabel metal2 957 -2916 957 -2916 0 net=9694
rlabel metal2 1199 -2916 1199 -2916 0 net=10115
rlabel metal2 1199 -2916 1199 -2916 0 net=10115
rlabel metal2 1227 -2916 1227 -2916 0 net=10261
rlabel metal2 1360 -2916 1360 -2916 0 net=12008
rlabel metal2 93 -2918 93 -2918 0 net=2502
rlabel metal2 128 -2918 128 -2918 0 net=5385
rlabel metal2 128 -2918 128 -2918 0 net=5385
rlabel metal2 166 -2918 166 -2918 0 net=7992
rlabel metal2 586 -2918 586 -2918 0 net=4630
rlabel metal2 754 -2918 754 -2918 0 net=6270
rlabel metal2 800 -2918 800 -2918 0 net=6252
rlabel metal2 1097 -2918 1097 -2918 0 net=10950
rlabel metal2 1360 -2918 1360 -2918 0 net=4181
rlabel metal2 93 -2920 93 -2920 0 net=8663
rlabel metal2 208 -2920 208 -2920 0 net=2886
rlabel metal2 436 -2920 436 -2920 0 net=5116
rlabel metal2 765 -2920 765 -2920 0 net=6309
rlabel metal2 828 -2920 828 -2920 0 net=7153
rlabel metal2 828 -2920 828 -2920 0 net=7153
rlabel metal2 838 -2920 838 -2920 0 net=7742
rlabel metal2 1227 -2920 1227 -2920 0 net=10013
rlabel metal2 1409 -2920 1409 -2920 0 net=10961
rlabel metal2 100 -2922 100 -2922 0 net=5613
rlabel metal2 184 -2922 184 -2922 0 net=2102
rlabel metal2 289 -2922 289 -2922 0 net=2788
rlabel metal2 310 -2922 310 -2922 0 net=3711
rlabel metal2 457 -2922 457 -2922 0 net=2910
rlabel metal2 838 -2922 838 -2922 0 net=7058
rlabel metal2 891 -2922 891 -2922 0 net=7667
rlabel metal2 912 -2922 912 -2922 0 net=9650
rlabel metal2 1178 -2922 1178 -2922 0 net=9959
rlabel metal2 1178 -2922 1178 -2922 0 net=9959
rlabel metal2 1185 -2922 1185 -2922 0 net=10171
rlabel metal2 1248 -2922 1248 -2922 0 net=10831
rlabel metal2 103 -2924 103 -2924 0 net=1274
rlabel metal2 768 -2924 768 -2924 0 net=9134
rlabel metal2 1136 -2924 1136 -2924 0 net=9833
rlabel metal2 1136 -2924 1136 -2924 0 net=9833
rlabel metal2 1192 -2924 1192 -2924 0 net=10285
rlabel metal2 1276 -2924 1276 -2924 0 net=10647
rlabel metal2 121 -2926 121 -2926 0 net=8068
rlabel metal2 884 -2926 884 -2926 0 net=7016
rlabel metal2 947 -2926 947 -2926 0 net=8274
rlabel metal2 996 -2926 996 -2926 0 net=8603
rlabel metal2 996 -2926 996 -2926 0 net=8603
rlabel metal2 1017 -2926 1017 -2926 0 net=8162
rlabel metal2 1076 -2926 1076 -2926 0 net=10102
rlabel metal2 1234 -2926 1234 -2926 0 net=10727
rlabel metal2 121 -2928 121 -2928 0 net=2511
rlabel metal2 219 -2928 219 -2928 0 net=4957
rlabel metal2 604 -2928 604 -2928 0 net=4667
rlabel metal2 667 -2928 667 -2928 0 net=5817
rlabel metal2 744 -2928 744 -2928 0 net=6023
rlabel metal2 789 -2928 789 -2928 0 net=9058
rlabel metal2 1087 -2928 1087 -2928 0 net=9669
rlabel metal2 1213 -2928 1213 -2928 0 net=10333
rlabel metal2 1269 -2928 1269 -2928 0 net=10459
rlabel metal2 142 -2930 142 -2930 0 net=4705
rlabel metal2 457 -2930 457 -2930 0 net=4947
rlabel metal2 604 -2930 604 -2930 0 net=5909
rlabel metal2 821 -2930 821 -2930 0 net=9087
rlabel metal2 1024 -2930 1024 -2930 0 net=9249
rlabel metal2 1080 -2930 1080 -2930 0 net=9411
rlabel metal2 1220 -2930 1220 -2930 0 net=10387
rlabel metal2 1269 -2930 1269 -2930 0 net=11241
rlabel metal2 107 -2932 107 -2932 0 net=6435
rlabel metal2 611 -2932 611 -2932 0 net=5874
rlabel metal2 646 -2932 646 -2932 0 net=5639
rlabel metal2 681 -2932 681 -2932 0 net=7317
rlabel metal2 891 -2932 891 -2932 0 net=7293
rlabel metal2 912 -2932 912 -2932 0 net=8218
rlabel metal2 1094 -2932 1094 -2932 0 net=9939
rlabel metal2 1206 -2932 1206 -2932 0 net=10907
rlabel metal2 107 -2934 107 -2934 0 net=5093
rlabel metal2 597 -2934 597 -2934 0 net=5053
rlabel metal2 691 -2934 691 -2934 0 net=9273
rlabel metal2 1101 -2934 1101 -2934 0 net=9711
rlabel metal2 1230 -2934 1230 -2934 0 net=1
rlabel metal2 1262 -2934 1262 -2934 0 net=11005
rlabel metal2 142 -2936 142 -2936 0 net=5625
rlabel metal2 709 -2936 709 -2936 0 net=6911
rlabel metal2 807 -2936 807 -2936 0 net=8875
rlabel metal2 1052 -2936 1052 -2936 0 net=9529
rlabel metal2 1241 -2936 1241 -2936 0 net=11275
rlabel metal2 184 -2938 184 -2938 0 net=1659
rlabel metal2 772 -2938 772 -2938 0 net=6601
rlabel metal2 821 -2938 821 -2938 0 net=7049
rlabel metal2 898 -2938 898 -2938 0 net=8037
rlabel metal2 954 -2938 954 -2938 0 net=8333
rlabel metal2 968 -2938 968 -2938 0 net=8455
rlabel metal2 968 -2938 968 -2938 0 net=8455
rlabel metal2 989 -2938 989 -2938 0 net=9157
rlabel metal2 1066 -2938 1066 -2938 0 net=9439
rlabel metal2 1129 -2938 1129 -2938 0 net=9899
rlabel metal2 1304 -2938 1304 -2938 0 net=10995
rlabel metal2 208 -2940 208 -2940 0 net=1768
rlabel metal2 240 -2940 240 -2940 0 net=6387
rlabel metal2 835 -2940 835 -2940 0 net=9227
rlabel metal2 1108 -2940 1108 -2940 0 net=9569
rlabel metal2 1311 -2940 1311 -2940 0 net=12045
rlabel metal2 212 -2942 212 -2942 0 net=3285
rlabel metal2 411 -2942 411 -2942 0 net=11327
rlabel metal2 1388 -2942 1388 -2942 0 net=7849
rlabel metal2 222 -2944 222 -2944 0 net=4786
rlabel metal2 492 -2944 492 -2944 0 net=2621
rlabel metal2 492 -2944 492 -2944 0 net=2621
rlabel metal2 495 -2944 495 -2944 0 net=7565
rlabel metal2 950 -2944 950 -2944 0 net=9209
rlabel metal2 1143 -2944 1143 -2944 0 net=7777
rlabel metal2 226 -2946 226 -2946 0 net=1655
rlabel metal2 275 -2946 275 -2946 0 net=8943
rlabel metal2 597 -2946 597 -2946 0 net=4301
rlabel metal2 639 -2946 639 -2946 0 net=1891
rlabel metal2 688 -2946 688 -2946 0 net=9868
rlabel metal2 842 -2946 842 -2946 0 net=4554
rlabel metal2 163 -2948 163 -2948 0 net=2021
rlabel metal2 275 -2948 275 -2948 0 net=3883
rlabel metal2 443 -2948 443 -2948 0 net=5333
rlabel metal2 751 -2948 751 -2948 0 net=9253
rlabel metal2 1143 -2948 1143 -2948 0 net=9879
rlabel metal2 163 -2950 163 -2950 0 net=3778
rlabel metal2 443 -2950 443 -2950 0 net=4497
rlabel metal2 513 -2950 513 -2950 0 net=5437
rlabel metal2 660 -2950 660 -2950 0 net=3665
rlabel metal2 135 -2952 135 -2952 0 net=3641
rlabel metal2 520 -2952 520 -2952 0 net=6468
rlabel metal2 772 -2952 772 -2952 0 net=6203
rlabel metal2 842 -2952 842 -2952 0 net=7135
rlabel metal2 870 -2952 870 -2952 0 net=10096
rlabel metal2 135 -2954 135 -2954 0 net=7331
rlabel metal2 898 -2954 898 -2954 0 net=7571
rlabel metal2 961 -2954 961 -2954 0 net=8381
rlabel metal2 1017 -2954 1017 -2954 0 net=9673
rlabel metal2 149 -2956 149 -2956 0 net=7503
rlabel metal2 915 -2956 915 -2956 0 net=9364
rlabel metal2 191 -2958 191 -2958 0 net=4847
rlabel metal2 464 -2958 464 -2958 0 net=9749
rlabel metal2 1031 -2958 1031 -2958 0 net=11409
rlabel metal2 191 -2960 191 -2960 0 net=5789
rlabel metal2 229 -2960 229 -2960 0 net=7978
rlabel metal2 786 -2960 786 -2960 0 net=8427
rlabel metal2 1038 -2960 1038 -2960 0 net=9609
rlabel metal2 86 -2962 86 -2962 0 net=7441
rlabel metal2 233 -2962 233 -2962 0 net=8665
rlabel metal2 296 -2962 296 -2962 0 net=6581
rlabel metal2 919 -2962 919 -2962 0 net=8280
rlabel metal2 1073 -2962 1073 -2962 0 net=10764
rlabel metal2 79 -2964 79 -2964 0 net=10463
rlabel metal2 219 -2964 219 -2964 0 net=369
rlabel metal2 940 -2964 940 -2964 0 net=9023
rlabel metal2 1283 -2964 1283 -2964 0 net=10701
rlabel metal2 240 -2966 240 -2966 0 net=2157
rlabel metal2 387 -2966 387 -2966 0 net=2707
rlabel metal2 674 -2966 674 -2966 0 net=8081
rlabel metal2 1003 -2966 1003 -2966 0 net=8707
rlabel metal2 1283 -2966 1283 -2966 0 net=11313
rlabel metal2 170 -2968 170 -2968 0 net=2331
rlabel metal2 401 -2968 401 -2968 0 net=4145
rlabel metal2 520 -2968 520 -2968 0 net=7381
rlabel metal2 1339 -2968 1339 -2968 0 net=11455
rlabel metal2 170 -2970 170 -2970 0 net=5797
rlabel metal2 1346 -2970 1346 -2970 0 net=2487
rlabel metal2 247 -2972 247 -2972 0 net=120
rlabel metal2 282 -2974 282 -2974 0 net=396
rlabel metal2 254 -2976 254 -2976 0 net=2215
rlabel metal2 289 -2976 289 -2976 0 net=2601
rlabel metal2 674 -2976 674 -2976 0 net=9445
rlabel metal2 254 -2978 254 -2978 0 net=3057
rlabel metal2 303 -2978 303 -2978 0 net=2413
rlabel metal2 373 -2978 373 -2978 0 net=3255
rlabel metal2 464 -2978 464 -2978 0 net=2745
rlabel metal2 534 -2978 534 -2978 0 net=5067
rlabel metal2 632 -2978 632 -2978 0 net=9465
rlabel metal2 261 -2980 261 -2980 0 net=3815
rlabel metal2 548 -2980 548 -2980 0 net=4789
rlabel metal2 261 -2982 261 -2982 0 net=2469
rlabel metal2 394 -2982 394 -2982 0 net=3405
rlabel metal2 485 -2982 485 -2982 0 net=3727
rlabel metal2 303 -2984 303 -2984 0 net=4811
rlabel metal2 324 -2984 324 -2984 0 net=2093
rlabel metal2 555 -2984 555 -2984 0 net=5339
rlabel metal2 317 -2986 317 -2986 0 net=2697
rlabel metal2 345 -2986 345 -2986 0 net=3089
rlabel metal2 562 -2986 562 -2986 0 net=4717
rlabel metal2 716 -2986 716 -2986 0 net=5995
rlabel metal2 145 -2988 145 -2988 0 net=4605
rlabel metal2 345 -2988 345 -2988 0 net=4869
rlabel metal2 695 -2988 695 -2988 0 net=5260
rlabel metal2 264 -2990 264 -2990 0 net=5763
rlabel metal2 698 -2990 698 -2990 0 net=8719
rlabel metal2 359 -2992 359 -2992 0 net=3491
rlabel metal2 408 -2992 408 -2992 0 net=7509
rlabel metal2 359 -2994 359 -2994 0 net=2391
rlabel metal2 499 -2994 499 -2994 0 net=3683
rlabel metal2 705 -2994 705 -2994 0 net=12127
rlabel metal2 429 -2996 429 -2996 0 net=2822
rlabel metal2 177 -2998 177 -2998 0 net=2807
rlabel metal2 478 -2998 478 -2998 0 net=4761
rlabel metal2 156 -3000 156 -3000 0 net=5017
rlabel metal2 541 -3000 541 -3000 0 net=7717
rlabel metal2 156 -3002 156 -3002 0 net=2855
rlabel metal2 723 -3002 723 -3002 0 net=5887
rlabel metal2 352 -3004 352 -3004 0 net=2345
rlabel metal2 730 -3004 730 -3004 0 net=6899
rlabel metal2 331 -3006 331 -3006 0 net=5453
rlabel metal2 779 -3006 779 -3006 0 net=6615
rlabel metal2 114 -3008 114 -3008 0 net=2875
rlabel metal2 779 -3008 779 -3008 0 net=5483
rlabel metal2 114 -3010 114 -3010 0 net=10131
rlabel metal2 922 -3012 922 -3012 0 net=11852
rlabel metal2 1353 -3014 1353 -3014 0 net=11563
rlabel metal2 1367 -3016 1367 -3016 0 net=11641
rlabel metal2 1374 -3018 1374 -3018 0 net=12097
rlabel metal2 758 -3020 758 -3020 0 net=4911
rlabel metal2 527 -3022 527 -3022 0 net=6155
rlabel metal2 527 -3024 527 -3024 0 net=3439
rlabel metal2 86 -3035 86 -3035 0 net=10464
rlabel metal2 156 -3035 156 -3035 0 net=2856
rlabel metal2 411 -3035 411 -3035 0 net=2708
rlabel metal2 660 -3035 660 -3035 0 net=9088
rlabel metal2 1017 -3035 1017 -3035 0 net=9211
rlabel metal2 1073 -3035 1073 -3035 0 net=4912
rlabel metal2 93 -3037 93 -3037 0 net=8664
rlabel metal2 835 -3037 835 -3037 0 net=9712
rlabel metal2 1283 -3037 1283 -3037 0 net=11315
rlabel metal2 1283 -3037 1283 -3037 0 net=11315
rlabel metal2 100 -3039 100 -3039 0 net=5614
rlabel metal2 198 -3039 198 -3039 0 net=7442
rlabel metal2 275 -3039 275 -3039 0 net=3885
rlabel metal2 289 -3039 289 -3039 0 net=2603
rlabel metal2 516 -3039 516 -3039 0 net=7718
rlabel metal2 555 -3039 555 -3039 0 net=5341
rlabel metal2 660 -3039 660 -3039 0 net=7511
rlabel metal2 919 -3039 919 -3039 0 net=10996
rlabel metal2 100 -3041 100 -3041 0 net=5387
rlabel metal2 135 -3041 135 -3041 0 net=7333
rlabel metal2 275 -3041 275 -3041 0 net=2415
rlabel metal2 422 -3041 422 -3041 0 net=4848
rlabel metal2 926 -3041 926 -3041 0 net=7566
rlabel metal2 107 -3043 107 -3043 0 net=5094
rlabel metal2 310 -3043 310 -3043 0 net=3712
rlabel metal2 450 -3043 450 -3043 0 net=3091
rlabel metal2 450 -3043 450 -3043 0 net=3091
rlabel metal2 471 -3043 471 -3043 0 net=3643
rlabel metal2 569 -3043 569 -3043 0 net=5069
rlabel metal2 569 -3043 569 -3043 0 net=5069
rlabel metal2 576 -3043 576 -3043 0 net=4959
rlabel metal2 681 -3043 681 -3043 0 net=5334
rlabel metal2 698 -3043 698 -3043 0 net=9158
rlabel metal2 1020 -3043 1020 -3043 0 net=10460
rlabel metal2 107 -3045 107 -3045 0 net=10291
rlabel metal2 310 -3045 310 -3045 0 net=1719
rlabel metal2 873 -3045 873 -3045 0 net=3666
rlabel metal2 114 -3047 114 -3047 0 net=10133
rlabel metal2 114 -3047 114 -3047 0 net=10133
rlabel metal2 128 -3047 128 -3047 0 net=8667
rlabel metal2 324 -3047 324 -3047 0 net=2094
rlabel metal2 863 -3047 863 -3047 0 net=10908
rlabel metal2 135 -3049 135 -3049 0 net=3373
rlabel metal2 1241 -3049 1241 -3049 0 net=11277
rlabel metal2 1325 -3049 1325 -3049 0 net=12129
rlabel metal2 142 -3051 142 -3051 0 net=5627
rlabel metal2 142 -3051 142 -3051 0 net=5627
rlabel metal2 149 -3051 149 -3051 0 net=2441
rlabel metal2 926 -3051 926 -3051 0 net=8605
rlabel metal2 1038 -3051 1038 -3051 0 net=9611
rlabel metal2 1136 -3051 1136 -3051 0 net=9835
rlabel metal2 1241 -3051 1241 -3051 0 net=11243
rlabel metal2 170 -3053 170 -3053 0 net=5799
rlabel metal2 229 -3053 229 -3053 0 net=6005
rlabel metal2 327 -3053 327 -3053 0 net=102
rlabel metal2 691 -3053 691 -3053 0 net=10262
rlabel metal2 170 -3055 170 -3055 0 net=8565
rlabel metal2 338 -3055 338 -3055 0 net=4607
rlabel metal2 513 -3055 513 -3055 0 net=4147
rlabel metal2 583 -3055 583 -3055 0 net=8945
rlabel metal2 1038 -3055 1038 -3055 0 net=9255
rlabel metal2 1115 -3055 1115 -3055 0 net=9671
rlabel metal2 1150 -3055 1150 -3055 0 net=10648
rlabel metal2 184 -3057 184 -3057 0 net=1661
rlabel metal2 338 -3057 338 -3057 0 net=3441
rlabel metal2 534 -3057 534 -3057 0 net=3816
rlabel metal2 618 -3057 618 -3057 0 net=4668
rlabel metal2 698 -3057 698 -3057 0 net=9960
rlabel metal2 1234 -3057 1234 -3057 0 net=10729
rlabel metal2 1297 -3057 1297 -3057 0 net=11389
rlabel metal2 184 -3059 184 -3059 0 net=1657
rlabel metal2 233 -3059 233 -3059 0 net=3059
rlabel metal2 345 -3059 345 -3059 0 net=4870
rlabel metal2 527 -3059 527 -3059 0 net=6437
rlabel metal2 618 -3059 618 -3059 0 net=8941
rlabel metal2 789 -3059 789 -3059 0 net=7979
rlabel metal2 877 -3059 877 -3059 0 net=10389
rlabel metal2 121 -3061 121 -3061 0 net=2512
rlabel metal2 345 -3061 345 -3061 0 net=4707
rlabel metal2 443 -3061 443 -3061 0 net=4499
rlabel metal2 590 -3061 590 -3061 0 net=9274
rlabel metal2 1150 -3061 1150 -3061 0 net=7779
rlabel metal2 1220 -3061 1220 -3061 0 net=10015
rlabel metal2 121 -3063 121 -3063 0 net=9807
rlabel metal2 331 -3063 331 -3063 0 net=2877
rlabel metal2 464 -3063 464 -3063 0 net=2746
rlabel metal2 534 -3063 534 -3063 0 net=4303
rlabel metal2 625 -3063 625 -3063 0 net=5439
rlabel metal2 625 -3063 625 -3063 0 net=5439
rlabel metal2 635 -3063 635 -3063 0 net=5501
rlabel metal2 730 -3063 730 -3063 0 net=6900
rlabel metal2 740 -3063 740 -3063 0 net=8038
rlabel metal2 982 -3063 982 -3063 0 net=8925
rlabel metal2 1213 -3063 1213 -3063 0 net=10335
rlabel metal2 166 -3065 166 -3065 0 net=1953
rlabel metal2 352 -3065 352 -3065 0 net=2347
rlabel metal2 380 -3065 380 -3065 0 net=2471
rlabel metal2 478 -3065 478 -3065 0 net=4763
rlabel metal2 597 -3065 597 -3065 0 net=5641
rlabel metal2 730 -3065 730 -3065 0 net=6311
rlabel metal2 796 -3065 796 -3065 0 net=10405
rlabel metal2 177 -3067 177 -3067 0 net=5018
rlabel metal2 257 -3067 257 -3067 0 net=3197
rlabel metal2 520 -3067 520 -3067 0 net=7383
rlabel metal2 744 -3067 744 -3067 0 net=6025
rlabel metal2 835 -3067 835 -3067 0 net=7137
rlabel metal2 863 -3067 863 -3067 0 net=7295
rlabel metal2 898 -3067 898 -3067 0 net=7573
rlabel metal2 1045 -3067 1045 -3067 0 net=9441
rlabel metal2 1178 -3067 1178 -3067 0 net=11643
rlabel metal2 177 -3069 177 -3069 0 net=3685
rlabel metal2 520 -3069 520 -3069 0 net=1893
rlabel metal2 649 -3069 649 -3069 0 net=9629
rlabel metal2 1101 -3069 1101 -3069 0 net=9675
rlabel metal2 1213 -3069 1213 -3069 0 net=11411
rlabel metal2 1367 -3069 1367 -3069 0 net=7851
rlabel metal2 380 -3071 380 -3071 0 net=4949
rlabel metal2 499 -3071 499 -3071 0 net=5911
rlabel metal2 611 -3071 611 -3071 0 net=5055
rlabel metal2 744 -3071 744 -3071 0 net=9530
rlabel metal2 1304 -3071 1304 -3071 0 net=11565
rlabel metal2 394 -3073 394 -3073 0 net=3407
rlabel metal2 429 -3073 429 -3073 0 net=2809
rlabel metal2 548 -3073 548 -3073 0 net=4791
rlabel metal2 733 -3073 733 -3073 0 net=1
rlabel metal2 842 -3073 842 -3073 0 net=7669
rlabel metal2 933 -3073 933 -3073 0 net=9751
rlabel metal2 1353 -3073 1353 -3073 0 net=4183
rlabel metal2 303 -3075 303 -3075 0 net=4813
rlabel metal2 747 -3075 747 -3075 0 net=11043
rlabel metal2 1360 -3075 1360 -3075 0 net=12099
rlabel metal2 303 -3077 303 -3077 0 net=2333
rlabel metal2 394 -3077 394 -3077 0 net=9295
rlabel metal2 887 -3077 887 -3077 0 net=10125
rlabel metal2 1059 -3077 1059 -3077 0 net=9251
rlabel metal2 1122 -3077 1122 -3077 0 net=9901
rlabel metal2 1374 -3077 1374 -3077 0 net=10963
rlabel metal2 401 -3079 401 -3079 0 net=3493
rlabel metal2 751 -3079 751 -3079 0 net=5485
rlabel metal2 891 -3079 891 -3079 0 net=8335
rlabel metal2 1059 -3079 1059 -3079 0 net=9413
rlabel metal2 1108 -3079 1108 -3079 0 net=9467
rlabel metal2 296 -3081 296 -3081 0 net=6583
rlabel metal2 415 -3081 415 -3081 0 net=5455
rlabel metal2 772 -3081 772 -3081 0 net=6205
rlabel metal2 898 -3081 898 -3081 0 net=10116
rlabel metal2 296 -3083 296 -3083 0 net=3257
rlabel metal2 415 -3083 415 -3083 0 net=2637
rlabel metal2 758 -3083 758 -3083 0 net=6157
rlabel metal2 901 -3083 901 -3083 0 net=9725
rlabel metal2 373 -3085 373 -3085 0 net=1865
rlabel metal2 905 -3085 905 -3085 0 net=8877
rlabel metal2 1080 -3085 1080 -3085 0 net=9881
rlabel metal2 688 -3087 688 -3087 0 net=5889
rlabel metal2 933 -3087 933 -3087 0 net=8383
rlabel metal2 1024 -3087 1024 -3087 0 net=9229
rlabel metal2 1108 -3087 1108 -3087 0 net=10287
rlabel metal2 674 -3089 674 -3089 0 net=9447
rlabel metal2 1143 -3089 1143 -3089 0 net=10173
rlabel metal2 1192 -3089 1192 -3089 0 net=11329
rlabel metal2 674 -3091 674 -3091 0 net=5819
rlabel metal2 716 -3091 716 -3091 0 net=5997
rlabel metal2 940 -3091 940 -3091 0 net=8083
rlabel metal2 1003 -3091 1003 -3091 0 net=8709
rlabel metal2 1290 -3091 1290 -3091 0 net=11457
rlabel metal2 485 -3093 485 -3093 0 net=3729
rlabel metal2 940 -3093 940 -3093 0 net=8457
rlabel metal2 1003 -3093 1003 -3093 0 net=9025
rlabel metal2 1339 -3093 1339 -3093 0 net=2489
rlabel metal2 317 -3095 317 -3095 0 net=2699
rlabel metal2 702 -3095 702 -3095 0 net=4719
rlabel metal2 912 -3095 912 -3095 0 net=8895
rlabel metal2 1031 -3095 1031 -3095 0 net=9941
rlabel metal2 163 -3097 163 -3097 0 net=9633
rlabel metal2 163 -3099 163 -3099 0 net=2023
rlabel metal2 317 -3099 317 -3099 0 net=2393
rlabel metal2 562 -3099 562 -3099 0 net=5765
rlabel metal2 912 -3099 912 -3099 0 net=9570
rlabel metal2 212 -3101 212 -3101 0 net=3287
rlabel metal2 324 -3101 324 -3101 0 net=6285
rlabel metal2 954 -3101 954 -3101 0 net=8429
rlabel metal2 1164 -3101 1164 -3101 0 net=11007
rlabel metal2 191 -3103 191 -3103 0 net=5791
rlabel metal2 240 -3103 240 -3103 0 net=2159
rlabel metal2 975 -3103 975 -3103 0 net=8721
rlabel metal2 1248 -3103 1248 -3103 0 net=10833
rlabel metal2 156 -3105 156 -3105 0 net=3619
rlabel metal2 240 -3105 240 -3105 0 net=3827
rlabel metal2 695 -3107 695 -3107 0 net=10547
rlabel metal2 1010 -3109 1010 -3109 0 net=10702
rlabel metal2 1311 -3111 1311 -3111 0 net=12047
rlabel metal2 884 -3113 884 -3113 0 net=11789
rlabel metal2 856 -3115 856 -3115 0 net=7505
rlabel metal2 849 -3117 849 -3117 0 net=7319
rlabel metal2 828 -3119 828 -3119 0 net=7155
rlabel metal2 814 -3121 814 -3121 0 net=6617
rlabel metal2 814 -3123 814 -3123 0 net=7051
rlabel metal2 737 -3125 737 -3125 0 net=6913
rlabel metal2 492 -3127 492 -3127 0 net=2622
rlabel metal2 492 -3129 492 -3129 0 net=3617
rlabel metal2 786 -3131 786 -3131 0 net=6389
rlabel metal2 800 -3133 800 -3133 0 net=6603
rlabel metal2 807 -3135 807 -3135 0 net=10237
rlabel metal2 100 -3146 100 -3146 0 net=5388
rlabel metal2 184 -3146 184 -3146 0 net=1658
rlabel metal2 331 -3146 331 -3146 0 net=1954
rlabel metal2 394 -3146 394 -3146 0 net=9296
rlabel metal2 758 -3146 758 -3146 0 net=7052
rlabel metal2 842 -3146 842 -3146 0 net=7671
rlabel metal2 842 -3146 842 -3146 0 net=7671
rlabel metal2 863 -3146 863 -3146 0 net=7297
rlabel metal2 863 -3146 863 -3146 0 net=7297
rlabel metal2 898 -3146 898 -3146 0 net=9836
rlabel metal2 1199 -3146 1199 -3146 0 net=10016
rlabel metal2 1293 -3146 1293 -3146 0 net=2490
rlabel metal2 1346 -3146 1346 -3146 0 net=12101
rlabel metal2 107 -3148 107 -3148 0 net=10292
rlabel metal2 296 -3148 296 -3148 0 net=3258
rlabel metal2 698 -3148 698 -3148 0 net=8896
rlabel metal2 1045 -3148 1045 -3148 0 net=9443
rlabel metal2 1045 -3148 1045 -3148 0 net=9443
rlabel metal2 1171 -3148 1171 -3148 0 net=11413
rlabel metal2 1297 -3148 1297 -3148 0 net=11391
rlabel metal2 1297 -3148 1297 -3148 0 net=11391
rlabel metal2 1335 -3148 1335 -3148 0 net=7852
rlabel metal2 114 -3150 114 -3150 0 net=10134
rlabel metal2 191 -3150 191 -3150 0 net=3620
rlabel metal2 254 -3150 254 -3150 0 net=1867
rlabel metal2 387 -3150 387 -3150 0 net=2700
rlabel metal2 492 -3150 492 -3150 0 net=3618
rlabel metal2 870 -3150 870 -3150 0 net=7981
rlabel metal2 912 -3150 912 -3150 0 net=5915
rlabel metal2 1206 -3150 1206 -3150 0 net=11244
rlabel metal2 1353 -3150 1353 -3150 0 net=4185
rlabel metal2 1353 -3150 1353 -3150 0 net=4185
rlabel metal2 1360 -3150 1360 -3150 0 net=10965
rlabel metal2 121 -3152 121 -3152 0 net=9808
rlabel metal2 247 -3152 247 -3152 0 net=2218
rlabel metal2 373 -3152 373 -3152 0 net=3495
rlabel metal2 460 -3152 460 -3152 0 net=6438
rlabel metal2 593 -3152 593 -3152 0 net=486
rlabel metal2 177 -3154 177 -3154 0 net=3687
rlabel metal2 394 -3154 394 -3154 0 net=2811
rlabel metal2 464 -3154 464 -3154 0 net=2472
rlabel metal2 607 -3154 607 -3154 0 net=9752
rlabel metal2 1206 -3154 1206 -3154 0 net=11279
rlabel metal2 177 -3156 177 -3156 0 net=2583
rlabel metal2 807 -3156 807 -3156 0 net=18
rlabel metal2 915 -3156 915 -3156 0 net=819
rlabel metal2 1241 -3156 1241 -3156 0 net=12049
rlabel metal2 191 -3158 191 -3158 0 net=6805
rlabel metal2 758 -3158 758 -3158 0 net=7157
rlabel metal2 870 -3158 870 -3158 0 net=7507
rlabel metal2 943 -3158 943 -3158 0 net=9672
rlabel metal2 1209 -3158 1209 -3158 0 net=12009
rlabel metal2 1276 -3158 1276 -3158 0 net=12131
rlabel metal2 198 -3160 198 -3160 0 net=5801
rlabel metal2 233 -3160 233 -3160 0 net=3061
rlabel metal2 268 -3160 268 -3160 0 net=3289
rlabel metal2 268 -3160 268 -3160 0 net=3289
rlabel metal2 275 -3160 275 -3160 0 net=2417
rlabel metal2 327 -3160 327 -3160 0 net=7595
rlabel metal2 492 -3160 492 -3160 0 net=4793
rlabel metal2 618 -3160 618 -3160 0 net=8942
rlabel metal2 1059 -3160 1059 -3160 0 net=9415
rlabel metal2 1213 -3160 1213 -3160 0 net=11567
rlabel metal2 128 -3162 128 -3162 0 net=8669
rlabel metal2 212 -3162 212 -3162 0 net=5793
rlabel metal2 212 -3162 212 -3162 0 net=5793
rlabel metal2 219 -3162 219 -3162 0 net=1663
rlabel metal2 331 -3162 331 -3162 0 net=4951
rlabel metal2 401 -3162 401 -3162 0 net=6585
rlabel metal2 635 -3162 635 -3162 0 net=6618
rlabel metal2 849 -3162 849 -3162 0 net=8723
rlabel metal2 1234 -3162 1234 -3162 0 net=10407
rlabel metal2 135 -3164 135 -3164 0 net=3375
rlabel metal2 338 -3164 338 -3164 0 net=3442
rlabel metal2 611 -3164 611 -3164 0 net=5503
rlabel metal2 695 -3164 695 -3164 0 net=6159
rlabel metal2 810 -3164 810 -3164 0 net=8710
rlabel metal2 1234 -3164 1234 -3164 0 net=11459
rlabel metal2 184 -3166 184 -3166 0 net=8181
rlabel metal2 338 -3166 338 -3166 0 net=2349
rlabel metal2 401 -3166 401 -3166 0 net=2879
rlabel metal2 464 -3166 464 -3166 0 net=3837
rlabel metal2 233 -3168 233 -3168 0 net=3887
rlabel metal2 345 -3168 345 -3168 0 net=4708
rlabel metal2 772 -3168 772 -3168 0 net=6391
rlabel metal2 877 -3168 877 -3168 0 net=10391
rlabel metal2 1108 -3168 1108 -3168 0 net=10289
rlabel metal2 282 -3170 282 -3170 0 net=2789
rlabel metal2 345 -3170 345 -3170 0 net=3093
rlabel metal2 506 -3170 506 -3170 0 net=2604
rlabel metal2 761 -3170 761 -3170 0 net=6925
rlabel metal2 877 -3170 877 -3170 0 net=8431
rlabel metal2 968 -3170 968 -3170 0 net=8927
rlabel metal2 1108 -3170 1108 -3170 0 net=10337
rlabel metal2 205 -3172 205 -3172 0 net=7335
rlabel metal2 471 -3172 471 -3172 0 net=4609
rlabel metal2 520 -3172 520 -3172 0 net=1894
rlabel metal2 740 -3172 740 -3172 0 net=11257
rlabel metal2 205 -3174 205 -3174 0 net=6007
rlabel metal2 352 -3174 352 -3174 0 net=4305
rlabel metal2 590 -3174 590 -3174 0 net=2793
rlabel metal2 884 -3174 884 -3174 0 net=8337
rlabel metal2 905 -3174 905 -3174 0 net=8879
rlabel metal2 975 -3174 975 -3174 0 net=9231
rlabel metal2 142 -3176 142 -3176 0 net=5629
rlabel metal2 317 -3176 317 -3176 0 net=2394
rlabel metal2 905 -3176 905 -3176 0 net=8385
rlabel metal2 982 -3176 982 -3176 0 net=9213
rlabel metal2 1024 -3176 1024 -3176 0 net=9677
rlabel metal2 240 -3178 240 -3178 0 net=3829
rlabel metal2 359 -3178 359 -3178 0 net=2161
rlabel metal2 415 -3178 415 -3178 0 net=2639
rlabel metal2 471 -3178 471 -3178 0 net=4149
rlabel metal2 625 -3178 625 -3178 0 net=5441
rlabel metal2 919 -3178 919 -3178 0 net=7575
rlabel metal2 1101 -3178 1101 -3178 0 net=10175
rlabel metal2 240 -3180 240 -3180 0 net=5735
rlabel metal2 646 -3180 646 -3180 0 net=6026
rlabel metal2 919 -3180 919 -3180 0 net=8545
rlabel metal2 359 -3182 359 -3182 0 net=3267
rlabel metal2 422 -3182 422 -3182 0 net=3409
rlabel metal2 443 -3182 443 -3182 0 net=5457
rlabel metal2 646 -3182 646 -3182 0 net=5767
rlabel metal2 716 -3182 716 -3182 0 net=3730
rlabel metal2 926 -3182 926 -3182 0 net=8607
rlabel metal2 996 -3182 996 -3182 0 net=10239
rlabel metal2 1143 -3182 1143 -3182 0 net=10835
rlabel metal2 366 -3184 366 -3184 0 net=5057
rlabel metal2 667 -3184 667 -3184 0 net=7385
rlabel metal2 926 -3184 926 -3184 0 net=9027
rlabel metal2 1150 -3184 1150 -3184 0 net=7780
rlabel metal2 408 -3186 408 -3186 0 net=3963
rlabel metal2 422 -3186 422 -3186 0 net=5913
rlabel metal2 513 -3186 513 -3186 0 net=5599
rlabel metal2 667 -3186 667 -3186 0 net=6469
rlabel metal2 961 -3186 961 -3186 0 net=8085
rlabel metal2 163 -3188 163 -3188 0 net=2025
rlabel metal2 443 -3188 443 -3188 0 net=3451
rlabel metal2 513 -3188 513 -3188 0 net=5343
rlabel metal2 681 -3188 681 -3188 0 net=5487
rlabel metal2 765 -3188 765 -3188 0 net=11790
rlabel metal2 156 -3190 156 -3190 0 net=6535
rlabel metal2 303 -3190 303 -3190 0 net=2335
rlabel metal2 520 -3190 520 -3190 0 net=4815
rlabel metal2 555 -3190 555 -3190 0 net=5071
rlabel metal2 597 -3190 597 -3190 0 net=5643
rlabel metal2 709 -3190 709 -3190 0 net=11644
rlabel metal2 303 -3192 303 -3192 0 net=1721
rlabel metal2 527 -3192 527 -3192 0 net=3645
rlabel metal2 548 -3192 548 -3192 0 net=4501
rlabel metal2 597 -3192 597 -3192 0 net=2395
rlabel metal2 996 -3192 996 -3192 0 net=9635
rlabel metal2 1150 -3192 1150 -3192 0 net=11045
rlabel metal2 149 -3194 149 -3194 0 net=2443
rlabel metal2 534 -3194 534 -3194 0 net=6915
rlabel metal2 947 -3194 947 -3194 0 net=10127
rlabel metal2 562 -3196 562 -3196 0 net=6287
rlabel metal2 716 -3196 716 -3196 0 net=6313
rlabel metal2 751 -3196 751 -3196 0 net=11479
rlabel metal2 562 -3198 562 -3198 0 net=4765
rlabel metal2 730 -3198 730 -3198 0 net=6207
rlabel metal2 793 -3198 793 -3198 0 net=6605
rlabel metal2 821 -3198 821 -3198 0 net=7139
rlabel metal2 940 -3198 940 -3198 0 net=8459
rlabel metal2 1003 -3198 1003 -3198 0 net=9613
rlabel metal2 170 -3200 170 -3200 0 net=8567
rlabel metal2 835 -3200 835 -3200 0 net=7321
rlabel metal2 940 -3200 940 -3200 0 net=9252
rlabel metal2 170 -3202 170 -3202 0 net=5999
rlabel metal2 856 -3202 856 -3202 0 net=8947
rlabel metal2 1031 -3202 1031 -3202 0 net=9943
rlabel metal2 478 -3204 478 -3204 0 net=3199
rlabel metal2 989 -3204 989 -3204 0 net=9257
rlabel metal2 1066 -3204 1066 -3204 0 net=10731
rlabel metal2 478 -3206 478 -3206 0 net=9468
rlabel metal2 516 -3208 516 -3208 0 net=6657
rlabel metal2 723 -3208 723 -3208 0 net=9631
rlabel metal2 1129 -3208 1129 -3208 0 net=10549
rlabel metal2 569 -3210 569 -3210 0 net=4961
rlabel metal2 814 -3210 814 -3210 0 net=3209
rlabel metal2 229 -3212 229 -3212 0 net=572
rlabel metal2 1031 -3212 1031 -3212 0 net=9727
rlabel metal2 1248 -3212 1248 -3212 0 net=11317
rlabel metal2 576 -3214 576 -3214 0 net=4720
rlabel metal2 961 -3214 961 -3214 0 net=10411
rlabel metal2 1269 -3214 1269 -3214 0 net=9915
rlabel metal2 688 -3216 688 -3216 0 net=5891
rlabel metal2 1038 -3216 1038 -3216 0 net=9449
rlabel metal2 1087 -3216 1087 -3216 0 net=10017
rlabel metal2 660 -3218 660 -3218 0 net=7513
rlabel metal2 1052 -3218 1052 -3218 0 net=9883
rlabel metal2 660 -3220 660 -3220 0 net=5821
rlabel metal2 1080 -3220 1080 -3220 0 net=9903
rlabel metal2 674 -3222 674 -3222 0 net=3297
rlabel metal2 1122 -3224 1122 -3224 0 net=11009
rlabel metal2 1164 -3226 1164 -3226 0 net=11330
rlabel metal2 796 -3228 796 -3228 0 net=10741
rlabel metal2 156 -3239 156 -3239 0 net=5795
rlabel metal2 219 -3239 219 -3239 0 net=1664
rlabel metal2 499 -3239 499 -3239 0 net=2336
rlabel metal2 712 -3239 712 -3239 0 net=721
rlabel metal2 1290 -3239 1290 -3239 0 net=10409
rlabel metal2 1339 -3239 1339 -3239 0 net=10967
rlabel metal2 163 -3241 163 -3241 0 net=6536
rlabel metal2 212 -3241 212 -3241 0 net=5737
rlabel metal2 243 -3241 243 -3241 0 net=2790
rlabel metal2 352 -3241 352 -3241 0 net=4306
rlabel metal2 702 -3241 702 -3241 0 net=5893
rlabel metal2 702 -3241 702 -3241 0 net=5893
rlabel metal2 733 -3241 733 -3241 0 net=3210
rlabel metal2 838 -3241 838 -3241 0 net=10742
rlabel metal2 1199 -3241 1199 -3241 0 net=11281
rlabel metal2 1227 -3241 1227 -3241 0 net=456
rlabel metal2 1293 -3241 1293 -3241 0 net=11392
rlabel metal2 1346 -3241 1346 -3241 0 net=12103
rlabel metal2 163 -3243 163 -3243 0 net=5059
rlabel metal2 373 -3243 373 -3243 0 net=3497
rlabel metal2 373 -3243 373 -3243 0 net=3497
rlabel metal2 394 -3243 394 -3243 0 net=2812
rlabel metal2 548 -3243 548 -3243 0 net=4503
rlabel metal2 632 -3243 632 -3243 0 net=5489
rlabel metal2 744 -3243 744 -3243 0 net=10732
rlabel metal2 1101 -3243 1101 -3243 0 net=10177
rlabel metal2 1101 -3243 1101 -3243 0 net=10177
rlabel metal2 1136 -3243 1136 -3243 0 net=9417
rlabel metal2 1346 -3243 1346 -3243 0 net=4187
rlabel metal2 170 -3245 170 -3245 0 net=6000
rlabel metal2 499 -3245 499 -3245 0 net=3465
rlabel metal2 751 -3245 751 -3245 0 net=6392
rlabel metal2 807 -3245 807 -3245 0 net=11589
rlabel metal2 1241 -3245 1241 -3245 0 net=12051
rlabel metal2 1241 -3245 1241 -3245 0 net=12051
rlabel metal2 170 -3247 170 -3247 0 net=2619
rlabel metal2 667 -3247 667 -3247 0 net=6471
rlabel metal2 758 -3247 758 -3247 0 net=7159
rlabel metal2 807 -3247 807 -3247 0 net=9115
rlabel metal2 933 -3247 933 -3247 0 net=8609
rlabel metal2 1164 -3247 1164 -3247 0 net=11460
rlabel metal2 177 -3249 177 -3249 0 net=2584
rlabel metal2 408 -3249 408 -3249 0 net=2026
rlabel metal2 527 -3249 527 -3249 0 net=3647
rlabel metal2 527 -3249 527 -3249 0 net=3647
rlabel metal2 541 -3249 541 -3249 0 net=5442
rlabel metal2 758 -3249 758 -3249 0 net=6606
rlabel metal2 810 -3249 810 -3249 0 net=9450
rlabel metal2 1045 -3249 1045 -3249 0 net=9444
rlabel metal2 177 -3251 177 -3251 0 net=8443
rlabel metal2 289 -3251 289 -3251 0 net=8183
rlabel metal2 863 -3251 863 -3251 0 net=7299
rlabel metal2 947 -3251 947 -3251 0 net=8461
rlabel metal2 1143 -3251 1143 -3251 0 net=10837
rlabel metal2 1178 -3251 1178 -3251 0 net=11481
rlabel metal2 1220 -3251 1220 -3251 0 net=12011
rlabel metal2 187 -3253 187 -3253 0 net=1868
rlabel metal2 268 -3253 268 -3253 0 net=3291
rlabel metal2 268 -3253 268 -3253 0 net=3291
rlabel metal2 282 -3253 282 -3253 0 net=2419
rlabel metal2 317 -3253 317 -3253 0 net=3831
rlabel metal2 408 -3253 408 -3253 0 net=3411
rlabel metal2 450 -3253 450 -3253 0 net=7336
rlabel metal2 618 -3253 618 -3253 0 net=6587
rlabel metal2 765 -3253 765 -3253 0 net=6927
rlabel metal2 793 -3253 793 -3253 0 net=7387
rlabel metal2 863 -3253 863 -3253 0 net=8339
rlabel metal2 891 -3253 891 -3253 0 net=9614
rlabel metal2 1024 -3253 1024 -3253 0 net=9679
rlabel metal2 1213 -3253 1213 -3253 0 net=11569
rlabel metal2 198 -3255 198 -3255 0 net=8671
rlabel metal2 247 -3255 247 -3255 0 net=3063
rlabel metal2 296 -3255 296 -3255 0 net=3453
rlabel metal2 450 -3255 450 -3255 0 net=4817
rlabel metal2 541 -3255 541 -3255 0 net=4963
rlabel metal2 618 -3255 618 -3255 0 net=5917
rlabel metal2 947 -3255 947 -3255 0 net=10019
rlabel metal2 1108 -3255 1108 -3255 0 net=10339
rlabel metal2 1213 -3255 1213 -3255 0 net=11319
rlabel metal2 205 -3257 205 -3257 0 net=6009
rlabel metal2 303 -3257 303 -3257 0 net=1723
rlabel metal2 324 -3257 324 -3257 0 net=3095
rlabel metal2 352 -3257 352 -3257 0 net=5345
rlabel metal2 548 -3257 548 -3257 0 net=4767
rlabel metal2 709 -3257 709 -3257 0 net=5415
rlabel metal2 1059 -3257 1059 -3257 0 net=10393
rlabel metal2 205 -3259 205 -3259 0 net=5803
rlabel metal2 247 -3259 247 -3259 0 net=5769
rlabel metal2 737 -3259 737 -3259 0 net=6505
rlabel metal2 198 -3261 198 -3261 0 net=3939
rlabel metal2 303 -3261 303 -3261 0 net=2163
rlabel metal2 387 -3261 387 -3261 0 net=3689
rlabel metal2 562 -3261 562 -3261 0 net=5021
rlabel metal2 768 -3261 768 -3261 0 net=7982
rlabel metal2 912 -3261 912 -3261 0 net=9029
rlabel metal2 954 -3261 954 -3261 0 net=8881
rlabel metal2 191 -3263 191 -3263 0 net=6807
rlabel metal2 387 -3263 387 -3263 0 net=3201
rlabel metal2 786 -3263 786 -3263 0 net=8547
rlabel metal2 954 -3263 954 -3263 0 net=8891
rlabel metal2 191 -3265 191 -3265 0 net=3377
rlabel metal2 331 -3265 331 -3265 0 net=4953
rlabel metal2 415 -3265 415 -3265 0 net=3964
rlabel metal2 779 -3265 779 -3265 0 net=7673
rlabel metal2 870 -3265 870 -3265 0 net=7508
rlabel metal2 964 -3265 964 -3265 0 net=10290
rlabel metal2 275 -3267 275 -3267 0 net=3269
rlabel metal2 415 -3267 415 -3267 0 net=5823
rlabel metal2 800 -3267 800 -3267 0 net=8569
rlabel metal2 996 -3267 996 -3267 0 net=9637
rlabel metal2 1059 -3267 1059 -3267 0 net=9945
rlabel metal2 1171 -3267 1171 -3267 0 net=11415
rlabel metal2 331 -3269 331 -3269 0 net=3839
rlabel metal2 478 -3269 478 -3269 0 net=5645
rlabel metal2 646 -3269 646 -3269 0 net=6161
rlabel metal2 828 -3269 828 -3269 0 net=8725
rlabel metal2 856 -3269 856 -3269 0 net=8949
rlabel metal2 996 -3269 996 -3269 0 net=9729
rlabel metal2 1052 -3269 1052 -3269 0 net=9885
rlabel metal2 1157 -3269 1157 -3269 0 net=11259
rlabel metal2 184 -3271 184 -3271 0 net=11539
rlabel metal2 842 -3271 842 -3271 0 net=8929
rlabel metal2 982 -3271 982 -3271 0 net=9215
rlabel metal2 1052 -3271 1052 -3271 0 net=11047
rlabel metal2 184 -3273 184 -3273 0 net=3889
rlabel metal2 310 -3273 310 -3273 0 net=2445
rlabel metal2 485 -3273 485 -3273 0 net=7597
rlabel metal2 614 -3273 614 -3273 0 net=6905
rlabel metal2 919 -3273 919 -3273 0 net=9233
rlabel metal2 982 -3273 982 -3273 0 net=9259
rlabel metal2 1010 -3273 1010 -3273 0 net=7577
rlabel metal2 233 -3275 233 -3275 0 net=3769
rlabel metal2 968 -3275 968 -3275 0 net=11011
rlabel metal2 1129 -3275 1129 -3275 0 net=10551
rlabel metal2 310 -3277 310 -3277 0 net=2397
rlabel metal2 625 -3277 625 -3277 0 net=5601
rlabel metal2 660 -3277 660 -3277 0 net=10475
rlabel metal2 359 -3279 359 -3279 0 net=2795
rlabel metal2 625 -3279 625 -3279 0 net=4631
rlabel metal2 821 -3279 821 -3279 0 net=7141
rlabel metal2 989 -3279 989 -3279 0 net=8483
rlabel metal2 422 -3281 422 -3281 0 net=5914
rlabel metal2 513 -3281 513 -3281 0 net=6289
rlabel metal2 667 -3281 667 -3281 0 net=7185
rlabel metal2 884 -3281 884 -3281 0 net=8387
rlabel metal2 940 -3281 940 -3281 0 net=8883
rlabel metal2 1017 -3281 1017 -3281 0 net=10241
rlabel metal2 1115 -3281 1115 -3281 0 net=10413
rlabel metal2 422 -3283 422 -3283 0 net=5073
rlabel metal2 583 -3283 583 -3283 0 net=6659
rlabel metal2 653 -3283 653 -3283 0 net=198
rlabel metal2 877 -3283 877 -3283 0 net=8433
rlabel metal2 1017 -3283 1017 -3283 0 net=9905
rlabel metal2 1094 -3283 1094 -3283 0 net=10129
rlabel metal2 429 -3285 429 -3285 0 net=2641
rlabel metal2 583 -3285 583 -3285 0 net=5505
rlabel metal2 681 -3285 681 -3285 0 net=3443
rlabel metal2 877 -3285 877 -3285 0 net=8087
rlabel metal2 429 -3287 429 -3287 0 net=5095
rlabel metal2 1006 -3287 1006 -3287 0 net=10117
rlabel metal2 1262 -3287 1262 -3287 0 net=12133
rlabel metal2 436 -3289 436 -3289 0 net=4795
rlabel metal2 534 -3289 534 -3289 0 net=6917
rlabel metal2 611 -3289 611 -3289 0 net=307
rlabel metal2 1027 -3289 1027 -3289 0 net=10823
rlabel metal2 1269 -3289 1269 -3289 0 net=9917
rlabel metal2 261 -3291 261 -3291 0 net=5631
rlabel metal2 688 -3291 688 -3291 0 net=7515
rlabel metal2 261 -3293 261 -3293 0 net=2881
rlabel metal2 443 -3293 443 -3293 0 net=4611
rlabel metal2 688 -3293 688 -3293 0 net=9779
rlabel metal2 338 -3295 338 -3295 0 net=2351
rlabel metal2 457 -3295 457 -3295 0 net=10139
rlabel metal2 338 -3297 338 -3297 0 net=4151
rlabel metal2 485 -3297 485 -3297 0 net=9632
rlabel metal2 457 -3299 457 -3299 0 net=5459
rlabel metal2 716 -3299 716 -3299 0 net=6315
rlabel metal2 471 -3301 471 -3301 0 net=2337
rlabel metal2 604 -3301 604 -3301 0 net=7323
rlabel metal2 506 -3303 506 -3303 0 net=3299
rlabel metal2 716 -3303 716 -3303 0 net=6209
rlabel metal2 674 -3305 674 -3305 0 net=4315
rlabel metal2 156 -3316 156 -3316 0 net=5796
rlabel metal2 303 -3316 303 -3316 0 net=2164
rlabel metal2 520 -3316 520 -3316 0 net=3690
rlabel metal2 576 -3316 576 -3316 0 net=4504
rlabel metal2 646 -3316 646 -3316 0 net=6163
rlabel metal2 646 -3316 646 -3316 0 net=6163
rlabel metal2 653 -3316 653 -3316 0 net=7516
rlabel metal2 856 -3316 856 -3316 0 net=10340
rlabel metal2 1181 -3316 1181 -3316 0 net=12134
rlabel metal2 1269 -3316 1269 -3316 0 net=10410
rlabel metal2 1339 -3316 1339 -3316 0 net=10969
rlabel metal2 1339 -3316 1339 -3316 0 net=10969
rlabel metal2 1346 -3316 1346 -3316 0 net=4189
rlabel metal2 1346 -3316 1346 -3316 0 net=4189
rlabel metal2 1353 -3316 1353 -3316 0 net=12105
rlabel metal2 1353 -3316 1353 -3316 0 net=12105
rlabel metal2 163 -3318 163 -3318 0 net=5060
rlabel metal2 436 -3318 436 -3318 0 net=4797
rlabel metal2 544 -3318 544 -3318 0 net=6472
rlabel metal2 761 -3318 761 -3318 0 net=8434
rlabel metal2 1003 -3318 1003 -3318 0 net=9886
rlabel metal2 1136 -3318 1136 -3318 0 net=12052
rlabel metal2 1272 -3318 1272 -3318 0 net=9918
rlabel metal2 177 -3320 177 -3320 0 net=8444
rlabel metal2 611 -3320 611 -3320 0 net=5603
rlabel metal2 660 -3320 660 -3320 0 net=7674
rlabel metal2 786 -3320 786 -3320 0 net=8549
rlabel metal2 824 -3320 824 -3320 0 net=8610
rlabel metal2 1073 -3320 1073 -3320 0 net=10553
rlabel metal2 184 -3322 184 -3322 0 net=3890
rlabel metal2 254 -3322 254 -3322 0 net=3065
rlabel metal2 254 -3322 254 -3322 0 net=3065
rlabel metal2 261 -3322 261 -3322 0 net=2882
rlabel metal2 411 -3322 411 -3322 0 net=294
rlabel metal2 891 -3322 891 -3322 0 net=9216
rlabel metal2 1038 -3322 1038 -3322 0 net=8462
rlabel metal2 1055 -3322 1055 -3322 0 net=10242
rlabel metal2 1139 -3322 1139 -3322 0 net=10824
rlabel metal2 198 -3324 198 -3324 0 net=8673
rlabel metal2 226 -3324 226 -3324 0 net=3941
rlabel metal2 282 -3324 282 -3324 0 net=2421
rlabel metal2 359 -3324 359 -3324 0 net=2796
rlabel metal2 670 -3324 670 -3324 0 net=8882
rlabel metal2 205 -3326 205 -3326 0 net=5805
rlabel metal2 205 -3326 205 -3326 0 net=5805
rlabel metal2 212 -3326 212 -3326 0 net=5739
rlabel metal2 212 -3326 212 -3326 0 net=5739
rlabel metal2 226 -3326 226 -3326 0 net=2399
rlabel metal2 387 -3326 387 -3326 0 net=3202
rlabel metal2 870 -3326 870 -3326 0 net=9680
rlabel metal2 275 -3328 275 -3328 0 net=3271
rlabel metal2 387 -3328 387 -3328 0 net=5647
rlabel metal2 513 -3328 513 -3328 0 net=6291
rlabel metal2 660 -3328 660 -3328 0 net=6507
rlabel metal2 751 -3328 751 -3328 0 net=7161
rlabel metal2 779 -3328 779 -3328 0 net=8185
rlabel metal2 828 -3328 828 -3328 0 net=8727
rlabel metal2 828 -3328 828 -3328 0 net=8727
rlabel metal2 835 -3328 835 -3328 0 net=7578
rlabel metal2 275 -3330 275 -3330 0 net=4954
rlabel metal2 394 -3330 394 -3330 0 net=3301
rlabel metal2 513 -3330 513 -3330 0 net=2165
rlabel metal2 667 -3330 667 -3330 0 net=6317
rlabel metal2 737 -3330 737 -3330 0 net=6929
rlabel metal2 807 -3330 807 -3330 0 net=9117
rlabel metal2 835 -3330 835 -3330 0 net=8571
rlabel metal2 947 -3330 947 -3330 0 net=10021
rlabel metal2 1192 -3330 1192 -3330 0 net=11321
rlabel metal2 282 -3332 282 -3332 0 net=3455
rlabel metal2 310 -3332 310 -3332 0 net=1725
rlabel metal2 345 -3332 345 -3332 0 net=3499
rlabel metal2 422 -3332 422 -3332 0 net=5074
rlabel metal2 569 -3332 569 -3332 0 net=7599
rlabel metal2 838 -3332 838 -3332 0 net=10130
rlabel metal2 219 -3334 219 -3334 0 net=3195
rlabel metal2 572 -3334 572 -3334 0 net=6409
rlabel metal2 761 -3334 761 -3334 0 net=9638
rlabel metal2 296 -3336 296 -3336 0 net=3097
rlabel metal2 373 -3336 373 -3336 0 net=2353
rlabel metal2 436 -3336 436 -3336 0 net=2447
rlabel metal2 478 -3336 478 -3336 0 net=4965
rlabel metal2 632 -3336 632 -3336 0 net=5491
rlabel metal2 842 -3336 842 -3336 0 net=8931
rlabel metal2 842 -3336 842 -3336 0 net=8931
rlabel metal2 849 -3336 849 -3336 0 net=8951
rlabel metal2 1003 -3336 1003 -3336 0 net=11049
rlabel metal2 317 -3338 317 -3338 0 net=3413
rlabel metal2 506 -3338 506 -3338 0 net=4335
rlabel metal2 632 -3338 632 -3338 0 net=6015
rlabel metal2 765 -3338 765 -3338 0 net=7389
rlabel metal2 856 -3338 856 -3338 0 net=8885
rlabel metal2 947 -3338 947 -3338 0 net=11013
rlabel metal2 1024 -3338 1024 -3338 0 net=12013
rlabel metal2 324 -3340 324 -3340 0 net=2339
rlabel metal2 534 -3340 534 -3340 0 net=8357
rlabel metal2 870 -3340 870 -3340 0 net=10141
rlabel metal2 170 -3342 170 -3342 0 net=2620
rlabel metal2 534 -3342 534 -3342 0 net=4769
rlabel metal2 681 -3342 681 -3342 0 net=3445
rlabel metal2 1027 -3342 1027 -3342 0 net=11416
rlabel metal2 331 -3344 331 -3344 0 net=3840
rlabel metal2 884 -3344 884 -3344 0 net=8389
rlabel metal2 1045 -3344 1045 -3344 0 net=10395
rlabel metal2 1185 -3344 1185 -3344 0 net=11283
rlabel metal2 331 -3346 331 -3346 0 net=4613
rlabel metal2 548 -3346 548 -3346 0 net=4633
rlabel metal2 688 -3346 688 -3346 0 net=5894
rlabel metal2 730 -3346 730 -3346 0 net=6589
rlabel metal2 884 -3346 884 -3346 0 net=9781
rlabel metal2 1052 -3346 1052 -3346 0 net=9418
rlabel metal2 380 -3348 380 -3348 0 net=6808
rlabel metal2 408 -3348 408 -3348 0 net=4319
rlabel metal2 492 -3348 492 -3348 0 net=5633
rlabel metal2 702 -3348 702 -3348 0 net=6211
rlabel metal2 744 -3348 744 -3348 0 net=8089
rlabel metal2 891 -3348 891 -3348 0 net=9031
rlabel metal2 926 -3348 926 -3348 0 net=11591
rlabel metal2 380 -3350 380 -3350 0 net=3467
rlabel metal2 597 -3350 597 -3350 0 net=6661
rlabel metal2 691 -3350 691 -3350 0 net=7585
rlabel metal2 877 -3350 877 -3350 0 net=9261
rlabel metal2 1094 -3350 1094 -3350 0 net=10415
rlabel metal2 443 -3352 443 -3352 0 net=3649
rlabel metal2 618 -3352 618 -3352 0 net=5919
rlabel metal2 894 -3352 894 -3352 0 net=7300
rlabel metal2 940 -3352 940 -3352 0 net=10119
rlabel metal2 1122 -3352 1122 -3352 0 net=11571
rlabel metal2 450 -3354 450 -3354 0 net=4819
rlabel metal2 527 -3354 527 -3354 0 net=4257
rlabel metal2 898 -3354 898 -3354 0 net=6906
rlabel metal2 1080 -3354 1080 -3354 0 net=10179
rlabel metal2 233 -3356 233 -3356 0 net=3771
rlabel metal2 457 -3356 457 -3356 0 net=5461
rlabel metal2 898 -3356 898 -3356 0 net=8893
rlabel metal2 961 -3356 961 -3356 0 net=11483
rlabel metal2 233 -3358 233 -3358 0 net=4153
rlabel metal2 422 -3358 422 -3358 0 net=3787
rlabel metal2 492 -3358 492 -3358 0 net=7325
rlabel metal2 758 -3358 758 -3358 0 net=322
rlabel metal2 975 -3358 975 -3358 0 net=7142
rlabel metal2 1017 -3358 1017 -3358 0 net=9907
rlabel metal2 338 -3360 338 -3360 0 net=5023
rlabel metal2 576 -3360 576 -3360 0 net=5573
rlabel metal2 674 -3360 674 -3360 0 net=4317
rlabel metal2 982 -3360 982 -3360 0 net=11261
rlabel metal2 247 -3362 247 -3362 0 net=5771
rlabel metal2 905 -3362 905 -3362 0 net=9235
rlabel metal2 933 -3362 933 -3362 0 net=8485
rlabel metal2 1013 -3362 1013 -3362 0 net=2473
rlabel metal2 191 -3364 191 -3364 0 net=3379
rlabel metal2 352 -3364 352 -3364 0 net=5347
rlabel metal2 583 -3364 583 -3364 0 net=5507
rlabel metal2 912 -3364 912 -3364 0 net=9731
rlabel metal2 352 -3366 352 -3366 0 net=2643
rlabel metal2 583 -3366 583 -3366 0 net=5417
rlabel metal2 800 -3366 800 -3366 0 net=7187
rlabel metal2 415 -3368 415 -3368 0 net=5824
rlabel metal2 590 -3368 590 -3368 0 net=6919
rlabel metal2 800 -3368 800 -3368 0 net=8341
rlabel metal2 919 -3368 919 -3368 0 net=11083
rlabel metal2 404 -3370 404 -3370 0 net=5463
rlabel metal2 695 -3370 695 -3370 0 net=11541
rlabel metal2 989 -3370 989 -3370 0 net=9947
rlabel metal2 415 -3372 415 -3372 0 net=5097
rlabel metal2 656 -3372 656 -3372 0 net=11717
rlabel metal2 1059 -3372 1059 -3372 0 net=10477
rlabel metal2 366 -3374 366 -3374 0 net=3833
rlabel metal2 520 -3374 520 -3374 0 net=4505
rlabel metal2 1129 -3374 1129 -3374 0 net=10839
rlabel metal2 289 -3376 289 -3376 0 net=6011
rlabel metal2 268 -3378 268 -3378 0 net=3293
rlabel metal2 198 -3389 198 -3389 0 net=8674
rlabel metal2 296 -3389 296 -3389 0 net=3098
rlabel metal2 457 -3389 457 -3389 0 net=3788
rlabel metal2 492 -3389 492 -3389 0 net=7326
rlabel metal2 681 -3389 681 -3389 0 net=6663
rlabel metal2 681 -3389 681 -3389 0 net=6663
rlabel metal2 723 -3389 723 -3389 0 net=6410
rlabel metal2 793 -3389 793 -3389 0 net=10142
rlabel metal2 1003 -3389 1003 -3389 0 net=11051
rlabel metal2 1003 -3389 1003 -3389 0 net=11051
rlabel metal2 1013 -3389 1013 -3389 0 net=10022
rlabel metal2 1101 -3389 1101 -3389 0 net=9909
rlabel metal2 1178 -3389 1178 -3389 0 net=11285
rlabel metal2 1339 -3389 1339 -3389 0 net=10971
rlabel metal2 1339 -3389 1339 -3389 0 net=10971
rlabel metal2 1346 -3389 1346 -3389 0 net=4191
rlabel metal2 205 -3391 205 -3391 0 net=5806
rlabel metal2 317 -3391 317 -3391 0 net=3414
rlabel metal2 422 -3391 422 -3391 0 net=10819
rlabel metal2 737 -3391 737 -3391 0 net=6931
rlabel metal2 807 -3391 807 -3391 0 net=5493
rlabel metal2 824 -3391 824 -3391 0 net=8894
rlabel metal2 1027 -3391 1027 -3391 0 net=11572
rlabel metal2 1181 -3391 1181 -3391 0 net=11322
rlabel metal2 1346 -3391 1346 -3391 0 net=12107
rlabel metal2 212 -3393 212 -3393 0 net=5740
rlabel metal2 271 -3393 271 -3393 0 net=548
rlabel metal2 737 -3393 737 -3393 0 net=4318
rlabel metal2 1066 -3393 1066 -3393 0 net=10180
rlabel metal2 1087 -3393 1087 -3393 0 net=10417
rlabel metal2 1115 -3393 1115 -3393 0 net=10841
rlabel metal2 219 -3395 219 -3395 0 net=3196
rlabel metal2 530 -3395 530 -3395 0 net=38
rlabel metal2 579 -3395 579 -3395 0 net=6164
rlabel metal2 649 -3395 649 -3395 0 net=11484
rlabel metal2 1010 -3395 1010 -3395 0 net=7467
rlabel metal2 247 -3397 247 -3397 0 net=3380
rlabel metal2 555 -3397 555 -3397 0 net=5465
rlabel metal2 597 -3397 597 -3397 0 net=5462
rlabel metal2 653 -3397 653 -3397 0 net=7189
rlabel metal2 1010 -3397 1010 -3397 0 net=10397
rlabel metal2 240 -3399 240 -3399 0 net=3943
rlabel metal2 261 -3399 261 -3399 0 net=3294
rlabel metal2 324 -3399 324 -3399 0 net=2340
rlabel metal2 366 -3399 366 -3399 0 net=6012
rlabel metal2 408 -3399 408 -3399 0 net=3835
rlabel metal2 450 -3399 450 -3399 0 net=3773
rlabel metal2 558 -3399 558 -3399 0 net=2887
rlabel metal2 667 -3399 667 -3399 0 net=6319
rlabel metal2 807 -3399 807 -3399 0 net=9263
rlabel metal2 933 -3399 933 -3399 0 net=8487
rlabel metal2 1031 -3399 1031 -3399 0 net=8391
rlabel metal2 226 -3401 226 -3401 0 net=2400
rlabel metal2 387 -3401 387 -3401 0 net=5649
rlabel metal2 450 -3401 450 -3401 0 net=5605
rlabel metal2 667 -3401 667 -3401 0 net=8359
rlabel metal2 859 -3401 859 -3401 0 net=1112
rlabel metal2 877 -3401 877 -3401 0 net=9033
rlabel metal2 961 -3401 961 -3401 0 net=12015
rlabel metal2 1031 -3401 1031 -3401 0 net=10479
rlabel metal2 254 -3403 254 -3403 0 net=3067
rlabel metal2 282 -3403 282 -3403 0 net=3457
rlabel metal2 359 -3403 359 -3403 0 net=3273
rlabel metal2 401 -3403 401 -3403 0 net=4967
rlabel metal2 485 -3403 485 -3403 0 net=4799
rlabel metal2 716 -3403 716 -3403 0 net=7587
rlabel metal2 968 -3403 968 -3403 0 net=3446
rlabel metal2 303 -3405 303 -3405 0 net=2423
rlabel metal2 345 -3405 345 -3405 0 net=3501
rlabel metal2 415 -3405 415 -3405 0 net=5099
rlabel metal2 457 -3405 457 -3405 0 net=4259
rlabel metal2 548 -3405 548 -3405 0 net=4635
rlabel metal2 716 -3405 716 -3405 0 net=7601
rlabel metal2 786 -3405 786 -3405 0 net=8343
rlabel metal2 863 -3405 863 -3405 0 net=11542
rlabel metal2 968 -3405 968 -3405 0 net=9949
rlabel metal2 233 -3407 233 -3407 0 net=4154
rlabel metal2 373 -3407 373 -3407 0 net=2355
rlabel metal2 478 -3407 478 -3407 0 net=4337
rlabel metal2 541 -3407 541 -3407 0 net=530
rlabel metal2 569 -3407 569 -3407 0 net=5508
rlabel metal2 660 -3407 660 -3407 0 net=6509
rlabel metal2 800 -3407 800 -3407 0 net=9119
rlabel metal2 863 -3407 863 -3407 0 net=11085
rlabel metal2 1349 -3407 1349 -3407 0 net=1
rlabel metal2 373 -3409 373 -3409 0 net=6455
rlabel metal2 919 -3409 919 -3409 0 net=11015
rlabel metal2 394 -3411 394 -3411 0 net=3303
rlabel metal2 572 -3411 572 -3411 0 net=1456
rlabel metal2 338 -3413 338 -3413 0 net=5025
rlabel metal2 485 -3413 485 -3413 0 net=4821
rlabel metal2 506 -3413 506 -3413 0 net=5575
rlabel metal2 618 -3413 618 -3413 0 net=11719
rlabel metal2 940 -3413 940 -3413 0 net=10121
rlabel metal2 310 -3415 310 -3415 0 net=1727
rlabel metal2 436 -3415 436 -3415 0 net=2449
rlabel metal2 632 -3415 632 -3415 0 net=6017
rlabel metal2 905 -3415 905 -3415 0 net=9237
rlabel metal2 310 -3417 310 -3417 0 net=4615
rlabel metal2 380 -3417 380 -3417 0 net=3469
rlabel metal2 499 -3417 499 -3417 0 net=8186
rlabel metal2 856 -3417 856 -3417 0 net=8887
rlabel metal2 331 -3419 331 -3419 0 net=2167
rlabel metal2 541 -3419 541 -3419 0 net=6293
rlabel metal2 674 -3419 674 -3419 0 net=5773
rlabel metal2 380 -3421 380 -3421 0 net=4321
rlabel metal2 513 -3421 513 -3421 0 net=4507
rlabel metal2 562 -3421 562 -3421 0 net=5349
rlabel metal2 674 -3421 674 -3421 0 net=7163
rlabel metal2 352 -3423 352 -3423 0 net=2645
rlabel metal2 576 -3423 576 -3423 0 net=5635
rlabel metal2 632 -3423 632 -3423 0 net=8573
rlabel metal2 352 -3425 352 -3425 0 net=9515
rlabel metal2 443 -3425 443 -3425 0 net=3651
rlabel metal2 625 -3425 625 -3425 0 net=6921
rlabel metal2 835 -3425 835 -3425 0 net=8933
rlabel metal2 464 -3427 464 -3427 0 net=5719
rlabel metal2 639 -3427 639 -3427 0 net=7391
rlabel metal2 842 -3427 842 -3427 0 net=11593
rlabel metal2 471 -3429 471 -3429 0 net=4771
rlabel metal2 688 -3429 688 -3429 0 net=5921
rlabel metal2 912 -3429 912 -3429 0 net=9733
rlabel metal2 534 -3431 534 -3431 0 net=5419
rlabel metal2 702 -3431 702 -3431 0 net=6213
rlabel metal2 765 -3431 765 -3431 0 net=8729
rlabel metal2 912 -3431 912 -3431 0 net=11263
rlabel metal2 583 -3433 583 -3433 0 net=8090
rlabel metal2 828 -3433 828 -3433 0 net=9783
rlabel metal2 982 -3433 982 -3433 0 net=11897
rlabel metal2 702 -3435 702 -3435 0 net=6591
rlabel metal2 744 -3435 744 -3435 0 net=2475
rlabel metal2 1038 -3435 1038 -3435 0 net=10555
rlabel metal2 709 -3437 709 -3437 0 net=8551
rlabel metal2 884 -3437 884 -3437 0 net=11217
rlabel metal2 730 -3439 730 -3439 0 net=8953
rlabel metal2 740 -3441 740 -3441 0 net=9639
rlabel metal2 247 -3452 247 -3452 0 net=3945
rlabel metal2 247 -3452 247 -3452 0 net=3945
rlabel metal2 261 -3452 261 -3452 0 net=3069
rlabel metal2 261 -3452 261 -3452 0 net=3069
rlabel metal2 275 -3452 275 -3452 0 net=7895
rlabel metal2 292 -3452 292 -3452 0 net=4616
rlabel metal2 331 -3452 331 -3452 0 net=2169
rlabel metal2 380 -3452 380 -3452 0 net=4323
rlabel metal2 464 -3452 464 -3452 0 net=5720
rlabel metal2 513 -3452 513 -3452 0 net=4508
rlabel metal2 611 -3452 611 -3452 0 net=4636
rlabel metal2 677 -3452 677 -3452 0 net=277
rlabel metal2 989 -3452 989 -3452 0 net=10399
rlabel metal2 1045 -3452 1045 -3452 0 net=8393
rlabel metal2 1080 -3452 1080 -3452 0 net=10419
rlabel metal2 1094 -3452 1094 -3452 0 net=7469
rlabel metal2 1136 -3452 1136 -3452 0 net=9911
rlabel metal2 1178 -3452 1178 -3452 0 net=11287
rlabel metal2 1178 -3452 1178 -3452 0 net=11287
rlabel metal2 1339 -3452 1339 -3452 0 net=10973
rlabel metal2 317 -3454 317 -3454 0 net=3459
rlabel metal2 338 -3454 338 -3454 0 net=1729
rlabel metal2 359 -3454 359 -3454 0 net=3503
rlabel metal2 380 -3454 380 -3454 0 net=3471
rlabel metal2 513 -3454 513 -3454 0 net=5421
rlabel metal2 611 -3454 611 -3454 0 net=8361
rlabel metal2 688 -3454 688 -3454 0 net=6592
rlabel metal2 726 -3454 726 -3454 0 net=9264
rlabel metal2 817 -3454 817 -3454 0 net=11086
rlabel metal2 870 -3454 870 -3454 0 net=536
rlabel metal2 898 -3454 898 -3454 0 net=11898
rlabel metal2 996 -3454 996 -3454 0 net=10556
rlabel metal2 1087 -3454 1087 -3454 0 net=5985
rlabel metal2 1339 -3454 1339 -3454 0 net=12109
rlabel metal2 324 -3456 324 -3456 0 net=2425
rlabel metal2 359 -3456 359 -3456 0 net=3275
rlabel metal2 408 -3456 408 -3456 0 net=3836
rlabel metal2 478 -3456 478 -3456 0 net=4338
rlabel metal2 604 -3456 604 -3456 0 net=2451
rlabel metal2 681 -3456 681 -3456 0 net=6665
rlabel metal2 691 -3456 691 -3456 0 net=11594
rlabel metal2 849 -3456 849 -3456 0 net=9640
rlabel metal2 905 -3456 905 -3456 0 net=8888
rlabel metal2 1003 -3456 1003 -3456 0 net=11053
rlabel metal2 1003 -3456 1003 -3456 0 net=11053
rlabel metal2 1010 -3456 1010 -3456 0 net=10481
rlabel metal2 1108 -3456 1108 -3456 0 net=10843
rlabel metal2 1346 -3456 1346 -3456 0 net=4192
rlabel metal2 408 -3458 408 -3458 0 net=5607
rlabel metal2 478 -3458 478 -3458 0 net=4651
rlabel metal2 597 -3458 597 -3458 0 net=4801
rlabel metal2 628 -3458 628 -3458 0 net=1222
rlabel metal2 422 -3460 422 -3460 0 net=5101
rlabel metal2 499 -3460 499 -3460 0 net=3803
rlabel metal2 562 -3460 562 -3460 0 net=2647
rlabel metal2 646 -3460 646 -3460 0 net=4289
rlabel metal2 744 -3460 744 -3460 0 net=2477
rlabel metal2 744 -3460 744 -3460 0 net=2477
rlabel metal2 751 -3460 751 -3460 0 net=6215
rlabel metal2 765 -3460 765 -3460 0 net=8731
rlabel metal2 765 -3460 765 -3460 0 net=8731
rlabel metal2 779 -3460 779 -3460 0 net=5923
rlabel metal2 877 -3460 877 -3460 0 net=9034
rlabel metal2 905 -3460 905 -3460 0 net=11265
rlabel metal2 919 -3460 919 -3460 0 net=11017
rlabel metal2 919 -3460 919 -3460 0 net=11017
rlabel metal2 926 -3460 926 -3460 0 net=9735
rlabel metal2 933 -3460 933 -3460 0 net=7589
rlabel metal2 940 -3460 940 -3460 0 net=9239
rlabel metal2 954 -3460 954 -3460 0 net=11219
rlabel metal2 436 -3462 436 -3462 0 net=4773
rlabel metal2 520 -3462 520 -3462 0 net=3652
rlabel metal2 653 -3462 653 -3462 0 net=7191
rlabel metal2 751 -3462 751 -3462 0 net=6321
rlabel metal2 779 -3462 779 -3462 0 net=4923
rlabel metal2 835 -3462 835 -3462 0 net=8934
rlabel metal2 891 -3462 891 -3462 0 net=5495
rlabel metal2 926 -3462 926 -3462 0 net=9951
rlabel metal2 527 -3464 527 -3464 0 net=5636
rlabel metal2 590 -3464 590 -3464 0 net=2889
rlabel metal2 660 -3464 660 -3464 0 net=5351
rlabel metal2 695 -3464 695 -3464 0 net=6018
rlabel metal2 772 -3464 772 -3464 0 net=6511
rlabel metal2 933 -3464 933 -3464 0 net=12017
rlabel metal2 425 -3466 425 -3466 0 net=7269
rlabel metal2 530 -3466 530 -3466 0 net=11737
rlabel metal2 674 -3466 674 -3466 0 net=7165
rlabel metal2 772 -3466 772 -3466 0 net=11081
rlabel metal2 940 -3466 940 -3466 0 net=10123
rlabel metal2 954 -3466 954 -3466 0 net=8488
rlabel metal2 443 -3468 443 -3468 0 net=11533
rlabel metal2 786 -3468 786 -3468 0 net=8345
rlabel metal2 1342 -3468 1342 -3468 0 net=1
rlabel metal2 443 -3470 443 -3470 0 net=4261
rlabel metal2 506 -3470 506 -3470 0 net=5577
rlabel metal2 562 -3470 562 -3470 0 net=11720
rlabel metal2 793 -3470 793 -3470 0 net=6932
rlabel metal2 828 -3470 828 -3470 0 net=9785
rlabel metal2 422 -3472 422 -3472 0 net=8821
rlabel metal2 618 -3472 618 -3472 0 net=6923
rlabel metal2 723 -3472 723 -3472 0 net=10821
rlabel metal2 446 -3474 446 -3474 0 net=5313
rlabel metal2 583 -3474 583 -3474 0 net=11115
rlabel metal2 800 -3474 800 -3474 0 net=9121
rlabel metal2 457 -3476 457 -3476 0 net=4823
rlabel metal2 709 -3476 709 -3476 0 net=8553
rlabel metal2 807 -3476 807 -3476 0 net=11791
rlabel metal2 485 -3478 485 -3478 0 net=6295
rlabel metal2 709 -3478 709 -3478 0 net=8955
rlabel metal2 814 -3478 814 -3478 0 net=5775
rlabel metal2 541 -3480 541 -3480 0 net=3305
rlabel metal2 695 -3480 695 -3480 0 net=7109
rlabel metal2 569 -3482 569 -3482 0 net=8575
rlabel metal2 716 -3482 716 -3482 0 net=7603
rlabel metal2 555 -3484 555 -3484 0 net=5467
rlabel metal2 639 -3484 639 -3484 0 net=7393
rlabel metal2 492 -3486 492 -3486 0 net=3775
rlabel metal2 639 -3486 639 -3486 0 net=6473
rlabel metal2 429 -3488 429 -3488 0 net=5650
rlabel metal2 394 -3490 394 -3490 0 net=5027
rlabel metal2 352 -3492 352 -3492 0 net=9517
rlabel metal2 352 -3494 352 -3494 0 net=6457
rlabel metal2 373 -3496 373 -3496 0 net=2357
rlabel metal2 415 -3498 415 -3498 0 net=1555
rlabel metal2 247 -3509 247 -3509 0 net=3947
rlabel metal2 247 -3509 247 -3509 0 net=3947
rlabel metal2 254 -3509 254 -3509 0 net=5731
rlabel metal2 352 -3509 352 -3509 0 net=6458
rlabel metal2 555 -3509 555 -3509 0 net=3776
rlabel metal2 639 -3509 639 -3509 0 net=6666
rlabel metal2 691 -3509 691 -3509 0 net=11082
rlabel metal2 821 -3509 821 -3509 0 net=10822
rlabel metal2 940 -3509 940 -3509 0 net=10124
rlabel metal2 940 -3509 940 -3509 0 net=10124
rlabel metal2 947 -3509 947 -3509 0 net=9240
rlabel metal2 968 -3509 968 -3509 0 net=9737
rlabel metal2 982 -3509 982 -3509 0 net=11220
rlabel metal2 1052 -3509 1052 -3509 0 net=8395
rlabel metal2 1052 -3509 1052 -3509 0 net=8395
rlabel metal2 1059 -3509 1059 -3509 0 net=5987
rlabel metal2 1108 -3509 1108 -3509 0 net=10845
rlabel metal2 1108 -3509 1108 -3509 0 net=10845
rlabel metal2 1122 -3509 1122 -3509 0 net=7470
rlabel metal2 1171 -3509 1171 -3509 0 net=11288
rlabel metal2 1339 -3509 1339 -3509 0 net=12110
rlabel metal2 261 -3511 261 -3511 0 net=3071
rlabel metal2 261 -3511 261 -3511 0 net=3071
rlabel metal2 268 -3511 268 -3511 0 net=7897
rlabel metal2 401 -3511 401 -3511 0 net=4324
rlabel metal2 429 -3511 429 -3511 0 net=5028
rlabel metal2 576 -3511 576 -3511 0 net=4802
rlabel metal2 611 -3511 611 -3511 0 net=8363
rlabel metal2 611 -3511 611 -3511 0 net=8363
rlabel metal2 618 -3511 618 -3511 0 net=6924
rlabel metal2 653 -3511 653 -3511 0 net=2890
rlabel metal2 702 -3511 702 -3511 0 net=7193
rlabel metal2 702 -3511 702 -3511 0 net=7193
rlabel metal2 709 -3511 709 -3511 0 net=8957
rlabel metal2 709 -3511 709 -3511 0 net=8957
rlabel metal2 730 -3511 730 -3511 0 net=7605
rlabel metal2 751 -3511 751 -3511 0 net=6323
rlabel metal2 751 -3511 751 -3511 0 net=6323
rlabel metal2 758 -3511 758 -3511 0 net=6217
rlabel metal2 758 -3511 758 -3511 0 net=6217
rlabel metal2 765 -3511 765 -3511 0 net=8733
rlabel metal2 765 -3511 765 -3511 0 net=8733
rlabel metal2 849 -3511 849 -3511 0 net=6475
rlabel metal2 905 -3511 905 -3511 0 net=11267
rlabel metal2 905 -3511 905 -3511 0 net=11267
rlabel metal2 933 -3511 933 -3511 0 net=12019
rlabel metal2 961 -3511 961 -3511 0 net=7591
rlabel metal2 989 -3511 989 -3511 0 net=10401
rlabel metal2 989 -3511 989 -3511 0 net=10401
rlabel metal2 996 -3511 996 -3511 0 net=10482
rlabel metal2 1080 -3511 1080 -3511 0 net=10421
rlabel metal2 1080 -3511 1080 -3511 0 net=10421
rlabel metal2 1150 -3511 1150 -3511 0 net=9913
rlabel metal2 1150 -3511 1150 -3511 0 net=9913
rlabel metal2 1346 -3511 1346 -3511 0 net=10974
rlabel metal2 387 -3513 387 -3513 0 net=3505
rlabel metal2 422 -3513 422 -3513 0 net=4652
rlabel metal2 495 -3513 495 -3513 0 net=1024
rlabel metal2 660 -3513 660 -3513 0 net=11739
rlabel metal2 730 -3513 730 -3513 0 net=2479
rlabel metal2 842 -3513 842 -3513 0 net=9123
rlabel metal2 870 -3513 870 -3513 0 net=8347
rlabel metal2 912 -3513 912 -3513 0 net=5496
rlabel metal2 1003 -3513 1003 -3513 0 net=11055
rlabel metal2 373 -3515 373 -3515 0 net=2359
rlabel metal2 429 -3515 429 -3515 0 net=2749
rlabel metal2 667 -3515 667 -3515 0 net=2452
rlabel metal2 737 -3515 737 -3515 0 net=7167
rlabel metal2 856 -3515 856 -3515 0 net=9787
rlabel metal2 877 -3515 877 -3515 0 net=5777
rlabel metal2 912 -3515 912 -3515 0 net=9953
rlabel metal2 450 -3517 450 -3517 0 net=5102
rlabel metal2 499 -3517 499 -3517 0 net=5315
rlabel metal2 548 -3517 548 -3517 0 net=3805
rlabel metal2 590 -3517 590 -3517 0 net=11535
rlabel metal2 667 -3517 667 -3517 0 net=11793
rlabel metal2 863 -3517 863 -3517 0 net=5925
rlabel metal2 919 -3517 919 -3517 0 net=11019
rlabel metal2 394 -3519 394 -3519 0 net=9518
rlabel metal2 453 -3519 453 -3519 0 net=2011
rlabel metal2 485 -3519 485 -3519 0 net=6297
rlabel metal2 499 -3519 499 -3519 0 net=11575
rlabel metal2 597 -3519 597 -3519 0 net=2648
rlabel metal2 674 -3519 674 -3519 0 net=5352
rlabel metal2 835 -3519 835 -3519 0 net=6513
rlabel metal2 359 -3521 359 -3521 0 net=3277
rlabel metal2 457 -3521 457 -3521 0 net=4825
rlabel metal2 555 -3521 555 -3521 0 net=8577
rlabel metal2 600 -3521 600 -3521 0 net=4290
rlabel metal2 677 -3521 677 -3521 0 net=1459
rlabel metal2 338 -3523 338 -3523 0 net=2427
rlabel metal2 408 -3523 408 -3523 0 net=5609
rlabel metal2 471 -3523 471 -3523 0 net=4971
rlabel metal2 471 -3523 471 -3523 0 net=4971
rlabel metal2 506 -3523 506 -3523 0 net=8823
rlabel metal2 506 -3523 506 -3523 0 net=8823
rlabel metal2 513 -3523 513 -3523 0 net=5423
rlabel metal2 569 -3523 569 -3523 0 net=11117
rlabel metal2 632 -3523 632 -3523 0 net=5469
rlabel metal2 800 -3523 800 -3523 0 net=8555
rlabel metal2 408 -3525 408 -3525 0 net=3691
rlabel metal2 467 -3525 467 -3525 0 net=5029
rlabel metal2 443 -3527 443 -3527 0 net=4263
rlabel metal2 520 -3527 520 -3527 0 net=7270
rlabel metal2 366 -3529 366 -3529 0 net=2170
rlabel metal2 464 -3529 464 -3529 0 net=2403
rlabel metal2 436 -3531 436 -3531 0 net=4775
rlabel metal2 527 -3531 527 -3531 0 net=5579
rlabel metal2 415 -3533 415 -3533 0 net=1557
rlabel metal2 527 -3533 527 -3533 0 net=3307
rlabel metal2 380 -3535 380 -3535 0 net=3473
rlabel metal2 541 -3535 541 -3535 0 net=7110
rlabel metal2 345 -3537 345 -3537 0 net=1731
rlabel metal2 695 -3537 695 -3537 0 net=7395
rlabel metal2 331 -3539 331 -3539 0 net=3461
rlabel metal2 716 -3539 716 -3539 0 net=4925
rlabel metal2 247 -3550 247 -3550 0 net=3948
rlabel metal2 261 -3550 261 -3550 0 net=3072
rlabel metal2 261 -3550 261 -3550 0 net=3072
rlabel metal2 268 -3550 268 -3550 0 net=7899
rlabel metal2 268 -3550 268 -3550 0 net=7899
rlabel metal2 296 -3550 296 -3550 0 net=5733
rlabel metal2 327 -3550 327 -3550 0 net=6933
rlabel metal2 394 -3550 394 -3550 0 net=3278
rlabel metal2 457 -3550 457 -3550 0 net=5610
rlabel metal2 604 -3550 604 -3550 0 net=2751
rlabel metal2 677 -3550 677 -3550 0 net=1871
rlabel metal2 968 -3550 968 -3550 0 net=7593
rlabel metal2 968 -3550 968 -3550 0 net=7593
rlabel metal2 975 -3550 975 -3550 0 net=9739
rlabel metal2 975 -3550 975 -3550 0 net=9739
rlabel metal2 989 -3550 989 -3550 0 net=10403
rlabel metal2 989 -3550 989 -3550 0 net=10403
rlabel metal2 1006 -3550 1006 -3550 0 net=11056
rlabel metal2 1038 -3550 1038 -3550 0 net=5989
rlabel metal2 1080 -3550 1080 -3550 0 net=10423
rlabel metal2 1108 -3550 1108 -3550 0 net=10847
rlabel metal2 1108 -3550 1108 -3550 0 net=10847
rlabel metal2 1150 -3550 1150 -3550 0 net=9914
rlabel metal2 345 -3552 345 -3552 0 net=3463
rlabel metal2 359 -3552 359 -3552 0 net=2429
rlabel metal2 359 -3552 359 -3552 0 net=2429
rlabel metal2 380 -3552 380 -3552 0 net=1733
rlabel metal2 401 -3552 401 -3552 0 net=3506
rlabel metal2 401 -3552 401 -3552 0 net=3506
rlabel metal2 443 -3552 443 -3552 0 net=5757
rlabel metal2 485 -3552 485 -3552 0 net=8824
rlabel metal2 520 -3552 520 -3552 0 net=4777
rlabel metal2 520 -3552 520 -3552 0 net=4777
rlabel metal2 544 -3552 544 -3552 0 net=3806
rlabel metal2 583 -3552 583 -3552 0 net=5031
rlabel metal2 611 -3552 611 -3552 0 net=8365
rlabel metal2 611 -3552 611 -3552 0 net=8365
rlabel metal2 618 -3552 618 -3552 0 net=11795
rlabel metal2 681 -3552 681 -3552 0 net=5471
rlabel metal2 695 -3552 695 -3552 0 net=7397
rlabel metal2 723 -3552 723 -3552 0 net=11741
rlabel metal2 765 -3552 765 -3552 0 net=8735
rlabel metal2 765 -3552 765 -3552 0 net=8735
rlabel metal2 849 -3552 849 -3552 0 net=9125
rlabel metal2 870 -3552 870 -3552 0 net=9788
rlabel metal2 905 -3552 905 -3552 0 net=11269
rlabel metal2 905 -3552 905 -3552 0 net=11269
rlabel metal2 912 -3552 912 -3552 0 net=9954
rlabel metal2 926 -3552 926 -3552 0 net=11021
rlabel metal2 926 -3552 926 -3552 0 net=11021
rlabel metal2 933 -3552 933 -3552 0 net=12020
rlabel metal2 1052 -3552 1052 -3552 0 net=8397
rlabel metal2 1052 -3552 1052 -3552 0 net=8397
rlabel metal2 488 -3554 488 -3554 0 net=5316
rlabel metal2 562 -3554 562 -3554 0 net=5424
rlabel metal2 639 -3554 639 -3554 0 net=11537
rlabel metal2 695 -3554 695 -3554 0 net=7195
rlabel metal2 723 -3554 723 -3554 0 net=2481
rlabel metal2 835 -3554 835 -3554 0 net=8557
rlabel metal2 863 -3554 863 -3554 0 net=6514
rlabel metal2 450 -3556 450 -3556 0 net=11215
rlabel metal2 702 -3556 702 -3556 0 net=4927
rlabel metal2 730 -3556 730 -3556 0 net=7607
rlabel metal2 884 -3556 884 -3556 0 net=8348
rlabel metal2 450 -3558 450 -3558 0 net=861
rlabel metal2 464 -3558 464 -3558 0 net=2404
rlabel metal2 492 -3558 492 -3558 0 net=6299
rlabel metal2 737 -3558 737 -3558 0 net=6325
rlabel metal2 891 -3558 891 -3558 0 net=5779
rlabel metal2 436 -3560 436 -3560 0 net=1559
rlabel metal2 478 -3560 478 -3560 0 net=2013
rlabel metal2 499 -3560 499 -3560 0 net=11577
rlabel metal2 751 -3560 751 -3560 0 net=6219
rlabel metal2 877 -3560 877 -3560 0 net=5927
rlabel metal2 898 -3560 898 -3560 0 net=6476
rlabel metal2 415 -3562 415 -3562 0 net=3475
rlabel metal2 471 -3562 471 -3562 0 net=4973
rlabel metal2 744 -3562 744 -3562 0 net=7169
rlabel metal2 408 -3564 408 -3564 0 net=3693
rlabel metal2 422 -3564 422 -3564 0 net=2361
rlabel metal2 478 -3564 478 -3564 0 net=8889
rlabel metal2 726 -3564 726 -3564 0 net=1
rlabel metal2 376 -3566 376 -3566 0 net=7705
rlabel metal2 541 -3566 541 -3566 0 net=8579
rlabel metal2 555 -3568 555 -3568 0 net=11119
rlabel metal2 548 -3570 548 -3570 0 net=4827
rlabel metal2 527 -3572 527 -3572 0 net=3309
rlabel metal2 513 -3574 513 -3574 0 net=4265
rlabel metal2 513 -3576 513 -3576 0 net=5580
rlabel metal2 264 -3587 264 -3587 0 net=7900
rlabel metal2 310 -3587 310 -3587 0 net=5734
rlabel metal2 352 -3587 352 -3587 0 net=3464
rlabel metal2 352 -3587 352 -3587 0 net=3464
rlabel metal2 359 -3587 359 -3587 0 net=2430
rlabel metal2 394 -3587 394 -3587 0 net=1735
rlabel metal2 408 -3587 408 -3587 0 net=7706
rlabel metal2 450 -3587 450 -3587 0 net=5758
rlabel metal2 492 -3587 492 -3587 0 net=2014
rlabel metal2 520 -3587 520 -3587 0 net=4778
rlabel metal2 562 -3587 562 -3587 0 net=11216
rlabel metal2 695 -3587 695 -3587 0 net=7197
rlabel metal2 695 -3587 695 -3587 0 net=7197
rlabel metal2 702 -3587 702 -3587 0 net=4929
rlabel metal2 702 -3587 702 -3587 0 net=4929
rlabel metal2 716 -3587 716 -3587 0 net=8961
rlabel metal2 716 -3587 716 -3587 0 net=8961
rlabel metal2 751 -3587 751 -3587 0 net=6221
rlabel metal2 758 -3587 758 -3587 0 net=7171
rlabel metal2 849 -3587 849 -3587 0 net=8559
rlabel metal2 905 -3587 905 -3587 0 net=11270
rlabel metal2 912 -3587 912 -3587 0 net=5781
rlabel metal2 926 -3587 926 -3587 0 net=11023
rlabel metal2 926 -3587 926 -3587 0 net=11023
rlabel metal2 940 -3587 940 -3587 0 net=1873
rlabel metal2 1052 -3587 1052 -3587 0 net=8399
rlabel metal2 1052 -3587 1052 -3587 0 net=8399
rlabel metal2 1083 -3587 1083 -3587 0 net=10424
rlabel metal2 1108 -3587 1108 -3587 0 net=10849
rlabel metal2 1108 -3587 1108 -3587 0 net=10849
rlabel metal2 324 -3589 324 -3589 0 net=1383
rlabel metal2 366 -3589 366 -3589 0 net=6934
rlabel metal2 408 -3589 408 -3589 0 net=3695
rlabel metal2 436 -3589 436 -3589 0 net=3477
rlabel metal2 471 -3589 471 -3589 0 net=2363
rlabel metal2 506 -3589 506 -3589 0 net=11579
rlabel metal2 534 -3589 534 -3589 0 net=6301
rlabel metal2 569 -3589 569 -3589 0 net=4829
rlabel metal2 597 -3589 597 -3589 0 net=5033
rlabel metal2 611 -3589 611 -3589 0 net=8366
rlabel metal2 646 -3589 646 -3589 0 net=2752
rlabel metal2 744 -3589 744 -3589 0 net=11742
rlabel metal2 856 -3589 856 -3589 0 net=9127
rlabel metal2 856 -3589 856 -3589 0 net=9127
rlabel metal2 891 -3589 891 -3589 0 net=5928
rlabel metal2 968 -3589 968 -3589 0 net=7594
rlabel metal2 985 -3589 985 -3589 0 net=10404
rlabel metal2 1031 -3589 1031 -3589 0 net=5991
rlabel metal2 443 -3591 443 -3591 0 net=8890
rlabel metal2 499 -3591 499 -3591 0 net=4975
rlabel metal2 516 -3591 516 -3591 0 net=8580
rlabel metal2 548 -3591 548 -3591 0 net=3311
rlabel metal2 597 -3591 597 -3591 0 net=11797
rlabel metal2 660 -3591 660 -3591 0 net=11538
rlabel metal2 737 -3591 737 -3591 0 net=6327
rlabel metal2 751 -3591 751 -3591 0 net=8737
rlabel metal2 975 -3591 975 -3591 0 net=9741
rlabel metal2 464 -3593 464 -3593 0 net=1561
rlabel metal2 548 -3593 548 -3593 0 net=11121
rlabel metal2 730 -3593 730 -3593 0 net=7609
rlabel metal2 901 -3593 901 -3593 0 net=3789
rlabel metal2 527 -3595 527 -3595 0 net=4267
rlabel metal2 723 -3595 723 -3595 0 net=2483
rlabel metal2 709 -3597 709 -3597 0 net=7399
rlabel metal2 688 -3599 688 -3599 0 net=5473
rlabel metal2 401 -3610 401 -3610 0 net=1737
rlabel metal2 457 -3610 457 -3610 0 net=3479
rlabel metal2 471 -3610 471 -3610 0 net=1563
rlabel metal2 471 -3610 471 -3610 0 net=1563
rlabel metal2 492 -3610 492 -3610 0 net=2364
rlabel metal2 520 -3610 520 -3610 0 net=11581
rlabel metal2 541 -3610 541 -3610 0 net=11122
rlabel metal2 555 -3610 555 -3610 0 net=4269
rlabel metal2 590 -3610 590 -3610 0 net=11799
rlabel metal2 604 -3610 604 -3610 0 net=5034
rlabel metal2 684 -3610 684 -3610 0 net=10675
rlabel metal2 856 -3610 856 -3610 0 net=9129
rlabel metal2 856 -3610 856 -3610 0 net=9129
rlabel metal2 863 -3610 863 -3610 0 net=8561
rlabel metal2 863 -3610 863 -3610 0 net=8561
rlabel metal2 926 -3610 926 -3610 0 net=11025
rlabel metal2 975 -3610 975 -3610 0 net=3791
rlabel metal2 1031 -3610 1031 -3610 0 net=5993
rlabel metal2 1031 -3610 1031 -3610 0 net=5993
rlabel metal2 1045 -3610 1045 -3610 0 net=1875
rlabel metal2 1108 -3610 1108 -3610 0 net=10851
rlabel metal2 1108 -3610 1108 -3610 0 net=10851
rlabel metal2 401 -3612 401 -3612 0 net=3697
rlabel metal2 506 -3612 506 -3612 0 net=4976
rlabel metal2 562 -3612 562 -3612 0 net=6303
rlabel metal2 562 -3612 562 -3612 0 net=6303
rlabel metal2 569 -3612 569 -3612 0 net=3313
rlabel metal2 569 -3612 569 -3612 0 net=3313
rlabel metal2 576 -3612 576 -3612 0 net=4831
rlabel metal2 576 -3612 576 -3612 0 net=4831
rlabel metal2 709 -3612 709 -3612 0 net=5475
rlabel metal2 730 -3612 730 -3612 0 net=2484
rlabel metal2 919 -3612 919 -3612 0 net=5783
rlabel metal2 982 -3612 982 -3612 0 net=9743
rlabel metal2 982 -3612 982 -3612 0 net=9743
rlabel metal2 1052 -3612 1052 -3612 0 net=8401
rlabel metal2 709 -3614 709 -3614 0 net=8963
rlabel metal2 751 -3614 751 -3614 0 net=8738
rlabel metal2 712 -3616 712 -3616 0 net=1
rlabel metal2 737 -3616 737 -3616 0 net=7611
rlabel metal2 758 -3616 758 -3616 0 net=6222
rlabel metal2 744 -3618 744 -3618 0 net=6329
rlabel metal2 765 -3618 765 -3618 0 net=7173
rlabel metal2 723 -3620 723 -3620 0 net=7401
rlabel metal2 702 -3622 702 -3622 0 net=4931
rlabel metal2 695 -3624 695 -3624 0 net=7199
rlabel metal2 401 -3635 401 -3635 0 net=3699
rlabel metal2 401 -3635 401 -3635 0 net=3699
rlabel metal2 408 -3635 408 -3635 0 net=1739
rlabel metal2 408 -3635 408 -3635 0 net=1739
rlabel metal2 464 -3635 464 -3635 0 net=3481
rlabel metal2 464 -3635 464 -3635 0 net=3481
rlabel metal2 471 -3635 471 -3635 0 net=1564
rlabel metal2 527 -3635 527 -3635 0 net=11583
rlabel metal2 527 -3635 527 -3635 0 net=11583
rlabel metal2 562 -3635 562 -3635 0 net=6304
rlabel metal2 583 -3635 583 -3635 0 net=4271
rlabel metal2 716 -3635 716 -3635 0 net=5476
rlabel metal2 716 -3635 716 -3635 0 net=5476
rlabel metal2 719 -3635 719 -3635 0 net=4932
rlabel metal2 744 -3635 744 -3635 0 net=7402
rlabel metal2 856 -3635 856 -3635 0 net=9130
rlabel metal2 863 -3635 863 -3635 0 net=8563
rlabel metal2 863 -3635 863 -3635 0 net=8563
rlabel metal2 926 -3635 926 -3635 0 net=5784
rlabel metal2 933 -3635 933 -3635 0 net=11027
rlabel metal2 933 -3635 933 -3635 0 net=11027
rlabel metal2 982 -3635 982 -3635 0 net=9745
rlabel metal2 1031 -3635 1031 -3635 0 net=5994
rlabel metal2 1055 -3635 1055 -3635 0 net=8402
rlabel metal2 1080 -3635 1080 -3635 0 net=1877
rlabel metal2 1108 -3635 1108 -3635 0 net=10852
rlabel metal2 576 -3637 576 -3637 0 net=4832
rlabel metal2 590 -3637 590 -3637 0 net=11801
rlabel metal2 590 -3637 590 -3637 0 net=11801
rlabel metal2 709 -3637 709 -3637 0 net=8965
rlabel metal2 751 -3637 751 -3637 0 net=7613
rlabel metal2 751 -3637 751 -3637 0 net=7613
rlabel metal2 758 -3637 758 -3637 0 net=6331
rlabel metal2 758 -3637 758 -3637 0 net=6331
rlabel metal2 765 -3637 765 -3637 0 net=7175
rlabel metal2 765 -3637 765 -3637 0 net=7175
rlabel metal2 800 -3637 800 -3637 0 net=10676
rlabel metal2 985 -3637 985 -3637 0 net=438
rlabel metal2 569 -3639 569 -3639 0 net=3315
rlabel metal2 702 -3639 702 -3639 0 net=7201
rlabel metal2 1003 -3639 1003 -3639 0 net=3792
rlabel metal2 401 -3650 401 -3650 0 net=3700
rlabel metal2 401 -3650 401 -3650 0 net=3700
rlabel metal2 408 -3650 408 -3650 0 net=1741
rlabel metal2 408 -3650 408 -3650 0 net=1741
rlabel metal2 464 -3650 464 -3650 0 net=3482
rlabel metal2 527 -3650 527 -3650 0 net=11585
rlabel metal2 569 -3650 569 -3650 0 net=3316
rlabel metal2 583 -3650 583 -3650 0 net=11802
rlabel metal2 709 -3650 709 -3650 0 net=7202
rlabel metal2 765 -3650 765 -3650 0 net=7177
rlabel metal2 856 -3650 856 -3650 0 net=8564
rlabel metal2 929 -3650 929 -3650 0 net=11028
rlabel metal2 985 -3650 985 -3650 0 net=9746
rlabel metal2 1094 -3650 1094 -3650 0 net=1878
rlabel metal2 586 -3652 586 -3652 0 net=4272
rlabel metal2 716 -3652 716 -3652 0 net=8966
rlabel metal2 758 -3652 758 -3652 0 net=6332
rlabel metal2 751 -3654 751 -3654 0 net=7615
rlabel metal2 404 -3665 404 -3665 0 net=1742
rlabel metal2 527 -3665 527 -3665 0 net=11586
rlabel metal2 758 -3665 758 -3665 0 net=7616
rlabel metal2 768 -3665 768 -3665 0 net=7178
<< end >>
