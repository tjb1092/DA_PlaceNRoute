magic
tech scmos
timestamp 1555017322 
<< pdiffusion >>
rect 155 -22 161 -16
rect 211 -22 217 -16
rect 239 -22 242 -16
rect 246 -22 249 -16
rect 260 -22 263 -16
rect 267 -22 273 -16
rect 274 -22 277 -16
rect 281 -22 287 -16
rect 337 -22 340 -16
rect 372 -22 375 -16
rect 379 -22 385 -16
rect 386 -22 389 -16
rect 393 -22 399 -16
rect 400 -22 406 -16
rect 407 -22 413 -16
rect 414 -22 417 -16
rect 421 -22 427 -16
rect 428 -22 431 -16
rect 456 -22 462 -16
rect 463 -22 469 -16
rect 477 -22 483 -16
rect 484 -22 487 -16
rect 498 -22 501 -16
rect 505 -22 508 -16
rect 512 -22 518 -16
rect 526 -22 529 -16
rect 547 -22 553 -16
rect 561 -22 567 -16
rect 568 -22 571 -16
rect 575 -22 578 -16
rect 582 -22 588 -16
rect 603 -22 609 -16
rect 638 -22 641 -16
rect 666 -22 669 -16
rect 680 -22 683 -16
rect 701 -22 707 -16
rect 708 -22 711 -16
rect 764 -22 767 -16
rect 799 -22 805 -16
rect 827 -22 830 -16
rect 148 -65 154 -59
rect 155 -65 161 -59
rect 162 -65 165 -59
rect 190 -65 193 -59
rect 218 -65 221 -59
rect 225 -65 228 -59
rect 232 -65 235 -59
rect 246 -65 249 -59
rect 253 -65 256 -59
rect 260 -65 263 -59
rect 267 -65 270 -59
rect 274 -65 277 -59
rect 281 -65 284 -59
rect 288 -65 294 -59
rect 295 -65 298 -59
rect 302 -65 305 -59
rect 309 -65 315 -59
rect 316 -65 319 -59
rect 323 -65 326 -59
rect 330 -65 333 -59
rect 337 -65 343 -59
rect 344 -65 350 -59
rect 351 -65 357 -59
rect 358 -65 361 -59
rect 365 -65 368 -59
rect 372 -65 375 -59
rect 379 -65 385 -59
rect 386 -65 389 -59
rect 393 -65 396 -59
rect 400 -65 403 -59
rect 407 -65 413 -59
rect 414 -65 420 -59
rect 421 -65 424 -59
rect 428 -65 431 -59
rect 435 -65 438 -59
rect 442 -65 445 -59
rect 449 -65 455 -59
rect 456 -65 459 -59
rect 463 -65 466 -59
rect 470 -65 473 -59
rect 477 -65 483 -59
rect 484 -65 487 -59
rect 491 -65 494 -59
rect 498 -65 504 -59
rect 505 -65 508 -59
rect 512 -65 515 -59
rect 519 -65 522 -59
rect 526 -65 529 -59
rect 533 -65 539 -59
rect 540 -65 543 -59
rect 547 -65 550 -59
rect 554 -65 560 -59
rect 561 -65 564 -59
rect 568 -65 571 -59
rect 575 -65 581 -59
rect 582 -65 585 -59
rect 589 -65 595 -59
rect 596 -65 599 -59
rect 603 -65 606 -59
rect 610 -65 613 -59
rect 617 -65 623 -59
rect 624 -65 627 -59
rect 631 -65 634 -59
rect 638 -65 641 -59
rect 645 -65 648 -59
rect 652 -65 655 -59
rect 659 -65 662 -59
rect 666 -65 672 -59
rect 673 -65 676 -59
rect 680 -65 683 -59
rect 687 -65 690 -59
rect 701 -65 704 -59
rect 715 -65 721 -59
rect 722 -65 725 -59
rect 750 -65 753 -59
rect 757 -65 760 -59
rect 771 -65 774 -59
rect 827 -65 830 -59
rect 848 -65 851 -59
rect 876 -65 879 -59
rect 904 -65 907 -59
rect 22 -126 25 -120
rect 29 -126 32 -120
rect 36 -126 39 -120
rect 43 -126 46 -120
rect 50 -126 53 -120
rect 57 -126 63 -120
rect 64 -126 70 -120
rect 71 -126 77 -120
rect 78 -126 81 -120
rect 85 -126 91 -120
rect 92 -126 95 -120
rect 99 -126 102 -120
rect 106 -126 109 -120
rect 113 -126 119 -120
rect 120 -126 123 -120
rect 127 -126 133 -120
rect 134 -126 137 -120
rect 141 -126 144 -120
rect 148 -126 151 -120
rect 155 -126 158 -120
rect 162 -126 165 -120
rect 169 -126 172 -120
rect 176 -126 179 -120
rect 183 -126 189 -120
rect 190 -126 196 -120
rect 197 -126 200 -120
rect 204 -126 207 -120
rect 211 -126 214 -120
rect 218 -126 221 -120
rect 225 -126 228 -120
rect 232 -126 235 -120
rect 239 -126 242 -120
rect 246 -126 249 -120
rect 253 -126 256 -120
rect 260 -126 263 -120
rect 267 -126 273 -120
rect 274 -126 277 -120
rect 281 -126 284 -120
rect 288 -126 291 -120
rect 295 -126 301 -120
rect 302 -126 305 -120
rect 309 -126 315 -120
rect 316 -126 319 -120
rect 323 -126 329 -120
rect 330 -126 333 -120
rect 337 -126 340 -120
rect 344 -126 347 -120
rect 351 -126 354 -120
rect 358 -126 364 -120
rect 365 -126 368 -120
rect 372 -126 375 -120
rect 379 -126 382 -120
rect 386 -126 389 -120
rect 393 -126 399 -120
rect 400 -126 406 -120
rect 407 -126 410 -120
rect 414 -126 417 -120
rect 421 -126 424 -120
rect 428 -126 431 -120
rect 435 -126 441 -120
rect 442 -126 445 -120
rect 449 -126 452 -120
rect 456 -126 459 -120
rect 463 -126 466 -120
rect 470 -126 473 -120
rect 477 -126 480 -120
rect 484 -126 487 -120
rect 491 -126 494 -120
rect 498 -126 501 -120
rect 505 -126 508 -120
rect 512 -126 515 -120
rect 519 -126 522 -120
rect 526 -126 532 -120
rect 533 -126 536 -120
rect 540 -126 543 -120
rect 547 -126 550 -120
rect 554 -126 557 -120
rect 561 -126 564 -120
rect 568 -126 571 -120
rect 575 -126 578 -120
rect 582 -126 585 -120
rect 589 -126 592 -120
rect 596 -126 599 -120
rect 603 -126 609 -120
rect 610 -126 613 -120
rect 617 -126 620 -120
rect 624 -126 627 -120
rect 631 -126 634 -120
rect 638 -126 641 -120
rect 645 -126 648 -120
rect 652 -126 655 -120
rect 659 -126 665 -120
rect 666 -126 669 -120
rect 673 -126 676 -120
rect 680 -126 683 -120
rect 687 -126 690 -120
rect 694 -126 697 -120
rect 701 -126 704 -120
rect 708 -126 711 -120
rect 715 -126 718 -120
rect 722 -126 725 -120
rect 729 -126 732 -120
rect 736 -126 739 -120
rect 743 -126 746 -120
rect 750 -126 753 -120
rect 757 -126 763 -120
rect 764 -126 767 -120
rect 771 -126 774 -120
rect 778 -126 781 -120
rect 785 -126 788 -120
rect 792 -126 795 -120
rect 799 -126 802 -120
rect 806 -126 809 -120
rect 813 -126 816 -120
rect 820 -126 823 -120
rect 848 -126 851 -120
rect 855 -126 858 -120
rect 869 -126 872 -120
rect 876 -126 879 -120
rect 939 -126 942 -120
rect 946 -126 949 -120
rect 1499 -126 1502 -120
rect 1506 -126 1512 -120
rect 8 -205 11 -199
rect 15 -205 18 -199
rect 22 -205 25 -199
rect 29 -205 32 -199
rect 36 -205 39 -199
rect 43 -205 46 -199
rect 50 -205 56 -199
rect 57 -205 60 -199
rect 64 -205 67 -199
rect 71 -205 74 -199
rect 78 -205 81 -199
rect 85 -205 88 -199
rect 92 -205 95 -199
rect 99 -205 105 -199
rect 106 -205 109 -199
rect 113 -205 116 -199
rect 120 -205 123 -199
rect 127 -205 130 -199
rect 134 -205 137 -199
rect 141 -205 147 -199
rect 148 -205 154 -199
rect 155 -205 161 -199
rect 162 -205 165 -199
rect 169 -205 172 -199
rect 176 -205 179 -199
rect 183 -205 186 -199
rect 190 -205 193 -199
rect 197 -205 200 -199
rect 204 -205 207 -199
rect 211 -205 214 -199
rect 218 -205 221 -199
rect 225 -205 228 -199
rect 232 -205 235 -199
rect 239 -205 245 -199
rect 246 -205 249 -199
rect 253 -205 256 -199
rect 260 -205 263 -199
rect 267 -205 273 -199
rect 274 -205 277 -199
rect 281 -205 284 -199
rect 288 -205 291 -199
rect 295 -205 298 -199
rect 302 -205 308 -199
rect 309 -205 312 -199
rect 316 -205 322 -199
rect 323 -205 326 -199
rect 330 -205 336 -199
rect 337 -205 340 -199
rect 344 -205 347 -199
rect 351 -205 354 -199
rect 358 -205 361 -199
rect 365 -205 368 -199
rect 372 -205 375 -199
rect 379 -205 382 -199
rect 386 -205 392 -199
rect 393 -205 396 -199
rect 400 -205 403 -199
rect 407 -205 410 -199
rect 414 -205 417 -199
rect 421 -205 424 -199
rect 428 -205 431 -199
rect 435 -205 441 -199
rect 442 -205 448 -199
rect 449 -205 452 -199
rect 456 -205 462 -199
rect 463 -205 466 -199
rect 470 -205 473 -199
rect 477 -205 480 -199
rect 484 -205 490 -199
rect 491 -205 494 -199
rect 498 -205 501 -199
rect 505 -205 508 -199
rect 512 -205 518 -199
rect 519 -205 522 -199
rect 526 -205 529 -199
rect 533 -205 539 -199
rect 540 -205 543 -199
rect 547 -205 550 -199
rect 554 -205 557 -199
rect 561 -205 564 -199
rect 568 -205 571 -199
rect 575 -205 578 -199
rect 582 -205 585 -199
rect 589 -205 592 -199
rect 596 -205 599 -199
rect 603 -205 609 -199
rect 610 -205 613 -199
rect 617 -205 620 -199
rect 624 -205 627 -199
rect 631 -205 634 -199
rect 638 -205 641 -199
rect 645 -205 648 -199
rect 652 -205 655 -199
rect 659 -205 662 -199
rect 666 -205 669 -199
rect 673 -205 676 -199
rect 680 -205 683 -199
rect 687 -205 690 -199
rect 694 -205 697 -199
rect 701 -205 704 -199
rect 708 -205 711 -199
rect 715 -205 721 -199
rect 722 -205 725 -199
rect 729 -205 732 -199
rect 736 -205 739 -199
rect 743 -205 746 -199
rect 750 -205 753 -199
rect 757 -205 760 -199
rect 764 -205 767 -199
rect 771 -205 774 -199
rect 778 -205 781 -199
rect 785 -205 788 -199
rect 792 -205 795 -199
rect 799 -205 802 -199
rect 806 -205 809 -199
rect 813 -205 816 -199
rect 820 -205 823 -199
rect 827 -205 830 -199
rect 834 -205 837 -199
rect 841 -205 844 -199
rect 848 -205 851 -199
rect 855 -205 858 -199
rect 862 -205 865 -199
rect 869 -205 872 -199
rect 876 -205 879 -199
rect 883 -205 886 -199
rect 890 -205 893 -199
rect 897 -205 900 -199
rect 904 -205 907 -199
rect 911 -205 914 -199
rect 918 -205 921 -199
rect 925 -205 928 -199
rect 932 -205 935 -199
rect 939 -205 942 -199
rect 946 -205 949 -199
rect 953 -205 956 -199
rect 960 -205 963 -199
rect 967 -205 970 -199
rect 974 -205 980 -199
rect 981 -205 987 -199
rect 988 -205 994 -199
rect 995 -205 998 -199
rect 1023 -205 1026 -199
rect 1499 -205 1502 -199
rect 1 -316 4 -310
rect 8 -316 11 -310
rect 15 -316 18 -310
rect 22 -316 28 -310
rect 29 -316 35 -310
rect 36 -316 42 -310
rect 43 -316 46 -310
rect 50 -316 56 -310
rect 57 -316 60 -310
rect 64 -316 70 -310
rect 71 -316 74 -310
rect 78 -316 84 -310
rect 85 -316 88 -310
rect 92 -316 98 -310
rect 99 -316 102 -310
rect 106 -316 109 -310
rect 113 -316 116 -310
rect 120 -316 126 -310
rect 127 -316 130 -310
rect 134 -316 137 -310
rect 141 -316 144 -310
rect 148 -316 151 -310
rect 155 -316 158 -310
rect 162 -316 165 -310
rect 169 -316 172 -310
rect 176 -316 179 -310
rect 183 -316 186 -310
rect 190 -316 193 -310
rect 197 -316 200 -310
rect 204 -316 207 -310
rect 211 -316 214 -310
rect 218 -316 221 -310
rect 225 -316 228 -310
rect 232 -316 235 -310
rect 239 -316 242 -310
rect 246 -316 249 -310
rect 253 -316 256 -310
rect 260 -316 263 -310
rect 267 -316 270 -310
rect 274 -316 277 -310
rect 281 -316 287 -310
rect 288 -316 291 -310
rect 295 -316 298 -310
rect 302 -316 305 -310
rect 309 -316 315 -310
rect 316 -316 322 -310
rect 323 -316 329 -310
rect 330 -316 333 -310
rect 337 -316 340 -310
rect 344 -316 347 -310
rect 351 -316 354 -310
rect 358 -316 364 -310
rect 365 -316 368 -310
rect 372 -316 375 -310
rect 379 -316 382 -310
rect 386 -316 389 -310
rect 393 -316 396 -310
rect 400 -316 403 -310
rect 407 -316 413 -310
rect 414 -316 417 -310
rect 421 -316 427 -310
rect 428 -316 431 -310
rect 435 -316 438 -310
rect 442 -316 445 -310
rect 449 -316 455 -310
rect 456 -316 459 -310
rect 463 -316 466 -310
rect 470 -316 473 -310
rect 477 -316 480 -310
rect 484 -316 487 -310
rect 491 -316 494 -310
rect 498 -316 501 -310
rect 505 -316 508 -310
rect 512 -316 515 -310
rect 519 -316 522 -310
rect 526 -316 529 -310
rect 533 -316 536 -310
rect 540 -316 546 -310
rect 547 -316 550 -310
rect 554 -316 557 -310
rect 561 -316 564 -310
rect 568 -316 571 -310
rect 575 -316 581 -310
rect 582 -316 588 -310
rect 589 -316 592 -310
rect 596 -316 599 -310
rect 603 -316 609 -310
rect 610 -316 613 -310
rect 617 -316 620 -310
rect 624 -316 627 -310
rect 631 -316 634 -310
rect 638 -316 641 -310
rect 645 -316 648 -310
rect 652 -316 655 -310
rect 659 -316 662 -310
rect 666 -316 669 -310
rect 673 -316 676 -310
rect 680 -316 683 -310
rect 687 -316 690 -310
rect 694 -316 700 -310
rect 701 -316 707 -310
rect 708 -316 711 -310
rect 715 -316 718 -310
rect 722 -316 725 -310
rect 729 -316 732 -310
rect 736 -316 739 -310
rect 743 -316 746 -310
rect 750 -316 753 -310
rect 757 -316 763 -310
rect 764 -316 767 -310
rect 771 -316 774 -310
rect 778 -316 781 -310
rect 785 -316 788 -310
rect 792 -316 795 -310
rect 799 -316 802 -310
rect 806 -316 809 -310
rect 813 -316 816 -310
rect 820 -316 823 -310
rect 827 -316 830 -310
rect 834 -316 837 -310
rect 841 -316 844 -310
rect 848 -316 851 -310
rect 855 -316 858 -310
rect 862 -316 865 -310
rect 869 -316 872 -310
rect 876 -316 879 -310
rect 883 -316 886 -310
rect 890 -316 893 -310
rect 897 -316 900 -310
rect 904 -316 907 -310
rect 911 -316 914 -310
rect 918 -316 921 -310
rect 925 -316 928 -310
rect 932 -316 935 -310
rect 939 -316 942 -310
rect 946 -316 949 -310
rect 953 -316 956 -310
rect 960 -316 963 -310
rect 967 -316 970 -310
rect 974 -316 977 -310
rect 981 -316 984 -310
rect 988 -316 991 -310
rect 995 -316 998 -310
rect 1002 -316 1005 -310
rect 1009 -316 1012 -310
rect 1016 -316 1019 -310
rect 1023 -316 1026 -310
rect 1030 -316 1033 -310
rect 1037 -316 1040 -310
rect 1044 -316 1047 -310
rect 1051 -316 1054 -310
rect 1058 -316 1061 -310
rect 1065 -316 1068 -310
rect 1072 -316 1075 -310
rect 1079 -316 1082 -310
rect 1086 -316 1089 -310
rect 1093 -316 1096 -310
rect 1100 -316 1103 -310
rect 1107 -316 1110 -310
rect 1114 -316 1117 -310
rect 1121 -316 1124 -310
rect 1128 -316 1131 -310
rect 1135 -316 1138 -310
rect 1142 -316 1145 -310
rect 1149 -316 1155 -310
rect 1177 -316 1180 -310
rect 1499 -316 1502 -310
rect 1 -405 4 -399
rect 8 -405 11 -399
rect 15 -405 18 -399
rect 22 -405 28 -399
rect 29 -405 32 -399
rect 36 -405 42 -399
rect 43 -405 49 -399
rect 50 -405 53 -399
rect 57 -405 63 -399
rect 64 -405 67 -399
rect 71 -405 77 -399
rect 78 -405 84 -399
rect 85 -405 91 -399
rect 92 -405 95 -399
rect 99 -405 102 -399
rect 106 -405 109 -399
rect 113 -405 116 -399
rect 120 -405 126 -399
rect 127 -405 130 -399
rect 134 -405 137 -399
rect 141 -405 144 -399
rect 148 -405 151 -399
rect 155 -405 158 -399
rect 162 -405 165 -399
rect 169 -405 172 -399
rect 176 -405 179 -399
rect 183 -405 186 -399
rect 190 -405 193 -399
rect 197 -405 200 -399
rect 204 -405 207 -399
rect 211 -405 214 -399
rect 218 -405 221 -399
rect 225 -405 228 -399
rect 232 -405 235 -399
rect 239 -405 242 -399
rect 246 -405 249 -399
rect 253 -405 256 -399
rect 260 -405 266 -399
rect 267 -405 270 -399
rect 274 -405 277 -399
rect 281 -405 284 -399
rect 288 -405 294 -399
rect 295 -405 298 -399
rect 302 -405 305 -399
rect 309 -405 312 -399
rect 316 -405 319 -399
rect 323 -405 326 -399
rect 330 -405 333 -399
rect 337 -405 340 -399
rect 344 -405 347 -399
rect 351 -405 354 -399
rect 358 -405 361 -399
rect 365 -405 368 -399
rect 372 -405 375 -399
rect 379 -405 382 -399
rect 386 -405 389 -399
rect 393 -405 399 -399
rect 400 -405 403 -399
rect 407 -405 413 -399
rect 414 -405 417 -399
rect 421 -405 424 -399
rect 428 -405 431 -399
rect 435 -405 438 -399
rect 442 -405 445 -399
rect 449 -405 452 -399
rect 456 -405 459 -399
rect 463 -405 466 -399
rect 470 -405 473 -399
rect 477 -405 480 -399
rect 484 -405 487 -399
rect 491 -405 494 -399
rect 498 -405 504 -399
rect 505 -405 511 -399
rect 512 -405 518 -399
rect 519 -405 522 -399
rect 526 -405 529 -399
rect 533 -405 536 -399
rect 540 -405 543 -399
rect 547 -405 553 -399
rect 554 -405 557 -399
rect 561 -405 567 -399
rect 568 -405 574 -399
rect 575 -405 578 -399
rect 582 -405 585 -399
rect 589 -405 595 -399
rect 596 -405 599 -399
rect 603 -405 606 -399
rect 610 -405 613 -399
rect 617 -405 620 -399
rect 624 -405 627 -399
rect 631 -405 634 -399
rect 638 -405 644 -399
rect 645 -405 648 -399
rect 652 -405 655 -399
rect 659 -405 665 -399
rect 666 -405 672 -399
rect 673 -405 676 -399
rect 680 -405 683 -399
rect 687 -405 690 -399
rect 694 -405 697 -399
rect 701 -405 704 -399
rect 708 -405 711 -399
rect 715 -405 718 -399
rect 722 -405 725 -399
rect 729 -405 732 -399
rect 736 -405 739 -399
rect 743 -405 746 -399
rect 750 -405 753 -399
rect 757 -405 760 -399
rect 764 -405 767 -399
rect 771 -405 774 -399
rect 778 -405 781 -399
rect 785 -405 788 -399
rect 792 -405 795 -399
rect 799 -405 802 -399
rect 806 -405 809 -399
rect 813 -405 816 -399
rect 820 -405 823 -399
rect 827 -405 830 -399
rect 834 -405 837 -399
rect 841 -405 844 -399
rect 848 -405 851 -399
rect 855 -405 858 -399
rect 862 -405 865 -399
rect 869 -405 872 -399
rect 876 -405 879 -399
rect 883 -405 886 -399
rect 890 -405 893 -399
rect 897 -405 900 -399
rect 904 -405 907 -399
rect 911 -405 914 -399
rect 918 -405 921 -399
rect 925 -405 928 -399
rect 932 -405 935 -399
rect 939 -405 942 -399
rect 946 -405 949 -399
rect 953 -405 956 -399
rect 960 -405 963 -399
rect 967 -405 970 -399
rect 974 -405 977 -399
rect 981 -405 984 -399
rect 988 -405 991 -399
rect 995 -405 998 -399
rect 1002 -405 1005 -399
rect 1009 -405 1012 -399
rect 1016 -405 1019 -399
rect 1023 -405 1026 -399
rect 1030 -405 1033 -399
rect 1037 -405 1040 -399
rect 1044 -405 1047 -399
rect 1051 -405 1054 -399
rect 1058 -405 1061 -399
rect 1065 -405 1068 -399
rect 1072 -405 1075 -399
rect 1079 -405 1082 -399
rect 1086 -405 1089 -399
rect 1093 -405 1096 -399
rect 1100 -405 1103 -399
rect 1107 -405 1110 -399
rect 1114 -405 1117 -399
rect 1121 -405 1124 -399
rect 1128 -405 1131 -399
rect 1135 -405 1138 -399
rect 1142 -405 1145 -399
rect 1149 -405 1152 -399
rect 1156 -405 1159 -399
rect 1163 -405 1166 -399
rect 1170 -405 1173 -399
rect 1177 -405 1180 -399
rect 1184 -405 1187 -399
rect 1191 -405 1194 -399
rect 1198 -405 1204 -399
rect 1205 -405 1211 -399
rect 1499 -405 1502 -399
rect 1 -520 7 -514
rect 8 -520 11 -514
rect 15 -520 18 -514
rect 22 -520 25 -514
rect 29 -520 35 -514
rect 36 -520 42 -514
rect 43 -520 46 -514
rect 50 -520 53 -514
rect 57 -520 60 -514
rect 64 -520 67 -514
rect 71 -520 77 -514
rect 78 -520 81 -514
rect 85 -520 91 -514
rect 92 -520 95 -514
rect 99 -520 102 -514
rect 106 -520 112 -514
rect 113 -520 116 -514
rect 120 -520 123 -514
rect 127 -520 130 -514
rect 134 -520 140 -514
rect 141 -520 147 -514
rect 148 -520 151 -514
rect 155 -520 161 -514
rect 162 -520 165 -514
rect 169 -520 172 -514
rect 176 -520 179 -514
rect 183 -520 186 -514
rect 190 -520 193 -514
rect 197 -520 203 -514
rect 204 -520 207 -514
rect 211 -520 214 -514
rect 218 -520 221 -514
rect 225 -520 228 -514
rect 232 -520 235 -514
rect 239 -520 242 -514
rect 246 -520 252 -514
rect 253 -520 259 -514
rect 260 -520 263 -514
rect 267 -520 270 -514
rect 274 -520 277 -514
rect 281 -520 284 -514
rect 288 -520 291 -514
rect 295 -520 298 -514
rect 302 -520 305 -514
rect 309 -520 312 -514
rect 316 -520 319 -514
rect 323 -520 326 -514
rect 330 -520 333 -514
rect 337 -520 340 -514
rect 344 -520 347 -514
rect 351 -520 354 -514
rect 358 -520 361 -514
rect 365 -520 368 -514
rect 372 -520 375 -514
rect 379 -520 385 -514
rect 386 -520 389 -514
rect 393 -520 396 -514
rect 400 -520 403 -514
rect 407 -520 410 -514
rect 414 -520 420 -514
rect 421 -520 427 -514
rect 428 -520 431 -514
rect 435 -520 438 -514
rect 442 -520 445 -514
rect 449 -520 452 -514
rect 456 -520 462 -514
rect 463 -520 466 -514
rect 470 -520 473 -514
rect 477 -520 480 -514
rect 484 -520 487 -514
rect 491 -520 494 -514
rect 498 -520 504 -514
rect 505 -520 511 -514
rect 512 -520 515 -514
rect 519 -520 522 -514
rect 526 -520 532 -514
rect 533 -520 539 -514
rect 540 -520 543 -514
rect 547 -520 550 -514
rect 554 -520 557 -514
rect 561 -520 564 -514
rect 568 -520 571 -514
rect 575 -520 578 -514
rect 582 -520 585 -514
rect 589 -520 592 -514
rect 596 -520 602 -514
rect 603 -520 606 -514
rect 610 -520 616 -514
rect 617 -520 620 -514
rect 624 -520 627 -514
rect 631 -520 634 -514
rect 638 -520 641 -514
rect 645 -520 648 -514
rect 652 -520 655 -514
rect 659 -520 665 -514
rect 666 -520 669 -514
rect 673 -520 676 -514
rect 680 -520 683 -514
rect 687 -520 690 -514
rect 694 -520 700 -514
rect 701 -520 707 -514
rect 708 -520 711 -514
rect 715 -520 718 -514
rect 722 -520 725 -514
rect 729 -520 732 -514
rect 736 -520 739 -514
rect 743 -520 746 -514
rect 750 -520 753 -514
rect 757 -520 760 -514
rect 764 -520 767 -514
rect 771 -520 774 -514
rect 778 -520 781 -514
rect 785 -520 788 -514
rect 792 -520 795 -514
rect 799 -520 802 -514
rect 806 -520 809 -514
rect 813 -520 816 -514
rect 820 -520 823 -514
rect 827 -520 830 -514
rect 834 -520 837 -514
rect 841 -520 844 -514
rect 848 -520 851 -514
rect 855 -520 858 -514
rect 862 -520 865 -514
rect 869 -520 872 -514
rect 876 -520 879 -514
rect 883 -520 886 -514
rect 890 -520 893 -514
rect 897 -520 900 -514
rect 904 -520 907 -514
rect 911 -520 914 -514
rect 918 -520 921 -514
rect 925 -520 928 -514
rect 932 -520 935 -514
rect 939 -520 942 -514
rect 946 -520 949 -514
rect 953 -520 956 -514
rect 960 -520 963 -514
rect 967 -520 970 -514
rect 974 -520 977 -514
rect 981 -520 984 -514
rect 988 -520 991 -514
rect 995 -520 998 -514
rect 1002 -520 1005 -514
rect 1009 -520 1012 -514
rect 1016 -520 1019 -514
rect 1023 -520 1026 -514
rect 1030 -520 1033 -514
rect 1037 -520 1040 -514
rect 1044 -520 1047 -514
rect 1051 -520 1054 -514
rect 1058 -520 1061 -514
rect 1065 -520 1068 -514
rect 1072 -520 1075 -514
rect 1079 -520 1082 -514
rect 1086 -520 1089 -514
rect 1093 -520 1096 -514
rect 1100 -520 1103 -514
rect 1107 -520 1110 -514
rect 1114 -520 1117 -514
rect 1121 -520 1124 -514
rect 1128 -520 1131 -514
rect 1135 -520 1138 -514
rect 1142 -520 1145 -514
rect 1149 -520 1152 -514
rect 1156 -520 1159 -514
rect 1163 -520 1166 -514
rect 1170 -520 1173 -514
rect 1177 -520 1180 -514
rect 1184 -520 1187 -514
rect 1191 -520 1194 -514
rect 1198 -520 1201 -514
rect 1205 -520 1208 -514
rect 1212 -520 1215 -514
rect 1219 -520 1222 -514
rect 1226 -520 1229 -514
rect 1233 -520 1236 -514
rect 1240 -520 1243 -514
rect 1247 -520 1250 -514
rect 1254 -520 1257 -514
rect 1261 -520 1264 -514
rect 1394 -520 1397 -514
rect 1499 -520 1502 -514
rect 1 -635 4 -629
rect 8 -635 11 -629
rect 15 -635 21 -629
rect 22 -635 25 -629
rect 29 -635 32 -629
rect 36 -635 42 -629
rect 43 -635 49 -629
rect 50 -635 53 -629
rect 57 -635 60 -629
rect 64 -635 67 -629
rect 71 -635 77 -629
rect 78 -635 81 -629
rect 85 -635 88 -629
rect 92 -635 98 -629
rect 99 -635 102 -629
rect 106 -635 109 -629
rect 113 -635 119 -629
rect 120 -635 123 -629
rect 127 -635 130 -629
rect 134 -635 137 -629
rect 141 -635 144 -629
rect 148 -635 151 -629
rect 155 -635 158 -629
rect 162 -635 165 -629
rect 169 -635 175 -629
rect 176 -635 179 -629
rect 183 -635 186 -629
rect 190 -635 193 -629
rect 197 -635 200 -629
rect 204 -635 207 -629
rect 211 -635 214 -629
rect 218 -635 221 -629
rect 225 -635 228 -629
rect 232 -635 235 -629
rect 239 -635 242 -629
rect 246 -635 249 -629
rect 253 -635 256 -629
rect 260 -635 263 -629
rect 267 -635 273 -629
rect 274 -635 277 -629
rect 281 -635 284 -629
rect 288 -635 291 -629
rect 295 -635 298 -629
rect 302 -635 305 -629
rect 309 -635 315 -629
rect 316 -635 319 -629
rect 323 -635 326 -629
rect 330 -635 333 -629
rect 337 -635 340 -629
rect 344 -635 350 -629
rect 351 -635 357 -629
rect 358 -635 361 -629
rect 365 -635 368 -629
rect 372 -635 375 -629
rect 379 -635 385 -629
rect 386 -635 392 -629
rect 393 -635 396 -629
rect 400 -635 403 -629
rect 407 -635 410 -629
rect 414 -635 420 -629
rect 421 -635 424 -629
rect 428 -635 431 -629
rect 435 -635 438 -629
rect 442 -635 448 -629
rect 449 -635 452 -629
rect 456 -635 459 -629
rect 463 -635 466 -629
rect 470 -635 473 -629
rect 477 -635 483 -629
rect 484 -635 487 -629
rect 491 -635 494 -629
rect 498 -635 501 -629
rect 505 -635 511 -629
rect 512 -635 515 -629
rect 519 -635 522 -629
rect 526 -635 529 -629
rect 533 -635 536 -629
rect 540 -635 543 -629
rect 547 -635 550 -629
rect 554 -635 557 -629
rect 561 -635 567 -629
rect 568 -635 571 -629
rect 575 -635 578 -629
rect 582 -635 585 -629
rect 589 -635 592 -629
rect 596 -635 599 -629
rect 603 -635 606 -629
rect 610 -635 616 -629
rect 617 -635 620 -629
rect 624 -635 630 -629
rect 631 -635 637 -629
rect 638 -635 641 -629
rect 645 -635 648 -629
rect 652 -635 655 -629
rect 659 -635 662 -629
rect 666 -635 672 -629
rect 673 -635 676 -629
rect 680 -635 683 -629
rect 687 -635 690 -629
rect 694 -635 697 -629
rect 701 -635 704 -629
rect 708 -635 711 -629
rect 715 -635 718 -629
rect 722 -635 725 -629
rect 729 -635 732 -629
rect 736 -635 739 -629
rect 743 -635 749 -629
rect 750 -635 753 -629
rect 757 -635 760 -629
rect 764 -635 767 -629
rect 771 -635 774 -629
rect 778 -635 781 -629
rect 785 -635 788 -629
rect 792 -635 795 -629
rect 799 -635 802 -629
rect 806 -635 809 -629
rect 813 -635 816 -629
rect 820 -635 823 -629
rect 827 -635 830 -629
rect 834 -635 837 -629
rect 841 -635 844 -629
rect 848 -635 851 -629
rect 855 -635 858 -629
rect 862 -635 865 -629
rect 869 -635 872 -629
rect 876 -635 879 -629
rect 883 -635 886 -629
rect 890 -635 893 -629
rect 897 -635 900 -629
rect 904 -635 907 -629
rect 911 -635 914 -629
rect 918 -635 921 -629
rect 925 -635 928 -629
rect 932 -635 935 -629
rect 939 -635 942 -629
rect 946 -635 949 -629
rect 953 -635 956 -629
rect 960 -635 966 -629
rect 967 -635 970 -629
rect 974 -635 977 -629
rect 981 -635 984 -629
rect 988 -635 991 -629
rect 995 -635 998 -629
rect 1002 -635 1005 -629
rect 1009 -635 1012 -629
rect 1016 -635 1019 -629
rect 1023 -635 1026 -629
rect 1030 -635 1036 -629
rect 1037 -635 1040 -629
rect 1044 -635 1047 -629
rect 1051 -635 1054 -629
rect 1058 -635 1061 -629
rect 1065 -635 1068 -629
rect 1072 -635 1075 -629
rect 1079 -635 1082 -629
rect 1086 -635 1089 -629
rect 1093 -635 1096 -629
rect 1100 -635 1103 -629
rect 1107 -635 1110 -629
rect 1114 -635 1117 -629
rect 1121 -635 1124 -629
rect 1128 -635 1131 -629
rect 1135 -635 1138 -629
rect 1142 -635 1145 -629
rect 1149 -635 1152 -629
rect 1156 -635 1159 -629
rect 1163 -635 1166 -629
rect 1170 -635 1173 -629
rect 1177 -635 1180 -629
rect 1184 -635 1187 -629
rect 1191 -635 1194 -629
rect 1198 -635 1201 -629
rect 1205 -635 1208 -629
rect 1212 -635 1215 -629
rect 1219 -635 1222 -629
rect 1226 -635 1229 -629
rect 1233 -635 1236 -629
rect 1240 -635 1243 -629
rect 1247 -635 1250 -629
rect 1254 -635 1257 -629
rect 1261 -635 1264 -629
rect 1268 -635 1271 -629
rect 1275 -635 1278 -629
rect 1282 -635 1285 -629
rect 1289 -635 1292 -629
rect 1296 -635 1299 -629
rect 1303 -635 1306 -629
rect 1310 -635 1313 -629
rect 1317 -635 1320 -629
rect 1324 -635 1327 -629
rect 1331 -635 1334 -629
rect 1338 -635 1341 -629
rect 1345 -635 1348 -629
rect 1352 -635 1355 -629
rect 1359 -635 1362 -629
rect 1366 -635 1369 -629
rect 1373 -635 1376 -629
rect 1471 -635 1474 -629
rect 1506 -635 1509 -629
rect 1 -754 7 -748
rect 8 -754 14 -748
rect 15 -754 18 -748
rect 22 -754 25 -748
rect 29 -754 32 -748
rect 36 -754 39 -748
rect 43 -754 46 -748
rect 50 -754 53 -748
rect 57 -754 63 -748
rect 64 -754 67 -748
rect 71 -754 77 -748
rect 78 -754 81 -748
rect 85 -754 88 -748
rect 92 -754 95 -748
rect 99 -754 105 -748
rect 106 -754 109 -748
rect 113 -754 119 -748
rect 120 -754 123 -748
rect 127 -754 130 -748
rect 134 -754 140 -748
rect 141 -754 144 -748
rect 148 -754 151 -748
rect 155 -754 158 -748
rect 162 -754 165 -748
rect 169 -754 172 -748
rect 176 -754 179 -748
rect 183 -754 186 -748
rect 190 -754 193 -748
rect 197 -754 200 -748
rect 204 -754 207 -748
rect 211 -754 214 -748
rect 218 -754 221 -748
rect 225 -754 228 -748
rect 232 -754 235 -748
rect 239 -754 242 -748
rect 246 -754 249 -748
rect 253 -754 256 -748
rect 260 -754 263 -748
rect 267 -754 273 -748
rect 274 -754 277 -748
rect 281 -754 284 -748
rect 288 -754 291 -748
rect 295 -754 298 -748
rect 302 -754 305 -748
rect 309 -754 312 -748
rect 316 -754 319 -748
rect 323 -754 326 -748
rect 330 -754 333 -748
rect 337 -754 340 -748
rect 344 -754 347 -748
rect 351 -754 357 -748
rect 358 -754 361 -748
rect 365 -754 371 -748
rect 372 -754 375 -748
rect 379 -754 382 -748
rect 386 -754 389 -748
rect 393 -754 396 -748
rect 400 -754 403 -748
rect 407 -754 410 -748
rect 414 -754 417 -748
rect 421 -754 427 -748
rect 428 -754 431 -748
rect 435 -754 438 -748
rect 442 -754 445 -748
rect 449 -754 452 -748
rect 456 -754 459 -748
rect 463 -754 466 -748
rect 470 -754 473 -748
rect 477 -754 480 -748
rect 484 -754 487 -748
rect 491 -754 494 -748
rect 498 -754 501 -748
rect 505 -754 508 -748
rect 512 -754 515 -748
rect 519 -754 525 -748
rect 526 -754 529 -748
rect 533 -754 539 -748
rect 540 -754 546 -748
rect 547 -754 550 -748
rect 554 -754 557 -748
rect 561 -754 567 -748
rect 568 -754 571 -748
rect 575 -754 578 -748
rect 582 -754 585 -748
rect 589 -754 592 -748
rect 596 -754 602 -748
rect 603 -754 606 -748
rect 610 -754 616 -748
rect 617 -754 623 -748
rect 624 -754 630 -748
rect 631 -754 634 -748
rect 638 -754 641 -748
rect 645 -754 648 -748
rect 652 -754 655 -748
rect 659 -754 665 -748
rect 666 -754 669 -748
rect 673 -754 676 -748
rect 680 -754 683 -748
rect 687 -754 690 -748
rect 694 -754 697 -748
rect 701 -754 704 -748
rect 708 -754 711 -748
rect 715 -754 718 -748
rect 722 -754 725 -748
rect 729 -754 732 -748
rect 736 -754 739 -748
rect 743 -754 749 -748
rect 750 -754 753 -748
rect 757 -754 763 -748
rect 764 -754 767 -748
rect 771 -754 777 -748
rect 778 -754 781 -748
rect 785 -754 788 -748
rect 792 -754 795 -748
rect 799 -754 802 -748
rect 806 -754 809 -748
rect 813 -754 816 -748
rect 820 -754 823 -748
rect 827 -754 830 -748
rect 834 -754 837 -748
rect 841 -754 844 -748
rect 848 -754 851 -748
rect 855 -754 858 -748
rect 862 -754 865 -748
rect 869 -754 872 -748
rect 876 -754 879 -748
rect 883 -754 889 -748
rect 890 -754 893 -748
rect 897 -754 900 -748
rect 904 -754 907 -748
rect 911 -754 914 -748
rect 918 -754 921 -748
rect 925 -754 928 -748
rect 932 -754 935 -748
rect 939 -754 945 -748
rect 946 -754 949 -748
rect 953 -754 956 -748
rect 960 -754 963 -748
rect 967 -754 970 -748
rect 974 -754 977 -748
rect 981 -754 984 -748
rect 988 -754 991 -748
rect 995 -754 998 -748
rect 1002 -754 1005 -748
rect 1009 -754 1012 -748
rect 1016 -754 1019 -748
rect 1023 -754 1026 -748
rect 1030 -754 1033 -748
rect 1037 -754 1040 -748
rect 1044 -754 1047 -748
rect 1051 -754 1054 -748
rect 1058 -754 1061 -748
rect 1065 -754 1068 -748
rect 1072 -754 1075 -748
rect 1079 -754 1082 -748
rect 1086 -754 1089 -748
rect 1093 -754 1096 -748
rect 1100 -754 1103 -748
rect 1107 -754 1110 -748
rect 1114 -754 1117 -748
rect 1121 -754 1124 -748
rect 1128 -754 1131 -748
rect 1135 -754 1138 -748
rect 1142 -754 1145 -748
rect 1149 -754 1152 -748
rect 1156 -754 1159 -748
rect 1163 -754 1166 -748
rect 1170 -754 1173 -748
rect 1177 -754 1180 -748
rect 1184 -754 1187 -748
rect 1191 -754 1194 -748
rect 1198 -754 1201 -748
rect 1205 -754 1208 -748
rect 1212 -754 1215 -748
rect 1219 -754 1222 -748
rect 1226 -754 1229 -748
rect 1233 -754 1236 -748
rect 1240 -754 1243 -748
rect 1247 -754 1250 -748
rect 1254 -754 1257 -748
rect 1261 -754 1264 -748
rect 1268 -754 1271 -748
rect 1275 -754 1278 -748
rect 1282 -754 1285 -748
rect 1289 -754 1292 -748
rect 1296 -754 1299 -748
rect 1303 -754 1306 -748
rect 1310 -754 1313 -748
rect 1317 -754 1320 -748
rect 1324 -754 1327 -748
rect 1331 -754 1334 -748
rect 1338 -754 1341 -748
rect 1345 -754 1348 -748
rect 1352 -754 1355 -748
rect 1359 -754 1362 -748
rect 1366 -754 1369 -748
rect 1373 -754 1376 -748
rect 1380 -754 1383 -748
rect 1387 -754 1390 -748
rect 1394 -754 1397 -748
rect 1401 -754 1404 -748
rect 1408 -754 1411 -748
rect 1415 -754 1418 -748
rect 1422 -754 1425 -748
rect 1429 -754 1432 -748
rect 1436 -754 1439 -748
rect 1443 -754 1446 -748
rect 1450 -754 1453 -748
rect 1457 -754 1460 -748
rect 1464 -754 1467 -748
rect 1471 -754 1474 -748
rect 1478 -754 1481 -748
rect 1485 -754 1488 -748
rect 1492 -754 1495 -748
rect 1499 -754 1502 -748
rect 1506 -754 1509 -748
rect 1513 -754 1516 -748
rect 1520 -754 1523 -748
rect 1527 -754 1530 -748
rect 1 -895 4 -889
rect 8 -895 11 -889
rect 15 -895 18 -889
rect 22 -895 25 -889
rect 29 -895 32 -889
rect 36 -895 42 -889
rect 43 -895 49 -889
rect 50 -895 53 -889
rect 57 -895 60 -889
rect 64 -895 67 -889
rect 71 -895 74 -889
rect 78 -895 81 -889
rect 85 -895 88 -889
rect 92 -895 95 -889
rect 99 -895 102 -889
rect 106 -895 109 -889
rect 113 -895 116 -889
rect 120 -895 123 -889
rect 127 -895 133 -889
rect 134 -895 137 -889
rect 141 -895 144 -889
rect 148 -895 151 -889
rect 155 -895 158 -889
rect 162 -895 168 -889
rect 169 -895 172 -889
rect 176 -895 179 -889
rect 183 -895 186 -889
rect 190 -895 193 -889
rect 197 -895 200 -889
rect 204 -895 207 -889
rect 211 -895 214 -889
rect 218 -895 221 -889
rect 225 -895 228 -889
rect 232 -895 238 -889
rect 239 -895 242 -889
rect 246 -895 249 -889
rect 253 -895 256 -889
rect 260 -895 263 -889
rect 267 -895 270 -889
rect 274 -895 277 -889
rect 281 -895 284 -889
rect 288 -895 291 -889
rect 295 -895 298 -889
rect 302 -895 305 -889
rect 309 -895 312 -889
rect 316 -895 319 -889
rect 323 -895 326 -889
rect 330 -895 333 -889
rect 337 -895 340 -889
rect 344 -895 347 -889
rect 351 -895 354 -889
rect 358 -895 361 -889
rect 365 -895 371 -889
rect 372 -895 375 -889
rect 379 -895 382 -889
rect 386 -895 389 -889
rect 393 -895 396 -889
rect 400 -895 403 -889
rect 407 -895 410 -889
rect 414 -895 417 -889
rect 421 -895 424 -889
rect 428 -895 431 -889
rect 435 -895 441 -889
rect 442 -895 445 -889
rect 449 -895 452 -889
rect 456 -895 462 -889
rect 463 -895 469 -889
rect 470 -895 473 -889
rect 477 -895 480 -889
rect 484 -895 487 -889
rect 491 -895 494 -889
rect 498 -895 501 -889
rect 505 -895 511 -889
rect 512 -895 515 -889
rect 519 -895 522 -889
rect 526 -895 529 -889
rect 533 -895 539 -889
rect 540 -895 546 -889
rect 547 -895 553 -889
rect 554 -895 557 -889
rect 561 -895 564 -889
rect 568 -895 571 -889
rect 575 -895 578 -889
rect 582 -895 585 -889
rect 589 -895 592 -889
rect 596 -895 599 -889
rect 603 -895 606 -889
rect 610 -895 613 -889
rect 617 -895 620 -889
rect 624 -895 627 -889
rect 631 -895 634 -889
rect 638 -895 644 -889
rect 645 -895 651 -889
rect 652 -895 658 -889
rect 659 -895 665 -889
rect 666 -895 669 -889
rect 673 -895 676 -889
rect 680 -895 683 -889
rect 687 -895 693 -889
rect 694 -895 697 -889
rect 701 -895 704 -889
rect 708 -895 714 -889
rect 715 -895 718 -889
rect 722 -895 725 -889
rect 729 -895 732 -889
rect 736 -895 739 -889
rect 743 -895 746 -889
rect 750 -895 753 -889
rect 757 -895 760 -889
rect 764 -895 770 -889
rect 771 -895 774 -889
rect 778 -895 781 -889
rect 785 -895 788 -889
rect 792 -895 795 -889
rect 799 -895 802 -889
rect 806 -895 812 -889
rect 813 -895 816 -889
rect 820 -895 823 -889
rect 827 -895 830 -889
rect 834 -895 840 -889
rect 841 -895 844 -889
rect 848 -895 851 -889
rect 855 -895 858 -889
rect 862 -895 865 -889
rect 869 -895 872 -889
rect 876 -895 879 -889
rect 883 -895 886 -889
rect 890 -895 893 -889
rect 897 -895 900 -889
rect 904 -895 907 -889
rect 911 -895 914 -889
rect 918 -895 921 -889
rect 925 -895 928 -889
rect 932 -895 935 -889
rect 939 -895 945 -889
rect 946 -895 949 -889
rect 953 -895 956 -889
rect 960 -895 963 -889
rect 967 -895 970 -889
rect 974 -895 977 -889
rect 981 -895 984 -889
rect 988 -895 991 -889
rect 995 -895 1001 -889
rect 1002 -895 1005 -889
rect 1009 -895 1012 -889
rect 1016 -895 1019 -889
rect 1023 -895 1026 -889
rect 1030 -895 1033 -889
rect 1037 -895 1040 -889
rect 1044 -895 1047 -889
rect 1051 -895 1054 -889
rect 1058 -895 1061 -889
rect 1065 -895 1068 -889
rect 1072 -895 1075 -889
rect 1079 -895 1082 -889
rect 1086 -895 1089 -889
rect 1093 -895 1096 -889
rect 1100 -895 1103 -889
rect 1107 -895 1110 -889
rect 1114 -895 1117 -889
rect 1121 -895 1124 -889
rect 1128 -895 1131 -889
rect 1135 -895 1138 -889
rect 1142 -895 1145 -889
rect 1149 -895 1152 -889
rect 1156 -895 1159 -889
rect 1163 -895 1166 -889
rect 1170 -895 1173 -889
rect 1177 -895 1180 -889
rect 1184 -895 1187 -889
rect 1191 -895 1194 -889
rect 1198 -895 1201 -889
rect 1205 -895 1208 -889
rect 1212 -895 1215 -889
rect 1219 -895 1222 -889
rect 1226 -895 1229 -889
rect 1233 -895 1236 -889
rect 1240 -895 1243 -889
rect 1247 -895 1250 -889
rect 1254 -895 1257 -889
rect 1261 -895 1264 -889
rect 1268 -895 1271 -889
rect 1275 -895 1278 -889
rect 1282 -895 1285 -889
rect 1289 -895 1292 -889
rect 1296 -895 1299 -889
rect 1303 -895 1306 -889
rect 1310 -895 1313 -889
rect 1317 -895 1320 -889
rect 1324 -895 1327 -889
rect 1331 -895 1334 -889
rect 1338 -895 1341 -889
rect 1345 -895 1348 -889
rect 1352 -895 1355 -889
rect 1359 -895 1362 -889
rect 1366 -895 1369 -889
rect 1373 -895 1376 -889
rect 1380 -895 1383 -889
rect 1387 -895 1390 -889
rect 1394 -895 1397 -889
rect 1401 -895 1404 -889
rect 1408 -895 1411 -889
rect 1415 -895 1418 -889
rect 1422 -895 1425 -889
rect 1429 -895 1432 -889
rect 1436 -895 1439 -889
rect 1443 -895 1446 -889
rect 1450 -895 1453 -889
rect 1457 -895 1460 -889
rect 1464 -895 1467 -889
rect 1471 -895 1474 -889
rect 1478 -895 1481 -889
rect 1485 -895 1488 -889
rect 1492 -895 1495 -889
rect 1499 -895 1505 -889
rect 1513 -895 1516 -889
rect 1 -1012 4 -1006
rect 8 -1012 11 -1006
rect 15 -1012 18 -1006
rect 22 -1012 25 -1006
rect 29 -1012 32 -1006
rect 36 -1012 39 -1006
rect 43 -1012 46 -1006
rect 50 -1012 53 -1006
rect 57 -1012 60 -1006
rect 64 -1012 67 -1006
rect 71 -1012 74 -1006
rect 78 -1012 81 -1006
rect 85 -1012 88 -1006
rect 92 -1012 98 -1006
rect 99 -1012 102 -1006
rect 106 -1012 109 -1006
rect 113 -1012 116 -1006
rect 120 -1012 123 -1006
rect 127 -1012 130 -1006
rect 134 -1012 137 -1006
rect 141 -1012 147 -1006
rect 148 -1012 151 -1006
rect 155 -1012 158 -1006
rect 162 -1012 165 -1006
rect 169 -1012 172 -1006
rect 176 -1012 179 -1006
rect 183 -1012 186 -1006
rect 190 -1012 193 -1006
rect 197 -1012 200 -1006
rect 204 -1012 207 -1006
rect 211 -1012 214 -1006
rect 218 -1012 221 -1006
rect 225 -1012 228 -1006
rect 232 -1012 235 -1006
rect 239 -1012 245 -1006
rect 246 -1012 249 -1006
rect 253 -1012 256 -1006
rect 260 -1012 263 -1006
rect 267 -1012 270 -1006
rect 274 -1012 277 -1006
rect 281 -1012 284 -1006
rect 288 -1012 291 -1006
rect 295 -1012 301 -1006
rect 302 -1012 305 -1006
rect 309 -1012 312 -1006
rect 316 -1012 319 -1006
rect 323 -1012 326 -1006
rect 330 -1012 336 -1006
rect 337 -1012 340 -1006
rect 344 -1012 347 -1006
rect 351 -1012 354 -1006
rect 358 -1012 361 -1006
rect 365 -1012 368 -1006
rect 372 -1012 378 -1006
rect 379 -1012 382 -1006
rect 386 -1012 389 -1006
rect 393 -1012 396 -1006
rect 400 -1012 403 -1006
rect 407 -1012 410 -1006
rect 414 -1012 417 -1006
rect 421 -1012 424 -1006
rect 428 -1012 431 -1006
rect 435 -1012 438 -1006
rect 442 -1012 445 -1006
rect 449 -1012 452 -1006
rect 456 -1012 459 -1006
rect 463 -1012 466 -1006
rect 470 -1012 473 -1006
rect 477 -1012 483 -1006
rect 484 -1012 487 -1006
rect 491 -1012 497 -1006
rect 498 -1012 501 -1006
rect 505 -1012 508 -1006
rect 512 -1012 515 -1006
rect 519 -1012 522 -1006
rect 526 -1012 529 -1006
rect 533 -1012 539 -1006
rect 540 -1012 546 -1006
rect 547 -1012 553 -1006
rect 554 -1012 557 -1006
rect 561 -1012 564 -1006
rect 568 -1012 571 -1006
rect 575 -1012 578 -1006
rect 582 -1012 585 -1006
rect 589 -1012 592 -1006
rect 596 -1012 602 -1006
rect 603 -1012 606 -1006
rect 610 -1012 613 -1006
rect 617 -1012 620 -1006
rect 624 -1012 627 -1006
rect 631 -1012 634 -1006
rect 638 -1012 641 -1006
rect 645 -1012 648 -1006
rect 652 -1012 655 -1006
rect 659 -1012 662 -1006
rect 666 -1012 669 -1006
rect 673 -1012 679 -1006
rect 680 -1012 683 -1006
rect 687 -1012 693 -1006
rect 694 -1012 697 -1006
rect 701 -1012 707 -1006
rect 708 -1012 711 -1006
rect 715 -1012 718 -1006
rect 722 -1012 725 -1006
rect 729 -1012 732 -1006
rect 736 -1012 739 -1006
rect 743 -1012 749 -1006
rect 750 -1012 756 -1006
rect 757 -1012 763 -1006
rect 764 -1012 767 -1006
rect 771 -1012 774 -1006
rect 778 -1012 781 -1006
rect 785 -1012 788 -1006
rect 792 -1012 795 -1006
rect 799 -1012 802 -1006
rect 806 -1012 809 -1006
rect 813 -1012 816 -1006
rect 820 -1012 826 -1006
rect 827 -1012 833 -1006
rect 834 -1012 837 -1006
rect 841 -1012 844 -1006
rect 848 -1012 851 -1006
rect 855 -1012 861 -1006
rect 862 -1012 865 -1006
rect 869 -1012 875 -1006
rect 876 -1012 879 -1006
rect 883 -1012 886 -1006
rect 890 -1012 893 -1006
rect 897 -1012 900 -1006
rect 904 -1012 910 -1006
rect 911 -1012 914 -1006
rect 918 -1012 921 -1006
rect 925 -1012 928 -1006
rect 932 -1012 935 -1006
rect 939 -1012 942 -1006
rect 946 -1012 949 -1006
rect 953 -1012 956 -1006
rect 960 -1012 963 -1006
rect 967 -1012 970 -1006
rect 974 -1012 977 -1006
rect 981 -1012 984 -1006
rect 988 -1012 994 -1006
rect 995 -1012 998 -1006
rect 1002 -1012 1005 -1006
rect 1009 -1012 1012 -1006
rect 1016 -1012 1019 -1006
rect 1023 -1012 1026 -1006
rect 1030 -1012 1033 -1006
rect 1037 -1012 1040 -1006
rect 1044 -1012 1047 -1006
rect 1051 -1012 1054 -1006
rect 1058 -1012 1061 -1006
rect 1065 -1012 1068 -1006
rect 1072 -1012 1075 -1006
rect 1079 -1012 1082 -1006
rect 1086 -1012 1089 -1006
rect 1093 -1012 1096 -1006
rect 1100 -1012 1103 -1006
rect 1107 -1012 1110 -1006
rect 1114 -1012 1117 -1006
rect 1121 -1012 1124 -1006
rect 1128 -1012 1131 -1006
rect 1135 -1012 1138 -1006
rect 1142 -1012 1145 -1006
rect 1149 -1012 1152 -1006
rect 1156 -1012 1159 -1006
rect 1163 -1012 1166 -1006
rect 1170 -1012 1173 -1006
rect 1177 -1012 1180 -1006
rect 1184 -1012 1187 -1006
rect 1191 -1012 1194 -1006
rect 1198 -1012 1201 -1006
rect 1205 -1012 1208 -1006
rect 1212 -1012 1215 -1006
rect 1219 -1012 1222 -1006
rect 1226 -1012 1229 -1006
rect 1233 -1012 1236 -1006
rect 1240 -1012 1243 -1006
rect 1247 -1012 1250 -1006
rect 1254 -1012 1257 -1006
rect 1261 -1012 1264 -1006
rect 1268 -1012 1271 -1006
rect 1275 -1012 1278 -1006
rect 1282 -1012 1285 -1006
rect 1289 -1012 1292 -1006
rect 1296 -1012 1299 -1006
rect 1303 -1012 1306 -1006
rect 1310 -1012 1313 -1006
rect 1317 -1012 1320 -1006
rect 1324 -1012 1327 -1006
rect 1331 -1012 1334 -1006
rect 1338 -1012 1341 -1006
rect 1345 -1012 1348 -1006
rect 1352 -1012 1355 -1006
rect 1359 -1012 1362 -1006
rect 1366 -1012 1369 -1006
rect 1373 -1012 1376 -1006
rect 1380 -1012 1383 -1006
rect 1387 -1012 1390 -1006
rect 1394 -1012 1397 -1006
rect 1401 -1012 1404 -1006
rect 1408 -1012 1411 -1006
rect 1415 -1012 1418 -1006
rect 1422 -1012 1428 -1006
rect 1429 -1012 1432 -1006
rect 1436 -1012 1439 -1006
rect 1443 -1012 1446 -1006
rect 1450 -1012 1453 -1006
rect 1457 -1012 1460 -1006
rect 1 -1159 4 -1153
rect 8 -1159 14 -1153
rect 15 -1159 18 -1153
rect 22 -1159 25 -1153
rect 29 -1159 35 -1153
rect 36 -1159 42 -1153
rect 43 -1159 46 -1153
rect 50 -1159 53 -1153
rect 57 -1159 60 -1153
rect 64 -1159 67 -1153
rect 71 -1159 74 -1153
rect 78 -1159 84 -1153
rect 85 -1159 88 -1153
rect 92 -1159 95 -1153
rect 99 -1159 102 -1153
rect 106 -1159 109 -1153
rect 113 -1159 116 -1153
rect 120 -1159 123 -1153
rect 127 -1159 130 -1153
rect 134 -1159 137 -1153
rect 141 -1159 144 -1153
rect 148 -1159 151 -1153
rect 155 -1159 158 -1153
rect 162 -1159 168 -1153
rect 169 -1159 172 -1153
rect 176 -1159 179 -1153
rect 183 -1159 186 -1153
rect 190 -1159 193 -1153
rect 197 -1159 203 -1153
rect 204 -1159 207 -1153
rect 211 -1159 214 -1153
rect 218 -1159 221 -1153
rect 225 -1159 228 -1153
rect 232 -1159 235 -1153
rect 239 -1159 242 -1153
rect 246 -1159 249 -1153
rect 253 -1159 256 -1153
rect 260 -1159 263 -1153
rect 267 -1159 270 -1153
rect 274 -1159 277 -1153
rect 281 -1159 284 -1153
rect 288 -1159 291 -1153
rect 295 -1159 298 -1153
rect 302 -1159 305 -1153
rect 309 -1159 312 -1153
rect 316 -1159 319 -1153
rect 323 -1159 326 -1153
rect 330 -1159 333 -1153
rect 337 -1159 340 -1153
rect 344 -1159 347 -1153
rect 351 -1159 357 -1153
rect 358 -1159 361 -1153
rect 365 -1159 368 -1153
rect 372 -1159 375 -1153
rect 379 -1159 382 -1153
rect 386 -1159 392 -1153
rect 393 -1159 396 -1153
rect 400 -1159 403 -1153
rect 407 -1159 410 -1153
rect 414 -1159 417 -1153
rect 421 -1159 424 -1153
rect 428 -1159 434 -1153
rect 435 -1159 438 -1153
rect 442 -1159 448 -1153
rect 449 -1159 452 -1153
rect 456 -1159 462 -1153
rect 463 -1159 466 -1153
rect 470 -1159 473 -1153
rect 477 -1159 480 -1153
rect 484 -1159 487 -1153
rect 491 -1159 494 -1153
rect 498 -1159 501 -1153
rect 505 -1159 508 -1153
rect 512 -1159 515 -1153
rect 519 -1159 522 -1153
rect 526 -1159 529 -1153
rect 533 -1159 536 -1153
rect 540 -1159 543 -1153
rect 547 -1159 550 -1153
rect 554 -1159 557 -1153
rect 561 -1159 564 -1153
rect 568 -1159 571 -1153
rect 575 -1159 578 -1153
rect 582 -1159 585 -1153
rect 589 -1159 595 -1153
rect 596 -1159 599 -1153
rect 603 -1159 609 -1153
rect 610 -1159 613 -1153
rect 617 -1159 620 -1153
rect 624 -1159 630 -1153
rect 631 -1159 634 -1153
rect 638 -1159 641 -1153
rect 645 -1159 648 -1153
rect 652 -1159 655 -1153
rect 659 -1159 665 -1153
rect 666 -1159 672 -1153
rect 673 -1159 676 -1153
rect 680 -1159 683 -1153
rect 687 -1159 690 -1153
rect 694 -1159 697 -1153
rect 701 -1159 704 -1153
rect 708 -1159 711 -1153
rect 715 -1159 721 -1153
rect 722 -1159 725 -1153
rect 729 -1159 735 -1153
rect 736 -1159 739 -1153
rect 743 -1159 746 -1153
rect 750 -1159 756 -1153
rect 757 -1159 760 -1153
rect 764 -1159 767 -1153
rect 771 -1159 774 -1153
rect 778 -1159 781 -1153
rect 785 -1159 788 -1153
rect 792 -1159 798 -1153
rect 799 -1159 802 -1153
rect 806 -1159 809 -1153
rect 813 -1159 816 -1153
rect 820 -1159 823 -1153
rect 827 -1159 833 -1153
rect 834 -1159 837 -1153
rect 841 -1159 844 -1153
rect 848 -1159 851 -1153
rect 855 -1159 861 -1153
rect 862 -1159 865 -1153
rect 869 -1159 872 -1153
rect 876 -1159 879 -1153
rect 883 -1159 886 -1153
rect 890 -1159 896 -1153
rect 897 -1159 900 -1153
rect 904 -1159 907 -1153
rect 911 -1159 914 -1153
rect 918 -1159 921 -1153
rect 925 -1159 928 -1153
rect 932 -1159 938 -1153
rect 939 -1159 942 -1153
rect 946 -1159 949 -1153
rect 953 -1159 959 -1153
rect 960 -1159 963 -1153
rect 967 -1159 970 -1153
rect 974 -1159 977 -1153
rect 981 -1159 984 -1153
rect 988 -1159 991 -1153
rect 995 -1159 998 -1153
rect 1002 -1159 1005 -1153
rect 1009 -1159 1012 -1153
rect 1016 -1159 1019 -1153
rect 1023 -1159 1026 -1153
rect 1030 -1159 1033 -1153
rect 1037 -1159 1040 -1153
rect 1044 -1159 1047 -1153
rect 1051 -1159 1054 -1153
rect 1058 -1159 1061 -1153
rect 1065 -1159 1068 -1153
rect 1072 -1159 1075 -1153
rect 1079 -1159 1082 -1153
rect 1086 -1159 1089 -1153
rect 1093 -1159 1096 -1153
rect 1100 -1159 1103 -1153
rect 1107 -1159 1110 -1153
rect 1114 -1159 1117 -1153
rect 1121 -1159 1124 -1153
rect 1128 -1159 1131 -1153
rect 1135 -1159 1138 -1153
rect 1142 -1159 1145 -1153
rect 1149 -1159 1152 -1153
rect 1156 -1159 1159 -1153
rect 1163 -1159 1166 -1153
rect 1170 -1159 1173 -1153
rect 1177 -1159 1180 -1153
rect 1184 -1159 1187 -1153
rect 1191 -1159 1194 -1153
rect 1198 -1159 1201 -1153
rect 1205 -1159 1208 -1153
rect 1212 -1159 1215 -1153
rect 1219 -1159 1222 -1153
rect 1226 -1159 1229 -1153
rect 1233 -1159 1236 -1153
rect 1240 -1159 1243 -1153
rect 1247 -1159 1250 -1153
rect 1254 -1159 1257 -1153
rect 1261 -1159 1264 -1153
rect 1268 -1159 1271 -1153
rect 1275 -1159 1278 -1153
rect 1282 -1159 1285 -1153
rect 1289 -1159 1292 -1153
rect 1296 -1159 1299 -1153
rect 1303 -1159 1306 -1153
rect 1310 -1159 1313 -1153
rect 1317 -1159 1320 -1153
rect 1324 -1159 1327 -1153
rect 1331 -1159 1334 -1153
rect 1338 -1159 1341 -1153
rect 1345 -1159 1348 -1153
rect 1352 -1159 1355 -1153
rect 1359 -1159 1362 -1153
rect 1366 -1159 1369 -1153
rect 1373 -1159 1376 -1153
rect 1380 -1159 1383 -1153
rect 1387 -1159 1390 -1153
rect 1394 -1159 1397 -1153
rect 1401 -1159 1404 -1153
rect 1408 -1159 1411 -1153
rect 1415 -1159 1418 -1153
rect 1422 -1159 1425 -1153
rect 1429 -1159 1432 -1153
rect 1436 -1159 1439 -1153
rect 1443 -1159 1446 -1153
rect 1450 -1159 1453 -1153
rect 1457 -1159 1460 -1153
rect 1464 -1159 1467 -1153
rect 1471 -1159 1474 -1153
rect 1478 -1159 1481 -1153
rect 1485 -1159 1488 -1153
rect 1492 -1159 1495 -1153
rect 1499 -1159 1502 -1153
rect 1506 -1159 1509 -1153
rect 1513 -1159 1516 -1153
rect 1520 -1159 1523 -1153
rect 1527 -1159 1530 -1153
rect 1534 -1159 1537 -1153
rect 1541 -1159 1544 -1153
rect 1548 -1159 1551 -1153
rect 1555 -1159 1558 -1153
rect 1562 -1159 1565 -1153
rect 1569 -1159 1572 -1153
rect 1576 -1159 1579 -1153
rect 1583 -1159 1586 -1153
rect 1590 -1159 1593 -1153
rect 1597 -1159 1600 -1153
rect 1 -1284 4 -1278
rect 8 -1284 11 -1278
rect 15 -1284 18 -1278
rect 22 -1284 25 -1278
rect 29 -1284 32 -1278
rect 36 -1284 39 -1278
rect 43 -1284 46 -1278
rect 50 -1284 53 -1278
rect 57 -1284 63 -1278
rect 64 -1284 67 -1278
rect 71 -1284 74 -1278
rect 78 -1284 81 -1278
rect 85 -1284 88 -1278
rect 92 -1284 95 -1278
rect 99 -1284 105 -1278
rect 106 -1284 109 -1278
rect 113 -1284 116 -1278
rect 120 -1284 123 -1278
rect 127 -1284 133 -1278
rect 134 -1284 137 -1278
rect 141 -1284 144 -1278
rect 148 -1284 151 -1278
rect 155 -1284 158 -1278
rect 162 -1284 165 -1278
rect 169 -1284 175 -1278
rect 176 -1284 179 -1278
rect 183 -1284 186 -1278
rect 190 -1284 193 -1278
rect 197 -1284 200 -1278
rect 204 -1284 207 -1278
rect 211 -1284 214 -1278
rect 218 -1284 221 -1278
rect 225 -1284 228 -1278
rect 232 -1284 235 -1278
rect 239 -1284 242 -1278
rect 246 -1284 249 -1278
rect 253 -1284 256 -1278
rect 260 -1284 263 -1278
rect 267 -1284 270 -1278
rect 274 -1284 277 -1278
rect 281 -1284 284 -1278
rect 288 -1284 291 -1278
rect 295 -1284 298 -1278
rect 302 -1284 305 -1278
rect 309 -1284 312 -1278
rect 316 -1284 322 -1278
rect 323 -1284 326 -1278
rect 330 -1284 333 -1278
rect 337 -1284 343 -1278
rect 344 -1284 347 -1278
rect 351 -1284 354 -1278
rect 358 -1284 364 -1278
rect 365 -1284 368 -1278
rect 372 -1284 375 -1278
rect 379 -1284 382 -1278
rect 386 -1284 389 -1278
rect 393 -1284 396 -1278
rect 400 -1284 403 -1278
rect 407 -1284 410 -1278
rect 414 -1284 417 -1278
rect 421 -1284 424 -1278
rect 428 -1284 431 -1278
rect 435 -1284 438 -1278
rect 442 -1284 445 -1278
rect 449 -1284 452 -1278
rect 456 -1284 459 -1278
rect 463 -1284 466 -1278
rect 470 -1284 473 -1278
rect 477 -1284 483 -1278
rect 484 -1284 487 -1278
rect 491 -1284 494 -1278
rect 498 -1284 501 -1278
rect 505 -1284 511 -1278
rect 512 -1284 515 -1278
rect 519 -1284 525 -1278
rect 526 -1284 532 -1278
rect 533 -1284 536 -1278
rect 540 -1284 543 -1278
rect 547 -1284 553 -1278
rect 554 -1284 560 -1278
rect 561 -1284 564 -1278
rect 568 -1284 571 -1278
rect 575 -1284 578 -1278
rect 582 -1284 585 -1278
rect 589 -1284 592 -1278
rect 596 -1284 599 -1278
rect 603 -1284 609 -1278
rect 610 -1284 613 -1278
rect 617 -1284 620 -1278
rect 624 -1284 627 -1278
rect 631 -1284 634 -1278
rect 638 -1284 641 -1278
rect 645 -1284 648 -1278
rect 652 -1284 655 -1278
rect 659 -1284 662 -1278
rect 666 -1284 669 -1278
rect 673 -1284 676 -1278
rect 680 -1284 683 -1278
rect 687 -1284 690 -1278
rect 694 -1284 697 -1278
rect 701 -1284 704 -1278
rect 708 -1284 711 -1278
rect 715 -1284 721 -1278
rect 722 -1284 728 -1278
rect 729 -1284 732 -1278
rect 736 -1284 739 -1278
rect 743 -1284 746 -1278
rect 750 -1284 756 -1278
rect 757 -1284 760 -1278
rect 764 -1284 770 -1278
rect 771 -1284 774 -1278
rect 778 -1284 784 -1278
rect 785 -1284 788 -1278
rect 792 -1284 795 -1278
rect 799 -1284 802 -1278
rect 806 -1284 809 -1278
rect 813 -1284 816 -1278
rect 820 -1284 823 -1278
rect 827 -1284 830 -1278
rect 834 -1284 840 -1278
rect 841 -1284 844 -1278
rect 848 -1284 851 -1278
rect 855 -1284 861 -1278
rect 862 -1284 865 -1278
rect 869 -1284 872 -1278
rect 876 -1284 879 -1278
rect 883 -1284 886 -1278
rect 890 -1284 893 -1278
rect 897 -1284 900 -1278
rect 904 -1284 907 -1278
rect 911 -1284 914 -1278
rect 918 -1284 924 -1278
rect 925 -1284 928 -1278
rect 932 -1284 938 -1278
rect 939 -1284 942 -1278
rect 946 -1284 949 -1278
rect 953 -1284 956 -1278
rect 960 -1284 963 -1278
rect 967 -1284 970 -1278
rect 974 -1284 977 -1278
rect 981 -1284 984 -1278
rect 988 -1284 991 -1278
rect 995 -1284 998 -1278
rect 1002 -1284 1005 -1278
rect 1009 -1284 1012 -1278
rect 1016 -1284 1019 -1278
rect 1023 -1284 1026 -1278
rect 1030 -1284 1033 -1278
rect 1037 -1284 1040 -1278
rect 1044 -1284 1047 -1278
rect 1051 -1284 1057 -1278
rect 1058 -1284 1061 -1278
rect 1065 -1284 1068 -1278
rect 1072 -1284 1075 -1278
rect 1079 -1284 1082 -1278
rect 1086 -1284 1089 -1278
rect 1093 -1284 1096 -1278
rect 1100 -1284 1103 -1278
rect 1107 -1284 1110 -1278
rect 1114 -1284 1117 -1278
rect 1121 -1284 1124 -1278
rect 1128 -1284 1131 -1278
rect 1135 -1284 1138 -1278
rect 1142 -1284 1145 -1278
rect 1149 -1284 1152 -1278
rect 1156 -1284 1159 -1278
rect 1163 -1284 1166 -1278
rect 1170 -1284 1176 -1278
rect 1177 -1284 1180 -1278
rect 1184 -1284 1187 -1278
rect 1191 -1284 1194 -1278
rect 1198 -1284 1201 -1278
rect 1205 -1284 1208 -1278
rect 1212 -1284 1215 -1278
rect 1219 -1284 1222 -1278
rect 1226 -1284 1229 -1278
rect 1233 -1284 1236 -1278
rect 1240 -1284 1243 -1278
rect 1247 -1284 1250 -1278
rect 1254 -1284 1257 -1278
rect 1261 -1284 1264 -1278
rect 1268 -1284 1271 -1278
rect 1275 -1284 1278 -1278
rect 1282 -1284 1285 -1278
rect 1289 -1284 1292 -1278
rect 1296 -1284 1299 -1278
rect 1303 -1284 1306 -1278
rect 1310 -1284 1313 -1278
rect 1317 -1284 1320 -1278
rect 1324 -1284 1327 -1278
rect 1331 -1284 1334 -1278
rect 1338 -1284 1341 -1278
rect 1345 -1284 1348 -1278
rect 1352 -1284 1355 -1278
rect 1359 -1284 1362 -1278
rect 1366 -1284 1369 -1278
rect 1373 -1284 1376 -1278
rect 1380 -1284 1383 -1278
rect 1387 -1284 1390 -1278
rect 1394 -1284 1397 -1278
rect 1401 -1284 1404 -1278
rect 1408 -1284 1411 -1278
rect 1415 -1284 1418 -1278
rect 1422 -1284 1425 -1278
rect 1429 -1284 1432 -1278
rect 1436 -1284 1439 -1278
rect 1443 -1284 1446 -1278
rect 1450 -1284 1453 -1278
rect 1457 -1284 1460 -1278
rect 1464 -1284 1467 -1278
rect 1471 -1284 1474 -1278
rect 1478 -1284 1481 -1278
rect 1485 -1284 1488 -1278
rect 1492 -1284 1495 -1278
rect 1499 -1284 1502 -1278
rect 1506 -1284 1509 -1278
rect 1513 -1284 1516 -1278
rect 1520 -1284 1523 -1278
rect 1527 -1284 1530 -1278
rect 1534 -1284 1537 -1278
rect 1541 -1284 1544 -1278
rect 1548 -1284 1551 -1278
rect 1555 -1284 1558 -1278
rect 1562 -1284 1565 -1278
rect 1 -1403 4 -1397
rect 8 -1403 11 -1397
rect 15 -1403 18 -1397
rect 22 -1403 25 -1397
rect 29 -1403 32 -1397
rect 36 -1403 39 -1397
rect 43 -1403 46 -1397
rect 50 -1403 53 -1397
rect 57 -1403 60 -1397
rect 64 -1403 70 -1397
rect 71 -1403 74 -1397
rect 78 -1403 84 -1397
rect 85 -1403 88 -1397
rect 92 -1403 95 -1397
rect 99 -1403 102 -1397
rect 106 -1403 112 -1397
rect 113 -1403 116 -1397
rect 120 -1403 123 -1397
rect 127 -1403 130 -1397
rect 134 -1403 137 -1397
rect 141 -1403 144 -1397
rect 148 -1403 151 -1397
rect 155 -1403 158 -1397
rect 162 -1403 165 -1397
rect 169 -1403 172 -1397
rect 176 -1403 179 -1397
rect 183 -1403 186 -1397
rect 190 -1403 193 -1397
rect 197 -1403 200 -1397
rect 204 -1403 207 -1397
rect 211 -1403 217 -1397
rect 218 -1403 221 -1397
rect 225 -1403 228 -1397
rect 232 -1403 235 -1397
rect 239 -1403 242 -1397
rect 246 -1403 249 -1397
rect 253 -1403 256 -1397
rect 260 -1403 263 -1397
rect 267 -1403 270 -1397
rect 274 -1403 277 -1397
rect 281 -1403 284 -1397
rect 288 -1403 291 -1397
rect 295 -1403 298 -1397
rect 302 -1403 305 -1397
rect 309 -1403 312 -1397
rect 316 -1403 322 -1397
rect 323 -1403 326 -1397
rect 330 -1403 333 -1397
rect 337 -1403 340 -1397
rect 344 -1403 347 -1397
rect 351 -1403 354 -1397
rect 358 -1403 361 -1397
rect 365 -1403 368 -1397
rect 372 -1403 375 -1397
rect 379 -1403 382 -1397
rect 386 -1403 392 -1397
rect 393 -1403 396 -1397
rect 400 -1403 406 -1397
rect 407 -1403 410 -1397
rect 414 -1403 420 -1397
rect 421 -1403 424 -1397
rect 428 -1403 431 -1397
rect 435 -1403 438 -1397
rect 442 -1403 445 -1397
rect 449 -1403 452 -1397
rect 456 -1403 459 -1397
rect 463 -1403 469 -1397
rect 470 -1403 473 -1397
rect 477 -1403 483 -1397
rect 484 -1403 490 -1397
rect 491 -1403 497 -1397
rect 498 -1403 501 -1397
rect 505 -1403 508 -1397
rect 512 -1403 518 -1397
rect 519 -1403 525 -1397
rect 526 -1403 529 -1397
rect 533 -1403 536 -1397
rect 540 -1403 543 -1397
rect 547 -1403 550 -1397
rect 554 -1403 557 -1397
rect 561 -1403 564 -1397
rect 568 -1403 571 -1397
rect 575 -1403 578 -1397
rect 582 -1403 585 -1397
rect 589 -1403 592 -1397
rect 596 -1403 599 -1397
rect 603 -1403 606 -1397
rect 610 -1403 613 -1397
rect 617 -1403 620 -1397
rect 624 -1403 627 -1397
rect 631 -1403 634 -1397
rect 638 -1403 641 -1397
rect 645 -1403 651 -1397
rect 652 -1403 655 -1397
rect 659 -1403 662 -1397
rect 666 -1403 669 -1397
rect 673 -1403 676 -1397
rect 680 -1403 683 -1397
rect 687 -1403 690 -1397
rect 694 -1403 697 -1397
rect 701 -1403 704 -1397
rect 708 -1403 714 -1397
rect 715 -1403 718 -1397
rect 722 -1403 725 -1397
rect 729 -1403 732 -1397
rect 736 -1403 739 -1397
rect 743 -1403 746 -1397
rect 750 -1403 753 -1397
rect 757 -1403 760 -1397
rect 764 -1403 767 -1397
rect 771 -1403 774 -1397
rect 778 -1403 781 -1397
rect 785 -1403 788 -1397
rect 792 -1403 795 -1397
rect 799 -1403 802 -1397
rect 806 -1403 809 -1397
rect 813 -1403 816 -1397
rect 820 -1403 823 -1397
rect 827 -1403 830 -1397
rect 834 -1403 837 -1397
rect 841 -1403 847 -1397
rect 848 -1403 851 -1397
rect 855 -1403 858 -1397
rect 862 -1403 865 -1397
rect 869 -1403 875 -1397
rect 876 -1403 882 -1397
rect 883 -1403 886 -1397
rect 890 -1403 893 -1397
rect 897 -1403 900 -1397
rect 904 -1403 907 -1397
rect 911 -1403 914 -1397
rect 918 -1403 924 -1397
rect 925 -1403 928 -1397
rect 932 -1403 935 -1397
rect 939 -1403 942 -1397
rect 946 -1403 952 -1397
rect 953 -1403 956 -1397
rect 960 -1403 963 -1397
rect 967 -1403 970 -1397
rect 974 -1403 980 -1397
rect 981 -1403 984 -1397
rect 988 -1403 991 -1397
rect 995 -1403 998 -1397
rect 1002 -1403 1008 -1397
rect 1009 -1403 1012 -1397
rect 1016 -1403 1022 -1397
rect 1023 -1403 1026 -1397
rect 1030 -1403 1033 -1397
rect 1037 -1403 1040 -1397
rect 1044 -1403 1047 -1397
rect 1051 -1403 1054 -1397
rect 1058 -1403 1061 -1397
rect 1065 -1403 1068 -1397
rect 1072 -1403 1075 -1397
rect 1079 -1403 1082 -1397
rect 1086 -1403 1089 -1397
rect 1093 -1403 1096 -1397
rect 1100 -1403 1103 -1397
rect 1107 -1403 1110 -1397
rect 1114 -1403 1117 -1397
rect 1121 -1403 1124 -1397
rect 1128 -1403 1131 -1397
rect 1135 -1403 1138 -1397
rect 1142 -1403 1145 -1397
rect 1149 -1403 1152 -1397
rect 1156 -1403 1159 -1397
rect 1163 -1403 1166 -1397
rect 1170 -1403 1173 -1397
rect 1177 -1403 1180 -1397
rect 1184 -1403 1187 -1397
rect 1191 -1403 1194 -1397
rect 1198 -1403 1201 -1397
rect 1205 -1403 1208 -1397
rect 1212 -1403 1215 -1397
rect 1219 -1403 1222 -1397
rect 1226 -1403 1229 -1397
rect 1233 -1403 1236 -1397
rect 1240 -1403 1243 -1397
rect 1247 -1403 1250 -1397
rect 1254 -1403 1257 -1397
rect 1261 -1403 1264 -1397
rect 1268 -1403 1271 -1397
rect 1275 -1403 1278 -1397
rect 1282 -1403 1285 -1397
rect 1289 -1403 1292 -1397
rect 1296 -1403 1299 -1397
rect 1303 -1403 1306 -1397
rect 1310 -1403 1313 -1397
rect 1317 -1403 1320 -1397
rect 1324 -1403 1327 -1397
rect 1331 -1403 1334 -1397
rect 1338 -1403 1341 -1397
rect 1345 -1403 1348 -1397
rect 1352 -1403 1355 -1397
rect 1359 -1403 1362 -1397
rect 1366 -1403 1369 -1397
rect 1373 -1403 1376 -1397
rect 1380 -1403 1383 -1397
rect 1387 -1403 1390 -1397
rect 1394 -1403 1397 -1397
rect 1401 -1403 1404 -1397
rect 1408 -1403 1411 -1397
rect 1415 -1403 1418 -1397
rect 1422 -1403 1425 -1397
rect 1429 -1403 1432 -1397
rect 1436 -1403 1439 -1397
rect 1443 -1403 1446 -1397
rect 1450 -1403 1453 -1397
rect 1457 -1403 1460 -1397
rect 1464 -1403 1467 -1397
rect 1471 -1403 1474 -1397
rect 1478 -1403 1481 -1397
rect 1485 -1403 1488 -1397
rect 1492 -1403 1495 -1397
rect 1499 -1403 1502 -1397
rect 1506 -1403 1509 -1397
rect 1513 -1403 1516 -1397
rect 1520 -1403 1526 -1397
rect 1527 -1403 1530 -1397
rect 1534 -1403 1537 -1397
rect 1 -1536 4 -1530
rect 8 -1536 11 -1530
rect 15 -1536 18 -1530
rect 22 -1536 25 -1530
rect 29 -1536 32 -1530
rect 36 -1536 39 -1530
rect 43 -1536 46 -1530
rect 50 -1536 56 -1530
rect 57 -1536 60 -1530
rect 64 -1536 67 -1530
rect 71 -1536 74 -1530
rect 78 -1536 84 -1530
rect 85 -1536 88 -1530
rect 92 -1536 95 -1530
rect 99 -1536 105 -1530
rect 106 -1536 109 -1530
rect 113 -1536 116 -1530
rect 120 -1536 123 -1530
rect 127 -1536 130 -1530
rect 134 -1536 137 -1530
rect 141 -1536 144 -1530
rect 148 -1536 151 -1530
rect 155 -1536 158 -1530
rect 162 -1536 165 -1530
rect 169 -1536 175 -1530
rect 176 -1536 179 -1530
rect 183 -1536 186 -1530
rect 190 -1536 193 -1530
rect 197 -1536 200 -1530
rect 204 -1536 207 -1530
rect 211 -1536 214 -1530
rect 218 -1536 221 -1530
rect 225 -1536 228 -1530
rect 232 -1536 235 -1530
rect 239 -1536 242 -1530
rect 246 -1536 249 -1530
rect 253 -1536 256 -1530
rect 260 -1536 263 -1530
rect 267 -1536 270 -1530
rect 274 -1536 277 -1530
rect 281 -1536 284 -1530
rect 288 -1536 291 -1530
rect 295 -1536 298 -1530
rect 302 -1536 305 -1530
rect 309 -1536 312 -1530
rect 316 -1536 319 -1530
rect 323 -1536 326 -1530
rect 330 -1536 333 -1530
rect 337 -1536 340 -1530
rect 344 -1536 347 -1530
rect 351 -1536 354 -1530
rect 358 -1536 361 -1530
rect 365 -1536 368 -1530
rect 372 -1536 375 -1530
rect 379 -1536 382 -1530
rect 386 -1536 389 -1530
rect 393 -1536 399 -1530
rect 400 -1536 403 -1530
rect 407 -1536 410 -1530
rect 414 -1536 417 -1530
rect 421 -1536 424 -1530
rect 428 -1536 434 -1530
rect 435 -1536 438 -1530
rect 442 -1536 445 -1530
rect 449 -1536 452 -1530
rect 456 -1536 459 -1530
rect 463 -1536 466 -1530
rect 470 -1536 476 -1530
rect 477 -1536 480 -1530
rect 484 -1536 487 -1530
rect 491 -1536 494 -1530
rect 498 -1536 504 -1530
rect 505 -1536 508 -1530
rect 512 -1536 515 -1530
rect 519 -1536 522 -1530
rect 526 -1536 529 -1530
rect 533 -1536 536 -1530
rect 540 -1536 543 -1530
rect 547 -1536 550 -1530
rect 554 -1536 557 -1530
rect 561 -1536 564 -1530
rect 568 -1536 571 -1530
rect 575 -1536 581 -1530
rect 582 -1536 585 -1530
rect 589 -1536 592 -1530
rect 596 -1536 602 -1530
rect 603 -1536 606 -1530
rect 610 -1536 613 -1530
rect 617 -1536 620 -1530
rect 624 -1536 627 -1530
rect 631 -1536 634 -1530
rect 638 -1536 641 -1530
rect 645 -1536 648 -1530
rect 652 -1536 655 -1530
rect 659 -1536 662 -1530
rect 666 -1536 669 -1530
rect 673 -1536 679 -1530
rect 680 -1536 686 -1530
rect 687 -1536 690 -1530
rect 694 -1536 697 -1530
rect 701 -1536 704 -1530
rect 708 -1536 711 -1530
rect 715 -1536 718 -1530
rect 722 -1536 728 -1530
rect 729 -1536 732 -1530
rect 736 -1536 739 -1530
rect 743 -1536 746 -1530
rect 750 -1536 753 -1530
rect 757 -1536 760 -1530
rect 764 -1536 770 -1530
rect 771 -1536 774 -1530
rect 778 -1536 781 -1530
rect 785 -1536 788 -1530
rect 792 -1536 795 -1530
rect 799 -1536 805 -1530
rect 806 -1536 809 -1530
rect 813 -1536 819 -1530
rect 820 -1536 823 -1530
rect 827 -1536 833 -1530
rect 834 -1536 840 -1530
rect 841 -1536 844 -1530
rect 848 -1536 851 -1530
rect 855 -1536 861 -1530
rect 862 -1536 865 -1530
rect 869 -1536 872 -1530
rect 876 -1536 882 -1530
rect 883 -1536 886 -1530
rect 890 -1536 893 -1530
rect 897 -1536 900 -1530
rect 904 -1536 907 -1530
rect 911 -1536 914 -1530
rect 918 -1536 921 -1530
rect 925 -1536 928 -1530
rect 932 -1536 935 -1530
rect 939 -1536 942 -1530
rect 946 -1536 949 -1530
rect 953 -1536 956 -1530
rect 960 -1536 963 -1530
rect 967 -1536 970 -1530
rect 974 -1536 977 -1530
rect 981 -1536 984 -1530
rect 988 -1536 994 -1530
rect 995 -1536 1001 -1530
rect 1002 -1536 1005 -1530
rect 1009 -1536 1012 -1530
rect 1016 -1536 1019 -1530
rect 1023 -1536 1026 -1530
rect 1030 -1536 1033 -1530
rect 1037 -1536 1040 -1530
rect 1044 -1536 1047 -1530
rect 1051 -1536 1054 -1530
rect 1058 -1536 1061 -1530
rect 1065 -1536 1068 -1530
rect 1072 -1536 1078 -1530
rect 1079 -1536 1082 -1530
rect 1086 -1536 1089 -1530
rect 1093 -1536 1096 -1530
rect 1100 -1536 1103 -1530
rect 1107 -1536 1110 -1530
rect 1114 -1536 1117 -1530
rect 1121 -1536 1127 -1530
rect 1128 -1536 1131 -1530
rect 1135 -1536 1138 -1530
rect 1142 -1536 1145 -1530
rect 1149 -1536 1152 -1530
rect 1156 -1536 1159 -1530
rect 1163 -1536 1166 -1530
rect 1170 -1536 1173 -1530
rect 1177 -1536 1180 -1530
rect 1184 -1536 1187 -1530
rect 1191 -1536 1194 -1530
rect 1198 -1536 1201 -1530
rect 1205 -1536 1208 -1530
rect 1212 -1536 1215 -1530
rect 1219 -1536 1222 -1530
rect 1226 -1536 1229 -1530
rect 1233 -1536 1236 -1530
rect 1240 -1536 1243 -1530
rect 1247 -1536 1250 -1530
rect 1254 -1536 1257 -1530
rect 1261 -1536 1264 -1530
rect 1268 -1536 1271 -1530
rect 1275 -1536 1278 -1530
rect 1282 -1536 1285 -1530
rect 1289 -1536 1292 -1530
rect 1296 -1536 1299 -1530
rect 1303 -1536 1306 -1530
rect 1310 -1536 1313 -1530
rect 1317 -1536 1320 -1530
rect 1324 -1536 1327 -1530
rect 1331 -1536 1334 -1530
rect 1338 -1536 1341 -1530
rect 1345 -1536 1348 -1530
rect 1352 -1536 1355 -1530
rect 1359 -1536 1362 -1530
rect 1366 -1536 1369 -1530
rect 1373 -1536 1376 -1530
rect 1380 -1536 1383 -1530
rect 1387 -1536 1390 -1530
rect 1394 -1536 1397 -1530
rect 1401 -1536 1404 -1530
rect 1408 -1536 1411 -1530
rect 1415 -1536 1418 -1530
rect 1422 -1536 1425 -1530
rect 1429 -1536 1432 -1530
rect 1436 -1536 1439 -1530
rect 1443 -1536 1446 -1530
rect 1450 -1536 1453 -1530
rect 1457 -1536 1460 -1530
rect 1464 -1536 1467 -1530
rect 1471 -1536 1474 -1530
rect 1478 -1536 1481 -1530
rect 1485 -1536 1488 -1530
rect 1492 -1536 1495 -1530
rect 1499 -1536 1502 -1530
rect 1506 -1536 1509 -1530
rect 1513 -1536 1516 -1530
rect 1520 -1536 1526 -1530
rect 1527 -1536 1530 -1530
rect 1534 -1536 1537 -1530
rect 1 -1643 4 -1637
rect 8 -1643 11 -1637
rect 15 -1643 18 -1637
rect 22 -1643 25 -1637
rect 29 -1643 32 -1637
rect 36 -1643 39 -1637
rect 43 -1643 46 -1637
rect 50 -1643 53 -1637
rect 57 -1643 60 -1637
rect 64 -1643 67 -1637
rect 71 -1643 77 -1637
rect 78 -1643 81 -1637
rect 85 -1643 88 -1637
rect 92 -1643 95 -1637
rect 99 -1643 102 -1637
rect 106 -1643 112 -1637
rect 113 -1643 116 -1637
rect 120 -1643 123 -1637
rect 127 -1643 133 -1637
rect 134 -1643 137 -1637
rect 141 -1643 147 -1637
rect 148 -1643 151 -1637
rect 155 -1643 158 -1637
rect 162 -1643 165 -1637
rect 169 -1643 172 -1637
rect 176 -1643 179 -1637
rect 183 -1643 186 -1637
rect 190 -1643 193 -1637
rect 197 -1643 200 -1637
rect 204 -1643 207 -1637
rect 211 -1643 214 -1637
rect 218 -1643 221 -1637
rect 225 -1643 228 -1637
rect 232 -1643 235 -1637
rect 239 -1643 242 -1637
rect 246 -1643 249 -1637
rect 253 -1643 256 -1637
rect 260 -1643 263 -1637
rect 267 -1643 273 -1637
rect 274 -1643 277 -1637
rect 281 -1643 284 -1637
rect 288 -1643 291 -1637
rect 295 -1643 298 -1637
rect 302 -1643 305 -1637
rect 309 -1643 312 -1637
rect 316 -1643 319 -1637
rect 323 -1643 326 -1637
rect 330 -1643 333 -1637
rect 337 -1643 340 -1637
rect 344 -1643 350 -1637
rect 351 -1643 354 -1637
rect 358 -1643 361 -1637
rect 365 -1643 371 -1637
rect 372 -1643 375 -1637
rect 379 -1643 382 -1637
rect 386 -1643 389 -1637
rect 393 -1643 396 -1637
rect 400 -1643 403 -1637
rect 407 -1643 410 -1637
rect 414 -1643 417 -1637
rect 421 -1643 424 -1637
rect 428 -1643 431 -1637
rect 435 -1643 441 -1637
rect 442 -1643 448 -1637
rect 449 -1643 452 -1637
rect 456 -1643 459 -1637
rect 463 -1643 466 -1637
rect 470 -1643 476 -1637
rect 477 -1643 480 -1637
rect 484 -1643 487 -1637
rect 491 -1643 494 -1637
rect 498 -1643 504 -1637
rect 505 -1643 508 -1637
rect 512 -1643 515 -1637
rect 519 -1643 522 -1637
rect 526 -1643 529 -1637
rect 533 -1643 536 -1637
rect 540 -1643 543 -1637
rect 547 -1643 550 -1637
rect 554 -1643 560 -1637
rect 561 -1643 567 -1637
rect 568 -1643 571 -1637
rect 575 -1643 578 -1637
rect 582 -1643 585 -1637
rect 589 -1643 592 -1637
rect 596 -1643 599 -1637
rect 603 -1643 606 -1637
rect 610 -1643 613 -1637
rect 617 -1643 623 -1637
rect 624 -1643 627 -1637
rect 631 -1643 634 -1637
rect 638 -1643 641 -1637
rect 645 -1643 651 -1637
rect 652 -1643 655 -1637
rect 659 -1643 662 -1637
rect 666 -1643 669 -1637
rect 673 -1643 676 -1637
rect 680 -1643 683 -1637
rect 687 -1643 690 -1637
rect 694 -1643 697 -1637
rect 701 -1643 704 -1637
rect 708 -1643 711 -1637
rect 715 -1643 718 -1637
rect 722 -1643 725 -1637
rect 729 -1643 732 -1637
rect 736 -1643 742 -1637
rect 743 -1643 746 -1637
rect 750 -1643 756 -1637
rect 757 -1643 760 -1637
rect 764 -1643 767 -1637
rect 771 -1643 774 -1637
rect 778 -1643 784 -1637
rect 785 -1643 788 -1637
rect 792 -1643 795 -1637
rect 799 -1643 802 -1637
rect 806 -1643 809 -1637
rect 813 -1643 819 -1637
rect 820 -1643 823 -1637
rect 827 -1643 833 -1637
rect 834 -1643 837 -1637
rect 841 -1643 844 -1637
rect 848 -1643 851 -1637
rect 855 -1643 858 -1637
rect 862 -1643 865 -1637
rect 869 -1643 872 -1637
rect 876 -1643 882 -1637
rect 883 -1643 886 -1637
rect 890 -1643 893 -1637
rect 897 -1643 900 -1637
rect 904 -1643 907 -1637
rect 911 -1643 914 -1637
rect 918 -1643 921 -1637
rect 925 -1643 928 -1637
rect 932 -1643 935 -1637
rect 939 -1643 942 -1637
rect 946 -1643 949 -1637
rect 953 -1643 959 -1637
rect 960 -1643 963 -1637
rect 967 -1643 970 -1637
rect 974 -1643 977 -1637
rect 981 -1643 984 -1637
rect 988 -1643 994 -1637
rect 995 -1643 998 -1637
rect 1002 -1643 1005 -1637
rect 1009 -1643 1012 -1637
rect 1016 -1643 1019 -1637
rect 1023 -1643 1026 -1637
rect 1030 -1643 1033 -1637
rect 1037 -1643 1040 -1637
rect 1044 -1643 1047 -1637
rect 1051 -1643 1054 -1637
rect 1058 -1643 1061 -1637
rect 1065 -1643 1068 -1637
rect 1072 -1643 1075 -1637
rect 1079 -1643 1082 -1637
rect 1086 -1643 1089 -1637
rect 1093 -1643 1096 -1637
rect 1100 -1643 1103 -1637
rect 1107 -1643 1110 -1637
rect 1114 -1643 1117 -1637
rect 1121 -1643 1124 -1637
rect 1128 -1643 1131 -1637
rect 1135 -1643 1138 -1637
rect 1142 -1643 1145 -1637
rect 1149 -1643 1152 -1637
rect 1156 -1643 1159 -1637
rect 1163 -1643 1166 -1637
rect 1170 -1643 1173 -1637
rect 1177 -1643 1180 -1637
rect 1184 -1643 1187 -1637
rect 1191 -1643 1194 -1637
rect 1198 -1643 1201 -1637
rect 1205 -1643 1208 -1637
rect 1212 -1643 1215 -1637
rect 1219 -1643 1222 -1637
rect 1226 -1643 1229 -1637
rect 1233 -1643 1236 -1637
rect 1240 -1643 1243 -1637
rect 1247 -1643 1250 -1637
rect 1254 -1643 1257 -1637
rect 1261 -1643 1264 -1637
rect 1268 -1643 1271 -1637
rect 1275 -1643 1278 -1637
rect 1282 -1643 1285 -1637
rect 1289 -1643 1292 -1637
rect 1296 -1643 1299 -1637
rect 1303 -1643 1306 -1637
rect 1310 -1643 1313 -1637
rect 1317 -1643 1320 -1637
rect 1324 -1643 1327 -1637
rect 1331 -1643 1334 -1637
rect 1338 -1643 1341 -1637
rect 1345 -1643 1351 -1637
rect 1352 -1643 1355 -1637
rect 1359 -1643 1362 -1637
rect 1366 -1643 1369 -1637
rect 1373 -1643 1376 -1637
rect 1380 -1643 1383 -1637
rect 1387 -1643 1390 -1637
rect 1394 -1643 1400 -1637
rect 1401 -1643 1404 -1637
rect 1408 -1643 1411 -1637
rect 1415 -1643 1418 -1637
rect 1422 -1643 1425 -1637
rect 1429 -1643 1432 -1637
rect 1436 -1643 1439 -1637
rect 1450 -1643 1453 -1637
rect 8 -1768 11 -1762
rect 15 -1768 18 -1762
rect 22 -1768 25 -1762
rect 29 -1768 32 -1762
rect 36 -1768 39 -1762
rect 43 -1768 46 -1762
rect 50 -1768 53 -1762
rect 57 -1768 60 -1762
rect 64 -1768 67 -1762
rect 71 -1768 77 -1762
rect 78 -1768 84 -1762
rect 85 -1768 88 -1762
rect 92 -1768 95 -1762
rect 99 -1768 102 -1762
rect 106 -1768 112 -1762
rect 113 -1768 116 -1762
rect 120 -1768 123 -1762
rect 127 -1768 130 -1762
rect 134 -1768 137 -1762
rect 141 -1768 144 -1762
rect 148 -1768 151 -1762
rect 155 -1768 158 -1762
rect 162 -1768 165 -1762
rect 169 -1768 172 -1762
rect 176 -1768 179 -1762
rect 183 -1768 186 -1762
rect 190 -1768 193 -1762
rect 197 -1768 200 -1762
rect 204 -1768 207 -1762
rect 211 -1768 214 -1762
rect 218 -1768 221 -1762
rect 225 -1768 228 -1762
rect 232 -1768 235 -1762
rect 239 -1768 242 -1762
rect 246 -1768 249 -1762
rect 253 -1768 256 -1762
rect 260 -1768 263 -1762
rect 267 -1768 270 -1762
rect 274 -1768 277 -1762
rect 281 -1768 284 -1762
rect 288 -1768 291 -1762
rect 295 -1768 298 -1762
rect 302 -1768 305 -1762
rect 309 -1768 312 -1762
rect 316 -1768 319 -1762
rect 323 -1768 326 -1762
rect 330 -1768 333 -1762
rect 337 -1768 343 -1762
rect 344 -1768 347 -1762
rect 351 -1768 354 -1762
rect 358 -1768 361 -1762
rect 365 -1768 371 -1762
rect 372 -1768 375 -1762
rect 379 -1768 382 -1762
rect 386 -1768 389 -1762
rect 393 -1768 396 -1762
rect 400 -1768 403 -1762
rect 407 -1768 410 -1762
rect 414 -1768 420 -1762
rect 421 -1768 427 -1762
rect 428 -1768 431 -1762
rect 435 -1768 438 -1762
rect 442 -1768 445 -1762
rect 449 -1768 452 -1762
rect 456 -1768 459 -1762
rect 463 -1768 466 -1762
rect 470 -1768 473 -1762
rect 477 -1768 480 -1762
rect 484 -1768 490 -1762
rect 491 -1768 494 -1762
rect 498 -1768 501 -1762
rect 505 -1768 511 -1762
rect 512 -1768 515 -1762
rect 519 -1768 525 -1762
rect 526 -1768 532 -1762
rect 533 -1768 536 -1762
rect 540 -1768 543 -1762
rect 547 -1768 550 -1762
rect 554 -1768 557 -1762
rect 561 -1768 564 -1762
rect 568 -1768 571 -1762
rect 575 -1768 578 -1762
rect 582 -1768 588 -1762
rect 589 -1768 592 -1762
rect 596 -1768 599 -1762
rect 603 -1768 606 -1762
rect 610 -1768 613 -1762
rect 617 -1768 620 -1762
rect 624 -1768 627 -1762
rect 631 -1768 637 -1762
rect 638 -1768 641 -1762
rect 645 -1768 648 -1762
rect 652 -1768 655 -1762
rect 659 -1768 662 -1762
rect 666 -1768 669 -1762
rect 673 -1768 676 -1762
rect 680 -1768 683 -1762
rect 687 -1768 690 -1762
rect 694 -1768 697 -1762
rect 701 -1768 704 -1762
rect 708 -1768 711 -1762
rect 715 -1768 721 -1762
rect 722 -1768 725 -1762
rect 729 -1768 732 -1762
rect 736 -1768 739 -1762
rect 743 -1768 746 -1762
rect 750 -1768 753 -1762
rect 757 -1768 760 -1762
rect 764 -1768 767 -1762
rect 771 -1768 777 -1762
rect 778 -1768 781 -1762
rect 785 -1768 788 -1762
rect 792 -1768 798 -1762
rect 799 -1768 802 -1762
rect 806 -1768 812 -1762
rect 813 -1768 816 -1762
rect 820 -1768 823 -1762
rect 827 -1768 830 -1762
rect 834 -1768 837 -1762
rect 841 -1768 847 -1762
rect 848 -1768 851 -1762
rect 855 -1768 858 -1762
rect 862 -1768 865 -1762
rect 869 -1768 875 -1762
rect 876 -1768 882 -1762
rect 883 -1768 886 -1762
rect 890 -1768 893 -1762
rect 897 -1768 903 -1762
rect 904 -1768 907 -1762
rect 911 -1768 914 -1762
rect 918 -1768 921 -1762
rect 925 -1768 928 -1762
rect 932 -1768 935 -1762
rect 939 -1768 942 -1762
rect 946 -1768 949 -1762
rect 953 -1768 956 -1762
rect 960 -1768 963 -1762
rect 967 -1768 970 -1762
rect 974 -1768 977 -1762
rect 981 -1768 984 -1762
rect 988 -1768 994 -1762
rect 995 -1768 998 -1762
rect 1002 -1768 1008 -1762
rect 1009 -1768 1012 -1762
rect 1016 -1768 1019 -1762
rect 1023 -1768 1026 -1762
rect 1030 -1768 1033 -1762
rect 1037 -1768 1040 -1762
rect 1044 -1768 1047 -1762
rect 1051 -1768 1054 -1762
rect 1058 -1768 1061 -1762
rect 1065 -1768 1068 -1762
rect 1072 -1768 1075 -1762
rect 1079 -1768 1082 -1762
rect 1086 -1768 1089 -1762
rect 1093 -1768 1096 -1762
rect 1100 -1768 1103 -1762
rect 1107 -1768 1110 -1762
rect 1114 -1768 1117 -1762
rect 1121 -1768 1124 -1762
rect 1128 -1768 1131 -1762
rect 1135 -1768 1138 -1762
rect 1142 -1768 1145 -1762
rect 1149 -1768 1152 -1762
rect 1156 -1768 1159 -1762
rect 1163 -1768 1166 -1762
rect 1170 -1768 1173 -1762
rect 1177 -1768 1180 -1762
rect 1184 -1768 1187 -1762
rect 1191 -1768 1194 -1762
rect 1198 -1768 1201 -1762
rect 1205 -1768 1208 -1762
rect 1212 -1768 1215 -1762
rect 1219 -1768 1222 -1762
rect 1226 -1768 1229 -1762
rect 1233 -1768 1236 -1762
rect 1240 -1768 1243 -1762
rect 1247 -1768 1250 -1762
rect 1254 -1768 1257 -1762
rect 1261 -1768 1264 -1762
rect 1268 -1768 1271 -1762
rect 1275 -1768 1278 -1762
rect 1282 -1768 1285 -1762
rect 1289 -1768 1292 -1762
rect 1296 -1768 1299 -1762
rect 1303 -1768 1306 -1762
rect 1310 -1768 1313 -1762
rect 1317 -1768 1320 -1762
rect 1324 -1768 1327 -1762
rect 1331 -1768 1334 -1762
rect 1338 -1768 1341 -1762
rect 1345 -1768 1348 -1762
rect 1352 -1768 1355 -1762
rect 1359 -1768 1362 -1762
rect 1366 -1768 1372 -1762
rect 1373 -1768 1379 -1762
rect 1380 -1768 1383 -1762
rect 1387 -1768 1390 -1762
rect 1394 -1768 1397 -1762
rect 1401 -1768 1404 -1762
rect 1408 -1768 1411 -1762
rect 1415 -1768 1418 -1762
rect 1422 -1768 1425 -1762
rect 1 -1865 4 -1859
rect 8 -1865 11 -1859
rect 15 -1865 21 -1859
rect 22 -1865 25 -1859
rect 29 -1865 32 -1859
rect 36 -1865 39 -1859
rect 43 -1865 46 -1859
rect 50 -1865 53 -1859
rect 57 -1865 63 -1859
rect 64 -1865 67 -1859
rect 71 -1865 74 -1859
rect 78 -1865 81 -1859
rect 85 -1865 91 -1859
rect 92 -1865 95 -1859
rect 99 -1865 102 -1859
rect 106 -1865 109 -1859
rect 113 -1865 116 -1859
rect 120 -1865 123 -1859
rect 127 -1865 130 -1859
rect 134 -1865 140 -1859
rect 141 -1865 144 -1859
rect 148 -1865 151 -1859
rect 155 -1865 158 -1859
rect 162 -1865 165 -1859
rect 169 -1865 172 -1859
rect 176 -1865 179 -1859
rect 183 -1865 186 -1859
rect 190 -1865 193 -1859
rect 197 -1865 200 -1859
rect 204 -1865 207 -1859
rect 211 -1865 214 -1859
rect 218 -1865 221 -1859
rect 225 -1865 228 -1859
rect 232 -1865 235 -1859
rect 239 -1865 242 -1859
rect 246 -1865 249 -1859
rect 253 -1865 256 -1859
rect 260 -1865 263 -1859
rect 267 -1865 270 -1859
rect 274 -1865 277 -1859
rect 281 -1865 284 -1859
rect 288 -1865 291 -1859
rect 295 -1865 301 -1859
rect 302 -1865 305 -1859
rect 309 -1865 312 -1859
rect 316 -1865 319 -1859
rect 323 -1865 326 -1859
rect 330 -1865 333 -1859
rect 337 -1865 340 -1859
rect 344 -1865 350 -1859
rect 351 -1865 354 -1859
rect 358 -1865 361 -1859
rect 365 -1865 368 -1859
rect 372 -1865 375 -1859
rect 379 -1865 382 -1859
rect 386 -1865 389 -1859
rect 393 -1865 399 -1859
rect 400 -1865 403 -1859
rect 407 -1865 410 -1859
rect 414 -1865 417 -1859
rect 421 -1865 424 -1859
rect 428 -1865 434 -1859
rect 435 -1865 438 -1859
rect 442 -1865 445 -1859
rect 449 -1865 452 -1859
rect 456 -1865 459 -1859
rect 463 -1865 466 -1859
rect 470 -1865 473 -1859
rect 477 -1865 480 -1859
rect 484 -1865 487 -1859
rect 491 -1865 494 -1859
rect 498 -1865 504 -1859
rect 505 -1865 508 -1859
rect 512 -1865 515 -1859
rect 519 -1865 522 -1859
rect 526 -1865 529 -1859
rect 533 -1865 536 -1859
rect 540 -1865 543 -1859
rect 547 -1865 550 -1859
rect 554 -1865 560 -1859
rect 561 -1865 564 -1859
rect 568 -1865 574 -1859
rect 575 -1865 578 -1859
rect 582 -1865 585 -1859
rect 589 -1865 595 -1859
rect 596 -1865 599 -1859
rect 603 -1865 606 -1859
rect 610 -1865 613 -1859
rect 617 -1865 620 -1859
rect 624 -1865 627 -1859
rect 631 -1865 634 -1859
rect 638 -1865 641 -1859
rect 645 -1865 648 -1859
rect 652 -1865 655 -1859
rect 659 -1865 665 -1859
rect 666 -1865 669 -1859
rect 673 -1865 676 -1859
rect 680 -1865 686 -1859
rect 687 -1865 693 -1859
rect 694 -1865 697 -1859
rect 701 -1865 704 -1859
rect 708 -1865 711 -1859
rect 715 -1865 721 -1859
rect 722 -1865 725 -1859
rect 729 -1865 732 -1859
rect 736 -1865 739 -1859
rect 743 -1865 746 -1859
rect 750 -1865 756 -1859
rect 757 -1865 760 -1859
rect 764 -1865 767 -1859
rect 771 -1865 777 -1859
rect 778 -1865 781 -1859
rect 785 -1865 788 -1859
rect 792 -1865 795 -1859
rect 799 -1865 805 -1859
rect 806 -1865 809 -1859
rect 813 -1865 816 -1859
rect 820 -1865 823 -1859
rect 827 -1865 830 -1859
rect 834 -1865 837 -1859
rect 841 -1865 844 -1859
rect 848 -1865 851 -1859
rect 855 -1865 858 -1859
rect 862 -1865 865 -1859
rect 869 -1865 872 -1859
rect 876 -1865 879 -1859
rect 883 -1865 889 -1859
rect 890 -1865 893 -1859
rect 897 -1865 900 -1859
rect 904 -1865 910 -1859
rect 911 -1865 914 -1859
rect 918 -1865 921 -1859
rect 925 -1865 928 -1859
rect 932 -1865 938 -1859
rect 939 -1865 942 -1859
rect 946 -1865 949 -1859
rect 953 -1865 956 -1859
rect 960 -1865 963 -1859
rect 967 -1865 970 -1859
rect 974 -1865 977 -1859
rect 981 -1865 984 -1859
rect 988 -1865 991 -1859
rect 995 -1865 998 -1859
rect 1002 -1865 1005 -1859
rect 1009 -1865 1012 -1859
rect 1016 -1865 1019 -1859
rect 1023 -1865 1026 -1859
rect 1030 -1865 1033 -1859
rect 1037 -1865 1040 -1859
rect 1044 -1865 1047 -1859
rect 1051 -1865 1054 -1859
rect 1058 -1865 1064 -1859
rect 1065 -1865 1071 -1859
rect 1072 -1865 1075 -1859
rect 1079 -1865 1082 -1859
rect 1086 -1865 1089 -1859
rect 1093 -1865 1096 -1859
rect 1100 -1865 1103 -1859
rect 1107 -1865 1110 -1859
rect 1114 -1865 1117 -1859
rect 1121 -1865 1124 -1859
rect 1128 -1865 1131 -1859
rect 1135 -1865 1138 -1859
rect 1142 -1865 1145 -1859
rect 1149 -1865 1152 -1859
rect 1156 -1865 1159 -1859
rect 1163 -1865 1166 -1859
rect 1170 -1865 1173 -1859
rect 1177 -1865 1180 -1859
rect 1184 -1865 1187 -1859
rect 1191 -1865 1194 -1859
rect 1198 -1865 1201 -1859
rect 1205 -1865 1208 -1859
rect 1212 -1865 1215 -1859
rect 1219 -1865 1222 -1859
rect 1226 -1865 1229 -1859
rect 1233 -1865 1236 -1859
rect 1240 -1865 1243 -1859
rect 1247 -1865 1250 -1859
rect 1254 -1865 1257 -1859
rect 1261 -1865 1264 -1859
rect 1268 -1865 1271 -1859
rect 1275 -1865 1278 -1859
rect 1282 -1865 1285 -1859
rect 1289 -1865 1292 -1859
rect 1296 -1865 1299 -1859
rect 1303 -1865 1306 -1859
rect 1310 -1865 1313 -1859
rect 1317 -1865 1320 -1859
rect 1324 -1865 1327 -1859
rect 1331 -1865 1334 -1859
rect 1338 -1865 1341 -1859
rect 1345 -1865 1348 -1859
rect 1352 -1865 1355 -1859
rect 1359 -1865 1362 -1859
rect 1366 -1865 1369 -1859
rect 1373 -1865 1376 -1859
rect 1380 -1865 1383 -1859
rect 1387 -1865 1390 -1859
rect 1394 -1865 1400 -1859
rect 1401 -1865 1404 -1859
rect 1408 -1865 1411 -1859
rect 1415 -1865 1418 -1859
rect 1422 -1865 1425 -1859
rect 1429 -1865 1432 -1859
rect 1 -1992 4 -1986
rect 8 -1992 11 -1986
rect 15 -1992 18 -1986
rect 22 -1992 28 -1986
rect 29 -1992 32 -1986
rect 36 -1992 42 -1986
rect 43 -1992 46 -1986
rect 50 -1992 53 -1986
rect 57 -1992 60 -1986
rect 64 -1992 70 -1986
rect 71 -1992 77 -1986
rect 78 -1992 81 -1986
rect 85 -1992 88 -1986
rect 92 -1992 95 -1986
rect 99 -1992 102 -1986
rect 106 -1992 109 -1986
rect 113 -1992 116 -1986
rect 120 -1992 123 -1986
rect 127 -1992 130 -1986
rect 134 -1992 137 -1986
rect 141 -1992 144 -1986
rect 148 -1992 151 -1986
rect 155 -1992 158 -1986
rect 162 -1992 165 -1986
rect 169 -1992 175 -1986
rect 176 -1992 179 -1986
rect 183 -1992 186 -1986
rect 190 -1992 193 -1986
rect 197 -1992 200 -1986
rect 204 -1992 207 -1986
rect 211 -1992 214 -1986
rect 218 -1992 221 -1986
rect 225 -1992 231 -1986
rect 232 -1992 235 -1986
rect 239 -1992 242 -1986
rect 246 -1992 249 -1986
rect 253 -1992 256 -1986
rect 260 -1992 263 -1986
rect 267 -1992 270 -1986
rect 274 -1992 277 -1986
rect 281 -1992 284 -1986
rect 288 -1992 291 -1986
rect 295 -1992 298 -1986
rect 302 -1992 305 -1986
rect 309 -1992 312 -1986
rect 316 -1992 319 -1986
rect 323 -1992 326 -1986
rect 330 -1992 333 -1986
rect 337 -1992 340 -1986
rect 344 -1992 347 -1986
rect 351 -1992 357 -1986
rect 358 -1992 361 -1986
rect 365 -1992 368 -1986
rect 372 -1992 378 -1986
rect 379 -1992 382 -1986
rect 386 -1992 389 -1986
rect 393 -1992 396 -1986
rect 400 -1992 403 -1986
rect 407 -1992 413 -1986
rect 414 -1992 417 -1986
rect 421 -1992 424 -1986
rect 428 -1992 431 -1986
rect 435 -1992 438 -1986
rect 442 -1992 445 -1986
rect 449 -1992 452 -1986
rect 456 -1992 459 -1986
rect 463 -1992 466 -1986
rect 470 -1992 473 -1986
rect 477 -1992 480 -1986
rect 484 -1992 487 -1986
rect 491 -1992 494 -1986
rect 498 -1992 501 -1986
rect 505 -1992 511 -1986
rect 512 -1992 518 -1986
rect 519 -1992 525 -1986
rect 526 -1992 529 -1986
rect 533 -1992 536 -1986
rect 540 -1992 543 -1986
rect 547 -1992 550 -1986
rect 554 -1992 557 -1986
rect 561 -1992 567 -1986
rect 568 -1992 571 -1986
rect 575 -1992 581 -1986
rect 582 -1992 588 -1986
rect 589 -1992 592 -1986
rect 596 -1992 599 -1986
rect 603 -1992 606 -1986
rect 610 -1992 616 -1986
rect 617 -1992 620 -1986
rect 624 -1992 627 -1986
rect 631 -1992 634 -1986
rect 638 -1992 644 -1986
rect 645 -1992 648 -1986
rect 652 -1992 655 -1986
rect 659 -1992 665 -1986
rect 666 -1992 669 -1986
rect 673 -1992 676 -1986
rect 680 -1992 683 -1986
rect 687 -1992 690 -1986
rect 694 -1992 697 -1986
rect 701 -1992 707 -1986
rect 708 -1992 711 -1986
rect 715 -1992 718 -1986
rect 722 -1992 728 -1986
rect 729 -1992 732 -1986
rect 736 -1992 739 -1986
rect 743 -1992 746 -1986
rect 750 -1992 756 -1986
rect 757 -1992 760 -1986
rect 764 -1992 767 -1986
rect 771 -1992 774 -1986
rect 778 -1992 784 -1986
rect 785 -1992 788 -1986
rect 792 -1992 795 -1986
rect 799 -1992 802 -1986
rect 806 -1992 812 -1986
rect 813 -1992 816 -1986
rect 820 -1992 823 -1986
rect 827 -1992 830 -1986
rect 834 -1992 837 -1986
rect 841 -1992 844 -1986
rect 848 -1992 854 -1986
rect 855 -1992 858 -1986
rect 862 -1992 865 -1986
rect 869 -1992 872 -1986
rect 876 -1992 879 -1986
rect 883 -1992 886 -1986
rect 890 -1992 893 -1986
rect 897 -1992 900 -1986
rect 904 -1992 907 -1986
rect 911 -1992 914 -1986
rect 918 -1992 921 -1986
rect 925 -1992 928 -1986
rect 932 -1992 935 -1986
rect 939 -1992 942 -1986
rect 946 -1992 952 -1986
rect 953 -1992 956 -1986
rect 960 -1992 963 -1986
rect 967 -1992 970 -1986
rect 974 -1992 977 -1986
rect 981 -1992 984 -1986
rect 988 -1992 991 -1986
rect 995 -1992 998 -1986
rect 1002 -1992 1005 -1986
rect 1009 -1992 1012 -1986
rect 1016 -1992 1019 -1986
rect 1023 -1992 1026 -1986
rect 1030 -1992 1033 -1986
rect 1037 -1992 1040 -1986
rect 1044 -1992 1047 -1986
rect 1051 -1992 1054 -1986
rect 1058 -1992 1061 -1986
rect 1065 -1992 1068 -1986
rect 1072 -1992 1075 -1986
rect 1079 -1992 1082 -1986
rect 1086 -1992 1089 -1986
rect 1093 -1992 1096 -1986
rect 1100 -1992 1103 -1986
rect 1107 -1992 1110 -1986
rect 1114 -1992 1117 -1986
rect 1121 -1992 1124 -1986
rect 1128 -1992 1131 -1986
rect 1135 -1992 1138 -1986
rect 1142 -1992 1145 -1986
rect 1149 -1992 1152 -1986
rect 1156 -1992 1159 -1986
rect 1163 -1992 1166 -1986
rect 1170 -1992 1173 -1986
rect 1177 -1992 1180 -1986
rect 1184 -1992 1187 -1986
rect 1191 -1992 1194 -1986
rect 1198 -1992 1201 -1986
rect 1205 -1992 1208 -1986
rect 1212 -1992 1215 -1986
rect 1219 -1992 1222 -1986
rect 1226 -1992 1229 -1986
rect 1233 -1992 1236 -1986
rect 1240 -1992 1243 -1986
rect 1247 -1992 1250 -1986
rect 1254 -1992 1257 -1986
rect 1261 -1992 1264 -1986
rect 1268 -1992 1271 -1986
rect 1275 -1992 1278 -1986
rect 1282 -1992 1285 -1986
rect 1289 -1992 1292 -1986
rect 1296 -1992 1299 -1986
rect 1303 -1992 1306 -1986
rect 1310 -1992 1313 -1986
rect 1317 -1992 1320 -1986
rect 1324 -1992 1327 -1986
rect 1331 -1992 1334 -1986
rect 1338 -1992 1341 -1986
rect 1345 -1992 1348 -1986
rect 1352 -1992 1355 -1986
rect 1359 -1992 1362 -1986
rect 1366 -1992 1369 -1986
rect 1373 -1992 1376 -1986
rect 1380 -1992 1383 -1986
rect 1387 -1992 1390 -1986
rect 1394 -1992 1397 -1986
rect 1401 -1992 1404 -1986
rect 1 -2111 7 -2105
rect 8 -2111 14 -2105
rect 15 -2111 18 -2105
rect 22 -2111 25 -2105
rect 29 -2111 32 -2105
rect 36 -2111 39 -2105
rect 43 -2111 46 -2105
rect 50 -2111 53 -2105
rect 57 -2111 60 -2105
rect 64 -2111 67 -2105
rect 71 -2111 74 -2105
rect 78 -2111 81 -2105
rect 85 -2111 88 -2105
rect 92 -2111 98 -2105
rect 99 -2111 102 -2105
rect 106 -2111 112 -2105
rect 113 -2111 116 -2105
rect 120 -2111 123 -2105
rect 127 -2111 133 -2105
rect 134 -2111 137 -2105
rect 141 -2111 144 -2105
rect 148 -2111 151 -2105
rect 155 -2111 158 -2105
rect 162 -2111 168 -2105
rect 169 -2111 175 -2105
rect 176 -2111 179 -2105
rect 183 -2111 186 -2105
rect 190 -2111 193 -2105
rect 197 -2111 200 -2105
rect 204 -2111 207 -2105
rect 211 -2111 214 -2105
rect 218 -2111 221 -2105
rect 225 -2111 228 -2105
rect 232 -2111 235 -2105
rect 239 -2111 242 -2105
rect 246 -2111 249 -2105
rect 253 -2111 256 -2105
rect 260 -2111 263 -2105
rect 267 -2111 270 -2105
rect 274 -2111 277 -2105
rect 281 -2111 284 -2105
rect 288 -2111 291 -2105
rect 295 -2111 298 -2105
rect 302 -2111 305 -2105
rect 309 -2111 312 -2105
rect 316 -2111 322 -2105
rect 323 -2111 326 -2105
rect 330 -2111 336 -2105
rect 337 -2111 340 -2105
rect 344 -2111 350 -2105
rect 351 -2111 354 -2105
rect 358 -2111 361 -2105
rect 365 -2111 368 -2105
rect 372 -2111 375 -2105
rect 379 -2111 382 -2105
rect 386 -2111 389 -2105
rect 393 -2111 396 -2105
rect 400 -2111 403 -2105
rect 407 -2111 410 -2105
rect 414 -2111 417 -2105
rect 421 -2111 424 -2105
rect 428 -2111 431 -2105
rect 435 -2111 438 -2105
rect 442 -2111 445 -2105
rect 449 -2111 455 -2105
rect 456 -2111 459 -2105
rect 463 -2111 466 -2105
rect 470 -2111 473 -2105
rect 477 -2111 480 -2105
rect 484 -2111 490 -2105
rect 491 -2111 494 -2105
rect 498 -2111 504 -2105
rect 505 -2111 508 -2105
rect 512 -2111 515 -2105
rect 519 -2111 522 -2105
rect 526 -2111 529 -2105
rect 533 -2111 536 -2105
rect 540 -2111 543 -2105
rect 547 -2111 550 -2105
rect 554 -2111 557 -2105
rect 561 -2111 564 -2105
rect 568 -2111 571 -2105
rect 575 -2111 581 -2105
rect 582 -2111 585 -2105
rect 589 -2111 592 -2105
rect 596 -2111 599 -2105
rect 603 -2111 606 -2105
rect 610 -2111 613 -2105
rect 617 -2111 623 -2105
rect 624 -2111 627 -2105
rect 631 -2111 634 -2105
rect 638 -2111 641 -2105
rect 645 -2111 648 -2105
rect 652 -2111 655 -2105
rect 659 -2111 662 -2105
rect 666 -2111 672 -2105
rect 673 -2111 676 -2105
rect 680 -2111 683 -2105
rect 687 -2111 693 -2105
rect 694 -2111 697 -2105
rect 701 -2111 704 -2105
rect 708 -2111 711 -2105
rect 715 -2111 718 -2105
rect 722 -2111 725 -2105
rect 729 -2111 732 -2105
rect 736 -2111 739 -2105
rect 743 -2111 746 -2105
rect 750 -2111 753 -2105
rect 757 -2111 760 -2105
rect 764 -2111 767 -2105
rect 771 -2111 774 -2105
rect 778 -2111 784 -2105
rect 785 -2111 788 -2105
rect 792 -2111 795 -2105
rect 799 -2111 802 -2105
rect 806 -2111 809 -2105
rect 813 -2111 819 -2105
rect 820 -2111 826 -2105
rect 827 -2111 830 -2105
rect 834 -2111 837 -2105
rect 841 -2111 844 -2105
rect 848 -2111 851 -2105
rect 855 -2111 858 -2105
rect 862 -2111 865 -2105
rect 869 -2111 872 -2105
rect 876 -2111 879 -2105
rect 883 -2111 886 -2105
rect 890 -2111 896 -2105
rect 897 -2111 900 -2105
rect 904 -2111 907 -2105
rect 911 -2111 914 -2105
rect 918 -2111 921 -2105
rect 925 -2111 928 -2105
rect 932 -2111 935 -2105
rect 939 -2111 942 -2105
rect 946 -2111 949 -2105
rect 953 -2111 956 -2105
rect 960 -2111 963 -2105
rect 967 -2111 973 -2105
rect 974 -2111 977 -2105
rect 981 -2111 984 -2105
rect 988 -2111 994 -2105
rect 995 -2111 998 -2105
rect 1002 -2111 1005 -2105
rect 1009 -2111 1012 -2105
rect 1016 -2111 1019 -2105
rect 1023 -2111 1026 -2105
rect 1030 -2111 1033 -2105
rect 1037 -2111 1040 -2105
rect 1044 -2111 1047 -2105
rect 1051 -2111 1054 -2105
rect 1058 -2111 1061 -2105
rect 1065 -2111 1068 -2105
rect 1072 -2111 1075 -2105
rect 1079 -2111 1082 -2105
rect 1086 -2111 1089 -2105
rect 1093 -2111 1096 -2105
rect 1100 -2111 1103 -2105
rect 1107 -2111 1110 -2105
rect 1114 -2111 1120 -2105
rect 1121 -2111 1124 -2105
rect 1128 -2111 1131 -2105
rect 1135 -2111 1141 -2105
rect 1142 -2111 1145 -2105
rect 1149 -2111 1152 -2105
rect 1156 -2111 1159 -2105
rect 1163 -2111 1166 -2105
rect 1170 -2111 1173 -2105
rect 1177 -2111 1180 -2105
rect 1184 -2111 1187 -2105
rect 1191 -2111 1194 -2105
rect 1198 -2111 1201 -2105
rect 1205 -2111 1208 -2105
rect 1212 -2111 1215 -2105
rect 1219 -2111 1222 -2105
rect 1226 -2111 1229 -2105
rect 1233 -2111 1236 -2105
rect 1240 -2111 1243 -2105
rect 1247 -2111 1250 -2105
rect 1254 -2111 1257 -2105
rect 1261 -2111 1264 -2105
rect 1268 -2111 1271 -2105
rect 1275 -2111 1278 -2105
rect 1282 -2111 1285 -2105
rect 1289 -2111 1292 -2105
rect 1296 -2111 1299 -2105
rect 1303 -2111 1306 -2105
rect 1310 -2111 1313 -2105
rect 1317 -2111 1320 -2105
rect 1324 -2111 1327 -2105
rect 1 -2244 4 -2238
rect 8 -2244 11 -2238
rect 15 -2244 18 -2238
rect 22 -2244 28 -2238
rect 29 -2244 35 -2238
rect 36 -2244 42 -2238
rect 43 -2244 46 -2238
rect 50 -2244 53 -2238
rect 57 -2244 60 -2238
rect 64 -2244 67 -2238
rect 71 -2244 77 -2238
rect 78 -2244 81 -2238
rect 85 -2244 88 -2238
rect 92 -2244 95 -2238
rect 99 -2244 102 -2238
rect 106 -2244 109 -2238
rect 113 -2244 119 -2238
rect 120 -2244 123 -2238
rect 127 -2244 130 -2238
rect 134 -2244 140 -2238
rect 141 -2244 144 -2238
rect 148 -2244 154 -2238
rect 155 -2244 158 -2238
rect 162 -2244 165 -2238
rect 169 -2244 172 -2238
rect 176 -2244 179 -2238
rect 183 -2244 186 -2238
rect 190 -2244 193 -2238
rect 197 -2244 200 -2238
rect 204 -2244 207 -2238
rect 211 -2244 214 -2238
rect 218 -2244 221 -2238
rect 225 -2244 228 -2238
rect 232 -2244 235 -2238
rect 239 -2244 242 -2238
rect 246 -2244 249 -2238
rect 253 -2244 256 -2238
rect 260 -2244 263 -2238
rect 267 -2244 270 -2238
rect 274 -2244 277 -2238
rect 281 -2244 284 -2238
rect 288 -2244 291 -2238
rect 295 -2244 301 -2238
rect 302 -2244 305 -2238
rect 309 -2244 312 -2238
rect 316 -2244 319 -2238
rect 323 -2244 326 -2238
rect 330 -2244 333 -2238
rect 337 -2244 343 -2238
rect 344 -2244 347 -2238
rect 351 -2244 354 -2238
rect 358 -2244 361 -2238
rect 365 -2244 368 -2238
rect 372 -2244 375 -2238
rect 379 -2244 382 -2238
rect 386 -2244 389 -2238
rect 393 -2244 399 -2238
rect 400 -2244 406 -2238
rect 407 -2244 413 -2238
rect 414 -2244 417 -2238
rect 421 -2244 427 -2238
rect 428 -2244 431 -2238
rect 435 -2244 438 -2238
rect 442 -2244 445 -2238
rect 449 -2244 455 -2238
rect 456 -2244 459 -2238
rect 463 -2244 466 -2238
rect 470 -2244 473 -2238
rect 477 -2244 480 -2238
rect 484 -2244 487 -2238
rect 491 -2244 494 -2238
rect 498 -2244 501 -2238
rect 505 -2244 508 -2238
rect 512 -2244 515 -2238
rect 519 -2244 525 -2238
rect 526 -2244 532 -2238
rect 533 -2244 536 -2238
rect 540 -2244 543 -2238
rect 547 -2244 550 -2238
rect 554 -2244 560 -2238
rect 561 -2244 564 -2238
rect 568 -2244 571 -2238
rect 575 -2244 578 -2238
rect 582 -2244 585 -2238
rect 589 -2244 592 -2238
rect 596 -2244 599 -2238
rect 603 -2244 606 -2238
rect 610 -2244 613 -2238
rect 617 -2244 623 -2238
rect 624 -2244 630 -2238
rect 631 -2244 634 -2238
rect 638 -2244 641 -2238
rect 645 -2244 651 -2238
rect 652 -2244 655 -2238
rect 659 -2244 662 -2238
rect 666 -2244 669 -2238
rect 673 -2244 679 -2238
rect 680 -2244 683 -2238
rect 687 -2244 690 -2238
rect 694 -2244 697 -2238
rect 701 -2244 704 -2238
rect 708 -2244 711 -2238
rect 715 -2244 718 -2238
rect 722 -2244 725 -2238
rect 729 -2244 732 -2238
rect 736 -2244 739 -2238
rect 743 -2244 746 -2238
rect 750 -2244 753 -2238
rect 757 -2244 760 -2238
rect 764 -2244 767 -2238
rect 771 -2244 774 -2238
rect 778 -2244 781 -2238
rect 785 -2244 788 -2238
rect 792 -2244 795 -2238
rect 799 -2244 802 -2238
rect 806 -2244 812 -2238
rect 813 -2244 816 -2238
rect 820 -2244 823 -2238
rect 827 -2244 830 -2238
rect 834 -2244 837 -2238
rect 841 -2244 844 -2238
rect 848 -2244 851 -2238
rect 855 -2244 858 -2238
rect 862 -2244 865 -2238
rect 869 -2244 875 -2238
rect 876 -2244 879 -2238
rect 883 -2244 886 -2238
rect 890 -2244 893 -2238
rect 897 -2244 900 -2238
rect 904 -2244 907 -2238
rect 911 -2244 914 -2238
rect 918 -2244 921 -2238
rect 925 -2244 928 -2238
rect 932 -2244 938 -2238
rect 939 -2244 942 -2238
rect 946 -2244 949 -2238
rect 953 -2244 956 -2238
rect 960 -2244 963 -2238
rect 967 -2244 970 -2238
rect 974 -2244 977 -2238
rect 981 -2244 987 -2238
rect 988 -2244 991 -2238
rect 995 -2244 998 -2238
rect 1002 -2244 1005 -2238
rect 1009 -2244 1012 -2238
rect 1016 -2244 1019 -2238
rect 1023 -2244 1026 -2238
rect 1030 -2244 1033 -2238
rect 1037 -2244 1040 -2238
rect 1044 -2244 1047 -2238
rect 1051 -2244 1054 -2238
rect 1058 -2244 1061 -2238
rect 1065 -2244 1068 -2238
rect 1072 -2244 1075 -2238
rect 1079 -2244 1082 -2238
rect 1086 -2244 1089 -2238
rect 1093 -2244 1096 -2238
rect 1100 -2244 1103 -2238
rect 1107 -2244 1110 -2238
rect 1114 -2244 1117 -2238
rect 1121 -2244 1124 -2238
rect 1128 -2244 1131 -2238
rect 1135 -2244 1138 -2238
rect 1142 -2244 1145 -2238
rect 1149 -2244 1152 -2238
rect 1156 -2244 1159 -2238
rect 1163 -2244 1166 -2238
rect 1170 -2244 1173 -2238
rect 1177 -2244 1180 -2238
rect 1184 -2244 1187 -2238
rect 1191 -2244 1194 -2238
rect 1198 -2244 1201 -2238
rect 1205 -2244 1208 -2238
rect 1212 -2244 1215 -2238
rect 1219 -2244 1222 -2238
rect 1226 -2244 1229 -2238
rect 1233 -2244 1236 -2238
rect 1240 -2244 1243 -2238
rect 1247 -2244 1250 -2238
rect 1254 -2244 1257 -2238
rect 1261 -2244 1264 -2238
rect 1268 -2244 1271 -2238
rect 1275 -2244 1278 -2238
rect 1282 -2244 1285 -2238
rect 1289 -2244 1292 -2238
rect 1296 -2244 1299 -2238
rect 1303 -2244 1306 -2238
rect 1310 -2244 1313 -2238
rect 1 -2369 7 -2363
rect 8 -2369 11 -2363
rect 15 -2369 18 -2363
rect 22 -2369 25 -2363
rect 29 -2369 32 -2363
rect 36 -2369 42 -2363
rect 43 -2369 46 -2363
rect 50 -2369 56 -2363
rect 57 -2369 63 -2363
rect 64 -2369 67 -2363
rect 71 -2369 74 -2363
rect 78 -2369 81 -2363
rect 85 -2369 88 -2363
rect 92 -2369 98 -2363
rect 99 -2369 102 -2363
rect 106 -2369 109 -2363
rect 113 -2369 116 -2363
rect 120 -2369 123 -2363
rect 127 -2369 130 -2363
rect 134 -2369 140 -2363
rect 141 -2369 144 -2363
rect 148 -2369 154 -2363
rect 155 -2369 158 -2363
rect 162 -2369 165 -2363
rect 169 -2369 172 -2363
rect 176 -2369 179 -2363
rect 183 -2369 186 -2363
rect 190 -2369 193 -2363
rect 197 -2369 200 -2363
rect 204 -2369 207 -2363
rect 211 -2369 214 -2363
rect 218 -2369 221 -2363
rect 225 -2369 228 -2363
rect 232 -2369 235 -2363
rect 239 -2369 242 -2363
rect 246 -2369 249 -2363
rect 253 -2369 256 -2363
rect 260 -2369 263 -2363
rect 267 -2369 270 -2363
rect 274 -2369 277 -2363
rect 281 -2369 284 -2363
rect 288 -2369 291 -2363
rect 295 -2369 298 -2363
rect 302 -2369 308 -2363
rect 309 -2369 312 -2363
rect 316 -2369 322 -2363
rect 323 -2369 326 -2363
rect 330 -2369 333 -2363
rect 337 -2369 343 -2363
rect 344 -2369 347 -2363
rect 351 -2369 354 -2363
rect 358 -2369 361 -2363
rect 365 -2369 368 -2363
rect 372 -2369 375 -2363
rect 379 -2369 382 -2363
rect 386 -2369 389 -2363
rect 393 -2369 399 -2363
rect 400 -2369 403 -2363
rect 407 -2369 410 -2363
rect 414 -2369 417 -2363
rect 421 -2369 427 -2363
rect 428 -2369 431 -2363
rect 435 -2369 441 -2363
rect 442 -2369 445 -2363
rect 449 -2369 452 -2363
rect 456 -2369 459 -2363
rect 463 -2369 466 -2363
rect 470 -2369 473 -2363
rect 477 -2369 480 -2363
rect 484 -2369 487 -2363
rect 491 -2369 494 -2363
rect 498 -2369 501 -2363
rect 505 -2369 508 -2363
rect 512 -2369 518 -2363
rect 519 -2369 522 -2363
rect 526 -2369 529 -2363
rect 533 -2369 536 -2363
rect 540 -2369 543 -2363
rect 547 -2369 550 -2363
rect 554 -2369 560 -2363
rect 561 -2369 564 -2363
rect 568 -2369 571 -2363
rect 575 -2369 581 -2363
rect 582 -2369 585 -2363
rect 589 -2369 595 -2363
rect 596 -2369 599 -2363
rect 603 -2369 606 -2363
rect 610 -2369 613 -2363
rect 617 -2369 620 -2363
rect 624 -2369 627 -2363
rect 631 -2369 637 -2363
rect 638 -2369 641 -2363
rect 645 -2369 648 -2363
rect 652 -2369 655 -2363
rect 659 -2369 665 -2363
rect 666 -2369 669 -2363
rect 673 -2369 676 -2363
rect 680 -2369 683 -2363
rect 687 -2369 690 -2363
rect 694 -2369 697 -2363
rect 701 -2369 704 -2363
rect 708 -2369 711 -2363
rect 715 -2369 718 -2363
rect 722 -2369 728 -2363
rect 729 -2369 732 -2363
rect 736 -2369 739 -2363
rect 743 -2369 749 -2363
rect 750 -2369 753 -2363
rect 757 -2369 763 -2363
rect 764 -2369 767 -2363
rect 771 -2369 774 -2363
rect 778 -2369 781 -2363
rect 785 -2369 788 -2363
rect 792 -2369 795 -2363
rect 799 -2369 802 -2363
rect 806 -2369 812 -2363
rect 813 -2369 816 -2363
rect 820 -2369 823 -2363
rect 827 -2369 830 -2363
rect 834 -2369 837 -2363
rect 841 -2369 844 -2363
rect 848 -2369 854 -2363
rect 855 -2369 858 -2363
rect 862 -2369 865 -2363
rect 869 -2369 872 -2363
rect 876 -2369 879 -2363
rect 883 -2369 886 -2363
rect 890 -2369 893 -2363
rect 897 -2369 900 -2363
rect 904 -2369 907 -2363
rect 911 -2369 914 -2363
rect 918 -2369 921 -2363
rect 925 -2369 928 -2363
rect 932 -2369 935 -2363
rect 939 -2369 942 -2363
rect 946 -2369 949 -2363
rect 953 -2369 956 -2363
rect 960 -2369 963 -2363
rect 967 -2369 970 -2363
rect 974 -2369 977 -2363
rect 981 -2369 984 -2363
rect 988 -2369 991 -2363
rect 995 -2369 998 -2363
rect 1002 -2369 1005 -2363
rect 1009 -2369 1012 -2363
rect 1016 -2369 1019 -2363
rect 1023 -2369 1026 -2363
rect 1030 -2369 1036 -2363
rect 1037 -2369 1040 -2363
rect 1044 -2369 1047 -2363
rect 1051 -2369 1054 -2363
rect 1058 -2369 1061 -2363
rect 1065 -2369 1068 -2363
rect 1072 -2369 1075 -2363
rect 1079 -2369 1082 -2363
rect 1086 -2369 1089 -2363
rect 1093 -2369 1096 -2363
rect 1100 -2369 1103 -2363
rect 1107 -2369 1110 -2363
rect 1114 -2369 1117 -2363
rect 1121 -2369 1124 -2363
rect 1128 -2369 1131 -2363
rect 1135 -2369 1138 -2363
rect 1142 -2369 1145 -2363
rect 1149 -2369 1152 -2363
rect 1156 -2369 1159 -2363
rect 1163 -2369 1166 -2363
rect 1170 -2369 1173 -2363
rect 1177 -2369 1180 -2363
rect 1184 -2369 1187 -2363
rect 1191 -2369 1194 -2363
rect 1198 -2369 1201 -2363
rect 1205 -2369 1208 -2363
rect 1212 -2369 1215 -2363
rect 1219 -2369 1222 -2363
rect 1226 -2369 1229 -2363
rect 1233 -2369 1236 -2363
rect 1240 -2369 1243 -2363
rect 1247 -2369 1250 -2363
rect 57 -2466 60 -2460
rect 64 -2466 67 -2460
rect 71 -2466 74 -2460
rect 78 -2466 81 -2460
rect 85 -2466 88 -2460
rect 92 -2466 95 -2460
rect 99 -2466 102 -2460
rect 106 -2466 109 -2460
rect 113 -2466 116 -2460
rect 120 -2466 126 -2460
rect 127 -2466 133 -2460
rect 134 -2466 137 -2460
rect 141 -2466 144 -2460
rect 148 -2466 151 -2460
rect 155 -2466 158 -2460
rect 162 -2466 168 -2460
rect 169 -2466 175 -2460
rect 176 -2466 179 -2460
rect 183 -2466 186 -2460
rect 190 -2466 193 -2460
rect 197 -2466 203 -2460
rect 204 -2466 207 -2460
rect 211 -2466 214 -2460
rect 218 -2466 221 -2460
rect 225 -2466 228 -2460
rect 232 -2466 235 -2460
rect 239 -2466 242 -2460
rect 246 -2466 249 -2460
rect 253 -2466 256 -2460
rect 260 -2466 263 -2460
rect 267 -2466 270 -2460
rect 274 -2466 277 -2460
rect 281 -2466 284 -2460
rect 288 -2466 291 -2460
rect 295 -2466 298 -2460
rect 302 -2466 305 -2460
rect 309 -2466 312 -2460
rect 316 -2466 319 -2460
rect 323 -2466 326 -2460
rect 330 -2466 333 -2460
rect 337 -2466 340 -2460
rect 344 -2466 347 -2460
rect 351 -2466 357 -2460
rect 358 -2466 361 -2460
rect 365 -2466 368 -2460
rect 372 -2466 378 -2460
rect 379 -2466 382 -2460
rect 386 -2466 389 -2460
rect 393 -2466 396 -2460
rect 400 -2466 403 -2460
rect 407 -2466 410 -2460
rect 414 -2466 417 -2460
rect 421 -2466 424 -2460
rect 428 -2466 431 -2460
rect 435 -2466 441 -2460
rect 442 -2466 448 -2460
rect 449 -2466 452 -2460
rect 456 -2466 459 -2460
rect 463 -2466 469 -2460
rect 470 -2466 473 -2460
rect 477 -2466 480 -2460
rect 484 -2466 487 -2460
rect 491 -2466 494 -2460
rect 498 -2466 501 -2460
rect 505 -2466 508 -2460
rect 512 -2466 518 -2460
rect 519 -2466 522 -2460
rect 526 -2466 529 -2460
rect 533 -2466 536 -2460
rect 540 -2466 543 -2460
rect 547 -2466 550 -2460
rect 554 -2466 557 -2460
rect 561 -2466 567 -2460
rect 568 -2466 574 -2460
rect 575 -2466 578 -2460
rect 582 -2466 585 -2460
rect 589 -2466 592 -2460
rect 596 -2466 599 -2460
rect 603 -2466 606 -2460
rect 610 -2466 616 -2460
rect 617 -2466 620 -2460
rect 624 -2466 627 -2460
rect 631 -2466 634 -2460
rect 638 -2466 641 -2460
rect 645 -2466 648 -2460
rect 652 -2466 655 -2460
rect 659 -2466 665 -2460
rect 666 -2466 669 -2460
rect 673 -2466 679 -2460
rect 680 -2466 683 -2460
rect 687 -2466 690 -2460
rect 694 -2466 700 -2460
rect 701 -2466 704 -2460
rect 708 -2466 711 -2460
rect 715 -2466 718 -2460
rect 722 -2466 728 -2460
rect 729 -2466 732 -2460
rect 736 -2466 739 -2460
rect 743 -2466 746 -2460
rect 750 -2466 753 -2460
rect 757 -2466 760 -2460
rect 764 -2466 767 -2460
rect 771 -2466 774 -2460
rect 778 -2466 781 -2460
rect 785 -2466 788 -2460
rect 792 -2466 798 -2460
rect 799 -2466 802 -2460
rect 806 -2466 809 -2460
rect 813 -2466 816 -2460
rect 820 -2466 823 -2460
rect 827 -2466 833 -2460
rect 834 -2466 837 -2460
rect 841 -2466 844 -2460
rect 848 -2466 851 -2460
rect 855 -2466 858 -2460
rect 862 -2466 865 -2460
rect 869 -2466 872 -2460
rect 876 -2466 879 -2460
rect 883 -2466 886 -2460
rect 890 -2466 893 -2460
rect 897 -2466 900 -2460
rect 904 -2466 910 -2460
rect 911 -2466 914 -2460
rect 918 -2466 921 -2460
rect 925 -2466 928 -2460
rect 932 -2466 935 -2460
rect 939 -2466 945 -2460
rect 946 -2466 949 -2460
rect 953 -2466 956 -2460
rect 960 -2466 963 -2460
rect 967 -2466 970 -2460
rect 974 -2466 977 -2460
rect 981 -2466 984 -2460
rect 988 -2466 991 -2460
rect 995 -2466 998 -2460
rect 1002 -2466 1005 -2460
rect 1009 -2466 1015 -2460
rect 1016 -2466 1019 -2460
rect 1023 -2466 1026 -2460
rect 1030 -2466 1033 -2460
rect 1058 -2466 1061 -2460
rect 1065 -2466 1068 -2460
rect 1072 -2466 1075 -2460
rect 1079 -2466 1082 -2460
rect 1086 -2466 1089 -2460
rect 1093 -2466 1096 -2460
rect 1100 -2466 1106 -2460
rect 1107 -2466 1110 -2460
rect 1128 -2466 1131 -2460
rect 1191 -2466 1194 -2460
rect 127 -2549 130 -2543
rect 134 -2549 137 -2543
rect 225 -2549 228 -2543
rect 232 -2549 235 -2543
rect 246 -2549 249 -2543
rect 253 -2549 256 -2543
rect 260 -2549 263 -2543
rect 267 -2549 270 -2543
rect 274 -2549 280 -2543
rect 281 -2549 284 -2543
rect 288 -2549 291 -2543
rect 295 -2549 298 -2543
rect 302 -2549 305 -2543
rect 309 -2549 312 -2543
rect 316 -2549 319 -2543
rect 323 -2549 329 -2543
rect 330 -2549 333 -2543
rect 337 -2549 340 -2543
rect 344 -2549 347 -2543
rect 351 -2549 354 -2543
rect 358 -2549 361 -2543
rect 365 -2549 371 -2543
rect 372 -2549 375 -2543
rect 379 -2549 382 -2543
rect 386 -2549 392 -2543
rect 393 -2549 396 -2543
rect 400 -2549 403 -2543
rect 407 -2549 410 -2543
rect 414 -2549 417 -2543
rect 421 -2549 424 -2543
rect 428 -2549 431 -2543
rect 435 -2549 438 -2543
rect 442 -2549 445 -2543
rect 449 -2549 452 -2543
rect 456 -2549 462 -2543
rect 463 -2549 466 -2543
rect 470 -2549 476 -2543
rect 477 -2549 480 -2543
rect 484 -2549 490 -2543
rect 491 -2549 494 -2543
rect 498 -2549 501 -2543
rect 505 -2549 511 -2543
rect 512 -2549 515 -2543
rect 519 -2549 525 -2543
rect 526 -2549 532 -2543
rect 533 -2549 536 -2543
rect 540 -2549 546 -2543
rect 547 -2549 553 -2543
rect 554 -2549 557 -2543
rect 561 -2549 564 -2543
rect 568 -2549 574 -2543
rect 575 -2549 578 -2543
rect 582 -2549 588 -2543
rect 589 -2549 595 -2543
rect 596 -2549 599 -2543
rect 603 -2549 606 -2543
rect 610 -2549 613 -2543
rect 617 -2549 623 -2543
rect 624 -2549 627 -2543
rect 631 -2549 634 -2543
rect 638 -2549 641 -2543
rect 645 -2549 648 -2543
rect 652 -2549 655 -2543
rect 659 -2549 662 -2543
rect 666 -2549 669 -2543
rect 673 -2549 676 -2543
rect 680 -2549 686 -2543
rect 687 -2549 693 -2543
rect 694 -2549 697 -2543
rect 701 -2549 704 -2543
rect 708 -2549 711 -2543
rect 715 -2549 718 -2543
rect 722 -2549 725 -2543
rect 729 -2549 732 -2543
rect 736 -2549 742 -2543
rect 743 -2549 749 -2543
rect 750 -2549 753 -2543
rect 757 -2549 760 -2543
rect 764 -2549 767 -2543
rect 771 -2549 774 -2543
rect 778 -2549 781 -2543
rect 785 -2549 788 -2543
rect 792 -2549 795 -2543
rect 799 -2549 802 -2543
rect 806 -2549 812 -2543
rect 827 -2549 830 -2543
rect 862 -2549 868 -2543
rect 869 -2549 872 -2543
rect 911 -2549 914 -2543
rect 925 -2549 928 -2543
rect 932 -2549 935 -2543
rect 946 -2549 949 -2543
rect 953 -2549 956 -2543
rect 974 -2549 977 -2543
rect 1016 -2549 1019 -2543
rect 1030 -2549 1033 -2543
rect 1037 -2549 1040 -2543
rect 1051 -2549 1054 -2543
rect 1065 -2549 1068 -2543
rect 1093 -2549 1099 -2543
rect 1142 -2549 1145 -2543
rect 1177 -2549 1183 -2543
rect 1184 -2549 1187 -2543
rect 127 -2594 133 -2588
rect 134 -2594 137 -2588
rect 253 -2594 259 -2588
rect 323 -2594 326 -2588
rect 330 -2594 333 -2588
rect 337 -2594 340 -2588
rect 344 -2594 350 -2588
rect 365 -2594 368 -2588
rect 372 -2594 378 -2588
rect 379 -2594 385 -2588
rect 442 -2594 445 -2588
rect 449 -2594 452 -2588
rect 470 -2594 473 -2588
rect 491 -2594 494 -2588
rect 498 -2594 501 -2588
rect 505 -2594 508 -2588
rect 512 -2594 518 -2588
rect 526 -2594 532 -2588
rect 533 -2594 536 -2588
rect 540 -2594 546 -2588
rect 547 -2594 553 -2588
rect 554 -2594 557 -2588
rect 561 -2594 567 -2588
rect 568 -2594 571 -2588
rect 575 -2594 578 -2588
rect 596 -2594 602 -2588
rect 645 -2594 651 -2588
rect 659 -2594 665 -2588
rect 666 -2594 669 -2588
rect 673 -2594 679 -2588
rect 680 -2594 686 -2588
rect 687 -2594 693 -2588
rect 708 -2594 714 -2588
rect 715 -2594 718 -2588
rect 722 -2594 725 -2588
rect 729 -2594 732 -2588
rect 750 -2594 753 -2588
rect 806 -2594 812 -2588
rect 813 -2594 816 -2588
rect 883 -2594 889 -2588
rect 897 -2594 900 -2588
rect 953 -2594 956 -2588
rect 960 -2594 966 -2588
rect 967 -2594 970 -2588
rect 1009 -2594 1015 -2588
rect 1016 -2594 1019 -2588
rect 1023 -2594 1026 -2588
rect 1044 -2594 1047 -2588
rect 1051 -2594 1057 -2588
rect 1058 -2594 1061 -2588
<< polysilicon >>
rect 156 -23 157 -21
rect 215 -17 216 -15
rect 215 -23 216 -21
rect 240 -17 241 -15
rect 240 -23 241 -21
rect 247 -17 248 -15
rect 247 -23 248 -21
rect 261 -17 262 -15
rect 261 -23 262 -21
rect 268 -17 269 -15
rect 275 -17 276 -15
rect 275 -23 276 -21
rect 282 -23 283 -21
rect 285 -23 286 -21
rect 338 -17 339 -15
rect 338 -23 339 -21
rect 373 -17 374 -15
rect 373 -23 374 -21
rect 380 -17 381 -15
rect 380 -23 381 -21
rect 383 -23 384 -21
rect 387 -17 388 -15
rect 387 -23 388 -21
rect 397 -17 398 -15
rect 397 -23 398 -21
rect 401 -17 402 -15
rect 401 -23 402 -21
rect 404 -23 405 -21
rect 408 -17 409 -15
rect 411 -17 412 -15
rect 408 -23 409 -21
rect 415 -17 416 -15
rect 415 -23 416 -21
rect 425 -17 426 -15
rect 425 -23 426 -21
rect 429 -17 430 -15
rect 429 -23 430 -21
rect 457 -17 458 -15
rect 457 -23 458 -21
rect 460 -23 461 -21
rect 464 -17 465 -15
rect 467 -17 468 -15
rect 467 -23 468 -21
rect 478 -17 479 -15
rect 478 -23 479 -21
rect 481 -23 482 -21
rect 485 -17 486 -15
rect 485 -23 486 -21
rect 499 -17 500 -15
rect 499 -23 500 -21
rect 506 -17 507 -15
rect 506 -23 507 -21
rect 516 -17 517 -15
rect 513 -23 514 -21
rect 516 -23 517 -21
rect 527 -17 528 -15
rect 527 -23 528 -21
rect 548 -23 549 -21
rect 551 -23 552 -21
rect 562 -17 563 -15
rect 562 -23 563 -21
rect 569 -17 570 -15
rect 569 -23 570 -21
rect 576 -17 577 -15
rect 576 -23 577 -21
rect 583 -17 584 -15
rect 586 -17 587 -15
rect 583 -23 584 -21
rect 604 -17 605 -15
rect 607 -17 608 -15
rect 607 -23 608 -21
rect 639 -17 640 -15
rect 639 -23 640 -21
rect 667 -17 668 -15
rect 667 -23 668 -21
rect 681 -17 682 -15
rect 681 -23 682 -21
rect 702 -17 703 -15
rect 702 -23 703 -21
rect 709 -17 710 -15
rect 709 -23 710 -21
rect 765 -17 766 -15
rect 765 -23 766 -21
rect 800 -17 801 -15
rect 803 -17 804 -15
rect 800 -23 801 -21
rect 828 -17 829 -15
rect 828 -23 829 -21
rect 149 -66 150 -64
rect 152 -66 153 -64
rect 156 -60 157 -58
rect 159 -66 160 -64
rect 163 -60 164 -58
rect 163 -66 164 -64
rect 191 -60 192 -58
rect 191 -66 192 -64
rect 219 -60 220 -58
rect 219 -66 220 -64
rect 226 -60 227 -58
rect 226 -66 227 -64
rect 233 -60 234 -58
rect 233 -66 234 -64
rect 247 -60 248 -58
rect 247 -66 248 -64
rect 254 -60 255 -58
rect 254 -66 255 -64
rect 261 -60 262 -58
rect 261 -66 262 -64
rect 268 -60 269 -58
rect 268 -66 269 -64
rect 275 -60 276 -58
rect 275 -66 276 -64
rect 282 -60 283 -58
rect 282 -66 283 -64
rect 292 -60 293 -58
rect 289 -66 290 -64
rect 292 -66 293 -64
rect 296 -60 297 -58
rect 296 -66 297 -64
rect 303 -60 304 -58
rect 303 -66 304 -64
rect 310 -60 311 -58
rect 310 -66 311 -64
rect 317 -60 318 -58
rect 317 -66 318 -64
rect 324 -60 325 -58
rect 324 -66 325 -64
rect 331 -60 332 -58
rect 331 -66 332 -64
rect 338 -66 339 -64
rect 341 -66 342 -64
rect 345 -60 346 -58
rect 345 -66 346 -64
rect 348 -66 349 -64
rect 355 -60 356 -58
rect 352 -66 353 -64
rect 355 -66 356 -64
rect 359 -60 360 -58
rect 359 -66 360 -64
rect 366 -60 367 -58
rect 366 -66 367 -64
rect 373 -60 374 -58
rect 373 -66 374 -64
rect 380 -60 381 -58
rect 383 -66 384 -64
rect 387 -60 388 -58
rect 387 -66 388 -64
rect 394 -60 395 -58
rect 394 -66 395 -64
rect 401 -60 402 -58
rect 401 -66 402 -64
rect 411 -60 412 -58
rect 411 -66 412 -64
rect 418 -60 419 -58
rect 415 -66 416 -64
rect 418 -66 419 -64
rect 422 -60 423 -58
rect 422 -66 423 -64
rect 429 -60 430 -58
rect 429 -66 430 -64
rect 436 -60 437 -58
rect 436 -66 437 -64
rect 443 -60 444 -58
rect 443 -66 444 -64
rect 450 -66 451 -64
rect 453 -66 454 -64
rect 457 -60 458 -58
rect 457 -66 458 -64
rect 464 -60 465 -58
rect 464 -66 465 -64
rect 471 -60 472 -58
rect 471 -66 472 -64
rect 478 -60 479 -58
rect 478 -66 479 -64
rect 481 -66 482 -64
rect 485 -60 486 -58
rect 485 -66 486 -64
rect 492 -60 493 -58
rect 492 -66 493 -64
rect 499 -60 500 -58
rect 502 -60 503 -58
rect 499 -66 500 -64
rect 506 -60 507 -58
rect 506 -66 507 -64
rect 513 -60 514 -58
rect 513 -66 514 -64
rect 520 -60 521 -58
rect 520 -66 521 -64
rect 527 -60 528 -58
rect 527 -66 528 -64
rect 534 -60 535 -58
rect 537 -60 538 -58
rect 537 -66 538 -64
rect 541 -60 542 -58
rect 541 -66 542 -64
rect 548 -60 549 -58
rect 548 -66 549 -64
rect 555 -60 556 -58
rect 555 -66 556 -64
rect 558 -66 559 -64
rect 562 -60 563 -58
rect 562 -66 563 -64
rect 569 -60 570 -58
rect 569 -66 570 -64
rect 579 -60 580 -58
rect 576 -66 577 -64
rect 579 -66 580 -64
rect 583 -60 584 -58
rect 583 -66 584 -64
rect 593 -60 594 -58
rect 590 -66 591 -64
rect 593 -66 594 -64
rect 597 -60 598 -58
rect 597 -66 598 -64
rect 604 -60 605 -58
rect 604 -66 605 -64
rect 611 -60 612 -58
rect 611 -66 612 -64
rect 618 -60 619 -58
rect 621 -60 622 -58
rect 618 -66 619 -64
rect 625 -60 626 -58
rect 625 -66 626 -64
rect 632 -60 633 -58
rect 632 -66 633 -64
rect 639 -60 640 -58
rect 639 -66 640 -64
rect 646 -60 647 -58
rect 646 -66 647 -64
rect 653 -60 654 -58
rect 653 -66 654 -64
rect 660 -60 661 -58
rect 660 -66 661 -64
rect 667 -60 668 -58
rect 670 -66 671 -64
rect 674 -60 675 -58
rect 674 -66 675 -64
rect 681 -60 682 -58
rect 681 -66 682 -64
rect 688 -60 689 -58
rect 688 -66 689 -64
rect 702 -60 703 -58
rect 702 -66 703 -64
rect 716 -60 717 -58
rect 719 -60 720 -58
rect 719 -66 720 -64
rect 723 -60 724 -58
rect 723 -66 724 -64
rect 751 -60 752 -58
rect 751 -66 752 -64
rect 758 -60 759 -58
rect 758 -66 759 -64
rect 772 -60 773 -58
rect 772 -66 773 -64
rect 828 -60 829 -58
rect 828 -66 829 -64
rect 849 -60 850 -58
rect 849 -66 850 -64
rect 877 -60 878 -58
rect 877 -66 878 -64
rect 905 -60 906 -58
rect 905 -66 906 -64
rect 23 -121 24 -119
rect 23 -127 24 -125
rect 30 -121 31 -119
rect 30 -127 31 -125
rect 37 -121 38 -119
rect 37 -127 38 -125
rect 44 -121 45 -119
rect 44 -127 45 -125
rect 51 -121 52 -119
rect 51 -127 52 -125
rect 58 -127 59 -125
rect 61 -127 62 -125
rect 65 -121 66 -119
rect 68 -127 69 -125
rect 75 -121 76 -119
rect 75 -127 76 -125
rect 79 -121 80 -119
rect 79 -127 80 -125
rect 86 -121 87 -119
rect 89 -121 90 -119
rect 89 -127 90 -125
rect 93 -121 94 -119
rect 93 -127 94 -125
rect 100 -121 101 -119
rect 100 -127 101 -125
rect 107 -121 108 -119
rect 107 -127 108 -125
rect 114 -121 115 -119
rect 117 -121 118 -119
rect 117 -127 118 -125
rect 121 -121 122 -119
rect 121 -127 122 -125
rect 128 -121 129 -119
rect 131 -127 132 -125
rect 135 -121 136 -119
rect 135 -127 136 -125
rect 142 -121 143 -119
rect 142 -127 143 -125
rect 149 -121 150 -119
rect 149 -127 150 -125
rect 156 -121 157 -119
rect 156 -127 157 -125
rect 163 -121 164 -119
rect 163 -127 164 -125
rect 170 -121 171 -119
rect 170 -127 171 -125
rect 177 -121 178 -119
rect 177 -127 178 -125
rect 184 -121 185 -119
rect 187 -121 188 -119
rect 187 -127 188 -125
rect 194 -121 195 -119
rect 191 -127 192 -125
rect 194 -127 195 -125
rect 198 -121 199 -119
rect 198 -127 199 -125
rect 205 -121 206 -119
rect 205 -127 206 -125
rect 212 -121 213 -119
rect 212 -127 213 -125
rect 219 -121 220 -119
rect 219 -127 220 -125
rect 226 -121 227 -119
rect 226 -127 227 -125
rect 233 -121 234 -119
rect 233 -127 234 -125
rect 240 -121 241 -119
rect 240 -127 241 -125
rect 247 -121 248 -119
rect 247 -127 248 -125
rect 254 -121 255 -119
rect 254 -127 255 -125
rect 261 -121 262 -119
rect 261 -127 262 -125
rect 268 -121 269 -119
rect 271 -121 272 -119
rect 268 -127 269 -125
rect 271 -127 272 -125
rect 275 -121 276 -119
rect 275 -127 276 -125
rect 282 -121 283 -119
rect 282 -127 283 -125
rect 289 -121 290 -119
rect 289 -127 290 -125
rect 299 -121 300 -119
rect 296 -127 297 -125
rect 299 -127 300 -125
rect 303 -121 304 -119
rect 303 -127 304 -125
rect 310 -121 311 -119
rect 313 -121 314 -119
rect 310 -127 311 -125
rect 317 -121 318 -119
rect 317 -127 318 -125
rect 327 -121 328 -119
rect 324 -127 325 -125
rect 327 -127 328 -125
rect 331 -121 332 -119
rect 331 -127 332 -125
rect 338 -121 339 -119
rect 338 -127 339 -125
rect 345 -121 346 -119
rect 345 -127 346 -125
rect 352 -121 353 -119
rect 352 -127 353 -125
rect 359 -121 360 -119
rect 362 -127 363 -125
rect 366 -121 367 -119
rect 366 -127 367 -125
rect 373 -121 374 -119
rect 373 -127 374 -125
rect 380 -121 381 -119
rect 380 -127 381 -125
rect 387 -121 388 -119
rect 387 -127 388 -125
rect 394 -121 395 -119
rect 397 -121 398 -119
rect 397 -127 398 -125
rect 401 -121 402 -119
rect 404 -121 405 -119
rect 401 -127 402 -125
rect 408 -121 409 -119
rect 408 -127 409 -125
rect 415 -121 416 -119
rect 415 -127 416 -125
rect 422 -121 423 -119
rect 422 -127 423 -125
rect 429 -121 430 -119
rect 429 -127 430 -125
rect 436 -121 437 -119
rect 439 -121 440 -119
rect 436 -127 437 -125
rect 439 -127 440 -125
rect 443 -121 444 -119
rect 443 -127 444 -125
rect 450 -121 451 -119
rect 450 -127 451 -125
rect 457 -121 458 -119
rect 457 -127 458 -125
rect 464 -121 465 -119
rect 464 -127 465 -125
rect 471 -121 472 -119
rect 471 -127 472 -125
rect 478 -121 479 -119
rect 478 -127 479 -125
rect 485 -121 486 -119
rect 485 -127 486 -125
rect 492 -121 493 -119
rect 492 -127 493 -125
rect 499 -121 500 -119
rect 499 -127 500 -125
rect 506 -121 507 -119
rect 506 -127 507 -125
rect 513 -121 514 -119
rect 513 -127 514 -125
rect 520 -121 521 -119
rect 520 -127 521 -125
rect 530 -121 531 -119
rect 527 -127 528 -125
rect 530 -127 531 -125
rect 534 -121 535 -119
rect 534 -127 535 -125
rect 541 -121 542 -119
rect 541 -127 542 -125
rect 548 -121 549 -119
rect 548 -127 549 -125
rect 555 -121 556 -119
rect 555 -127 556 -125
rect 562 -121 563 -119
rect 562 -127 563 -125
rect 569 -121 570 -119
rect 569 -127 570 -125
rect 576 -121 577 -119
rect 576 -127 577 -125
rect 583 -121 584 -119
rect 583 -127 584 -125
rect 590 -121 591 -119
rect 590 -127 591 -125
rect 597 -121 598 -119
rect 597 -127 598 -125
rect 604 -121 605 -119
rect 607 -121 608 -119
rect 607 -127 608 -125
rect 611 -121 612 -119
rect 611 -127 612 -125
rect 618 -121 619 -119
rect 618 -127 619 -125
rect 625 -121 626 -119
rect 625 -127 626 -125
rect 632 -121 633 -119
rect 632 -127 633 -125
rect 639 -121 640 -119
rect 639 -127 640 -125
rect 646 -121 647 -119
rect 646 -127 647 -125
rect 653 -121 654 -119
rect 653 -127 654 -125
rect 660 -121 661 -119
rect 663 -121 664 -119
rect 663 -127 664 -125
rect 667 -121 668 -119
rect 667 -127 668 -125
rect 674 -121 675 -119
rect 674 -127 675 -125
rect 681 -121 682 -119
rect 681 -127 682 -125
rect 688 -121 689 -119
rect 688 -127 689 -125
rect 695 -121 696 -119
rect 695 -127 696 -125
rect 702 -121 703 -119
rect 702 -127 703 -125
rect 709 -121 710 -119
rect 709 -127 710 -125
rect 716 -121 717 -119
rect 716 -127 717 -125
rect 723 -121 724 -119
rect 723 -127 724 -125
rect 730 -121 731 -119
rect 730 -127 731 -125
rect 737 -121 738 -119
rect 737 -127 738 -125
rect 744 -121 745 -119
rect 744 -127 745 -125
rect 751 -121 752 -119
rect 751 -127 752 -125
rect 761 -121 762 -119
rect 765 -121 766 -119
rect 765 -127 766 -125
rect 772 -121 773 -119
rect 772 -127 773 -125
rect 779 -121 780 -119
rect 779 -127 780 -125
rect 786 -121 787 -119
rect 786 -127 787 -125
rect 793 -121 794 -119
rect 793 -127 794 -125
rect 800 -121 801 -119
rect 800 -127 801 -125
rect 807 -121 808 -119
rect 807 -127 808 -125
rect 814 -121 815 -119
rect 814 -127 815 -125
rect 821 -121 822 -119
rect 821 -127 822 -125
rect 849 -121 850 -119
rect 849 -127 850 -125
rect 856 -121 857 -119
rect 856 -127 857 -125
rect 870 -121 871 -119
rect 870 -127 871 -125
rect 877 -121 878 -119
rect 877 -127 878 -125
rect 940 -121 941 -119
rect 940 -127 941 -125
rect 947 -121 948 -119
rect 947 -127 948 -125
rect 1500 -121 1501 -119
rect 1500 -127 1501 -125
rect 1507 -121 1508 -119
rect 9 -200 10 -198
rect 9 -206 10 -204
rect 16 -200 17 -198
rect 16 -206 17 -204
rect 23 -200 24 -198
rect 23 -206 24 -204
rect 30 -200 31 -198
rect 30 -206 31 -204
rect 37 -200 38 -198
rect 37 -206 38 -204
rect 44 -200 45 -198
rect 44 -206 45 -204
rect 51 -200 52 -198
rect 54 -200 55 -198
rect 51 -206 52 -204
rect 54 -206 55 -204
rect 58 -200 59 -198
rect 58 -206 59 -204
rect 65 -200 66 -198
rect 65 -206 66 -204
rect 72 -200 73 -198
rect 72 -206 73 -204
rect 79 -200 80 -198
rect 79 -206 80 -204
rect 86 -200 87 -198
rect 86 -206 87 -204
rect 93 -200 94 -198
rect 93 -206 94 -204
rect 100 -200 101 -198
rect 103 -200 104 -198
rect 103 -206 104 -204
rect 107 -200 108 -198
rect 107 -206 108 -204
rect 114 -200 115 -198
rect 114 -206 115 -204
rect 121 -200 122 -198
rect 121 -206 122 -204
rect 128 -200 129 -198
rect 128 -206 129 -204
rect 135 -200 136 -198
rect 135 -206 136 -204
rect 142 -200 143 -198
rect 145 -200 146 -198
rect 142 -206 143 -204
rect 149 -200 150 -198
rect 152 -200 153 -198
rect 149 -206 150 -204
rect 156 -200 157 -198
rect 156 -206 157 -204
rect 159 -206 160 -204
rect 163 -200 164 -198
rect 163 -206 164 -204
rect 170 -200 171 -198
rect 170 -206 171 -204
rect 177 -200 178 -198
rect 177 -206 178 -204
rect 184 -200 185 -198
rect 184 -206 185 -204
rect 191 -200 192 -198
rect 191 -206 192 -204
rect 198 -200 199 -198
rect 198 -206 199 -204
rect 205 -200 206 -198
rect 205 -206 206 -204
rect 212 -200 213 -198
rect 212 -206 213 -204
rect 219 -200 220 -198
rect 219 -206 220 -204
rect 226 -200 227 -198
rect 226 -206 227 -204
rect 233 -200 234 -198
rect 233 -206 234 -204
rect 240 -200 241 -198
rect 240 -206 241 -204
rect 243 -206 244 -204
rect 247 -200 248 -198
rect 247 -206 248 -204
rect 254 -200 255 -198
rect 254 -206 255 -204
rect 261 -200 262 -198
rect 261 -206 262 -204
rect 268 -200 269 -198
rect 271 -200 272 -198
rect 268 -206 269 -204
rect 271 -206 272 -204
rect 275 -200 276 -198
rect 275 -206 276 -204
rect 282 -200 283 -198
rect 282 -206 283 -204
rect 289 -200 290 -198
rect 289 -206 290 -204
rect 296 -200 297 -198
rect 296 -206 297 -204
rect 303 -200 304 -198
rect 306 -200 307 -198
rect 303 -206 304 -204
rect 310 -200 311 -198
rect 310 -206 311 -204
rect 317 -200 318 -198
rect 320 -200 321 -198
rect 317 -206 318 -204
rect 320 -206 321 -204
rect 324 -200 325 -198
rect 324 -206 325 -204
rect 331 -200 332 -198
rect 334 -200 335 -198
rect 334 -206 335 -204
rect 338 -200 339 -198
rect 338 -206 339 -204
rect 345 -200 346 -198
rect 345 -206 346 -204
rect 352 -200 353 -198
rect 352 -206 353 -204
rect 359 -200 360 -198
rect 359 -206 360 -204
rect 366 -200 367 -198
rect 366 -206 367 -204
rect 373 -200 374 -198
rect 373 -206 374 -204
rect 380 -200 381 -198
rect 380 -206 381 -204
rect 387 -200 388 -198
rect 390 -200 391 -198
rect 387 -206 388 -204
rect 390 -206 391 -204
rect 394 -200 395 -198
rect 394 -206 395 -204
rect 401 -200 402 -198
rect 401 -206 402 -204
rect 408 -200 409 -198
rect 408 -206 409 -204
rect 415 -200 416 -198
rect 415 -206 416 -204
rect 422 -200 423 -198
rect 422 -206 423 -204
rect 429 -200 430 -198
rect 429 -206 430 -204
rect 436 -200 437 -198
rect 439 -200 440 -198
rect 436 -206 437 -204
rect 439 -206 440 -204
rect 443 -200 444 -198
rect 443 -206 444 -204
rect 446 -206 447 -204
rect 450 -200 451 -198
rect 450 -206 451 -204
rect 457 -200 458 -198
rect 460 -200 461 -198
rect 457 -206 458 -204
rect 464 -200 465 -198
rect 464 -206 465 -204
rect 471 -200 472 -198
rect 471 -206 472 -204
rect 478 -200 479 -198
rect 478 -206 479 -204
rect 485 -200 486 -198
rect 488 -200 489 -198
rect 485 -206 486 -204
rect 492 -200 493 -198
rect 492 -206 493 -204
rect 499 -200 500 -198
rect 499 -206 500 -204
rect 506 -200 507 -198
rect 506 -206 507 -204
rect 516 -200 517 -198
rect 513 -206 514 -204
rect 516 -206 517 -204
rect 520 -200 521 -198
rect 520 -206 521 -204
rect 527 -200 528 -198
rect 527 -206 528 -204
rect 534 -200 535 -198
rect 537 -200 538 -198
rect 534 -206 535 -204
rect 537 -206 538 -204
rect 541 -200 542 -198
rect 541 -206 542 -204
rect 548 -200 549 -198
rect 548 -206 549 -204
rect 555 -200 556 -198
rect 555 -206 556 -204
rect 562 -200 563 -198
rect 562 -206 563 -204
rect 569 -200 570 -198
rect 569 -206 570 -204
rect 576 -200 577 -198
rect 576 -206 577 -204
rect 583 -200 584 -198
rect 583 -206 584 -204
rect 590 -200 591 -198
rect 590 -206 591 -204
rect 597 -200 598 -198
rect 597 -206 598 -204
rect 604 -200 605 -198
rect 607 -200 608 -198
rect 604 -206 605 -204
rect 607 -206 608 -204
rect 611 -200 612 -198
rect 611 -206 612 -204
rect 618 -200 619 -198
rect 618 -206 619 -204
rect 625 -200 626 -198
rect 625 -206 626 -204
rect 632 -200 633 -198
rect 632 -206 633 -204
rect 639 -200 640 -198
rect 639 -206 640 -204
rect 646 -200 647 -198
rect 646 -206 647 -204
rect 653 -200 654 -198
rect 653 -206 654 -204
rect 660 -200 661 -198
rect 660 -206 661 -204
rect 667 -200 668 -198
rect 667 -206 668 -204
rect 674 -200 675 -198
rect 674 -206 675 -204
rect 681 -200 682 -198
rect 681 -206 682 -204
rect 688 -200 689 -198
rect 688 -206 689 -204
rect 695 -200 696 -198
rect 695 -206 696 -204
rect 702 -200 703 -198
rect 702 -206 703 -204
rect 709 -200 710 -198
rect 709 -206 710 -204
rect 719 -200 720 -198
rect 716 -206 717 -204
rect 719 -206 720 -204
rect 723 -200 724 -198
rect 723 -206 724 -204
rect 730 -200 731 -198
rect 730 -206 731 -204
rect 737 -200 738 -198
rect 737 -206 738 -204
rect 744 -200 745 -198
rect 744 -206 745 -204
rect 751 -200 752 -198
rect 751 -206 752 -204
rect 758 -200 759 -198
rect 758 -206 759 -204
rect 765 -200 766 -198
rect 765 -206 766 -204
rect 772 -200 773 -198
rect 772 -206 773 -204
rect 779 -200 780 -198
rect 779 -206 780 -204
rect 786 -200 787 -198
rect 786 -206 787 -204
rect 793 -200 794 -198
rect 793 -206 794 -204
rect 800 -200 801 -198
rect 800 -206 801 -204
rect 807 -200 808 -198
rect 807 -206 808 -204
rect 814 -200 815 -198
rect 814 -206 815 -204
rect 821 -200 822 -198
rect 821 -206 822 -204
rect 828 -200 829 -198
rect 828 -206 829 -204
rect 835 -200 836 -198
rect 835 -206 836 -204
rect 842 -200 843 -198
rect 842 -206 843 -204
rect 849 -200 850 -198
rect 849 -206 850 -204
rect 856 -200 857 -198
rect 856 -206 857 -204
rect 863 -200 864 -198
rect 863 -206 864 -204
rect 870 -200 871 -198
rect 870 -206 871 -204
rect 877 -200 878 -198
rect 877 -206 878 -204
rect 884 -200 885 -198
rect 884 -206 885 -204
rect 891 -200 892 -198
rect 891 -206 892 -204
rect 898 -200 899 -198
rect 898 -206 899 -204
rect 905 -200 906 -198
rect 905 -206 906 -204
rect 912 -200 913 -198
rect 912 -206 913 -204
rect 919 -200 920 -198
rect 919 -206 920 -204
rect 926 -200 927 -198
rect 926 -206 927 -204
rect 933 -200 934 -198
rect 933 -206 934 -204
rect 940 -200 941 -198
rect 940 -206 941 -204
rect 947 -200 948 -198
rect 947 -206 948 -204
rect 954 -200 955 -198
rect 954 -206 955 -204
rect 961 -200 962 -198
rect 961 -206 962 -204
rect 968 -200 969 -198
rect 968 -206 969 -204
rect 975 -200 976 -198
rect 978 -200 979 -198
rect 975 -206 976 -204
rect 978 -206 979 -204
rect 982 -200 983 -198
rect 985 -200 986 -198
rect 982 -206 983 -204
rect 989 -200 990 -198
rect 992 -206 993 -204
rect 996 -200 997 -198
rect 996 -206 997 -204
rect 1024 -200 1025 -198
rect 1024 -206 1025 -204
rect 1500 -200 1501 -198
rect 1500 -206 1501 -204
rect 2 -311 3 -309
rect 2 -317 3 -315
rect 9 -311 10 -309
rect 9 -317 10 -315
rect 16 -311 17 -309
rect 16 -317 17 -315
rect 26 -311 27 -309
rect 23 -317 24 -315
rect 26 -317 27 -315
rect 30 -311 31 -309
rect 33 -311 34 -309
rect 33 -317 34 -315
rect 37 -311 38 -309
rect 40 -311 41 -309
rect 37 -317 38 -315
rect 44 -311 45 -309
rect 44 -317 45 -315
rect 51 -311 52 -309
rect 54 -311 55 -309
rect 51 -317 52 -315
rect 58 -311 59 -309
rect 58 -317 59 -315
rect 65 -311 66 -309
rect 68 -311 69 -309
rect 68 -317 69 -315
rect 72 -311 73 -309
rect 72 -317 73 -315
rect 82 -311 83 -309
rect 79 -317 80 -315
rect 82 -317 83 -315
rect 86 -311 87 -309
rect 86 -317 87 -315
rect 93 -311 94 -309
rect 96 -311 97 -309
rect 93 -317 94 -315
rect 96 -317 97 -315
rect 100 -311 101 -309
rect 100 -317 101 -315
rect 107 -311 108 -309
rect 107 -317 108 -315
rect 114 -311 115 -309
rect 114 -317 115 -315
rect 121 -311 122 -309
rect 124 -311 125 -309
rect 121 -317 122 -315
rect 124 -317 125 -315
rect 128 -311 129 -309
rect 128 -317 129 -315
rect 135 -311 136 -309
rect 135 -317 136 -315
rect 142 -311 143 -309
rect 142 -317 143 -315
rect 149 -311 150 -309
rect 149 -317 150 -315
rect 156 -311 157 -309
rect 156 -317 157 -315
rect 163 -311 164 -309
rect 163 -317 164 -315
rect 170 -311 171 -309
rect 170 -317 171 -315
rect 177 -311 178 -309
rect 177 -317 178 -315
rect 184 -311 185 -309
rect 184 -317 185 -315
rect 191 -311 192 -309
rect 191 -317 192 -315
rect 198 -311 199 -309
rect 198 -317 199 -315
rect 205 -311 206 -309
rect 205 -317 206 -315
rect 212 -311 213 -309
rect 212 -317 213 -315
rect 219 -311 220 -309
rect 219 -317 220 -315
rect 226 -311 227 -309
rect 226 -317 227 -315
rect 233 -311 234 -309
rect 233 -317 234 -315
rect 240 -311 241 -309
rect 240 -317 241 -315
rect 247 -311 248 -309
rect 247 -317 248 -315
rect 254 -311 255 -309
rect 254 -317 255 -315
rect 261 -311 262 -309
rect 261 -317 262 -315
rect 268 -311 269 -309
rect 268 -317 269 -315
rect 275 -311 276 -309
rect 275 -317 276 -315
rect 282 -311 283 -309
rect 285 -311 286 -309
rect 282 -317 283 -315
rect 285 -317 286 -315
rect 289 -311 290 -309
rect 289 -317 290 -315
rect 296 -311 297 -309
rect 296 -317 297 -315
rect 303 -311 304 -309
rect 303 -317 304 -315
rect 310 -311 311 -309
rect 313 -311 314 -309
rect 313 -317 314 -315
rect 317 -311 318 -309
rect 320 -311 321 -309
rect 317 -317 318 -315
rect 320 -317 321 -315
rect 324 -311 325 -309
rect 327 -311 328 -309
rect 324 -317 325 -315
rect 327 -317 328 -315
rect 331 -311 332 -309
rect 331 -317 332 -315
rect 338 -311 339 -309
rect 338 -317 339 -315
rect 345 -311 346 -309
rect 345 -317 346 -315
rect 352 -311 353 -309
rect 352 -317 353 -315
rect 359 -311 360 -309
rect 362 -311 363 -309
rect 359 -317 360 -315
rect 366 -311 367 -309
rect 366 -317 367 -315
rect 373 -311 374 -309
rect 373 -317 374 -315
rect 380 -311 381 -309
rect 380 -317 381 -315
rect 387 -311 388 -309
rect 387 -317 388 -315
rect 394 -311 395 -309
rect 394 -317 395 -315
rect 401 -311 402 -309
rect 401 -317 402 -315
rect 408 -311 409 -309
rect 408 -317 409 -315
rect 411 -317 412 -315
rect 415 -311 416 -309
rect 415 -317 416 -315
rect 422 -311 423 -309
rect 425 -311 426 -309
rect 422 -317 423 -315
rect 429 -311 430 -309
rect 429 -317 430 -315
rect 436 -311 437 -309
rect 436 -317 437 -315
rect 443 -311 444 -309
rect 443 -317 444 -315
rect 450 -311 451 -309
rect 453 -311 454 -309
rect 450 -317 451 -315
rect 453 -317 454 -315
rect 457 -311 458 -309
rect 457 -317 458 -315
rect 464 -311 465 -309
rect 464 -317 465 -315
rect 471 -311 472 -309
rect 471 -317 472 -315
rect 478 -311 479 -309
rect 478 -317 479 -315
rect 485 -311 486 -309
rect 485 -317 486 -315
rect 492 -311 493 -309
rect 492 -317 493 -315
rect 499 -311 500 -309
rect 499 -317 500 -315
rect 506 -311 507 -309
rect 506 -317 507 -315
rect 513 -311 514 -309
rect 513 -317 514 -315
rect 520 -311 521 -309
rect 520 -317 521 -315
rect 527 -311 528 -309
rect 527 -317 528 -315
rect 534 -311 535 -309
rect 534 -317 535 -315
rect 541 -311 542 -309
rect 544 -311 545 -309
rect 544 -317 545 -315
rect 548 -311 549 -309
rect 548 -317 549 -315
rect 555 -311 556 -309
rect 555 -317 556 -315
rect 562 -311 563 -309
rect 562 -317 563 -315
rect 569 -311 570 -309
rect 569 -317 570 -315
rect 576 -311 577 -309
rect 579 -311 580 -309
rect 576 -317 577 -315
rect 579 -317 580 -315
rect 583 -311 584 -309
rect 583 -317 584 -315
rect 586 -317 587 -315
rect 590 -311 591 -309
rect 590 -317 591 -315
rect 597 -311 598 -309
rect 597 -317 598 -315
rect 604 -311 605 -309
rect 607 -311 608 -309
rect 611 -311 612 -309
rect 611 -317 612 -315
rect 618 -311 619 -309
rect 618 -317 619 -315
rect 625 -311 626 -309
rect 625 -317 626 -315
rect 632 -311 633 -309
rect 632 -317 633 -315
rect 639 -311 640 -309
rect 639 -317 640 -315
rect 646 -311 647 -309
rect 646 -317 647 -315
rect 653 -311 654 -309
rect 653 -317 654 -315
rect 660 -311 661 -309
rect 660 -317 661 -315
rect 667 -311 668 -309
rect 667 -317 668 -315
rect 674 -311 675 -309
rect 674 -317 675 -315
rect 681 -311 682 -309
rect 681 -317 682 -315
rect 688 -311 689 -309
rect 688 -317 689 -315
rect 695 -311 696 -309
rect 698 -311 699 -309
rect 695 -317 696 -315
rect 698 -317 699 -315
rect 705 -311 706 -309
rect 702 -317 703 -315
rect 709 -311 710 -309
rect 709 -317 710 -315
rect 716 -311 717 -309
rect 716 -317 717 -315
rect 723 -311 724 -309
rect 723 -317 724 -315
rect 730 -311 731 -309
rect 730 -317 731 -315
rect 737 -311 738 -309
rect 737 -317 738 -315
rect 744 -311 745 -309
rect 744 -317 745 -315
rect 751 -311 752 -309
rect 751 -317 752 -315
rect 758 -311 759 -309
rect 758 -317 759 -315
rect 765 -311 766 -309
rect 765 -317 766 -315
rect 772 -311 773 -309
rect 772 -317 773 -315
rect 779 -311 780 -309
rect 779 -317 780 -315
rect 786 -311 787 -309
rect 786 -317 787 -315
rect 793 -311 794 -309
rect 793 -317 794 -315
rect 800 -311 801 -309
rect 800 -317 801 -315
rect 807 -311 808 -309
rect 807 -317 808 -315
rect 814 -311 815 -309
rect 814 -317 815 -315
rect 821 -311 822 -309
rect 821 -317 822 -315
rect 828 -311 829 -309
rect 828 -317 829 -315
rect 835 -311 836 -309
rect 835 -317 836 -315
rect 842 -311 843 -309
rect 842 -317 843 -315
rect 849 -311 850 -309
rect 849 -317 850 -315
rect 856 -311 857 -309
rect 856 -317 857 -315
rect 863 -311 864 -309
rect 863 -317 864 -315
rect 870 -311 871 -309
rect 870 -317 871 -315
rect 877 -311 878 -309
rect 877 -317 878 -315
rect 884 -311 885 -309
rect 884 -317 885 -315
rect 891 -311 892 -309
rect 891 -317 892 -315
rect 898 -311 899 -309
rect 898 -317 899 -315
rect 905 -311 906 -309
rect 905 -317 906 -315
rect 912 -311 913 -309
rect 912 -317 913 -315
rect 919 -311 920 -309
rect 919 -317 920 -315
rect 926 -311 927 -309
rect 926 -317 927 -315
rect 933 -311 934 -309
rect 933 -317 934 -315
rect 940 -311 941 -309
rect 940 -317 941 -315
rect 947 -311 948 -309
rect 947 -317 948 -315
rect 954 -311 955 -309
rect 954 -317 955 -315
rect 961 -311 962 -309
rect 961 -317 962 -315
rect 968 -311 969 -309
rect 968 -317 969 -315
rect 975 -311 976 -309
rect 975 -317 976 -315
rect 982 -311 983 -309
rect 982 -317 983 -315
rect 989 -311 990 -309
rect 989 -317 990 -315
rect 996 -311 997 -309
rect 996 -317 997 -315
rect 1003 -311 1004 -309
rect 1003 -317 1004 -315
rect 1010 -311 1011 -309
rect 1010 -317 1011 -315
rect 1017 -311 1018 -309
rect 1017 -317 1018 -315
rect 1024 -311 1025 -309
rect 1024 -317 1025 -315
rect 1031 -311 1032 -309
rect 1031 -317 1032 -315
rect 1038 -311 1039 -309
rect 1038 -317 1039 -315
rect 1045 -311 1046 -309
rect 1045 -317 1046 -315
rect 1052 -311 1053 -309
rect 1052 -317 1053 -315
rect 1059 -311 1060 -309
rect 1059 -317 1060 -315
rect 1066 -311 1067 -309
rect 1066 -317 1067 -315
rect 1073 -311 1074 -309
rect 1073 -317 1074 -315
rect 1080 -311 1081 -309
rect 1080 -317 1081 -315
rect 1087 -311 1088 -309
rect 1087 -317 1088 -315
rect 1094 -311 1095 -309
rect 1094 -317 1095 -315
rect 1101 -311 1102 -309
rect 1101 -317 1102 -315
rect 1108 -311 1109 -309
rect 1108 -317 1109 -315
rect 1115 -311 1116 -309
rect 1115 -317 1116 -315
rect 1122 -311 1123 -309
rect 1122 -317 1123 -315
rect 1129 -311 1130 -309
rect 1129 -317 1130 -315
rect 1136 -311 1137 -309
rect 1136 -317 1137 -315
rect 1143 -311 1144 -309
rect 1143 -317 1144 -315
rect 1150 -311 1151 -309
rect 1153 -311 1154 -309
rect 1178 -311 1179 -309
rect 1178 -317 1179 -315
rect 1500 -311 1501 -309
rect 1500 -317 1501 -315
rect 2 -400 3 -398
rect 2 -406 3 -404
rect 9 -400 10 -398
rect 9 -406 10 -404
rect 16 -400 17 -398
rect 16 -406 17 -404
rect 23 -400 24 -398
rect 26 -400 27 -398
rect 23 -406 24 -404
rect 26 -406 27 -404
rect 30 -400 31 -398
rect 30 -406 31 -404
rect 37 -400 38 -398
rect 40 -400 41 -398
rect 37 -406 38 -404
rect 44 -400 45 -398
rect 47 -400 48 -398
rect 44 -406 45 -404
rect 47 -406 48 -404
rect 51 -400 52 -398
rect 51 -406 52 -404
rect 58 -400 59 -398
rect 61 -400 62 -398
rect 58 -406 59 -404
rect 61 -406 62 -404
rect 65 -400 66 -398
rect 65 -406 66 -404
rect 72 -400 73 -398
rect 75 -400 76 -398
rect 75 -406 76 -404
rect 79 -400 80 -398
rect 82 -400 83 -398
rect 79 -406 80 -404
rect 82 -406 83 -404
rect 86 -400 87 -398
rect 89 -400 90 -398
rect 86 -406 87 -404
rect 89 -406 90 -404
rect 93 -400 94 -398
rect 93 -406 94 -404
rect 100 -400 101 -398
rect 100 -406 101 -404
rect 107 -400 108 -398
rect 107 -406 108 -404
rect 114 -400 115 -398
rect 114 -406 115 -404
rect 121 -400 122 -398
rect 124 -400 125 -398
rect 124 -406 125 -404
rect 128 -400 129 -398
rect 128 -406 129 -404
rect 135 -400 136 -398
rect 135 -406 136 -404
rect 142 -400 143 -398
rect 142 -406 143 -404
rect 149 -400 150 -398
rect 149 -406 150 -404
rect 156 -400 157 -398
rect 156 -406 157 -404
rect 163 -400 164 -398
rect 163 -406 164 -404
rect 170 -400 171 -398
rect 170 -406 171 -404
rect 177 -400 178 -398
rect 177 -406 178 -404
rect 184 -400 185 -398
rect 184 -406 185 -404
rect 191 -400 192 -398
rect 191 -406 192 -404
rect 198 -400 199 -398
rect 198 -406 199 -404
rect 205 -400 206 -398
rect 205 -406 206 -404
rect 212 -400 213 -398
rect 212 -406 213 -404
rect 219 -400 220 -398
rect 219 -406 220 -404
rect 226 -400 227 -398
rect 226 -406 227 -404
rect 233 -400 234 -398
rect 233 -406 234 -404
rect 240 -400 241 -398
rect 240 -406 241 -404
rect 247 -400 248 -398
rect 247 -406 248 -404
rect 254 -400 255 -398
rect 254 -406 255 -404
rect 261 -400 262 -398
rect 264 -400 265 -398
rect 261 -406 262 -404
rect 264 -406 265 -404
rect 268 -400 269 -398
rect 268 -406 269 -404
rect 275 -400 276 -398
rect 275 -406 276 -404
rect 282 -400 283 -398
rect 282 -406 283 -404
rect 289 -400 290 -398
rect 289 -406 290 -404
rect 296 -400 297 -398
rect 296 -406 297 -404
rect 303 -400 304 -398
rect 303 -406 304 -404
rect 310 -400 311 -398
rect 310 -406 311 -404
rect 317 -400 318 -398
rect 317 -406 318 -404
rect 324 -400 325 -398
rect 324 -406 325 -404
rect 331 -400 332 -398
rect 331 -406 332 -404
rect 338 -400 339 -398
rect 338 -406 339 -404
rect 345 -400 346 -398
rect 345 -406 346 -404
rect 352 -400 353 -398
rect 352 -406 353 -404
rect 359 -400 360 -398
rect 359 -406 360 -404
rect 366 -400 367 -398
rect 366 -406 367 -404
rect 373 -400 374 -398
rect 373 -406 374 -404
rect 380 -400 381 -398
rect 380 -406 381 -404
rect 387 -400 388 -398
rect 387 -406 388 -404
rect 397 -400 398 -398
rect 394 -406 395 -404
rect 397 -406 398 -404
rect 401 -400 402 -398
rect 401 -406 402 -404
rect 408 -400 409 -398
rect 411 -400 412 -398
rect 408 -406 409 -404
rect 411 -406 412 -404
rect 415 -400 416 -398
rect 415 -406 416 -404
rect 422 -400 423 -398
rect 422 -406 423 -404
rect 429 -400 430 -398
rect 429 -406 430 -404
rect 436 -400 437 -398
rect 436 -406 437 -404
rect 443 -400 444 -398
rect 443 -406 444 -404
rect 450 -400 451 -398
rect 450 -406 451 -404
rect 457 -400 458 -398
rect 457 -406 458 -404
rect 464 -400 465 -398
rect 464 -406 465 -404
rect 471 -400 472 -398
rect 471 -406 472 -404
rect 478 -400 479 -398
rect 478 -406 479 -404
rect 485 -400 486 -398
rect 485 -406 486 -404
rect 492 -400 493 -398
rect 492 -406 493 -404
rect 499 -400 500 -398
rect 502 -400 503 -398
rect 499 -406 500 -404
rect 502 -406 503 -404
rect 506 -400 507 -398
rect 509 -400 510 -398
rect 513 -400 514 -398
rect 516 -400 517 -398
rect 516 -406 517 -404
rect 520 -400 521 -398
rect 520 -406 521 -404
rect 527 -400 528 -398
rect 527 -406 528 -404
rect 534 -400 535 -398
rect 534 -406 535 -404
rect 541 -400 542 -398
rect 541 -406 542 -404
rect 548 -400 549 -398
rect 551 -400 552 -398
rect 548 -406 549 -404
rect 551 -406 552 -404
rect 555 -400 556 -398
rect 555 -406 556 -404
rect 565 -400 566 -398
rect 562 -406 563 -404
rect 565 -406 566 -404
rect 569 -400 570 -398
rect 572 -400 573 -398
rect 569 -406 570 -404
rect 572 -406 573 -404
rect 576 -400 577 -398
rect 576 -406 577 -404
rect 583 -400 584 -398
rect 583 -406 584 -404
rect 590 -400 591 -398
rect 590 -406 591 -404
rect 593 -406 594 -404
rect 597 -400 598 -398
rect 597 -406 598 -404
rect 604 -400 605 -398
rect 604 -406 605 -404
rect 611 -400 612 -398
rect 611 -406 612 -404
rect 618 -400 619 -398
rect 618 -406 619 -404
rect 625 -400 626 -398
rect 625 -406 626 -404
rect 632 -400 633 -398
rect 632 -406 633 -404
rect 639 -400 640 -398
rect 642 -400 643 -398
rect 642 -406 643 -404
rect 646 -400 647 -398
rect 646 -406 647 -404
rect 653 -400 654 -398
rect 653 -406 654 -404
rect 660 -400 661 -398
rect 660 -406 661 -404
rect 663 -406 664 -404
rect 667 -400 668 -398
rect 670 -400 671 -398
rect 667 -406 668 -404
rect 670 -406 671 -404
rect 674 -400 675 -398
rect 674 -406 675 -404
rect 681 -400 682 -398
rect 681 -406 682 -404
rect 688 -400 689 -398
rect 688 -406 689 -404
rect 695 -400 696 -398
rect 695 -406 696 -404
rect 702 -400 703 -398
rect 702 -406 703 -404
rect 709 -400 710 -398
rect 709 -406 710 -404
rect 716 -400 717 -398
rect 716 -406 717 -404
rect 723 -400 724 -398
rect 723 -406 724 -404
rect 730 -400 731 -398
rect 730 -406 731 -404
rect 737 -400 738 -398
rect 737 -406 738 -404
rect 744 -400 745 -398
rect 744 -406 745 -404
rect 751 -400 752 -398
rect 751 -406 752 -404
rect 758 -400 759 -398
rect 758 -406 759 -404
rect 765 -400 766 -398
rect 765 -406 766 -404
rect 772 -400 773 -398
rect 772 -406 773 -404
rect 779 -400 780 -398
rect 779 -406 780 -404
rect 786 -400 787 -398
rect 786 -406 787 -404
rect 793 -400 794 -398
rect 793 -406 794 -404
rect 800 -400 801 -398
rect 800 -406 801 -404
rect 807 -400 808 -398
rect 807 -406 808 -404
rect 814 -400 815 -398
rect 814 -406 815 -404
rect 821 -400 822 -398
rect 821 -406 822 -404
rect 828 -400 829 -398
rect 828 -406 829 -404
rect 835 -400 836 -398
rect 835 -406 836 -404
rect 842 -400 843 -398
rect 842 -406 843 -404
rect 849 -400 850 -398
rect 849 -406 850 -404
rect 856 -400 857 -398
rect 856 -406 857 -404
rect 863 -400 864 -398
rect 863 -406 864 -404
rect 870 -400 871 -398
rect 870 -406 871 -404
rect 877 -400 878 -398
rect 877 -406 878 -404
rect 884 -400 885 -398
rect 884 -406 885 -404
rect 891 -400 892 -398
rect 891 -406 892 -404
rect 898 -400 899 -398
rect 898 -406 899 -404
rect 905 -400 906 -398
rect 905 -406 906 -404
rect 912 -400 913 -398
rect 912 -406 913 -404
rect 919 -400 920 -398
rect 919 -406 920 -404
rect 926 -400 927 -398
rect 926 -406 927 -404
rect 933 -400 934 -398
rect 933 -406 934 -404
rect 940 -400 941 -398
rect 940 -406 941 -404
rect 947 -400 948 -398
rect 947 -406 948 -404
rect 954 -400 955 -398
rect 954 -406 955 -404
rect 961 -400 962 -398
rect 961 -406 962 -404
rect 968 -400 969 -398
rect 968 -406 969 -404
rect 975 -400 976 -398
rect 975 -406 976 -404
rect 982 -400 983 -398
rect 982 -406 983 -404
rect 989 -400 990 -398
rect 989 -406 990 -404
rect 996 -400 997 -398
rect 996 -406 997 -404
rect 1003 -400 1004 -398
rect 1003 -406 1004 -404
rect 1010 -400 1011 -398
rect 1010 -406 1011 -404
rect 1017 -400 1018 -398
rect 1017 -406 1018 -404
rect 1024 -400 1025 -398
rect 1024 -406 1025 -404
rect 1031 -400 1032 -398
rect 1031 -406 1032 -404
rect 1038 -400 1039 -398
rect 1038 -406 1039 -404
rect 1045 -400 1046 -398
rect 1045 -406 1046 -404
rect 1052 -400 1053 -398
rect 1052 -406 1053 -404
rect 1059 -400 1060 -398
rect 1059 -406 1060 -404
rect 1066 -400 1067 -398
rect 1066 -406 1067 -404
rect 1073 -400 1074 -398
rect 1073 -406 1074 -404
rect 1080 -400 1081 -398
rect 1080 -406 1081 -404
rect 1087 -400 1088 -398
rect 1087 -406 1088 -404
rect 1094 -400 1095 -398
rect 1094 -406 1095 -404
rect 1101 -400 1102 -398
rect 1101 -406 1102 -404
rect 1108 -400 1109 -398
rect 1108 -406 1109 -404
rect 1115 -400 1116 -398
rect 1115 -406 1116 -404
rect 1122 -400 1123 -398
rect 1122 -406 1123 -404
rect 1129 -400 1130 -398
rect 1129 -406 1130 -404
rect 1136 -400 1137 -398
rect 1136 -406 1137 -404
rect 1143 -400 1144 -398
rect 1143 -406 1144 -404
rect 1150 -400 1151 -398
rect 1150 -406 1151 -404
rect 1157 -400 1158 -398
rect 1157 -406 1158 -404
rect 1164 -400 1165 -398
rect 1164 -406 1165 -404
rect 1171 -400 1172 -398
rect 1171 -406 1172 -404
rect 1178 -400 1179 -398
rect 1178 -406 1179 -404
rect 1185 -400 1186 -398
rect 1185 -406 1186 -404
rect 1192 -400 1193 -398
rect 1192 -406 1193 -404
rect 1202 -400 1203 -398
rect 1199 -406 1200 -404
rect 1202 -406 1203 -404
rect 1209 -400 1210 -398
rect 1209 -406 1210 -404
rect 1500 -400 1501 -398
rect 1500 -406 1501 -404
rect 2 -521 3 -519
rect 5 -521 6 -519
rect 9 -515 10 -513
rect 9 -521 10 -519
rect 16 -515 17 -513
rect 16 -521 17 -519
rect 23 -515 24 -513
rect 23 -521 24 -519
rect 30 -515 31 -513
rect 33 -515 34 -513
rect 33 -521 34 -519
rect 37 -515 38 -513
rect 40 -515 41 -513
rect 37 -521 38 -519
rect 40 -521 41 -519
rect 44 -515 45 -513
rect 44 -521 45 -519
rect 51 -515 52 -513
rect 51 -521 52 -519
rect 58 -515 59 -513
rect 58 -521 59 -519
rect 65 -515 66 -513
rect 65 -521 66 -519
rect 72 -515 73 -513
rect 75 -515 76 -513
rect 72 -521 73 -519
rect 79 -515 80 -513
rect 79 -521 80 -519
rect 86 -515 87 -513
rect 89 -515 90 -513
rect 86 -521 87 -519
rect 89 -521 90 -519
rect 93 -515 94 -513
rect 93 -521 94 -519
rect 100 -515 101 -513
rect 100 -521 101 -519
rect 107 -515 108 -513
rect 110 -515 111 -513
rect 107 -521 108 -519
rect 110 -521 111 -519
rect 114 -515 115 -513
rect 114 -521 115 -519
rect 121 -515 122 -513
rect 121 -521 122 -519
rect 128 -515 129 -513
rect 128 -521 129 -519
rect 135 -515 136 -513
rect 138 -515 139 -513
rect 135 -521 136 -519
rect 138 -521 139 -519
rect 142 -515 143 -513
rect 145 -515 146 -513
rect 142 -521 143 -519
rect 145 -521 146 -519
rect 149 -515 150 -513
rect 149 -521 150 -519
rect 159 -515 160 -513
rect 156 -521 157 -519
rect 159 -521 160 -519
rect 163 -515 164 -513
rect 163 -521 164 -519
rect 170 -515 171 -513
rect 170 -521 171 -519
rect 177 -515 178 -513
rect 177 -521 178 -519
rect 184 -515 185 -513
rect 184 -521 185 -519
rect 191 -515 192 -513
rect 191 -521 192 -519
rect 198 -515 199 -513
rect 201 -515 202 -513
rect 198 -521 199 -519
rect 201 -521 202 -519
rect 205 -515 206 -513
rect 205 -521 206 -519
rect 212 -515 213 -513
rect 212 -521 213 -519
rect 219 -515 220 -513
rect 219 -521 220 -519
rect 226 -515 227 -513
rect 226 -521 227 -519
rect 233 -515 234 -513
rect 233 -521 234 -519
rect 240 -515 241 -513
rect 240 -521 241 -519
rect 247 -521 248 -519
rect 250 -521 251 -519
rect 254 -521 255 -519
rect 257 -521 258 -519
rect 261 -515 262 -513
rect 261 -521 262 -519
rect 268 -515 269 -513
rect 268 -521 269 -519
rect 275 -515 276 -513
rect 275 -521 276 -519
rect 282 -515 283 -513
rect 282 -521 283 -519
rect 289 -515 290 -513
rect 289 -521 290 -519
rect 296 -515 297 -513
rect 296 -521 297 -519
rect 303 -515 304 -513
rect 303 -521 304 -519
rect 310 -515 311 -513
rect 310 -521 311 -519
rect 317 -515 318 -513
rect 317 -521 318 -519
rect 324 -515 325 -513
rect 324 -521 325 -519
rect 331 -515 332 -513
rect 331 -521 332 -519
rect 338 -515 339 -513
rect 338 -521 339 -519
rect 345 -515 346 -513
rect 345 -521 346 -519
rect 352 -515 353 -513
rect 352 -521 353 -519
rect 359 -515 360 -513
rect 359 -521 360 -519
rect 366 -515 367 -513
rect 366 -521 367 -519
rect 373 -515 374 -513
rect 373 -521 374 -519
rect 380 -515 381 -513
rect 383 -515 384 -513
rect 380 -521 381 -519
rect 383 -521 384 -519
rect 387 -515 388 -513
rect 387 -521 388 -519
rect 394 -515 395 -513
rect 394 -521 395 -519
rect 401 -515 402 -513
rect 401 -521 402 -519
rect 408 -515 409 -513
rect 408 -521 409 -519
rect 415 -515 416 -513
rect 415 -521 416 -519
rect 418 -521 419 -519
rect 422 -515 423 -513
rect 425 -515 426 -513
rect 422 -521 423 -519
rect 425 -521 426 -519
rect 429 -515 430 -513
rect 429 -521 430 -519
rect 436 -515 437 -513
rect 436 -521 437 -519
rect 443 -515 444 -513
rect 443 -521 444 -519
rect 450 -515 451 -513
rect 450 -521 451 -519
rect 457 -515 458 -513
rect 460 -515 461 -513
rect 457 -521 458 -519
rect 460 -521 461 -519
rect 464 -515 465 -513
rect 464 -521 465 -519
rect 471 -515 472 -513
rect 471 -521 472 -519
rect 478 -515 479 -513
rect 478 -521 479 -519
rect 485 -515 486 -513
rect 485 -521 486 -519
rect 492 -515 493 -513
rect 492 -521 493 -519
rect 499 -515 500 -513
rect 502 -515 503 -513
rect 499 -521 500 -519
rect 502 -521 503 -519
rect 506 -515 507 -513
rect 509 -515 510 -513
rect 506 -521 507 -519
rect 509 -521 510 -519
rect 513 -515 514 -513
rect 513 -521 514 -519
rect 520 -515 521 -513
rect 520 -521 521 -519
rect 527 -515 528 -513
rect 530 -515 531 -513
rect 530 -521 531 -519
rect 534 -515 535 -513
rect 537 -515 538 -513
rect 534 -521 535 -519
rect 541 -515 542 -513
rect 541 -521 542 -519
rect 548 -515 549 -513
rect 548 -521 549 -519
rect 555 -515 556 -513
rect 555 -521 556 -519
rect 562 -515 563 -513
rect 562 -521 563 -519
rect 569 -515 570 -513
rect 569 -521 570 -519
rect 576 -515 577 -513
rect 576 -521 577 -519
rect 583 -515 584 -513
rect 583 -521 584 -519
rect 590 -515 591 -513
rect 590 -521 591 -519
rect 597 -515 598 -513
rect 600 -515 601 -513
rect 597 -521 598 -519
rect 600 -521 601 -519
rect 604 -515 605 -513
rect 604 -521 605 -519
rect 611 -515 612 -513
rect 614 -515 615 -513
rect 611 -521 612 -519
rect 614 -521 615 -519
rect 618 -515 619 -513
rect 618 -521 619 -519
rect 625 -515 626 -513
rect 625 -521 626 -519
rect 632 -515 633 -513
rect 632 -521 633 -519
rect 639 -515 640 -513
rect 639 -521 640 -519
rect 646 -515 647 -513
rect 646 -521 647 -519
rect 653 -515 654 -513
rect 653 -521 654 -519
rect 660 -515 661 -513
rect 663 -515 664 -513
rect 660 -521 661 -519
rect 663 -521 664 -519
rect 667 -515 668 -513
rect 667 -521 668 -519
rect 674 -515 675 -513
rect 674 -521 675 -519
rect 681 -515 682 -513
rect 681 -521 682 -519
rect 688 -515 689 -513
rect 688 -521 689 -519
rect 698 -515 699 -513
rect 695 -521 696 -519
rect 698 -521 699 -519
rect 702 -515 703 -513
rect 705 -515 706 -513
rect 702 -521 703 -519
rect 705 -521 706 -519
rect 709 -515 710 -513
rect 709 -521 710 -519
rect 716 -515 717 -513
rect 716 -521 717 -519
rect 723 -515 724 -513
rect 723 -521 724 -519
rect 730 -515 731 -513
rect 730 -521 731 -519
rect 737 -515 738 -513
rect 737 -521 738 -519
rect 744 -515 745 -513
rect 744 -521 745 -519
rect 751 -515 752 -513
rect 751 -521 752 -519
rect 758 -515 759 -513
rect 758 -521 759 -519
rect 765 -515 766 -513
rect 765 -521 766 -519
rect 772 -515 773 -513
rect 772 -521 773 -519
rect 779 -515 780 -513
rect 779 -521 780 -519
rect 786 -515 787 -513
rect 786 -521 787 -519
rect 793 -515 794 -513
rect 793 -521 794 -519
rect 800 -515 801 -513
rect 800 -521 801 -519
rect 807 -515 808 -513
rect 807 -521 808 -519
rect 814 -515 815 -513
rect 814 -521 815 -519
rect 821 -515 822 -513
rect 821 -521 822 -519
rect 828 -515 829 -513
rect 828 -521 829 -519
rect 835 -515 836 -513
rect 835 -521 836 -519
rect 842 -515 843 -513
rect 842 -521 843 -519
rect 849 -515 850 -513
rect 849 -521 850 -519
rect 856 -515 857 -513
rect 856 -521 857 -519
rect 863 -515 864 -513
rect 863 -521 864 -519
rect 870 -515 871 -513
rect 870 -521 871 -519
rect 877 -515 878 -513
rect 877 -521 878 -519
rect 884 -515 885 -513
rect 884 -521 885 -519
rect 891 -515 892 -513
rect 891 -521 892 -519
rect 898 -515 899 -513
rect 898 -521 899 -519
rect 905 -515 906 -513
rect 905 -521 906 -519
rect 912 -515 913 -513
rect 912 -521 913 -519
rect 919 -515 920 -513
rect 919 -521 920 -519
rect 926 -515 927 -513
rect 926 -521 927 -519
rect 933 -515 934 -513
rect 933 -521 934 -519
rect 940 -515 941 -513
rect 940 -521 941 -519
rect 947 -515 948 -513
rect 947 -521 948 -519
rect 954 -515 955 -513
rect 954 -521 955 -519
rect 961 -515 962 -513
rect 961 -521 962 -519
rect 968 -515 969 -513
rect 968 -521 969 -519
rect 975 -515 976 -513
rect 975 -521 976 -519
rect 982 -515 983 -513
rect 982 -521 983 -519
rect 989 -515 990 -513
rect 989 -521 990 -519
rect 996 -515 997 -513
rect 996 -521 997 -519
rect 1003 -515 1004 -513
rect 1003 -521 1004 -519
rect 1010 -515 1011 -513
rect 1010 -521 1011 -519
rect 1017 -515 1018 -513
rect 1017 -521 1018 -519
rect 1024 -515 1025 -513
rect 1024 -521 1025 -519
rect 1031 -515 1032 -513
rect 1031 -521 1032 -519
rect 1038 -515 1039 -513
rect 1038 -521 1039 -519
rect 1045 -515 1046 -513
rect 1045 -521 1046 -519
rect 1052 -515 1053 -513
rect 1052 -521 1053 -519
rect 1059 -515 1060 -513
rect 1059 -521 1060 -519
rect 1066 -515 1067 -513
rect 1066 -521 1067 -519
rect 1073 -515 1074 -513
rect 1073 -521 1074 -519
rect 1080 -515 1081 -513
rect 1080 -521 1081 -519
rect 1087 -515 1088 -513
rect 1087 -521 1088 -519
rect 1094 -515 1095 -513
rect 1094 -521 1095 -519
rect 1101 -515 1102 -513
rect 1101 -521 1102 -519
rect 1108 -515 1109 -513
rect 1108 -521 1109 -519
rect 1115 -515 1116 -513
rect 1115 -521 1116 -519
rect 1122 -515 1123 -513
rect 1122 -521 1123 -519
rect 1129 -515 1130 -513
rect 1129 -521 1130 -519
rect 1136 -515 1137 -513
rect 1136 -521 1137 -519
rect 1143 -515 1144 -513
rect 1143 -521 1144 -519
rect 1150 -515 1151 -513
rect 1150 -521 1151 -519
rect 1157 -515 1158 -513
rect 1157 -521 1158 -519
rect 1164 -515 1165 -513
rect 1164 -521 1165 -519
rect 1171 -515 1172 -513
rect 1171 -521 1172 -519
rect 1178 -515 1179 -513
rect 1178 -521 1179 -519
rect 1185 -515 1186 -513
rect 1185 -521 1186 -519
rect 1192 -515 1193 -513
rect 1192 -521 1193 -519
rect 1199 -515 1200 -513
rect 1199 -521 1200 -519
rect 1206 -515 1207 -513
rect 1206 -521 1207 -519
rect 1213 -515 1214 -513
rect 1213 -521 1214 -519
rect 1220 -515 1221 -513
rect 1220 -521 1221 -519
rect 1227 -515 1228 -513
rect 1227 -521 1228 -519
rect 1234 -515 1235 -513
rect 1234 -521 1235 -519
rect 1241 -515 1242 -513
rect 1241 -521 1242 -519
rect 1248 -515 1249 -513
rect 1248 -521 1249 -519
rect 1255 -515 1256 -513
rect 1255 -521 1256 -519
rect 1262 -515 1263 -513
rect 1262 -521 1263 -519
rect 1395 -515 1396 -513
rect 1395 -521 1396 -519
rect 1500 -515 1501 -513
rect 1500 -521 1501 -519
rect 2 -630 3 -628
rect 2 -636 3 -634
rect 9 -630 10 -628
rect 9 -636 10 -634
rect 19 -630 20 -628
rect 16 -636 17 -634
rect 19 -636 20 -634
rect 23 -630 24 -628
rect 23 -636 24 -634
rect 30 -630 31 -628
rect 30 -636 31 -634
rect 37 -630 38 -628
rect 40 -630 41 -628
rect 44 -630 45 -628
rect 47 -630 48 -628
rect 44 -636 45 -634
rect 47 -636 48 -634
rect 51 -630 52 -628
rect 51 -636 52 -634
rect 58 -630 59 -628
rect 58 -636 59 -634
rect 65 -630 66 -628
rect 65 -636 66 -634
rect 72 -630 73 -628
rect 75 -630 76 -628
rect 72 -636 73 -634
rect 75 -636 76 -634
rect 79 -630 80 -628
rect 79 -636 80 -634
rect 86 -630 87 -628
rect 86 -636 87 -634
rect 93 -630 94 -628
rect 96 -630 97 -628
rect 93 -636 94 -634
rect 96 -636 97 -634
rect 100 -630 101 -628
rect 100 -636 101 -634
rect 107 -630 108 -628
rect 107 -636 108 -634
rect 114 -630 115 -628
rect 117 -630 118 -628
rect 114 -636 115 -634
rect 117 -636 118 -634
rect 121 -630 122 -628
rect 121 -636 122 -634
rect 128 -630 129 -628
rect 128 -636 129 -634
rect 135 -630 136 -628
rect 135 -636 136 -634
rect 142 -630 143 -628
rect 142 -636 143 -634
rect 149 -630 150 -628
rect 149 -636 150 -634
rect 156 -630 157 -628
rect 156 -636 157 -634
rect 163 -630 164 -628
rect 163 -636 164 -634
rect 170 -630 171 -628
rect 170 -636 171 -634
rect 173 -636 174 -634
rect 177 -630 178 -628
rect 177 -636 178 -634
rect 184 -630 185 -628
rect 184 -636 185 -634
rect 191 -630 192 -628
rect 191 -636 192 -634
rect 198 -630 199 -628
rect 198 -636 199 -634
rect 205 -630 206 -628
rect 205 -636 206 -634
rect 212 -630 213 -628
rect 212 -636 213 -634
rect 219 -630 220 -628
rect 219 -636 220 -634
rect 226 -630 227 -628
rect 226 -636 227 -634
rect 233 -630 234 -628
rect 233 -636 234 -634
rect 240 -630 241 -628
rect 240 -636 241 -634
rect 247 -630 248 -628
rect 247 -636 248 -634
rect 254 -630 255 -628
rect 254 -636 255 -634
rect 261 -630 262 -628
rect 261 -636 262 -634
rect 268 -630 269 -628
rect 271 -630 272 -628
rect 271 -636 272 -634
rect 275 -630 276 -628
rect 275 -636 276 -634
rect 282 -630 283 -628
rect 282 -636 283 -634
rect 289 -630 290 -628
rect 289 -636 290 -634
rect 296 -630 297 -628
rect 296 -636 297 -634
rect 303 -630 304 -628
rect 303 -636 304 -634
rect 310 -636 311 -634
rect 313 -636 314 -634
rect 317 -630 318 -628
rect 317 -636 318 -634
rect 324 -630 325 -628
rect 324 -636 325 -634
rect 331 -630 332 -628
rect 331 -636 332 -634
rect 338 -630 339 -628
rect 338 -636 339 -634
rect 348 -630 349 -628
rect 345 -636 346 -634
rect 348 -636 349 -634
rect 352 -630 353 -628
rect 355 -636 356 -634
rect 359 -630 360 -628
rect 359 -636 360 -634
rect 366 -630 367 -628
rect 366 -636 367 -634
rect 373 -630 374 -628
rect 373 -636 374 -634
rect 380 -630 381 -628
rect 380 -636 381 -634
rect 383 -636 384 -634
rect 387 -630 388 -628
rect 390 -630 391 -628
rect 387 -636 388 -634
rect 390 -636 391 -634
rect 394 -630 395 -628
rect 394 -636 395 -634
rect 401 -630 402 -628
rect 401 -636 402 -634
rect 408 -630 409 -628
rect 408 -636 409 -634
rect 415 -630 416 -628
rect 418 -630 419 -628
rect 415 -636 416 -634
rect 418 -636 419 -634
rect 422 -630 423 -628
rect 422 -636 423 -634
rect 429 -630 430 -628
rect 429 -636 430 -634
rect 436 -630 437 -628
rect 436 -636 437 -634
rect 443 -630 444 -628
rect 446 -630 447 -628
rect 443 -636 444 -634
rect 446 -636 447 -634
rect 450 -630 451 -628
rect 450 -636 451 -634
rect 457 -630 458 -628
rect 457 -636 458 -634
rect 464 -630 465 -628
rect 464 -636 465 -634
rect 471 -630 472 -628
rect 471 -636 472 -634
rect 481 -630 482 -628
rect 478 -636 479 -634
rect 481 -636 482 -634
rect 485 -630 486 -628
rect 485 -636 486 -634
rect 492 -630 493 -628
rect 492 -636 493 -634
rect 499 -630 500 -628
rect 499 -636 500 -634
rect 506 -630 507 -628
rect 509 -630 510 -628
rect 506 -636 507 -634
rect 509 -636 510 -634
rect 513 -630 514 -628
rect 513 -636 514 -634
rect 520 -630 521 -628
rect 520 -636 521 -634
rect 527 -630 528 -628
rect 527 -636 528 -634
rect 534 -630 535 -628
rect 534 -636 535 -634
rect 541 -630 542 -628
rect 541 -636 542 -634
rect 548 -630 549 -628
rect 548 -636 549 -634
rect 555 -630 556 -628
rect 555 -636 556 -634
rect 562 -630 563 -628
rect 565 -630 566 -628
rect 562 -636 563 -634
rect 569 -630 570 -628
rect 569 -636 570 -634
rect 576 -630 577 -628
rect 576 -636 577 -634
rect 583 -630 584 -628
rect 583 -636 584 -634
rect 590 -630 591 -628
rect 590 -636 591 -634
rect 597 -630 598 -628
rect 597 -636 598 -634
rect 604 -630 605 -628
rect 604 -636 605 -634
rect 611 -630 612 -628
rect 614 -630 615 -628
rect 611 -636 612 -634
rect 614 -636 615 -634
rect 618 -630 619 -628
rect 618 -636 619 -634
rect 625 -630 626 -628
rect 628 -630 629 -628
rect 625 -636 626 -634
rect 628 -636 629 -634
rect 632 -630 633 -628
rect 635 -630 636 -628
rect 632 -636 633 -634
rect 635 -636 636 -634
rect 639 -630 640 -628
rect 639 -636 640 -634
rect 646 -630 647 -628
rect 646 -636 647 -634
rect 653 -630 654 -628
rect 653 -636 654 -634
rect 660 -630 661 -628
rect 660 -636 661 -634
rect 667 -630 668 -628
rect 670 -630 671 -628
rect 667 -636 668 -634
rect 674 -630 675 -628
rect 674 -636 675 -634
rect 681 -630 682 -628
rect 681 -636 682 -634
rect 688 -630 689 -628
rect 688 -636 689 -634
rect 695 -630 696 -628
rect 695 -636 696 -634
rect 702 -630 703 -628
rect 702 -636 703 -634
rect 709 -630 710 -628
rect 709 -636 710 -634
rect 716 -630 717 -628
rect 716 -636 717 -634
rect 723 -630 724 -628
rect 723 -636 724 -634
rect 730 -630 731 -628
rect 730 -636 731 -634
rect 737 -630 738 -628
rect 737 -636 738 -634
rect 747 -630 748 -628
rect 744 -636 745 -634
rect 747 -636 748 -634
rect 751 -630 752 -628
rect 751 -636 752 -634
rect 758 -630 759 -628
rect 758 -636 759 -634
rect 765 -630 766 -628
rect 765 -636 766 -634
rect 772 -630 773 -628
rect 772 -636 773 -634
rect 779 -630 780 -628
rect 779 -636 780 -634
rect 786 -630 787 -628
rect 786 -636 787 -634
rect 793 -630 794 -628
rect 793 -636 794 -634
rect 800 -630 801 -628
rect 800 -636 801 -634
rect 807 -630 808 -628
rect 807 -636 808 -634
rect 814 -630 815 -628
rect 814 -636 815 -634
rect 821 -630 822 -628
rect 821 -636 822 -634
rect 828 -630 829 -628
rect 828 -636 829 -634
rect 835 -630 836 -628
rect 835 -636 836 -634
rect 842 -630 843 -628
rect 842 -636 843 -634
rect 849 -630 850 -628
rect 849 -636 850 -634
rect 856 -630 857 -628
rect 856 -636 857 -634
rect 863 -630 864 -628
rect 863 -636 864 -634
rect 870 -630 871 -628
rect 870 -636 871 -634
rect 877 -630 878 -628
rect 877 -636 878 -634
rect 884 -630 885 -628
rect 884 -636 885 -634
rect 891 -630 892 -628
rect 891 -636 892 -634
rect 898 -630 899 -628
rect 898 -636 899 -634
rect 905 -630 906 -628
rect 905 -636 906 -634
rect 912 -630 913 -628
rect 912 -636 913 -634
rect 919 -630 920 -628
rect 919 -636 920 -634
rect 926 -630 927 -628
rect 926 -636 927 -634
rect 933 -630 934 -628
rect 933 -636 934 -634
rect 940 -630 941 -628
rect 940 -636 941 -634
rect 947 -630 948 -628
rect 947 -636 948 -634
rect 954 -630 955 -628
rect 954 -636 955 -634
rect 961 -630 962 -628
rect 961 -636 962 -634
rect 964 -636 965 -634
rect 968 -630 969 -628
rect 968 -636 969 -634
rect 975 -630 976 -628
rect 975 -636 976 -634
rect 982 -630 983 -628
rect 982 -636 983 -634
rect 989 -630 990 -628
rect 989 -636 990 -634
rect 996 -630 997 -628
rect 996 -636 997 -634
rect 1003 -630 1004 -628
rect 1003 -636 1004 -634
rect 1010 -630 1011 -628
rect 1010 -636 1011 -634
rect 1017 -630 1018 -628
rect 1017 -636 1018 -634
rect 1024 -630 1025 -628
rect 1024 -636 1025 -634
rect 1031 -630 1032 -628
rect 1034 -630 1035 -628
rect 1034 -636 1035 -634
rect 1038 -630 1039 -628
rect 1038 -636 1039 -634
rect 1045 -630 1046 -628
rect 1045 -636 1046 -634
rect 1052 -630 1053 -628
rect 1052 -636 1053 -634
rect 1059 -630 1060 -628
rect 1059 -636 1060 -634
rect 1066 -630 1067 -628
rect 1066 -636 1067 -634
rect 1073 -630 1074 -628
rect 1073 -636 1074 -634
rect 1080 -630 1081 -628
rect 1080 -636 1081 -634
rect 1087 -630 1088 -628
rect 1087 -636 1088 -634
rect 1094 -630 1095 -628
rect 1094 -636 1095 -634
rect 1101 -630 1102 -628
rect 1101 -636 1102 -634
rect 1108 -630 1109 -628
rect 1108 -636 1109 -634
rect 1115 -630 1116 -628
rect 1115 -636 1116 -634
rect 1122 -630 1123 -628
rect 1122 -636 1123 -634
rect 1129 -630 1130 -628
rect 1129 -636 1130 -634
rect 1136 -630 1137 -628
rect 1136 -636 1137 -634
rect 1143 -630 1144 -628
rect 1143 -636 1144 -634
rect 1150 -630 1151 -628
rect 1150 -636 1151 -634
rect 1157 -630 1158 -628
rect 1157 -636 1158 -634
rect 1164 -630 1165 -628
rect 1164 -636 1165 -634
rect 1171 -630 1172 -628
rect 1171 -636 1172 -634
rect 1178 -630 1179 -628
rect 1178 -636 1179 -634
rect 1185 -630 1186 -628
rect 1185 -636 1186 -634
rect 1192 -630 1193 -628
rect 1192 -636 1193 -634
rect 1199 -630 1200 -628
rect 1199 -636 1200 -634
rect 1206 -630 1207 -628
rect 1206 -636 1207 -634
rect 1213 -630 1214 -628
rect 1213 -636 1214 -634
rect 1220 -630 1221 -628
rect 1220 -636 1221 -634
rect 1227 -630 1228 -628
rect 1227 -636 1228 -634
rect 1234 -630 1235 -628
rect 1234 -636 1235 -634
rect 1241 -630 1242 -628
rect 1241 -636 1242 -634
rect 1248 -630 1249 -628
rect 1248 -636 1249 -634
rect 1255 -630 1256 -628
rect 1255 -636 1256 -634
rect 1262 -630 1263 -628
rect 1262 -636 1263 -634
rect 1269 -630 1270 -628
rect 1269 -636 1270 -634
rect 1276 -630 1277 -628
rect 1276 -636 1277 -634
rect 1283 -630 1284 -628
rect 1283 -636 1284 -634
rect 1290 -630 1291 -628
rect 1290 -636 1291 -634
rect 1297 -630 1298 -628
rect 1297 -636 1298 -634
rect 1304 -630 1305 -628
rect 1304 -636 1305 -634
rect 1311 -630 1312 -628
rect 1311 -636 1312 -634
rect 1318 -630 1319 -628
rect 1318 -636 1319 -634
rect 1325 -630 1326 -628
rect 1325 -636 1326 -634
rect 1332 -630 1333 -628
rect 1332 -636 1333 -634
rect 1339 -630 1340 -628
rect 1339 -636 1340 -634
rect 1346 -630 1347 -628
rect 1346 -636 1347 -634
rect 1353 -630 1354 -628
rect 1353 -636 1354 -634
rect 1360 -630 1361 -628
rect 1360 -636 1361 -634
rect 1367 -630 1368 -628
rect 1367 -636 1368 -634
rect 1374 -630 1375 -628
rect 1374 -636 1375 -634
rect 1472 -630 1473 -628
rect 1472 -636 1473 -634
rect 1507 -630 1508 -628
rect 1507 -636 1508 -634
rect 5 -749 6 -747
rect 2 -755 3 -753
rect 12 -749 13 -747
rect 9 -755 10 -753
rect 12 -755 13 -753
rect 16 -749 17 -747
rect 16 -755 17 -753
rect 23 -749 24 -747
rect 23 -755 24 -753
rect 30 -749 31 -747
rect 30 -755 31 -753
rect 37 -749 38 -747
rect 37 -755 38 -753
rect 44 -749 45 -747
rect 44 -755 45 -753
rect 51 -749 52 -747
rect 51 -755 52 -753
rect 58 -749 59 -747
rect 61 -749 62 -747
rect 58 -755 59 -753
rect 61 -755 62 -753
rect 65 -749 66 -747
rect 65 -755 66 -753
rect 72 -749 73 -747
rect 75 -749 76 -747
rect 72 -755 73 -753
rect 75 -755 76 -753
rect 79 -749 80 -747
rect 79 -755 80 -753
rect 86 -749 87 -747
rect 86 -755 87 -753
rect 93 -749 94 -747
rect 93 -755 94 -753
rect 100 -749 101 -747
rect 103 -749 104 -747
rect 100 -755 101 -753
rect 103 -755 104 -753
rect 107 -749 108 -747
rect 107 -755 108 -753
rect 114 -749 115 -747
rect 117 -749 118 -747
rect 114 -755 115 -753
rect 117 -755 118 -753
rect 121 -749 122 -747
rect 121 -755 122 -753
rect 128 -749 129 -747
rect 128 -755 129 -753
rect 135 -755 136 -753
rect 138 -755 139 -753
rect 142 -749 143 -747
rect 142 -755 143 -753
rect 149 -749 150 -747
rect 149 -755 150 -753
rect 156 -749 157 -747
rect 156 -755 157 -753
rect 163 -749 164 -747
rect 163 -755 164 -753
rect 170 -749 171 -747
rect 170 -755 171 -753
rect 177 -749 178 -747
rect 177 -755 178 -753
rect 184 -749 185 -747
rect 184 -755 185 -753
rect 191 -749 192 -747
rect 191 -755 192 -753
rect 198 -749 199 -747
rect 198 -755 199 -753
rect 205 -749 206 -747
rect 205 -755 206 -753
rect 212 -749 213 -747
rect 212 -755 213 -753
rect 219 -749 220 -747
rect 219 -755 220 -753
rect 226 -749 227 -747
rect 226 -755 227 -753
rect 233 -749 234 -747
rect 233 -755 234 -753
rect 240 -749 241 -747
rect 240 -755 241 -753
rect 247 -749 248 -747
rect 247 -755 248 -753
rect 254 -749 255 -747
rect 254 -755 255 -753
rect 261 -749 262 -747
rect 261 -755 262 -753
rect 268 -749 269 -747
rect 271 -749 272 -747
rect 268 -755 269 -753
rect 271 -755 272 -753
rect 275 -749 276 -747
rect 275 -755 276 -753
rect 282 -749 283 -747
rect 282 -755 283 -753
rect 289 -749 290 -747
rect 289 -755 290 -753
rect 296 -749 297 -747
rect 296 -755 297 -753
rect 303 -749 304 -747
rect 303 -755 304 -753
rect 310 -749 311 -747
rect 310 -755 311 -753
rect 317 -749 318 -747
rect 317 -755 318 -753
rect 324 -749 325 -747
rect 324 -755 325 -753
rect 331 -749 332 -747
rect 331 -755 332 -753
rect 338 -749 339 -747
rect 338 -755 339 -753
rect 345 -749 346 -747
rect 345 -755 346 -753
rect 352 -749 353 -747
rect 355 -749 356 -747
rect 352 -755 353 -753
rect 355 -755 356 -753
rect 359 -749 360 -747
rect 359 -755 360 -753
rect 366 -749 367 -747
rect 366 -755 367 -753
rect 369 -755 370 -753
rect 373 -749 374 -747
rect 373 -755 374 -753
rect 380 -749 381 -747
rect 380 -755 381 -753
rect 387 -749 388 -747
rect 387 -755 388 -753
rect 394 -749 395 -747
rect 394 -755 395 -753
rect 401 -749 402 -747
rect 401 -755 402 -753
rect 408 -749 409 -747
rect 408 -755 409 -753
rect 415 -749 416 -747
rect 422 -749 423 -747
rect 425 -749 426 -747
rect 422 -755 423 -753
rect 425 -755 426 -753
rect 429 -749 430 -747
rect 429 -755 430 -753
rect 436 -749 437 -747
rect 436 -755 437 -753
rect 443 -749 444 -747
rect 443 -755 444 -753
rect 450 -749 451 -747
rect 450 -755 451 -753
rect 457 -749 458 -747
rect 457 -755 458 -753
rect 464 -749 465 -747
rect 464 -755 465 -753
rect 471 -749 472 -747
rect 471 -755 472 -753
rect 478 -749 479 -747
rect 478 -755 479 -753
rect 485 -749 486 -747
rect 485 -755 486 -753
rect 492 -749 493 -747
rect 492 -755 493 -753
rect 499 -749 500 -747
rect 499 -755 500 -753
rect 506 -749 507 -747
rect 506 -755 507 -753
rect 513 -749 514 -747
rect 513 -755 514 -753
rect 523 -749 524 -747
rect 520 -755 521 -753
rect 523 -755 524 -753
rect 527 -749 528 -747
rect 527 -755 528 -753
rect 530 -755 531 -753
rect 534 -749 535 -747
rect 537 -749 538 -747
rect 534 -755 535 -753
rect 537 -755 538 -753
rect 541 -749 542 -747
rect 544 -749 545 -747
rect 541 -755 542 -753
rect 544 -755 545 -753
rect 548 -749 549 -747
rect 548 -755 549 -753
rect 555 -749 556 -747
rect 555 -755 556 -753
rect 562 -749 563 -747
rect 565 -749 566 -747
rect 562 -755 563 -753
rect 569 -749 570 -747
rect 569 -755 570 -753
rect 576 -749 577 -747
rect 576 -755 577 -753
rect 583 -749 584 -747
rect 583 -755 584 -753
rect 590 -749 591 -747
rect 590 -755 591 -753
rect 600 -749 601 -747
rect 597 -755 598 -753
rect 600 -755 601 -753
rect 604 -749 605 -747
rect 604 -755 605 -753
rect 611 -749 612 -747
rect 614 -749 615 -747
rect 611 -755 612 -753
rect 614 -755 615 -753
rect 618 -749 619 -747
rect 621 -749 622 -747
rect 618 -755 619 -753
rect 628 -749 629 -747
rect 625 -755 626 -753
rect 632 -749 633 -747
rect 632 -755 633 -753
rect 639 -749 640 -747
rect 639 -755 640 -753
rect 646 -749 647 -747
rect 646 -755 647 -753
rect 653 -749 654 -747
rect 653 -755 654 -753
rect 660 -749 661 -747
rect 663 -749 664 -747
rect 660 -755 661 -753
rect 663 -755 664 -753
rect 667 -749 668 -747
rect 667 -755 668 -753
rect 674 -749 675 -747
rect 674 -755 675 -753
rect 681 -749 682 -747
rect 681 -755 682 -753
rect 688 -749 689 -747
rect 688 -755 689 -753
rect 695 -749 696 -747
rect 695 -755 696 -753
rect 702 -749 703 -747
rect 702 -755 703 -753
rect 709 -749 710 -747
rect 709 -755 710 -753
rect 716 -749 717 -747
rect 716 -755 717 -753
rect 723 -749 724 -747
rect 723 -755 724 -753
rect 730 -749 731 -747
rect 730 -755 731 -753
rect 737 -749 738 -747
rect 737 -755 738 -753
rect 744 -749 745 -747
rect 747 -749 748 -747
rect 744 -755 745 -753
rect 747 -755 748 -753
rect 751 -749 752 -747
rect 751 -755 752 -753
rect 758 -749 759 -747
rect 761 -749 762 -747
rect 758 -755 759 -753
rect 761 -755 762 -753
rect 765 -749 766 -747
rect 765 -755 766 -753
rect 772 -749 773 -747
rect 772 -755 773 -753
rect 775 -755 776 -753
rect 779 -749 780 -747
rect 779 -755 780 -753
rect 786 -749 787 -747
rect 786 -755 787 -753
rect 793 -749 794 -747
rect 793 -755 794 -753
rect 800 -749 801 -747
rect 800 -755 801 -753
rect 807 -749 808 -747
rect 807 -755 808 -753
rect 814 -749 815 -747
rect 814 -755 815 -753
rect 821 -749 822 -747
rect 821 -755 822 -753
rect 828 -749 829 -747
rect 828 -755 829 -753
rect 835 -749 836 -747
rect 835 -755 836 -753
rect 842 -749 843 -747
rect 842 -755 843 -753
rect 849 -749 850 -747
rect 849 -755 850 -753
rect 856 -749 857 -747
rect 856 -755 857 -753
rect 863 -749 864 -747
rect 863 -755 864 -753
rect 870 -749 871 -747
rect 870 -755 871 -753
rect 877 -749 878 -747
rect 877 -755 878 -753
rect 884 -749 885 -747
rect 887 -749 888 -747
rect 884 -755 885 -753
rect 887 -755 888 -753
rect 891 -749 892 -747
rect 891 -755 892 -753
rect 898 -749 899 -747
rect 898 -755 899 -753
rect 905 -749 906 -747
rect 905 -755 906 -753
rect 912 -749 913 -747
rect 912 -755 913 -753
rect 919 -749 920 -747
rect 919 -755 920 -753
rect 926 -749 927 -747
rect 926 -755 927 -753
rect 933 -749 934 -747
rect 933 -755 934 -753
rect 940 -749 941 -747
rect 943 -749 944 -747
rect 940 -755 941 -753
rect 943 -755 944 -753
rect 947 -749 948 -747
rect 947 -755 948 -753
rect 954 -749 955 -747
rect 954 -755 955 -753
rect 961 -749 962 -747
rect 961 -755 962 -753
rect 968 -749 969 -747
rect 968 -755 969 -753
rect 975 -749 976 -747
rect 975 -755 976 -753
rect 982 -749 983 -747
rect 982 -755 983 -753
rect 989 -749 990 -747
rect 989 -755 990 -753
rect 996 -749 997 -747
rect 996 -755 997 -753
rect 1003 -749 1004 -747
rect 1003 -755 1004 -753
rect 1010 -749 1011 -747
rect 1010 -755 1011 -753
rect 1017 -749 1018 -747
rect 1017 -755 1018 -753
rect 1024 -749 1025 -747
rect 1024 -755 1025 -753
rect 1031 -749 1032 -747
rect 1031 -755 1032 -753
rect 1038 -749 1039 -747
rect 1038 -755 1039 -753
rect 1045 -749 1046 -747
rect 1045 -755 1046 -753
rect 1052 -749 1053 -747
rect 1052 -755 1053 -753
rect 1059 -749 1060 -747
rect 1059 -755 1060 -753
rect 1066 -749 1067 -747
rect 1066 -755 1067 -753
rect 1073 -749 1074 -747
rect 1073 -755 1074 -753
rect 1080 -749 1081 -747
rect 1080 -755 1081 -753
rect 1087 -749 1088 -747
rect 1087 -755 1088 -753
rect 1094 -749 1095 -747
rect 1094 -755 1095 -753
rect 1101 -749 1102 -747
rect 1101 -755 1102 -753
rect 1108 -749 1109 -747
rect 1108 -755 1109 -753
rect 1115 -749 1116 -747
rect 1115 -755 1116 -753
rect 1122 -749 1123 -747
rect 1122 -755 1123 -753
rect 1129 -749 1130 -747
rect 1129 -755 1130 -753
rect 1136 -749 1137 -747
rect 1136 -755 1137 -753
rect 1143 -749 1144 -747
rect 1143 -755 1144 -753
rect 1150 -749 1151 -747
rect 1150 -755 1151 -753
rect 1157 -749 1158 -747
rect 1157 -755 1158 -753
rect 1164 -749 1165 -747
rect 1164 -755 1165 -753
rect 1171 -749 1172 -747
rect 1171 -755 1172 -753
rect 1178 -749 1179 -747
rect 1178 -755 1179 -753
rect 1185 -749 1186 -747
rect 1185 -755 1186 -753
rect 1192 -749 1193 -747
rect 1192 -755 1193 -753
rect 1199 -749 1200 -747
rect 1199 -755 1200 -753
rect 1206 -749 1207 -747
rect 1206 -755 1207 -753
rect 1213 -749 1214 -747
rect 1213 -755 1214 -753
rect 1220 -749 1221 -747
rect 1220 -755 1221 -753
rect 1227 -749 1228 -747
rect 1227 -755 1228 -753
rect 1234 -749 1235 -747
rect 1234 -755 1235 -753
rect 1241 -749 1242 -747
rect 1241 -755 1242 -753
rect 1248 -749 1249 -747
rect 1248 -755 1249 -753
rect 1255 -749 1256 -747
rect 1255 -755 1256 -753
rect 1262 -749 1263 -747
rect 1262 -755 1263 -753
rect 1269 -749 1270 -747
rect 1269 -755 1270 -753
rect 1276 -749 1277 -747
rect 1276 -755 1277 -753
rect 1283 -749 1284 -747
rect 1283 -755 1284 -753
rect 1290 -749 1291 -747
rect 1290 -755 1291 -753
rect 1297 -749 1298 -747
rect 1297 -755 1298 -753
rect 1304 -749 1305 -747
rect 1304 -755 1305 -753
rect 1311 -749 1312 -747
rect 1311 -755 1312 -753
rect 1318 -749 1319 -747
rect 1318 -755 1319 -753
rect 1325 -749 1326 -747
rect 1325 -755 1326 -753
rect 1332 -749 1333 -747
rect 1332 -755 1333 -753
rect 1339 -749 1340 -747
rect 1339 -755 1340 -753
rect 1346 -749 1347 -747
rect 1346 -755 1347 -753
rect 1353 -749 1354 -747
rect 1353 -755 1354 -753
rect 1360 -749 1361 -747
rect 1360 -755 1361 -753
rect 1367 -749 1368 -747
rect 1367 -755 1368 -753
rect 1374 -749 1375 -747
rect 1374 -755 1375 -753
rect 1381 -749 1382 -747
rect 1381 -755 1382 -753
rect 1388 -749 1389 -747
rect 1388 -755 1389 -753
rect 1395 -749 1396 -747
rect 1395 -755 1396 -753
rect 1402 -749 1403 -747
rect 1402 -755 1403 -753
rect 1409 -749 1410 -747
rect 1409 -755 1410 -753
rect 1416 -749 1417 -747
rect 1416 -755 1417 -753
rect 1423 -749 1424 -747
rect 1423 -755 1424 -753
rect 1430 -749 1431 -747
rect 1430 -755 1431 -753
rect 1437 -749 1438 -747
rect 1437 -755 1438 -753
rect 1444 -749 1445 -747
rect 1444 -755 1445 -753
rect 1451 -749 1452 -747
rect 1451 -755 1452 -753
rect 1458 -749 1459 -747
rect 1458 -755 1459 -753
rect 1465 -749 1466 -747
rect 1465 -755 1466 -753
rect 1472 -749 1473 -747
rect 1472 -755 1473 -753
rect 1479 -749 1480 -747
rect 1479 -755 1480 -753
rect 1486 -749 1487 -747
rect 1486 -755 1487 -753
rect 1493 -749 1494 -747
rect 1493 -755 1494 -753
rect 1500 -749 1501 -747
rect 1500 -755 1501 -753
rect 1507 -749 1508 -747
rect 1507 -755 1508 -753
rect 1514 -749 1515 -747
rect 1514 -755 1515 -753
rect 1521 -749 1522 -747
rect 1521 -755 1522 -753
rect 1528 -749 1529 -747
rect 1528 -755 1529 -753
rect 2 -890 3 -888
rect 2 -896 3 -894
rect 9 -890 10 -888
rect 9 -896 10 -894
rect 16 -890 17 -888
rect 16 -896 17 -894
rect 23 -890 24 -888
rect 23 -896 24 -894
rect 30 -890 31 -888
rect 30 -896 31 -894
rect 40 -890 41 -888
rect 37 -896 38 -894
rect 40 -896 41 -894
rect 44 -890 45 -888
rect 47 -890 48 -888
rect 44 -896 45 -894
rect 51 -890 52 -888
rect 51 -896 52 -894
rect 58 -890 59 -888
rect 58 -896 59 -894
rect 65 -890 66 -888
rect 65 -896 66 -894
rect 72 -890 73 -888
rect 72 -896 73 -894
rect 79 -890 80 -888
rect 79 -896 80 -894
rect 86 -890 87 -888
rect 86 -896 87 -894
rect 93 -890 94 -888
rect 93 -896 94 -894
rect 100 -890 101 -888
rect 100 -896 101 -894
rect 107 -890 108 -888
rect 107 -896 108 -894
rect 114 -890 115 -888
rect 114 -896 115 -894
rect 121 -890 122 -888
rect 121 -896 122 -894
rect 128 -890 129 -888
rect 131 -890 132 -888
rect 128 -896 129 -894
rect 131 -896 132 -894
rect 135 -890 136 -888
rect 135 -896 136 -894
rect 142 -890 143 -888
rect 142 -896 143 -894
rect 149 -890 150 -888
rect 149 -896 150 -894
rect 156 -890 157 -888
rect 156 -896 157 -894
rect 163 -890 164 -888
rect 166 -890 167 -888
rect 163 -896 164 -894
rect 170 -890 171 -888
rect 170 -896 171 -894
rect 177 -890 178 -888
rect 177 -896 178 -894
rect 184 -890 185 -888
rect 184 -896 185 -894
rect 191 -890 192 -888
rect 191 -896 192 -894
rect 198 -890 199 -888
rect 198 -896 199 -894
rect 205 -890 206 -888
rect 205 -896 206 -894
rect 212 -890 213 -888
rect 212 -896 213 -894
rect 219 -890 220 -888
rect 219 -896 220 -894
rect 226 -890 227 -888
rect 226 -896 227 -894
rect 233 -890 234 -888
rect 236 -890 237 -888
rect 233 -896 234 -894
rect 236 -896 237 -894
rect 240 -890 241 -888
rect 240 -896 241 -894
rect 247 -890 248 -888
rect 247 -896 248 -894
rect 254 -890 255 -888
rect 254 -896 255 -894
rect 261 -890 262 -888
rect 261 -896 262 -894
rect 268 -890 269 -888
rect 268 -896 269 -894
rect 275 -890 276 -888
rect 275 -896 276 -894
rect 282 -890 283 -888
rect 282 -896 283 -894
rect 289 -890 290 -888
rect 289 -896 290 -894
rect 296 -890 297 -888
rect 296 -896 297 -894
rect 303 -890 304 -888
rect 303 -896 304 -894
rect 310 -890 311 -888
rect 310 -896 311 -894
rect 317 -890 318 -888
rect 317 -896 318 -894
rect 324 -890 325 -888
rect 324 -896 325 -894
rect 331 -890 332 -888
rect 331 -896 332 -894
rect 338 -890 339 -888
rect 338 -896 339 -894
rect 345 -890 346 -888
rect 345 -896 346 -894
rect 352 -890 353 -888
rect 352 -896 353 -894
rect 359 -890 360 -888
rect 359 -896 360 -894
rect 366 -890 367 -888
rect 369 -890 370 -888
rect 366 -896 367 -894
rect 369 -896 370 -894
rect 373 -890 374 -888
rect 373 -896 374 -894
rect 380 -890 381 -888
rect 380 -896 381 -894
rect 387 -890 388 -888
rect 387 -896 388 -894
rect 394 -890 395 -888
rect 394 -896 395 -894
rect 401 -890 402 -888
rect 401 -896 402 -894
rect 408 -890 409 -888
rect 408 -896 409 -894
rect 415 -896 416 -894
rect 422 -890 423 -888
rect 422 -896 423 -894
rect 429 -890 430 -888
rect 429 -896 430 -894
rect 436 -890 437 -888
rect 439 -890 440 -888
rect 436 -896 437 -894
rect 443 -890 444 -888
rect 443 -896 444 -894
rect 450 -890 451 -888
rect 450 -896 451 -894
rect 457 -890 458 -888
rect 460 -890 461 -888
rect 457 -896 458 -894
rect 460 -896 461 -894
rect 464 -890 465 -888
rect 467 -890 468 -888
rect 464 -896 465 -894
rect 467 -896 468 -894
rect 471 -890 472 -888
rect 471 -896 472 -894
rect 478 -890 479 -888
rect 478 -896 479 -894
rect 485 -890 486 -888
rect 485 -896 486 -894
rect 492 -890 493 -888
rect 492 -896 493 -894
rect 499 -890 500 -888
rect 499 -896 500 -894
rect 506 -890 507 -888
rect 509 -890 510 -888
rect 506 -896 507 -894
rect 509 -896 510 -894
rect 513 -890 514 -888
rect 513 -896 514 -894
rect 520 -890 521 -888
rect 520 -896 521 -894
rect 527 -890 528 -888
rect 530 -890 531 -888
rect 527 -896 528 -894
rect 534 -890 535 -888
rect 537 -890 538 -888
rect 534 -896 535 -894
rect 537 -896 538 -894
rect 541 -890 542 -888
rect 541 -896 542 -894
rect 544 -896 545 -894
rect 548 -890 549 -888
rect 551 -890 552 -888
rect 548 -896 549 -894
rect 551 -896 552 -894
rect 555 -890 556 -888
rect 555 -896 556 -894
rect 562 -890 563 -888
rect 562 -896 563 -894
rect 569 -890 570 -888
rect 569 -896 570 -894
rect 576 -890 577 -888
rect 576 -896 577 -894
rect 583 -890 584 -888
rect 583 -896 584 -894
rect 590 -890 591 -888
rect 590 -896 591 -894
rect 597 -890 598 -888
rect 597 -896 598 -894
rect 604 -890 605 -888
rect 604 -896 605 -894
rect 611 -890 612 -888
rect 611 -896 612 -894
rect 618 -890 619 -888
rect 618 -896 619 -894
rect 625 -890 626 -888
rect 625 -896 626 -894
rect 632 -890 633 -888
rect 632 -896 633 -894
rect 639 -890 640 -888
rect 642 -890 643 -888
rect 639 -896 640 -894
rect 642 -896 643 -894
rect 646 -890 647 -888
rect 649 -890 650 -888
rect 646 -896 647 -894
rect 649 -896 650 -894
rect 653 -890 654 -888
rect 656 -890 657 -888
rect 653 -896 654 -894
rect 656 -896 657 -894
rect 660 -890 661 -888
rect 663 -890 664 -888
rect 660 -896 661 -894
rect 667 -890 668 -888
rect 667 -896 668 -894
rect 674 -890 675 -888
rect 674 -896 675 -894
rect 681 -890 682 -888
rect 681 -896 682 -894
rect 691 -890 692 -888
rect 688 -896 689 -894
rect 691 -896 692 -894
rect 695 -890 696 -888
rect 695 -896 696 -894
rect 702 -890 703 -888
rect 702 -896 703 -894
rect 709 -890 710 -888
rect 712 -890 713 -888
rect 709 -896 710 -894
rect 712 -896 713 -894
rect 716 -890 717 -888
rect 716 -896 717 -894
rect 723 -890 724 -888
rect 723 -896 724 -894
rect 730 -890 731 -888
rect 730 -896 731 -894
rect 737 -890 738 -888
rect 737 -896 738 -894
rect 744 -890 745 -888
rect 744 -896 745 -894
rect 751 -890 752 -888
rect 751 -896 752 -894
rect 758 -890 759 -888
rect 758 -896 759 -894
rect 765 -890 766 -888
rect 768 -890 769 -888
rect 765 -896 766 -894
rect 768 -896 769 -894
rect 772 -890 773 -888
rect 772 -896 773 -894
rect 779 -890 780 -888
rect 779 -896 780 -894
rect 786 -890 787 -888
rect 786 -896 787 -894
rect 793 -890 794 -888
rect 793 -896 794 -894
rect 800 -890 801 -888
rect 800 -896 801 -894
rect 807 -890 808 -888
rect 807 -896 808 -894
rect 810 -896 811 -894
rect 814 -890 815 -888
rect 814 -896 815 -894
rect 821 -890 822 -888
rect 821 -896 822 -894
rect 828 -890 829 -888
rect 828 -896 829 -894
rect 835 -890 836 -888
rect 838 -890 839 -888
rect 835 -896 836 -894
rect 838 -896 839 -894
rect 842 -890 843 -888
rect 842 -896 843 -894
rect 849 -890 850 -888
rect 849 -896 850 -894
rect 856 -890 857 -888
rect 856 -896 857 -894
rect 863 -890 864 -888
rect 863 -896 864 -894
rect 870 -890 871 -888
rect 870 -896 871 -894
rect 877 -890 878 -888
rect 877 -896 878 -894
rect 884 -890 885 -888
rect 884 -896 885 -894
rect 891 -890 892 -888
rect 891 -896 892 -894
rect 898 -890 899 -888
rect 898 -896 899 -894
rect 905 -890 906 -888
rect 905 -896 906 -894
rect 912 -890 913 -888
rect 912 -896 913 -894
rect 919 -890 920 -888
rect 919 -896 920 -894
rect 926 -890 927 -888
rect 926 -896 927 -894
rect 933 -890 934 -888
rect 933 -896 934 -894
rect 943 -890 944 -888
rect 943 -896 944 -894
rect 947 -890 948 -888
rect 947 -896 948 -894
rect 954 -890 955 -888
rect 954 -896 955 -894
rect 961 -890 962 -888
rect 961 -896 962 -894
rect 968 -890 969 -888
rect 968 -896 969 -894
rect 975 -890 976 -888
rect 975 -896 976 -894
rect 982 -890 983 -888
rect 989 -890 990 -888
rect 989 -896 990 -894
rect 996 -890 997 -888
rect 999 -890 1000 -888
rect 996 -896 997 -894
rect 1003 -890 1004 -888
rect 1003 -896 1004 -894
rect 1010 -890 1011 -888
rect 1010 -896 1011 -894
rect 1017 -890 1018 -888
rect 1017 -896 1018 -894
rect 1024 -890 1025 -888
rect 1024 -896 1025 -894
rect 1031 -890 1032 -888
rect 1031 -896 1032 -894
rect 1038 -890 1039 -888
rect 1038 -896 1039 -894
rect 1045 -890 1046 -888
rect 1045 -896 1046 -894
rect 1052 -890 1053 -888
rect 1052 -896 1053 -894
rect 1059 -890 1060 -888
rect 1059 -896 1060 -894
rect 1066 -890 1067 -888
rect 1066 -896 1067 -894
rect 1069 -896 1070 -894
rect 1073 -890 1074 -888
rect 1073 -896 1074 -894
rect 1080 -890 1081 -888
rect 1080 -896 1081 -894
rect 1087 -890 1088 -888
rect 1087 -896 1088 -894
rect 1094 -890 1095 -888
rect 1094 -896 1095 -894
rect 1101 -890 1102 -888
rect 1101 -896 1102 -894
rect 1108 -890 1109 -888
rect 1108 -896 1109 -894
rect 1115 -890 1116 -888
rect 1115 -896 1116 -894
rect 1122 -890 1123 -888
rect 1122 -896 1123 -894
rect 1129 -890 1130 -888
rect 1129 -896 1130 -894
rect 1136 -890 1137 -888
rect 1136 -896 1137 -894
rect 1143 -890 1144 -888
rect 1143 -896 1144 -894
rect 1150 -890 1151 -888
rect 1150 -896 1151 -894
rect 1157 -890 1158 -888
rect 1157 -896 1158 -894
rect 1164 -890 1165 -888
rect 1164 -896 1165 -894
rect 1171 -890 1172 -888
rect 1171 -896 1172 -894
rect 1178 -890 1179 -888
rect 1178 -896 1179 -894
rect 1185 -890 1186 -888
rect 1185 -896 1186 -894
rect 1192 -890 1193 -888
rect 1192 -896 1193 -894
rect 1199 -890 1200 -888
rect 1199 -896 1200 -894
rect 1206 -890 1207 -888
rect 1206 -896 1207 -894
rect 1213 -890 1214 -888
rect 1213 -896 1214 -894
rect 1220 -890 1221 -888
rect 1220 -896 1221 -894
rect 1227 -890 1228 -888
rect 1227 -896 1228 -894
rect 1234 -890 1235 -888
rect 1234 -896 1235 -894
rect 1241 -890 1242 -888
rect 1241 -896 1242 -894
rect 1248 -890 1249 -888
rect 1248 -896 1249 -894
rect 1255 -890 1256 -888
rect 1255 -896 1256 -894
rect 1262 -890 1263 -888
rect 1262 -896 1263 -894
rect 1269 -890 1270 -888
rect 1269 -896 1270 -894
rect 1276 -890 1277 -888
rect 1276 -896 1277 -894
rect 1283 -890 1284 -888
rect 1283 -896 1284 -894
rect 1290 -890 1291 -888
rect 1290 -896 1291 -894
rect 1297 -890 1298 -888
rect 1297 -896 1298 -894
rect 1304 -890 1305 -888
rect 1304 -896 1305 -894
rect 1311 -890 1312 -888
rect 1311 -896 1312 -894
rect 1318 -890 1319 -888
rect 1318 -896 1319 -894
rect 1325 -890 1326 -888
rect 1325 -896 1326 -894
rect 1332 -890 1333 -888
rect 1332 -896 1333 -894
rect 1339 -890 1340 -888
rect 1339 -896 1340 -894
rect 1346 -890 1347 -888
rect 1346 -896 1347 -894
rect 1353 -890 1354 -888
rect 1353 -896 1354 -894
rect 1360 -890 1361 -888
rect 1360 -896 1361 -894
rect 1367 -890 1368 -888
rect 1367 -896 1368 -894
rect 1374 -890 1375 -888
rect 1374 -896 1375 -894
rect 1381 -890 1382 -888
rect 1381 -896 1382 -894
rect 1388 -890 1389 -888
rect 1388 -896 1389 -894
rect 1395 -890 1396 -888
rect 1395 -896 1396 -894
rect 1402 -890 1403 -888
rect 1402 -896 1403 -894
rect 1409 -890 1410 -888
rect 1409 -896 1410 -894
rect 1416 -890 1417 -888
rect 1416 -896 1417 -894
rect 1423 -890 1424 -888
rect 1423 -896 1424 -894
rect 1430 -890 1431 -888
rect 1430 -896 1431 -894
rect 1437 -890 1438 -888
rect 1437 -896 1438 -894
rect 1444 -890 1445 -888
rect 1444 -896 1445 -894
rect 1451 -890 1452 -888
rect 1451 -896 1452 -894
rect 1458 -890 1459 -888
rect 1458 -896 1459 -894
rect 1465 -890 1466 -888
rect 1465 -896 1466 -894
rect 1472 -890 1473 -888
rect 1472 -896 1473 -894
rect 1479 -890 1480 -888
rect 1479 -896 1480 -894
rect 1486 -890 1487 -888
rect 1486 -896 1487 -894
rect 1493 -890 1494 -888
rect 1493 -896 1494 -894
rect 1500 -890 1501 -888
rect 1503 -890 1504 -888
rect 1500 -896 1501 -894
rect 1503 -896 1504 -894
rect 1514 -890 1515 -888
rect 1514 -896 1515 -894
rect 2 -1007 3 -1005
rect 2 -1013 3 -1011
rect 9 -1007 10 -1005
rect 9 -1013 10 -1011
rect 16 -1007 17 -1005
rect 16 -1013 17 -1011
rect 23 -1007 24 -1005
rect 23 -1013 24 -1011
rect 30 -1007 31 -1005
rect 30 -1013 31 -1011
rect 37 -1007 38 -1005
rect 37 -1013 38 -1011
rect 44 -1007 45 -1005
rect 44 -1013 45 -1011
rect 51 -1007 52 -1005
rect 51 -1013 52 -1011
rect 58 -1007 59 -1005
rect 58 -1013 59 -1011
rect 65 -1007 66 -1005
rect 65 -1013 66 -1011
rect 72 -1007 73 -1005
rect 72 -1013 73 -1011
rect 79 -1007 80 -1005
rect 79 -1013 80 -1011
rect 86 -1007 87 -1005
rect 86 -1013 87 -1011
rect 93 -1007 94 -1005
rect 96 -1007 97 -1005
rect 93 -1013 94 -1011
rect 96 -1013 97 -1011
rect 100 -1007 101 -1005
rect 100 -1013 101 -1011
rect 107 -1007 108 -1005
rect 107 -1013 108 -1011
rect 114 -1007 115 -1005
rect 114 -1013 115 -1011
rect 121 -1007 122 -1005
rect 121 -1013 122 -1011
rect 128 -1007 129 -1005
rect 128 -1013 129 -1011
rect 135 -1007 136 -1005
rect 135 -1013 136 -1011
rect 142 -1007 143 -1005
rect 145 -1007 146 -1005
rect 142 -1013 143 -1011
rect 145 -1013 146 -1011
rect 149 -1007 150 -1005
rect 149 -1013 150 -1011
rect 156 -1007 157 -1005
rect 156 -1013 157 -1011
rect 163 -1007 164 -1005
rect 163 -1013 164 -1011
rect 170 -1007 171 -1005
rect 170 -1013 171 -1011
rect 177 -1007 178 -1005
rect 177 -1013 178 -1011
rect 184 -1007 185 -1005
rect 184 -1013 185 -1011
rect 191 -1007 192 -1005
rect 191 -1013 192 -1011
rect 198 -1007 199 -1005
rect 198 -1013 199 -1011
rect 205 -1007 206 -1005
rect 205 -1013 206 -1011
rect 212 -1007 213 -1005
rect 212 -1013 213 -1011
rect 219 -1007 220 -1005
rect 219 -1013 220 -1011
rect 226 -1007 227 -1005
rect 226 -1013 227 -1011
rect 233 -1007 234 -1005
rect 233 -1013 234 -1011
rect 243 -1007 244 -1005
rect 240 -1013 241 -1011
rect 243 -1013 244 -1011
rect 247 -1007 248 -1005
rect 247 -1013 248 -1011
rect 254 -1007 255 -1005
rect 254 -1013 255 -1011
rect 261 -1007 262 -1005
rect 261 -1013 262 -1011
rect 268 -1007 269 -1005
rect 268 -1013 269 -1011
rect 275 -1007 276 -1005
rect 275 -1013 276 -1011
rect 282 -1007 283 -1005
rect 282 -1013 283 -1011
rect 289 -1007 290 -1005
rect 289 -1013 290 -1011
rect 296 -1007 297 -1005
rect 299 -1007 300 -1005
rect 296 -1013 297 -1011
rect 299 -1013 300 -1011
rect 303 -1007 304 -1005
rect 303 -1013 304 -1011
rect 310 -1007 311 -1005
rect 310 -1013 311 -1011
rect 317 -1007 318 -1005
rect 317 -1013 318 -1011
rect 324 -1007 325 -1005
rect 324 -1013 325 -1011
rect 334 -1007 335 -1005
rect 331 -1013 332 -1011
rect 334 -1013 335 -1011
rect 338 -1007 339 -1005
rect 338 -1013 339 -1011
rect 345 -1007 346 -1005
rect 345 -1013 346 -1011
rect 352 -1007 353 -1005
rect 352 -1013 353 -1011
rect 359 -1007 360 -1005
rect 359 -1013 360 -1011
rect 366 -1007 367 -1005
rect 366 -1013 367 -1011
rect 373 -1007 374 -1005
rect 376 -1007 377 -1005
rect 373 -1013 374 -1011
rect 376 -1013 377 -1011
rect 380 -1007 381 -1005
rect 380 -1013 381 -1011
rect 387 -1007 388 -1005
rect 387 -1013 388 -1011
rect 394 -1007 395 -1005
rect 394 -1013 395 -1011
rect 401 -1007 402 -1005
rect 401 -1013 402 -1011
rect 408 -1007 409 -1005
rect 408 -1013 409 -1011
rect 415 -1007 416 -1005
rect 415 -1013 416 -1011
rect 422 -1007 423 -1005
rect 422 -1013 423 -1011
rect 429 -1007 430 -1005
rect 429 -1013 430 -1011
rect 436 -1007 437 -1005
rect 436 -1013 437 -1011
rect 443 -1007 444 -1005
rect 443 -1013 444 -1011
rect 450 -1007 451 -1005
rect 450 -1013 451 -1011
rect 457 -1007 458 -1005
rect 457 -1013 458 -1011
rect 464 -1007 465 -1005
rect 464 -1013 465 -1011
rect 471 -1007 472 -1005
rect 471 -1013 472 -1011
rect 478 -1007 479 -1005
rect 478 -1013 479 -1011
rect 481 -1013 482 -1011
rect 485 -1007 486 -1005
rect 485 -1013 486 -1011
rect 492 -1007 493 -1005
rect 495 -1007 496 -1005
rect 492 -1013 493 -1011
rect 495 -1013 496 -1011
rect 499 -1007 500 -1005
rect 499 -1013 500 -1011
rect 506 -1007 507 -1005
rect 506 -1013 507 -1011
rect 513 -1007 514 -1005
rect 513 -1013 514 -1011
rect 520 -1007 521 -1005
rect 520 -1013 521 -1011
rect 527 -1007 528 -1005
rect 527 -1013 528 -1011
rect 534 -1007 535 -1005
rect 537 -1007 538 -1005
rect 534 -1013 535 -1011
rect 537 -1013 538 -1011
rect 541 -1007 542 -1005
rect 544 -1007 545 -1005
rect 541 -1013 542 -1011
rect 544 -1013 545 -1011
rect 548 -1007 549 -1005
rect 551 -1007 552 -1005
rect 548 -1013 549 -1011
rect 551 -1013 552 -1011
rect 555 -1007 556 -1005
rect 555 -1013 556 -1011
rect 562 -1007 563 -1005
rect 562 -1013 563 -1011
rect 569 -1007 570 -1005
rect 569 -1013 570 -1011
rect 576 -1007 577 -1005
rect 576 -1013 577 -1011
rect 583 -1007 584 -1005
rect 583 -1013 584 -1011
rect 590 -1007 591 -1005
rect 590 -1013 591 -1011
rect 597 -1007 598 -1005
rect 600 -1007 601 -1005
rect 597 -1013 598 -1011
rect 600 -1013 601 -1011
rect 604 -1007 605 -1005
rect 604 -1013 605 -1011
rect 611 -1007 612 -1005
rect 611 -1013 612 -1011
rect 618 -1007 619 -1005
rect 618 -1013 619 -1011
rect 625 -1007 626 -1005
rect 625 -1013 626 -1011
rect 632 -1007 633 -1005
rect 632 -1013 633 -1011
rect 639 -1007 640 -1005
rect 639 -1013 640 -1011
rect 646 -1007 647 -1005
rect 646 -1013 647 -1011
rect 653 -1007 654 -1005
rect 653 -1013 654 -1011
rect 660 -1007 661 -1005
rect 660 -1013 661 -1011
rect 667 -1007 668 -1005
rect 667 -1013 668 -1011
rect 674 -1007 675 -1005
rect 677 -1007 678 -1005
rect 674 -1013 675 -1011
rect 677 -1013 678 -1011
rect 681 -1007 682 -1005
rect 681 -1013 682 -1011
rect 688 -1007 689 -1005
rect 691 -1007 692 -1005
rect 691 -1013 692 -1011
rect 695 -1007 696 -1005
rect 695 -1013 696 -1011
rect 702 -1007 703 -1005
rect 705 -1007 706 -1005
rect 702 -1013 703 -1011
rect 705 -1013 706 -1011
rect 709 -1007 710 -1005
rect 709 -1013 710 -1011
rect 716 -1007 717 -1005
rect 716 -1013 717 -1011
rect 723 -1007 724 -1005
rect 723 -1013 724 -1011
rect 730 -1007 731 -1005
rect 730 -1013 731 -1011
rect 737 -1007 738 -1005
rect 737 -1013 738 -1011
rect 744 -1007 745 -1005
rect 747 -1007 748 -1005
rect 744 -1013 745 -1011
rect 747 -1013 748 -1011
rect 751 -1007 752 -1005
rect 754 -1007 755 -1005
rect 751 -1013 752 -1011
rect 754 -1013 755 -1011
rect 758 -1007 759 -1005
rect 761 -1007 762 -1005
rect 758 -1013 759 -1011
rect 761 -1013 762 -1011
rect 765 -1007 766 -1005
rect 765 -1013 766 -1011
rect 772 -1007 773 -1005
rect 772 -1013 773 -1011
rect 779 -1007 780 -1005
rect 779 -1013 780 -1011
rect 786 -1007 787 -1005
rect 786 -1013 787 -1011
rect 793 -1007 794 -1005
rect 793 -1013 794 -1011
rect 800 -1007 801 -1005
rect 800 -1013 801 -1011
rect 807 -1007 808 -1005
rect 807 -1013 808 -1011
rect 814 -1007 815 -1005
rect 814 -1013 815 -1011
rect 821 -1007 822 -1005
rect 824 -1007 825 -1005
rect 821 -1013 822 -1011
rect 824 -1013 825 -1011
rect 828 -1007 829 -1005
rect 831 -1007 832 -1005
rect 828 -1013 829 -1011
rect 831 -1013 832 -1011
rect 835 -1007 836 -1005
rect 835 -1013 836 -1011
rect 842 -1007 843 -1005
rect 842 -1013 843 -1011
rect 849 -1007 850 -1005
rect 849 -1013 850 -1011
rect 856 -1007 857 -1005
rect 859 -1007 860 -1005
rect 856 -1013 857 -1011
rect 859 -1013 860 -1011
rect 863 -1007 864 -1005
rect 863 -1013 864 -1011
rect 870 -1007 871 -1005
rect 870 -1013 871 -1011
rect 873 -1013 874 -1011
rect 877 -1007 878 -1005
rect 877 -1013 878 -1011
rect 884 -1007 885 -1005
rect 884 -1013 885 -1011
rect 891 -1007 892 -1005
rect 891 -1013 892 -1011
rect 898 -1007 899 -1005
rect 898 -1013 899 -1011
rect 905 -1007 906 -1005
rect 908 -1007 909 -1005
rect 908 -1013 909 -1011
rect 912 -1007 913 -1005
rect 912 -1013 913 -1011
rect 919 -1007 920 -1005
rect 919 -1013 920 -1011
rect 926 -1007 927 -1005
rect 926 -1013 927 -1011
rect 933 -1007 934 -1005
rect 933 -1013 934 -1011
rect 940 -1007 941 -1005
rect 940 -1013 941 -1011
rect 947 -1007 948 -1005
rect 947 -1013 948 -1011
rect 954 -1007 955 -1005
rect 954 -1013 955 -1011
rect 961 -1007 962 -1005
rect 961 -1013 962 -1011
rect 968 -1007 969 -1005
rect 968 -1013 969 -1011
rect 975 -1007 976 -1005
rect 975 -1013 976 -1011
rect 982 -1013 983 -1011
rect 992 -1007 993 -1005
rect 989 -1013 990 -1011
rect 992 -1013 993 -1011
rect 996 -1007 997 -1005
rect 996 -1013 997 -1011
rect 1003 -1007 1004 -1005
rect 1003 -1013 1004 -1011
rect 1010 -1007 1011 -1005
rect 1010 -1013 1011 -1011
rect 1017 -1007 1018 -1005
rect 1017 -1013 1018 -1011
rect 1024 -1007 1025 -1005
rect 1024 -1013 1025 -1011
rect 1031 -1007 1032 -1005
rect 1031 -1013 1032 -1011
rect 1038 -1007 1039 -1005
rect 1038 -1013 1039 -1011
rect 1045 -1007 1046 -1005
rect 1045 -1013 1046 -1011
rect 1052 -1007 1053 -1005
rect 1052 -1013 1053 -1011
rect 1059 -1007 1060 -1005
rect 1059 -1013 1060 -1011
rect 1066 -1007 1067 -1005
rect 1069 -1007 1070 -1005
rect 1066 -1013 1067 -1011
rect 1073 -1007 1074 -1005
rect 1073 -1013 1074 -1011
rect 1080 -1007 1081 -1005
rect 1080 -1013 1081 -1011
rect 1087 -1007 1088 -1005
rect 1087 -1013 1088 -1011
rect 1094 -1007 1095 -1005
rect 1094 -1013 1095 -1011
rect 1101 -1007 1102 -1005
rect 1101 -1013 1102 -1011
rect 1108 -1007 1109 -1005
rect 1108 -1013 1109 -1011
rect 1115 -1007 1116 -1005
rect 1115 -1013 1116 -1011
rect 1122 -1007 1123 -1005
rect 1122 -1013 1123 -1011
rect 1129 -1007 1130 -1005
rect 1129 -1013 1130 -1011
rect 1136 -1007 1137 -1005
rect 1136 -1013 1137 -1011
rect 1143 -1007 1144 -1005
rect 1143 -1013 1144 -1011
rect 1150 -1007 1151 -1005
rect 1150 -1013 1151 -1011
rect 1157 -1007 1158 -1005
rect 1157 -1013 1158 -1011
rect 1164 -1007 1165 -1005
rect 1164 -1013 1165 -1011
rect 1171 -1007 1172 -1005
rect 1171 -1013 1172 -1011
rect 1178 -1007 1179 -1005
rect 1178 -1013 1179 -1011
rect 1185 -1007 1186 -1005
rect 1185 -1013 1186 -1011
rect 1192 -1007 1193 -1005
rect 1192 -1013 1193 -1011
rect 1199 -1007 1200 -1005
rect 1199 -1013 1200 -1011
rect 1206 -1007 1207 -1005
rect 1206 -1013 1207 -1011
rect 1213 -1007 1214 -1005
rect 1213 -1013 1214 -1011
rect 1220 -1007 1221 -1005
rect 1220 -1013 1221 -1011
rect 1227 -1007 1228 -1005
rect 1227 -1013 1228 -1011
rect 1234 -1007 1235 -1005
rect 1234 -1013 1235 -1011
rect 1241 -1007 1242 -1005
rect 1241 -1013 1242 -1011
rect 1248 -1007 1249 -1005
rect 1248 -1013 1249 -1011
rect 1255 -1007 1256 -1005
rect 1255 -1013 1256 -1011
rect 1262 -1007 1263 -1005
rect 1262 -1013 1263 -1011
rect 1269 -1007 1270 -1005
rect 1269 -1013 1270 -1011
rect 1276 -1007 1277 -1005
rect 1276 -1013 1277 -1011
rect 1283 -1007 1284 -1005
rect 1283 -1013 1284 -1011
rect 1290 -1007 1291 -1005
rect 1290 -1013 1291 -1011
rect 1297 -1007 1298 -1005
rect 1297 -1013 1298 -1011
rect 1304 -1007 1305 -1005
rect 1304 -1013 1305 -1011
rect 1311 -1007 1312 -1005
rect 1311 -1013 1312 -1011
rect 1318 -1007 1319 -1005
rect 1318 -1013 1319 -1011
rect 1325 -1007 1326 -1005
rect 1325 -1013 1326 -1011
rect 1332 -1007 1333 -1005
rect 1332 -1013 1333 -1011
rect 1339 -1007 1340 -1005
rect 1339 -1013 1340 -1011
rect 1346 -1007 1347 -1005
rect 1346 -1013 1347 -1011
rect 1353 -1007 1354 -1005
rect 1353 -1013 1354 -1011
rect 1360 -1007 1361 -1005
rect 1360 -1013 1361 -1011
rect 1367 -1007 1368 -1005
rect 1367 -1013 1368 -1011
rect 1374 -1007 1375 -1005
rect 1374 -1013 1375 -1011
rect 1381 -1007 1382 -1005
rect 1381 -1013 1382 -1011
rect 1388 -1007 1389 -1005
rect 1388 -1013 1389 -1011
rect 1395 -1007 1396 -1005
rect 1395 -1013 1396 -1011
rect 1402 -1007 1403 -1005
rect 1402 -1013 1403 -1011
rect 1409 -1007 1410 -1005
rect 1409 -1013 1410 -1011
rect 1416 -1007 1417 -1005
rect 1416 -1013 1417 -1011
rect 1423 -1007 1424 -1005
rect 1426 -1007 1427 -1005
rect 1423 -1013 1424 -1011
rect 1426 -1013 1427 -1011
rect 1430 -1007 1431 -1005
rect 1430 -1013 1431 -1011
rect 1437 -1007 1438 -1005
rect 1437 -1013 1438 -1011
rect 1444 -1007 1445 -1005
rect 1444 -1013 1445 -1011
rect 1451 -1007 1452 -1005
rect 1451 -1013 1452 -1011
rect 1458 -1007 1459 -1005
rect 1458 -1013 1459 -1011
rect 2 -1154 3 -1152
rect 2 -1160 3 -1158
rect 9 -1154 10 -1152
rect 9 -1160 10 -1158
rect 12 -1160 13 -1158
rect 16 -1154 17 -1152
rect 16 -1160 17 -1158
rect 23 -1154 24 -1152
rect 23 -1160 24 -1158
rect 30 -1154 31 -1152
rect 33 -1154 34 -1152
rect 33 -1160 34 -1158
rect 37 -1154 38 -1152
rect 40 -1154 41 -1152
rect 37 -1160 38 -1158
rect 40 -1160 41 -1158
rect 44 -1154 45 -1152
rect 44 -1160 45 -1158
rect 51 -1154 52 -1152
rect 51 -1160 52 -1158
rect 58 -1154 59 -1152
rect 58 -1160 59 -1158
rect 65 -1154 66 -1152
rect 65 -1160 66 -1158
rect 72 -1154 73 -1152
rect 72 -1160 73 -1158
rect 79 -1154 80 -1152
rect 82 -1154 83 -1152
rect 79 -1160 80 -1158
rect 82 -1160 83 -1158
rect 86 -1154 87 -1152
rect 86 -1160 87 -1158
rect 93 -1154 94 -1152
rect 93 -1160 94 -1158
rect 100 -1154 101 -1152
rect 100 -1160 101 -1158
rect 107 -1154 108 -1152
rect 107 -1160 108 -1158
rect 114 -1154 115 -1152
rect 114 -1160 115 -1158
rect 121 -1154 122 -1152
rect 121 -1160 122 -1158
rect 128 -1154 129 -1152
rect 128 -1160 129 -1158
rect 135 -1154 136 -1152
rect 135 -1160 136 -1158
rect 142 -1154 143 -1152
rect 142 -1160 143 -1158
rect 149 -1154 150 -1152
rect 149 -1160 150 -1158
rect 156 -1154 157 -1152
rect 156 -1160 157 -1158
rect 166 -1154 167 -1152
rect 163 -1160 164 -1158
rect 166 -1160 167 -1158
rect 170 -1154 171 -1152
rect 170 -1160 171 -1158
rect 177 -1154 178 -1152
rect 177 -1160 178 -1158
rect 184 -1154 185 -1152
rect 184 -1160 185 -1158
rect 191 -1154 192 -1152
rect 191 -1160 192 -1158
rect 198 -1154 199 -1152
rect 201 -1154 202 -1152
rect 198 -1160 199 -1158
rect 205 -1154 206 -1152
rect 205 -1160 206 -1158
rect 212 -1154 213 -1152
rect 212 -1160 213 -1158
rect 219 -1154 220 -1152
rect 219 -1160 220 -1158
rect 226 -1154 227 -1152
rect 226 -1160 227 -1158
rect 233 -1154 234 -1152
rect 233 -1160 234 -1158
rect 240 -1154 241 -1152
rect 240 -1160 241 -1158
rect 247 -1154 248 -1152
rect 247 -1160 248 -1158
rect 254 -1154 255 -1152
rect 254 -1160 255 -1158
rect 261 -1154 262 -1152
rect 261 -1160 262 -1158
rect 268 -1154 269 -1152
rect 268 -1160 269 -1158
rect 275 -1154 276 -1152
rect 275 -1160 276 -1158
rect 282 -1154 283 -1152
rect 282 -1160 283 -1158
rect 289 -1154 290 -1152
rect 289 -1160 290 -1158
rect 296 -1154 297 -1152
rect 296 -1160 297 -1158
rect 303 -1154 304 -1152
rect 303 -1160 304 -1158
rect 310 -1154 311 -1152
rect 310 -1160 311 -1158
rect 317 -1154 318 -1152
rect 317 -1160 318 -1158
rect 324 -1154 325 -1152
rect 324 -1160 325 -1158
rect 331 -1154 332 -1152
rect 331 -1160 332 -1158
rect 338 -1154 339 -1152
rect 338 -1160 339 -1158
rect 345 -1154 346 -1152
rect 345 -1160 346 -1158
rect 352 -1154 353 -1152
rect 355 -1154 356 -1152
rect 352 -1160 353 -1158
rect 355 -1160 356 -1158
rect 359 -1154 360 -1152
rect 359 -1160 360 -1158
rect 366 -1154 367 -1152
rect 366 -1160 367 -1158
rect 373 -1154 374 -1152
rect 373 -1160 374 -1158
rect 380 -1154 381 -1152
rect 380 -1160 381 -1158
rect 387 -1154 388 -1152
rect 390 -1154 391 -1152
rect 387 -1160 388 -1158
rect 390 -1160 391 -1158
rect 394 -1154 395 -1152
rect 394 -1160 395 -1158
rect 401 -1154 402 -1152
rect 401 -1160 402 -1158
rect 408 -1154 409 -1152
rect 408 -1160 409 -1158
rect 415 -1154 416 -1152
rect 415 -1160 416 -1158
rect 422 -1154 423 -1152
rect 422 -1160 423 -1158
rect 432 -1154 433 -1152
rect 429 -1160 430 -1158
rect 436 -1154 437 -1152
rect 436 -1160 437 -1158
rect 443 -1154 444 -1152
rect 446 -1154 447 -1152
rect 443 -1160 444 -1158
rect 446 -1160 447 -1158
rect 450 -1154 451 -1152
rect 450 -1160 451 -1158
rect 457 -1154 458 -1152
rect 460 -1154 461 -1152
rect 457 -1160 458 -1158
rect 460 -1160 461 -1158
rect 464 -1154 465 -1152
rect 464 -1160 465 -1158
rect 471 -1154 472 -1152
rect 471 -1160 472 -1158
rect 478 -1154 479 -1152
rect 478 -1160 479 -1158
rect 485 -1154 486 -1152
rect 485 -1160 486 -1158
rect 492 -1154 493 -1152
rect 492 -1160 493 -1158
rect 499 -1154 500 -1152
rect 499 -1160 500 -1158
rect 506 -1154 507 -1152
rect 506 -1160 507 -1158
rect 513 -1154 514 -1152
rect 513 -1160 514 -1158
rect 520 -1154 521 -1152
rect 520 -1160 521 -1158
rect 527 -1154 528 -1152
rect 527 -1160 528 -1158
rect 534 -1154 535 -1152
rect 534 -1160 535 -1158
rect 541 -1154 542 -1152
rect 541 -1160 542 -1158
rect 548 -1154 549 -1152
rect 548 -1160 549 -1158
rect 555 -1154 556 -1152
rect 555 -1160 556 -1158
rect 562 -1154 563 -1152
rect 562 -1160 563 -1158
rect 569 -1154 570 -1152
rect 569 -1160 570 -1158
rect 576 -1154 577 -1152
rect 576 -1160 577 -1158
rect 583 -1154 584 -1152
rect 583 -1160 584 -1158
rect 590 -1154 591 -1152
rect 593 -1154 594 -1152
rect 590 -1160 591 -1158
rect 593 -1160 594 -1158
rect 597 -1154 598 -1152
rect 597 -1160 598 -1158
rect 604 -1154 605 -1152
rect 607 -1154 608 -1152
rect 604 -1160 605 -1158
rect 611 -1154 612 -1152
rect 611 -1160 612 -1158
rect 618 -1154 619 -1152
rect 618 -1160 619 -1158
rect 625 -1154 626 -1152
rect 628 -1154 629 -1152
rect 625 -1160 626 -1158
rect 628 -1160 629 -1158
rect 632 -1154 633 -1152
rect 632 -1160 633 -1158
rect 639 -1154 640 -1152
rect 639 -1160 640 -1158
rect 646 -1154 647 -1152
rect 646 -1160 647 -1158
rect 653 -1154 654 -1152
rect 653 -1160 654 -1158
rect 660 -1154 661 -1152
rect 663 -1154 664 -1152
rect 660 -1160 661 -1158
rect 663 -1160 664 -1158
rect 667 -1154 668 -1152
rect 670 -1154 671 -1152
rect 667 -1160 668 -1158
rect 670 -1160 671 -1158
rect 674 -1154 675 -1152
rect 674 -1160 675 -1158
rect 681 -1154 682 -1152
rect 681 -1160 682 -1158
rect 688 -1154 689 -1152
rect 688 -1160 689 -1158
rect 695 -1154 696 -1152
rect 695 -1160 696 -1158
rect 702 -1154 703 -1152
rect 702 -1160 703 -1158
rect 709 -1154 710 -1152
rect 709 -1160 710 -1158
rect 716 -1154 717 -1152
rect 719 -1154 720 -1152
rect 716 -1160 717 -1158
rect 719 -1160 720 -1158
rect 723 -1154 724 -1152
rect 723 -1160 724 -1158
rect 730 -1154 731 -1152
rect 733 -1154 734 -1152
rect 730 -1160 731 -1158
rect 733 -1160 734 -1158
rect 737 -1154 738 -1152
rect 737 -1160 738 -1158
rect 744 -1154 745 -1152
rect 744 -1160 745 -1158
rect 751 -1154 752 -1152
rect 754 -1154 755 -1152
rect 751 -1160 752 -1158
rect 754 -1160 755 -1158
rect 758 -1154 759 -1152
rect 758 -1160 759 -1158
rect 765 -1154 766 -1152
rect 765 -1160 766 -1158
rect 772 -1154 773 -1152
rect 772 -1160 773 -1158
rect 779 -1154 780 -1152
rect 779 -1160 780 -1158
rect 786 -1154 787 -1152
rect 786 -1160 787 -1158
rect 793 -1154 794 -1152
rect 796 -1154 797 -1152
rect 793 -1160 794 -1158
rect 796 -1160 797 -1158
rect 800 -1154 801 -1152
rect 800 -1160 801 -1158
rect 807 -1154 808 -1152
rect 807 -1160 808 -1158
rect 814 -1154 815 -1152
rect 814 -1160 815 -1158
rect 821 -1154 822 -1152
rect 821 -1160 822 -1158
rect 828 -1154 829 -1152
rect 831 -1154 832 -1152
rect 828 -1160 829 -1158
rect 831 -1160 832 -1158
rect 835 -1154 836 -1152
rect 835 -1160 836 -1158
rect 842 -1154 843 -1152
rect 842 -1160 843 -1158
rect 849 -1154 850 -1152
rect 849 -1160 850 -1158
rect 856 -1154 857 -1152
rect 859 -1154 860 -1152
rect 856 -1160 857 -1158
rect 859 -1160 860 -1158
rect 863 -1154 864 -1152
rect 863 -1160 864 -1158
rect 870 -1154 871 -1152
rect 870 -1160 871 -1158
rect 877 -1154 878 -1152
rect 877 -1160 878 -1158
rect 884 -1154 885 -1152
rect 884 -1160 885 -1158
rect 894 -1154 895 -1152
rect 891 -1160 892 -1158
rect 894 -1160 895 -1158
rect 898 -1154 899 -1152
rect 898 -1160 899 -1158
rect 905 -1154 906 -1152
rect 905 -1160 906 -1158
rect 912 -1154 913 -1152
rect 912 -1160 913 -1158
rect 919 -1154 920 -1152
rect 919 -1160 920 -1158
rect 926 -1154 927 -1152
rect 926 -1160 927 -1158
rect 933 -1154 934 -1152
rect 936 -1154 937 -1152
rect 933 -1160 934 -1158
rect 936 -1160 937 -1158
rect 940 -1154 941 -1152
rect 940 -1160 941 -1158
rect 947 -1154 948 -1152
rect 947 -1160 948 -1158
rect 954 -1154 955 -1152
rect 957 -1154 958 -1152
rect 954 -1160 955 -1158
rect 957 -1160 958 -1158
rect 961 -1154 962 -1152
rect 961 -1160 962 -1158
rect 968 -1154 969 -1152
rect 968 -1160 969 -1158
rect 975 -1154 976 -1152
rect 975 -1160 976 -1158
rect 982 -1154 983 -1152
rect 982 -1160 983 -1158
rect 989 -1154 990 -1152
rect 989 -1160 990 -1158
rect 996 -1154 997 -1152
rect 996 -1160 997 -1158
rect 1003 -1154 1004 -1152
rect 1003 -1160 1004 -1158
rect 1010 -1154 1011 -1152
rect 1010 -1160 1011 -1158
rect 1017 -1154 1018 -1152
rect 1017 -1160 1018 -1158
rect 1024 -1154 1025 -1152
rect 1024 -1160 1025 -1158
rect 1031 -1154 1032 -1152
rect 1038 -1154 1039 -1152
rect 1038 -1160 1039 -1158
rect 1045 -1154 1046 -1152
rect 1045 -1160 1046 -1158
rect 1052 -1154 1053 -1152
rect 1052 -1160 1053 -1158
rect 1059 -1154 1060 -1152
rect 1059 -1160 1060 -1158
rect 1066 -1154 1067 -1152
rect 1066 -1160 1067 -1158
rect 1073 -1154 1074 -1152
rect 1073 -1160 1074 -1158
rect 1080 -1154 1081 -1152
rect 1080 -1160 1081 -1158
rect 1087 -1154 1088 -1152
rect 1087 -1160 1088 -1158
rect 1094 -1154 1095 -1152
rect 1094 -1160 1095 -1158
rect 1101 -1154 1102 -1152
rect 1101 -1160 1102 -1158
rect 1108 -1154 1109 -1152
rect 1108 -1160 1109 -1158
rect 1115 -1154 1116 -1152
rect 1115 -1160 1116 -1158
rect 1122 -1154 1123 -1152
rect 1122 -1160 1123 -1158
rect 1129 -1154 1130 -1152
rect 1129 -1160 1130 -1158
rect 1136 -1154 1137 -1152
rect 1136 -1160 1137 -1158
rect 1143 -1154 1144 -1152
rect 1143 -1160 1144 -1158
rect 1150 -1154 1151 -1152
rect 1150 -1160 1151 -1158
rect 1157 -1154 1158 -1152
rect 1157 -1160 1158 -1158
rect 1164 -1154 1165 -1152
rect 1164 -1160 1165 -1158
rect 1171 -1154 1172 -1152
rect 1171 -1160 1172 -1158
rect 1178 -1154 1179 -1152
rect 1178 -1160 1179 -1158
rect 1185 -1154 1186 -1152
rect 1185 -1160 1186 -1158
rect 1192 -1154 1193 -1152
rect 1192 -1160 1193 -1158
rect 1199 -1154 1200 -1152
rect 1199 -1160 1200 -1158
rect 1206 -1154 1207 -1152
rect 1206 -1160 1207 -1158
rect 1213 -1154 1214 -1152
rect 1213 -1160 1214 -1158
rect 1220 -1154 1221 -1152
rect 1220 -1160 1221 -1158
rect 1227 -1154 1228 -1152
rect 1227 -1160 1228 -1158
rect 1234 -1154 1235 -1152
rect 1234 -1160 1235 -1158
rect 1241 -1154 1242 -1152
rect 1241 -1160 1242 -1158
rect 1248 -1154 1249 -1152
rect 1248 -1160 1249 -1158
rect 1251 -1160 1252 -1158
rect 1255 -1154 1256 -1152
rect 1255 -1160 1256 -1158
rect 1262 -1154 1263 -1152
rect 1262 -1160 1263 -1158
rect 1269 -1154 1270 -1152
rect 1269 -1160 1270 -1158
rect 1276 -1154 1277 -1152
rect 1276 -1160 1277 -1158
rect 1283 -1154 1284 -1152
rect 1283 -1160 1284 -1158
rect 1290 -1154 1291 -1152
rect 1290 -1160 1291 -1158
rect 1297 -1154 1298 -1152
rect 1297 -1160 1298 -1158
rect 1304 -1154 1305 -1152
rect 1304 -1160 1305 -1158
rect 1311 -1154 1312 -1152
rect 1311 -1160 1312 -1158
rect 1318 -1154 1319 -1152
rect 1318 -1160 1319 -1158
rect 1325 -1154 1326 -1152
rect 1325 -1160 1326 -1158
rect 1332 -1154 1333 -1152
rect 1332 -1160 1333 -1158
rect 1339 -1154 1340 -1152
rect 1339 -1160 1340 -1158
rect 1346 -1154 1347 -1152
rect 1346 -1160 1347 -1158
rect 1353 -1154 1354 -1152
rect 1353 -1160 1354 -1158
rect 1360 -1154 1361 -1152
rect 1360 -1160 1361 -1158
rect 1367 -1154 1368 -1152
rect 1367 -1160 1368 -1158
rect 1374 -1154 1375 -1152
rect 1374 -1160 1375 -1158
rect 1381 -1154 1382 -1152
rect 1381 -1160 1382 -1158
rect 1388 -1154 1389 -1152
rect 1388 -1160 1389 -1158
rect 1395 -1154 1396 -1152
rect 1395 -1160 1396 -1158
rect 1402 -1154 1403 -1152
rect 1402 -1160 1403 -1158
rect 1409 -1154 1410 -1152
rect 1409 -1160 1410 -1158
rect 1416 -1154 1417 -1152
rect 1416 -1160 1417 -1158
rect 1423 -1154 1424 -1152
rect 1423 -1160 1424 -1158
rect 1430 -1154 1431 -1152
rect 1430 -1160 1431 -1158
rect 1437 -1154 1438 -1152
rect 1437 -1160 1438 -1158
rect 1444 -1154 1445 -1152
rect 1444 -1160 1445 -1158
rect 1451 -1154 1452 -1152
rect 1451 -1160 1452 -1158
rect 1458 -1154 1459 -1152
rect 1458 -1160 1459 -1158
rect 1465 -1154 1466 -1152
rect 1465 -1160 1466 -1158
rect 1472 -1154 1473 -1152
rect 1472 -1160 1473 -1158
rect 1479 -1154 1480 -1152
rect 1479 -1160 1480 -1158
rect 1486 -1154 1487 -1152
rect 1486 -1160 1487 -1158
rect 1493 -1154 1494 -1152
rect 1493 -1160 1494 -1158
rect 1500 -1154 1501 -1152
rect 1500 -1160 1501 -1158
rect 1507 -1154 1508 -1152
rect 1507 -1160 1508 -1158
rect 1514 -1154 1515 -1152
rect 1514 -1160 1515 -1158
rect 1521 -1154 1522 -1152
rect 1521 -1160 1522 -1158
rect 1528 -1154 1529 -1152
rect 1528 -1160 1529 -1158
rect 1535 -1154 1536 -1152
rect 1535 -1160 1536 -1158
rect 1542 -1154 1543 -1152
rect 1542 -1160 1543 -1158
rect 1549 -1154 1550 -1152
rect 1549 -1160 1550 -1158
rect 1556 -1154 1557 -1152
rect 1556 -1160 1557 -1158
rect 1563 -1154 1564 -1152
rect 1563 -1160 1564 -1158
rect 1570 -1154 1571 -1152
rect 1570 -1160 1571 -1158
rect 1577 -1154 1578 -1152
rect 1577 -1160 1578 -1158
rect 1584 -1154 1585 -1152
rect 1584 -1160 1585 -1158
rect 1591 -1154 1592 -1152
rect 1591 -1160 1592 -1158
rect 1598 -1154 1599 -1152
rect 1598 -1160 1599 -1158
rect 2 -1279 3 -1277
rect 2 -1285 3 -1283
rect 9 -1279 10 -1277
rect 9 -1285 10 -1283
rect 16 -1279 17 -1277
rect 16 -1285 17 -1283
rect 23 -1279 24 -1277
rect 23 -1285 24 -1283
rect 30 -1279 31 -1277
rect 30 -1285 31 -1283
rect 37 -1279 38 -1277
rect 37 -1285 38 -1283
rect 44 -1279 45 -1277
rect 44 -1285 45 -1283
rect 51 -1279 52 -1277
rect 51 -1285 52 -1283
rect 58 -1279 59 -1277
rect 61 -1279 62 -1277
rect 58 -1285 59 -1283
rect 61 -1285 62 -1283
rect 65 -1279 66 -1277
rect 65 -1285 66 -1283
rect 72 -1279 73 -1277
rect 72 -1285 73 -1283
rect 79 -1279 80 -1277
rect 79 -1285 80 -1283
rect 86 -1279 87 -1277
rect 86 -1285 87 -1283
rect 93 -1279 94 -1277
rect 93 -1285 94 -1283
rect 100 -1279 101 -1277
rect 103 -1279 104 -1277
rect 100 -1285 101 -1283
rect 103 -1285 104 -1283
rect 107 -1279 108 -1277
rect 107 -1285 108 -1283
rect 114 -1279 115 -1277
rect 114 -1285 115 -1283
rect 121 -1279 122 -1277
rect 121 -1285 122 -1283
rect 128 -1279 129 -1277
rect 131 -1279 132 -1277
rect 128 -1285 129 -1283
rect 131 -1285 132 -1283
rect 135 -1279 136 -1277
rect 135 -1285 136 -1283
rect 142 -1279 143 -1277
rect 142 -1285 143 -1283
rect 149 -1279 150 -1277
rect 149 -1285 150 -1283
rect 156 -1279 157 -1277
rect 156 -1285 157 -1283
rect 163 -1279 164 -1277
rect 163 -1285 164 -1283
rect 170 -1279 171 -1277
rect 173 -1279 174 -1277
rect 170 -1285 171 -1283
rect 177 -1279 178 -1277
rect 177 -1285 178 -1283
rect 184 -1279 185 -1277
rect 184 -1285 185 -1283
rect 191 -1279 192 -1277
rect 191 -1285 192 -1283
rect 198 -1279 199 -1277
rect 198 -1285 199 -1283
rect 205 -1279 206 -1277
rect 205 -1285 206 -1283
rect 212 -1279 213 -1277
rect 212 -1285 213 -1283
rect 219 -1279 220 -1277
rect 219 -1285 220 -1283
rect 226 -1279 227 -1277
rect 226 -1285 227 -1283
rect 233 -1279 234 -1277
rect 233 -1285 234 -1283
rect 240 -1279 241 -1277
rect 240 -1285 241 -1283
rect 247 -1279 248 -1277
rect 247 -1285 248 -1283
rect 254 -1279 255 -1277
rect 254 -1285 255 -1283
rect 261 -1279 262 -1277
rect 261 -1285 262 -1283
rect 268 -1279 269 -1277
rect 268 -1285 269 -1283
rect 275 -1279 276 -1277
rect 275 -1285 276 -1283
rect 282 -1279 283 -1277
rect 282 -1285 283 -1283
rect 289 -1279 290 -1277
rect 289 -1285 290 -1283
rect 296 -1279 297 -1277
rect 296 -1285 297 -1283
rect 303 -1279 304 -1277
rect 303 -1285 304 -1283
rect 310 -1279 311 -1277
rect 310 -1285 311 -1283
rect 317 -1279 318 -1277
rect 320 -1279 321 -1277
rect 317 -1285 318 -1283
rect 320 -1285 321 -1283
rect 324 -1279 325 -1277
rect 324 -1285 325 -1283
rect 331 -1279 332 -1277
rect 331 -1285 332 -1283
rect 338 -1279 339 -1277
rect 341 -1279 342 -1277
rect 345 -1279 346 -1277
rect 345 -1285 346 -1283
rect 352 -1279 353 -1277
rect 352 -1285 353 -1283
rect 359 -1279 360 -1277
rect 362 -1279 363 -1277
rect 359 -1285 360 -1283
rect 362 -1285 363 -1283
rect 366 -1279 367 -1277
rect 366 -1285 367 -1283
rect 373 -1279 374 -1277
rect 373 -1285 374 -1283
rect 380 -1279 381 -1277
rect 380 -1285 381 -1283
rect 387 -1279 388 -1277
rect 387 -1285 388 -1283
rect 394 -1279 395 -1277
rect 394 -1285 395 -1283
rect 401 -1279 402 -1277
rect 401 -1285 402 -1283
rect 408 -1279 409 -1277
rect 408 -1285 409 -1283
rect 415 -1279 416 -1277
rect 415 -1285 416 -1283
rect 422 -1279 423 -1277
rect 422 -1285 423 -1283
rect 429 -1279 430 -1277
rect 429 -1285 430 -1283
rect 436 -1279 437 -1277
rect 436 -1285 437 -1283
rect 443 -1279 444 -1277
rect 443 -1285 444 -1283
rect 450 -1279 451 -1277
rect 450 -1285 451 -1283
rect 457 -1279 458 -1277
rect 457 -1285 458 -1283
rect 464 -1279 465 -1277
rect 464 -1285 465 -1283
rect 471 -1279 472 -1277
rect 471 -1285 472 -1283
rect 478 -1279 479 -1277
rect 481 -1279 482 -1277
rect 478 -1285 479 -1283
rect 481 -1285 482 -1283
rect 485 -1279 486 -1277
rect 485 -1285 486 -1283
rect 492 -1279 493 -1277
rect 492 -1285 493 -1283
rect 499 -1279 500 -1277
rect 499 -1285 500 -1283
rect 506 -1279 507 -1277
rect 509 -1279 510 -1277
rect 506 -1285 507 -1283
rect 509 -1285 510 -1283
rect 513 -1279 514 -1277
rect 513 -1285 514 -1283
rect 520 -1279 521 -1277
rect 520 -1285 521 -1283
rect 523 -1285 524 -1283
rect 527 -1279 528 -1277
rect 530 -1279 531 -1277
rect 527 -1285 528 -1283
rect 530 -1285 531 -1283
rect 534 -1279 535 -1277
rect 534 -1285 535 -1283
rect 541 -1279 542 -1277
rect 541 -1285 542 -1283
rect 548 -1279 549 -1277
rect 548 -1285 549 -1283
rect 551 -1285 552 -1283
rect 555 -1279 556 -1277
rect 558 -1279 559 -1277
rect 555 -1285 556 -1283
rect 558 -1285 559 -1283
rect 562 -1279 563 -1277
rect 562 -1285 563 -1283
rect 569 -1279 570 -1277
rect 569 -1285 570 -1283
rect 576 -1279 577 -1277
rect 576 -1285 577 -1283
rect 583 -1279 584 -1277
rect 583 -1285 584 -1283
rect 590 -1279 591 -1277
rect 590 -1285 591 -1283
rect 597 -1279 598 -1277
rect 597 -1285 598 -1283
rect 604 -1279 605 -1277
rect 607 -1279 608 -1277
rect 604 -1285 605 -1283
rect 607 -1285 608 -1283
rect 611 -1279 612 -1277
rect 611 -1285 612 -1283
rect 618 -1279 619 -1277
rect 618 -1285 619 -1283
rect 625 -1279 626 -1277
rect 625 -1285 626 -1283
rect 632 -1279 633 -1277
rect 632 -1285 633 -1283
rect 639 -1279 640 -1277
rect 639 -1285 640 -1283
rect 646 -1279 647 -1277
rect 646 -1285 647 -1283
rect 653 -1279 654 -1277
rect 653 -1285 654 -1283
rect 660 -1279 661 -1277
rect 660 -1285 661 -1283
rect 667 -1279 668 -1277
rect 667 -1285 668 -1283
rect 674 -1279 675 -1277
rect 674 -1285 675 -1283
rect 681 -1279 682 -1277
rect 681 -1285 682 -1283
rect 688 -1279 689 -1277
rect 688 -1285 689 -1283
rect 695 -1279 696 -1277
rect 695 -1285 696 -1283
rect 702 -1279 703 -1277
rect 702 -1285 703 -1283
rect 709 -1279 710 -1277
rect 709 -1285 710 -1283
rect 716 -1279 717 -1277
rect 719 -1279 720 -1277
rect 716 -1285 717 -1283
rect 719 -1285 720 -1283
rect 723 -1279 724 -1277
rect 726 -1279 727 -1277
rect 723 -1285 724 -1283
rect 726 -1285 727 -1283
rect 730 -1279 731 -1277
rect 730 -1285 731 -1283
rect 737 -1279 738 -1277
rect 737 -1285 738 -1283
rect 744 -1279 745 -1277
rect 744 -1285 745 -1283
rect 751 -1279 752 -1277
rect 754 -1279 755 -1277
rect 751 -1285 752 -1283
rect 754 -1285 755 -1283
rect 758 -1279 759 -1277
rect 758 -1285 759 -1283
rect 765 -1279 766 -1277
rect 768 -1279 769 -1277
rect 765 -1285 766 -1283
rect 768 -1285 769 -1283
rect 772 -1279 773 -1277
rect 772 -1285 773 -1283
rect 779 -1279 780 -1277
rect 782 -1279 783 -1277
rect 779 -1285 780 -1283
rect 782 -1285 783 -1283
rect 786 -1279 787 -1277
rect 786 -1285 787 -1283
rect 793 -1279 794 -1277
rect 793 -1285 794 -1283
rect 800 -1279 801 -1277
rect 800 -1285 801 -1283
rect 807 -1279 808 -1277
rect 807 -1285 808 -1283
rect 814 -1279 815 -1277
rect 814 -1285 815 -1283
rect 821 -1279 822 -1277
rect 821 -1285 822 -1283
rect 828 -1279 829 -1277
rect 828 -1285 829 -1283
rect 835 -1279 836 -1277
rect 838 -1279 839 -1277
rect 835 -1285 836 -1283
rect 838 -1285 839 -1283
rect 842 -1279 843 -1277
rect 842 -1285 843 -1283
rect 849 -1279 850 -1277
rect 849 -1285 850 -1283
rect 856 -1279 857 -1277
rect 859 -1279 860 -1277
rect 856 -1285 857 -1283
rect 859 -1285 860 -1283
rect 863 -1279 864 -1277
rect 863 -1285 864 -1283
rect 870 -1279 871 -1277
rect 870 -1285 871 -1283
rect 877 -1279 878 -1277
rect 877 -1285 878 -1283
rect 884 -1279 885 -1277
rect 884 -1285 885 -1283
rect 891 -1279 892 -1277
rect 891 -1285 892 -1283
rect 898 -1279 899 -1277
rect 898 -1285 899 -1283
rect 905 -1279 906 -1277
rect 905 -1285 906 -1283
rect 912 -1279 913 -1277
rect 912 -1285 913 -1283
rect 919 -1279 920 -1277
rect 922 -1279 923 -1277
rect 922 -1285 923 -1283
rect 926 -1279 927 -1277
rect 926 -1285 927 -1283
rect 933 -1279 934 -1277
rect 936 -1279 937 -1277
rect 933 -1285 934 -1283
rect 940 -1279 941 -1277
rect 940 -1285 941 -1283
rect 947 -1279 948 -1277
rect 947 -1285 948 -1283
rect 954 -1279 955 -1277
rect 954 -1285 955 -1283
rect 961 -1279 962 -1277
rect 961 -1285 962 -1283
rect 968 -1279 969 -1277
rect 968 -1285 969 -1283
rect 975 -1279 976 -1277
rect 975 -1285 976 -1283
rect 982 -1279 983 -1277
rect 982 -1285 983 -1283
rect 989 -1279 990 -1277
rect 989 -1285 990 -1283
rect 996 -1279 997 -1277
rect 996 -1285 997 -1283
rect 1003 -1279 1004 -1277
rect 1003 -1285 1004 -1283
rect 1010 -1279 1011 -1277
rect 1010 -1285 1011 -1283
rect 1017 -1279 1018 -1277
rect 1017 -1285 1018 -1283
rect 1024 -1279 1025 -1277
rect 1024 -1285 1025 -1283
rect 1031 -1285 1032 -1283
rect 1038 -1279 1039 -1277
rect 1038 -1285 1039 -1283
rect 1045 -1279 1046 -1277
rect 1045 -1285 1046 -1283
rect 1052 -1279 1053 -1277
rect 1055 -1279 1056 -1277
rect 1052 -1285 1053 -1283
rect 1055 -1285 1056 -1283
rect 1059 -1279 1060 -1277
rect 1059 -1285 1060 -1283
rect 1066 -1279 1067 -1277
rect 1066 -1285 1067 -1283
rect 1073 -1279 1074 -1277
rect 1073 -1285 1074 -1283
rect 1080 -1279 1081 -1277
rect 1080 -1285 1081 -1283
rect 1087 -1279 1088 -1277
rect 1087 -1285 1088 -1283
rect 1094 -1279 1095 -1277
rect 1094 -1285 1095 -1283
rect 1101 -1279 1102 -1277
rect 1101 -1285 1102 -1283
rect 1108 -1279 1109 -1277
rect 1108 -1285 1109 -1283
rect 1115 -1279 1116 -1277
rect 1115 -1285 1116 -1283
rect 1122 -1279 1123 -1277
rect 1122 -1285 1123 -1283
rect 1129 -1279 1130 -1277
rect 1129 -1285 1130 -1283
rect 1136 -1279 1137 -1277
rect 1136 -1285 1137 -1283
rect 1143 -1279 1144 -1277
rect 1143 -1285 1144 -1283
rect 1150 -1279 1151 -1277
rect 1150 -1285 1151 -1283
rect 1157 -1279 1158 -1277
rect 1157 -1285 1158 -1283
rect 1164 -1279 1165 -1277
rect 1164 -1285 1165 -1283
rect 1174 -1279 1175 -1277
rect 1171 -1285 1172 -1283
rect 1178 -1279 1179 -1277
rect 1178 -1285 1179 -1283
rect 1185 -1279 1186 -1277
rect 1185 -1285 1186 -1283
rect 1192 -1279 1193 -1277
rect 1192 -1285 1193 -1283
rect 1199 -1279 1200 -1277
rect 1199 -1285 1200 -1283
rect 1206 -1279 1207 -1277
rect 1206 -1285 1207 -1283
rect 1213 -1279 1214 -1277
rect 1213 -1285 1214 -1283
rect 1220 -1279 1221 -1277
rect 1220 -1285 1221 -1283
rect 1227 -1279 1228 -1277
rect 1227 -1285 1228 -1283
rect 1234 -1279 1235 -1277
rect 1234 -1285 1235 -1283
rect 1241 -1279 1242 -1277
rect 1241 -1285 1242 -1283
rect 1248 -1279 1249 -1277
rect 1251 -1279 1252 -1277
rect 1248 -1285 1249 -1283
rect 1255 -1279 1256 -1277
rect 1255 -1285 1256 -1283
rect 1262 -1279 1263 -1277
rect 1262 -1285 1263 -1283
rect 1269 -1279 1270 -1277
rect 1269 -1285 1270 -1283
rect 1276 -1279 1277 -1277
rect 1276 -1285 1277 -1283
rect 1283 -1279 1284 -1277
rect 1283 -1285 1284 -1283
rect 1290 -1279 1291 -1277
rect 1290 -1285 1291 -1283
rect 1297 -1279 1298 -1277
rect 1297 -1285 1298 -1283
rect 1304 -1279 1305 -1277
rect 1304 -1285 1305 -1283
rect 1311 -1279 1312 -1277
rect 1311 -1285 1312 -1283
rect 1318 -1279 1319 -1277
rect 1318 -1285 1319 -1283
rect 1325 -1279 1326 -1277
rect 1325 -1285 1326 -1283
rect 1332 -1279 1333 -1277
rect 1332 -1285 1333 -1283
rect 1339 -1279 1340 -1277
rect 1339 -1285 1340 -1283
rect 1346 -1279 1347 -1277
rect 1346 -1285 1347 -1283
rect 1353 -1279 1354 -1277
rect 1353 -1285 1354 -1283
rect 1360 -1279 1361 -1277
rect 1360 -1285 1361 -1283
rect 1367 -1279 1368 -1277
rect 1367 -1285 1368 -1283
rect 1374 -1279 1375 -1277
rect 1374 -1285 1375 -1283
rect 1381 -1279 1382 -1277
rect 1381 -1285 1382 -1283
rect 1388 -1279 1389 -1277
rect 1388 -1285 1389 -1283
rect 1395 -1279 1396 -1277
rect 1395 -1285 1396 -1283
rect 1402 -1279 1403 -1277
rect 1402 -1285 1403 -1283
rect 1409 -1279 1410 -1277
rect 1409 -1285 1410 -1283
rect 1416 -1279 1417 -1277
rect 1416 -1285 1417 -1283
rect 1423 -1279 1424 -1277
rect 1423 -1285 1424 -1283
rect 1430 -1279 1431 -1277
rect 1430 -1285 1431 -1283
rect 1437 -1279 1438 -1277
rect 1437 -1285 1438 -1283
rect 1444 -1279 1445 -1277
rect 1444 -1285 1445 -1283
rect 1451 -1279 1452 -1277
rect 1451 -1285 1452 -1283
rect 1458 -1279 1459 -1277
rect 1458 -1285 1459 -1283
rect 1465 -1279 1466 -1277
rect 1465 -1285 1466 -1283
rect 1472 -1279 1473 -1277
rect 1472 -1285 1473 -1283
rect 1479 -1279 1480 -1277
rect 1479 -1285 1480 -1283
rect 1486 -1279 1487 -1277
rect 1486 -1285 1487 -1283
rect 1493 -1279 1494 -1277
rect 1493 -1285 1494 -1283
rect 1500 -1279 1501 -1277
rect 1500 -1285 1501 -1283
rect 1507 -1279 1508 -1277
rect 1507 -1285 1508 -1283
rect 1514 -1279 1515 -1277
rect 1514 -1285 1515 -1283
rect 1521 -1279 1522 -1277
rect 1521 -1285 1522 -1283
rect 1528 -1279 1529 -1277
rect 1528 -1285 1529 -1283
rect 1535 -1279 1536 -1277
rect 1535 -1285 1536 -1283
rect 1542 -1279 1543 -1277
rect 1542 -1285 1543 -1283
rect 1549 -1279 1550 -1277
rect 1549 -1285 1550 -1283
rect 1556 -1279 1557 -1277
rect 1556 -1285 1557 -1283
rect 1563 -1279 1564 -1277
rect 1563 -1285 1564 -1283
rect 2 -1398 3 -1396
rect 2 -1404 3 -1402
rect 9 -1398 10 -1396
rect 9 -1404 10 -1402
rect 16 -1398 17 -1396
rect 16 -1404 17 -1402
rect 23 -1398 24 -1396
rect 23 -1404 24 -1402
rect 30 -1398 31 -1396
rect 30 -1404 31 -1402
rect 37 -1398 38 -1396
rect 37 -1404 38 -1402
rect 44 -1398 45 -1396
rect 44 -1404 45 -1402
rect 51 -1398 52 -1396
rect 51 -1404 52 -1402
rect 58 -1398 59 -1396
rect 58 -1404 59 -1402
rect 65 -1398 66 -1396
rect 68 -1398 69 -1396
rect 65 -1404 66 -1402
rect 68 -1404 69 -1402
rect 72 -1398 73 -1396
rect 72 -1404 73 -1402
rect 79 -1398 80 -1396
rect 82 -1398 83 -1396
rect 79 -1404 80 -1402
rect 82 -1404 83 -1402
rect 86 -1398 87 -1396
rect 86 -1404 87 -1402
rect 93 -1398 94 -1396
rect 93 -1404 94 -1402
rect 100 -1398 101 -1396
rect 100 -1404 101 -1402
rect 107 -1398 108 -1396
rect 110 -1398 111 -1396
rect 107 -1404 108 -1402
rect 110 -1404 111 -1402
rect 114 -1398 115 -1396
rect 114 -1404 115 -1402
rect 121 -1398 122 -1396
rect 121 -1404 122 -1402
rect 128 -1398 129 -1396
rect 128 -1404 129 -1402
rect 135 -1398 136 -1396
rect 135 -1404 136 -1402
rect 142 -1398 143 -1396
rect 142 -1404 143 -1402
rect 149 -1398 150 -1396
rect 149 -1404 150 -1402
rect 156 -1398 157 -1396
rect 156 -1404 157 -1402
rect 163 -1398 164 -1396
rect 163 -1404 164 -1402
rect 170 -1398 171 -1396
rect 170 -1404 171 -1402
rect 177 -1398 178 -1396
rect 177 -1404 178 -1402
rect 184 -1398 185 -1396
rect 184 -1404 185 -1402
rect 191 -1398 192 -1396
rect 191 -1404 192 -1402
rect 198 -1398 199 -1396
rect 198 -1404 199 -1402
rect 205 -1398 206 -1396
rect 205 -1404 206 -1402
rect 212 -1398 213 -1396
rect 215 -1398 216 -1396
rect 212 -1404 213 -1402
rect 219 -1398 220 -1396
rect 219 -1404 220 -1402
rect 226 -1398 227 -1396
rect 226 -1404 227 -1402
rect 233 -1398 234 -1396
rect 233 -1404 234 -1402
rect 240 -1398 241 -1396
rect 240 -1404 241 -1402
rect 247 -1398 248 -1396
rect 247 -1404 248 -1402
rect 254 -1398 255 -1396
rect 254 -1404 255 -1402
rect 261 -1398 262 -1396
rect 261 -1404 262 -1402
rect 268 -1398 269 -1396
rect 268 -1404 269 -1402
rect 275 -1398 276 -1396
rect 275 -1404 276 -1402
rect 282 -1398 283 -1396
rect 282 -1404 283 -1402
rect 289 -1398 290 -1396
rect 289 -1404 290 -1402
rect 296 -1398 297 -1396
rect 296 -1404 297 -1402
rect 303 -1398 304 -1396
rect 303 -1404 304 -1402
rect 310 -1398 311 -1396
rect 310 -1404 311 -1402
rect 317 -1398 318 -1396
rect 320 -1398 321 -1396
rect 317 -1404 318 -1402
rect 320 -1404 321 -1402
rect 324 -1398 325 -1396
rect 324 -1404 325 -1402
rect 331 -1398 332 -1396
rect 331 -1404 332 -1402
rect 338 -1398 339 -1396
rect 338 -1404 339 -1402
rect 345 -1398 346 -1396
rect 345 -1404 346 -1402
rect 352 -1398 353 -1396
rect 352 -1404 353 -1402
rect 359 -1398 360 -1396
rect 359 -1404 360 -1402
rect 366 -1398 367 -1396
rect 366 -1404 367 -1402
rect 373 -1398 374 -1396
rect 373 -1404 374 -1402
rect 380 -1398 381 -1396
rect 380 -1404 381 -1402
rect 387 -1398 388 -1396
rect 390 -1398 391 -1396
rect 387 -1404 388 -1402
rect 390 -1404 391 -1402
rect 394 -1398 395 -1396
rect 394 -1404 395 -1402
rect 404 -1398 405 -1396
rect 401 -1404 402 -1402
rect 404 -1404 405 -1402
rect 408 -1398 409 -1396
rect 408 -1404 409 -1402
rect 418 -1398 419 -1396
rect 415 -1404 416 -1402
rect 418 -1404 419 -1402
rect 422 -1398 423 -1396
rect 422 -1404 423 -1402
rect 429 -1398 430 -1396
rect 429 -1404 430 -1402
rect 436 -1398 437 -1396
rect 436 -1404 437 -1402
rect 443 -1398 444 -1396
rect 443 -1404 444 -1402
rect 450 -1398 451 -1396
rect 450 -1404 451 -1402
rect 457 -1398 458 -1396
rect 457 -1404 458 -1402
rect 464 -1398 465 -1396
rect 467 -1398 468 -1396
rect 464 -1404 465 -1402
rect 467 -1404 468 -1402
rect 471 -1398 472 -1396
rect 471 -1404 472 -1402
rect 478 -1398 479 -1396
rect 481 -1398 482 -1396
rect 478 -1404 479 -1402
rect 481 -1404 482 -1402
rect 485 -1398 486 -1396
rect 488 -1398 489 -1396
rect 485 -1404 486 -1402
rect 488 -1404 489 -1402
rect 492 -1398 493 -1396
rect 495 -1398 496 -1396
rect 492 -1404 493 -1402
rect 495 -1404 496 -1402
rect 499 -1398 500 -1396
rect 499 -1404 500 -1402
rect 506 -1398 507 -1396
rect 506 -1404 507 -1402
rect 513 -1398 514 -1396
rect 516 -1398 517 -1396
rect 513 -1404 514 -1402
rect 516 -1404 517 -1402
rect 520 -1398 521 -1396
rect 523 -1398 524 -1396
rect 520 -1404 521 -1402
rect 523 -1404 524 -1402
rect 527 -1398 528 -1396
rect 527 -1404 528 -1402
rect 534 -1398 535 -1396
rect 534 -1404 535 -1402
rect 541 -1398 542 -1396
rect 541 -1404 542 -1402
rect 548 -1398 549 -1396
rect 548 -1404 549 -1402
rect 555 -1398 556 -1396
rect 555 -1404 556 -1402
rect 562 -1398 563 -1396
rect 562 -1404 563 -1402
rect 569 -1398 570 -1396
rect 569 -1404 570 -1402
rect 576 -1398 577 -1396
rect 576 -1404 577 -1402
rect 583 -1398 584 -1396
rect 583 -1404 584 -1402
rect 590 -1398 591 -1396
rect 590 -1404 591 -1402
rect 597 -1398 598 -1396
rect 597 -1404 598 -1402
rect 604 -1398 605 -1396
rect 604 -1404 605 -1402
rect 611 -1398 612 -1396
rect 611 -1404 612 -1402
rect 618 -1398 619 -1396
rect 618 -1404 619 -1402
rect 625 -1398 626 -1396
rect 625 -1404 626 -1402
rect 632 -1398 633 -1396
rect 632 -1404 633 -1402
rect 639 -1398 640 -1396
rect 639 -1404 640 -1402
rect 646 -1398 647 -1396
rect 649 -1398 650 -1396
rect 646 -1404 647 -1402
rect 649 -1404 650 -1402
rect 653 -1398 654 -1396
rect 653 -1404 654 -1402
rect 660 -1398 661 -1396
rect 660 -1404 661 -1402
rect 667 -1398 668 -1396
rect 667 -1404 668 -1402
rect 674 -1398 675 -1396
rect 674 -1404 675 -1402
rect 681 -1398 682 -1396
rect 681 -1404 682 -1402
rect 688 -1398 689 -1396
rect 688 -1404 689 -1402
rect 695 -1398 696 -1396
rect 695 -1404 696 -1402
rect 702 -1398 703 -1396
rect 702 -1404 703 -1402
rect 709 -1398 710 -1396
rect 712 -1398 713 -1396
rect 709 -1404 710 -1402
rect 712 -1404 713 -1402
rect 716 -1398 717 -1396
rect 716 -1404 717 -1402
rect 723 -1398 724 -1396
rect 723 -1404 724 -1402
rect 730 -1398 731 -1396
rect 730 -1404 731 -1402
rect 737 -1398 738 -1396
rect 737 -1404 738 -1402
rect 744 -1398 745 -1396
rect 744 -1404 745 -1402
rect 751 -1398 752 -1396
rect 751 -1404 752 -1402
rect 758 -1398 759 -1396
rect 758 -1404 759 -1402
rect 765 -1398 766 -1396
rect 765 -1404 766 -1402
rect 772 -1398 773 -1396
rect 772 -1404 773 -1402
rect 779 -1398 780 -1396
rect 779 -1404 780 -1402
rect 786 -1398 787 -1396
rect 786 -1404 787 -1402
rect 793 -1398 794 -1396
rect 793 -1404 794 -1402
rect 800 -1398 801 -1396
rect 800 -1404 801 -1402
rect 807 -1398 808 -1396
rect 807 -1404 808 -1402
rect 814 -1398 815 -1396
rect 814 -1404 815 -1402
rect 821 -1398 822 -1396
rect 821 -1404 822 -1402
rect 828 -1398 829 -1396
rect 828 -1404 829 -1402
rect 835 -1398 836 -1396
rect 835 -1404 836 -1402
rect 842 -1398 843 -1396
rect 845 -1398 846 -1396
rect 842 -1404 843 -1402
rect 845 -1404 846 -1402
rect 849 -1398 850 -1396
rect 849 -1404 850 -1402
rect 856 -1398 857 -1396
rect 856 -1404 857 -1402
rect 863 -1398 864 -1396
rect 863 -1404 864 -1402
rect 870 -1398 871 -1396
rect 873 -1398 874 -1396
rect 870 -1404 871 -1402
rect 873 -1404 874 -1402
rect 877 -1398 878 -1396
rect 880 -1398 881 -1396
rect 877 -1404 878 -1402
rect 880 -1404 881 -1402
rect 884 -1398 885 -1396
rect 884 -1404 885 -1402
rect 891 -1398 892 -1396
rect 891 -1404 892 -1402
rect 898 -1398 899 -1396
rect 898 -1404 899 -1402
rect 905 -1398 906 -1396
rect 905 -1404 906 -1402
rect 912 -1398 913 -1396
rect 912 -1404 913 -1402
rect 919 -1398 920 -1396
rect 922 -1398 923 -1396
rect 919 -1404 920 -1402
rect 922 -1404 923 -1402
rect 926 -1398 927 -1396
rect 926 -1404 927 -1402
rect 933 -1398 934 -1396
rect 933 -1404 934 -1402
rect 940 -1398 941 -1396
rect 940 -1404 941 -1402
rect 947 -1398 948 -1396
rect 950 -1398 951 -1396
rect 947 -1404 948 -1402
rect 950 -1404 951 -1402
rect 954 -1398 955 -1396
rect 954 -1404 955 -1402
rect 961 -1398 962 -1396
rect 961 -1404 962 -1402
rect 968 -1398 969 -1396
rect 968 -1404 969 -1402
rect 975 -1398 976 -1396
rect 978 -1398 979 -1396
rect 975 -1404 976 -1402
rect 978 -1404 979 -1402
rect 982 -1398 983 -1396
rect 982 -1404 983 -1402
rect 989 -1398 990 -1396
rect 989 -1404 990 -1402
rect 996 -1398 997 -1396
rect 996 -1404 997 -1402
rect 1003 -1398 1004 -1396
rect 1006 -1398 1007 -1396
rect 1006 -1404 1007 -1402
rect 1010 -1398 1011 -1396
rect 1010 -1404 1011 -1402
rect 1017 -1398 1018 -1396
rect 1017 -1404 1018 -1402
rect 1020 -1404 1021 -1402
rect 1024 -1398 1025 -1396
rect 1024 -1404 1025 -1402
rect 1031 -1398 1032 -1396
rect 1031 -1404 1032 -1402
rect 1038 -1398 1039 -1396
rect 1038 -1404 1039 -1402
rect 1045 -1398 1046 -1396
rect 1045 -1404 1046 -1402
rect 1052 -1398 1053 -1396
rect 1052 -1404 1053 -1402
rect 1059 -1398 1060 -1396
rect 1059 -1404 1060 -1402
rect 1066 -1398 1067 -1396
rect 1066 -1404 1067 -1402
rect 1073 -1398 1074 -1396
rect 1073 -1404 1074 -1402
rect 1080 -1398 1081 -1396
rect 1080 -1404 1081 -1402
rect 1087 -1398 1088 -1396
rect 1087 -1404 1088 -1402
rect 1094 -1398 1095 -1396
rect 1094 -1404 1095 -1402
rect 1101 -1398 1102 -1396
rect 1101 -1404 1102 -1402
rect 1108 -1398 1109 -1396
rect 1108 -1404 1109 -1402
rect 1115 -1398 1116 -1396
rect 1115 -1404 1116 -1402
rect 1122 -1398 1123 -1396
rect 1122 -1404 1123 -1402
rect 1129 -1398 1130 -1396
rect 1129 -1404 1130 -1402
rect 1136 -1398 1137 -1396
rect 1136 -1404 1137 -1402
rect 1143 -1398 1144 -1396
rect 1143 -1404 1144 -1402
rect 1150 -1398 1151 -1396
rect 1150 -1404 1151 -1402
rect 1157 -1398 1158 -1396
rect 1157 -1404 1158 -1402
rect 1164 -1398 1165 -1396
rect 1164 -1404 1165 -1402
rect 1171 -1398 1172 -1396
rect 1171 -1404 1172 -1402
rect 1178 -1398 1179 -1396
rect 1178 -1404 1179 -1402
rect 1185 -1398 1186 -1396
rect 1185 -1404 1186 -1402
rect 1192 -1398 1193 -1396
rect 1192 -1404 1193 -1402
rect 1199 -1398 1200 -1396
rect 1199 -1404 1200 -1402
rect 1206 -1398 1207 -1396
rect 1206 -1404 1207 -1402
rect 1213 -1398 1214 -1396
rect 1213 -1404 1214 -1402
rect 1220 -1398 1221 -1396
rect 1220 -1404 1221 -1402
rect 1227 -1398 1228 -1396
rect 1227 -1404 1228 -1402
rect 1234 -1398 1235 -1396
rect 1234 -1404 1235 -1402
rect 1241 -1398 1242 -1396
rect 1241 -1404 1242 -1402
rect 1248 -1398 1249 -1396
rect 1248 -1404 1249 -1402
rect 1255 -1398 1256 -1396
rect 1255 -1404 1256 -1402
rect 1262 -1398 1263 -1396
rect 1262 -1404 1263 -1402
rect 1269 -1398 1270 -1396
rect 1269 -1404 1270 -1402
rect 1276 -1398 1277 -1396
rect 1276 -1404 1277 -1402
rect 1283 -1398 1284 -1396
rect 1283 -1404 1284 -1402
rect 1290 -1398 1291 -1396
rect 1290 -1404 1291 -1402
rect 1297 -1398 1298 -1396
rect 1297 -1404 1298 -1402
rect 1304 -1398 1305 -1396
rect 1304 -1404 1305 -1402
rect 1311 -1398 1312 -1396
rect 1311 -1404 1312 -1402
rect 1318 -1398 1319 -1396
rect 1318 -1404 1319 -1402
rect 1325 -1398 1326 -1396
rect 1325 -1404 1326 -1402
rect 1332 -1398 1333 -1396
rect 1332 -1404 1333 -1402
rect 1339 -1398 1340 -1396
rect 1339 -1404 1340 -1402
rect 1346 -1398 1347 -1396
rect 1346 -1404 1347 -1402
rect 1353 -1398 1354 -1396
rect 1353 -1404 1354 -1402
rect 1360 -1398 1361 -1396
rect 1360 -1404 1361 -1402
rect 1367 -1398 1368 -1396
rect 1367 -1404 1368 -1402
rect 1374 -1398 1375 -1396
rect 1374 -1404 1375 -1402
rect 1381 -1398 1382 -1396
rect 1381 -1404 1382 -1402
rect 1388 -1398 1389 -1396
rect 1388 -1404 1389 -1402
rect 1395 -1398 1396 -1396
rect 1395 -1404 1396 -1402
rect 1402 -1398 1403 -1396
rect 1402 -1404 1403 -1402
rect 1409 -1398 1410 -1396
rect 1409 -1404 1410 -1402
rect 1416 -1398 1417 -1396
rect 1416 -1404 1417 -1402
rect 1423 -1398 1424 -1396
rect 1423 -1404 1424 -1402
rect 1430 -1398 1431 -1396
rect 1430 -1404 1431 -1402
rect 1437 -1398 1438 -1396
rect 1437 -1404 1438 -1402
rect 1444 -1398 1445 -1396
rect 1444 -1404 1445 -1402
rect 1451 -1398 1452 -1396
rect 1451 -1404 1452 -1402
rect 1458 -1398 1459 -1396
rect 1458 -1404 1459 -1402
rect 1465 -1398 1466 -1396
rect 1465 -1404 1466 -1402
rect 1472 -1398 1473 -1396
rect 1472 -1404 1473 -1402
rect 1479 -1398 1480 -1396
rect 1479 -1404 1480 -1402
rect 1486 -1398 1487 -1396
rect 1486 -1404 1487 -1402
rect 1493 -1398 1494 -1396
rect 1493 -1404 1494 -1402
rect 1500 -1398 1501 -1396
rect 1500 -1404 1501 -1402
rect 1507 -1398 1508 -1396
rect 1507 -1404 1508 -1402
rect 1514 -1398 1515 -1396
rect 1514 -1404 1515 -1402
rect 1521 -1398 1522 -1396
rect 1521 -1404 1522 -1402
rect 1524 -1404 1525 -1402
rect 1528 -1398 1529 -1396
rect 1528 -1404 1529 -1402
rect 1535 -1398 1536 -1396
rect 1535 -1404 1536 -1402
rect 2 -1531 3 -1529
rect 2 -1537 3 -1535
rect 9 -1531 10 -1529
rect 9 -1537 10 -1535
rect 16 -1531 17 -1529
rect 16 -1537 17 -1535
rect 23 -1531 24 -1529
rect 23 -1537 24 -1535
rect 30 -1531 31 -1529
rect 30 -1537 31 -1535
rect 37 -1531 38 -1529
rect 37 -1537 38 -1535
rect 44 -1531 45 -1529
rect 44 -1537 45 -1535
rect 51 -1531 52 -1529
rect 54 -1531 55 -1529
rect 51 -1537 52 -1535
rect 54 -1537 55 -1535
rect 58 -1531 59 -1529
rect 58 -1537 59 -1535
rect 65 -1531 66 -1529
rect 65 -1537 66 -1535
rect 72 -1531 73 -1529
rect 72 -1537 73 -1535
rect 79 -1531 80 -1529
rect 82 -1531 83 -1529
rect 82 -1537 83 -1535
rect 86 -1531 87 -1529
rect 86 -1537 87 -1535
rect 93 -1531 94 -1529
rect 93 -1537 94 -1535
rect 100 -1531 101 -1529
rect 103 -1531 104 -1529
rect 100 -1537 101 -1535
rect 103 -1537 104 -1535
rect 107 -1531 108 -1529
rect 107 -1537 108 -1535
rect 114 -1531 115 -1529
rect 114 -1537 115 -1535
rect 121 -1531 122 -1529
rect 121 -1537 122 -1535
rect 128 -1531 129 -1529
rect 128 -1537 129 -1535
rect 135 -1531 136 -1529
rect 135 -1537 136 -1535
rect 142 -1531 143 -1529
rect 142 -1537 143 -1535
rect 149 -1531 150 -1529
rect 149 -1537 150 -1535
rect 156 -1531 157 -1529
rect 156 -1537 157 -1535
rect 163 -1531 164 -1529
rect 163 -1537 164 -1535
rect 173 -1531 174 -1529
rect 170 -1537 171 -1535
rect 173 -1537 174 -1535
rect 177 -1531 178 -1529
rect 177 -1537 178 -1535
rect 184 -1531 185 -1529
rect 184 -1537 185 -1535
rect 191 -1531 192 -1529
rect 191 -1537 192 -1535
rect 198 -1531 199 -1529
rect 198 -1537 199 -1535
rect 205 -1531 206 -1529
rect 205 -1537 206 -1535
rect 212 -1531 213 -1529
rect 212 -1537 213 -1535
rect 219 -1531 220 -1529
rect 219 -1537 220 -1535
rect 226 -1531 227 -1529
rect 226 -1537 227 -1535
rect 233 -1531 234 -1529
rect 233 -1537 234 -1535
rect 240 -1531 241 -1529
rect 240 -1537 241 -1535
rect 247 -1531 248 -1529
rect 247 -1537 248 -1535
rect 254 -1531 255 -1529
rect 254 -1537 255 -1535
rect 261 -1531 262 -1529
rect 261 -1537 262 -1535
rect 268 -1531 269 -1529
rect 268 -1537 269 -1535
rect 275 -1531 276 -1529
rect 275 -1537 276 -1535
rect 282 -1531 283 -1529
rect 282 -1537 283 -1535
rect 289 -1531 290 -1529
rect 289 -1537 290 -1535
rect 296 -1531 297 -1529
rect 296 -1537 297 -1535
rect 303 -1531 304 -1529
rect 303 -1537 304 -1535
rect 310 -1531 311 -1529
rect 310 -1537 311 -1535
rect 317 -1531 318 -1529
rect 317 -1537 318 -1535
rect 324 -1531 325 -1529
rect 324 -1537 325 -1535
rect 331 -1531 332 -1529
rect 331 -1537 332 -1535
rect 338 -1531 339 -1529
rect 338 -1537 339 -1535
rect 345 -1531 346 -1529
rect 345 -1537 346 -1535
rect 352 -1531 353 -1529
rect 352 -1537 353 -1535
rect 359 -1531 360 -1529
rect 359 -1537 360 -1535
rect 366 -1531 367 -1529
rect 366 -1537 367 -1535
rect 373 -1531 374 -1529
rect 373 -1537 374 -1535
rect 380 -1531 381 -1529
rect 380 -1537 381 -1535
rect 387 -1531 388 -1529
rect 387 -1537 388 -1535
rect 394 -1531 395 -1529
rect 397 -1531 398 -1529
rect 394 -1537 395 -1535
rect 397 -1537 398 -1535
rect 401 -1531 402 -1529
rect 401 -1537 402 -1535
rect 408 -1531 409 -1529
rect 408 -1537 409 -1535
rect 415 -1531 416 -1529
rect 415 -1537 416 -1535
rect 422 -1531 423 -1529
rect 422 -1537 423 -1535
rect 429 -1531 430 -1529
rect 432 -1531 433 -1529
rect 432 -1537 433 -1535
rect 436 -1531 437 -1529
rect 436 -1537 437 -1535
rect 443 -1531 444 -1529
rect 443 -1537 444 -1535
rect 450 -1531 451 -1529
rect 450 -1537 451 -1535
rect 457 -1531 458 -1529
rect 457 -1537 458 -1535
rect 464 -1531 465 -1529
rect 464 -1537 465 -1535
rect 471 -1531 472 -1529
rect 474 -1531 475 -1529
rect 471 -1537 472 -1535
rect 474 -1537 475 -1535
rect 478 -1531 479 -1529
rect 478 -1537 479 -1535
rect 485 -1531 486 -1529
rect 485 -1537 486 -1535
rect 492 -1531 493 -1529
rect 492 -1537 493 -1535
rect 499 -1531 500 -1529
rect 502 -1531 503 -1529
rect 499 -1537 500 -1535
rect 502 -1537 503 -1535
rect 506 -1531 507 -1529
rect 506 -1537 507 -1535
rect 513 -1531 514 -1529
rect 513 -1537 514 -1535
rect 520 -1531 521 -1529
rect 520 -1537 521 -1535
rect 527 -1531 528 -1529
rect 527 -1537 528 -1535
rect 534 -1531 535 -1529
rect 534 -1537 535 -1535
rect 541 -1531 542 -1529
rect 541 -1537 542 -1535
rect 548 -1531 549 -1529
rect 548 -1537 549 -1535
rect 555 -1531 556 -1529
rect 555 -1537 556 -1535
rect 562 -1531 563 -1529
rect 562 -1537 563 -1535
rect 569 -1531 570 -1529
rect 569 -1537 570 -1535
rect 576 -1531 577 -1529
rect 579 -1531 580 -1529
rect 576 -1537 577 -1535
rect 579 -1537 580 -1535
rect 583 -1531 584 -1529
rect 583 -1537 584 -1535
rect 590 -1531 591 -1529
rect 590 -1537 591 -1535
rect 597 -1531 598 -1529
rect 600 -1531 601 -1529
rect 600 -1537 601 -1535
rect 604 -1531 605 -1529
rect 604 -1537 605 -1535
rect 611 -1531 612 -1529
rect 611 -1537 612 -1535
rect 618 -1531 619 -1529
rect 618 -1537 619 -1535
rect 625 -1531 626 -1529
rect 625 -1537 626 -1535
rect 632 -1531 633 -1529
rect 632 -1537 633 -1535
rect 639 -1531 640 -1529
rect 639 -1537 640 -1535
rect 646 -1531 647 -1529
rect 646 -1537 647 -1535
rect 653 -1531 654 -1529
rect 653 -1537 654 -1535
rect 660 -1531 661 -1529
rect 660 -1537 661 -1535
rect 667 -1531 668 -1529
rect 667 -1537 668 -1535
rect 674 -1531 675 -1529
rect 677 -1531 678 -1529
rect 674 -1537 675 -1535
rect 677 -1537 678 -1535
rect 681 -1531 682 -1529
rect 684 -1531 685 -1529
rect 681 -1537 682 -1535
rect 684 -1537 685 -1535
rect 688 -1531 689 -1529
rect 688 -1537 689 -1535
rect 695 -1531 696 -1529
rect 695 -1537 696 -1535
rect 702 -1531 703 -1529
rect 702 -1537 703 -1535
rect 709 -1531 710 -1529
rect 709 -1537 710 -1535
rect 716 -1531 717 -1529
rect 716 -1537 717 -1535
rect 723 -1531 724 -1529
rect 726 -1531 727 -1529
rect 723 -1537 724 -1535
rect 726 -1537 727 -1535
rect 730 -1531 731 -1529
rect 730 -1537 731 -1535
rect 737 -1531 738 -1529
rect 737 -1537 738 -1535
rect 744 -1531 745 -1529
rect 744 -1537 745 -1535
rect 751 -1531 752 -1529
rect 751 -1537 752 -1535
rect 758 -1531 759 -1529
rect 758 -1537 759 -1535
rect 765 -1531 766 -1529
rect 768 -1531 769 -1529
rect 765 -1537 766 -1535
rect 768 -1537 769 -1535
rect 772 -1531 773 -1529
rect 772 -1537 773 -1535
rect 779 -1531 780 -1529
rect 779 -1537 780 -1535
rect 786 -1531 787 -1529
rect 786 -1537 787 -1535
rect 793 -1531 794 -1529
rect 793 -1537 794 -1535
rect 800 -1531 801 -1529
rect 803 -1531 804 -1529
rect 800 -1537 801 -1535
rect 803 -1537 804 -1535
rect 807 -1531 808 -1529
rect 807 -1537 808 -1535
rect 814 -1531 815 -1529
rect 817 -1531 818 -1529
rect 814 -1537 815 -1535
rect 817 -1537 818 -1535
rect 821 -1531 822 -1529
rect 821 -1537 822 -1535
rect 828 -1531 829 -1529
rect 831 -1531 832 -1529
rect 828 -1537 829 -1535
rect 831 -1537 832 -1535
rect 835 -1531 836 -1529
rect 838 -1531 839 -1529
rect 835 -1537 836 -1535
rect 838 -1537 839 -1535
rect 842 -1531 843 -1529
rect 842 -1537 843 -1535
rect 849 -1531 850 -1529
rect 849 -1537 850 -1535
rect 856 -1531 857 -1529
rect 859 -1531 860 -1529
rect 859 -1537 860 -1535
rect 863 -1531 864 -1529
rect 863 -1537 864 -1535
rect 870 -1531 871 -1529
rect 870 -1537 871 -1535
rect 877 -1531 878 -1529
rect 880 -1531 881 -1529
rect 877 -1537 878 -1535
rect 884 -1531 885 -1529
rect 884 -1537 885 -1535
rect 891 -1531 892 -1529
rect 891 -1537 892 -1535
rect 898 -1531 899 -1529
rect 898 -1537 899 -1535
rect 905 -1531 906 -1529
rect 905 -1537 906 -1535
rect 912 -1531 913 -1529
rect 912 -1537 913 -1535
rect 919 -1531 920 -1529
rect 919 -1537 920 -1535
rect 926 -1531 927 -1529
rect 926 -1537 927 -1535
rect 933 -1531 934 -1529
rect 933 -1537 934 -1535
rect 940 -1531 941 -1529
rect 940 -1537 941 -1535
rect 947 -1531 948 -1529
rect 947 -1537 948 -1535
rect 954 -1531 955 -1529
rect 954 -1537 955 -1535
rect 961 -1531 962 -1529
rect 961 -1537 962 -1535
rect 968 -1531 969 -1529
rect 968 -1537 969 -1535
rect 975 -1531 976 -1529
rect 975 -1537 976 -1535
rect 982 -1531 983 -1529
rect 982 -1537 983 -1535
rect 989 -1531 990 -1529
rect 992 -1531 993 -1529
rect 989 -1537 990 -1535
rect 992 -1537 993 -1535
rect 999 -1531 1000 -1529
rect 996 -1537 997 -1535
rect 999 -1537 1000 -1535
rect 1003 -1531 1004 -1529
rect 1003 -1537 1004 -1535
rect 1010 -1531 1011 -1529
rect 1010 -1537 1011 -1535
rect 1017 -1531 1018 -1529
rect 1017 -1537 1018 -1535
rect 1024 -1531 1025 -1529
rect 1024 -1537 1025 -1535
rect 1031 -1531 1032 -1529
rect 1031 -1537 1032 -1535
rect 1038 -1531 1039 -1529
rect 1038 -1537 1039 -1535
rect 1045 -1531 1046 -1529
rect 1045 -1537 1046 -1535
rect 1052 -1531 1053 -1529
rect 1052 -1537 1053 -1535
rect 1059 -1531 1060 -1529
rect 1059 -1537 1060 -1535
rect 1066 -1531 1067 -1529
rect 1066 -1537 1067 -1535
rect 1073 -1531 1074 -1529
rect 1076 -1531 1077 -1529
rect 1073 -1537 1074 -1535
rect 1076 -1537 1077 -1535
rect 1080 -1531 1081 -1529
rect 1080 -1537 1081 -1535
rect 1087 -1531 1088 -1529
rect 1087 -1537 1088 -1535
rect 1094 -1531 1095 -1529
rect 1094 -1537 1095 -1535
rect 1101 -1531 1102 -1529
rect 1101 -1537 1102 -1535
rect 1108 -1531 1109 -1529
rect 1108 -1537 1109 -1535
rect 1115 -1531 1116 -1529
rect 1115 -1537 1116 -1535
rect 1122 -1531 1123 -1529
rect 1125 -1531 1126 -1529
rect 1122 -1537 1123 -1535
rect 1129 -1531 1130 -1529
rect 1129 -1537 1130 -1535
rect 1136 -1531 1137 -1529
rect 1136 -1537 1137 -1535
rect 1143 -1531 1144 -1529
rect 1143 -1537 1144 -1535
rect 1150 -1531 1151 -1529
rect 1150 -1537 1151 -1535
rect 1153 -1537 1154 -1535
rect 1157 -1531 1158 -1529
rect 1157 -1537 1158 -1535
rect 1164 -1531 1165 -1529
rect 1164 -1537 1165 -1535
rect 1171 -1531 1172 -1529
rect 1171 -1537 1172 -1535
rect 1178 -1531 1179 -1529
rect 1178 -1537 1179 -1535
rect 1185 -1531 1186 -1529
rect 1185 -1537 1186 -1535
rect 1192 -1531 1193 -1529
rect 1192 -1537 1193 -1535
rect 1199 -1531 1200 -1529
rect 1199 -1537 1200 -1535
rect 1206 -1531 1207 -1529
rect 1206 -1537 1207 -1535
rect 1213 -1531 1214 -1529
rect 1213 -1537 1214 -1535
rect 1220 -1531 1221 -1529
rect 1220 -1537 1221 -1535
rect 1227 -1531 1228 -1529
rect 1227 -1537 1228 -1535
rect 1234 -1531 1235 -1529
rect 1234 -1537 1235 -1535
rect 1241 -1531 1242 -1529
rect 1241 -1537 1242 -1535
rect 1248 -1531 1249 -1529
rect 1248 -1537 1249 -1535
rect 1255 -1531 1256 -1529
rect 1255 -1537 1256 -1535
rect 1262 -1531 1263 -1529
rect 1262 -1537 1263 -1535
rect 1269 -1531 1270 -1529
rect 1269 -1537 1270 -1535
rect 1276 -1531 1277 -1529
rect 1276 -1537 1277 -1535
rect 1283 -1531 1284 -1529
rect 1283 -1537 1284 -1535
rect 1290 -1531 1291 -1529
rect 1290 -1537 1291 -1535
rect 1297 -1531 1298 -1529
rect 1297 -1537 1298 -1535
rect 1304 -1531 1305 -1529
rect 1304 -1537 1305 -1535
rect 1311 -1531 1312 -1529
rect 1311 -1537 1312 -1535
rect 1318 -1531 1319 -1529
rect 1318 -1537 1319 -1535
rect 1325 -1531 1326 -1529
rect 1325 -1537 1326 -1535
rect 1332 -1531 1333 -1529
rect 1332 -1537 1333 -1535
rect 1339 -1531 1340 -1529
rect 1339 -1537 1340 -1535
rect 1346 -1531 1347 -1529
rect 1346 -1537 1347 -1535
rect 1353 -1531 1354 -1529
rect 1353 -1537 1354 -1535
rect 1360 -1531 1361 -1529
rect 1360 -1537 1361 -1535
rect 1367 -1531 1368 -1529
rect 1367 -1537 1368 -1535
rect 1374 -1531 1375 -1529
rect 1374 -1537 1375 -1535
rect 1381 -1531 1382 -1529
rect 1381 -1537 1382 -1535
rect 1388 -1531 1389 -1529
rect 1388 -1537 1389 -1535
rect 1395 -1531 1396 -1529
rect 1395 -1537 1396 -1535
rect 1402 -1531 1403 -1529
rect 1402 -1537 1403 -1535
rect 1409 -1531 1410 -1529
rect 1409 -1537 1410 -1535
rect 1416 -1531 1417 -1529
rect 1416 -1537 1417 -1535
rect 1423 -1531 1424 -1529
rect 1423 -1537 1424 -1535
rect 1430 -1531 1431 -1529
rect 1430 -1537 1431 -1535
rect 1437 -1531 1438 -1529
rect 1437 -1537 1438 -1535
rect 1444 -1531 1445 -1529
rect 1444 -1537 1445 -1535
rect 1451 -1531 1452 -1529
rect 1451 -1537 1452 -1535
rect 1458 -1531 1459 -1529
rect 1458 -1537 1459 -1535
rect 1465 -1531 1466 -1529
rect 1465 -1537 1466 -1535
rect 1472 -1531 1473 -1529
rect 1472 -1537 1473 -1535
rect 1479 -1531 1480 -1529
rect 1479 -1537 1480 -1535
rect 1486 -1531 1487 -1529
rect 1486 -1537 1487 -1535
rect 1493 -1531 1494 -1529
rect 1493 -1537 1494 -1535
rect 1500 -1531 1501 -1529
rect 1500 -1537 1501 -1535
rect 1507 -1531 1508 -1529
rect 1507 -1537 1508 -1535
rect 1514 -1531 1515 -1529
rect 1514 -1537 1515 -1535
rect 1521 -1531 1522 -1529
rect 1524 -1531 1525 -1529
rect 1521 -1537 1522 -1535
rect 1524 -1537 1525 -1535
rect 1528 -1531 1529 -1529
rect 1528 -1537 1529 -1535
rect 1535 -1531 1536 -1529
rect 1535 -1537 1536 -1535
rect 2 -1638 3 -1636
rect 2 -1644 3 -1642
rect 9 -1638 10 -1636
rect 9 -1644 10 -1642
rect 16 -1638 17 -1636
rect 16 -1644 17 -1642
rect 23 -1638 24 -1636
rect 23 -1644 24 -1642
rect 30 -1638 31 -1636
rect 30 -1644 31 -1642
rect 37 -1638 38 -1636
rect 37 -1644 38 -1642
rect 44 -1638 45 -1636
rect 44 -1644 45 -1642
rect 51 -1638 52 -1636
rect 51 -1644 52 -1642
rect 58 -1638 59 -1636
rect 58 -1644 59 -1642
rect 65 -1638 66 -1636
rect 65 -1644 66 -1642
rect 72 -1638 73 -1636
rect 75 -1638 76 -1636
rect 72 -1644 73 -1642
rect 75 -1644 76 -1642
rect 79 -1638 80 -1636
rect 79 -1644 80 -1642
rect 86 -1638 87 -1636
rect 86 -1644 87 -1642
rect 93 -1638 94 -1636
rect 93 -1644 94 -1642
rect 100 -1638 101 -1636
rect 100 -1644 101 -1642
rect 107 -1638 108 -1636
rect 107 -1644 108 -1642
rect 110 -1644 111 -1642
rect 114 -1638 115 -1636
rect 114 -1644 115 -1642
rect 121 -1638 122 -1636
rect 121 -1644 122 -1642
rect 128 -1638 129 -1636
rect 131 -1638 132 -1636
rect 128 -1644 129 -1642
rect 131 -1644 132 -1642
rect 135 -1638 136 -1636
rect 135 -1644 136 -1642
rect 142 -1638 143 -1636
rect 145 -1638 146 -1636
rect 142 -1644 143 -1642
rect 145 -1644 146 -1642
rect 149 -1638 150 -1636
rect 149 -1644 150 -1642
rect 156 -1638 157 -1636
rect 156 -1644 157 -1642
rect 163 -1638 164 -1636
rect 163 -1644 164 -1642
rect 170 -1638 171 -1636
rect 170 -1644 171 -1642
rect 177 -1638 178 -1636
rect 177 -1644 178 -1642
rect 184 -1638 185 -1636
rect 184 -1644 185 -1642
rect 191 -1638 192 -1636
rect 191 -1644 192 -1642
rect 198 -1638 199 -1636
rect 198 -1644 199 -1642
rect 205 -1638 206 -1636
rect 205 -1644 206 -1642
rect 212 -1638 213 -1636
rect 212 -1644 213 -1642
rect 219 -1638 220 -1636
rect 219 -1644 220 -1642
rect 226 -1638 227 -1636
rect 226 -1644 227 -1642
rect 233 -1638 234 -1636
rect 233 -1644 234 -1642
rect 240 -1638 241 -1636
rect 240 -1644 241 -1642
rect 247 -1638 248 -1636
rect 247 -1644 248 -1642
rect 254 -1638 255 -1636
rect 254 -1644 255 -1642
rect 261 -1638 262 -1636
rect 261 -1644 262 -1642
rect 268 -1638 269 -1636
rect 271 -1638 272 -1636
rect 268 -1644 269 -1642
rect 271 -1644 272 -1642
rect 275 -1638 276 -1636
rect 275 -1644 276 -1642
rect 282 -1638 283 -1636
rect 282 -1644 283 -1642
rect 289 -1638 290 -1636
rect 289 -1644 290 -1642
rect 296 -1638 297 -1636
rect 296 -1644 297 -1642
rect 303 -1638 304 -1636
rect 303 -1644 304 -1642
rect 310 -1638 311 -1636
rect 310 -1644 311 -1642
rect 317 -1638 318 -1636
rect 317 -1644 318 -1642
rect 324 -1638 325 -1636
rect 324 -1644 325 -1642
rect 331 -1638 332 -1636
rect 331 -1644 332 -1642
rect 338 -1638 339 -1636
rect 338 -1644 339 -1642
rect 348 -1638 349 -1636
rect 345 -1644 346 -1642
rect 352 -1638 353 -1636
rect 352 -1644 353 -1642
rect 359 -1638 360 -1636
rect 359 -1644 360 -1642
rect 366 -1638 367 -1636
rect 369 -1638 370 -1636
rect 366 -1644 367 -1642
rect 369 -1644 370 -1642
rect 373 -1638 374 -1636
rect 373 -1644 374 -1642
rect 380 -1638 381 -1636
rect 380 -1644 381 -1642
rect 387 -1638 388 -1636
rect 387 -1644 388 -1642
rect 394 -1638 395 -1636
rect 394 -1644 395 -1642
rect 401 -1638 402 -1636
rect 401 -1644 402 -1642
rect 408 -1638 409 -1636
rect 408 -1644 409 -1642
rect 415 -1638 416 -1636
rect 415 -1644 416 -1642
rect 422 -1638 423 -1636
rect 422 -1644 423 -1642
rect 429 -1638 430 -1636
rect 429 -1644 430 -1642
rect 439 -1638 440 -1636
rect 436 -1644 437 -1642
rect 443 -1638 444 -1636
rect 446 -1638 447 -1636
rect 446 -1644 447 -1642
rect 450 -1638 451 -1636
rect 450 -1644 451 -1642
rect 457 -1638 458 -1636
rect 457 -1644 458 -1642
rect 464 -1638 465 -1636
rect 464 -1644 465 -1642
rect 471 -1638 472 -1636
rect 474 -1638 475 -1636
rect 471 -1644 472 -1642
rect 474 -1644 475 -1642
rect 478 -1638 479 -1636
rect 478 -1644 479 -1642
rect 485 -1638 486 -1636
rect 485 -1644 486 -1642
rect 492 -1638 493 -1636
rect 492 -1644 493 -1642
rect 499 -1638 500 -1636
rect 502 -1638 503 -1636
rect 499 -1644 500 -1642
rect 502 -1644 503 -1642
rect 506 -1638 507 -1636
rect 506 -1644 507 -1642
rect 513 -1638 514 -1636
rect 513 -1644 514 -1642
rect 520 -1638 521 -1636
rect 520 -1644 521 -1642
rect 527 -1638 528 -1636
rect 527 -1644 528 -1642
rect 534 -1638 535 -1636
rect 534 -1644 535 -1642
rect 541 -1638 542 -1636
rect 541 -1644 542 -1642
rect 548 -1638 549 -1636
rect 548 -1644 549 -1642
rect 555 -1638 556 -1636
rect 558 -1638 559 -1636
rect 555 -1644 556 -1642
rect 562 -1638 563 -1636
rect 565 -1638 566 -1636
rect 562 -1644 563 -1642
rect 565 -1644 566 -1642
rect 569 -1638 570 -1636
rect 569 -1644 570 -1642
rect 576 -1638 577 -1636
rect 576 -1644 577 -1642
rect 583 -1638 584 -1636
rect 583 -1644 584 -1642
rect 590 -1638 591 -1636
rect 590 -1644 591 -1642
rect 597 -1644 598 -1642
rect 604 -1638 605 -1636
rect 604 -1644 605 -1642
rect 611 -1638 612 -1636
rect 611 -1644 612 -1642
rect 618 -1638 619 -1636
rect 621 -1638 622 -1636
rect 618 -1644 619 -1642
rect 621 -1644 622 -1642
rect 625 -1638 626 -1636
rect 625 -1644 626 -1642
rect 632 -1638 633 -1636
rect 632 -1644 633 -1642
rect 639 -1638 640 -1636
rect 639 -1644 640 -1642
rect 646 -1638 647 -1636
rect 649 -1638 650 -1636
rect 646 -1644 647 -1642
rect 649 -1644 650 -1642
rect 653 -1638 654 -1636
rect 653 -1644 654 -1642
rect 660 -1638 661 -1636
rect 660 -1644 661 -1642
rect 667 -1638 668 -1636
rect 667 -1644 668 -1642
rect 674 -1638 675 -1636
rect 674 -1644 675 -1642
rect 681 -1638 682 -1636
rect 681 -1644 682 -1642
rect 688 -1638 689 -1636
rect 688 -1644 689 -1642
rect 695 -1638 696 -1636
rect 695 -1644 696 -1642
rect 702 -1638 703 -1636
rect 702 -1644 703 -1642
rect 709 -1638 710 -1636
rect 709 -1644 710 -1642
rect 716 -1638 717 -1636
rect 716 -1644 717 -1642
rect 723 -1638 724 -1636
rect 723 -1644 724 -1642
rect 730 -1638 731 -1636
rect 730 -1644 731 -1642
rect 737 -1638 738 -1636
rect 740 -1638 741 -1636
rect 737 -1644 738 -1642
rect 740 -1644 741 -1642
rect 744 -1638 745 -1636
rect 744 -1644 745 -1642
rect 751 -1638 752 -1636
rect 754 -1638 755 -1636
rect 751 -1644 752 -1642
rect 754 -1644 755 -1642
rect 758 -1638 759 -1636
rect 758 -1644 759 -1642
rect 765 -1638 766 -1636
rect 765 -1644 766 -1642
rect 772 -1638 773 -1636
rect 772 -1644 773 -1642
rect 779 -1638 780 -1636
rect 782 -1638 783 -1636
rect 779 -1644 780 -1642
rect 782 -1644 783 -1642
rect 786 -1638 787 -1636
rect 786 -1644 787 -1642
rect 793 -1638 794 -1636
rect 793 -1644 794 -1642
rect 800 -1638 801 -1636
rect 800 -1644 801 -1642
rect 807 -1638 808 -1636
rect 807 -1644 808 -1642
rect 814 -1638 815 -1636
rect 817 -1638 818 -1636
rect 817 -1644 818 -1642
rect 821 -1638 822 -1636
rect 821 -1644 822 -1642
rect 828 -1638 829 -1636
rect 831 -1638 832 -1636
rect 828 -1644 829 -1642
rect 831 -1644 832 -1642
rect 835 -1638 836 -1636
rect 835 -1644 836 -1642
rect 842 -1638 843 -1636
rect 842 -1644 843 -1642
rect 849 -1638 850 -1636
rect 849 -1644 850 -1642
rect 856 -1638 857 -1636
rect 856 -1644 857 -1642
rect 863 -1638 864 -1636
rect 863 -1644 864 -1642
rect 870 -1638 871 -1636
rect 870 -1644 871 -1642
rect 877 -1638 878 -1636
rect 880 -1638 881 -1636
rect 877 -1644 878 -1642
rect 880 -1644 881 -1642
rect 884 -1638 885 -1636
rect 884 -1644 885 -1642
rect 891 -1638 892 -1636
rect 891 -1644 892 -1642
rect 898 -1638 899 -1636
rect 898 -1644 899 -1642
rect 905 -1638 906 -1636
rect 905 -1644 906 -1642
rect 912 -1638 913 -1636
rect 912 -1644 913 -1642
rect 919 -1638 920 -1636
rect 919 -1644 920 -1642
rect 926 -1638 927 -1636
rect 926 -1644 927 -1642
rect 933 -1638 934 -1636
rect 933 -1644 934 -1642
rect 940 -1638 941 -1636
rect 940 -1644 941 -1642
rect 947 -1638 948 -1636
rect 947 -1644 948 -1642
rect 954 -1638 955 -1636
rect 957 -1638 958 -1636
rect 954 -1644 955 -1642
rect 961 -1638 962 -1636
rect 961 -1644 962 -1642
rect 968 -1638 969 -1636
rect 968 -1644 969 -1642
rect 975 -1638 976 -1636
rect 975 -1644 976 -1642
rect 982 -1638 983 -1636
rect 982 -1644 983 -1642
rect 989 -1638 990 -1636
rect 992 -1638 993 -1636
rect 992 -1644 993 -1642
rect 996 -1638 997 -1636
rect 996 -1644 997 -1642
rect 1003 -1638 1004 -1636
rect 1003 -1644 1004 -1642
rect 1010 -1638 1011 -1636
rect 1010 -1644 1011 -1642
rect 1017 -1638 1018 -1636
rect 1017 -1644 1018 -1642
rect 1024 -1638 1025 -1636
rect 1024 -1644 1025 -1642
rect 1031 -1638 1032 -1636
rect 1031 -1644 1032 -1642
rect 1038 -1638 1039 -1636
rect 1038 -1644 1039 -1642
rect 1045 -1638 1046 -1636
rect 1045 -1644 1046 -1642
rect 1052 -1638 1053 -1636
rect 1052 -1644 1053 -1642
rect 1059 -1638 1060 -1636
rect 1059 -1644 1060 -1642
rect 1066 -1638 1067 -1636
rect 1066 -1644 1067 -1642
rect 1073 -1638 1074 -1636
rect 1073 -1644 1074 -1642
rect 1080 -1638 1081 -1636
rect 1080 -1644 1081 -1642
rect 1087 -1638 1088 -1636
rect 1087 -1644 1088 -1642
rect 1094 -1638 1095 -1636
rect 1094 -1644 1095 -1642
rect 1101 -1638 1102 -1636
rect 1101 -1644 1102 -1642
rect 1108 -1638 1109 -1636
rect 1108 -1644 1109 -1642
rect 1115 -1638 1116 -1636
rect 1115 -1644 1116 -1642
rect 1122 -1638 1123 -1636
rect 1122 -1644 1123 -1642
rect 1129 -1638 1130 -1636
rect 1129 -1644 1130 -1642
rect 1136 -1638 1137 -1636
rect 1136 -1644 1137 -1642
rect 1143 -1638 1144 -1636
rect 1143 -1644 1144 -1642
rect 1150 -1638 1151 -1636
rect 1153 -1638 1154 -1636
rect 1150 -1644 1151 -1642
rect 1157 -1638 1158 -1636
rect 1157 -1644 1158 -1642
rect 1164 -1638 1165 -1636
rect 1164 -1644 1165 -1642
rect 1171 -1638 1172 -1636
rect 1171 -1644 1172 -1642
rect 1178 -1638 1179 -1636
rect 1178 -1644 1179 -1642
rect 1185 -1638 1186 -1636
rect 1185 -1644 1186 -1642
rect 1192 -1638 1193 -1636
rect 1192 -1644 1193 -1642
rect 1199 -1638 1200 -1636
rect 1199 -1644 1200 -1642
rect 1206 -1638 1207 -1636
rect 1206 -1644 1207 -1642
rect 1213 -1638 1214 -1636
rect 1213 -1644 1214 -1642
rect 1220 -1638 1221 -1636
rect 1220 -1644 1221 -1642
rect 1227 -1638 1228 -1636
rect 1227 -1644 1228 -1642
rect 1234 -1638 1235 -1636
rect 1234 -1644 1235 -1642
rect 1241 -1638 1242 -1636
rect 1241 -1644 1242 -1642
rect 1248 -1638 1249 -1636
rect 1248 -1644 1249 -1642
rect 1255 -1638 1256 -1636
rect 1255 -1644 1256 -1642
rect 1262 -1638 1263 -1636
rect 1262 -1644 1263 -1642
rect 1269 -1638 1270 -1636
rect 1269 -1644 1270 -1642
rect 1276 -1638 1277 -1636
rect 1276 -1644 1277 -1642
rect 1283 -1638 1284 -1636
rect 1283 -1644 1284 -1642
rect 1290 -1638 1291 -1636
rect 1290 -1644 1291 -1642
rect 1297 -1638 1298 -1636
rect 1297 -1644 1298 -1642
rect 1304 -1638 1305 -1636
rect 1304 -1644 1305 -1642
rect 1311 -1638 1312 -1636
rect 1311 -1644 1312 -1642
rect 1318 -1638 1319 -1636
rect 1318 -1644 1319 -1642
rect 1325 -1638 1326 -1636
rect 1325 -1644 1326 -1642
rect 1332 -1638 1333 -1636
rect 1332 -1644 1333 -1642
rect 1339 -1638 1340 -1636
rect 1339 -1644 1340 -1642
rect 1346 -1638 1347 -1636
rect 1349 -1638 1350 -1636
rect 1346 -1644 1347 -1642
rect 1349 -1644 1350 -1642
rect 1353 -1638 1354 -1636
rect 1353 -1644 1354 -1642
rect 1360 -1638 1361 -1636
rect 1360 -1644 1361 -1642
rect 1367 -1638 1368 -1636
rect 1367 -1644 1368 -1642
rect 1374 -1638 1375 -1636
rect 1374 -1644 1375 -1642
rect 1381 -1638 1382 -1636
rect 1381 -1644 1382 -1642
rect 1388 -1638 1389 -1636
rect 1388 -1644 1389 -1642
rect 1395 -1638 1396 -1636
rect 1395 -1644 1396 -1642
rect 1402 -1638 1403 -1636
rect 1402 -1644 1403 -1642
rect 1409 -1638 1410 -1636
rect 1409 -1644 1410 -1642
rect 1416 -1638 1417 -1636
rect 1416 -1644 1417 -1642
rect 1423 -1638 1424 -1636
rect 1423 -1644 1424 -1642
rect 1430 -1638 1431 -1636
rect 1430 -1644 1431 -1642
rect 1437 -1638 1438 -1636
rect 1437 -1644 1438 -1642
rect 1451 -1638 1452 -1636
rect 1451 -1644 1452 -1642
rect 9 -1763 10 -1761
rect 9 -1769 10 -1767
rect 16 -1763 17 -1761
rect 16 -1769 17 -1767
rect 23 -1763 24 -1761
rect 23 -1769 24 -1767
rect 30 -1763 31 -1761
rect 30 -1769 31 -1767
rect 37 -1763 38 -1761
rect 37 -1769 38 -1767
rect 44 -1763 45 -1761
rect 44 -1769 45 -1767
rect 51 -1763 52 -1761
rect 51 -1769 52 -1767
rect 58 -1763 59 -1761
rect 58 -1769 59 -1767
rect 65 -1763 66 -1761
rect 65 -1769 66 -1767
rect 72 -1763 73 -1761
rect 75 -1763 76 -1761
rect 72 -1769 73 -1767
rect 75 -1769 76 -1767
rect 79 -1763 80 -1761
rect 82 -1763 83 -1761
rect 79 -1769 80 -1767
rect 82 -1769 83 -1767
rect 86 -1763 87 -1761
rect 86 -1769 87 -1767
rect 93 -1763 94 -1761
rect 93 -1769 94 -1767
rect 100 -1763 101 -1761
rect 100 -1769 101 -1767
rect 107 -1763 108 -1761
rect 110 -1763 111 -1761
rect 107 -1769 108 -1767
rect 114 -1763 115 -1761
rect 114 -1769 115 -1767
rect 121 -1763 122 -1761
rect 121 -1769 122 -1767
rect 128 -1763 129 -1761
rect 128 -1769 129 -1767
rect 135 -1763 136 -1761
rect 135 -1769 136 -1767
rect 142 -1763 143 -1761
rect 142 -1769 143 -1767
rect 149 -1763 150 -1761
rect 149 -1769 150 -1767
rect 156 -1763 157 -1761
rect 156 -1769 157 -1767
rect 163 -1763 164 -1761
rect 163 -1769 164 -1767
rect 170 -1763 171 -1761
rect 170 -1769 171 -1767
rect 177 -1763 178 -1761
rect 177 -1769 178 -1767
rect 184 -1763 185 -1761
rect 184 -1769 185 -1767
rect 191 -1763 192 -1761
rect 191 -1769 192 -1767
rect 198 -1763 199 -1761
rect 198 -1769 199 -1767
rect 205 -1763 206 -1761
rect 205 -1769 206 -1767
rect 212 -1763 213 -1761
rect 212 -1769 213 -1767
rect 219 -1763 220 -1761
rect 219 -1769 220 -1767
rect 226 -1763 227 -1761
rect 226 -1769 227 -1767
rect 233 -1763 234 -1761
rect 233 -1769 234 -1767
rect 240 -1763 241 -1761
rect 240 -1769 241 -1767
rect 247 -1763 248 -1761
rect 247 -1769 248 -1767
rect 254 -1763 255 -1761
rect 254 -1769 255 -1767
rect 261 -1763 262 -1761
rect 261 -1769 262 -1767
rect 268 -1763 269 -1761
rect 268 -1769 269 -1767
rect 275 -1763 276 -1761
rect 275 -1769 276 -1767
rect 282 -1763 283 -1761
rect 282 -1769 283 -1767
rect 289 -1763 290 -1761
rect 289 -1769 290 -1767
rect 296 -1763 297 -1761
rect 296 -1769 297 -1767
rect 303 -1763 304 -1761
rect 303 -1769 304 -1767
rect 310 -1763 311 -1761
rect 310 -1769 311 -1767
rect 317 -1763 318 -1761
rect 317 -1769 318 -1767
rect 324 -1763 325 -1761
rect 324 -1769 325 -1767
rect 331 -1763 332 -1761
rect 331 -1769 332 -1767
rect 338 -1763 339 -1761
rect 341 -1763 342 -1761
rect 338 -1769 339 -1767
rect 341 -1769 342 -1767
rect 345 -1763 346 -1761
rect 345 -1769 346 -1767
rect 352 -1763 353 -1761
rect 352 -1769 353 -1767
rect 359 -1763 360 -1761
rect 359 -1769 360 -1767
rect 366 -1763 367 -1761
rect 369 -1763 370 -1761
rect 366 -1769 367 -1767
rect 369 -1769 370 -1767
rect 373 -1763 374 -1761
rect 373 -1769 374 -1767
rect 380 -1763 381 -1761
rect 380 -1769 381 -1767
rect 387 -1763 388 -1761
rect 387 -1769 388 -1767
rect 394 -1763 395 -1761
rect 394 -1769 395 -1767
rect 401 -1763 402 -1761
rect 401 -1769 402 -1767
rect 408 -1763 409 -1761
rect 408 -1769 409 -1767
rect 415 -1763 416 -1761
rect 418 -1763 419 -1761
rect 415 -1769 416 -1767
rect 418 -1769 419 -1767
rect 422 -1763 423 -1761
rect 425 -1763 426 -1761
rect 422 -1769 423 -1767
rect 429 -1763 430 -1761
rect 429 -1769 430 -1767
rect 436 -1763 437 -1761
rect 436 -1769 437 -1767
rect 443 -1763 444 -1761
rect 443 -1769 444 -1767
rect 450 -1763 451 -1761
rect 450 -1769 451 -1767
rect 457 -1763 458 -1761
rect 464 -1763 465 -1761
rect 464 -1769 465 -1767
rect 471 -1763 472 -1761
rect 471 -1769 472 -1767
rect 478 -1763 479 -1761
rect 478 -1769 479 -1767
rect 488 -1763 489 -1761
rect 485 -1769 486 -1767
rect 488 -1769 489 -1767
rect 492 -1763 493 -1761
rect 492 -1769 493 -1767
rect 499 -1763 500 -1761
rect 499 -1769 500 -1767
rect 506 -1763 507 -1761
rect 509 -1763 510 -1761
rect 506 -1769 507 -1767
rect 509 -1769 510 -1767
rect 513 -1763 514 -1761
rect 513 -1769 514 -1767
rect 520 -1763 521 -1761
rect 523 -1763 524 -1761
rect 527 -1763 528 -1761
rect 530 -1763 531 -1761
rect 527 -1769 528 -1767
rect 530 -1769 531 -1767
rect 534 -1763 535 -1761
rect 534 -1769 535 -1767
rect 541 -1763 542 -1761
rect 541 -1769 542 -1767
rect 548 -1763 549 -1761
rect 548 -1769 549 -1767
rect 555 -1763 556 -1761
rect 555 -1769 556 -1767
rect 562 -1763 563 -1761
rect 562 -1769 563 -1767
rect 569 -1763 570 -1761
rect 569 -1769 570 -1767
rect 576 -1763 577 -1761
rect 576 -1769 577 -1767
rect 583 -1763 584 -1761
rect 586 -1763 587 -1761
rect 583 -1769 584 -1767
rect 586 -1769 587 -1767
rect 590 -1763 591 -1761
rect 590 -1769 591 -1767
rect 597 -1763 598 -1761
rect 597 -1769 598 -1767
rect 604 -1763 605 -1761
rect 604 -1769 605 -1767
rect 611 -1763 612 -1761
rect 611 -1769 612 -1767
rect 618 -1763 619 -1761
rect 618 -1769 619 -1767
rect 625 -1763 626 -1761
rect 625 -1769 626 -1767
rect 632 -1763 633 -1761
rect 635 -1763 636 -1761
rect 632 -1769 633 -1767
rect 635 -1769 636 -1767
rect 639 -1763 640 -1761
rect 639 -1769 640 -1767
rect 646 -1763 647 -1761
rect 646 -1769 647 -1767
rect 653 -1763 654 -1761
rect 653 -1769 654 -1767
rect 660 -1763 661 -1761
rect 660 -1769 661 -1767
rect 667 -1763 668 -1761
rect 667 -1769 668 -1767
rect 674 -1763 675 -1761
rect 674 -1769 675 -1767
rect 681 -1763 682 -1761
rect 681 -1769 682 -1767
rect 688 -1763 689 -1761
rect 688 -1769 689 -1767
rect 695 -1763 696 -1761
rect 695 -1769 696 -1767
rect 702 -1763 703 -1761
rect 702 -1769 703 -1767
rect 709 -1763 710 -1761
rect 709 -1769 710 -1767
rect 716 -1763 717 -1761
rect 719 -1763 720 -1761
rect 716 -1769 717 -1767
rect 719 -1769 720 -1767
rect 723 -1763 724 -1761
rect 723 -1769 724 -1767
rect 730 -1763 731 -1761
rect 730 -1769 731 -1767
rect 737 -1763 738 -1761
rect 737 -1769 738 -1767
rect 744 -1763 745 -1761
rect 744 -1769 745 -1767
rect 751 -1763 752 -1761
rect 751 -1769 752 -1767
rect 758 -1763 759 -1761
rect 758 -1769 759 -1767
rect 765 -1763 766 -1761
rect 765 -1769 766 -1767
rect 772 -1763 773 -1761
rect 775 -1763 776 -1761
rect 772 -1769 773 -1767
rect 775 -1769 776 -1767
rect 779 -1763 780 -1761
rect 779 -1769 780 -1767
rect 786 -1763 787 -1761
rect 786 -1769 787 -1767
rect 793 -1763 794 -1761
rect 796 -1763 797 -1761
rect 793 -1769 794 -1767
rect 796 -1769 797 -1767
rect 800 -1763 801 -1761
rect 800 -1769 801 -1767
rect 810 -1763 811 -1761
rect 807 -1769 808 -1767
rect 810 -1769 811 -1767
rect 814 -1763 815 -1761
rect 814 -1769 815 -1767
rect 821 -1763 822 -1761
rect 821 -1769 822 -1767
rect 828 -1763 829 -1761
rect 828 -1769 829 -1767
rect 835 -1763 836 -1761
rect 835 -1769 836 -1767
rect 842 -1763 843 -1761
rect 845 -1763 846 -1761
rect 842 -1769 843 -1767
rect 845 -1769 846 -1767
rect 849 -1763 850 -1761
rect 849 -1769 850 -1767
rect 856 -1763 857 -1761
rect 856 -1769 857 -1767
rect 863 -1763 864 -1761
rect 863 -1769 864 -1767
rect 870 -1763 871 -1761
rect 873 -1763 874 -1761
rect 870 -1769 871 -1767
rect 873 -1769 874 -1767
rect 877 -1763 878 -1761
rect 880 -1763 881 -1761
rect 877 -1769 878 -1767
rect 880 -1769 881 -1767
rect 884 -1763 885 -1761
rect 884 -1769 885 -1767
rect 891 -1763 892 -1761
rect 891 -1769 892 -1767
rect 898 -1763 899 -1761
rect 901 -1763 902 -1761
rect 898 -1769 899 -1767
rect 901 -1769 902 -1767
rect 905 -1763 906 -1761
rect 905 -1769 906 -1767
rect 912 -1763 913 -1761
rect 912 -1769 913 -1767
rect 919 -1763 920 -1761
rect 919 -1769 920 -1767
rect 926 -1763 927 -1761
rect 926 -1769 927 -1767
rect 933 -1763 934 -1761
rect 933 -1769 934 -1767
rect 940 -1763 941 -1761
rect 940 -1769 941 -1767
rect 947 -1763 948 -1761
rect 947 -1769 948 -1767
rect 954 -1763 955 -1761
rect 954 -1769 955 -1767
rect 961 -1763 962 -1761
rect 961 -1769 962 -1767
rect 968 -1763 969 -1761
rect 968 -1769 969 -1767
rect 975 -1763 976 -1761
rect 975 -1769 976 -1767
rect 982 -1763 983 -1761
rect 982 -1769 983 -1767
rect 989 -1763 990 -1761
rect 992 -1763 993 -1761
rect 989 -1769 990 -1767
rect 996 -1763 997 -1761
rect 996 -1769 997 -1767
rect 1003 -1763 1004 -1761
rect 1006 -1763 1007 -1761
rect 1003 -1769 1004 -1767
rect 1006 -1769 1007 -1767
rect 1010 -1763 1011 -1761
rect 1010 -1769 1011 -1767
rect 1017 -1763 1018 -1761
rect 1017 -1769 1018 -1767
rect 1024 -1763 1025 -1761
rect 1024 -1769 1025 -1767
rect 1031 -1763 1032 -1761
rect 1031 -1769 1032 -1767
rect 1038 -1763 1039 -1761
rect 1038 -1769 1039 -1767
rect 1045 -1763 1046 -1761
rect 1045 -1769 1046 -1767
rect 1052 -1763 1053 -1761
rect 1052 -1769 1053 -1767
rect 1059 -1763 1060 -1761
rect 1059 -1769 1060 -1767
rect 1066 -1763 1067 -1761
rect 1066 -1769 1067 -1767
rect 1073 -1763 1074 -1761
rect 1073 -1769 1074 -1767
rect 1080 -1763 1081 -1761
rect 1080 -1769 1081 -1767
rect 1087 -1763 1088 -1761
rect 1087 -1769 1088 -1767
rect 1094 -1763 1095 -1761
rect 1094 -1769 1095 -1767
rect 1101 -1763 1102 -1761
rect 1101 -1769 1102 -1767
rect 1108 -1763 1109 -1761
rect 1108 -1769 1109 -1767
rect 1115 -1763 1116 -1761
rect 1115 -1769 1116 -1767
rect 1122 -1763 1123 -1761
rect 1122 -1769 1123 -1767
rect 1129 -1763 1130 -1761
rect 1129 -1769 1130 -1767
rect 1136 -1763 1137 -1761
rect 1136 -1769 1137 -1767
rect 1143 -1763 1144 -1761
rect 1143 -1769 1144 -1767
rect 1150 -1763 1151 -1761
rect 1150 -1769 1151 -1767
rect 1157 -1763 1158 -1761
rect 1157 -1769 1158 -1767
rect 1164 -1763 1165 -1761
rect 1164 -1769 1165 -1767
rect 1171 -1763 1172 -1761
rect 1171 -1769 1172 -1767
rect 1178 -1763 1179 -1761
rect 1178 -1769 1179 -1767
rect 1185 -1763 1186 -1761
rect 1185 -1769 1186 -1767
rect 1192 -1763 1193 -1761
rect 1192 -1769 1193 -1767
rect 1199 -1763 1200 -1761
rect 1199 -1769 1200 -1767
rect 1206 -1763 1207 -1761
rect 1206 -1769 1207 -1767
rect 1213 -1763 1214 -1761
rect 1213 -1769 1214 -1767
rect 1220 -1763 1221 -1761
rect 1220 -1769 1221 -1767
rect 1227 -1763 1228 -1761
rect 1227 -1769 1228 -1767
rect 1234 -1763 1235 -1761
rect 1234 -1769 1235 -1767
rect 1241 -1763 1242 -1761
rect 1241 -1769 1242 -1767
rect 1248 -1763 1249 -1761
rect 1248 -1769 1249 -1767
rect 1255 -1763 1256 -1761
rect 1255 -1769 1256 -1767
rect 1258 -1769 1259 -1767
rect 1262 -1763 1263 -1761
rect 1262 -1769 1263 -1767
rect 1269 -1763 1270 -1761
rect 1269 -1769 1270 -1767
rect 1276 -1763 1277 -1761
rect 1276 -1769 1277 -1767
rect 1283 -1763 1284 -1761
rect 1283 -1769 1284 -1767
rect 1290 -1763 1291 -1761
rect 1290 -1769 1291 -1767
rect 1297 -1763 1298 -1761
rect 1297 -1769 1298 -1767
rect 1304 -1763 1305 -1761
rect 1304 -1769 1305 -1767
rect 1311 -1763 1312 -1761
rect 1311 -1769 1312 -1767
rect 1318 -1763 1319 -1761
rect 1318 -1769 1319 -1767
rect 1325 -1763 1326 -1761
rect 1325 -1769 1326 -1767
rect 1332 -1763 1333 -1761
rect 1332 -1769 1333 -1767
rect 1339 -1763 1340 -1761
rect 1339 -1769 1340 -1767
rect 1346 -1763 1347 -1761
rect 1346 -1769 1347 -1767
rect 1353 -1763 1354 -1761
rect 1353 -1769 1354 -1767
rect 1360 -1763 1361 -1761
rect 1360 -1769 1361 -1767
rect 1367 -1763 1368 -1761
rect 1370 -1763 1371 -1761
rect 1367 -1769 1368 -1767
rect 1370 -1769 1371 -1767
rect 1374 -1763 1375 -1761
rect 1377 -1763 1378 -1761
rect 1374 -1769 1375 -1767
rect 1377 -1769 1378 -1767
rect 1381 -1763 1382 -1761
rect 1381 -1769 1382 -1767
rect 1388 -1763 1389 -1761
rect 1388 -1769 1389 -1767
rect 1395 -1763 1396 -1761
rect 1395 -1769 1396 -1767
rect 1402 -1763 1403 -1761
rect 1402 -1769 1403 -1767
rect 1409 -1763 1410 -1761
rect 1409 -1769 1410 -1767
rect 1416 -1763 1417 -1761
rect 1416 -1769 1417 -1767
rect 1423 -1763 1424 -1761
rect 1423 -1769 1424 -1767
rect 2 -1860 3 -1858
rect 2 -1866 3 -1864
rect 9 -1860 10 -1858
rect 9 -1866 10 -1864
rect 19 -1860 20 -1858
rect 16 -1866 17 -1864
rect 19 -1866 20 -1864
rect 23 -1860 24 -1858
rect 23 -1866 24 -1864
rect 30 -1860 31 -1858
rect 30 -1866 31 -1864
rect 37 -1860 38 -1858
rect 37 -1866 38 -1864
rect 44 -1860 45 -1858
rect 44 -1866 45 -1864
rect 51 -1860 52 -1858
rect 51 -1866 52 -1864
rect 58 -1860 59 -1858
rect 61 -1860 62 -1858
rect 58 -1866 59 -1864
rect 61 -1866 62 -1864
rect 65 -1860 66 -1858
rect 65 -1866 66 -1864
rect 72 -1860 73 -1858
rect 72 -1866 73 -1864
rect 79 -1860 80 -1858
rect 79 -1866 80 -1864
rect 86 -1860 87 -1858
rect 89 -1860 90 -1858
rect 86 -1866 87 -1864
rect 89 -1866 90 -1864
rect 93 -1860 94 -1858
rect 93 -1866 94 -1864
rect 100 -1860 101 -1858
rect 100 -1866 101 -1864
rect 107 -1860 108 -1858
rect 107 -1866 108 -1864
rect 114 -1860 115 -1858
rect 114 -1866 115 -1864
rect 121 -1860 122 -1858
rect 121 -1866 122 -1864
rect 128 -1860 129 -1858
rect 128 -1866 129 -1864
rect 135 -1860 136 -1858
rect 138 -1860 139 -1858
rect 135 -1866 136 -1864
rect 138 -1866 139 -1864
rect 142 -1860 143 -1858
rect 142 -1866 143 -1864
rect 149 -1860 150 -1858
rect 149 -1866 150 -1864
rect 156 -1860 157 -1858
rect 156 -1866 157 -1864
rect 163 -1860 164 -1858
rect 163 -1866 164 -1864
rect 170 -1860 171 -1858
rect 170 -1866 171 -1864
rect 177 -1860 178 -1858
rect 177 -1866 178 -1864
rect 184 -1860 185 -1858
rect 184 -1866 185 -1864
rect 191 -1860 192 -1858
rect 191 -1866 192 -1864
rect 198 -1860 199 -1858
rect 198 -1866 199 -1864
rect 205 -1860 206 -1858
rect 205 -1866 206 -1864
rect 212 -1860 213 -1858
rect 212 -1866 213 -1864
rect 219 -1860 220 -1858
rect 219 -1866 220 -1864
rect 226 -1860 227 -1858
rect 226 -1866 227 -1864
rect 233 -1860 234 -1858
rect 233 -1866 234 -1864
rect 240 -1860 241 -1858
rect 240 -1866 241 -1864
rect 247 -1860 248 -1858
rect 247 -1866 248 -1864
rect 254 -1860 255 -1858
rect 254 -1866 255 -1864
rect 261 -1860 262 -1858
rect 261 -1866 262 -1864
rect 268 -1860 269 -1858
rect 268 -1866 269 -1864
rect 275 -1860 276 -1858
rect 275 -1866 276 -1864
rect 282 -1860 283 -1858
rect 282 -1866 283 -1864
rect 289 -1860 290 -1858
rect 289 -1866 290 -1864
rect 296 -1860 297 -1858
rect 299 -1860 300 -1858
rect 296 -1866 297 -1864
rect 299 -1866 300 -1864
rect 303 -1860 304 -1858
rect 303 -1866 304 -1864
rect 310 -1860 311 -1858
rect 310 -1866 311 -1864
rect 317 -1860 318 -1858
rect 317 -1866 318 -1864
rect 324 -1860 325 -1858
rect 324 -1866 325 -1864
rect 331 -1860 332 -1858
rect 331 -1866 332 -1864
rect 338 -1860 339 -1858
rect 338 -1866 339 -1864
rect 345 -1860 346 -1858
rect 345 -1866 346 -1864
rect 348 -1866 349 -1864
rect 352 -1860 353 -1858
rect 352 -1866 353 -1864
rect 359 -1860 360 -1858
rect 359 -1866 360 -1864
rect 366 -1860 367 -1858
rect 366 -1866 367 -1864
rect 373 -1860 374 -1858
rect 373 -1866 374 -1864
rect 380 -1860 381 -1858
rect 380 -1866 381 -1864
rect 387 -1860 388 -1858
rect 387 -1866 388 -1864
rect 394 -1860 395 -1858
rect 397 -1860 398 -1858
rect 394 -1866 395 -1864
rect 397 -1866 398 -1864
rect 401 -1860 402 -1858
rect 401 -1866 402 -1864
rect 408 -1860 409 -1858
rect 408 -1866 409 -1864
rect 415 -1860 416 -1858
rect 415 -1866 416 -1864
rect 422 -1860 423 -1858
rect 422 -1866 423 -1864
rect 432 -1860 433 -1858
rect 429 -1866 430 -1864
rect 432 -1866 433 -1864
rect 436 -1860 437 -1858
rect 436 -1866 437 -1864
rect 443 -1860 444 -1858
rect 443 -1866 444 -1864
rect 450 -1860 451 -1858
rect 450 -1866 451 -1864
rect 457 -1866 458 -1864
rect 464 -1860 465 -1858
rect 464 -1866 465 -1864
rect 471 -1860 472 -1858
rect 471 -1866 472 -1864
rect 478 -1860 479 -1858
rect 478 -1866 479 -1864
rect 485 -1860 486 -1858
rect 485 -1866 486 -1864
rect 492 -1860 493 -1858
rect 492 -1866 493 -1864
rect 499 -1860 500 -1858
rect 502 -1860 503 -1858
rect 499 -1866 500 -1864
rect 502 -1866 503 -1864
rect 506 -1860 507 -1858
rect 506 -1866 507 -1864
rect 513 -1860 514 -1858
rect 513 -1866 514 -1864
rect 520 -1860 521 -1858
rect 520 -1866 521 -1864
rect 527 -1860 528 -1858
rect 527 -1866 528 -1864
rect 534 -1860 535 -1858
rect 534 -1866 535 -1864
rect 541 -1860 542 -1858
rect 541 -1866 542 -1864
rect 548 -1860 549 -1858
rect 548 -1866 549 -1864
rect 555 -1860 556 -1858
rect 558 -1860 559 -1858
rect 558 -1866 559 -1864
rect 562 -1860 563 -1858
rect 562 -1866 563 -1864
rect 569 -1860 570 -1858
rect 572 -1860 573 -1858
rect 569 -1866 570 -1864
rect 572 -1866 573 -1864
rect 576 -1860 577 -1858
rect 576 -1866 577 -1864
rect 583 -1860 584 -1858
rect 583 -1866 584 -1864
rect 590 -1860 591 -1858
rect 593 -1860 594 -1858
rect 590 -1866 591 -1864
rect 593 -1866 594 -1864
rect 597 -1860 598 -1858
rect 597 -1866 598 -1864
rect 604 -1860 605 -1858
rect 604 -1866 605 -1864
rect 611 -1860 612 -1858
rect 611 -1866 612 -1864
rect 618 -1860 619 -1858
rect 618 -1866 619 -1864
rect 625 -1860 626 -1858
rect 625 -1866 626 -1864
rect 632 -1860 633 -1858
rect 632 -1866 633 -1864
rect 639 -1860 640 -1858
rect 639 -1866 640 -1864
rect 646 -1860 647 -1858
rect 646 -1866 647 -1864
rect 653 -1860 654 -1858
rect 653 -1866 654 -1864
rect 660 -1860 661 -1858
rect 663 -1860 664 -1858
rect 660 -1866 661 -1864
rect 663 -1866 664 -1864
rect 667 -1860 668 -1858
rect 667 -1866 668 -1864
rect 674 -1860 675 -1858
rect 674 -1866 675 -1864
rect 681 -1860 682 -1858
rect 684 -1860 685 -1858
rect 681 -1866 682 -1864
rect 684 -1866 685 -1864
rect 688 -1860 689 -1858
rect 691 -1860 692 -1858
rect 688 -1866 689 -1864
rect 691 -1866 692 -1864
rect 695 -1860 696 -1858
rect 695 -1866 696 -1864
rect 702 -1860 703 -1858
rect 702 -1866 703 -1864
rect 709 -1860 710 -1858
rect 709 -1866 710 -1864
rect 716 -1860 717 -1858
rect 719 -1860 720 -1858
rect 716 -1866 717 -1864
rect 719 -1866 720 -1864
rect 723 -1860 724 -1858
rect 723 -1866 724 -1864
rect 730 -1860 731 -1858
rect 730 -1866 731 -1864
rect 737 -1860 738 -1858
rect 737 -1866 738 -1864
rect 744 -1860 745 -1858
rect 744 -1866 745 -1864
rect 751 -1860 752 -1858
rect 754 -1860 755 -1858
rect 751 -1866 752 -1864
rect 754 -1866 755 -1864
rect 758 -1860 759 -1858
rect 758 -1866 759 -1864
rect 765 -1860 766 -1858
rect 765 -1866 766 -1864
rect 772 -1860 773 -1858
rect 772 -1866 773 -1864
rect 775 -1866 776 -1864
rect 779 -1860 780 -1858
rect 779 -1866 780 -1864
rect 786 -1860 787 -1858
rect 786 -1866 787 -1864
rect 793 -1860 794 -1858
rect 793 -1866 794 -1864
rect 800 -1860 801 -1858
rect 803 -1860 804 -1858
rect 800 -1866 801 -1864
rect 803 -1866 804 -1864
rect 807 -1860 808 -1858
rect 807 -1866 808 -1864
rect 814 -1860 815 -1858
rect 814 -1866 815 -1864
rect 821 -1860 822 -1858
rect 821 -1866 822 -1864
rect 828 -1860 829 -1858
rect 828 -1866 829 -1864
rect 835 -1860 836 -1858
rect 835 -1866 836 -1864
rect 842 -1860 843 -1858
rect 842 -1866 843 -1864
rect 849 -1860 850 -1858
rect 849 -1866 850 -1864
rect 856 -1860 857 -1858
rect 856 -1866 857 -1864
rect 863 -1860 864 -1858
rect 863 -1866 864 -1864
rect 870 -1860 871 -1858
rect 870 -1866 871 -1864
rect 877 -1860 878 -1858
rect 877 -1866 878 -1864
rect 884 -1860 885 -1858
rect 887 -1860 888 -1858
rect 884 -1866 885 -1864
rect 887 -1866 888 -1864
rect 891 -1860 892 -1858
rect 891 -1866 892 -1864
rect 898 -1860 899 -1858
rect 898 -1866 899 -1864
rect 905 -1860 906 -1858
rect 908 -1860 909 -1858
rect 908 -1866 909 -1864
rect 912 -1860 913 -1858
rect 912 -1866 913 -1864
rect 919 -1860 920 -1858
rect 919 -1866 920 -1864
rect 926 -1860 927 -1858
rect 926 -1866 927 -1864
rect 933 -1860 934 -1858
rect 936 -1860 937 -1858
rect 933 -1866 934 -1864
rect 936 -1866 937 -1864
rect 940 -1860 941 -1858
rect 940 -1866 941 -1864
rect 947 -1860 948 -1858
rect 947 -1866 948 -1864
rect 954 -1860 955 -1858
rect 954 -1866 955 -1864
rect 961 -1860 962 -1858
rect 961 -1866 962 -1864
rect 968 -1860 969 -1858
rect 968 -1866 969 -1864
rect 975 -1860 976 -1858
rect 975 -1866 976 -1864
rect 982 -1860 983 -1858
rect 982 -1866 983 -1864
rect 989 -1860 990 -1858
rect 989 -1866 990 -1864
rect 996 -1860 997 -1858
rect 996 -1866 997 -1864
rect 1003 -1860 1004 -1858
rect 1003 -1866 1004 -1864
rect 1010 -1860 1011 -1858
rect 1010 -1866 1011 -1864
rect 1017 -1860 1018 -1858
rect 1017 -1866 1018 -1864
rect 1024 -1860 1025 -1858
rect 1024 -1866 1025 -1864
rect 1031 -1860 1032 -1858
rect 1031 -1866 1032 -1864
rect 1038 -1860 1039 -1858
rect 1038 -1866 1039 -1864
rect 1045 -1860 1046 -1858
rect 1045 -1866 1046 -1864
rect 1052 -1860 1053 -1858
rect 1052 -1866 1053 -1864
rect 1062 -1860 1063 -1858
rect 1059 -1866 1060 -1864
rect 1062 -1866 1063 -1864
rect 1066 -1860 1067 -1858
rect 1066 -1866 1067 -1864
rect 1073 -1860 1074 -1858
rect 1073 -1866 1074 -1864
rect 1080 -1860 1081 -1858
rect 1080 -1866 1081 -1864
rect 1087 -1860 1088 -1858
rect 1087 -1866 1088 -1864
rect 1094 -1860 1095 -1858
rect 1094 -1866 1095 -1864
rect 1101 -1860 1102 -1858
rect 1101 -1866 1102 -1864
rect 1108 -1860 1109 -1858
rect 1108 -1866 1109 -1864
rect 1115 -1860 1116 -1858
rect 1115 -1866 1116 -1864
rect 1122 -1860 1123 -1858
rect 1122 -1866 1123 -1864
rect 1129 -1860 1130 -1858
rect 1129 -1866 1130 -1864
rect 1136 -1860 1137 -1858
rect 1136 -1866 1137 -1864
rect 1143 -1860 1144 -1858
rect 1143 -1866 1144 -1864
rect 1150 -1860 1151 -1858
rect 1150 -1866 1151 -1864
rect 1157 -1860 1158 -1858
rect 1157 -1866 1158 -1864
rect 1164 -1860 1165 -1858
rect 1164 -1866 1165 -1864
rect 1171 -1860 1172 -1858
rect 1171 -1866 1172 -1864
rect 1178 -1860 1179 -1858
rect 1178 -1866 1179 -1864
rect 1185 -1860 1186 -1858
rect 1185 -1866 1186 -1864
rect 1192 -1860 1193 -1858
rect 1192 -1866 1193 -1864
rect 1199 -1860 1200 -1858
rect 1199 -1866 1200 -1864
rect 1206 -1860 1207 -1858
rect 1206 -1866 1207 -1864
rect 1213 -1860 1214 -1858
rect 1213 -1866 1214 -1864
rect 1220 -1860 1221 -1858
rect 1220 -1866 1221 -1864
rect 1227 -1860 1228 -1858
rect 1227 -1866 1228 -1864
rect 1234 -1860 1235 -1858
rect 1234 -1866 1235 -1864
rect 1241 -1860 1242 -1858
rect 1241 -1866 1242 -1864
rect 1248 -1860 1249 -1858
rect 1248 -1866 1249 -1864
rect 1255 -1860 1256 -1858
rect 1258 -1860 1259 -1858
rect 1255 -1866 1256 -1864
rect 1262 -1860 1263 -1858
rect 1262 -1866 1263 -1864
rect 1269 -1860 1270 -1858
rect 1269 -1866 1270 -1864
rect 1276 -1860 1277 -1858
rect 1276 -1866 1277 -1864
rect 1283 -1860 1284 -1858
rect 1283 -1866 1284 -1864
rect 1290 -1860 1291 -1858
rect 1290 -1866 1291 -1864
rect 1297 -1860 1298 -1858
rect 1297 -1866 1298 -1864
rect 1304 -1860 1305 -1858
rect 1304 -1866 1305 -1864
rect 1311 -1860 1312 -1858
rect 1311 -1866 1312 -1864
rect 1318 -1860 1319 -1858
rect 1318 -1866 1319 -1864
rect 1325 -1860 1326 -1858
rect 1325 -1866 1326 -1864
rect 1332 -1860 1333 -1858
rect 1332 -1866 1333 -1864
rect 1339 -1860 1340 -1858
rect 1339 -1866 1340 -1864
rect 1346 -1860 1347 -1858
rect 1346 -1866 1347 -1864
rect 1353 -1860 1354 -1858
rect 1353 -1866 1354 -1864
rect 1360 -1860 1361 -1858
rect 1360 -1866 1361 -1864
rect 1367 -1860 1368 -1858
rect 1367 -1866 1368 -1864
rect 1374 -1860 1375 -1858
rect 1374 -1866 1375 -1864
rect 1381 -1860 1382 -1858
rect 1381 -1866 1382 -1864
rect 1388 -1860 1389 -1858
rect 1388 -1866 1389 -1864
rect 1395 -1860 1396 -1858
rect 1395 -1866 1396 -1864
rect 1398 -1866 1399 -1864
rect 1402 -1860 1403 -1858
rect 1402 -1866 1403 -1864
rect 1409 -1860 1410 -1858
rect 1409 -1866 1410 -1864
rect 1416 -1860 1417 -1858
rect 1416 -1866 1417 -1864
rect 1423 -1860 1424 -1858
rect 1423 -1866 1424 -1864
rect 1430 -1860 1431 -1858
rect 1430 -1866 1431 -1864
rect 2 -1987 3 -1985
rect 2 -1993 3 -1991
rect 9 -1987 10 -1985
rect 9 -1993 10 -1991
rect 16 -1987 17 -1985
rect 16 -1993 17 -1991
rect 23 -1987 24 -1985
rect 26 -1987 27 -1985
rect 23 -1993 24 -1991
rect 30 -1987 31 -1985
rect 30 -1993 31 -1991
rect 37 -1987 38 -1985
rect 40 -1987 41 -1985
rect 37 -1993 38 -1991
rect 40 -1993 41 -1991
rect 44 -1987 45 -1985
rect 44 -1993 45 -1991
rect 51 -1987 52 -1985
rect 51 -1993 52 -1991
rect 58 -1987 59 -1985
rect 58 -1993 59 -1991
rect 65 -1987 66 -1985
rect 68 -1987 69 -1985
rect 65 -1993 66 -1991
rect 68 -1993 69 -1991
rect 72 -1987 73 -1985
rect 75 -1987 76 -1985
rect 72 -1993 73 -1991
rect 75 -1993 76 -1991
rect 79 -1987 80 -1985
rect 79 -1993 80 -1991
rect 86 -1987 87 -1985
rect 86 -1993 87 -1991
rect 93 -1987 94 -1985
rect 93 -1993 94 -1991
rect 100 -1987 101 -1985
rect 100 -1993 101 -1991
rect 107 -1987 108 -1985
rect 107 -1993 108 -1991
rect 114 -1987 115 -1985
rect 114 -1993 115 -1991
rect 121 -1987 122 -1985
rect 121 -1993 122 -1991
rect 128 -1987 129 -1985
rect 128 -1993 129 -1991
rect 135 -1987 136 -1985
rect 135 -1993 136 -1991
rect 142 -1987 143 -1985
rect 142 -1993 143 -1991
rect 149 -1987 150 -1985
rect 149 -1993 150 -1991
rect 156 -1987 157 -1985
rect 156 -1993 157 -1991
rect 163 -1987 164 -1985
rect 163 -1993 164 -1991
rect 170 -1987 171 -1985
rect 173 -1987 174 -1985
rect 170 -1993 171 -1991
rect 173 -1993 174 -1991
rect 177 -1987 178 -1985
rect 177 -1993 178 -1991
rect 184 -1987 185 -1985
rect 184 -1993 185 -1991
rect 191 -1987 192 -1985
rect 191 -1993 192 -1991
rect 198 -1987 199 -1985
rect 198 -1993 199 -1991
rect 205 -1987 206 -1985
rect 205 -1993 206 -1991
rect 212 -1987 213 -1985
rect 212 -1993 213 -1991
rect 219 -1987 220 -1985
rect 219 -1993 220 -1991
rect 226 -1987 227 -1985
rect 229 -1987 230 -1985
rect 226 -1993 227 -1991
rect 229 -1993 230 -1991
rect 233 -1987 234 -1985
rect 233 -1993 234 -1991
rect 240 -1987 241 -1985
rect 240 -1993 241 -1991
rect 247 -1987 248 -1985
rect 247 -1993 248 -1991
rect 254 -1987 255 -1985
rect 254 -1993 255 -1991
rect 261 -1987 262 -1985
rect 261 -1993 262 -1991
rect 268 -1987 269 -1985
rect 268 -1993 269 -1991
rect 275 -1987 276 -1985
rect 275 -1993 276 -1991
rect 282 -1987 283 -1985
rect 282 -1993 283 -1991
rect 289 -1987 290 -1985
rect 289 -1993 290 -1991
rect 296 -1987 297 -1985
rect 296 -1993 297 -1991
rect 303 -1987 304 -1985
rect 303 -1993 304 -1991
rect 310 -1987 311 -1985
rect 310 -1993 311 -1991
rect 317 -1987 318 -1985
rect 317 -1993 318 -1991
rect 324 -1987 325 -1985
rect 324 -1993 325 -1991
rect 331 -1987 332 -1985
rect 331 -1993 332 -1991
rect 338 -1987 339 -1985
rect 338 -1993 339 -1991
rect 345 -1987 346 -1985
rect 345 -1993 346 -1991
rect 352 -1987 353 -1985
rect 355 -1987 356 -1985
rect 352 -1993 353 -1991
rect 355 -1993 356 -1991
rect 359 -1987 360 -1985
rect 359 -1993 360 -1991
rect 366 -1987 367 -1985
rect 366 -1993 367 -1991
rect 373 -1987 374 -1985
rect 373 -1993 374 -1991
rect 376 -1993 377 -1991
rect 380 -1987 381 -1985
rect 380 -1993 381 -1991
rect 387 -1987 388 -1985
rect 387 -1993 388 -1991
rect 394 -1987 395 -1985
rect 394 -1993 395 -1991
rect 401 -1987 402 -1985
rect 401 -1993 402 -1991
rect 408 -1987 409 -1985
rect 411 -1987 412 -1985
rect 408 -1993 409 -1991
rect 411 -1993 412 -1991
rect 415 -1987 416 -1985
rect 415 -1993 416 -1991
rect 422 -1987 423 -1985
rect 422 -1993 423 -1991
rect 429 -1987 430 -1985
rect 429 -1993 430 -1991
rect 436 -1987 437 -1985
rect 436 -1993 437 -1991
rect 443 -1987 444 -1985
rect 443 -1993 444 -1991
rect 450 -1987 451 -1985
rect 450 -1993 451 -1991
rect 457 -1987 458 -1985
rect 457 -1993 458 -1991
rect 464 -1987 465 -1985
rect 464 -1993 465 -1991
rect 471 -1987 472 -1985
rect 471 -1993 472 -1991
rect 478 -1987 479 -1985
rect 478 -1993 479 -1991
rect 485 -1987 486 -1985
rect 485 -1993 486 -1991
rect 492 -1987 493 -1985
rect 492 -1993 493 -1991
rect 499 -1987 500 -1985
rect 499 -1993 500 -1991
rect 506 -1987 507 -1985
rect 509 -1987 510 -1985
rect 506 -1993 507 -1991
rect 509 -1993 510 -1991
rect 513 -1987 514 -1985
rect 516 -1987 517 -1985
rect 513 -1993 514 -1991
rect 516 -1993 517 -1991
rect 520 -1987 521 -1985
rect 523 -1987 524 -1985
rect 520 -1993 521 -1991
rect 523 -1993 524 -1991
rect 527 -1987 528 -1985
rect 527 -1993 528 -1991
rect 534 -1987 535 -1985
rect 534 -1993 535 -1991
rect 541 -1987 542 -1985
rect 541 -1993 542 -1991
rect 548 -1987 549 -1985
rect 548 -1993 549 -1991
rect 555 -1987 556 -1985
rect 555 -1993 556 -1991
rect 562 -1987 563 -1985
rect 565 -1987 566 -1985
rect 562 -1993 563 -1991
rect 569 -1987 570 -1985
rect 569 -1993 570 -1991
rect 576 -1987 577 -1985
rect 579 -1987 580 -1985
rect 576 -1993 577 -1991
rect 579 -1993 580 -1991
rect 583 -1987 584 -1985
rect 583 -1993 584 -1991
rect 586 -1993 587 -1991
rect 590 -1987 591 -1985
rect 590 -1993 591 -1991
rect 597 -1987 598 -1985
rect 597 -1993 598 -1991
rect 604 -1987 605 -1985
rect 604 -1993 605 -1991
rect 611 -1987 612 -1985
rect 614 -1987 615 -1985
rect 611 -1993 612 -1991
rect 614 -1993 615 -1991
rect 618 -1987 619 -1985
rect 618 -1993 619 -1991
rect 625 -1987 626 -1985
rect 625 -1993 626 -1991
rect 632 -1987 633 -1985
rect 632 -1993 633 -1991
rect 639 -1987 640 -1985
rect 642 -1987 643 -1985
rect 639 -1993 640 -1991
rect 642 -1993 643 -1991
rect 646 -1987 647 -1985
rect 646 -1993 647 -1991
rect 653 -1987 654 -1985
rect 653 -1993 654 -1991
rect 660 -1987 661 -1985
rect 663 -1987 664 -1985
rect 660 -1993 661 -1991
rect 663 -1993 664 -1991
rect 667 -1987 668 -1985
rect 667 -1993 668 -1991
rect 674 -1987 675 -1985
rect 674 -1993 675 -1991
rect 681 -1987 682 -1985
rect 681 -1993 682 -1991
rect 688 -1987 689 -1985
rect 688 -1993 689 -1991
rect 695 -1987 696 -1985
rect 695 -1993 696 -1991
rect 702 -1987 703 -1985
rect 705 -1987 706 -1985
rect 702 -1993 703 -1991
rect 705 -1993 706 -1991
rect 709 -1987 710 -1985
rect 709 -1993 710 -1991
rect 716 -1987 717 -1985
rect 716 -1993 717 -1991
rect 723 -1987 724 -1985
rect 726 -1987 727 -1985
rect 723 -1993 724 -1991
rect 726 -1993 727 -1991
rect 730 -1987 731 -1985
rect 730 -1993 731 -1991
rect 737 -1987 738 -1985
rect 737 -1993 738 -1991
rect 744 -1987 745 -1985
rect 744 -1993 745 -1991
rect 751 -1987 752 -1985
rect 754 -1987 755 -1985
rect 751 -1993 752 -1991
rect 754 -1993 755 -1991
rect 758 -1987 759 -1985
rect 758 -1993 759 -1991
rect 765 -1987 766 -1985
rect 765 -1993 766 -1991
rect 772 -1987 773 -1985
rect 772 -1993 773 -1991
rect 779 -1987 780 -1985
rect 782 -1987 783 -1985
rect 779 -1993 780 -1991
rect 782 -1993 783 -1991
rect 786 -1987 787 -1985
rect 786 -1993 787 -1991
rect 793 -1987 794 -1985
rect 793 -1993 794 -1991
rect 800 -1987 801 -1985
rect 800 -1993 801 -1991
rect 807 -1987 808 -1985
rect 807 -1993 808 -1991
rect 810 -1993 811 -1991
rect 814 -1987 815 -1985
rect 814 -1993 815 -1991
rect 821 -1987 822 -1985
rect 821 -1993 822 -1991
rect 828 -1987 829 -1985
rect 828 -1993 829 -1991
rect 835 -1987 836 -1985
rect 835 -1993 836 -1991
rect 842 -1987 843 -1985
rect 842 -1993 843 -1991
rect 852 -1987 853 -1985
rect 849 -1993 850 -1991
rect 852 -1993 853 -1991
rect 856 -1987 857 -1985
rect 856 -1993 857 -1991
rect 863 -1987 864 -1985
rect 863 -1993 864 -1991
rect 870 -1987 871 -1985
rect 870 -1993 871 -1991
rect 877 -1987 878 -1985
rect 877 -1993 878 -1991
rect 884 -1987 885 -1985
rect 884 -1993 885 -1991
rect 891 -1987 892 -1985
rect 891 -1993 892 -1991
rect 898 -1987 899 -1985
rect 898 -1993 899 -1991
rect 905 -1987 906 -1985
rect 905 -1993 906 -1991
rect 912 -1987 913 -1985
rect 912 -1993 913 -1991
rect 919 -1987 920 -1985
rect 919 -1993 920 -1991
rect 926 -1987 927 -1985
rect 926 -1993 927 -1991
rect 933 -1987 934 -1985
rect 933 -1993 934 -1991
rect 940 -1987 941 -1985
rect 940 -1993 941 -1991
rect 947 -1987 948 -1985
rect 947 -1993 948 -1991
rect 954 -1987 955 -1985
rect 954 -1993 955 -1991
rect 961 -1987 962 -1985
rect 961 -1993 962 -1991
rect 968 -1987 969 -1985
rect 968 -1993 969 -1991
rect 975 -1987 976 -1985
rect 975 -1993 976 -1991
rect 982 -1987 983 -1985
rect 982 -1993 983 -1991
rect 989 -1987 990 -1985
rect 989 -1993 990 -1991
rect 996 -1987 997 -1985
rect 996 -1993 997 -1991
rect 1003 -1987 1004 -1985
rect 1003 -1993 1004 -1991
rect 1010 -1987 1011 -1985
rect 1010 -1993 1011 -1991
rect 1017 -1987 1018 -1985
rect 1017 -1993 1018 -1991
rect 1024 -1987 1025 -1985
rect 1024 -1993 1025 -1991
rect 1031 -1987 1032 -1985
rect 1031 -1993 1032 -1991
rect 1038 -1987 1039 -1985
rect 1038 -1993 1039 -1991
rect 1045 -1987 1046 -1985
rect 1045 -1993 1046 -1991
rect 1052 -1987 1053 -1985
rect 1052 -1993 1053 -1991
rect 1059 -1987 1060 -1985
rect 1059 -1993 1060 -1991
rect 1066 -1987 1067 -1985
rect 1066 -1993 1067 -1991
rect 1073 -1987 1074 -1985
rect 1073 -1993 1074 -1991
rect 1080 -1987 1081 -1985
rect 1080 -1993 1081 -1991
rect 1087 -1987 1088 -1985
rect 1087 -1993 1088 -1991
rect 1094 -1987 1095 -1985
rect 1094 -1993 1095 -1991
rect 1101 -1987 1102 -1985
rect 1101 -1993 1102 -1991
rect 1108 -1987 1109 -1985
rect 1108 -1993 1109 -1991
rect 1115 -1987 1116 -1985
rect 1115 -1993 1116 -1991
rect 1122 -1987 1123 -1985
rect 1122 -1993 1123 -1991
rect 1129 -1987 1130 -1985
rect 1129 -1993 1130 -1991
rect 1136 -1987 1137 -1985
rect 1136 -1993 1137 -1991
rect 1143 -1987 1144 -1985
rect 1143 -1993 1144 -1991
rect 1150 -1987 1151 -1985
rect 1150 -1993 1151 -1991
rect 1157 -1987 1158 -1985
rect 1157 -1993 1158 -1991
rect 1164 -1987 1165 -1985
rect 1164 -1993 1165 -1991
rect 1171 -1987 1172 -1985
rect 1171 -1993 1172 -1991
rect 1178 -1987 1179 -1985
rect 1178 -1993 1179 -1991
rect 1185 -1987 1186 -1985
rect 1185 -1993 1186 -1991
rect 1192 -1987 1193 -1985
rect 1192 -1993 1193 -1991
rect 1199 -1987 1200 -1985
rect 1199 -1993 1200 -1991
rect 1206 -1987 1207 -1985
rect 1206 -1993 1207 -1991
rect 1213 -1987 1214 -1985
rect 1213 -1993 1214 -1991
rect 1220 -1987 1221 -1985
rect 1220 -1993 1221 -1991
rect 1227 -1987 1228 -1985
rect 1227 -1993 1228 -1991
rect 1234 -1987 1235 -1985
rect 1234 -1993 1235 -1991
rect 1241 -1987 1242 -1985
rect 1241 -1993 1242 -1991
rect 1248 -1987 1249 -1985
rect 1248 -1993 1249 -1991
rect 1255 -1987 1256 -1985
rect 1255 -1993 1256 -1991
rect 1262 -1987 1263 -1985
rect 1262 -1993 1263 -1991
rect 1269 -1987 1270 -1985
rect 1269 -1993 1270 -1991
rect 1276 -1987 1277 -1985
rect 1276 -1993 1277 -1991
rect 1283 -1987 1284 -1985
rect 1283 -1993 1284 -1991
rect 1290 -1987 1291 -1985
rect 1290 -1993 1291 -1991
rect 1297 -1987 1298 -1985
rect 1297 -1993 1298 -1991
rect 1304 -1987 1305 -1985
rect 1304 -1993 1305 -1991
rect 1311 -1987 1312 -1985
rect 1311 -1993 1312 -1991
rect 1318 -1987 1319 -1985
rect 1318 -1993 1319 -1991
rect 1325 -1987 1326 -1985
rect 1325 -1993 1326 -1991
rect 1332 -1987 1333 -1985
rect 1332 -1993 1333 -1991
rect 1339 -1987 1340 -1985
rect 1339 -1993 1340 -1991
rect 1346 -1987 1347 -1985
rect 1346 -1993 1347 -1991
rect 1353 -1987 1354 -1985
rect 1353 -1993 1354 -1991
rect 1360 -1987 1361 -1985
rect 1360 -1993 1361 -1991
rect 1367 -1987 1368 -1985
rect 1367 -1993 1368 -1991
rect 1374 -1987 1375 -1985
rect 1374 -1993 1375 -1991
rect 1381 -1987 1382 -1985
rect 1381 -1993 1382 -1991
rect 1388 -1987 1389 -1985
rect 1388 -1993 1389 -1991
rect 1395 -1987 1396 -1985
rect 1395 -1993 1396 -1991
rect 1402 -1987 1403 -1985
rect 1402 -1993 1403 -1991
rect 2 -2106 3 -2104
rect 5 -2106 6 -2104
rect 5 -2112 6 -2110
rect 9 -2106 10 -2104
rect 9 -2112 10 -2110
rect 16 -2106 17 -2104
rect 16 -2112 17 -2110
rect 23 -2106 24 -2104
rect 23 -2112 24 -2110
rect 30 -2106 31 -2104
rect 30 -2112 31 -2110
rect 37 -2106 38 -2104
rect 37 -2112 38 -2110
rect 44 -2106 45 -2104
rect 44 -2112 45 -2110
rect 51 -2106 52 -2104
rect 51 -2112 52 -2110
rect 58 -2106 59 -2104
rect 58 -2112 59 -2110
rect 65 -2106 66 -2104
rect 65 -2112 66 -2110
rect 72 -2106 73 -2104
rect 72 -2112 73 -2110
rect 79 -2106 80 -2104
rect 79 -2112 80 -2110
rect 86 -2106 87 -2104
rect 86 -2112 87 -2110
rect 93 -2106 94 -2104
rect 96 -2106 97 -2104
rect 93 -2112 94 -2110
rect 100 -2106 101 -2104
rect 100 -2112 101 -2110
rect 107 -2106 108 -2104
rect 110 -2106 111 -2104
rect 107 -2112 108 -2110
rect 110 -2112 111 -2110
rect 114 -2106 115 -2104
rect 114 -2112 115 -2110
rect 121 -2106 122 -2104
rect 121 -2112 122 -2110
rect 128 -2106 129 -2104
rect 131 -2106 132 -2104
rect 128 -2112 129 -2110
rect 131 -2112 132 -2110
rect 135 -2106 136 -2104
rect 135 -2112 136 -2110
rect 142 -2106 143 -2104
rect 142 -2112 143 -2110
rect 149 -2106 150 -2104
rect 149 -2112 150 -2110
rect 156 -2106 157 -2104
rect 156 -2112 157 -2110
rect 163 -2106 164 -2104
rect 166 -2106 167 -2104
rect 170 -2106 171 -2104
rect 173 -2106 174 -2104
rect 170 -2112 171 -2110
rect 177 -2106 178 -2104
rect 177 -2112 178 -2110
rect 184 -2106 185 -2104
rect 184 -2112 185 -2110
rect 191 -2106 192 -2104
rect 191 -2112 192 -2110
rect 198 -2106 199 -2104
rect 198 -2112 199 -2110
rect 205 -2106 206 -2104
rect 205 -2112 206 -2110
rect 212 -2106 213 -2104
rect 212 -2112 213 -2110
rect 219 -2106 220 -2104
rect 219 -2112 220 -2110
rect 226 -2106 227 -2104
rect 226 -2112 227 -2110
rect 233 -2106 234 -2104
rect 240 -2106 241 -2104
rect 240 -2112 241 -2110
rect 247 -2106 248 -2104
rect 247 -2112 248 -2110
rect 254 -2106 255 -2104
rect 254 -2112 255 -2110
rect 261 -2106 262 -2104
rect 261 -2112 262 -2110
rect 268 -2106 269 -2104
rect 268 -2112 269 -2110
rect 275 -2106 276 -2104
rect 275 -2112 276 -2110
rect 282 -2106 283 -2104
rect 282 -2112 283 -2110
rect 289 -2106 290 -2104
rect 289 -2112 290 -2110
rect 296 -2106 297 -2104
rect 296 -2112 297 -2110
rect 303 -2106 304 -2104
rect 303 -2112 304 -2110
rect 310 -2106 311 -2104
rect 310 -2112 311 -2110
rect 317 -2106 318 -2104
rect 320 -2106 321 -2104
rect 317 -2112 318 -2110
rect 320 -2112 321 -2110
rect 324 -2106 325 -2104
rect 324 -2112 325 -2110
rect 331 -2106 332 -2104
rect 334 -2106 335 -2104
rect 331 -2112 332 -2110
rect 334 -2112 335 -2110
rect 338 -2106 339 -2104
rect 338 -2112 339 -2110
rect 345 -2106 346 -2104
rect 348 -2112 349 -2110
rect 352 -2106 353 -2104
rect 352 -2112 353 -2110
rect 359 -2106 360 -2104
rect 359 -2112 360 -2110
rect 366 -2106 367 -2104
rect 366 -2112 367 -2110
rect 373 -2106 374 -2104
rect 373 -2112 374 -2110
rect 380 -2106 381 -2104
rect 380 -2112 381 -2110
rect 387 -2106 388 -2104
rect 387 -2112 388 -2110
rect 394 -2106 395 -2104
rect 394 -2112 395 -2110
rect 401 -2106 402 -2104
rect 401 -2112 402 -2110
rect 408 -2106 409 -2104
rect 408 -2112 409 -2110
rect 415 -2106 416 -2104
rect 415 -2112 416 -2110
rect 422 -2106 423 -2104
rect 422 -2112 423 -2110
rect 429 -2106 430 -2104
rect 429 -2112 430 -2110
rect 436 -2106 437 -2104
rect 436 -2112 437 -2110
rect 443 -2106 444 -2104
rect 443 -2112 444 -2110
rect 450 -2106 451 -2104
rect 453 -2106 454 -2104
rect 450 -2112 451 -2110
rect 453 -2112 454 -2110
rect 457 -2106 458 -2104
rect 457 -2112 458 -2110
rect 464 -2106 465 -2104
rect 464 -2112 465 -2110
rect 471 -2106 472 -2104
rect 471 -2112 472 -2110
rect 478 -2106 479 -2104
rect 478 -2112 479 -2110
rect 485 -2106 486 -2104
rect 488 -2106 489 -2104
rect 485 -2112 486 -2110
rect 488 -2112 489 -2110
rect 492 -2106 493 -2104
rect 492 -2112 493 -2110
rect 499 -2106 500 -2104
rect 502 -2106 503 -2104
rect 499 -2112 500 -2110
rect 502 -2112 503 -2110
rect 506 -2106 507 -2104
rect 506 -2112 507 -2110
rect 513 -2106 514 -2104
rect 513 -2112 514 -2110
rect 520 -2106 521 -2104
rect 520 -2112 521 -2110
rect 527 -2106 528 -2104
rect 527 -2112 528 -2110
rect 534 -2106 535 -2104
rect 534 -2112 535 -2110
rect 541 -2106 542 -2104
rect 541 -2112 542 -2110
rect 548 -2106 549 -2104
rect 548 -2112 549 -2110
rect 555 -2106 556 -2104
rect 555 -2112 556 -2110
rect 562 -2106 563 -2104
rect 562 -2112 563 -2110
rect 569 -2106 570 -2104
rect 569 -2112 570 -2110
rect 576 -2106 577 -2104
rect 579 -2106 580 -2104
rect 576 -2112 577 -2110
rect 579 -2112 580 -2110
rect 583 -2106 584 -2104
rect 583 -2112 584 -2110
rect 590 -2106 591 -2104
rect 590 -2112 591 -2110
rect 597 -2106 598 -2104
rect 597 -2112 598 -2110
rect 604 -2106 605 -2104
rect 604 -2112 605 -2110
rect 611 -2106 612 -2104
rect 611 -2112 612 -2110
rect 618 -2106 619 -2104
rect 621 -2106 622 -2104
rect 618 -2112 619 -2110
rect 621 -2112 622 -2110
rect 625 -2106 626 -2104
rect 625 -2112 626 -2110
rect 632 -2106 633 -2104
rect 632 -2112 633 -2110
rect 639 -2106 640 -2104
rect 639 -2112 640 -2110
rect 646 -2106 647 -2104
rect 646 -2112 647 -2110
rect 653 -2106 654 -2104
rect 653 -2112 654 -2110
rect 660 -2106 661 -2104
rect 660 -2112 661 -2110
rect 667 -2106 668 -2104
rect 670 -2106 671 -2104
rect 667 -2112 668 -2110
rect 674 -2106 675 -2104
rect 674 -2112 675 -2110
rect 681 -2106 682 -2104
rect 681 -2112 682 -2110
rect 688 -2106 689 -2104
rect 691 -2106 692 -2104
rect 688 -2112 689 -2110
rect 691 -2112 692 -2110
rect 695 -2106 696 -2104
rect 695 -2112 696 -2110
rect 702 -2106 703 -2104
rect 702 -2112 703 -2110
rect 709 -2106 710 -2104
rect 709 -2112 710 -2110
rect 716 -2106 717 -2104
rect 716 -2112 717 -2110
rect 723 -2106 724 -2104
rect 723 -2112 724 -2110
rect 730 -2106 731 -2104
rect 730 -2112 731 -2110
rect 737 -2106 738 -2104
rect 737 -2112 738 -2110
rect 744 -2106 745 -2104
rect 744 -2112 745 -2110
rect 751 -2106 752 -2104
rect 751 -2112 752 -2110
rect 758 -2106 759 -2104
rect 758 -2112 759 -2110
rect 765 -2106 766 -2104
rect 765 -2112 766 -2110
rect 768 -2112 769 -2110
rect 772 -2106 773 -2104
rect 772 -2112 773 -2110
rect 779 -2106 780 -2104
rect 782 -2106 783 -2104
rect 782 -2112 783 -2110
rect 786 -2106 787 -2104
rect 786 -2112 787 -2110
rect 793 -2106 794 -2104
rect 793 -2112 794 -2110
rect 800 -2106 801 -2104
rect 800 -2112 801 -2110
rect 807 -2106 808 -2104
rect 807 -2112 808 -2110
rect 814 -2106 815 -2104
rect 817 -2106 818 -2104
rect 814 -2112 815 -2110
rect 817 -2112 818 -2110
rect 821 -2106 822 -2104
rect 824 -2106 825 -2104
rect 824 -2112 825 -2110
rect 828 -2106 829 -2104
rect 828 -2112 829 -2110
rect 835 -2106 836 -2104
rect 835 -2112 836 -2110
rect 842 -2106 843 -2104
rect 842 -2112 843 -2110
rect 849 -2106 850 -2104
rect 849 -2112 850 -2110
rect 856 -2106 857 -2104
rect 856 -2112 857 -2110
rect 863 -2106 864 -2104
rect 863 -2112 864 -2110
rect 870 -2106 871 -2104
rect 870 -2112 871 -2110
rect 877 -2106 878 -2104
rect 877 -2112 878 -2110
rect 884 -2106 885 -2104
rect 884 -2112 885 -2110
rect 894 -2106 895 -2104
rect 891 -2112 892 -2110
rect 894 -2112 895 -2110
rect 898 -2106 899 -2104
rect 898 -2112 899 -2110
rect 905 -2106 906 -2104
rect 905 -2112 906 -2110
rect 912 -2106 913 -2104
rect 912 -2112 913 -2110
rect 919 -2106 920 -2104
rect 919 -2112 920 -2110
rect 926 -2106 927 -2104
rect 926 -2112 927 -2110
rect 933 -2106 934 -2104
rect 933 -2112 934 -2110
rect 940 -2106 941 -2104
rect 940 -2112 941 -2110
rect 947 -2106 948 -2104
rect 947 -2112 948 -2110
rect 954 -2106 955 -2104
rect 954 -2112 955 -2110
rect 961 -2106 962 -2104
rect 961 -2112 962 -2110
rect 968 -2106 969 -2104
rect 971 -2106 972 -2104
rect 968 -2112 969 -2110
rect 971 -2112 972 -2110
rect 975 -2106 976 -2104
rect 975 -2112 976 -2110
rect 982 -2106 983 -2104
rect 982 -2112 983 -2110
rect 992 -2106 993 -2104
rect 989 -2112 990 -2110
rect 992 -2112 993 -2110
rect 996 -2106 997 -2104
rect 996 -2112 997 -2110
rect 1003 -2106 1004 -2104
rect 1003 -2112 1004 -2110
rect 1010 -2106 1011 -2104
rect 1010 -2112 1011 -2110
rect 1017 -2106 1018 -2104
rect 1017 -2112 1018 -2110
rect 1024 -2106 1025 -2104
rect 1024 -2112 1025 -2110
rect 1031 -2106 1032 -2104
rect 1031 -2112 1032 -2110
rect 1038 -2106 1039 -2104
rect 1038 -2112 1039 -2110
rect 1045 -2106 1046 -2104
rect 1045 -2112 1046 -2110
rect 1052 -2106 1053 -2104
rect 1052 -2112 1053 -2110
rect 1059 -2106 1060 -2104
rect 1059 -2112 1060 -2110
rect 1066 -2106 1067 -2104
rect 1066 -2112 1067 -2110
rect 1073 -2106 1074 -2104
rect 1073 -2112 1074 -2110
rect 1080 -2106 1081 -2104
rect 1080 -2112 1081 -2110
rect 1087 -2106 1088 -2104
rect 1087 -2112 1088 -2110
rect 1094 -2106 1095 -2104
rect 1094 -2112 1095 -2110
rect 1101 -2106 1102 -2104
rect 1101 -2112 1102 -2110
rect 1108 -2106 1109 -2104
rect 1108 -2112 1109 -2110
rect 1115 -2106 1116 -2104
rect 1115 -2112 1116 -2110
rect 1118 -2112 1119 -2110
rect 1122 -2106 1123 -2104
rect 1122 -2112 1123 -2110
rect 1129 -2106 1130 -2104
rect 1129 -2112 1130 -2110
rect 1139 -2106 1140 -2104
rect 1136 -2112 1137 -2110
rect 1139 -2112 1140 -2110
rect 1143 -2106 1144 -2104
rect 1143 -2112 1144 -2110
rect 1150 -2106 1151 -2104
rect 1150 -2112 1151 -2110
rect 1157 -2106 1158 -2104
rect 1157 -2112 1158 -2110
rect 1164 -2106 1165 -2104
rect 1164 -2112 1165 -2110
rect 1171 -2106 1172 -2104
rect 1171 -2112 1172 -2110
rect 1178 -2106 1179 -2104
rect 1178 -2112 1179 -2110
rect 1185 -2106 1186 -2104
rect 1185 -2112 1186 -2110
rect 1192 -2106 1193 -2104
rect 1192 -2112 1193 -2110
rect 1199 -2106 1200 -2104
rect 1199 -2112 1200 -2110
rect 1206 -2106 1207 -2104
rect 1206 -2112 1207 -2110
rect 1213 -2106 1214 -2104
rect 1213 -2112 1214 -2110
rect 1220 -2106 1221 -2104
rect 1220 -2112 1221 -2110
rect 1227 -2106 1228 -2104
rect 1227 -2112 1228 -2110
rect 1234 -2106 1235 -2104
rect 1234 -2112 1235 -2110
rect 1241 -2106 1242 -2104
rect 1241 -2112 1242 -2110
rect 1248 -2106 1249 -2104
rect 1248 -2112 1249 -2110
rect 1255 -2106 1256 -2104
rect 1255 -2112 1256 -2110
rect 1262 -2106 1263 -2104
rect 1262 -2112 1263 -2110
rect 1269 -2106 1270 -2104
rect 1269 -2112 1270 -2110
rect 1276 -2106 1277 -2104
rect 1276 -2112 1277 -2110
rect 1283 -2106 1284 -2104
rect 1283 -2112 1284 -2110
rect 1290 -2106 1291 -2104
rect 1290 -2112 1291 -2110
rect 1297 -2106 1298 -2104
rect 1297 -2112 1298 -2110
rect 1304 -2106 1305 -2104
rect 1304 -2112 1305 -2110
rect 1311 -2106 1312 -2104
rect 1311 -2112 1312 -2110
rect 1318 -2106 1319 -2104
rect 1318 -2112 1319 -2110
rect 1325 -2106 1326 -2104
rect 1325 -2112 1326 -2110
rect 2 -2239 3 -2237
rect 2 -2245 3 -2243
rect 9 -2239 10 -2237
rect 9 -2245 10 -2243
rect 16 -2239 17 -2237
rect 16 -2245 17 -2243
rect 23 -2239 24 -2237
rect 26 -2239 27 -2237
rect 23 -2245 24 -2243
rect 30 -2245 31 -2243
rect 33 -2245 34 -2243
rect 37 -2239 38 -2237
rect 40 -2239 41 -2237
rect 37 -2245 38 -2243
rect 40 -2245 41 -2243
rect 44 -2239 45 -2237
rect 44 -2245 45 -2243
rect 51 -2239 52 -2237
rect 51 -2245 52 -2243
rect 58 -2239 59 -2237
rect 58 -2245 59 -2243
rect 65 -2239 66 -2237
rect 65 -2245 66 -2243
rect 72 -2239 73 -2237
rect 75 -2239 76 -2237
rect 72 -2245 73 -2243
rect 75 -2245 76 -2243
rect 79 -2239 80 -2237
rect 79 -2245 80 -2243
rect 86 -2239 87 -2237
rect 86 -2245 87 -2243
rect 93 -2239 94 -2237
rect 93 -2245 94 -2243
rect 100 -2239 101 -2237
rect 100 -2245 101 -2243
rect 107 -2239 108 -2237
rect 107 -2245 108 -2243
rect 117 -2239 118 -2237
rect 114 -2245 115 -2243
rect 117 -2245 118 -2243
rect 121 -2239 122 -2237
rect 121 -2245 122 -2243
rect 128 -2239 129 -2237
rect 128 -2245 129 -2243
rect 135 -2239 136 -2237
rect 138 -2239 139 -2237
rect 135 -2245 136 -2243
rect 138 -2245 139 -2243
rect 142 -2239 143 -2237
rect 142 -2245 143 -2243
rect 149 -2239 150 -2237
rect 152 -2239 153 -2237
rect 149 -2245 150 -2243
rect 156 -2239 157 -2237
rect 156 -2245 157 -2243
rect 163 -2239 164 -2237
rect 163 -2245 164 -2243
rect 170 -2239 171 -2237
rect 170 -2245 171 -2243
rect 177 -2239 178 -2237
rect 177 -2245 178 -2243
rect 184 -2239 185 -2237
rect 184 -2245 185 -2243
rect 191 -2239 192 -2237
rect 191 -2245 192 -2243
rect 198 -2239 199 -2237
rect 198 -2245 199 -2243
rect 205 -2239 206 -2237
rect 205 -2245 206 -2243
rect 212 -2239 213 -2237
rect 212 -2245 213 -2243
rect 219 -2239 220 -2237
rect 219 -2245 220 -2243
rect 226 -2239 227 -2237
rect 226 -2245 227 -2243
rect 233 -2245 234 -2243
rect 240 -2239 241 -2237
rect 240 -2245 241 -2243
rect 247 -2239 248 -2237
rect 247 -2245 248 -2243
rect 254 -2239 255 -2237
rect 254 -2245 255 -2243
rect 261 -2239 262 -2237
rect 261 -2245 262 -2243
rect 268 -2239 269 -2237
rect 268 -2245 269 -2243
rect 275 -2239 276 -2237
rect 275 -2245 276 -2243
rect 282 -2239 283 -2237
rect 282 -2245 283 -2243
rect 289 -2239 290 -2237
rect 289 -2245 290 -2243
rect 296 -2239 297 -2237
rect 299 -2239 300 -2237
rect 296 -2245 297 -2243
rect 299 -2245 300 -2243
rect 303 -2239 304 -2237
rect 303 -2245 304 -2243
rect 310 -2239 311 -2237
rect 310 -2245 311 -2243
rect 317 -2239 318 -2237
rect 317 -2245 318 -2243
rect 324 -2239 325 -2237
rect 324 -2245 325 -2243
rect 331 -2239 332 -2237
rect 331 -2245 332 -2243
rect 338 -2239 339 -2237
rect 338 -2245 339 -2243
rect 341 -2245 342 -2243
rect 345 -2239 346 -2237
rect 345 -2245 346 -2243
rect 352 -2239 353 -2237
rect 352 -2245 353 -2243
rect 359 -2239 360 -2237
rect 359 -2245 360 -2243
rect 366 -2239 367 -2237
rect 366 -2245 367 -2243
rect 373 -2239 374 -2237
rect 373 -2245 374 -2243
rect 380 -2239 381 -2237
rect 380 -2245 381 -2243
rect 387 -2239 388 -2237
rect 387 -2245 388 -2243
rect 394 -2239 395 -2237
rect 397 -2239 398 -2237
rect 394 -2245 395 -2243
rect 397 -2245 398 -2243
rect 401 -2239 402 -2237
rect 404 -2239 405 -2237
rect 401 -2245 402 -2243
rect 404 -2245 405 -2243
rect 408 -2239 409 -2237
rect 411 -2239 412 -2237
rect 408 -2245 409 -2243
rect 411 -2245 412 -2243
rect 415 -2239 416 -2237
rect 415 -2245 416 -2243
rect 425 -2239 426 -2237
rect 422 -2245 423 -2243
rect 425 -2245 426 -2243
rect 429 -2239 430 -2237
rect 429 -2245 430 -2243
rect 436 -2239 437 -2237
rect 436 -2245 437 -2243
rect 443 -2239 444 -2237
rect 443 -2245 444 -2243
rect 450 -2239 451 -2237
rect 453 -2239 454 -2237
rect 450 -2245 451 -2243
rect 453 -2245 454 -2243
rect 457 -2239 458 -2237
rect 457 -2245 458 -2243
rect 464 -2239 465 -2237
rect 464 -2245 465 -2243
rect 471 -2239 472 -2237
rect 471 -2245 472 -2243
rect 478 -2239 479 -2237
rect 478 -2245 479 -2243
rect 485 -2239 486 -2237
rect 485 -2245 486 -2243
rect 492 -2239 493 -2237
rect 492 -2245 493 -2243
rect 499 -2239 500 -2237
rect 499 -2245 500 -2243
rect 506 -2239 507 -2237
rect 506 -2245 507 -2243
rect 513 -2239 514 -2237
rect 513 -2245 514 -2243
rect 520 -2239 521 -2237
rect 523 -2239 524 -2237
rect 520 -2245 521 -2243
rect 523 -2245 524 -2243
rect 527 -2239 528 -2237
rect 530 -2239 531 -2237
rect 527 -2245 528 -2243
rect 530 -2245 531 -2243
rect 534 -2239 535 -2237
rect 534 -2245 535 -2243
rect 541 -2239 542 -2237
rect 541 -2245 542 -2243
rect 548 -2239 549 -2237
rect 548 -2245 549 -2243
rect 555 -2239 556 -2237
rect 555 -2245 556 -2243
rect 558 -2245 559 -2243
rect 562 -2239 563 -2237
rect 562 -2245 563 -2243
rect 569 -2239 570 -2237
rect 569 -2245 570 -2243
rect 576 -2239 577 -2237
rect 576 -2245 577 -2243
rect 583 -2239 584 -2237
rect 583 -2245 584 -2243
rect 590 -2239 591 -2237
rect 590 -2245 591 -2243
rect 597 -2239 598 -2237
rect 597 -2245 598 -2243
rect 604 -2239 605 -2237
rect 604 -2245 605 -2243
rect 611 -2239 612 -2237
rect 611 -2245 612 -2243
rect 618 -2239 619 -2237
rect 621 -2239 622 -2237
rect 618 -2245 619 -2243
rect 621 -2245 622 -2243
rect 625 -2239 626 -2237
rect 628 -2239 629 -2237
rect 628 -2245 629 -2243
rect 632 -2239 633 -2237
rect 632 -2245 633 -2243
rect 639 -2239 640 -2237
rect 639 -2245 640 -2243
rect 646 -2239 647 -2237
rect 649 -2239 650 -2237
rect 646 -2245 647 -2243
rect 653 -2239 654 -2237
rect 653 -2245 654 -2243
rect 660 -2239 661 -2237
rect 660 -2245 661 -2243
rect 667 -2239 668 -2237
rect 667 -2245 668 -2243
rect 677 -2239 678 -2237
rect 677 -2245 678 -2243
rect 681 -2239 682 -2237
rect 681 -2245 682 -2243
rect 688 -2239 689 -2237
rect 688 -2245 689 -2243
rect 695 -2239 696 -2237
rect 695 -2245 696 -2243
rect 702 -2239 703 -2237
rect 702 -2245 703 -2243
rect 709 -2239 710 -2237
rect 709 -2245 710 -2243
rect 716 -2239 717 -2237
rect 716 -2245 717 -2243
rect 723 -2239 724 -2237
rect 723 -2245 724 -2243
rect 730 -2239 731 -2237
rect 730 -2245 731 -2243
rect 737 -2239 738 -2237
rect 737 -2245 738 -2243
rect 744 -2239 745 -2237
rect 744 -2245 745 -2243
rect 751 -2239 752 -2237
rect 751 -2245 752 -2243
rect 758 -2239 759 -2237
rect 758 -2245 759 -2243
rect 765 -2239 766 -2237
rect 768 -2239 769 -2237
rect 765 -2245 766 -2243
rect 772 -2239 773 -2237
rect 772 -2245 773 -2243
rect 779 -2239 780 -2237
rect 779 -2245 780 -2243
rect 786 -2239 787 -2237
rect 786 -2245 787 -2243
rect 793 -2239 794 -2237
rect 793 -2245 794 -2243
rect 800 -2239 801 -2237
rect 800 -2245 801 -2243
rect 807 -2239 808 -2237
rect 810 -2239 811 -2237
rect 807 -2245 808 -2243
rect 810 -2245 811 -2243
rect 814 -2239 815 -2237
rect 814 -2245 815 -2243
rect 821 -2239 822 -2237
rect 821 -2245 822 -2243
rect 828 -2239 829 -2237
rect 828 -2245 829 -2243
rect 835 -2239 836 -2237
rect 835 -2245 836 -2243
rect 842 -2239 843 -2237
rect 842 -2245 843 -2243
rect 849 -2239 850 -2237
rect 849 -2245 850 -2243
rect 856 -2239 857 -2237
rect 856 -2245 857 -2243
rect 863 -2239 864 -2237
rect 863 -2245 864 -2243
rect 870 -2239 871 -2237
rect 870 -2245 871 -2243
rect 873 -2245 874 -2243
rect 877 -2239 878 -2237
rect 877 -2245 878 -2243
rect 884 -2239 885 -2237
rect 884 -2245 885 -2243
rect 891 -2239 892 -2237
rect 891 -2245 892 -2243
rect 898 -2239 899 -2237
rect 898 -2245 899 -2243
rect 905 -2239 906 -2237
rect 905 -2245 906 -2243
rect 912 -2239 913 -2237
rect 912 -2245 913 -2243
rect 919 -2239 920 -2237
rect 919 -2245 920 -2243
rect 926 -2239 927 -2237
rect 926 -2245 927 -2243
rect 933 -2239 934 -2237
rect 936 -2239 937 -2237
rect 933 -2245 934 -2243
rect 940 -2239 941 -2237
rect 940 -2245 941 -2243
rect 947 -2239 948 -2237
rect 947 -2245 948 -2243
rect 954 -2239 955 -2237
rect 954 -2245 955 -2243
rect 961 -2239 962 -2237
rect 961 -2245 962 -2243
rect 968 -2239 969 -2237
rect 968 -2245 969 -2243
rect 975 -2239 976 -2237
rect 975 -2245 976 -2243
rect 982 -2239 983 -2237
rect 985 -2239 986 -2237
rect 982 -2245 983 -2243
rect 985 -2245 986 -2243
rect 989 -2239 990 -2237
rect 989 -2245 990 -2243
rect 996 -2239 997 -2237
rect 996 -2245 997 -2243
rect 1003 -2239 1004 -2237
rect 1003 -2245 1004 -2243
rect 1010 -2239 1011 -2237
rect 1010 -2245 1011 -2243
rect 1017 -2239 1018 -2237
rect 1017 -2245 1018 -2243
rect 1024 -2239 1025 -2237
rect 1024 -2245 1025 -2243
rect 1031 -2239 1032 -2237
rect 1031 -2245 1032 -2243
rect 1038 -2239 1039 -2237
rect 1038 -2245 1039 -2243
rect 1045 -2239 1046 -2237
rect 1045 -2245 1046 -2243
rect 1052 -2239 1053 -2237
rect 1052 -2245 1053 -2243
rect 1059 -2239 1060 -2237
rect 1059 -2245 1060 -2243
rect 1066 -2239 1067 -2237
rect 1066 -2245 1067 -2243
rect 1073 -2239 1074 -2237
rect 1073 -2245 1074 -2243
rect 1080 -2239 1081 -2237
rect 1080 -2245 1081 -2243
rect 1087 -2239 1088 -2237
rect 1087 -2245 1088 -2243
rect 1094 -2239 1095 -2237
rect 1094 -2245 1095 -2243
rect 1101 -2239 1102 -2237
rect 1101 -2245 1102 -2243
rect 1108 -2239 1109 -2237
rect 1108 -2245 1109 -2243
rect 1115 -2239 1116 -2237
rect 1115 -2245 1116 -2243
rect 1122 -2239 1123 -2237
rect 1122 -2245 1123 -2243
rect 1129 -2239 1130 -2237
rect 1129 -2245 1130 -2243
rect 1136 -2239 1137 -2237
rect 1136 -2245 1137 -2243
rect 1143 -2239 1144 -2237
rect 1143 -2245 1144 -2243
rect 1150 -2239 1151 -2237
rect 1150 -2245 1151 -2243
rect 1157 -2239 1158 -2237
rect 1157 -2245 1158 -2243
rect 1164 -2239 1165 -2237
rect 1164 -2245 1165 -2243
rect 1171 -2239 1172 -2237
rect 1171 -2245 1172 -2243
rect 1178 -2239 1179 -2237
rect 1178 -2245 1179 -2243
rect 1185 -2239 1186 -2237
rect 1185 -2245 1186 -2243
rect 1192 -2239 1193 -2237
rect 1192 -2245 1193 -2243
rect 1199 -2239 1200 -2237
rect 1199 -2245 1200 -2243
rect 1206 -2239 1207 -2237
rect 1206 -2245 1207 -2243
rect 1213 -2239 1214 -2237
rect 1213 -2245 1214 -2243
rect 1220 -2239 1221 -2237
rect 1220 -2245 1221 -2243
rect 1227 -2239 1228 -2237
rect 1227 -2245 1228 -2243
rect 1234 -2239 1235 -2237
rect 1234 -2245 1235 -2243
rect 1241 -2239 1242 -2237
rect 1241 -2245 1242 -2243
rect 1248 -2239 1249 -2237
rect 1248 -2245 1249 -2243
rect 1255 -2239 1256 -2237
rect 1255 -2245 1256 -2243
rect 1262 -2239 1263 -2237
rect 1262 -2245 1263 -2243
rect 1269 -2239 1270 -2237
rect 1269 -2245 1270 -2243
rect 1276 -2239 1277 -2237
rect 1276 -2245 1277 -2243
rect 1283 -2239 1284 -2237
rect 1283 -2245 1284 -2243
rect 1290 -2239 1291 -2237
rect 1290 -2245 1291 -2243
rect 1297 -2239 1298 -2237
rect 1297 -2245 1298 -2243
rect 1304 -2239 1305 -2237
rect 1304 -2245 1305 -2243
rect 1311 -2239 1312 -2237
rect 1311 -2245 1312 -2243
rect 2 -2364 3 -2362
rect 5 -2364 6 -2362
rect 9 -2364 10 -2362
rect 9 -2370 10 -2368
rect 16 -2364 17 -2362
rect 16 -2370 17 -2368
rect 23 -2364 24 -2362
rect 23 -2370 24 -2368
rect 30 -2364 31 -2362
rect 30 -2370 31 -2368
rect 37 -2364 38 -2362
rect 40 -2364 41 -2362
rect 37 -2370 38 -2368
rect 40 -2370 41 -2368
rect 44 -2364 45 -2362
rect 44 -2370 45 -2368
rect 51 -2364 52 -2362
rect 51 -2370 52 -2368
rect 54 -2370 55 -2368
rect 58 -2364 59 -2362
rect 61 -2364 62 -2362
rect 58 -2370 59 -2368
rect 61 -2370 62 -2368
rect 65 -2364 66 -2362
rect 65 -2370 66 -2368
rect 72 -2364 73 -2362
rect 72 -2370 73 -2368
rect 79 -2364 80 -2362
rect 79 -2370 80 -2368
rect 86 -2364 87 -2362
rect 86 -2370 87 -2368
rect 93 -2364 94 -2362
rect 96 -2364 97 -2362
rect 93 -2370 94 -2368
rect 100 -2364 101 -2362
rect 100 -2370 101 -2368
rect 107 -2364 108 -2362
rect 107 -2370 108 -2368
rect 114 -2364 115 -2362
rect 114 -2370 115 -2368
rect 121 -2364 122 -2362
rect 121 -2370 122 -2368
rect 128 -2364 129 -2362
rect 128 -2370 129 -2368
rect 135 -2364 136 -2362
rect 138 -2364 139 -2362
rect 135 -2370 136 -2368
rect 138 -2370 139 -2368
rect 142 -2364 143 -2362
rect 142 -2370 143 -2368
rect 149 -2364 150 -2362
rect 152 -2364 153 -2362
rect 156 -2364 157 -2362
rect 156 -2370 157 -2368
rect 163 -2364 164 -2362
rect 163 -2370 164 -2368
rect 170 -2364 171 -2362
rect 170 -2370 171 -2368
rect 177 -2364 178 -2362
rect 177 -2370 178 -2368
rect 184 -2364 185 -2362
rect 184 -2370 185 -2368
rect 191 -2364 192 -2362
rect 191 -2370 192 -2368
rect 198 -2364 199 -2362
rect 198 -2370 199 -2368
rect 205 -2364 206 -2362
rect 205 -2370 206 -2368
rect 212 -2364 213 -2362
rect 212 -2370 213 -2368
rect 219 -2364 220 -2362
rect 219 -2370 220 -2368
rect 226 -2364 227 -2362
rect 226 -2370 227 -2368
rect 233 -2364 234 -2362
rect 233 -2370 234 -2368
rect 240 -2364 241 -2362
rect 240 -2370 241 -2368
rect 247 -2364 248 -2362
rect 247 -2370 248 -2368
rect 254 -2364 255 -2362
rect 254 -2370 255 -2368
rect 261 -2364 262 -2362
rect 261 -2370 262 -2368
rect 268 -2364 269 -2362
rect 268 -2370 269 -2368
rect 275 -2364 276 -2362
rect 275 -2370 276 -2368
rect 282 -2364 283 -2362
rect 282 -2370 283 -2368
rect 289 -2364 290 -2362
rect 289 -2370 290 -2368
rect 296 -2364 297 -2362
rect 296 -2370 297 -2368
rect 306 -2364 307 -2362
rect 303 -2370 304 -2368
rect 306 -2370 307 -2368
rect 310 -2364 311 -2362
rect 310 -2370 311 -2368
rect 317 -2364 318 -2362
rect 320 -2364 321 -2362
rect 317 -2370 318 -2368
rect 320 -2370 321 -2368
rect 324 -2364 325 -2362
rect 324 -2370 325 -2368
rect 331 -2364 332 -2362
rect 331 -2370 332 -2368
rect 338 -2364 339 -2362
rect 341 -2364 342 -2362
rect 341 -2370 342 -2368
rect 345 -2364 346 -2362
rect 345 -2370 346 -2368
rect 352 -2364 353 -2362
rect 352 -2370 353 -2368
rect 359 -2364 360 -2362
rect 359 -2370 360 -2368
rect 366 -2364 367 -2362
rect 366 -2370 367 -2368
rect 373 -2364 374 -2362
rect 373 -2370 374 -2368
rect 380 -2364 381 -2362
rect 380 -2370 381 -2368
rect 387 -2364 388 -2362
rect 387 -2370 388 -2368
rect 394 -2364 395 -2362
rect 397 -2364 398 -2362
rect 394 -2370 395 -2368
rect 397 -2370 398 -2368
rect 401 -2364 402 -2362
rect 401 -2370 402 -2368
rect 408 -2364 409 -2362
rect 408 -2370 409 -2368
rect 415 -2364 416 -2362
rect 415 -2370 416 -2368
rect 425 -2364 426 -2362
rect 422 -2370 423 -2368
rect 425 -2370 426 -2368
rect 429 -2364 430 -2362
rect 429 -2370 430 -2368
rect 436 -2364 437 -2362
rect 436 -2370 437 -2368
rect 439 -2370 440 -2368
rect 443 -2364 444 -2362
rect 443 -2370 444 -2368
rect 450 -2364 451 -2362
rect 450 -2370 451 -2368
rect 457 -2364 458 -2362
rect 457 -2370 458 -2368
rect 464 -2364 465 -2362
rect 464 -2370 465 -2368
rect 471 -2364 472 -2362
rect 471 -2370 472 -2368
rect 478 -2364 479 -2362
rect 478 -2370 479 -2368
rect 485 -2364 486 -2362
rect 485 -2370 486 -2368
rect 492 -2364 493 -2362
rect 492 -2370 493 -2368
rect 499 -2364 500 -2362
rect 499 -2370 500 -2368
rect 506 -2364 507 -2362
rect 506 -2370 507 -2368
rect 513 -2364 514 -2362
rect 516 -2364 517 -2362
rect 513 -2370 514 -2368
rect 516 -2370 517 -2368
rect 520 -2364 521 -2362
rect 520 -2370 521 -2368
rect 527 -2364 528 -2362
rect 527 -2370 528 -2368
rect 534 -2364 535 -2362
rect 534 -2370 535 -2368
rect 541 -2364 542 -2362
rect 541 -2370 542 -2368
rect 548 -2364 549 -2362
rect 548 -2370 549 -2368
rect 555 -2364 556 -2362
rect 558 -2370 559 -2368
rect 562 -2364 563 -2362
rect 562 -2370 563 -2368
rect 569 -2364 570 -2362
rect 569 -2370 570 -2368
rect 576 -2364 577 -2362
rect 579 -2364 580 -2362
rect 576 -2370 577 -2368
rect 579 -2370 580 -2368
rect 583 -2364 584 -2362
rect 583 -2370 584 -2368
rect 590 -2364 591 -2362
rect 593 -2364 594 -2362
rect 590 -2370 591 -2368
rect 593 -2370 594 -2368
rect 597 -2364 598 -2362
rect 597 -2370 598 -2368
rect 604 -2364 605 -2362
rect 604 -2370 605 -2368
rect 611 -2364 612 -2362
rect 611 -2370 612 -2368
rect 618 -2364 619 -2362
rect 618 -2370 619 -2368
rect 625 -2364 626 -2362
rect 625 -2370 626 -2368
rect 632 -2364 633 -2362
rect 635 -2364 636 -2362
rect 632 -2370 633 -2368
rect 635 -2370 636 -2368
rect 639 -2364 640 -2362
rect 639 -2370 640 -2368
rect 646 -2364 647 -2362
rect 646 -2370 647 -2368
rect 653 -2364 654 -2362
rect 653 -2370 654 -2368
rect 660 -2364 661 -2362
rect 663 -2364 664 -2362
rect 660 -2370 661 -2368
rect 667 -2364 668 -2362
rect 667 -2370 668 -2368
rect 674 -2364 675 -2362
rect 674 -2370 675 -2368
rect 681 -2364 682 -2362
rect 681 -2370 682 -2368
rect 688 -2364 689 -2362
rect 688 -2370 689 -2368
rect 695 -2364 696 -2362
rect 695 -2370 696 -2368
rect 702 -2364 703 -2362
rect 702 -2370 703 -2368
rect 709 -2364 710 -2362
rect 709 -2370 710 -2368
rect 716 -2364 717 -2362
rect 716 -2370 717 -2368
rect 726 -2364 727 -2362
rect 723 -2370 724 -2368
rect 726 -2370 727 -2368
rect 730 -2364 731 -2362
rect 730 -2370 731 -2368
rect 737 -2364 738 -2362
rect 737 -2370 738 -2368
rect 744 -2364 745 -2362
rect 747 -2364 748 -2362
rect 744 -2370 745 -2368
rect 751 -2364 752 -2362
rect 751 -2370 752 -2368
rect 758 -2364 759 -2362
rect 761 -2364 762 -2362
rect 758 -2370 759 -2368
rect 761 -2370 762 -2368
rect 765 -2364 766 -2362
rect 765 -2370 766 -2368
rect 772 -2364 773 -2362
rect 772 -2370 773 -2368
rect 779 -2364 780 -2362
rect 779 -2370 780 -2368
rect 786 -2364 787 -2362
rect 786 -2370 787 -2368
rect 793 -2364 794 -2362
rect 793 -2370 794 -2368
rect 800 -2364 801 -2362
rect 800 -2370 801 -2368
rect 807 -2364 808 -2362
rect 810 -2364 811 -2362
rect 807 -2370 808 -2368
rect 810 -2370 811 -2368
rect 814 -2364 815 -2362
rect 814 -2370 815 -2368
rect 821 -2364 822 -2362
rect 821 -2370 822 -2368
rect 828 -2364 829 -2362
rect 828 -2370 829 -2368
rect 835 -2364 836 -2362
rect 835 -2370 836 -2368
rect 842 -2364 843 -2362
rect 842 -2370 843 -2368
rect 849 -2364 850 -2362
rect 849 -2370 850 -2368
rect 852 -2370 853 -2368
rect 856 -2364 857 -2362
rect 856 -2370 857 -2368
rect 863 -2364 864 -2362
rect 863 -2370 864 -2368
rect 870 -2364 871 -2362
rect 870 -2370 871 -2368
rect 877 -2364 878 -2362
rect 877 -2370 878 -2368
rect 884 -2364 885 -2362
rect 884 -2370 885 -2368
rect 891 -2364 892 -2362
rect 891 -2370 892 -2368
rect 898 -2364 899 -2362
rect 898 -2370 899 -2368
rect 905 -2364 906 -2362
rect 905 -2370 906 -2368
rect 912 -2364 913 -2362
rect 912 -2370 913 -2368
rect 919 -2364 920 -2362
rect 919 -2370 920 -2368
rect 926 -2364 927 -2362
rect 926 -2370 927 -2368
rect 933 -2364 934 -2362
rect 933 -2370 934 -2368
rect 940 -2364 941 -2362
rect 940 -2370 941 -2368
rect 947 -2364 948 -2362
rect 947 -2370 948 -2368
rect 954 -2364 955 -2362
rect 954 -2370 955 -2368
rect 961 -2364 962 -2362
rect 961 -2370 962 -2368
rect 968 -2364 969 -2362
rect 968 -2370 969 -2368
rect 975 -2364 976 -2362
rect 975 -2370 976 -2368
rect 982 -2364 983 -2362
rect 982 -2370 983 -2368
rect 989 -2364 990 -2362
rect 989 -2370 990 -2368
rect 996 -2364 997 -2362
rect 996 -2370 997 -2368
rect 1003 -2364 1004 -2362
rect 1003 -2370 1004 -2368
rect 1010 -2364 1011 -2362
rect 1010 -2370 1011 -2368
rect 1017 -2364 1018 -2362
rect 1017 -2370 1018 -2368
rect 1024 -2364 1025 -2362
rect 1024 -2370 1025 -2368
rect 1031 -2364 1032 -2362
rect 1034 -2364 1035 -2362
rect 1034 -2370 1035 -2368
rect 1038 -2364 1039 -2362
rect 1038 -2370 1039 -2368
rect 1045 -2364 1046 -2362
rect 1045 -2370 1046 -2368
rect 1052 -2364 1053 -2362
rect 1052 -2370 1053 -2368
rect 1059 -2364 1060 -2362
rect 1059 -2370 1060 -2368
rect 1066 -2364 1067 -2362
rect 1066 -2370 1067 -2368
rect 1073 -2364 1074 -2362
rect 1073 -2370 1074 -2368
rect 1080 -2364 1081 -2362
rect 1080 -2370 1081 -2368
rect 1087 -2364 1088 -2362
rect 1087 -2370 1088 -2368
rect 1094 -2364 1095 -2362
rect 1094 -2370 1095 -2368
rect 1101 -2364 1102 -2362
rect 1101 -2370 1102 -2368
rect 1108 -2364 1109 -2362
rect 1108 -2370 1109 -2368
rect 1115 -2364 1116 -2362
rect 1115 -2370 1116 -2368
rect 1122 -2364 1123 -2362
rect 1122 -2370 1123 -2368
rect 1129 -2364 1130 -2362
rect 1129 -2370 1130 -2368
rect 1136 -2364 1137 -2362
rect 1136 -2370 1137 -2368
rect 1143 -2364 1144 -2362
rect 1143 -2370 1144 -2368
rect 1150 -2364 1151 -2362
rect 1150 -2370 1151 -2368
rect 1157 -2364 1158 -2362
rect 1157 -2370 1158 -2368
rect 1164 -2364 1165 -2362
rect 1164 -2370 1165 -2368
rect 1171 -2364 1172 -2362
rect 1171 -2370 1172 -2368
rect 1178 -2364 1179 -2362
rect 1178 -2370 1179 -2368
rect 1185 -2364 1186 -2362
rect 1185 -2370 1186 -2368
rect 1192 -2364 1193 -2362
rect 1192 -2370 1193 -2368
rect 1199 -2364 1200 -2362
rect 1199 -2370 1200 -2368
rect 1206 -2364 1207 -2362
rect 1206 -2370 1207 -2368
rect 1213 -2364 1214 -2362
rect 1213 -2370 1214 -2368
rect 1220 -2364 1221 -2362
rect 1220 -2370 1221 -2368
rect 1227 -2364 1228 -2362
rect 1227 -2370 1228 -2368
rect 1234 -2364 1235 -2362
rect 1234 -2370 1235 -2368
rect 1241 -2364 1242 -2362
rect 1241 -2370 1242 -2368
rect 1248 -2364 1249 -2362
rect 1248 -2370 1249 -2368
rect 58 -2461 59 -2459
rect 58 -2467 59 -2465
rect 65 -2461 66 -2459
rect 65 -2467 66 -2465
rect 72 -2461 73 -2459
rect 72 -2467 73 -2465
rect 79 -2461 80 -2459
rect 79 -2467 80 -2465
rect 86 -2461 87 -2459
rect 86 -2467 87 -2465
rect 93 -2461 94 -2459
rect 93 -2467 94 -2465
rect 100 -2461 101 -2459
rect 100 -2467 101 -2465
rect 107 -2461 108 -2459
rect 107 -2467 108 -2465
rect 114 -2461 115 -2459
rect 114 -2467 115 -2465
rect 124 -2461 125 -2459
rect 121 -2467 122 -2465
rect 124 -2467 125 -2465
rect 128 -2461 129 -2459
rect 131 -2461 132 -2459
rect 128 -2467 129 -2465
rect 131 -2467 132 -2465
rect 135 -2461 136 -2459
rect 135 -2467 136 -2465
rect 142 -2461 143 -2459
rect 142 -2467 143 -2465
rect 149 -2461 150 -2459
rect 149 -2467 150 -2465
rect 156 -2461 157 -2459
rect 156 -2467 157 -2465
rect 163 -2461 164 -2459
rect 166 -2467 167 -2465
rect 170 -2461 171 -2459
rect 170 -2467 171 -2465
rect 173 -2467 174 -2465
rect 177 -2461 178 -2459
rect 177 -2467 178 -2465
rect 184 -2461 185 -2459
rect 184 -2467 185 -2465
rect 191 -2461 192 -2459
rect 191 -2467 192 -2465
rect 198 -2461 199 -2459
rect 201 -2461 202 -2459
rect 201 -2467 202 -2465
rect 205 -2461 206 -2459
rect 205 -2467 206 -2465
rect 212 -2461 213 -2459
rect 212 -2467 213 -2465
rect 219 -2461 220 -2459
rect 219 -2467 220 -2465
rect 226 -2461 227 -2459
rect 226 -2467 227 -2465
rect 233 -2461 234 -2459
rect 233 -2467 234 -2465
rect 240 -2461 241 -2459
rect 240 -2467 241 -2465
rect 247 -2461 248 -2459
rect 247 -2467 248 -2465
rect 254 -2461 255 -2459
rect 254 -2467 255 -2465
rect 261 -2461 262 -2459
rect 261 -2467 262 -2465
rect 268 -2461 269 -2459
rect 268 -2467 269 -2465
rect 275 -2461 276 -2459
rect 275 -2467 276 -2465
rect 282 -2461 283 -2459
rect 282 -2467 283 -2465
rect 289 -2461 290 -2459
rect 289 -2467 290 -2465
rect 296 -2461 297 -2459
rect 296 -2467 297 -2465
rect 303 -2461 304 -2459
rect 303 -2467 304 -2465
rect 310 -2461 311 -2459
rect 310 -2467 311 -2465
rect 317 -2461 318 -2459
rect 317 -2467 318 -2465
rect 324 -2461 325 -2459
rect 324 -2467 325 -2465
rect 331 -2461 332 -2459
rect 331 -2467 332 -2465
rect 338 -2461 339 -2459
rect 338 -2467 339 -2465
rect 345 -2461 346 -2459
rect 345 -2467 346 -2465
rect 352 -2461 353 -2459
rect 352 -2467 353 -2465
rect 355 -2467 356 -2465
rect 359 -2461 360 -2459
rect 359 -2467 360 -2465
rect 366 -2461 367 -2459
rect 366 -2467 367 -2465
rect 373 -2461 374 -2459
rect 376 -2461 377 -2459
rect 373 -2467 374 -2465
rect 376 -2467 377 -2465
rect 380 -2461 381 -2459
rect 380 -2467 381 -2465
rect 387 -2461 388 -2459
rect 387 -2467 388 -2465
rect 394 -2461 395 -2459
rect 394 -2467 395 -2465
rect 401 -2461 402 -2459
rect 401 -2467 402 -2465
rect 408 -2461 409 -2459
rect 408 -2467 409 -2465
rect 415 -2461 416 -2459
rect 415 -2467 416 -2465
rect 422 -2461 423 -2459
rect 422 -2467 423 -2465
rect 429 -2461 430 -2459
rect 429 -2467 430 -2465
rect 439 -2461 440 -2459
rect 436 -2467 437 -2465
rect 439 -2467 440 -2465
rect 443 -2461 444 -2459
rect 446 -2461 447 -2459
rect 443 -2467 444 -2465
rect 446 -2467 447 -2465
rect 450 -2461 451 -2459
rect 450 -2467 451 -2465
rect 457 -2461 458 -2459
rect 457 -2467 458 -2465
rect 464 -2461 465 -2459
rect 467 -2461 468 -2459
rect 467 -2467 468 -2465
rect 471 -2461 472 -2459
rect 471 -2467 472 -2465
rect 478 -2461 479 -2459
rect 478 -2467 479 -2465
rect 485 -2461 486 -2459
rect 485 -2467 486 -2465
rect 492 -2461 493 -2459
rect 492 -2467 493 -2465
rect 499 -2461 500 -2459
rect 499 -2467 500 -2465
rect 506 -2461 507 -2459
rect 506 -2467 507 -2465
rect 513 -2461 514 -2459
rect 516 -2461 517 -2459
rect 513 -2467 514 -2465
rect 520 -2461 521 -2459
rect 520 -2467 521 -2465
rect 527 -2461 528 -2459
rect 527 -2467 528 -2465
rect 534 -2461 535 -2459
rect 534 -2467 535 -2465
rect 541 -2461 542 -2459
rect 541 -2467 542 -2465
rect 548 -2461 549 -2459
rect 548 -2467 549 -2465
rect 555 -2461 556 -2459
rect 555 -2467 556 -2465
rect 562 -2461 563 -2459
rect 562 -2467 563 -2465
rect 565 -2467 566 -2465
rect 569 -2461 570 -2459
rect 572 -2461 573 -2459
rect 569 -2467 570 -2465
rect 572 -2467 573 -2465
rect 576 -2461 577 -2459
rect 576 -2467 577 -2465
rect 583 -2461 584 -2459
rect 583 -2467 584 -2465
rect 590 -2461 591 -2459
rect 590 -2467 591 -2465
rect 597 -2461 598 -2459
rect 597 -2467 598 -2465
rect 604 -2461 605 -2459
rect 604 -2467 605 -2465
rect 611 -2461 612 -2459
rect 614 -2461 615 -2459
rect 611 -2467 612 -2465
rect 618 -2461 619 -2459
rect 618 -2467 619 -2465
rect 625 -2461 626 -2459
rect 625 -2467 626 -2465
rect 632 -2461 633 -2459
rect 632 -2467 633 -2465
rect 639 -2461 640 -2459
rect 639 -2467 640 -2465
rect 646 -2461 647 -2459
rect 646 -2467 647 -2465
rect 653 -2461 654 -2459
rect 653 -2467 654 -2465
rect 660 -2461 661 -2459
rect 663 -2461 664 -2459
rect 660 -2467 661 -2465
rect 667 -2461 668 -2459
rect 667 -2467 668 -2465
rect 674 -2461 675 -2459
rect 674 -2467 675 -2465
rect 677 -2467 678 -2465
rect 681 -2461 682 -2459
rect 681 -2467 682 -2465
rect 688 -2461 689 -2459
rect 688 -2467 689 -2465
rect 695 -2461 696 -2459
rect 695 -2467 696 -2465
rect 702 -2461 703 -2459
rect 702 -2467 703 -2465
rect 709 -2461 710 -2459
rect 709 -2467 710 -2465
rect 716 -2461 717 -2459
rect 716 -2467 717 -2465
rect 723 -2461 724 -2459
rect 726 -2461 727 -2459
rect 723 -2467 724 -2465
rect 730 -2461 731 -2459
rect 730 -2467 731 -2465
rect 737 -2461 738 -2459
rect 737 -2467 738 -2465
rect 744 -2461 745 -2459
rect 744 -2467 745 -2465
rect 751 -2461 752 -2459
rect 751 -2467 752 -2465
rect 758 -2461 759 -2459
rect 758 -2467 759 -2465
rect 765 -2461 766 -2459
rect 765 -2467 766 -2465
rect 772 -2461 773 -2459
rect 772 -2467 773 -2465
rect 779 -2461 780 -2459
rect 779 -2467 780 -2465
rect 786 -2461 787 -2459
rect 786 -2467 787 -2465
rect 796 -2461 797 -2459
rect 793 -2467 794 -2465
rect 800 -2461 801 -2459
rect 800 -2467 801 -2465
rect 807 -2461 808 -2459
rect 807 -2467 808 -2465
rect 814 -2461 815 -2459
rect 814 -2467 815 -2465
rect 821 -2461 822 -2459
rect 821 -2467 822 -2465
rect 828 -2461 829 -2459
rect 828 -2467 829 -2465
rect 835 -2461 836 -2459
rect 835 -2467 836 -2465
rect 842 -2461 843 -2459
rect 842 -2467 843 -2465
rect 849 -2461 850 -2459
rect 849 -2467 850 -2465
rect 856 -2461 857 -2459
rect 856 -2467 857 -2465
rect 863 -2461 864 -2459
rect 863 -2467 864 -2465
rect 870 -2461 871 -2459
rect 870 -2467 871 -2465
rect 877 -2461 878 -2459
rect 877 -2467 878 -2465
rect 884 -2461 885 -2459
rect 884 -2467 885 -2465
rect 891 -2461 892 -2459
rect 891 -2467 892 -2465
rect 898 -2461 899 -2459
rect 898 -2467 899 -2465
rect 905 -2461 906 -2459
rect 908 -2461 909 -2459
rect 905 -2467 906 -2465
rect 912 -2461 913 -2459
rect 912 -2467 913 -2465
rect 919 -2461 920 -2459
rect 919 -2467 920 -2465
rect 926 -2461 927 -2459
rect 926 -2467 927 -2465
rect 933 -2461 934 -2459
rect 933 -2467 934 -2465
rect 940 -2461 941 -2459
rect 943 -2461 944 -2459
rect 943 -2467 944 -2465
rect 947 -2461 948 -2459
rect 947 -2467 948 -2465
rect 954 -2461 955 -2459
rect 954 -2467 955 -2465
rect 961 -2461 962 -2459
rect 961 -2467 962 -2465
rect 968 -2461 969 -2459
rect 968 -2467 969 -2465
rect 975 -2461 976 -2459
rect 975 -2467 976 -2465
rect 982 -2461 983 -2459
rect 982 -2467 983 -2465
rect 989 -2461 990 -2459
rect 989 -2467 990 -2465
rect 996 -2461 997 -2459
rect 996 -2467 997 -2465
rect 1003 -2461 1004 -2459
rect 1003 -2467 1004 -2465
rect 1010 -2461 1011 -2459
rect 1013 -2461 1014 -2459
rect 1013 -2467 1014 -2465
rect 1017 -2461 1018 -2459
rect 1017 -2467 1018 -2465
rect 1024 -2461 1025 -2459
rect 1024 -2467 1025 -2465
rect 1031 -2461 1032 -2459
rect 1031 -2467 1032 -2465
rect 1059 -2461 1060 -2459
rect 1059 -2467 1060 -2465
rect 1066 -2461 1067 -2459
rect 1066 -2467 1067 -2465
rect 1073 -2461 1074 -2459
rect 1073 -2467 1074 -2465
rect 1080 -2461 1081 -2459
rect 1080 -2467 1081 -2465
rect 1087 -2461 1088 -2459
rect 1087 -2467 1088 -2465
rect 1094 -2461 1095 -2459
rect 1094 -2467 1095 -2465
rect 1101 -2461 1102 -2459
rect 1104 -2461 1105 -2459
rect 1101 -2467 1102 -2465
rect 1104 -2467 1105 -2465
rect 1108 -2461 1109 -2459
rect 1108 -2467 1109 -2465
rect 1129 -2461 1130 -2459
rect 1129 -2467 1130 -2465
rect 1192 -2461 1193 -2459
rect 1192 -2467 1193 -2465
rect 128 -2544 129 -2542
rect 128 -2550 129 -2548
rect 135 -2544 136 -2542
rect 135 -2550 136 -2548
rect 226 -2544 227 -2542
rect 226 -2550 227 -2548
rect 233 -2544 234 -2542
rect 233 -2550 234 -2548
rect 247 -2544 248 -2542
rect 247 -2550 248 -2548
rect 254 -2544 255 -2542
rect 254 -2550 255 -2548
rect 261 -2544 262 -2542
rect 261 -2550 262 -2548
rect 268 -2544 269 -2542
rect 268 -2550 269 -2548
rect 278 -2544 279 -2542
rect 275 -2550 276 -2548
rect 282 -2544 283 -2542
rect 282 -2550 283 -2548
rect 289 -2544 290 -2542
rect 289 -2550 290 -2548
rect 296 -2544 297 -2542
rect 296 -2550 297 -2548
rect 303 -2544 304 -2542
rect 303 -2550 304 -2548
rect 310 -2544 311 -2542
rect 310 -2550 311 -2548
rect 317 -2544 318 -2542
rect 317 -2550 318 -2548
rect 327 -2544 328 -2542
rect 324 -2550 325 -2548
rect 331 -2544 332 -2542
rect 331 -2550 332 -2548
rect 338 -2544 339 -2542
rect 338 -2550 339 -2548
rect 345 -2544 346 -2542
rect 345 -2550 346 -2548
rect 352 -2544 353 -2542
rect 352 -2550 353 -2548
rect 359 -2544 360 -2542
rect 359 -2550 360 -2548
rect 366 -2544 367 -2542
rect 366 -2550 367 -2548
rect 373 -2544 374 -2542
rect 373 -2550 374 -2548
rect 380 -2544 381 -2542
rect 380 -2550 381 -2548
rect 387 -2544 388 -2542
rect 390 -2544 391 -2542
rect 387 -2550 388 -2548
rect 394 -2544 395 -2542
rect 394 -2550 395 -2548
rect 401 -2544 402 -2542
rect 401 -2550 402 -2548
rect 408 -2544 409 -2542
rect 408 -2550 409 -2548
rect 415 -2544 416 -2542
rect 415 -2550 416 -2548
rect 422 -2544 423 -2542
rect 422 -2550 423 -2548
rect 429 -2544 430 -2542
rect 429 -2550 430 -2548
rect 436 -2544 437 -2542
rect 436 -2550 437 -2548
rect 443 -2544 444 -2542
rect 443 -2550 444 -2548
rect 450 -2544 451 -2542
rect 450 -2550 451 -2548
rect 457 -2544 458 -2542
rect 460 -2544 461 -2542
rect 460 -2550 461 -2548
rect 464 -2544 465 -2542
rect 464 -2550 465 -2548
rect 471 -2544 472 -2542
rect 474 -2544 475 -2542
rect 478 -2544 479 -2542
rect 478 -2550 479 -2548
rect 485 -2544 486 -2542
rect 485 -2550 486 -2548
rect 488 -2550 489 -2548
rect 492 -2544 493 -2542
rect 492 -2550 493 -2548
rect 499 -2544 500 -2542
rect 499 -2550 500 -2548
rect 506 -2544 507 -2542
rect 509 -2544 510 -2542
rect 506 -2550 507 -2548
rect 513 -2544 514 -2542
rect 513 -2550 514 -2548
rect 520 -2544 521 -2542
rect 523 -2544 524 -2542
rect 523 -2550 524 -2548
rect 530 -2544 531 -2542
rect 527 -2550 528 -2548
rect 530 -2550 531 -2548
rect 534 -2544 535 -2542
rect 534 -2550 535 -2548
rect 544 -2544 545 -2542
rect 541 -2550 542 -2548
rect 548 -2544 549 -2542
rect 551 -2544 552 -2542
rect 548 -2550 549 -2548
rect 555 -2544 556 -2542
rect 555 -2550 556 -2548
rect 562 -2544 563 -2542
rect 562 -2550 563 -2548
rect 569 -2544 570 -2542
rect 572 -2544 573 -2542
rect 569 -2550 570 -2548
rect 576 -2544 577 -2542
rect 576 -2550 577 -2548
rect 583 -2544 584 -2542
rect 586 -2544 587 -2542
rect 590 -2544 591 -2542
rect 590 -2550 591 -2548
rect 593 -2550 594 -2548
rect 597 -2544 598 -2542
rect 597 -2550 598 -2548
rect 604 -2544 605 -2542
rect 604 -2550 605 -2548
rect 611 -2544 612 -2542
rect 611 -2550 612 -2548
rect 618 -2544 619 -2542
rect 621 -2550 622 -2548
rect 625 -2544 626 -2542
rect 625 -2550 626 -2548
rect 632 -2544 633 -2542
rect 632 -2550 633 -2548
rect 639 -2544 640 -2542
rect 639 -2550 640 -2548
rect 646 -2544 647 -2542
rect 646 -2550 647 -2548
rect 653 -2544 654 -2542
rect 653 -2550 654 -2548
rect 660 -2544 661 -2542
rect 660 -2550 661 -2548
rect 667 -2544 668 -2542
rect 667 -2550 668 -2548
rect 674 -2544 675 -2542
rect 674 -2550 675 -2548
rect 681 -2544 682 -2542
rect 684 -2544 685 -2542
rect 681 -2550 682 -2548
rect 684 -2550 685 -2548
rect 691 -2544 692 -2542
rect 688 -2550 689 -2548
rect 691 -2550 692 -2548
rect 695 -2544 696 -2542
rect 695 -2550 696 -2548
rect 702 -2544 703 -2542
rect 702 -2550 703 -2548
rect 709 -2544 710 -2542
rect 709 -2550 710 -2548
rect 716 -2544 717 -2542
rect 716 -2550 717 -2548
rect 723 -2544 724 -2542
rect 723 -2550 724 -2548
rect 730 -2544 731 -2542
rect 730 -2550 731 -2548
rect 737 -2544 738 -2542
rect 740 -2544 741 -2542
rect 744 -2544 745 -2542
rect 744 -2550 745 -2548
rect 747 -2550 748 -2548
rect 751 -2544 752 -2542
rect 751 -2550 752 -2548
rect 758 -2544 759 -2542
rect 758 -2550 759 -2548
rect 765 -2544 766 -2542
rect 765 -2550 766 -2548
rect 772 -2544 773 -2542
rect 772 -2550 773 -2548
rect 779 -2544 780 -2542
rect 779 -2550 780 -2548
rect 786 -2544 787 -2542
rect 786 -2550 787 -2548
rect 793 -2544 794 -2542
rect 793 -2550 794 -2548
rect 800 -2544 801 -2542
rect 800 -2550 801 -2548
rect 807 -2544 808 -2542
rect 810 -2544 811 -2542
rect 807 -2550 808 -2548
rect 828 -2544 829 -2542
rect 828 -2550 829 -2548
rect 863 -2544 864 -2542
rect 866 -2544 867 -2542
rect 866 -2550 867 -2548
rect 870 -2544 871 -2542
rect 870 -2550 871 -2548
rect 912 -2544 913 -2542
rect 912 -2550 913 -2548
rect 926 -2544 927 -2542
rect 926 -2550 927 -2548
rect 933 -2544 934 -2542
rect 933 -2550 934 -2548
rect 947 -2544 948 -2542
rect 947 -2550 948 -2548
rect 954 -2544 955 -2542
rect 954 -2550 955 -2548
rect 975 -2544 976 -2542
rect 975 -2550 976 -2548
rect 1017 -2544 1018 -2542
rect 1017 -2550 1018 -2548
rect 1031 -2544 1032 -2542
rect 1031 -2550 1032 -2548
rect 1038 -2544 1039 -2542
rect 1038 -2550 1039 -2548
rect 1052 -2544 1053 -2542
rect 1052 -2550 1053 -2548
rect 1066 -2544 1067 -2542
rect 1066 -2550 1067 -2548
rect 1094 -2544 1095 -2542
rect 1143 -2544 1144 -2542
rect 1143 -2550 1144 -2548
rect 1178 -2544 1179 -2542
rect 1178 -2550 1179 -2548
rect 1181 -2550 1182 -2548
rect 1185 -2544 1186 -2542
rect 1185 -2550 1186 -2548
rect 131 -2589 132 -2587
rect 131 -2595 132 -2593
rect 135 -2589 136 -2587
rect 135 -2595 136 -2593
rect 254 -2589 255 -2587
rect 257 -2589 258 -2587
rect 324 -2589 325 -2587
rect 324 -2595 325 -2593
rect 331 -2589 332 -2587
rect 331 -2595 332 -2593
rect 338 -2589 339 -2587
rect 338 -2595 339 -2593
rect 348 -2595 349 -2593
rect 366 -2589 367 -2587
rect 366 -2595 367 -2593
rect 373 -2589 374 -2587
rect 373 -2595 374 -2593
rect 383 -2589 384 -2587
rect 380 -2595 381 -2593
rect 383 -2595 384 -2593
rect 443 -2589 444 -2587
rect 443 -2595 444 -2593
rect 450 -2589 451 -2587
rect 450 -2595 451 -2593
rect 471 -2589 472 -2587
rect 471 -2595 472 -2593
rect 492 -2589 493 -2587
rect 492 -2595 493 -2593
rect 499 -2589 500 -2587
rect 499 -2595 500 -2593
rect 506 -2589 507 -2587
rect 506 -2595 507 -2593
rect 513 -2589 514 -2587
rect 513 -2595 514 -2593
rect 516 -2595 517 -2593
rect 527 -2589 528 -2587
rect 530 -2589 531 -2587
rect 534 -2589 535 -2587
rect 534 -2595 535 -2593
rect 541 -2589 542 -2587
rect 544 -2589 545 -2587
rect 544 -2595 545 -2593
rect 551 -2589 552 -2587
rect 548 -2595 549 -2593
rect 551 -2595 552 -2593
rect 555 -2589 556 -2587
rect 555 -2595 556 -2593
rect 562 -2589 563 -2587
rect 565 -2589 566 -2587
rect 565 -2595 566 -2593
rect 569 -2589 570 -2587
rect 569 -2595 570 -2593
rect 576 -2589 577 -2587
rect 576 -2595 577 -2593
rect 597 -2589 598 -2587
rect 600 -2589 601 -2587
rect 600 -2595 601 -2593
rect 646 -2589 647 -2587
rect 649 -2589 650 -2587
rect 649 -2595 650 -2593
rect 663 -2589 664 -2587
rect 660 -2595 661 -2593
rect 663 -2595 664 -2593
rect 667 -2589 668 -2587
rect 667 -2595 668 -2593
rect 677 -2589 678 -2587
rect 674 -2595 675 -2593
rect 681 -2589 682 -2587
rect 681 -2595 682 -2593
rect 684 -2595 685 -2593
rect 691 -2589 692 -2587
rect 709 -2589 710 -2587
rect 712 -2589 713 -2587
rect 709 -2595 710 -2593
rect 716 -2589 717 -2587
rect 716 -2595 717 -2593
rect 723 -2589 724 -2587
rect 723 -2595 724 -2593
rect 730 -2589 731 -2587
rect 730 -2595 731 -2593
rect 751 -2589 752 -2587
rect 751 -2595 752 -2593
rect 810 -2589 811 -2587
rect 807 -2595 808 -2593
rect 810 -2595 811 -2593
rect 814 -2589 815 -2587
rect 814 -2595 815 -2593
rect 884 -2589 885 -2587
rect 887 -2589 888 -2587
rect 884 -2595 885 -2593
rect 898 -2589 899 -2587
rect 898 -2595 899 -2593
rect 954 -2589 955 -2587
rect 954 -2595 955 -2593
rect 964 -2589 965 -2587
rect 961 -2595 962 -2593
rect 964 -2595 965 -2593
rect 968 -2589 969 -2587
rect 968 -2595 969 -2593
rect 1013 -2589 1014 -2587
rect 1010 -2595 1011 -2593
rect 1013 -2595 1014 -2593
rect 1017 -2589 1018 -2587
rect 1017 -2595 1018 -2593
rect 1024 -2589 1025 -2587
rect 1024 -2595 1025 -2593
rect 1045 -2589 1046 -2587
rect 1045 -2595 1046 -2593
rect 1052 -2595 1053 -2593
rect 1055 -2595 1056 -2593
rect 1059 -2589 1060 -2587
rect 1059 -2595 1060 -2593
<< metal1 >>
rect 215 0 241 1
rect 247 0 479 1
rect 562 0 640 1
rect 667 0 703 1
rect 800 0 829 1
rect 261 -2 269 -1
rect 275 -2 409 -1
rect 411 -2 507 -1
rect 576 -2 608 -1
rect 681 -2 804 -1
rect 338 -4 381 -3
rect 387 -4 584 -3
rect 586 -4 710 -3
rect 373 -6 402 -5
rect 415 -6 458 -5
rect 464 -6 528 -5
rect 604 -6 766 -5
rect 397 -8 486 -7
rect 425 -10 570 -9
rect 429 -12 517 -11
rect 467 -14 500 -13
rect 163 -25 286 -24
rect 292 -25 339 -24
rect 359 -25 468 -24
rect 478 -25 605 -24
rect 621 -25 724 -24
rect 800 -25 906 -24
rect 191 -27 248 -26
rect 254 -27 402 -26
rect 404 -27 444 -26
rect 464 -27 608 -26
rect 639 -27 689 -26
rect 702 -27 752 -26
rect 828 -27 850 -26
rect 215 -29 220 -28
rect 226 -29 276 -28
rect 282 -29 395 -28
rect 401 -29 412 -28
rect 436 -29 461 -28
rect 481 -29 661 -28
rect 667 -29 675 -28
rect 709 -29 759 -28
rect 765 -29 829 -28
rect 233 -31 241 -30
rect 247 -31 262 -30
rect 268 -31 384 -30
rect 408 -31 472 -30
rect 485 -31 521 -30
rect 527 -31 542 -30
rect 551 -31 598 -30
rect 639 -31 682 -30
rect 719 -31 878 -30
rect 261 -33 388 -32
rect 492 -33 549 -32
rect 555 -33 682 -32
rect 275 -35 356 -34
rect 366 -35 514 -34
rect 516 -35 633 -34
rect 653 -35 717 -34
rect 282 -37 426 -36
rect 499 -37 514 -36
rect 534 -37 703 -36
rect 296 -39 430 -38
rect 502 -39 528 -38
rect 548 -39 619 -38
rect 303 -41 398 -40
rect 429 -41 538 -40
rect 569 -41 626 -40
rect 310 -43 423 -42
rect 457 -43 570 -42
rect 576 -43 612 -42
rect 317 -45 580 -44
rect 583 -45 647 -44
rect 324 -47 374 -46
rect 380 -47 486 -46
rect 506 -47 584 -46
rect 593 -47 773 -46
rect 331 -49 419 -48
rect 457 -49 479 -48
rect 506 -49 563 -48
rect 345 -51 668 -50
rect 373 -53 416 -52
rect 380 -55 563 -54
rect 387 -57 500 -56
rect 23 -68 356 -67
rect 415 -68 549 -67
rect 562 -68 710 -67
rect 723 -68 780 -67
rect 828 -68 871 -67
rect 877 -68 941 -67
rect 1500 -68 1508 -67
rect 30 -70 153 -69
rect 156 -70 293 -69
rect 313 -70 398 -69
rect 422 -70 549 -69
rect 562 -70 640 -69
rect 663 -70 857 -69
rect 905 -70 948 -69
rect 37 -72 332 -71
rect 373 -72 416 -71
rect 478 -72 696 -71
rect 702 -72 801 -71
rect 849 -72 878 -71
rect 44 -74 160 -73
rect 170 -74 311 -73
rect 324 -74 381 -73
rect 394 -74 479 -73
rect 481 -74 486 -73
rect 499 -74 535 -73
rect 541 -74 580 -73
rect 604 -74 724 -73
rect 751 -74 815 -73
rect 51 -76 367 -75
rect 373 -76 430 -75
rect 471 -76 542 -75
rect 576 -76 822 -75
rect 75 -78 101 -77
rect 107 -78 118 -77
rect 121 -78 451 -77
rect 471 -78 556 -77
rect 576 -78 594 -77
rect 604 -78 752 -77
rect 758 -78 787 -77
rect 79 -80 384 -79
rect 429 -80 458 -79
rect 485 -80 612 -79
rect 618 -80 717 -79
rect 772 -80 850 -79
rect 86 -82 90 -81
rect 93 -82 276 -81
rect 296 -82 423 -81
rect 436 -82 458 -81
rect 499 -82 559 -81
rect 618 -82 675 -81
rect 681 -82 731 -81
rect 114 -84 276 -83
rect 299 -84 437 -83
rect 450 -84 598 -83
rect 632 -84 682 -83
rect 688 -84 745 -83
rect 128 -86 213 -85
rect 219 -86 332 -85
rect 352 -86 556 -85
rect 625 -86 633 -85
rect 646 -86 773 -85
rect 135 -88 318 -87
rect 352 -88 360 -87
rect 366 -88 388 -87
rect 404 -88 647 -87
rect 660 -88 675 -87
rect 142 -90 164 -89
rect 177 -90 342 -89
rect 359 -90 703 -89
rect 163 -92 328 -91
rect 338 -92 388 -91
rect 453 -92 689 -91
rect 184 -94 283 -93
rect 338 -94 395 -93
rect 506 -94 612 -93
rect 625 -94 654 -93
rect 660 -94 738 -93
rect 187 -96 227 -95
rect 254 -96 318 -95
rect 464 -96 507 -95
rect 513 -96 598 -95
rect 667 -96 720 -95
rect 149 -98 227 -97
rect 254 -98 262 -97
rect 268 -98 409 -97
rect 411 -98 514 -97
rect 520 -98 640 -97
rect 670 -98 808 -97
rect 149 -100 195 -99
rect 198 -100 234 -99
rect 247 -100 269 -99
rect 271 -100 311 -99
rect 520 -100 608 -99
rect 191 -102 241 -101
rect 247 -102 419 -101
rect 527 -102 766 -101
rect 205 -104 349 -103
rect 530 -104 794 -103
rect 219 -106 346 -105
rect 569 -106 654 -105
rect 233 -108 290 -107
rect 345 -108 591 -107
rect 65 -110 290 -109
rect 443 -110 570 -109
rect 261 -112 402 -111
rect 439 -112 444 -111
rect 492 -112 591 -111
rect 282 -114 538 -113
rect 401 -116 465 -115
rect 492 -116 584 -115
rect 583 -118 762 -117
rect 16 -129 440 -128
rect 488 -129 766 -128
rect 793 -129 829 -128
rect 849 -129 885 -128
rect 940 -129 969 -128
rect 975 -129 1025 -128
rect 9 -131 440 -130
rect 516 -131 598 -130
rect 604 -131 773 -130
rect 800 -131 913 -130
rect 947 -131 979 -130
rect 30 -133 55 -132
rect 58 -133 66 -132
rect 72 -133 76 -132
rect 86 -133 367 -132
rect 394 -133 986 -132
rect 30 -135 62 -134
rect 107 -135 115 -134
rect 117 -135 391 -134
rect 537 -135 836 -134
rect 849 -135 983 -134
rect 44 -137 272 -136
rect 275 -137 360 -136
rect 541 -137 598 -136
rect 607 -137 920 -136
rect 51 -139 402 -138
rect 464 -139 608 -138
rect 611 -139 843 -138
rect 856 -139 962 -138
rect 51 -141 143 -140
rect 145 -141 300 -140
rect 310 -141 402 -140
rect 443 -141 465 -140
rect 478 -141 612 -140
rect 646 -141 794 -140
rect 807 -141 892 -140
rect 58 -143 80 -142
rect 93 -143 276 -142
rect 289 -143 528 -142
rect 555 -143 997 -142
rect 79 -145 164 -144
rect 226 -145 297 -144
rect 327 -145 353 -144
rect 422 -145 479 -144
rect 513 -145 542 -144
rect 562 -145 773 -144
rect 779 -145 857 -144
rect 870 -145 927 -144
rect 121 -147 185 -146
rect 226 -147 363 -146
rect 422 -147 500 -146
rect 520 -147 528 -146
rect 646 -147 682 -146
rect 688 -147 759 -146
rect 779 -147 815 -146
rect 821 -147 955 -146
rect 89 -149 521 -148
rect 639 -149 822 -148
rect 877 -149 948 -148
rect 100 -151 122 -150
rect 131 -151 311 -150
rect 324 -151 353 -150
rect 429 -151 556 -150
rect 583 -151 640 -150
rect 653 -151 878 -150
rect 68 -153 101 -152
rect 135 -153 297 -152
rect 443 -153 710 -152
rect 716 -153 906 -152
rect 135 -155 171 -154
rect 233 -155 367 -154
rect 485 -155 584 -154
rect 590 -155 710 -154
rect 719 -155 801 -154
rect 807 -155 990 -154
rect 142 -157 192 -156
rect 194 -157 234 -156
rect 247 -157 325 -156
rect 415 -157 591 -156
rect 625 -157 654 -156
rect 660 -157 787 -156
rect 149 -159 188 -158
rect 247 -159 398 -158
rect 415 -159 472 -158
rect 485 -159 563 -158
rect 576 -159 626 -158
rect 667 -159 815 -158
rect 44 -161 150 -160
rect 152 -161 192 -160
rect 254 -161 321 -160
rect 387 -161 472 -160
rect 492 -161 577 -160
rect 663 -161 668 -160
rect 674 -161 766 -160
rect 163 -163 178 -162
rect 219 -163 255 -162
rect 271 -163 318 -162
rect 373 -163 388 -162
rect 457 -163 493 -162
rect 569 -163 675 -162
rect 688 -163 696 -162
rect 702 -163 899 -162
rect 170 -165 206 -164
rect 219 -165 307 -164
rect 317 -165 682 -164
rect 723 -165 934 -164
rect 177 -167 213 -166
rect 268 -167 703 -166
rect 730 -167 787 -166
rect 107 -169 269 -168
rect 282 -169 290 -168
rect 303 -169 374 -168
rect 457 -169 696 -168
rect 737 -169 871 -168
rect 198 -171 206 -170
rect 240 -171 283 -170
rect 303 -171 430 -170
rect 530 -171 738 -170
rect 744 -171 864 -170
rect 128 -173 241 -172
rect 331 -173 570 -172
rect 618 -173 724 -172
rect 751 -173 941 -172
rect 93 -175 332 -174
rect 334 -175 731 -174
rect 156 -177 199 -176
rect 436 -177 745 -176
rect 156 -179 213 -178
rect 436 -179 500 -178
rect 534 -179 619 -178
rect 450 -181 535 -180
rect 548 -181 752 -180
rect 408 -183 451 -182
rect 506 -183 549 -182
rect 103 -185 507 -184
rect 380 -187 409 -186
rect 338 -189 381 -188
rect 338 -191 346 -190
rect 37 -193 346 -192
rect 37 -195 262 -194
rect 261 -197 461 -196
rect 2 -208 31 -207
rect 37 -208 388 -207
rect 436 -208 591 -207
rect 604 -208 1081 -207
rect 1150 -208 1179 -207
rect 37 -210 388 -209
rect 394 -210 437 -209
rect 439 -210 843 -209
rect 849 -210 1060 -209
rect 44 -212 286 -211
rect 303 -212 314 -211
rect 446 -212 794 -211
rect 835 -212 1088 -211
rect 44 -214 66 -213
rect 72 -214 83 -213
rect 103 -214 241 -213
rect 243 -214 538 -213
rect 544 -214 822 -213
rect 863 -214 1109 -213
rect 51 -216 990 -215
rect 1024 -216 1046 -215
rect 51 -218 101 -217
rect 107 -218 304 -217
rect 310 -218 395 -217
rect 453 -218 878 -217
rect 891 -218 1018 -217
rect 65 -220 73 -219
rect 107 -220 444 -219
rect 485 -220 815 -219
rect 821 -220 829 -219
rect 870 -220 1102 -219
rect 96 -222 871 -221
rect 912 -222 1123 -221
rect 205 -224 272 -223
rect 282 -224 1067 -223
rect 159 -226 283 -225
rect 310 -226 332 -225
rect 362 -226 836 -225
rect 926 -226 1053 -225
rect 198 -228 206 -227
rect 233 -228 321 -227
rect 415 -228 444 -227
rect 457 -228 913 -227
rect 947 -228 1130 -227
rect 177 -230 199 -229
rect 233 -230 335 -229
rect 408 -230 416 -229
rect 425 -230 829 -229
rect 947 -230 976 -229
rect 54 -232 976 -231
rect 177 -234 318 -233
rect 320 -234 1137 -233
rect 240 -236 318 -235
rect 429 -236 458 -235
rect 506 -236 591 -235
rect 607 -236 1074 -235
rect 124 -238 430 -237
rect 513 -238 1116 -237
rect 268 -240 556 -239
rect 579 -240 1144 -239
rect 128 -242 269 -241
rect 373 -242 507 -241
rect 513 -242 549 -241
rect 607 -242 941 -241
rect 954 -242 1095 -241
rect 26 -244 955 -243
rect 961 -244 1011 -243
rect 128 -246 213 -245
rect 219 -246 374 -245
rect 408 -246 556 -245
rect 639 -246 878 -245
rect 919 -246 962 -245
rect 968 -246 983 -245
rect 170 -248 213 -247
rect 219 -248 227 -247
rect 401 -248 640 -247
rect 674 -248 794 -247
rect 800 -248 969 -247
rect 978 -248 983 -247
rect 40 -250 171 -249
rect 345 -250 402 -249
rect 492 -250 549 -249
rect 576 -250 675 -249
rect 688 -250 717 -249
rect 719 -250 1004 -249
rect 86 -252 493 -251
rect 516 -252 993 -251
rect 58 -254 87 -253
rect 163 -254 227 -253
rect 327 -254 689 -253
rect 695 -254 815 -253
rect 58 -256 290 -255
rect 345 -256 367 -255
rect 534 -256 934 -255
rect 23 -258 290 -257
rect 359 -258 367 -257
rect 534 -258 1154 -257
rect 163 -260 423 -259
rect 576 -260 906 -259
rect 191 -262 360 -261
rect 618 -262 717 -261
rect 737 -262 920 -261
rect 33 -264 192 -263
rect 562 -264 619 -263
rect 625 -264 738 -263
rect 744 -264 941 -263
rect 541 -266 563 -265
rect 583 -266 745 -265
rect 758 -266 1025 -265
rect 380 -268 584 -267
rect 611 -268 626 -267
rect 667 -268 801 -267
rect 884 -268 934 -267
rect 121 -270 381 -269
rect 527 -270 612 -269
rect 698 -270 843 -269
rect 121 -272 486 -271
rect 499 -272 528 -271
rect 541 -272 1032 -271
rect 142 -274 885 -273
rect 114 -276 143 -275
rect 296 -276 500 -275
rect 702 -276 927 -275
rect 114 -278 136 -277
rect 296 -278 605 -277
rect 705 -278 899 -277
rect 135 -280 423 -279
rect 709 -280 850 -279
rect 352 -282 668 -281
rect 730 -282 899 -281
rect 93 -284 353 -283
rect 520 -284 731 -283
rect 758 -284 1039 -283
rect 9 -286 94 -285
rect 478 -286 521 -285
rect 597 -286 710 -285
rect 765 -286 864 -285
rect 9 -288 80 -287
rect 184 -288 598 -287
rect 779 -288 892 -287
rect 184 -290 248 -289
rect 390 -290 766 -289
rect 779 -290 997 -289
rect 247 -292 276 -291
rect 450 -292 479 -291
rect 786 -292 906 -291
rect 254 -294 276 -293
rect 450 -294 752 -293
rect 856 -294 997 -293
rect 254 -296 325 -295
rect 646 -296 787 -295
rect 324 -298 339 -297
rect 569 -298 647 -297
rect 681 -298 857 -297
rect 68 -300 339 -299
rect 653 -300 682 -299
rect 723 -300 752 -299
rect 156 -302 570 -301
rect 653 -302 661 -301
rect 723 -302 808 -301
rect 149 -304 157 -303
rect 660 -304 696 -303
rect 772 -304 808 -303
rect 30 -306 773 -305
rect 54 -308 150 -307
rect 2 -319 41 -318
rect 65 -319 87 -318
rect 93 -319 227 -318
rect 264 -319 276 -318
rect 285 -319 1193 -318
rect 2 -321 45 -320
rect 58 -321 276 -320
rect 310 -321 451 -320
rect 471 -321 545 -320
rect 586 -321 1060 -320
rect 1101 -321 1172 -320
rect 1178 -321 1203 -320
rect 9 -323 31 -322
rect 37 -323 573 -322
rect 604 -323 619 -322
rect 695 -323 1102 -322
rect 1115 -323 1179 -322
rect 9 -325 234 -324
rect 317 -325 500 -324
rect 527 -325 542 -324
rect 702 -325 1165 -324
rect 16 -327 90 -326
rect 93 -327 178 -326
rect 184 -327 503 -326
rect 702 -327 710 -326
rect 758 -327 885 -326
rect 961 -327 1186 -326
rect 16 -329 314 -328
rect 327 -329 598 -328
rect 667 -329 759 -328
rect 884 -329 906 -328
rect 1031 -329 1060 -328
rect 1129 -329 1151 -328
rect 26 -331 192 -330
rect 198 -331 321 -330
rect 359 -331 668 -330
rect 709 -331 724 -330
rect 891 -331 906 -330
rect 996 -331 1032 -330
rect 1052 -331 1116 -330
rect 1136 -331 1158 -330
rect 37 -333 990 -332
rect 1087 -333 1130 -332
rect 44 -335 48 -334
rect 61 -335 234 -334
rect 254 -335 360 -334
rect 394 -335 412 -334
rect 422 -335 479 -334
rect 485 -335 619 -334
rect 653 -335 724 -334
rect 765 -335 997 -334
rect 1024 -335 1088 -334
rect 1094 -335 1137 -334
rect 68 -337 731 -336
rect 786 -337 892 -336
rect 947 -337 1053 -336
rect 72 -339 83 -338
rect 107 -339 111 -338
rect 121 -339 591 -338
rect 625 -339 766 -338
rect 786 -339 815 -338
rect 940 -339 948 -338
rect 982 -339 990 -338
rect 1045 -339 1095 -338
rect 75 -341 1144 -340
rect 79 -343 1025 -342
rect 1122 -343 1144 -342
rect 82 -345 1067 -344
rect 1073 -345 1123 -344
rect 107 -347 136 -346
rect 156 -347 454 -346
rect 471 -347 493 -346
rect 499 -347 563 -346
rect 569 -347 731 -346
rect 814 -347 822 -346
rect 898 -347 941 -346
rect 968 -347 983 -346
rect 1017 -347 1046 -346
rect 110 -349 136 -348
rect 163 -349 479 -348
rect 516 -349 899 -348
rect 954 -349 969 -348
rect 975 -349 1018 -348
rect 1038 -349 1067 -348
rect 96 -351 955 -350
rect 1003 -351 1039 -350
rect 100 -353 164 -352
rect 177 -353 283 -352
rect 303 -353 318 -352
rect 331 -353 423 -352
rect 429 -353 528 -352
rect 555 -353 598 -352
rect 625 -353 633 -352
rect 653 -353 675 -352
rect 800 -353 822 -352
rect 926 -353 976 -352
rect 51 -355 101 -354
rect 114 -355 122 -354
rect 128 -355 185 -354
rect 191 -355 213 -354
rect 219 -355 227 -354
rect 282 -355 374 -354
rect 380 -355 486 -354
rect 509 -355 633 -354
rect 674 -355 780 -354
rect 800 -355 1210 -354
rect 72 -357 115 -356
rect 128 -357 612 -356
rect 779 -357 808 -356
rect 919 -357 927 -356
rect 933 -357 1004 -356
rect 142 -359 220 -358
rect 303 -359 353 -358
rect 366 -359 381 -358
rect 397 -359 1081 -358
rect 86 -361 143 -360
rect 198 -361 206 -360
rect 212 -361 699 -360
rect 772 -361 808 -360
rect 849 -361 934 -360
rect 1010 -361 1081 -360
rect 149 -363 206 -362
rect 289 -363 353 -362
rect 366 -363 643 -362
rect 772 -363 794 -362
rect 828 -363 850 -362
rect 870 -363 920 -362
rect 1010 -363 1109 -362
rect 79 -365 829 -364
rect 149 -367 248 -366
rect 289 -367 552 -366
rect 569 -367 878 -366
rect 247 -369 269 -368
rect 373 -369 521 -368
rect 583 -369 794 -368
rect 835 -369 878 -368
rect 23 -371 836 -370
rect 23 -373 34 -372
rect 261 -373 269 -372
rect 387 -373 1109 -372
rect 261 -375 507 -374
rect 513 -375 556 -374
rect 583 -375 661 -374
rect 751 -375 871 -374
rect 331 -377 661 -376
rect 737 -377 752 -376
rect 345 -379 388 -378
rect 408 -379 962 -378
rect 51 -381 409 -380
rect 415 -381 430 -380
rect 436 -381 696 -380
rect 296 -383 346 -382
rect 415 -383 671 -382
rect 124 -385 297 -384
rect 338 -385 437 -384
rect 450 -385 458 -384
rect 464 -385 493 -384
rect 506 -385 745 -384
rect 124 -387 157 -386
rect 338 -387 577 -386
rect 579 -387 738 -386
rect 324 -389 577 -388
rect 590 -389 1074 -388
rect 240 -391 325 -390
rect 443 -391 458 -390
rect 464 -391 514 -390
rect 520 -391 535 -390
rect 611 -391 647 -390
rect 716 -391 745 -390
rect 58 -393 241 -392
rect 411 -393 717 -392
rect 170 -395 444 -394
rect 534 -395 549 -394
rect 639 -395 647 -394
rect 26 -397 171 -396
rect 254 -397 549 -396
rect 565 -397 640 -396
rect 23 -408 1109 -407
rect 1129 -408 1214 -407
rect 23 -410 265 -409
rect 331 -410 538 -409
rect 548 -410 1172 -409
rect 1209 -410 1396 -409
rect 26 -412 976 -411
rect 1017 -412 1207 -411
rect 30 -414 59 -413
rect 75 -414 122 -413
rect 128 -414 384 -413
rect 408 -414 430 -413
rect 460 -414 920 -413
rect 975 -414 1203 -413
rect 30 -416 941 -415
rect 1038 -416 1130 -415
rect 1136 -416 1221 -415
rect 40 -418 283 -417
rect 331 -418 654 -417
rect 663 -418 1179 -417
rect 44 -420 178 -419
rect 201 -420 206 -419
rect 261 -420 388 -419
rect 401 -420 430 -419
rect 471 -420 514 -419
rect 551 -420 808 -419
rect 814 -420 818 -419
rect 870 -420 941 -419
rect 968 -420 1039 -419
rect 1045 -420 1137 -419
rect 1143 -420 1228 -419
rect 2 -422 45 -421
rect 58 -422 66 -421
rect 79 -422 920 -421
rect 961 -422 1046 -421
rect 1059 -422 1144 -421
rect 1150 -422 1235 -421
rect 9 -424 80 -423
rect 86 -424 178 -423
rect 198 -424 206 -423
rect 261 -424 374 -423
rect 401 -424 612 -423
rect 625 -424 640 -423
rect 670 -424 1053 -423
rect 1066 -424 1151 -423
rect 1157 -424 1256 -423
rect 61 -426 1179 -425
rect 65 -428 556 -427
rect 562 -428 878 -427
rect 898 -428 962 -427
rect 982 -428 1067 -427
rect 1073 -428 1158 -427
rect 47 -430 878 -429
rect 884 -430 899 -429
rect 905 -430 969 -429
rect 1003 -430 1060 -429
rect 1080 -430 1172 -429
rect 86 -432 220 -431
rect 275 -432 388 -431
rect 411 -432 465 -431
rect 478 -432 517 -431
rect 520 -432 556 -431
rect 569 -432 934 -431
rect 1003 -432 1011 -431
rect 89 -434 1242 -433
rect 89 -436 822 -435
rect 828 -436 983 -435
rect 989 -436 1011 -435
rect 93 -438 125 -437
rect 138 -438 1193 -437
rect 72 -440 94 -439
rect 100 -440 409 -439
rect 422 -440 465 -439
rect 478 -440 759 -439
rect 772 -440 822 -439
rect 835 -440 906 -439
rect 1122 -440 1193 -439
rect 33 -442 773 -441
rect 779 -442 836 -441
rect 849 -442 871 -441
rect 1031 -442 1123 -441
rect 100 -444 143 -443
rect 145 -444 829 -443
rect 863 -444 934 -443
rect 107 -446 129 -445
rect 142 -446 185 -445
rect 198 -446 577 -445
rect 590 -446 664 -445
rect 698 -446 1018 -445
rect 107 -448 885 -447
rect 156 -450 549 -449
rect 572 -450 864 -449
rect 163 -452 283 -451
rect 338 -452 563 -451
rect 576 -452 619 -451
rect 632 -452 654 -451
rect 705 -452 1186 -451
rect 170 -454 570 -453
rect 593 -454 696 -453
rect 716 -454 780 -453
rect 793 -454 1032 -453
rect 1101 -454 1186 -453
rect 149 -456 171 -455
rect 184 -456 311 -455
rect 338 -456 493 -455
rect 509 -456 766 -455
rect 800 -456 850 -455
rect 114 -458 766 -457
rect 814 -458 927 -457
rect 114 -460 290 -459
rect 310 -460 318 -459
rect 345 -460 808 -459
rect 856 -460 927 -459
rect 51 -462 290 -461
rect 296 -462 346 -461
rect 373 -462 451 -461
rect 457 -462 472 -461
rect 485 -462 493 -461
rect 520 -462 584 -461
rect 597 -462 633 -461
rect 642 -462 990 -461
rect 51 -464 381 -463
rect 422 -464 794 -463
rect 817 -464 857 -463
rect 149 -466 241 -465
rect 268 -466 276 -465
rect 296 -466 398 -465
rect 425 -466 1074 -465
rect 212 -468 269 -467
rect 366 -468 451 -467
rect 457 -468 591 -467
rect 597 -468 1249 -467
rect 212 -470 234 -469
rect 366 -470 507 -469
rect 534 -470 584 -469
rect 600 -470 997 -469
rect 219 -472 325 -471
rect 380 -472 1081 -471
rect 226 -474 241 -473
rect 303 -474 325 -473
rect 436 -474 486 -473
rect 604 -474 626 -473
rect 646 -474 1102 -473
rect 16 -476 304 -475
rect 317 -476 535 -475
rect 611 -476 1088 -475
rect 16 -478 248 -477
rect 352 -478 437 -477
rect 527 -478 605 -477
rect 614 -478 1053 -477
rect 82 -480 647 -479
rect 681 -480 717 -479
rect 737 -480 759 -479
rect 912 -480 997 -479
rect 1024 -480 1088 -479
rect 159 -482 913 -481
rect 947 -482 1025 -481
rect 191 -484 227 -483
rect 233 -484 395 -483
rect 499 -484 682 -483
rect 751 -484 801 -483
rect 891 -484 948 -483
rect 135 -486 192 -485
rect 254 -486 395 -485
rect 527 -486 1109 -485
rect 135 -488 955 -487
rect 37 -490 955 -489
rect 37 -492 76 -491
rect 163 -492 500 -491
rect 565 -492 738 -491
rect 842 -492 892 -491
rect 352 -494 360 -493
rect 618 -494 675 -493
rect 702 -494 752 -493
rect 786 -494 843 -493
rect 110 -496 360 -495
rect 415 -496 703 -495
rect 730 -496 787 -495
rect 415 -498 1165 -497
rect 502 -500 675 -499
rect 688 -500 731 -499
rect 1094 -500 1165 -499
rect 9 -502 503 -501
rect 688 -502 724 -501
rect 1094 -502 1116 -501
rect 723 -504 745 -503
rect 1115 -504 1200 -503
rect 667 -506 1200 -505
rect 660 -508 668 -507
rect 709 -508 745 -507
rect 443 -510 710 -509
rect 443 -512 531 -511
rect 660 -512 1263 -511
rect 2 -523 1242 -522
rect 1248 -523 1361 -522
rect 1395 -523 1473 -522
rect 1500 -523 1508 -522
rect 2 -525 566 -524
rect 600 -525 1270 -524
rect 16 -527 255 -526
rect 261 -527 458 -526
rect 460 -527 920 -526
rect 1003 -527 1340 -526
rect 30 -529 584 -528
rect 635 -529 759 -528
rect 828 -529 920 -528
rect 940 -529 1004 -528
rect 1094 -529 1284 -528
rect 33 -531 73 -530
rect 75 -531 220 -530
rect 226 -531 381 -530
rect 425 -531 615 -530
rect 660 -531 815 -530
rect 870 -531 941 -530
rect 1024 -531 1095 -530
rect 1150 -531 1242 -530
rect 1255 -531 1375 -530
rect 40 -533 1207 -532
rect 1213 -533 1305 -532
rect 40 -535 1074 -534
rect 1080 -535 1151 -534
rect 1157 -535 1249 -534
rect 1262 -535 1368 -534
rect 47 -537 199 -536
rect 226 -537 276 -536
rect 317 -537 612 -536
rect 614 -537 822 -536
rect 954 -537 1025 -536
rect 1136 -537 1214 -536
rect 1220 -537 1312 -536
rect 72 -539 234 -538
rect 240 -539 262 -538
rect 271 -539 808 -538
rect 912 -539 955 -538
rect 996 -539 1074 -538
rect 1164 -539 1207 -538
rect 1227 -539 1333 -538
rect 110 -541 493 -540
rect 499 -541 1158 -540
rect 1171 -541 1277 -540
rect 114 -543 318 -542
rect 331 -543 510 -542
rect 520 -543 528 -542
rect 530 -543 752 -542
rect 779 -543 829 -542
rect 842 -543 913 -542
rect 933 -543 997 -542
rect 1017 -543 1081 -542
rect 1108 -543 1165 -542
rect 1178 -543 1256 -542
rect 114 -545 1326 -544
rect 117 -547 402 -546
rect 408 -547 500 -546
rect 502 -547 1102 -546
rect 1122 -547 1172 -546
rect 1185 -547 1263 -546
rect 135 -549 1046 -548
rect 1192 -549 1291 -548
rect 121 -551 136 -550
rect 142 -551 878 -550
rect 898 -551 1193 -550
rect 1199 -551 1298 -550
rect 121 -553 248 -552
rect 275 -553 384 -552
rect 401 -553 570 -552
rect 611 -553 1137 -552
rect 1234 -553 1354 -552
rect 44 -555 570 -554
rect 625 -555 752 -554
rect 765 -555 1179 -554
rect 142 -557 202 -556
rect 212 -557 332 -556
rect 338 -557 416 -556
rect 443 -557 493 -556
rect 509 -557 843 -556
rect 849 -557 899 -556
rect 968 -557 1046 -556
rect 1129 -557 1200 -556
rect 58 -559 416 -558
rect 450 -559 454 -558
rect 457 -559 563 -558
rect 625 -559 1319 -558
rect 37 -561 59 -560
rect 138 -561 213 -560
rect 233 -561 311 -560
rect 338 -561 374 -560
rect 450 -561 514 -560
rect 534 -561 1186 -560
rect 79 -563 535 -562
rect 548 -563 584 -562
rect 628 -563 1109 -562
rect 1143 -563 1235 -562
rect 65 -565 549 -564
rect 660 -565 906 -564
rect 1031 -565 1102 -564
rect 65 -567 164 -566
rect 170 -567 255 -566
rect 345 -567 423 -566
rect 464 -567 521 -566
rect 663 -567 780 -566
rect 786 -567 822 -566
rect 835 -567 906 -566
rect 1031 -567 1347 -566
rect 5 -569 423 -568
rect 481 -569 983 -568
rect 1052 -569 1130 -568
rect 23 -571 465 -570
rect 485 -571 514 -570
rect 670 -571 1116 -570
rect 23 -573 325 -572
rect 348 -573 969 -572
rect 1010 -573 1053 -572
rect 1059 -573 1144 -572
rect 79 -575 101 -574
rect 107 -575 983 -574
rect 989 -575 1060 -574
rect 96 -577 101 -576
rect 107 -577 160 -576
rect 163 -577 185 -576
rect 191 -577 199 -576
rect 240 -577 269 -576
rect 324 -577 472 -576
rect 506 -577 850 -576
rect 863 -577 934 -576
rect 947 -577 1011 -576
rect 19 -579 185 -578
rect 191 -579 206 -578
rect 247 -579 258 -578
rect 268 -579 706 -578
rect 723 -579 871 -578
rect 884 -579 948 -578
rect 145 -581 794 -580
rect 800 -581 878 -580
rect 926 -581 990 -580
rect 170 -583 220 -582
rect 250 -583 787 -582
rect 856 -583 927 -582
rect 86 -585 857 -584
rect 86 -587 556 -586
rect 618 -587 1116 -586
rect 205 -589 304 -588
rect 352 -589 447 -588
rect 453 -589 486 -588
rect 506 -589 976 -588
rect 282 -591 619 -590
rect 674 -591 1221 -590
rect 51 -593 283 -592
rect 303 -593 353 -592
rect 359 -593 409 -592
rect 436 -593 675 -592
rect 681 -593 759 -592
rect 765 -593 1039 -592
rect 359 -595 388 -594
rect 418 -595 437 -594
rect 471 -595 563 -594
rect 590 -595 682 -594
rect 688 -595 724 -594
rect 730 -595 801 -594
rect 891 -595 976 -594
rect 89 -597 892 -596
rect 961 -597 1039 -596
rect 289 -599 388 -598
rect 418 -599 1123 -598
rect 289 -601 395 -600
rect 443 -601 591 -600
rect 646 -601 731 -600
rect 737 -601 808 -600
rect 863 -601 962 -600
rect 373 -603 598 -602
rect 653 -603 738 -602
rect 744 -603 815 -602
rect 394 -605 430 -604
rect 478 -605 598 -604
rect 653 -605 710 -604
rect 716 -605 794 -604
rect 44 -607 710 -606
rect 747 -607 885 -606
rect 149 -609 430 -608
rect 541 -609 556 -608
rect 576 -609 647 -608
rect 667 -609 689 -608
rect 695 -609 1067 -608
rect 37 -611 577 -610
rect 632 -611 717 -610
rect 772 -611 836 -610
rect 149 -613 381 -612
rect 390 -613 1067 -612
rect 366 -615 542 -614
rect 632 -615 696 -614
rect 702 -615 1228 -614
rect 156 -617 703 -616
rect 772 -617 1035 -616
rect 128 -619 157 -618
rect 296 -619 367 -618
rect 667 -619 1018 -618
rect 9 -621 297 -620
rect 9 -623 605 -622
rect 93 -625 129 -624
rect 604 -625 699 -624
rect 51 -627 94 -626
rect 37 -638 325 -637
rect 383 -638 731 -637
rect 747 -638 997 -637
rect 1034 -638 1375 -637
rect 1472 -638 1529 -637
rect 2 -640 325 -639
rect 387 -640 451 -639
rect 506 -640 773 -639
rect 807 -640 1438 -639
rect 1507 -640 1515 -639
rect 5 -642 1473 -641
rect 44 -644 1179 -643
rect 1206 -644 1382 -643
rect 44 -646 234 -645
rect 282 -646 346 -645
rect 387 -646 542 -645
rect 544 -646 1452 -645
rect 47 -648 423 -647
rect 443 -648 549 -647
rect 614 -648 752 -647
rect 807 -648 927 -647
rect 940 -648 997 -647
rect 1101 -648 1179 -647
rect 1255 -648 1389 -647
rect 30 -650 423 -649
rect 429 -650 444 -649
rect 446 -650 1459 -649
rect 30 -652 353 -651
rect 408 -652 451 -651
rect 471 -652 773 -651
rect 870 -652 1032 -651
rect 1059 -652 1102 -651
rect 1150 -652 1256 -651
rect 1262 -652 1396 -651
rect 65 -654 94 -653
rect 100 -654 171 -653
rect 233 -654 391 -653
rect 415 -654 661 -653
rect 663 -654 1340 -653
rect 1346 -654 1494 -653
rect 65 -656 220 -655
rect 261 -656 283 -655
rect 296 -656 752 -655
rect 870 -656 1095 -655
rect 1150 -656 1165 -655
rect 1227 -656 1340 -655
rect 1353 -656 1501 -655
rect 23 -658 262 -657
rect 296 -658 395 -657
rect 401 -658 1095 -657
rect 1157 -658 1263 -657
rect 1283 -658 1403 -657
rect 23 -660 311 -659
rect 345 -660 465 -659
rect 506 -660 682 -659
rect 730 -660 738 -659
rect 744 -660 1375 -659
rect 9 -662 682 -661
rect 702 -662 738 -661
rect 744 -662 1046 -661
rect 1052 -662 1284 -661
rect 1290 -662 1410 -661
rect 79 -664 402 -663
rect 415 -664 622 -663
rect 628 -664 1116 -663
rect 1171 -664 1291 -663
rect 1304 -664 1417 -663
rect 79 -666 122 -665
rect 128 -666 171 -665
rect 219 -666 318 -665
rect 348 -666 409 -665
rect 436 -666 472 -665
rect 509 -666 535 -665
rect 548 -666 584 -665
rect 597 -666 927 -665
rect 940 -666 1207 -665
rect 1248 -666 1347 -665
rect 1360 -666 1445 -665
rect 58 -668 584 -667
rect 614 -668 1165 -667
rect 1171 -668 1235 -667
rect 1297 -668 1361 -667
rect 1367 -668 1522 -667
rect 58 -670 157 -669
rect 268 -670 1368 -669
rect 61 -672 1298 -671
rect 1311 -672 1424 -671
rect 86 -674 430 -673
rect 436 -674 605 -673
rect 628 -674 1270 -673
rect 1318 -674 1431 -673
rect 86 -676 332 -675
rect 359 -676 395 -675
rect 604 -676 696 -675
rect 702 -676 794 -675
rect 842 -676 1270 -675
rect 1325 -676 1480 -675
rect 93 -678 601 -677
rect 635 -678 1004 -677
rect 1010 -678 1053 -677
rect 1073 -678 1116 -677
rect 1129 -678 1235 -677
rect 1332 -678 1487 -677
rect 19 -680 1074 -679
rect 1080 -680 1130 -679
rect 1143 -680 1249 -679
rect 72 -682 1144 -681
rect 1199 -682 1312 -681
rect 72 -684 524 -683
rect 747 -684 1186 -683
rect 1199 -684 1242 -683
rect 96 -686 1228 -685
rect 100 -688 619 -687
rect 761 -688 1158 -687
rect 1213 -688 1319 -687
rect 114 -690 374 -689
rect 380 -690 465 -689
rect 478 -690 1081 -689
rect 1108 -690 1214 -689
rect 1220 -690 1326 -689
rect 114 -692 920 -691
rect 943 -692 1277 -691
rect 121 -694 482 -693
rect 618 -694 1305 -693
rect 128 -696 419 -695
rect 425 -696 696 -695
rect 765 -696 1354 -695
rect 135 -698 174 -697
rect 247 -698 332 -697
rect 359 -698 486 -697
rect 513 -698 766 -697
rect 779 -698 794 -697
rect 856 -698 1186 -697
rect 12 -700 857 -699
rect 877 -700 1046 -699
rect 1066 -700 1109 -699
rect 1136 -700 1242 -699
rect 107 -702 248 -701
rect 310 -702 528 -701
rect 537 -702 780 -701
rect 849 -702 878 -701
rect 919 -702 990 -701
rect 1017 -702 1060 -701
rect 1087 -702 1277 -701
rect 107 -704 241 -703
rect 313 -704 479 -703
rect 485 -704 493 -703
rect 499 -704 528 -703
rect 653 -704 1221 -703
rect 149 -706 157 -705
rect 177 -706 241 -705
rect 317 -706 717 -705
rect 835 -706 990 -705
rect 1024 -706 1333 -705
rect 149 -708 626 -707
rect 639 -708 654 -707
rect 667 -708 1018 -707
rect 1038 -708 1088 -707
rect 103 -710 640 -709
rect 667 -710 710 -709
rect 716 -710 801 -709
rect 814 -710 836 -709
rect 849 -710 892 -709
rect 947 -710 1004 -709
rect 177 -712 185 -711
rect 338 -712 514 -711
rect 565 -712 1039 -711
rect 184 -714 213 -713
rect 338 -714 675 -713
rect 709 -714 724 -713
rect 786 -714 801 -713
rect 814 -714 822 -713
rect 954 -714 1011 -713
rect 163 -716 213 -715
rect 355 -716 948 -715
rect 961 -716 1067 -715
rect 142 -718 164 -717
rect 355 -718 458 -717
rect 492 -718 661 -717
rect 786 -718 1123 -717
rect 142 -720 272 -719
rect 366 -720 724 -719
rect 758 -720 1123 -719
rect 75 -722 272 -721
rect 373 -722 521 -721
rect 632 -722 892 -721
rect 898 -722 955 -721
rect 964 -722 1466 -721
rect 289 -724 633 -723
rect 646 -724 675 -723
rect 758 -724 1193 -723
rect 226 -726 290 -725
rect 457 -726 577 -725
rect 590 -726 647 -725
rect 821 -726 888 -725
rect 905 -726 962 -725
rect 968 -726 1025 -725
rect 226 -728 255 -727
rect 499 -728 542 -727
rect 555 -728 591 -727
rect 611 -728 1193 -727
rect 205 -730 255 -729
rect 534 -730 556 -729
rect 569 -730 577 -729
rect 611 -730 1137 -729
rect 205 -732 276 -731
rect 562 -732 570 -731
rect 863 -732 899 -731
rect 905 -732 976 -731
rect 982 -732 1508 -731
rect 117 -734 983 -733
rect 275 -736 304 -735
rect 366 -736 976 -735
rect 198 -738 304 -737
rect 380 -738 563 -737
rect 863 -738 934 -737
rect 51 -740 199 -739
rect 828 -740 934 -739
rect 51 -742 76 -741
rect 117 -742 829 -741
rect 912 -742 969 -741
rect 884 -744 913 -743
rect 842 -746 885 -745
rect 2 -757 1095 -756
rect 2 -759 612 -758
rect 614 -759 1438 -758
rect 9 -761 339 -760
rect 369 -761 944 -760
rect 1066 -761 1095 -760
rect 1437 -761 1459 -760
rect 9 -763 643 -762
rect 649 -763 1298 -762
rect 1458 -763 1473 -762
rect 12 -765 969 -764
rect 1066 -765 1214 -764
rect 1472 -765 1494 -764
rect 23 -767 272 -766
rect 310 -767 713 -766
rect 747 -767 1214 -766
rect 16 -769 24 -768
rect 47 -769 633 -768
rect 653 -769 664 -768
rect 775 -769 1522 -768
rect 16 -771 185 -770
rect 226 -771 367 -770
rect 394 -771 398 -770
rect 485 -771 489 -770
rect 509 -771 1046 -770
rect 1164 -771 1298 -770
rect 58 -773 1508 -772
rect 58 -775 80 -774
rect 117 -775 724 -774
rect 884 -775 1249 -774
rect 51 -777 80 -776
rect 121 -777 311 -776
rect 324 -777 423 -776
rect 485 -777 528 -776
rect 534 -777 1333 -776
rect 51 -779 297 -778
rect 324 -779 440 -778
rect 520 -779 531 -778
rect 537 -779 752 -778
rect 887 -779 1445 -778
rect 61 -781 1074 -780
rect 1164 -781 1326 -780
rect 1332 -781 1347 -780
rect 1444 -781 1487 -780
rect 65 -783 461 -782
rect 520 -783 605 -782
rect 611 -783 899 -782
rect 940 -783 1424 -782
rect 65 -785 318 -784
rect 338 -785 353 -784
rect 394 -785 402 -784
rect 422 -785 577 -784
rect 583 -785 605 -784
rect 618 -785 703 -784
rect 723 -785 801 -784
rect 856 -785 899 -784
rect 943 -785 1256 -784
rect 72 -787 1361 -786
rect 72 -789 262 -788
rect 296 -789 769 -788
rect 800 -789 822 -788
rect 856 -789 948 -788
rect 968 -789 1102 -788
rect 1150 -789 1256 -788
rect 1360 -789 1410 -788
rect 75 -791 1186 -790
rect 1199 -791 1347 -790
rect 1409 -791 1431 -790
rect 100 -793 1424 -792
rect 1430 -793 1452 -792
rect 100 -795 360 -794
rect 401 -795 409 -794
rect 464 -795 577 -794
rect 597 -795 962 -794
rect 1017 -795 1074 -794
rect 1101 -795 1130 -794
rect 1199 -795 1235 -794
rect 1248 -795 1284 -794
rect 1451 -795 1466 -794
rect 114 -797 1326 -796
rect 1465 -797 1480 -796
rect 114 -799 283 -798
rect 408 -799 416 -798
rect 464 -799 1123 -798
rect 1129 -799 1193 -798
rect 1234 -799 1270 -798
rect 1283 -799 1312 -798
rect 1479 -799 1501 -798
rect 121 -801 178 -800
rect 184 -801 304 -800
rect 425 -801 1123 -800
rect 1171 -801 1312 -800
rect 1500 -801 1515 -800
rect 131 -803 171 -802
rect 177 -803 213 -802
rect 226 -803 381 -802
rect 523 -803 990 -802
rect 1017 -803 1263 -802
rect 1269 -803 1305 -802
rect 1514 -803 1529 -802
rect 107 -805 171 -804
rect 205 -805 318 -804
rect 380 -805 556 -804
rect 569 -805 885 -804
rect 891 -805 1151 -804
rect 1192 -805 1228 -804
rect 107 -807 220 -806
rect 236 -807 283 -806
rect 289 -807 304 -806
rect 436 -807 556 -806
rect 618 -807 927 -806
rect 989 -807 1053 -806
rect 1115 -807 1172 -806
rect 1227 -807 1291 -806
rect 30 -809 1053 -808
rect 30 -811 451 -810
rect 467 -811 1291 -810
rect 135 -813 692 -812
rect 695 -813 703 -812
rect 779 -813 1305 -812
rect 135 -815 164 -814
rect 205 -815 1504 -814
rect 138 -817 773 -816
rect 779 -817 794 -816
rect 814 -817 822 -816
rect 905 -817 927 -816
rect 1038 -817 1487 -816
rect 93 -819 815 -818
rect 905 -819 955 -818
rect 1038 -819 1081 -818
rect 93 -821 507 -820
rect 534 -821 598 -820
rect 632 -821 675 -820
rect 681 -821 696 -820
rect 730 -821 773 -820
rect 786 -821 1186 -820
rect 142 -823 360 -822
rect 429 -823 675 -822
rect 688 -823 731 -822
rect 758 -823 955 -822
rect 1045 -823 1088 -822
rect 86 -825 430 -824
rect 436 -825 892 -824
rect 919 -825 962 -824
rect 1080 -825 1137 -824
rect 86 -827 710 -826
rect 758 -827 808 -826
rect 919 -827 997 -826
rect 1087 -827 1207 -826
rect 103 -829 143 -828
rect 163 -829 1494 -828
rect 212 -831 367 -830
rect 450 -831 717 -830
rect 793 -831 836 -830
rect 947 -831 997 -830
rect 1136 -831 1179 -830
rect 1206 -831 1242 -830
rect 219 -833 269 -832
rect 492 -833 682 -832
rect 709 -833 1025 -832
rect 1241 -833 1277 -832
rect 240 -835 290 -834
rect 331 -835 493 -834
rect 506 -835 745 -834
rect 1024 -835 1109 -834
rect 1276 -835 1340 -834
rect 233 -837 241 -836
rect 254 -837 353 -836
rect 541 -837 1032 -836
rect 1108 -837 1144 -836
rect 191 -839 234 -838
rect 261 -839 664 -838
rect 667 -839 752 -838
rect 912 -839 1032 -838
rect 1143 -839 1319 -838
rect 191 -841 276 -840
rect 331 -841 374 -840
rect 541 -841 808 -840
rect 863 -841 913 -840
rect 999 -841 1340 -840
rect 128 -843 276 -842
rect 373 -843 514 -842
rect 544 -843 766 -842
rect 1157 -843 1319 -842
rect 37 -845 514 -844
rect 548 -845 584 -844
rect 600 -845 787 -844
rect 838 -845 1158 -844
rect 128 -847 1354 -846
rect 198 -849 255 -848
rect 268 -849 346 -848
rect 530 -849 549 -848
rect 551 -849 983 -848
rect 1353 -849 1368 -848
rect 198 -851 248 -850
rect 345 -851 356 -850
rect 562 -851 1179 -850
rect 1367 -851 1375 -850
rect 44 -853 248 -852
rect 562 -853 591 -852
rect 639 -853 983 -852
rect 1374 -853 1382 -852
rect 44 -855 717 -854
rect 737 -855 745 -854
rect 765 -855 934 -854
rect 1381 -855 1389 -854
rect 166 -857 591 -856
rect 646 -857 668 -856
rect 737 -857 878 -856
rect 933 -857 1004 -856
rect 1388 -857 1396 -856
rect 457 -859 878 -858
rect 1395 -859 1403 -858
rect 457 -861 1221 -860
rect 1402 -861 1417 -860
rect 569 -863 836 -862
rect 625 -865 1004 -864
rect 40 -867 626 -866
rect 646 -867 1263 -866
rect 653 -869 1116 -868
rect 656 -871 871 -870
rect 660 -873 864 -872
rect 870 -873 976 -872
rect 149 -875 661 -874
rect 761 -875 1221 -874
rect 149 -877 157 -876
rect 828 -877 1417 -876
rect 156 -879 388 -878
rect 639 -879 829 -878
rect 975 -879 1011 -878
rect 369 -881 388 -880
rect 1010 -881 1060 -880
rect 842 -883 1060 -882
rect 842 -885 850 -884
rect 537 -887 850 -886
rect 40 -898 360 -897
rect 376 -898 1179 -897
rect 1318 -898 1427 -897
rect 1503 -898 1515 -897
rect 44 -900 1102 -899
rect 1178 -900 1235 -899
rect 51 -902 465 -901
rect 467 -902 1074 -901
rect 1234 -902 1256 -901
rect 51 -904 297 -903
rect 334 -904 339 -903
rect 352 -904 360 -903
rect 387 -904 552 -903
rect 646 -904 1039 -903
rect 1066 -904 1070 -903
rect 1073 -904 1501 -903
rect 30 -906 388 -905
rect 429 -906 437 -905
rect 443 -906 465 -905
rect 492 -906 650 -905
rect 656 -906 731 -905
rect 747 -906 759 -905
rect 761 -906 1298 -905
rect 30 -908 171 -907
rect 184 -908 244 -907
rect 296 -908 1053 -907
rect 1066 -908 1109 -907
rect 1297 -908 1375 -907
rect 16 -910 171 -909
rect 184 -910 192 -909
rect 198 -910 370 -909
rect 436 -910 528 -909
rect 534 -910 563 -909
rect 660 -910 1046 -909
rect 1094 -910 1256 -909
rect 1374 -910 1438 -909
rect 65 -912 643 -911
rect 691 -912 1011 -911
rect 1017 -912 1319 -911
rect 1437 -912 1494 -911
rect 65 -914 80 -913
rect 100 -914 493 -913
rect 495 -914 647 -913
rect 705 -914 1165 -913
rect 79 -916 94 -915
rect 100 -916 206 -915
rect 212 -916 430 -915
rect 450 -916 601 -915
rect 639 -916 1095 -915
rect 16 -918 94 -917
rect 114 -918 234 -917
rect 240 -918 444 -917
rect 509 -918 675 -917
rect 709 -918 1410 -917
rect 9 -920 675 -919
rect 712 -920 1305 -919
rect 9 -922 73 -921
rect 96 -922 234 -921
rect 338 -922 619 -921
rect 639 -922 993 -921
rect 1045 -922 1123 -921
rect 1143 -922 1410 -921
rect 72 -924 143 -923
rect 145 -924 1053 -923
rect 1122 -924 1137 -923
rect 1143 -924 1200 -923
rect 1290 -924 1305 -923
rect 114 -926 311 -925
rect 352 -926 461 -925
rect 513 -926 528 -925
rect 534 -926 619 -925
rect 667 -926 710 -925
rect 730 -926 801 -925
rect 807 -926 1361 -925
rect 142 -928 1431 -927
rect 163 -930 227 -929
rect 310 -930 416 -929
rect 513 -930 633 -929
rect 754 -930 1228 -929
rect 1290 -930 1354 -929
rect 1360 -930 1424 -929
rect 37 -932 1228 -931
rect 1353 -932 1417 -931
rect 37 -934 157 -933
rect 163 -934 479 -933
rect 520 -934 668 -933
rect 758 -934 1277 -933
rect 1416 -934 1466 -933
rect 2 -936 521 -935
rect 537 -936 1326 -935
rect 2 -938 696 -937
rect 768 -938 1445 -937
rect 131 -940 696 -939
rect 800 -940 892 -939
rect 908 -940 1333 -939
rect 1444 -940 1473 -939
rect 156 -942 654 -941
rect 807 -942 857 -941
rect 891 -942 906 -941
rect 940 -942 955 -941
rect 975 -942 979 -941
rect 989 -942 1039 -941
rect 1129 -942 1137 -941
rect 1199 -942 1249 -941
rect 1325 -942 1382 -941
rect 177 -944 227 -943
rect 380 -944 451 -943
rect 478 -944 878 -943
rect 943 -944 1165 -943
rect 1248 -944 1284 -943
rect 1332 -944 1389 -943
rect 128 -946 178 -945
rect 191 -946 262 -945
rect 275 -946 381 -945
rect 415 -946 1186 -945
rect 1283 -946 1347 -945
rect 1381 -946 1452 -945
rect 121 -948 129 -947
rect 198 -948 237 -947
rect 254 -948 276 -947
rect 373 -948 1452 -947
rect 121 -950 150 -949
rect 205 -950 374 -949
rect 537 -950 1172 -949
rect 1185 -950 1242 -949
rect 1388 -950 1459 -949
rect 149 -952 811 -951
rect 824 -952 927 -951
rect 975 -952 983 -951
rect 1010 -952 1424 -951
rect 212 -954 304 -953
rect 541 -954 1221 -953
rect 1241 -954 1270 -953
rect 254 -956 325 -955
rect 541 -956 563 -955
rect 576 -956 661 -955
rect 677 -956 1221 -955
rect 1269 -956 1312 -955
rect 261 -958 290 -957
rect 303 -958 395 -957
rect 544 -958 591 -957
rect 828 -958 906 -957
rect 926 -958 934 -957
rect 1059 -958 1459 -957
rect 44 -960 545 -959
rect 548 -960 1431 -959
rect 289 -962 409 -961
rect 551 -962 1347 -961
rect 324 -964 346 -963
rect 394 -964 752 -963
rect 828 -964 1277 -963
rect 1311 -964 1340 -963
rect 247 -966 346 -965
rect 401 -966 409 -965
rect 555 -966 577 -965
rect 590 -966 598 -965
rect 831 -966 1032 -965
rect 1059 -966 1081 -965
rect 1129 -966 1193 -965
rect 1339 -966 1396 -965
rect 86 -968 556 -967
rect 597 -968 738 -967
rect 838 -968 1480 -967
rect 86 -970 108 -969
rect 219 -970 402 -969
rect 723 -970 738 -969
rect 849 -970 860 -969
rect 877 -970 885 -969
rect 933 -970 948 -969
rect 996 -970 1396 -969
rect 107 -972 136 -971
rect 219 -972 507 -971
rect 625 -972 850 -971
rect 856 -972 955 -971
rect 968 -972 997 -971
rect 1003 -972 1032 -971
rect 1069 -972 1109 -971
rect 1171 -972 1214 -971
rect 135 -974 458 -973
rect 583 -974 626 -973
rect 884 -974 913 -973
rect 947 -974 962 -973
rect 1003 -974 1116 -973
rect 1192 -974 1368 -973
rect 247 -976 300 -975
rect 331 -976 458 -975
rect 611 -976 969 -975
rect 1080 -976 1151 -975
rect 1213 -976 1263 -975
rect 1367 -976 1487 -975
rect 282 -978 507 -977
rect 611 -978 703 -977
rect 716 -978 1263 -977
rect 282 -980 570 -979
rect 632 -980 703 -979
rect 863 -980 962 -979
rect 1087 -980 1116 -979
rect 1150 -980 1207 -979
rect 366 -982 724 -981
rect 835 -982 1207 -981
rect 268 -984 367 -983
rect 422 -984 584 -983
rect 688 -984 913 -983
rect 1087 -984 1158 -983
rect 268 -986 318 -985
rect 422 -986 745 -985
rect 751 -986 1158 -985
rect 317 -988 689 -987
rect 691 -988 717 -987
rect 744 -988 1102 -987
rect 569 -990 766 -989
rect 786 -990 836 -989
rect 863 -990 871 -989
rect 653 -992 871 -991
rect 765 -994 773 -993
rect 786 -994 815 -993
rect 548 -996 773 -995
rect 793 -996 815 -995
rect 779 -998 794 -997
rect 779 -1000 843 -999
rect 821 -1002 843 -1001
rect 821 -1004 1018 -1003
rect 72 -1015 759 -1014
rect 796 -1015 1039 -1014
rect 1164 -1015 1592 -1014
rect 72 -1017 83 -1016
rect 93 -1017 969 -1016
rect 989 -1017 1235 -1016
rect 1276 -1017 1571 -1016
rect 93 -1019 220 -1018
rect 226 -1019 300 -1018
rect 310 -1019 538 -1018
rect 541 -1019 1312 -1018
rect 1325 -1019 1487 -1018
rect 2 -1021 542 -1020
rect 548 -1021 794 -1020
rect 821 -1021 1410 -1020
rect 1423 -1021 1445 -1020
rect 1451 -1021 1536 -1020
rect 2 -1023 269 -1022
rect 310 -1023 895 -1022
rect 908 -1023 1515 -1022
rect 44 -1025 227 -1024
rect 240 -1025 251 -1024
rect 254 -1025 703 -1024
rect 705 -1025 1452 -1024
rect 23 -1027 45 -1026
rect 96 -1027 584 -1026
rect 590 -1027 689 -1026
rect 691 -1027 969 -1026
rect 992 -1027 1060 -1026
rect 1108 -1027 1235 -1026
rect 1255 -1027 1410 -1026
rect 1437 -1027 1599 -1026
rect 23 -1029 41 -1028
rect 107 -1029 143 -1028
rect 184 -1029 335 -1028
rect 376 -1029 570 -1028
rect 576 -1029 598 -1028
rect 600 -1029 1256 -1028
rect 1283 -1029 1445 -1028
rect 37 -1031 598 -1030
rect 607 -1031 1053 -1030
rect 1143 -1031 1284 -1030
rect 1297 -1031 1480 -1030
rect 37 -1033 59 -1032
rect 107 -1033 178 -1032
rect 184 -1033 353 -1032
rect 390 -1033 1067 -1032
rect 1192 -1033 1473 -1032
rect 33 -1035 178 -1034
rect 201 -1035 220 -1034
rect 240 -1035 755 -1034
rect 842 -1035 906 -1034
rect 940 -1035 1060 -1034
rect 1192 -1035 1214 -1034
rect 1304 -1035 1424 -1034
rect 58 -1037 199 -1036
rect 247 -1037 577 -1036
rect 593 -1037 1319 -1036
rect 1332 -1037 1501 -1036
rect 79 -1039 843 -1038
rect 856 -1039 892 -1038
rect 940 -1039 997 -1038
rect 1052 -1039 1459 -1038
rect 86 -1041 199 -1040
rect 247 -1041 276 -1040
rect 394 -1041 552 -1040
rect 569 -1041 696 -1040
rect 702 -1041 710 -1040
rect 716 -1041 755 -1040
rect 758 -1041 857 -1040
rect 859 -1041 1417 -1040
rect 114 -1043 269 -1042
rect 275 -1043 353 -1042
rect 415 -1043 584 -1042
rect 611 -1043 717 -1042
rect 719 -1043 1326 -1042
rect 1339 -1043 1508 -1042
rect 114 -1045 297 -1044
rect 331 -1045 696 -1044
rect 733 -1045 1039 -1044
rect 1136 -1045 1214 -1044
rect 1290 -1045 1459 -1044
rect 30 -1047 332 -1046
rect 408 -1047 416 -1046
rect 432 -1047 661 -1046
rect 663 -1047 1578 -1046
rect 30 -1049 87 -1048
rect 142 -1049 206 -1048
rect 254 -1049 633 -1048
rect 660 -1049 815 -1048
rect 859 -1049 1438 -1048
rect 156 -1051 297 -1050
rect 338 -1051 633 -1050
rect 667 -1051 822 -1050
rect 863 -1051 990 -1050
rect 996 -1051 1025 -1050
rect 1171 -1051 1319 -1050
rect 1346 -1051 1522 -1050
rect 135 -1053 157 -1052
rect 205 -1053 825 -1052
rect 870 -1053 1403 -1052
rect 121 -1055 136 -1054
rect 261 -1055 374 -1054
rect 408 -1055 682 -1054
rect 730 -1055 815 -1054
rect 936 -1055 1291 -1054
rect 1311 -1055 1431 -1054
rect 121 -1057 192 -1056
rect 212 -1057 262 -1056
rect 338 -1057 482 -1056
rect 485 -1057 549 -1056
rect 562 -1057 710 -1056
rect 747 -1057 808 -1056
rect 954 -1057 1067 -1056
rect 1178 -1057 1333 -1056
rect 1353 -1057 1529 -1056
rect 9 -1059 213 -1058
rect 359 -1059 374 -1058
rect 394 -1059 731 -1058
rect 793 -1059 1403 -1058
rect 145 -1061 192 -1060
rect 359 -1061 381 -1060
rect 446 -1061 1025 -1060
rect 1045 -1061 1172 -1060
rect 1185 -1061 1340 -1060
rect 1367 -1061 1564 -1060
rect 163 -1063 381 -1062
rect 460 -1063 1277 -1062
rect 1374 -1063 1543 -1062
rect 166 -1065 1179 -1064
rect 1199 -1065 1354 -1064
rect 1381 -1065 1550 -1064
rect 464 -1067 871 -1066
rect 933 -1067 1046 -1066
rect 1073 -1067 1186 -1066
rect 1220 -1067 1375 -1066
rect 1388 -1067 1557 -1066
rect 9 -1069 1221 -1068
rect 1227 -1069 1382 -1068
rect 1395 -1069 1585 -1068
rect 243 -1071 465 -1070
rect 478 -1071 521 -1070
rect 534 -1071 1417 -1070
rect 429 -1073 479 -1072
rect 485 -1073 829 -1072
rect 933 -1073 1270 -1072
rect 492 -1075 1347 -1074
rect 355 -1077 493 -1076
rect 495 -1077 864 -1076
rect 947 -1077 1074 -1076
rect 1080 -1077 1368 -1076
rect 499 -1079 535 -1078
rect 544 -1079 682 -1078
rect 828 -1079 1137 -1078
rect 1241 -1079 1389 -1078
rect 471 -1081 500 -1080
rect 555 -1081 808 -1080
rect 877 -1081 948 -1080
rect 954 -1081 1494 -1080
rect 443 -1083 472 -1082
rect 555 -1083 874 -1082
rect 957 -1083 1158 -1082
rect 1248 -1083 1396 -1082
rect 443 -1085 1144 -1084
rect 1248 -1085 1361 -1084
rect 562 -1087 832 -1086
rect 835 -1087 878 -1086
rect 975 -1087 1109 -1086
rect 1115 -1087 1228 -1086
rect 1262 -1087 1431 -1086
rect 79 -1089 1263 -1088
rect 611 -1091 773 -1090
rect 779 -1091 1116 -1090
rect 1129 -1091 1270 -1090
rect 250 -1093 773 -1092
rect 831 -1093 1305 -1092
rect 628 -1095 1298 -1094
rect 653 -1097 1081 -1096
rect 1087 -1097 1242 -1096
rect 604 -1099 654 -1098
rect 670 -1099 1165 -1098
rect 1206 -1099 1361 -1098
rect 674 -1101 1466 -1100
rect 674 -1103 745 -1102
rect 751 -1103 780 -1102
rect 835 -1103 983 -1102
rect 1003 -1103 1158 -1102
rect 513 -1105 745 -1104
rect 751 -1105 1123 -1104
rect 401 -1107 514 -1106
rect 639 -1107 983 -1106
rect 1003 -1107 1018 -1106
rect 1094 -1107 1200 -1106
rect 401 -1109 451 -1108
rect 457 -1109 640 -1108
rect 884 -1109 1130 -1108
rect 450 -1111 647 -1110
rect 737 -1111 885 -1110
rect 912 -1111 1018 -1110
rect 1031 -1111 1095 -1110
rect 1101 -1111 1207 -1110
rect 457 -1113 521 -1112
rect 604 -1113 913 -1112
rect 919 -1113 1123 -1112
rect 625 -1115 647 -1114
rect 723 -1115 1032 -1114
rect 282 -1117 724 -1116
rect 737 -1117 762 -1116
rect 849 -1117 1102 -1116
rect 282 -1119 591 -1118
rect 849 -1119 1011 -1118
rect 317 -1121 626 -1120
rect 898 -1121 920 -1120
rect 926 -1121 1011 -1120
rect 100 -1123 318 -1122
rect 436 -1123 899 -1122
rect 961 -1123 1088 -1122
rect 100 -1125 304 -1124
rect 387 -1125 437 -1124
rect 786 -1125 927 -1124
rect 975 -1125 1427 -1124
rect 65 -1127 304 -1126
rect 667 -1127 787 -1126
rect 800 -1127 962 -1126
rect 51 -1129 66 -1128
rect 765 -1129 801 -1128
rect 16 -1131 766 -1130
rect 16 -1133 290 -1132
rect 51 -1135 507 -1134
rect 233 -1137 290 -1136
rect 506 -1137 678 -1136
rect 149 -1139 234 -1138
rect 128 -1141 150 -1140
rect 128 -1143 619 -1142
rect 527 -1145 619 -1144
rect 366 -1147 528 -1146
rect 324 -1149 367 -1148
rect 324 -1151 388 -1150
rect 9 -1162 304 -1161
rect 341 -1162 346 -1161
rect 352 -1162 668 -1161
rect 670 -1162 801 -1161
rect 828 -1162 1123 -1161
rect 1248 -1162 1252 -1161
rect 9 -1164 608 -1163
rect 667 -1164 773 -1163
rect 782 -1164 808 -1163
rect 828 -1164 864 -1163
rect 894 -1164 1368 -1163
rect 12 -1166 45 -1165
rect 61 -1166 598 -1165
rect 719 -1166 1130 -1165
rect 1248 -1166 1452 -1165
rect 30 -1168 703 -1167
rect 719 -1168 1459 -1167
rect 33 -1170 290 -1169
rect 310 -1170 346 -1169
rect 408 -1170 955 -1169
rect 957 -1170 1529 -1169
rect 37 -1172 724 -1171
rect 730 -1172 1473 -1171
rect 1528 -1172 1564 -1171
rect 37 -1174 759 -1173
rect 772 -1174 934 -1173
rect 954 -1174 983 -1173
rect 989 -1174 993 -1173
rect 1055 -1174 1564 -1173
rect 40 -1176 584 -1175
rect 597 -1176 640 -1175
rect 702 -1176 1270 -1175
rect 1367 -1176 1403 -1175
rect 1451 -1176 1501 -1175
rect 44 -1178 94 -1177
rect 103 -1178 423 -1177
rect 457 -1178 619 -1177
rect 625 -1178 983 -1177
rect 989 -1178 1032 -1177
rect 1122 -1178 1144 -1177
rect 1171 -1178 1473 -1177
rect 51 -1180 458 -1179
rect 481 -1180 1298 -1179
rect 1381 -1180 1459 -1179
rect 51 -1182 178 -1181
rect 184 -1182 734 -1181
rect 754 -1182 1060 -1181
rect 1143 -1182 1165 -1181
rect 1251 -1182 1501 -1181
rect 79 -1184 101 -1183
rect 107 -1184 594 -1183
rect 618 -1184 752 -1183
rect 758 -1184 822 -1183
rect 831 -1184 1109 -1183
rect 1164 -1184 1207 -1183
rect 1297 -1184 1326 -1183
rect 1381 -1184 1438 -1183
rect 79 -1186 388 -1185
rect 408 -1186 486 -1185
rect 506 -1186 860 -1185
rect 863 -1186 878 -1185
rect 922 -1186 1375 -1185
rect 1402 -1186 1424 -1185
rect 82 -1188 465 -1187
rect 485 -1188 563 -1187
rect 569 -1188 822 -1187
rect 835 -1188 937 -1187
rect 996 -1188 1109 -1187
rect 1192 -1188 1326 -1187
rect 1374 -1188 1431 -1187
rect 86 -1190 108 -1189
rect 114 -1190 507 -1189
rect 509 -1190 871 -1189
rect 877 -1190 906 -1189
rect 1059 -1190 1137 -1189
rect 1192 -1190 1389 -1189
rect 1430 -1190 1480 -1189
rect 86 -1192 199 -1191
rect 205 -1192 304 -1191
rect 310 -1192 664 -1191
rect 723 -1192 1018 -1191
rect 1136 -1192 1158 -1191
rect 1206 -1192 1228 -1191
rect 1262 -1192 1424 -1191
rect 1479 -1192 1550 -1191
rect 93 -1194 717 -1193
rect 730 -1194 1081 -1193
rect 1157 -1194 1175 -1193
rect 1227 -1194 1256 -1193
rect 1262 -1194 1487 -1193
rect 100 -1196 997 -1195
rect 1080 -1196 1095 -1195
rect 1255 -1196 1312 -1195
rect 1360 -1196 1487 -1195
rect 114 -1198 479 -1197
rect 513 -1198 605 -1197
rect 611 -1198 871 -1197
rect 905 -1198 920 -1197
rect 940 -1198 1018 -1197
rect 1311 -1198 1333 -1197
rect 1360 -1198 1396 -1197
rect 2 -1200 479 -1199
rect 541 -1200 626 -1199
rect 639 -1200 647 -1199
rect 653 -1200 1550 -1199
rect 2 -1202 976 -1201
rect 1003 -1202 1095 -1201
rect 1220 -1202 1333 -1201
rect 1388 -1202 1543 -1201
rect 121 -1204 531 -1203
rect 541 -1204 556 -1203
rect 583 -1204 766 -1203
rect 786 -1204 808 -1203
rect 856 -1204 1508 -1203
rect 1542 -1204 1599 -1203
rect 121 -1206 269 -1205
rect 289 -1206 339 -1205
rect 366 -1206 388 -1205
rect 394 -1206 717 -1205
rect 751 -1206 1130 -1205
rect 1395 -1206 1445 -1205
rect 1507 -1206 1571 -1205
rect 131 -1208 920 -1207
rect 936 -1208 1221 -1207
rect 1276 -1208 1445 -1207
rect 166 -1210 899 -1209
rect 940 -1210 962 -1209
rect 975 -1210 1074 -1209
rect 1150 -1210 1277 -1209
rect 177 -1212 248 -1211
rect 254 -1212 934 -1211
rect 961 -1212 1046 -1211
rect 1150 -1212 1179 -1211
rect 16 -1214 248 -1213
rect 261 -1214 269 -1213
rect 362 -1214 1046 -1213
rect 1178 -1214 1319 -1213
rect 16 -1216 276 -1215
rect 366 -1216 374 -1215
rect 394 -1216 416 -1215
rect 422 -1216 461 -1215
rect 520 -1216 647 -1215
rect 653 -1216 738 -1215
rect 765 -1216 1116 -1215
rect 1318 -1216 1347 -1215
rect 65 -1218 255 -1217
rect 275 -1218 430 -1217
rect 436 -1218 465 -1217
rect 520 -1218 1536 -1217
rect 65 -1220 528 -1219
rect 548 -1220 563 -1219
rect 590 -1220 1347 -1219
rect 1535 -1220 1585 -1219
rect 170 -1222 262 -1221
rect 317 -1222 437 -1221
rect 527 -1222 1270 -1221
rect 170 -1224 353 -1223
rect 373 -1224 500 -1223
rect 548 -1224 612 -1223
rect 628 -1224 1004 -1223
rect 184 -1226 559 -1225
rect 590 -1226 682 -1225
rect 744 -1226 1116 -1225
rect 191 -1228 206 -1227
rect 212 -1228 447 -1227
rect 555 -1228 1592 -1227
rect 191 -1230 234 -1229
rect 240 -1230 416 -1229
rect 429 -1230 472 -1229
rect 604 -1230 1284 -1229
rect 58 -1232 241 -1231
rect 338 -1232 745 -1231
rect 786 -1232 843 -1231
rect 859 -1232 1354 -1231
rect 149 -1234 234 -1233
rect 380 -1234 500 -1233
rect 681 -1234 689 -1233
rect 796 -1234 1011 -1233
rect 1199 -1234 1284 -1233
rect 1353 -1234 1494 -1233
rect 128 -1236 689 -1235
rect 768 -1236 1200 -1235
rect 1409 -1236 1494 -1235
rect 149 -1238 661 -1237
rect 800 -1238 850 -1237
rect 898 -1238 948 -1237
rect 1010 -1238 1067 -1237
rect 1409 -1238 1417 -1237
rect 198 -1240 318 -1239
rect 401 -1240 570 -1239
rect 660 -1240 727 -1239
rect 814 -1240 857 -1239
rect 947 -1240 969 -1239
rect 1066 -1240 1088 -1239
rect 1416 -1240 1466 -1239
rect 212 -1242 360 -1241
rect 401 -1242 577 -1241
rect 632 -1242 815 -1241
rect 838 -1242 1074 -1241
rect 1087 -1242 1102 -1241
rect 1465 -1242 1515 -1241
rect 219 -1244 514 -1243
rect 576 -1244 927 -1243
rect 968 -1244 1025 -1243
rect 1514 -1244 1578 -1243
rect 142 -1246 220 -1245
rect 226 -1246 391 -1245
rect 450 -1246 843 -1245
rect 849 -1246 885 -1245
rect 912 -1246 1102 -1245
rect 58 -1248 885 -1247
rect 926 -1248 1053 -1247
rect 128 -1250 143 -1249
rect 226 -1250 325 -1249
rect 450 -1250 535 -1249
rect 632 -1250 696 -1249
rect 737 -1250 1053 -1249
rect 296 -1252 381 -1251
rect 471 -1252 710 -1251
rect 779 -1252 913 -1251
rect 1024 -1252 1039 -1251
rect 163 -1254 710 -1253
rect 779 -1254 1438 -1253
rect 156 -1256 164 -1255
rect 296 -1256 493 -1255
rect 534 -1256 794 -1255
rect 1038 -1256 1186 -1255
rect 135 -1258 157 -1257
rect 173 -1258 794 -1257
rect 1185 -1258 1214 -1257
rect 135 -1260 360 -1259
rect 492 -1260 836 -1259
rect 1213 -1260 1235 -1259
rect 320 -1262 696 -1261
rect 1234 -1262 1242 -1261
rect 324 -1264 332 -1263
rect 1241 -1264 1291 -1263
rect 331 -1266 444 -1265
rect 1290 -1266 1305 -1265
rect 443 -1268 755 -1267
rect 1304 -1268 1340 -1267
rect 1339 -1270 1522 -1269
rect 1521 -1272 1557 -1271
rect 891 -1274 1557 -1273
rect 355 -1276 892 -1275
rect 2 -1287 556 -1286
rect 562 -1287 605 -1286
rect 649 -1287 1487 -1286
rect 2 -1289 374 -1288
rect 478 -1289 1291 -1288
rect 1451 -1289 1455 -1288
rect 1486 -1289 1515 -1288
rect 30 -1291 755 -1290
rect 765 -1291 1347 -1290
rect 1451 -1291 1466 -1290
rect 1514 -1291 1543 -1290
rect 30 -1293 45 -1292
rect 61 -1293 1473 -1292
rect 37 -1295 521 -1294
rect 527 -1295 542 -1294
rect 548 -1295 1550 -1294
rect 37 -1297 444 -1296
rect 488 -1297 500 -1296
rect 509 -1297 983 -1296
rect 1052 -1297 1459 -1296
rect 1472 -1297 1480 -1296
rect 44 -1299 241 -1298
rect 338 -1299 409 -1298
rect 422 -1299 444 -1298
rect 467 -1299 500 -1298
rect 548 -1299 780 -1298
rect 782 -1299 1522 -1298
rect 68 -1301 815 -1300
rect 835 -1301 1235 -1300
rect 1346 -1301 1368 -1300
rect 1388 -1301 1459 -1300
rect 1479 -1301 1508 -1300
rect 100 -1303 430 -1302
rect 555 -1303 675 -1302
rect 719 -1303 1522 -1302
rect 100 -1305 150 -1304
rect 177 -1305 321 -1304
rect 345 -1305 374 -1304
rect 387 -1305 430 -1304
rect 562 -1305 787 -1304
rect 793 -1305 1007 -1304
rect 1055 -1305 1529 -1304
rect 79 -1307 388 -1306
rect 401 -1307 542 -1306
rect 674 -1307 682 -1306
rect 723 -1307 1032 -1306
rect 1171 -1307 1403 -1306
rect 1454 -1307 1466 -1306
rect 1507 -1307 1536 -1306
rect 79 -1309 199 -1308
rect 233 -1309 360 -1308
rect 418 -1309 1368 -1308
rect 1388 -1309 1431 -1308
rect 1528 -1309 1557 -1308
rect 82 -1311 178 -1310
rect 198 -1311 531 -1310
rect 632 -1311 682 -1310
rect 723 -1311 769 -1310
rect 779 -1311 829 -1310
rect 835 -1311 843 -1310
rect 880 -1311 1501 -1310
rect 86 -1313 321 -1312
rect 345 -1313 363 -1312
rect 422 -1313 451 -1312
rect 481 -1313 794 -1312
rect 828 -1313 857 -1312
rect 922 -1313 1445 -1312
rect 86 -1315 416 -1314
rect 450 -1315 486 -1314
rect 604 -1315 923 -1314
rect 933 -1315 1494 -1314
rect 9 -1317 486 -1316
rect 737 -1317 874 -1316
rect 933 -1317 955 -1316
rect 975 -1317 1053 -1316
rect 1101 -1317 1536 -1316
rect 9 -1319 66 -1318
rect 93 -1319 150 -1318
rect 212 -1319 482 -1318
rect 667 -1319 738 -1318
rect 744 -1319 815 -1318
rect 838 -1319 864 -1318
rect 898 -1319 955 -1318
rect 982 -1319 997 -1318
rect 1024 -1319 1032 -1318
rect 1101 -1319 1214 -1318
rect 1234 -1319 1263 -1318
rect 1339 -1319 1494 -1318
rect 93 -1321 570 -1320
rect 618 -1321 668 -1320
rect 688 -1321 745 -1320
rect 751 -1321 1312 -1320
rect 1353 -1321 1431 -1320
rect 103 -1323 1424 -1322
rect 110 -1325 297 -1324
rect 303 -1325 752 -1324
rect 765 -1325 801 -1324
rect 849 -1325 899 -1324
rect 961 -1325 1025 -1324
rect 1038 -1325 1214 -1324
rect 1255 -1325 1501 -1324
rect 128 -1327 860 -1326
rect 863 -1327 927 -1326
rect 940 -1327 962 -1326
rect 996 -1327 1004 -1326
rect 1010 -1327 1039 -1326
rect 1087 -1327 1340 -1326
rect 1395 -1327 1403 -1326
rect 1416 -1327 1424 -1326
rect 107 -1329 129 -1328
rect 131 -1329 703 -1328
rect 712 -1329 1263 -1328
rect 1311 -1329 1361 -1328
rect 1395 -1329 1438 -1328
rect 107 -1331 115 -1330
rect 215 -1331 297 -1330
rect 303 -1331 325 -1330
rect 352 -1331 528 -1330
rect 618 -1331 640 -1330
rect 730 -1331 1088 -1330
rect 1143 -1331 1172 -1330
rect 1178 -1331 1291 -1330
rect 1332 -1331 1438 -1330
rect 16 -1333 353 -1332
rect 436 -1333 570 -1332
rect 639 -1333 913 -1332
rect 926 -1333 990 -1332
rect 1059 -1333 1144 -1332
rect 1157 -1333 1445 -1332
rect 16 -1335 206 -1334
rect 233 -1335 311 -1334
rect 436 -1335 465 -1334
rect 471 -1335 689 -1334
rect 786 -1335 871 -1334
rect 940 -1335 979 -1334
rect 989 -1335 1151 -1334
rect 1164 -1335 1179 -1334
rect 1192 -1335 1354 -1334
rect 1360 -1335 1375 -1334
rect 51 -1337 115 -1336
rect 170 -1337 325 -1336
rect 457 -1337 703 -1336
rect 800 -1337 808 -1336
rect 842 -1337 850 -1336
rect 856 -1337 878 -1336
rect 947 -1337 1011 -1336
rect 1122 -1337 1158 -1336
rect 1255 -1337 1277 -1336
rect 1374 -1337 1382 -1336
rect 51 -1339 262 -1338
rect 275 -1339 311 -1338
rect 317 -1339 808 -1338
rect 877 -1339 892 -1338
rect 905 -1339 948 -1338
rect 1003 -1339 1060 -1338
rect 1122 -1339 1228 -1338
rect 1248 -1339 1382 -1338
rect 65 -1341 913 -1340
rect 1080 -1341 1249 -1340
rect 1269 -1341 1277 -1340
rect 142 -1343 171 -1342
rect 184 -1343 276 -1342
rect 317 -1343 633 -1342
rect 695 -1343 1270 -1342
rect 58 -1345 696 -1344
rect 884 -1345 906 -1344
rect 1073 -1345 1081 -1344
rect 1129 -1345 1333 -1344
rect 58 -1347 626 -1346
rect 884 -1347 969 -1346
rect 1066 -1347 1074 -1346
rect 1136 -1347 1165 -1346
rect 1227 -1347 1319 -1346
rect 135 -1349 1130 -1348
rect 1136 -1349 1200 -1348
rect 1297 -1349 1319 -1348
rect 72 -1351 136 -1350
rect 142 -1351 290 -1350
rect 457 -1351 493 -1350
rect 495 -1351 871 -1350
rect 891 -1351 920 -1350
rect 1045 -1351 1067 -1350
rect 1150 -1351 1186 -1350
rect 1199 -1351 1207 -1350
rect 1297 -1351 1326 -1350
rect 72 -1353 220 -1352
rect 226 -1353 472 -1352
rect 478 -1353 731 -1352
rect 1108 -1353 1207 -1352
rect 1304 -1353 1326 -1352
rect 121 -1355 290 -1354
rect 464 -1355 598 -1354
rect 625 -1355 661 -1354
rect 709 -1355 1109 -1354
rect 1185 -1355 1564 -1354
rect 121 -1357 332 -1356
rect 492 -1357 521 -1356
rect 523 -1357 1046 -1356
rect 163 -1359 185 -1358
rect 205 -1359 559 -1358
rect 597 -1359 951 -1358
rect 1017 -1359 1305 -1358
rect 163 -1361 405 -1360
rect 506 -1361 1417 -1360
rect 219 -1363 535 -1362
rect 611 -1363 661 -1362
rect 709 -1363 1116 -1362
rect 226 -1365 717 -1364
rect 845 -1365 1116 -1364
rect 240 -1367 381 -1366
rect 390 -1367 535 -1366
rect 551 -1367 717 -1366
rect 247 -1369 409 -1368
rect 506 -1369 976 -1368
rect 247 -1371 584 -1370
rect 590 -1371 612 -1370
rect 254 -1373 360 -1372
rect 380 -1373 395 -1372
rect 513 -1373 584 -1372
rect 590 -1373 727 -1372
rect 212 -1375 255 -1374
rect 261 -1375 608 -1374
rect 331 -1377 1018 -1376
rect 394 -1379 654 -1378
rect 513 -1381 1284 -1380
rect 516 -1383 1284 -1382
rect 523 -1385 1193 -1384
rect 576 -1387 654 -1386
rect 576 -1389 822 -1388
rect 758 -1391 822 -1390
rect 646 -1393 759 -1392
rect 646 -1395 969 -1394
rect 44 -1406 650 -1405
rect 684 -1406 731 -1405
rect 800 -1406 839 -1405
rect 842 -1406 1354 -1405
rect 44 -1408 115 -1407
rect 121 -1408 468 -1407
rect 471 -1408 496 -1407
rect 520 -1408 528 -1407
rect 646 -1408 1270 -1407
rect 1353 -1408 1361 -1407
rect 51 -1410 419 -1409
rect 478 -1410 1193 -1409
rect 1311 -1410 1361 -1409
rect 51 -1412 318 -1411
rect 320 -1412 409 -1411
rect 478 -1412 1144 -1411
rect 1192 -1412 1298 -1411
rect 65 -1414 297 -1413
rect 366 -1414 398 -1413
rect 408 -1414 493 -1413
rect 499 -1414 521 -1413
rect 646 -1414 1116 -1413
rect 1276 -1414 1312 -1413
rect 65 -1416 570 -1415
rect 712 -1416 780 -1415
rect 800 -1416 1305 -1415
rect 82 -1418 276 -1417
rect 296 -1418 339 -1417
rect 390 -1418 524 -1417
rect 562 -1418 780 -1417
rect 807 -1418 1270 -1417
rect 68 -1420 339 -1419
rect 394 -1420 832 -1419
rect 842 -1420 857 -1419
rect 873 -1420 1235 -1419
rect 1262 -1420 1277 -1419
rect 82 -1422 122 -1421
rect 184 -1422 514 -1421
rect 562 -1422 661 -1421
rect 723 -1422 727 -1421
rect 730 -1422 836 -1421
rect 856 -1422 1207 -1421
rect 1234 -1422 1522 -1421
rect 93 -1424 493 -1423
rect 513 -1424 542 -1423
rect 569 -1424 993 -1423
rect 1003 -1424 1046 -1423
rect 1076 -1424 1319 -1423
rect 1332 -1424 1522 -1423
rect 37 -1426 94 -1425
rect 100 -1426 405 -1425
rect 464 -1426 1144 -1425
rect 1164 -1426 1263 -1425
rect 37 -1428 836 -1427
rect 880 -1428 934 -1427
rect 950 -1428 1466 -1427
rect 100 -1430 255 -1429
rect 275 -1430 689 -1429
rect 723 -1430 1214 -1429
rect 1444 -1430 1466 -1429
rect 103 -1432 433 -1431
rect 436 -1432 465 -1431
rect 481 -1432 1298 -1431
rect 1416 -1432 1445 -1431
rect 114 -1434 262 -1433
rect 324 -1434 367 -1433
rect 436 -1434 633 -1433
rect 660 -1434 745 -1433
rect 768 -1434 808 -1433
rect 880 -1434 1326 -1433
rect 1381 -1434 1417 -1433
rect 135 -1436 255 -1435
rect 261 -1436 360 -1435
rect 541 -1436 850 -1435
rect 884 -1436 888 -1435
rect 919 -1436 1508 -1435
rect 79 -1438 1508 -1437
rect 135 -1440 174 -1439
rect 184 -1440 192 -1439
rect 205 -1440 528 -1439
rect 555 -1440 1165 -1439
rect 1178 -1440 1333 -1439
rect 1381 -1440 1410 -1439
rect 72 -1442 206 -1441
rect 219 -1442 601 -1441
rect 688 -1442 696 -1441
rect 744 -1442 773 -1441
rect 803 -1442 1046 -1441
rect 1080 -1442 1207 -1441
rect 1213 -1442 1221 -1441
rect 1409 -1442 1459 -1441
rect 72 -1444 654 -1443
rect 772 -1444 899 -1443
rect 905 -1444 1081 -1443
rect 1129 -1444 1326 -1443
rect 191 -1446 584 -1445
rect 653 -1446 675 -1445
rect 849 -1446 1039 -1445
rect 1129 -1446 1256 -1445
rect 219 -1448 517 -1447
rect 583 -1448 619 -1447
rect 859 -1448 1459 -1447
rect 233 -1450 318 -1449
rect 324 -1450 549 -1449
rect 884 -1450 962 -1449
rect 975 -1450 1515 -1449
rect 177 -1452 234 -1451
rect 240 -1452 678 -1451
rect 887 -1452 962 -1451
rect 978 -1452 1249 -1451
rect 1514 -1452 1525 -1451
rect 177 -1454 591 -1453
rect 674 -1454 1249 -1453
rect 1437 -1454 1525 -1453
rect 198 -1456 549 -1455
rect 898 -1456 955 -1455
rect 1006 -1456 1424 -1455
rect 16 -1458 199 -1457
rect 226 -1458 591 -1457
rect 905 -1458 941 -1457
rect 947 -1458 1256 -1457
rect 1388 -1458 1424 -1457
rect 16 -1460 31 -1459
rect 226 -1460 346 -1459
rect 359 -1460 444 -1459
rect 485 -1460 556 -1459
rect 919 -1460 969 -1459
rect 1017 -1460 1088 -1459
rect 1136 -1460 1305 -1459
rect 1374 -1460 1389 -1459
rect 30 -1462 507 -1461
rect 877 -1462 969 -1461
rect 989 -1462 1137 -1461
rect 1150 -1462 1179 -1461
rect 1220 -1462 1228 -1461
rect 107 -1464 507 -1463
rect 758 -1464 878 -1463
rect 926 -1464 976 -1463
rect 989 -1464 1403 -1463
rect 107 -1466 164 -1465
rect 240 -1466 458 -1465
rect 488 -1466 1375 -1465
rect 128 -1468 164 -1467
rect 247 -1468 846 -1467
rect 933 -1468 1000 -1467
rect 1017 -1468 1074 -1467
rect 1087 -1468 1095 -1467
rect 1122 -1468 1228 -1467
rect 128 -1470 871 -1469
rect 940 -1470 983 -1469
rect 1020 -1470 1494 -1469
rect 79 -1472 871 -1471
rect 947 -1472 1067 -1471
rect 1094 -1472 1109 -1471
rect 1150 -1472 1291 -1471
rect 1486 -1472 1494 -1471
rect 247 -1474 290 -1473
rect 331 -1474 619 -1473
rect 632 -1474 1123 -1473
rect 1283 -1474 1291 -1473
rect 1479 -1474 1487 -1473
rect 282 -1476 290 -1475
rect 331 -1476 423 -1475
rect 443 -1476 580 -1475
rect 695 -1476 1074 -1475
rect 1283 -1476 1501 -1475
rect 282 -1478 304 -1477
rect 345 -1478 500 -1477
rect 502 -1478 927 -1477
rect 954 -1478 1011 -1477
rect 1024 -1478 1067 -1477
rect 1472 -1478 1501 -1477
rect 303 -1480 311 -1479
rect 352 -1480 458 -1479
rect 709 -1480 1480 -1479
rect 9 -1482 353 -1481
rect 387 -1482 423 -1481
rect 450 -1482 486 -1481
rect 716 -1482 1403 -1481
rect 1451 -1482 1473 -1481
rect 9 -1484 682 -1483
rect 758 -1484 766 -1483
rect 982 -1484 997 -1483
rect 1010 -1484 1060 -1483
rect 1430 -1484 1452 -1483
rect 54 -1486 710 -1485
rect 765 -1486 923 -1485
rect 1024 -1486 1053 -1485
rect 1059 -1486 1172 -1485
rect 1395 -1486 1431 -1485
rect 58 -1488 717 -1487
rect 751 -1488 1053 -1487
rect 1367 -1488 1396 -1487
rect 58 -1490 815 -1489
rect 1031 -1490 1116 -1489
rect 212 -1492 451 -1491
rect 471 -1492 1172 -1491
rect 149 -1494 213 -1493
rect 310 -1494 475 -1493
rect 751 -1494 822 -1493
rect 1031 -1494 1158 -1493
rect 149 -1496 171 -1495
rect 387 -1496 430 -1495
rect 681 -1496 1158 -1495
rect 401 -1498 1109 -1497
rect 2 -1500 402 -1499
rect 415 -1500 1368 -1499
rect 2 -1502 143 -1501
rect 373 -1502 416 -1501
rect 429 -1502 892 -1501
rect 1038 -1502 1186 -1501
rect 142 -1504 157 -1503
rect 373 -1504 381 -1503
rect 814 -1504 1340 -1503
rect 86 -1506 381 -1505
rect 821 -1506 864 -1505
rect 891 -1506 913 -1505
rect 1101 -1506 1186 -1505
rect 86 -1508 605 -1507
rect 639 -1508 864 -1507
rect 1101 -1508 1200 -1507
rect 110 -1510 1340 -1509
rect 156 -1512 577 -1511
rect 604 -1512 626 -1511
rect 639 -1512 668 -1511
rect 786 -1512 913 -1511
rect 534 -1514 668 -1513
rect 786 -1514 829 -1513
rect 534 -1516 598 -1515
rect 611 -1516 626 -1515
rect 817 -1516 1200 -1515
rect 576 -1518 1126 -1517
rect 597 -1520 1438 -1519
rect 611 -1522 703 -1521
rect 828 -1522 1319 -1521
rect 702 -1524 738 -1523
rect 737 -1526 794 -1525
rect 394 -1528 794 -1527
rect 2 -1539 132 -1538
rect 142 -1539 174 -1538
rect 212 -1539 433 -1538
rect 471 -1539 668 -1538
rect 674 -1539 1326 -1538
rect 1349 -1539 1536 -1538
rect 2 -1541 276 -1540
rect 345 -1541 857 -1540
rect 859 -1541 1515 -1540
rect 9 -1543 13 -1542
rect 30 -1543 447 -1542
rect 474 -1543 818 -1542
rect 838 -1543 1221 -1542
rect 1325 -1543 1396 -1542
rect 9 -1545 486 -1544
rect 502 -1545 626 -1544
rect 639 -1545 755 -1544
rect 758 -1545 769 -1544
rect 782 -1545 850 -1544
rect 880 -1545 1186 -1544
rect 1220 -1545 1298 -1544
rect 30 -1547 136 -1546
rect 142 -1547 633 -1546
rect 639 -1547 654 -1546
rect 667 -1547 808 -1546
rect 849 -1547 864 -1546
rect 947 -1547 951 -1546
rect 992 -1547 1333 -1546
rect 44 -1549 276 -1548
rect 366 -1549 633 -1548
rect 653 -1549 717 -1548
rect 765 -1549 1172 -1548
rect 1185 -1549 1249 -1548
rect 1297 -1549 1375 -1548
rect 44 -1551 612 -1550
rect 618 -1551 675 -1550
rect 677 -1551 1522 -1550
rect 51 -1553 108 -1552
rect 128 -1553 213 -1552
rect 397 -1553 1403 -1552
rect 51 -1555 563 -1554
rect 579 -1555 731 -1554
rect 765 -1555 958 -1554
rect 996 -1555 1116 -1554
rect 1122 -1555 1410 -1554
rect 54 -1557 773 -1556
rect 863 -1557 920 -1556
rect 947 -1557 1004 -1556
rect 1073 -1557 1501 -1556
rect 65 -1559 503 -1558
rect 506 -1559 808 -1558
rect 919 -1559 983 -1558
rect 992 -1559 1074 -1558
rect 1115 -1559 1144 -1558
rect 1150 -1559 1154 -1558
rect 1171 -1559 1235 -1558
rect 1374 -1559 1452 -1558
rect 65 -1561 73 -1560
rect 75 -1561 528 -1560
rect 583 -1561 650 -1560
rect 681 -1561 1081 -1560
rect 1101 -1561 1144 -1560
rect 1150 -1561 1200 -1560
rect 1234 -1561 1417 -1560
rect 1451 -1561 1529 -1560
rect 58 -1563 528 -1562
rect 583 -1563 591 -1562
rect 600 -1563 752 -1562
rect 800 -1563 1081 -1562
rect 1101 -1563 1109 -1562
rect 1192 -1563 1249 -1562
rect 1283 -1563 1417 -1562
rect 58 -1565 374 -1564
rect 394 -1565 1410 -1564
rect 72 -1567 255 -1566
rect 373 -1567 458 -1566
rect 478 -1567 832 -1566
rect 982 -1567 1018 -1566
rect 1059 -1567 1109 -1566
rect 1192 -1567 1270 -1566
rect 1283 -1567 1312 -1566
rect 1402 -1567 1480 -1566
rect 79 -1569 115 -1568
rect 135 -1569 724 -1568
rect 730 -1569 794 -1568
rect 800 -1569 843 -1568
rect 989 -1569 1018 -1568
rect 1024 -1569 1270 -1568
rect 1311 -1569 1459 -1568
rect 82 -1571 493 -1570
rect 506 -1571 871 -1570
rect 898 -1571 1025 -1570
rect 1059 -1571 1396 -1570
rect 103 -1573 227 -1572
rect 380 -1573 479 -1572
rect 492 -1573 521 -1572
rect 590 -1573 703 -1572
rect 716 -1573 738 -1572
rect 751 -1573 1032 -1572
rect 107 -1575 339 -1574
rect 348 -1575 381 -1574
rect 394 -1575 556 -1574
rect 611 -1575 661 -1574
rect 681 -1575 696 -1574
rect 702 -1575 787 -1574
rect 793 -1575 1525 -1574
rect 114 -1577 262 -1576
rect 338 -1577 727 -1576
rect 737 -1577 1263 -1576
rect 145 -1579 745 -1578
rect 786 -1579 815 -1578
rect 870 -1579 927 -1578
rect 933 -1579 1032 -1578
rect 1262 -1579 1340 -1578
rect 128 -1581 934 -1580
rect 996 -1581 1077 -1580
rect 1255 -1581 1340 -1580
rect 156 -1583 626 -1582
rect 646 -1583 832 -1582
rect 898 -1583 976 -1582
rect 999 -1583 1130 -1582
rect 156 -1585 272 -1584
rect 408 -1585 773 -1584
rect 814 -1585 885 -1584
rect 975 -1585 1039 -1584
rect 1045 -1585 1256 -1584
rect 163 -1587 843 -1586
rect 884 -1587 962 -1586
rect 1038 -1587 1088 -1586
rect 1129 -1587 1158 -1586
rect 163 -1589 402 -1588
rect 429 -1589 465 -1588
rect 474 -1589 521 -1588
rect 555 -1589 1368 -1588
rect 170 -1591 440 -1590
rect 450 -1591 759 -1590
rect 817 -1591 927 -1590
rect 1045 -1591 1095 -1590
rect 1157 -1591 1214 -1590
rect 1367 -1591 1445 -1590
rect 170 -1593 206 -1592
rect 261 -1593 311 -1592
rect 352 -1593 402 -1592
rect 415 -1593 465 -1592
rect 499 -1593 962 -1592
rect 1094 -1593 1277 -1592
rect 100 -1595 206 -1594
rect 240 -1595 311 -1594
rect 331 -1595 416 -1594
rect 450 -1595 804 -1594
rect 1213 -1595 1431 -1594
rect 100 -1597 122 -1596
rect 177 -1597 486 -1596
rect 499 -1597 1333 -1596
rect 93 -1599 122 -1598
rect 177 -1599 598 -1598
rect 621 -1599 913 -1598
rect 1052 -1599 1431 -1598
rect 93 -1601 220 -1600
rect 240 -1601 388 -1600
rect 457 -1601 514 -1600
rect 646 -1601 1137 -1600
rect 1153 -1601 1200 -1600
rect 1276 -1601 1347 -1600
rect 86 -1603 514 -1602
rect 660 -1603 689 -1602
rect 695 -1603 780 -1602
rect 912 -1603 969 -1602
rect 989 -1603 1347 -1602
rect 86 -1605 283 -1604
rect 296 -1605 353 -1604
rect 369 -1605 388 -1604
rect 471 -1605 689 -1604
rect 723 -1605 822 -1604
rect 968 -1605 1165 -1604
rect 184 -1607 367 -1606
rect 684 -1607 1508 -1606
rect 184 -1609 234 -1608
rect 282 -1609 290 -1608
rect 331 -1609 566 -1608
rect 740 -1609 1088 -1608
rect 1136 -1609 1179 -1608
rect 191 -1611 409 -1610
rect 744 -1611 836 -1610
rect 1052 -1611 1319 -1610
rect 191 -1613 619 -1612
rect 709 -1613 1319 -1612
rect 198 -1615 255 -1614
rect 289 -1615 360 -1614
rect 548 -1615 710 -1614
rect 779 -1615 1067 -1614
rect 1164 -1615 1228 -1614
rect 198 -1617 269 -1616
rect 359 -1617 577 -1616
rect 821 -1617 829 -1616
rect 835 -1617 892 -1616
rect 905 -1617 1067 -1616
rect 1178 -1617 1242 -1616
rect 219 -1619 248 -1618
rect 541 -1619 577 -1618
rect 828 -1619 1123 -1618
rect 1227 -1619 1354 -1618
rect 226 -1621 269 -1620
rect 422 -1621 542 -1620
rect 548 -1621 605 -1620
rect 891 -1621 955 -1620
rect 1241 -1621 1305 -1620
rect 1353 -1621 1382 -1620
rect 233 -1623 559 -1622
rect 569 -1623 605 -1622
rect 905 -1623 941 -1622
rect 954 -1623 1361 -1622
rect 1381 -1623 1466 -1622
rect 247 -1625 444 -1624
rect 877 -1625 941 -1624
rect 1304 -1625 1389 -1624
rect 296 -1627 444 -1626
rect 877 -1627 1207 -1626
rect 1360 -1627 1438 -1626
rect 324 -1629 423 -1628
rect 436 -1629 570 -1628
rect 1206 -1629 1291 -1628
rect 1388 -1629 1473 -1628
rect 317 -1631 325 -1630
rect 1290 -1631 1424 -1630
rect 1437 -1631 1487 -1630
rect 37 -1633 318 -1632
rect 1423 -1633 1494 -1632
rect 37 -1635 563 -1634
rect 2 -1646 437 -1645
rect 446 -1646 475 -1645
rect 488 -1646 1207 -1645
rect 1283 -1646 1347 -1645
rect 1377 -1646 1452 -1645
rect 37 -1648 342 -1647
rect 429 -1648 444 -1647
rect 471 -1648 598 -1647
rect 621 -1648 766 -1647
rect 814 -1648 1018 -1647
rect 1206 -1648 1298 -1647
rect 37 -1650 388 -1649
rect 429 -1650 521 -1649
rect 555 -1650 668 -1649
rect 709 -1650 874 -1649
rect 877 -1650 1004 -1649
rect 1017 -1650 1151 -1649
rect 1283 -1650 1368 -1649
rect 65 -1652 587 -1651
rect 597 -1652 864 -1651
rect 877 -1652 1298 -1651
rect 1367 -1652 1431 -1651
rect 65 -1654 150 -1653
rect 163 -1654 419 -1653
rect 436 -1654 783 -1653
rect 828 -1654 1095 -1653
rect 1150 -1654 1200 -1653
rect 72 -1656 507 -1655
rect 513 -1656 741 -1655
rect 744 -1656 776 -1655
rect 817 -1656 1200 -1655
rect 82 -1658 626 -1657
rect 635 -1658 787 -1657
rect 828 -1658 934 -1657
rect 1094 -1658 1305 -1657
rect 128 -1660 633 -1659
rect 653 -1660 657 -1659
rect 667 -1660 675 -1659
rect 709 -1660 717 -1659
rect 719 -1660 969 -1659
rect 1006 -1660 1305 -1659
rect 128 -1662 136 -1661
rect 149 -1662 234 -1661
rect 240 -1662 370 -1661
rect 387 -1662 493 -1661
rect 513 -1662 524 -1661
rect 555 -1662 591 -1661
rect 604 -1662 675 -1661
rect 723 -1662 881 -1661
rect 933 -1662 1081 -1661
rect 9 -1664 370 -1663
rect 471 -1664 738 -1663
rect 751 -1664 1347 -1663
rect 9 -1666 94 -1665
rect 121 -1666 136 -1665
rect 142 -1666 234 -1665
rect 240 -1666 255 -1665
rect 303 -1666 346 -1665
rect 359 -1666 633 -1665
rect 653 -1666 689 -1665
rect 751 -1666 822 -1665
rect 863 -1666 892 -1665
rect 968 -1666 1039 -1665
rect 1080 -1666 1186 -1665
rect 93 -1668 549 -1667
rect 562 -1668 1256 -1667
rect 114 -1670 304 -1669
rect 310 -1670 521 -1669
rect 527 -1670 563 -1669
rect 565 -1670 808 -1669
rect 821 -1670 885 -1669
rect 891 -1670 948 -1669
rect 1038 -1670 1144 -1669
rect 1255 -1670 1291 -1669
rect 79 -1672 115 -1671
rect 121 -1672 157 -1671
rect 163 -1672 185 -1671
rect 198 -1672 272 -1671
rect 310 -1672 402 -1671
rect 408 -1672 549 -1671
rect 590 -1672 661 -1671
rect 758 -1672 832 -1671
rect 845 -1672 1186 -1671
rect 1290 -1672 1375 -1671
rect 58 -1674 157 -1673
rect 177 -1674 500 -1673
rect 604 -1674 780 -1673
rect 786 -1674 990 -1673
rect 58 -1676 542 -1675
rect 625 -1676 640 -1675
rect 656 -1676 689 -1675
rect 758 -1676 1032 -1675
rect 79 -1678 325 -1677
rect 345 -1678 416 -1677
rect 485 -1678 738 -1677
rect 765 -1678 962 -1677
rect 1031 -1678 1158 -1677
rect 110 -1680 409 -1679
rect 492 -1680 650 -1679
rect 660 -1680 731 -1679
rect 779 -1680 836 -1679
rect 880 -1680 1011 -1679
rect 1157 -1680 1242 -1679
rect 110 -1682 843 -1681
rect 884 -1682 906 -1681
rect 926 -1682 1144 -1681
rect 142 -1684 696 -1683
rect 730 -1684 850 -1683
rect 905 -1684 1350 -1683
rect 177 -1686 755 -1685
rect 835 -1686 871 -1685
rect 926 -1686 1102 -1685
rect 184 -1688 426 -1687
rect 506 -1688 1242 -1687
rect 198 -1690 955 -1689
rect 961 -1690 983 -1689
rect 1010 -1690 1172 -1689
rect 205 -1692 528 -1691
rect 576 -1692 696 -1691
rect 842 -1692 1228 -1691
rect 205 -1694 262 -1693
rect 268 -1694 500 -1693
rect 576 -1694 1004 -1693
rect 1101 -1694 1221 -1693
rect 1227 -1694 1410 -1693
rect 219 -1696 262 -1695
rect 268 -1696 318 -1695
rect 359 -1696 465 -1695
rect 611 -1696 640 -1695
rect 849 -1696 920 -1695
rect 947 -1696 1046 -1695
rect 1220 -1696 1319 -1695
rect 219 -1698 797 -1697
rect 870 -1698 1235 -1697
rect 1248 -1698 1319 -1697
rect 254 -1700 416 -1699
rect 464 -1700 479 -1699
rect 611 -1700 857 -1699
rect 901 -1700 1249 -1699
rect 289 -1702 318 -1701
rect 366 -1702 745 -1701
rect 856 -1702 899 -1701
rect 919 -1702 1088 -1701
rect 1234 -1702 1389 -1701
rect 212 -1704 367 -1703
rect 394 -1704 542 -1703
rect 898 -1704 941 -1703
rect 954 -1704 1130 -1703
rect 131 -1706 1130 -1705
rect 212 -1708 276 -1707
rect 282 -1708 290 -1707
rect 296 -1708 325 -1707
rect 394 -1708 423 -1707
rect 478 -1708 535 -1707
rect 940 -1708 976 -1707
rect 982 -1708 1074 -1707
rect 1087 -1708 1193 -1707
rect 75 -1710 297 -1709
rect 401 -1710 570 -1709
rect 975 -1710 1123 -1709
rect 1192 -1710 1263 -1709
rect 75 -1712 724 -1711
rect 996 -1712 1172 -1711
rect 1262 -1712 1333 -1711
rect 107 -1714 276 -1713
rect 282 -1714 374 -1713
rect 380 -1714 570 -1713
rect 996 -1714 1109 -1713
rect 1332 -1714 1403 -1713
rect 72 -1716 381 -1715
rect 422 -1716 584 -1715
rect 1024 -1716 1410 -1715
rect 107 -1718 451 -1717
rect 502 -1718 1025 -1717
rect 1045 -1718 1165 -1717
rect 1402 -1718 1424 -1717
rect 247 -1720 374 -1719
rect 534 -1720 794 -1719
rect 1052 -1720 1123 -1719
rect 1164 -1720 1277 -1719
rect 1423 -1720 1438 -1719
rect 145 -1722 248 -1721
rect 331 -1722 451 -1721
rect 793 -1722 1312 -1721
rect 331 -1724 353 -1723
rect 810 -1724 1053 -1723
rect 1066 -1724 1389 -1723
rect 338 -1726 353 -1725
rect 992 -1726 1312 -1725
rect 30 -1728 339 -1727
rect 992 -1728 1340 -1727
rect 16 -1730 31 -1729
rect 646 -1730 1340 -1729
rect 16 -1732 101 -1731
rect 646 -1732 682 -1731
rect 1066 -1732 1116 -1731
rect 1276 -1732 1361 -1731
rect 100 -1734 192 -1733
rect 530 -1734 1116 -1733
rect 191 -1736 510 -1735
rect 681 -1736 703 -1735
rect 716 -1736 1361 -1735
rect 702 -1738 773 -1737
rect 1073 -1738 1179 -1737
rect 772 -1740 1270 -1739
rect 1108 -1742 1137 -1741
rect 1178 -1742 1382 -1741
rect 1136 -1744 1326 -1743
rect 1374 -1744 1382 -1743
rect 618 -1746 1326 -1745
rect 44 -1748 619 -1747
rect 1213 -1748 1270 -1747
rect 44 -1750 227 -1749
rect 1213 -1750 1396 -1749
rect 86 -1752 227 -1751
rect 1353 -1752 1396 -1751
rect 86 -1754 171 -1753
rect 1353 -1754 1417 -1753
rect 170 -1756 458 -1755
rect 912 -1756 1417 -1755
rect 457 -1758 584 -1757
rect 912 -1758 1060 -1757
rect 1059 -1760 1371 -1759
rect 2 -1771 591 -1770
rect 667 -1771 843 -1770
rect 877 -1771 1158 -1770
rect 1255 -1771 1259 -1770
rect 1360 -1771 1371 -1770
rect 1377 -1771 1396 -1770
rect 19 -1773 535 -1772
rect 562 -1773 591 -1772
rect 667 -1773 682 -1772
rect 684 -1773 787 -1772
rect 793 -1773 836 -1772
rect 842 -1773 864 -1772
rect 887 -1773 969 -1772
rect 1003 -1773 1067 -1772
rect 1255 -1773 1263 -1772
rect 1367 -1773 1403 -1772
rect 61 -1775 1228 -1774
rect 1346 -1775 1368 -1774
rect 1381 -1775 1431 -1774
rect 72 -1777 797 -1776
rect 800 -1777 808 -1776
rect 814 -1777 836 -1776
rect 849 -1777 878 -1776
rect 898 -1777 1193 -1776
rect 1339 -1777 1347 -1776
rect 1353 -1777 1382 -1776
rect 30 -1779 73 -1778
rect 75 -1779 143 -1778
rect 247 -1779 881 -1778
rect 898 -1779 941 -1778
rect 968 -1779 1060 -1778
rect 1066 -1779 1109 -1778
rect 1332 -1779 1340 -1778
rect 1353 -1779 1375 -1778
rect 23 -1781 31 -1780
rect 89 -1781 311 -1780
rect 324 -1781 370 -1780
rect 373 -1781 503 -1780
rect 513 -1781 787 -1780
rect 793 -1781 1396 -1780
rect 23 -1783 633 -1782
rect 635 -1783 1193 -1782
rect 1234 -1783 1333 -1782
rect 51 -1785 633 -1784
rect 691 -1785 1249 -1784
rect 1325 -1785 1375 -1784
rect 51 -1787 122 -1786
rect 138 -1787 416 -1786
rect 436 -1787 440 -1786
rect 464 -1787 510 -1786
rect 513 -1787 542 -1786
rect 569 -1787 815 -1786
rect 849 -1787 857 -1786
rect 863 -1787 892 -1786
rect 908 -1787 1151 -1786
rect 1178 -1787 1326 -1786
rect 58 -1789 122 -1788
rect 191 -1789 374 -1788
rect 380 -1789 563 -1788
rect 569 -1789 766 -1788
rect 800 -1789 1011 -1788
rect 1129 -1789 1151 -1788
rect 1234 -1789 1389 -1788
rect 9 -1791 59 -1790
rect 82 -1791 892 -1790
rect 926 -1791 1158 -1790
rect 1241 -1791 1249 -1790
rect 9 -1793 157 -1792
rect 191 -1793 269 -1792
rect 275 -1793 664 -1792
rect 716 -1793 1109 -1792
rect 1136 -1793 1242 -1792
rect 37 -1795 157 -1794
rect 212 -1795 269 -1794
rect 289 -1795 300 -1794
rect 310 -1795 423 -1794
rect 436 -1795 458 -1794
rect 464 -1795 696 -1794
rect 719 -1795 983 -1794
rect 989 -1795 1130 -1794
rect 107 -1797 398 -1796
rect 415 -1797 605 -1796
rect 611 -1797 808 -1796
rect 810 -1797 1389 -1796
rect 100 -1799 108 -1798
rect 114 -1799 143 -1798
rect 212 -1799 367 -1798
rect 380 -1799 444 -1798
rect 527 -1799 752 -1798
rect 765 -1799 780 -1798
rect 803 -1799 1228 -1798
rect 1258 -1799 1263 -1798
rect 100 -1801 185 -1800
rect 226 -1801 276 -1800
rect 296 -1801 367 -1800
rect 387 -1801 521 -1800
rect 527 -1801 703 -1800
rect 719 -1801 829 -1800
rect 856 -1801 885 -1800
rect 926 -1801 962 -1800
rect 989 -1801 1172 -1800
rect 65 -1803 185 -1802
rect 247 -1803 255 -1802
rect 261 -1803 486 -1802
rect 534 -1803 731 -1802
rect 737 -1803 755 -1802
rect 779 -1803 1221 -1802
rect 65 -1805 87 -1804
rect 114 -1805 150 -1804
rect 163 -1805 227 -1804
rect 233 -1805 262 -1804
rect 296 -1805 1063 -1804
rect 1094 -1805 1221 -1804
rect 135 -1807 150 -1806
rect 163 -1807 171 -1806
rect 233 -1807 346 -1806
rect 352 -1807 444 -1806
rect 485 -1807 885 -1806
rect 919 -1807 1172 -1806
rect 37 -1809 136 -1808
rect 240 -1809 255 -1808
rect 324 -1809 577 -1808
rect 604 -1809 619 -1808
rect 695 -1809 724 -1808
rect 737 -1809 1018 -1808
rect 1087 -1809 1095 -1808
rect 1122 -1809 1137 -1808
rect 44 -1811 346 -1810
rect 352 -1811 472 -1810
rect 488 -1811 577 -1810
rect 611 -1811 647 -1810
rect 702 -1811 710 -1810
rect 723 -1811 937 -1810
rect 940 -1811 1417 -1810
rect 44 -1813 409 -1812
rect 492 -1813 731 -1812
rect 744 -1813 983 -1812
rect 996 -1813 1004 -1812
rect 1006 -1813 1319 -1812
rect 93 -1815 171 -1814
rect 240 -1815 451 -1814
rect 530 -1815 745 -1814
rect 751 -1815 962 -1814
rect 975 -1815 1018 -1814
rect 1073 -1815 1088 -1814
rect 1311 -1815 1319 -1814
rect 93 -1817 419 -1816
rect 450 -1817 776 -1816
rect 821 -1817 829 -1816
rect 870 -1817 1417 -1816
rect 128 -1819 472 -1818
rect 506 -1819 976 -1818
rect 996 -1819 1144 -1818
rect 1304 -1819 1312 -1818
rect 128 -1821 594 -1820
rect 597 -1821 822 -1820
rect 870 -1821 913 -1820
rect 919 -1821 1081 -1820
rect 1115 -1821 1144 -1820
rect 1297 -1821 1305 -1820
rect 317 -1823 409 -1822
rect 478 -1823 507 -1822
rect 541 -1823 549 -1822
rect 555 -1823 598 -1822
rect 618 -1823 1025 -1822
rect 1045 -1823 1074 -1822
rect 1290 -1823 1298 -1822
rect 282 -1825 318 -1824
rect 331 -1825 423 -1824
rect 432 -1825 1046 -1824
rect 1052 -1825 1081 -1824
rect 1283 -1825 1291 -1824
rect 282 -1827 360 -1826
rect 387 -1827 654 -1826
rect 681 -1827 1116 -1826
rect 219 -1829 360 -1828
rect 401 -1829 549 -1828
rect 555 -1829 689 -1828
rect 709 -1829 906 -1828
rect 933 -1829 1025 -1828
rect 1031 -1829 1053 -1828
rect 1101 -1829 1284 -1828
rect 79 -1831 220 -1830
rect 303 -1831 332 -1830
rect 338 -1831 493 -1830
rect 558 -1831 913 -1830
rect 1010 -1831 1207 -1830
rect 16 -1833 80 -1832
rect 303 -1833 395 -1832
rect 401 -1833 846 -1832
rect 873 -1833 1123 -1832
rect 1185 -1833 1207 -1832
rect 86 -1835 1186 -1834
rect 338 -1837 584 -1836
rect 586 -1837 906 -1836
rect 1031 -1837 1039 -1836
rect 1101 -1837 1410 -1836
rect 341 -1839 1214 -1838
rect 394 -1841 1361 -1840
rect 478 -1843 500 -1842
rect 583 -1843 640 -1842
rect 653 -1843 759 -1842
rect 901 -1843 1410 -1842
rect 289 -1845 500 -1844
rect 625 -1845 647 -1844
rect 688 -1845 1179 -1844
rect 1199 -1845 1214 -1844
rect 625 -1847 661 -1846
rect 716 -1847 759 -1846
rect 954 -1847 1200 -1846
rect 639 -1849 934 -1848
rect 947 -1849 955 -1848
rect 1038 -1849 1277 -1848
rect 572 -1851 948 -1850
rect 1269 -1851 1277 -1850
rect 660 -1853 1403 -1852
rect 772 -1855 1270 -1854
rect 429 -1857 773 -1856
rect 2 -1868 6 -1867
rect 9 -1868 398 -1867
rect 432 -1868 745 -1867
rect 751 -1868 1284 -1867
rect 1395 -1868 1424 -1867
rect 2 -1870 52 -1869
rect 100 -1870 300 -1869
rect 373 -1870 559 -1869
rect 565 -1870 913 -1869
rect 933 -1870 1382 -1869
rect 9 -1872 262 -1871
rect 282 -1872 346 -1871
rect 471 -1872 615 -1871
rect 618 -1872 773 -1871
rect 775 -1872 969 -1871
rect 1062 -1872 1263 -1871
rect 19 -1874 76 -1873
rect 100 -1874 115 -1873
rect 128 -1874 937 -1873
rect 968 -1874 976 -1873
rect 1234 -1874 1396 -1873
rect 26 -1876 31 -1875
rect 37 -1876 395 -1875
rect 401 -1876 472 -1875
rect 499 -1876 598 -1875
rect 618 -1876 804 -1875
rect 856 -1876 906 -1875
rect 912 -1876 927 -1875
rect 933 -1876 1004 -1875
rect 1066 -1876 1235 -1875
rect 30 -1878 458 -1877
rect 502 -1878 1382 -1877
rect 37 -1880 1200 -1879
rect 44 -1882 510 -1881
rect 523 -1882 1207 -1881
rect 44 -1884 605 -1883
rect 646 -1884 664 -1883
rect 681 -1884 1399 -1883
rect 51 -1886 213 -1885
rect 219 -1886 402 -1885
rect 527 -1886 598 -1885
rect 604 -1886 1060 -1885
rect 1199 -1886 1242 -1885
rect 58 -1888 857 -1887
rect 884 -1888 1431 -1887
rect 58 -1890 514 -1889
rect 555 -1890 626 -1889
rect 660 -1890 1158 -1889
rect 1206 -1890 1298 -1889
rect 40 -1892 1158 -1891
rect 1241 -1892 1256 -1891
rect 1297 -1892 1333 -1891
rect 61 -1894 262 -1893
rect 282 -1894 409 -1893
rect 513 -1894 724 -1893
rect 726 -1894 1263 -1893
rect 1332 -1894 1368 -1893
rect 79 -1896 213 -1895
rect 219 -1896 353 -1895
rect 355 -1896 976 -1895
rect 996 -1896 1067 -1895
rect 1122 -1896 1368 -1895
rect 79 -1898 143 -1897
rect 170 -1898 643 -1897
rect 688 -1898 1172 -1897
rect 1255 -1898 1312 -1897
rect 89 -1900 647 -1899
rect 660 -1900 689 -1899
rect 691 -1900 1172 -1899
rect 1311 -1900 1340 -1899
rect 121 -1902 500 -1901
rect 625 -1902 710 -1901
rect 737 -1902 997 -1901
rect 1003 -1902 1074 -1901
rect 1122 -1902 1221 -1901
rect 1339 -1902 1389 -1901
rect 121 -1904 507 -1903
rect 702 -1904 720 -1903
rect 737 -1904 808 -1903
rect 870 -1904 885 -1903
rect 926 -1904 1018 -1903
rect 1038 -1904 1221 -1903
rect 1388 -1904 1417 -1903
rect 128 -1906 444 -1905
rect 506 -1906 1249 -1905
rect 135 -1908 1144 -1907
rect 1248 -1908 1305 -1907
rect 135 -1910 150 -1909
rect 170 -1910 1375 -1909
rect 142 -1912 297 -1911
rect 338 -1912 1018 -1911
rect 1038 -1912 1109 -1911
rect 1143 -1912 1193 -1911
rect 1374 -1912 1410 -1911
rect 149 -1914 668 -1913
rect 716 -1914 1305 -1913
rect 205 -1916 570 -1915
rect 611 -1916 703 -1915
rect 716 -1916 759 -1915
rect 772 -1916 829 -1915
rect 870 -1916 892 -1915
rect 1059 -1916 1130 -1915
rect 1192 -1916 1277 -1915
rect 205 -1918 332 -1917
rect 338 -1918 367 -1917
rect 387 -1918 664 -1917
rect 744 -1918 822 -1917
rect 828 -1918 864 -1917
rect 891 -1918 948 -1917
rect 1108 -1918 1403 -1917
rect 93 -1920 864 -1919
rect 898 -1920 948 -1919
rect 1024 -1920 1403 -1919
rect 93 -1922 199 -1921
rect 233 -1922 430 -1921
rect 492 -1922 668 -1921
rect 751 -1922 1074 -1921
rect 1129 -1922 1326 -1921
rect 198 -1924 787 -1923
rect 800 -1924 955 -1923
rect 1024 -1924 1088 -1923
rect 1276 -1924 1319 -1923
rect 1325 -1924 1354 -1923
rect 86 -1926 1354 -1925
rect 86 -1928 349 -1927
rect 352 -1928 388 -1927
rect 408 -1928 528 -1927
rect 569 -1928 577 -1927
rect 611 -1928 710 -1927
rect 723 -1928 787 -1927
rect 800 -1928 941 -1927
rect 954 -1928 1046 -1927
rect 1087 -1928 1270 -1927
rect 1318 -1928 1347 -1927
rect 138 -1930 1046 -1929
rect 1346 -1930 1361 -1929
rect 233 -1932 633 -1931
rect 653 -1932 899 -1931
rect 940 -1932 1116 -1931
rect 240 -1934 685 -1933
rect 754 -1934 878 -1933
rect 989 -1934 1361 -1933
rect 240 -1936 423 -1935
rect 429 -1936 909 -1935
rect 989 -1936 1053 -1935
rect 1115 -1936 1186 -1935
rect 191 -1938 423 -1937
rect 464 -1938 493 -1937
rect 520 -1938 577 -1937
rect 674 -1938 755 -1937
rect 758 -1938 766 -1937
rect 782 -1938 1102 -1937
rect 1150 -1938 1186 -1937
rect 72 -1940 192 -1939
rect 247 -1940 395 -1939
rect 464 -1940 794 -1939
rect 807 -1940 1284 -1939
rect 72 -1942 174 -1941
rect 268 -1942 444 -1941
rect 485 -1942 794 -1941
rect 821 -1942 850 -1941
rect 1010 -1942 1151 -1941
rect 107 -1944 248 -1943
rect 268 -1944 276 -1943
rect 289 -1944 633 -1943
rect 765 -1944 815 -1943
rect 835 -1944 878 -1943
rect 1010 -1944 1081 -1943
rect 1101 -1944 1179 -1943
rect 16 -1946 108 -1945
rect 163 -1946 290 -1945
rect 296 -1946 542 -1945
rect 572 -1946 815 -1945
rect 835 -1946 843 -1945
rect 1052 -1946 1095 -1945
rect 1178 -1946 1228 -1945
rect 16 -1948 24 -1947
rect 163 -1948 594 -1947
rect 842 -1948 962 -1947
rect 1080 -1948 1137 -1947
rect 23 -1950 1214 -1949
rect 229 -1952 276 -1951
rect 310 -1952 486 -1951
rect 579 -1952 675 -1951
rect 705 -1952 1137 -1951
rect 1213 -1952 1291 -1951
rect 310 -1954 325 -1953
rect 331 -1954 549 -1953
rect 887 -1954 1291 -1953
rect 65 -1956 325 -1955
rect 345 -1956 517 -1955
rect 548 -1956 563 -1955
rect 961 -1956 983 -1955
rect 1094 -1956 1165 -1955
rect 65 -1958 115 -1957
rect 317 -1958 563 -1957
rect 779 -1958 1165 -1957
rect 317 -1960 437 -1959
rect 478 -1960 542 -1959
rect 681 -1960 780 -1959
rect 982 -1960 1032 -1959
rect 359 -1962 458 -1961
rect 919 -1962 1032 -1961
rect 359 -1964 451 -1963
rect 590 -1964 920 -1963
rect 177 -1966 451 -1965
rect 583 -1966 591 -1965
rect 177 -1968 227 -1967
rect 366 -1968 640 -1967
rect 184 -1970 227 -1969
rect 373 -1970 1270 -1969
rect 68 -1972 185 -1971
rect 380 -1972 521 -1971
rect 583 -1972 1228 -1971
rect 156 -1974 381 -1973
rect 415 -1974 479 -1973
rect 639 -1974 654 -1973
rect 5 -1976 416 -1975
rect 436 -1976 853 -1975
rect 156 -1978 696 -1977
rect 695 -1980 731 -1979
rect 534 -1982 731 -1981
rect 411 -1984 535 -1983
rect 2 -1995 38 -1994
rect 51 -1995 661 -1994
rect 663 -1995 997 -1994
rect 1139 -1995 1368 -1994
rect 5 -1997 192 -1996
rect 205 -1997 321 -1996
rect 324 -1997 377 -1996
rect 408 -1997 1263 -1996
rect 37 -1999 339 -1998
rect 408 -1999 542 -1998
rect 579 -1999 1186 -1998
rect 1262 -1999 1284 -1998
rect 51 -2001 262 -2000
rect 268 -2001 356 -2000
rect 373 -2001 1186 -2000
rect 1283 -2001 1326 -2000
rect 58 -2003 489 -2002
rect 502 -2003 1305 -2002
rect 1325 -2003 1389 -2002
rect 58 -2005 248 -2004
rect 261 -2005 388 -2004
rect 411 -2005 1235 -2004
rect 65 -2007 290 -2006
rect 334 -2007 1277 -2006
rect 65 -2009 304 -2008
rect 338 -2009 395 -2008
rect 415 -2009 542 -2008
rect 614 -2009 1242 -2008
rect 68 -2011 325 -2010
rect 373 -2011 479 -2010
rect 513 -2011 1291 -2010
rect 72 -2013 1228 -2012
rect 1290 -2013 1333 -2012
rect 72 -2015 332 -2014
rect 387 -2015 486 -2014
rect 513 -2015 626 -2014
rect 639 -2015 1081 -2014
rect 1108 -2015 1305 -2014
rect 93 -2017 206 -2016
rect 268 -2017 430 -2016
rect 453 -2017 1242 -2016
rect 93 -2019 640 -2018
rect 646 -2019 661 -2018
rect 691 -2019 1361 -2018
rect 96 -2021 101 -2020
rect 107 -2021 248 -2020
rect 289 -2021 437 -2020
rect 478 -2021 528 -2020
rect 604 -2021 626 -2020
rect 646 -2021 682 -2020
rect 705 -2021 773 -2020
rect 782 -2021 822 -2020
rect 849 -2021 934 -2020
rect 947 -2021 1144 -2020
rect 1213 -2021 1277 -2020
rect 100 -2023 174 -2022
rect 177 -2023 332 -2022
rect 415 -2023 493 -2022
rect 516 -2023 766 -2022
rect 807 -2023 1046 -2022
rect 1059 -2023 1081 -2022
rect 1129 -2023 1235 -2022
rect 121 -2025 493 -2024
rect 499 -2025 808 -2024
rect 821 -2025 1200 -2024
rect 1206 -2025 1214 -2024
rect 1227 -2025 1256 -2024
rect 23 -2027 122 -2026
rect 128 -2027 682 -2026
rect 726 -2027 1403 -2026
rect 16 -2029 129 -2028
rect 131 -2029 395 -2028
rect 422 -2029 510 -2028
rect 520 -2029 591 -2028
rect 621 -2029 1354 -2028
rect 16 -2031 241 -2030
rect 296 -2031 500 -2030
rect 520 -2031 818 -2030
rect 849 -2031 857 -2030
rect 912 -2031 1109 -2030
rect 1129 -2031 1137 -2030
rect 1143 -2031 1165 -2030
rect 1199 -2031 1221 -2030
rect 23 -2033 157 -2032
rect 163 -2033 227 -2032
rect 296 -2033 612 -2032
rect 730 -2033 734 -2032
rect 737 -2033 773 -2032
rect 779 -2033 1165 -2032
rect 1206 -2033 1319 -2032
rect 9 -2035 164 -2034
rect 166 -2035 1018 -2034
rect 1059 -2035 1095 -2034
rect 1220 -2035 1249 -2034
rect 1318 -2035 1382 -2034
rect 9 -2037 1256 -2036
rect 135 -2039 157 -2038
rect 173 -2039 213 -2038
rect 219 -2039 241 -2038
rect 303 -2039 311 -2038
rect 422 -2039 451 -2038
rect 527 -2039 549 -2038
rect 555 -2039 605 -2038
rect 716 -2039 738 -2038
rect 754 -2039 899 -2038
rect 933 -2039 993 -2038
rect 996 -2039 1123 -2038
rect 1248 -2039 1270 -2038
rect 110 -2041 213 -2040
rect 219 -2041 535 -2040
rect 548 -2041 783 -2040
rect 842 -2041 913 -2040
rect 968 -2041 1046 -2040
rect 1094 -2041 1193 -2040
rect 1269 -2041 1312 -2040
rect 135 -2043 671 -2042
rect 730 -2043 801 -2042
rect 828 -2043 843 -2042
rect 852 -2043 906 -2042
rect 971 -2043 1298 -2042
rect 1311 -2043 1375 -2042
rect 142 -2045 311 -2044
rect 429 -2045 825 -2044
rect 856 -2045 955 -2044
rect 1017 -2045 1088 -2044
rect 1101 -2045 1193 -2044
rect 1297 -2045 1340 -2044
rect 142 -2047 360 -2046
rect 436 -2047 472 -2046
rect 485 -2047 717 -2046
rect 765 -2047 864 -2046
rect 870 -2047 899 -2046
rect 954 -2047 990 -2046
rect 1073 -2047 1088 -2046
rect 1101 -2047 1116 -2046
rect 30 -2049 360 -2048
rect 443 -2049 451 -2048
rect 457 -2049 472 -2048
rect 555 -2049 587 -2048
rect 590 -2049 633 -2048
rect 779 -2049 1347 -2048
rect 30 -2051 41 -2050
rect 170 -2051 444 -2050
rect 457 -2051 465 -2050
rect 569 -2051 612 -2050
rect 786 -2051 801 -2050
rect 863 -2051 895 -2050
rect 1066 -2051 1074 -2050
rect 75 -2053 171 -2052
rect 177 -2053 724 -2052
rect 744 -2053 787 -2052
rect 870 -2053 1116 -2052
rect 191 -2055 619 -2054
rect 674 -2055 724 -2054
rect 733 -2055 745 -2054
rect 891 -2055 906 -2054
rect 149 -2057 619 -2056
rect 674 -2057 696 -2056
rect 149 -2059 1158 -2058
rect 198 -2061 465 -2060
rect 506 -2061 1067 -2060
rect 184 -2063 199 -2062
rect 226 -2063 752 -2062
rect 184 -2065 255 -2064
rect 562 -2065 1158 -2064
rect 229 -2067 507 -2066
rect 562 -2067 976 -2066
rect 233 -2069 535 -2068
rect 569 -2069 668 -2068
rect 695 -2069 794 -2068
rect 975 -2069 983 -2068
rect 86 -2071 234 -2070
rect 254 -2071 283 -2070
rect 576 -2071 633 -2070
rect 667 -2071 1151 -2070
rect 86 -2073 108 -2072
rect 282 -2073 346 -2072
rect 576 -2073 962 -2072
rect 982 -2073 1396 -2072
rect 345 -2075 402 -2074
rect 579 -2075 948 -2074
rect 1150 -2075 1172 -2074
rect 401 -2077 643 -2076
rect 751 -2077 759 -2076
rect 793 -2077 1004 -2076
rect 1171 -2077 1179 -2076
rect 597 -2079 829 -2078
rect 835 -2079 1004 -2078
rect 523 -2081 598 -2080
rect 688 -2081 759 -2080
rect 814 -2081 836 -2080
rect 926 -2081 962 -2080
rect 583 -2083 689 -2082
rect 709 -2083 1179 -2082
rect 380 -2085 710 -2084
rect 814 -2085 1053 -2084
rect 44 -2087 381 -2086
rect 583 -2087 654 -2086
rect 919 -2087 927 -2086
rect 940 -2087 1053 -2086
rect 2 -2089 654 -2088
rect 940 -2089 1039 -2088
rect 44 -2091 80 -2090
rect 352 -2091 920 -2090
rect 968 -2091 1039 -2090
rect 79 -2093 318 -2092
rect 275 -2095 353 -2094
rect 275 -2097 367 -2096
rect 317 -2099 1123 -2098
rect 366 -2101 703 -2100
rect 702 -2103 811 -2102
rect 9 -2114 45 -2113
rect 51 -2114 668 -2113
rect 765 -2114 769 -2113
rect 793 -2114 892 -2113
rect 936 -2114 976 -2113
rect 989 -2114 1046 -2113
rect 1115 -2114 1263 -2113
rect 9 -2116 472 -2115
rect 478 -2116 692 -2115
rect 695 -2116 794 -2115
rect 814 -2116 906 -2115
rect 968 -2116 1116 -2115
rect 1118 -2116 1214 -2115
rect 1262 -2116 1284 -2115
rect 30 -2118 45 -2117
rect 51 -2118 661 -2117
rect 667 -2118 738 -2117
rect 765 -2118 836 -2117
rect 891 -2118 1053 -2117
rect 1139 -2118 1277 -2117
rect 75 -2120 710 -2119
rect 814 -2120 899 -2119
rect 905 -2120 955 -2119
rect 985 -2120 1284 -2119
rect 107 -2122 1193 -2121
rect 1213 -2122 1242 -2121
rect 1276 -2122 1291 -2121
rect 107 -2124 412 -2123
rect 450 -2124 1081 -2123
rect 1192 -2124 1221 -2123
rect 1241 -2124 1256 -2123
rect 1290 -2124 1298 -2123
rect 40 -2126 1221 -2125
rect 1297 -2126 1319 -2125
rect 110 -2128 269 -2127
rect 320 -2128 486 -2127
rect 488 -2128 899 -2127
rect 989 -2128 1011 -2127
rect 1045 -2128 1088 -2127
rect 1206 -2128 1256 -2127
rect 131 -2130 157 -2129
rect 170 -2130 178 -2129
rect 184 -2130 335 -2129
rect 345 -2130 556 -2129
rect 579 -2130 682 -2129
rect 695 -2130 983 -2129
rect 992 -2130 1312 -2129
rect 37 -2132 185 -2131
rect 191 -2132 678 -2131
rect 821 -2132 850 -2131
rect 856 -2132 955 -2131
rect 996 -2132 1088 -2131
rect 1206 -2132 1235 -2131
rect 79 -2134 178 -2133
rect 191 -2134 318 -2133
rect 331 -2134 976 -2133
rect 996 -2134 1032 -2133
rect 1080 -2134 1123 -2133
rect 79 -2136 542 -2135
rect 555 -2136 654 -2135
rect 660 -2136 731 -2135
rect 849 -2136 885 -2135
rect 940 -2136 1011 -2135
rect 1031 -2136 1039 -2135
rect 138 -2138 157 -2137
rect 163 -2138 983 -2137
rect 1003 -2138 1312 -2137
rect 170 -2140 622 -2139
rect 628 -2140 1235 -2139
rect 205 -2142 209 -2141
rect 219 -2142 972 -2141
rect 1003 -2142 1025 -2141
rect 1038 -2142 1095 -2141
rect 205 -2144 234 -2143
rect 247 -2144 472 -2143
rect 478 -2144 640 -2143
rect 649 -2144 745 -2143
rect 884 -2144 920 -2143
rect 1094 -2144 1130 -2143
rect 247 -2146 300 -2145
rect 317 -2146 339 -2145
rect 352 -2146 426 -2145
rect 450 -2146 783 -2145
rect 1129 -2146 1165 -2145
rect 5 -2148 353 -2147
rect 373 -2148 682 -2147
rect 702 -2148 857 -2147
rect 1164 -2148 1186 -2147
rect 72 -2150 339 -2149
rect 394 -2150 969 -2149
rect 1185 -2150 1200 -2149
rect 72 -2152 150 -2151
rect 254 -2152 349 -2151
rect 394 -2152 423 -2151
rect 464 -2152 710 -2151
rect 730 -2152 825 -2151
rect 1199 -2152 1228 -2151
rect 2 -2154 150 -2153
rect 261 -2154 269 -2153
rect 310 -2154 374 -2153
rect 397 -2154 454 -2153
rect 464 -2154 531 -2153
rect 541 -2154 591 -2153
rect 597 -2154 738 -2153
rect 744 -2154 948 -2153
rect 1227 -2154 1249 -2153
rect 65 -2156 255 -2155
rect 261 -2156 276 -2155
rect 296 -2156 311 -2155
rect 404 -2156 689 -2155
rect 702 -2156 724 -2155
rect 768 -2156 836 -2155
rect 1248 -2156 1270 -2155
rect 65 -2158 87 -2157
rect 275 -2158 304 -2157
rect 453 -2158 808 -2157
rect 1269 -2158 1305 -2157
rect 86 -2160 227 -2159
rect 240 -2160 304 -2159
rect 485 -2160 528 -2159
rect 548 -2160 948 -2159
rect 1304 -2160 1326 -2159
rect 198 -2162 227 -2161
rect 240 -2162 360 -2161
rect 443 -2162 549 -2161
rect 590 -2162 717 -2161
rect 723 -2162 759 -2161
rect 772 -2162 920 -2161
rect 198 -2164 388 -2163
rect 436 -2164 444 -2163
rect 499 -2164 1179 -2163
rect 128 -2166 1179 -2165
rect 114 -2168 129 -2167
rect 219 -2168 528 -2167
rect 576 -2168 773 -2167
rect 807 -2168 1123 -2167
rect 296 -2170 332 -2169
rect 359 -2170 895 -2169
rect 324 -2172 388 -2171
rect 415 -2172 437 -2171
rect 499 -2172 811 -2171
rect 212 -2174 416 -2173
rect 502 -2174 780 -2173
rect 212 -2176 493 -2175
rect 520 -2176 640 -2175
rect 653 -2176 818 -2175
rect 324 -2178 402 -2177
rect 492 -2178 927 -2177
rect 401 -2180 1025 -2179
rect 523 -2182 941 -2181
rect 576 -2184 675 -2183
rect 716 -2184 752 -2183
rect 758 -2184 787 -2183
rect 597 -2186 619 -2185
rect 621 -2186 829 -2185
rect 506 -2188 619 -2187
rect 632 -2188 927 -2187
rect 93 -2190 507 -2189
rect 611 -2190 689 -2189
rect 751 -2190 801 -2189
rect 828 -2190 864 -2189
rect 93 -2192 283 -2191
rect 583 -2192 612 -2191
rect 786 -2192 1137 -2191
rect 117 -2194 633 -2193
rect 800 -2194 843 -2193
rect 863 -2194 913 -2193
rect 1136 -2194 1158 -2193
rect 282 -2196 514 -2195
rect 534 -2196 584 -2195
rect 842 -2196 878 -2195
rect 912 -2196 934 -2195
rect 1017 -2196 1158 -2195
rect 37 -2198 878 -2197
rect 933 -2198 1109 -2197
rect 380 -2200 514 -2199
rect 534 -2200 570 -2199
rect 1017 -2200 1060 -2199
rect 1108 -2200 1151 -2199
rect 135 -2202 381 -2201
rect 520 -2202 1060 -2201
rect 135 -2204 367 -2203
rect 569 -2204 626 -2203
rect 16 -2206 367 -2205
rect 562 -2206 626 -2205
rect 16 -2208 458 -2207
rect 562 -2208 605 -2207
rect 58 -2210 458 -2209
rect 604 -2210 647 -2209
rect 58 -2212 143 -2211
rect 152 -2212 1151 -2211
rect 100 -2214 647 -2213
rect 100 -2216 290 -2215
rect 121 -2218 143 -2217
rect 289 -2218 430 -2217
rect 23 -2220 430 -2219
rect 23 -2222 27 -2221
rect 121 -2222 409 -2221
rect 408 -2224 1067 -2223
rect 1066 -2226 1102 -2225
rect 1101 -2228 1144 -2227
rect 1143 -2230 1172 -2229
rect 1073 -2232 1172 -2231
rect 870 -2234 1074 -2233
rect 870 -2236 1053 -2235
rect 5 -2247 45 -2246
rect 61 -2247 493 -2246
rect 516 -2247 727 -2246
rect 747 -2247 1088 -2246
rect 23 -2249 1025 -2248
rect 1034 -2249 1291 -2248
rect 23 -2251 402 -2250
rect 408 -2251 416 -2250
rect 425 -2251 689 -2250
rect 761 -2251 857 -2250
rect 870 -2251 1235 -2250
rect 33 -2253 199 -2252
rect 205 -2253 339 -2252
rect 387 -2253 524 -2252
rect 527 -2253 738 -2252
rect 810 -2253 962 -2252
rect 982 -2253 1277 -2252
rect 9 -2255 199 -2254
rect 205 -2255 374 -2254
rect 387 -2255 423 -2254
rect 520 -2255 563 -2254
rect 579 -2255 969 -2254
rect 982 -2255 986 -2254
rect 1024 -2255 1095 -2254
rect 9 -2257 360 -2256
rect 411 -2257 465 -2256
rect 527 -2257 934 -2256
rect 961 -2257 1018 -2256
rect 1094 -2257 1151 -2256
rect 37 -2259 976 -2258
rect 1017 -2259 1081 -2258
rect 1150 -2259 1221 -2258
rect 37 -2261 342 -2260
rect 359 -2261 486 -2260
rect 530 -2261 927 -2260
rect 933 -2261 1060 -2260
rect 1080 -2261 1298 -2260
rect 40 -2263 353 -2262
rect 464 -2263 850 -2262
rect 856 -2263 1011 -2262
rect 1059 -2263 1123 -2262
rect 40 -2265 927 -2264
rect 975 -2265 1270 -2264
rect 44 -2267 381 -2266
rect 485 -2267 514 -2266
rect 548 -2267 689 -2266
rect 695 -2267 850 -2266
rect 870 -2267 941 -2266
rect 1122 -2267 1193 -2266
rect 79 -2269 416 -2268
rect 548 -2269 605 -2268
rect 625 -2269 640 -2268
rect 674 -2269 773 -2268
rect 873 -2269 1032 -2268
rect 1192 -2269 1242 -2268
rect 16 -2271 80 -2270
rect 86 -2271 297 -2270
rect 306 -2271 409 -2270
rect 492 -2271 1032 -2270
rect 1129 -2271 1242 -2270
rect 16 -2273 318 -2272
rect 320 -2273 1235 -2272
rect 86 -2275 724 -2274
rect 737 -2275 745 -2274
rect 772 -2275 801 -2274
rect 96 -2277 619 -2276
rect 628 -2277 969 -2276
rect 100 -2279 115 -2278
rect 117 -2279 1179 -2278
rect 100 -2281 346 -2280
rect 352 -2281 479 -2280
rect 513 -2281 1130 -2280
rect 1178 -2281 1256 -2280
rect 114 -2283 192 -2282
rect 240 -2283 521 -2282
rect 558 -2283 682 -2282
rect 695 -2283 794 -2282
rect 800 -2283 815 -2282
rect 121 -2285 745 -2284
rect 793 -2285 811 -2284
rect 814 -2285 878 -2284
rect 121 -2287 451 -2286
rect 555 -2287 682 -2286
rect 877 -2287 948 -2286
rect 149 -2289 920 -2288
rect 947 -2289 1046 -2288
rect 149 -2291 437 -2290
rect 450 -2291 584 -2290
rect 593 -2291 836 -2290
rect 919 -2291 990 -2290
rect 1045 -2291 1305 -2290
rect 152 -2293 808 -2292
rect 989 -2293 1067 -2292
rect 156 -2295 297 -2294
rect 331 -2295 941 -2294
rect 1066 -2295 1165 -2294
rect 2 -2297 332 -2296
rect 341 -2297 458 -2296
rect 562 -2297 661 -2296
rect 677 -2297 1137 -2296
rect 2 -2299 479 -2298
rect 569 -2299 584 -2298
rect 604 -2299 703 -2298
rect 786 -2299 836 -2298
rect 107 -2301 458 -2300
rect 471 -2301 570 -2300
rect 611 -2301 619 -2300
rect 635 -2301 759 -2300
rect 807 -2301 1004 -2300
rect 107 -2303 129 -2302
rect 156 -2303 185 -2302
rect 191 -2303 290 -2302
rect 380 -2303 577 -2302
rect 611 -2303 633 -2302
rect 639 -2303 710 -2302
rect 758 -2303 1172 -2302
rect 75 -2305 633 -2304
rect 646 -2305 1165 -2304
rect 128 -2307 395 -2306
rect 471 -2307 507 -2306
rect 576 -2307 1221 -2306
rect 51 -2309 395 -2308
rect 499 -2309 507 -2308
rect 597 -2309 647 -2308
rect 660 -2309 1284 -2308
rect 51 -2311 139 -2310
rect 163 -2311 290 -2310
rect 338 -2311 1172 -2310
rect 138 -2313 1088 -2312
rect 163 -2315 405 -2314
rect 499 -2315 535 -2314
rect 590 -2315 598 -2314
rect 702 -2315 752 -2314
rect 1003 -2315 1207 -2314
rect 177 -2317 346 -2316
rect 534 -2317 864 -2316
rect 1206 -2317 1249 -2316
rect 170 -2319 178 -2318
rect 184 -2319 234 -2318
rect 254 -2319 374 -2318
rect 590 -2319 1137 -2318
rect 1248 -2319 1312 -2318
rect 93 -2321 255 -2320
rect 261 -2321 402 -2320
rect 709 -2321 717 -2320
rect 751 -2321 843 -2320
rect 863 -2321 955 -2320
rect 65 -2323 94 -2322
rect 170 -2323 318 -2322
rect 397 -2323 843 -2322
rect 954 -2323 1109 -2322
rect 30 -2325 66 -2324
rect 219 -2325 241 -2324
rect 261 -2325 556 -2324
rect 716 -2325 766 -2324
rect 1108 -2325 1186 -2324
rect 30 -2327 426 -2326
rect 1185 -2327 1228 -2326
rect 135 -2329 766 -2328
rect 891 -2329 1228 -2328
rect 135 -2331 367 -2330
rect 397 -2331 731 -2330
rect 891 -2331 997 -2330
rect 219 -2333 325 -2332
rect 366 -2333 542 -2332
rect 730 -2333 822 -2332
rect 996 -2333 1074 -2332
rect 226 -2335 787 -2334
rect 821 -2335 885 -2334
rect 1073 -2335 1144 -2334
rect 142 -2337 227 -2336
rect 233 -2337 269 -2336
rect 282 -2337 664 -2336
rect 779 -2337 885 -2336
rect 1143 -2337 1200 -2336
rect 142 -2339 829 -2338
rect 268 -2341 311 -2340
rect 324 -2341 444 -2340
rect 541 -2341 654 -2340
rect 779 -2341 913 -2340
rect 275 -2343 311 -2342
rect 443 -2343 454 -2342
rect 621 -2343 1200 -2342
rect 275 -2345 430 -2344
rect 653 -2345 668 -2344
rect 828 -2345 899 -2344
rect 912 -2345 1053 -2344
rect 72 -2347 668 -2346
rect 898 -2347 906 -2346
rect 72 -2349 248 -2348
rect 282 -2349 300 -2348
rect 436 -2349 1053 -2348
rect 58 -2351 248 -2350
rect 905 -2351 1116 -2350
rect 58 -2353 1011 -2352
rect 1038 -2353 1116 -2352
rect 212 -2355 430 -2354
rect 1038 -2355 1102 -2354
rect 212 -2357 304 -2356
rect 1101 -2357 1158 -2356
rect 1157 -2359 1214 -2358
rect 1213 -2361 1263 -2360
rect 9 -2372 377 -2371
rect 394 -2372 1235 -2371
rect 23 -2374 342 -2373
rect 352 -2374 437 -2373
rect 446 -2374 780 -2373
rect 796 -2374 955 -2373
rect 1031 -2374 1074 -2373
rect 1104 -2374 1116 -2373
rect 30 -2376 202 -2375
rect 303 -2376 843 -2375
rect 849 -2376 920 -2375
rect 954 -2376 1046 -2375
rect 1073 -2376 1200 -2375
rect 37 -2378 297 -2377
rect 303 -2378 426 -2377
rect 464 -2378 759 -2377
rect 779 -2378 1011 -2377
rect 1034 -2378 1179 -2377
rect 40 -2380 941 -2379
rect 1010 -2380 1060 -2379
rect 54 -2382 255 -2381
rect 320 -2382 787 -2381
rect 807 -2382 1144 -2381
rect 61 -2384 570 -2383
rect 576 -2384 906 -2383
rect 908 -2384 1221 -2383
rect 72 -2386 514 -2385
rect 520 -2386 811 -2385
rect 842 -2386 1109 -2385
rect 72 -2388 171 -2387
rect 184 -2388 307 -2387
rect 338 -2388 444 -2387
rect 485 -2388 850 -2387
rect 898 -2388 1014 -2387
rect 1059 -2388 1081 -2387
rect 79 -2390 150 -2389
rect 163 -2390 297 -2389
rect 359 -2390 363 -2389
rect 366 -2390 517 -2389
rect 520 -2390 594 -2389
rect 614 -2390 864 -2389
rect 898 -2390 1158 -2389
rect 44 -2392 80 -2391
rect 86 -2392 367 -2391
rect 394 -2392 472 -2391
rect 516 -2392 1165 -2391
rect 86 -2394 283 -2393
rect 359 -2394 409 -2393
rect 422 -2394 689 -2393
rect 723 -2394 773 -2393
rect 786 -2394 853 -2393
rect 905 -2394 1242 -2393
rect 93 -2396 423 -2395
rect 450 -2396 864 -2395
rect 919 -2396 997 -2395
rect 1080 -2396 1137 -2395
rect 93 -2398 398 -2397
rect 450 -2398 871 -2397
rect 884 -2398 997 -2397
rect 100 -2400 745 -2399
rect 751 -2400 759 -2399
rect 765 -2400 808 -2399
rect 870 -2400 913 -2399
rect 940 -2400 1123 -2399
rect 100 -2402 143 -2401
rect 184 -2402 563 -2401
rect 569 -2402 626 -2401
rect 635 -2402 703 -2401
rect 709 -2402 885 -2401
rect 912 -2402 1172 -2401
rect 107 -2404 171 -2403
rect 198 -2404 440 -2403
rect 457 -2404 486 -2403
rect 548 -2404 577 -2403
rect 590 -2404 654 -2403
rect 660 -2404 1228 -2403
rect 107 -2406 598 -2405
rect 611 -2406 654 -2405
rect 663 -2406 1067 -2405
rect 58 -2408 598 -2407
rect 646 -2408 745 -2407
rect 751 -2408 892 -2407
rect 961 -2408 1109 -2407
rect 58 -2410 248 -2409
rect 261 -2410 591 -2409
rect 646 -2410 934 -2409
rect 1066 -2410 1130 -2409
rect 121 -2412 255 -2411
rect 261 -2412 507 -2411
rect 555 -2412 731 -2411
rect 765 -2412 976 -2411
rect 1129 -2412 1249 -2411
rect 124 -2414 969 -2413
rect 128 -2416 164 -2415
rect 198 -2416 227 -2415
rect 247 -2416 325 -2415
rect 362 -2416 409 -2415
rect 415 -2416 661 -2415
rect 667 -2416 703 -2415
rect 709 -2416 990 -2415
rect 128 -2418 139 -2417
rect 142 -2418 318 -2417
rect 387 -2418 626 -2417
rect 667 -2418 829 -2417
rect 877 -2418 934 -2417
rect 989 -2418 1193 -2417
rect 131 -2420 549 -2419
rect 558 -2420 640 -2419
rect 674 -2420 976 -2419
rect 1192 -2420 1207 -2419
rect 226 -2422 332 -2421
rect 380 -2422 675 -2421
rect 681 -2422 724 -2421
rect 726 -2422 962 -2421
rect 51 -2424 381 -2423
rect 387 -2424 430 -2423
rect 439 -2424 762 -2423
rect 772 -2424 857 -2423
rect 877 -2424 1018 -2423
rect 275 -2426 727 -2425
rect 814 -2426 892 -2425
rect 1017 -2426 1214 -2425
rect 212 -2428 276 -2427
rect 282 -2428 402 -2427
rect 415 -2428 465 -2427
rect 471 -2428 605 -2427
rect 611 -2428 969 -2427
rect 212 -2430 241 -2429
rect 289 -2430 325 -2429
rect 331 -2430 374 -2429
rect 401 -2430 514 -2429
rect 579 -2430 731 -2429
rect 814 -2430 1095 -2429
rect 177 -2432 241 -2431
rect 289 -2432 353 -2431
rect 373 -2432 829 -2431
rect 856 -2432 1039 -2431
rect 156 -2434 178 -2433
rect 317 -2434 346 -2433
rect 429 -2434 535 -2433
rect 604 -2434 1088 -2433
rect 156 -2436 234 -2435
rect 345 -2436 468 -2435
rect 478 -2436 563 -2435
rect 618 -2436 682 -2435
rect 688 -2436 927 -2435
rect 982 -2436 1088 -2435
rect 233 -2438 528 -2437
rect 534 -2438 633 -2437
rect 639 -2438 738 -2437
rect 926 -2438 1004 -2437
rect 457 -2440 493 -2439
rect 499 -2440 507 -2439
rect 527 -2440 696 -2439
rect 737 -2440 944 -2439
rect 982 -2440 1102 -2439
rect 478 -2442 584 -2441
rect 618 -2442 717 -2441
rect 821 -2442 1004 -2441
rect 1094 -2442 1102 -2441
rect 268 -2444 584 -2443
rect 632 -2444 801 -2443
rect 821 -2444 1053 -2443
rect 205 -2446 269 -2445
rect 492 -2446 794 -2445
rect 205 -2448 220 -2447
rect 499 -2448 573 -2447
rect 695 -2448 1151 -2447
rect 191 -2450 220 -2449
rect 541 -2450 801 -2449
rect 16 -2452 192 -2451
rect 443 -2452 542 -2451
rect 716 -2452 836 -2451
rect 835 -2454 1025 -2453
rect 947 -2456 1025 -2455
rect 947 -2458 1186 -2457
rect 58 -2469 461 -2468
rect 471 -2469 524 -2468
rect 530 -2469 584 -2468
rect 625 -2469 867 -2468
rect 961 -2469 1102 -2468
rect 1108 -2469 1144 -2468
rect 1185 -2469 1193 -2468
rect 65 -2471 353 -2470
rect 366 -2471 587 -2470
rect 625 -2471 822 -2470
rect 828 -2471 871 -2470
rect 1013 -2471 1130 -2470
rect 72 -2473 132 -2472
rect 149 -2473 353 -2472
rect 366 -2473 605 -2472
rect 639 -2473 643 -2472
rect 674 -2473 759 -2472
rect 793 -2473 808 -2472
rect 828 -2473 857 -2472
rect 863 -2473 871 -2472
rect 1024 -2473 1105 -2472
rect 79 -2475 472 -2474
rect 478 -2475 696 -2474
rect 723 -2475 948 -2474
rect 1038 -2475 1074 -2474
rect 1087 -2475 1179 -2474
rect 86 -2477 167 -2476
rect 191 -2477 692 -2476
rect 740 -2477 878 -2476
rect 926 -2477 948 -2476
rect 1052 -2477 1060 -2476
rect 107 -2479 468 -2478
rect 492 -2479 605 -2478
rect 618 -2479 724 -2478
rect 758 -2479 843 -2478
rect 863 -2479 983 -2478
rect 124 -2481 227 -2480
rect 247 -2481 493 -2480
rect 499 -2481 584 -2480
rect 639 -2481 787 -2480
rect 800 -2481 811 -2480
rect 926 -2481 997 -2480
rect 173 -2483 248 -2482
rect 278 -2483 360 -2482
rect 373 -2483 444 -2482
rect 446 -2483 850 -2482
rect 201 -2485 227 -2484
rect 282 -2485 479 -2484
rect 499 -2485 745 -2484
rect 772 -2485 794 -2484
rect 800 -2485 913 -2484
rect 212 -2487 552 -2486
rect 565 -2487 976 -2486
rect 219 -2489 356 -2488
rect 359 -2489 377 -2488
rect 380 -2489 685 -2488
rect 730 -2489 787 -2488
rect 807 -2489 990 -2488
rect 205 -2491 381 -2490
rect 390 -2491 514 -2490
rect 520 -2491 696 -2490
rect 730 -2491 752 -2490
rect 772 -2491 836 -2490
rect 912 -2491 955 -2490
rect 975 -2491 1004 -2490
rect 93 -2493 521 -2492
rect 544 -2493 573 -2492
rect 597 -2493 745 -2492
rect 954 -2493 1018 -2492
rect 114 -2495 573 -2494
rect 597 -2495 738 -2494
rect 1017 -2495 1032 -2494
rect 282 -2497 346 -2496
rect 373 -2497 535 -2496
rect 548 -2497 944 -2496
rect 1031 -2497 1067 -2496
rect 289 -2499 612 -2498
rect 646 -2499 752 -2498
rect 1066 -2499 1081 -2498
rect 233 -2501 290 -2500
rect 296 -2501 678 -2500
rect 170 -2503 234 -2502
rect 296 -2503 304 -2502
rect 317 -2503 440 -2502
rect 443 -2503 556 -2502
rect 569 -2503 780 -2502
rect 100 -2505 304 -2504
rect 327 -2505 402 -2504
rect 415 -2505 535 -2504
rect 541 -2505 612 -2504
rect 642 -2505 647 -2504
rect 653 -2505 738 -2504
rect 240 -2507 416 -2506
rect 422 -2507 619 -2506
rect 653 -2507 703 -2506
rect 275 -2509 318 -2508
rect 331 -2509 465 -2508
rect 509 -2509 969 -2508
rect 128 -2511 332 -2510
rect 345 -2511 486 -2510
rect 513 -2511 710 -2510
rect 121 -2513 129 -2512
rect 310 -2513 402 -2512
rect 429 -2513 661 -2512
rect 667 -2513 675 -2512
rect 702 -2513 717 -2512
rect 184 -2515 311 -2514
rect 408 -2515 430 -2514
rect 436 -2515 906 -2514
rect 268 -2517 409 -2516
rect 450 -2517 475 -2516
rect 485 -2517 815 -2516
rect 142 -2519 269 -2518
rect 387 -2519 437 -2518
rect 527 -2519 710 -2518
rect 177 -2521 451 -2520
rect 548 -2521 920 -2520
rect 387 -2523 395 -2522
rect 555 -2523 689 -2522
rect 324 -2525 395 -2524
rect 569 -2525 682 -2524
rect 576 -2527 668 -2526
rect 681 -2527 934 -2526
rect 457 -2529 577 -2528
rect 590 -2529 780 -2528
rect 884 -2529 934 -2528
rect 422 -2531 458 -2530
rect 590 -2531 892 -2530
rect 632 -2533 717 -2532
rect 562 -2535 633 -2534
rect 660 -2535 766 -2534
rect 506 -2537 563 -2536
rect 765 -2537 899 -2536
rect 261 -2539 507 -2538
rect 156 -2541 262 -2540
rect 131 -2552 136 -2551
rect 226 -2552 258 -2551
rect 261 -2552 367 -2551
rect 380 -2552 528 -2551
rect 530 -2552 703 -2551
rect 716 -2552 808 -2551
rect 814 -2552 829 -2551
rect 866 -2552 927 -2551
rect 933 -2552 965 -2551
rect 968 -2552 976 -2551
rect 1013 -2552 1039 -2551
rect 1045 -2552 1053 -2551
rect 1059 -2552 1067 -2551
rect 1143 -2552 1179 -2551
rect 1181 -2552 1186 -2551
rect 128 -2554 136 -2553
rect 233 -2554 276 -2553
rect 282 -2554 388 -2553
rect 394 -2554 472 -2553
rect 478 -2554 678 -2553
rect 681 -2554 773 -2553
rect 870 -2554 888 -2553
rect 898 -2554 913 -2553
rect 1024 -2554 1032 -2553
rect 247 -2556 325 -2555
rect 331 -2556 486 -2555
rect 492 -2556 685 -2555
rect 688 -2556 731 -2555
rect 744 -2556 794 -2555
rect 884 -2556 955 -2555
rect 268 -2558 325 -2557
rect 345 -2558 367 -2557
rect 401 -2558 549 -2557
rect 551 -2558 654 -2557
rect 663 -2558 668 -2557
rect 681 -2558 780 -2557
rect 947 -2558 955 -2557
rect 289 -2560 384 -2559
rect 415 -2560 493 -2559
rect 506 -2560 612 -2559
rect 621 -2560 801 -2559
rect 303 -2562 594 -2561
rect 600 -2562 647 -2561
rect 660 -2562 668 -2561
rect 716 -2562 759 -2561
rect 310 -2564 650 -2563
rect 723 -2564 811 -2563
rect 317 -2566 332 -2565
rect 359 -2566 507 -2565
rect 523 -2566 542 -2565
rect 565 -2566 640 -2565
rect 723 -2566 766 -2565
rect 429 -2568 489 -2567
rect 527 -2568 556 -2567
rect 569 -2568 675 -2567
rect 730 -2568 752 -2567
rect 436 -2570 545 -2569
rect 576 -2570 591 -2569
rect 632 -2570 713 -2569
rect 747 -2570 787 -2569
rect 443 -2572 461 -2571
rect 513 -2572 556 -2571
rect 576 -2572 598 -2571
rect 695 -2572 752 -2571
rect 338 -2574 514 -2573
rect 530 -2574 563 -2573
rect 296 -2576 339 -2575
rect 373 -2576 444 -2575
rect 450 -2576 570 -2575
rect 352 -2578 451 -2577
rect 464 -2578 598 -2577
rect 373 -2580 423 -2579
rect 534 -2580 647 -2579
rect 408 -2582 535 -2581
rect 541 -2582 710 -2581
rect 562 -2584 626 -2583
rect 604 -2586 710 -2585
rect 131 -2597 136 -2596
rect 324 -2597 384 -2596
rect 443 -2597 517 -2596
rect 534 -2597 664 -2596
rect 674 -2597 724 -2596
rect 751 -2597 808 -2596
rect 810 -2597 815 -2596
rect 884 -2597 899 -2596
rect 954 -2597 965 -2596
rect 1010 -2597 1018 -2596
rect 1045 -2597 1053 -2596
rect 1055 -2597 1060 -2596
rect 331 -2599 349 -2598
rect 366 -2599 381 -2598
rect 450 -2599 545 -2598
rect 548 -2599 577 -2598
rect 660 -2599 668 -2598
rect 684 -2599 717 -2598
rect 961 -2599 969 -2598
rect 1013 -2599 1025 -2598
rect 338 -2601 374 -2600
rect 471 -2601 552 -2600
rect 555 -2601 601 -2600
rect 709 -2601 731 -2600
rect 492 -2603 566 -2602
rect 569 -2603 682 -2602
rect 499 -2605 514 -2604
rect 506 -2607 650 -2606
<< m2contact >>
rect 215 0 216 1
rect 240 0 241 1
rect 247 0 248 1
rect 478 0 479 1
rect 562 0 563 1
rect 639 0 640 1
rect 667 0 668 1
rect 702 0 703 1
rect 800 0 801 1
rect 828 0 829 1
rect 261 -2 262 -1
rect 268 -2 269 -1
rect 275 -2 276 -1
rect 408 -2 409 -1
rect 411 -2 412 -1
rect 506 -2 507 -1
rect 576 -2 577 -1
rect 607 -2 608 -1
rect 681 -2 682 -1
rect 803 -2 804 -1
rect 338 -4 339 -3
rect 380 -4 381 -3
rect 387 -4 388 -3
rect 583 -4 584 -3
rect 586 -4 587 -3
rect 709 -4 710 -3
rect 373 -6 374 -5
rect 401 -6 402 -5
rect 415 -6 416 -5
rect 457 -6 458 -5
rect 464 -6 465 -5
rect 527 -6 528 -5
rect 604 -6 605 -5
rect 765 -6 766 -5
rect 397 -8 398 -7
rect 485 -8 486 -7
rect 425 -10 426 -9
rect 569 -10 570 -9
rect 429 -12 430 -11
rect 516 -12 517 -11
rect 467 -14 468 -13
rect 499 -14 500 -13
rect 163 -25 164 -24
rect 285 -25 286 -24
rect 292 -25 293 -24
rect 338 -25 339 -24
rect 359 -25 360 -24
rect 467 -25 468 -24
rect 478 -25 479 -24
rect 604 -25 605 -24
rect 621 -25 622 -24
rect 723 -25 724 -24
rect 800 -25 801 -24
rect 905 -25 906 -24
rect 191 -27 192 -26
rect 247 -27 248 -26
rect 254 -27 255 -26
rect 401 -27 402 -26
rect 404 -27 405 -26
rect 443 -27 444 -26
rect 464 -27 465 -26
rect 607 -27 608 -26
rect 639 -27 640 -26
rect 688 -27 689 -26
rect 702 -27 703 -26
rect 751 -27 752 -26
rect 828 -27 829 -26
rect 849 -27 850 -26
rect 215 -29 216 -28
rect 219 -29 220 -28
rect 226 -29 227 -28
rect 275 -29 276 -28
rect 282 -29 283 -28
rect 394 -29 395 -28
rect 401 -29 402 -28
rect 411 -29 412 -28
rect 436 -29 437 -28
rect 460 -29 461 -28
rect 481 -29 482 -28
rect 660 -29 661 -28
rect 667 -29 668 -28
rect 674 -29 675 -28
rect 709 -29 710 -28
rect 758 -29 759 -28
rect 765 -29 766 -28
rect 828 -29 829 -28
rect 233 -31 234 -30
rect 240 -31 241 -30
rect 247 -31 248 -30
rect 261 -31 262 -30
rect 268 -31 269 -30
rect 383 -31 384 -30
rect 408 -31 409 -30
rect 471 -31 472 -30
rect 485 -31 486 -30
rect 520 -31 521 -30
rect 527 -31 528 -30
rect 541 -31 542 -30
rect 551 -31 552 -30
rect 597 -31 598 -30
rect 639 -31 640 -30
rect 681 -31 682 -30
rect 719 -31 720 -30
rect 877 -31 878 -30
rect 261 -33 262 -32
rect 387 -33 388 -32
rect 492 -33 493 -32
rect 548 -33 549 -32
rect 555 -33 556 -32
rect 681 -33 682 -32
rect 275 -35 276 -34
rect 355 -35 356 -34
rect 366 -35 367 -34
rect 513 -35 514 -34
rect 516 -35 517 -34
rect 632 -35 633 -34
rect 653 -35 654 -34
rect 716 -35 717 -34
rect 282 -37 283 -36
rect 425 -37 426 -36
rect 499 -37 500 -36
rect 513 -37 514 -36
rect 534 -37 535 -36
rect 702 -37 703 -36
rect 296 -39 297 -38
rect 429 -39 430 -38
rect 502 -39 503 -38
rect 527 -39 528 -38
rect 548 -39 549 -38
rect 618 -39 619 -38
rect 303 -41 304 -40
rect 397 -41 398 -40
rect 429 -41 430 -40
rect 537 -41 538 -40
rect 569 -41 570 -40
rect 625 -41 626 -40
rect 310 -43 311 -42
rect 422 -43 423 -42
rect 457 -43 458 -42
rect 569 -43 570 -42
rect 576 -43 577 -42
rect 611 -43 612 -42
rect 317 -45 318 -44
rect 579 -45 580 -44
rect 583 -45 584 -44
rect 646 -45 647 -44
rect 324 -47 325 -46
rect 373 -47 374 -46
rect 380 -47 381 -46
rect 485 -47 486 -46
rect 506 -47 507 -46
rect 583 -47 584 -46
rect 593 -47 594 -46
rect 772 -47 773 -46
rect 331 -49 332 -48
rect 418 -49 419 -48
rect 457 -49 458 -48
rect 478 -49 479 -48
rect 506 -49 507 -48
rect 562 -49 563 -48
rect 345 -51 346 -50
rect 667 -51 668 -50
rect 373 -53 374 -52
rect 415 -53 416 -52
rect 380 -55 381 -54
rect 562 -55 563 -54
rect 387 -57 388 -56
rect 499 -57 500 -56
rect 23 -68 24 -67
rect 355 -68 356 -67
rect 415 -68 416 -67
rect 548 -68 549 -67
rect 562 -68 563 -67
rect 709 -68 710 -67
rect 723 -68 724 -67
rect 779 -68 780 -67
rect 828 -68 829 -67
rect 870 -68 871 -67
rect 877 -68 878 -67
rect 940 -68 941 -67
rect 1500 -68 1501 -67
rect 1507 -68 1508 -67
rect 30 -70 31 -69
rect 152 -70 153 -69
rect 156 -70 157 -69
rect 292 -70 293 -69
rect 313 -70 314 -69
rect 397 -70 398 -69
rect 422 -70 423 -69
rect 548 -70 549 -69
rect 562 -70 563 -69
rect 639 -70 640 -69
rect 663 -70 664 -69
rect 856 -70 857 -69
rect 905 -70 906 -69
rect 947 -70 948 -69
rect 37 -72 38 -71
rect 331 -72 332 -71
rect 373 -72 374 -71
rect 415 -72 416 -71
rect 478 -72 479 -71
rect 695 -72 696 -71
rect 702 -72 703 -71
rect 800 -72 801 -71
rect 849 -72 850 -71
rect 877 -72 878 -71
rect 44 -74 45 -73
rect 159 -74 160 -73
rect 170 -74 171 -73
rect 310 -74 311 -73
rect 324 -74 325 -73
rect 380 -74 381 -73
rect 394 -74 395 -73
rect 478 -74 479 -73
rect 481 -74 482 -73
rect 485 -74 486 -73
rect 499 -74 500 -73
rect 534 -74 535 -73
rect 541 -74 542 -73
rect 579 -74 580 -73
rect 604 -74 605 -73
rect 723 -74 724 -73
rect 751 -74 752 -73
rect 814 -74 815 -73
rect 51 -76 52 -75
rect 366 -76 367 -75
rect 373 -76 374 -75
rect 429 -76 430 -75
rect 471 -76 472 -75
rect 541 -76 542 -75
rect 576 -76 577 -75
rect 821 -76 822 -75
rect 75 -78 76 -77
rect 100 -78 101 -77
rect 107 -78 108 -77
rect 117 -78 118 -77
rect 121 -78 122 -77
rect 450 -78 451 -77
rect 471 -78 472 -77
rect 555 -78 556 -77
rect 576 -78 577 -77
rect 593 -78 594 -77
rect 604 -78 605 -77
rect 751 -78 752 -77
rect 758 -78 759 -77
rect 786 -78 787 -77
rect 79 -80 80 -79
rect 383 -80 384 -79
rect 429 -80 430 -79
rect 457 -80 458 -79
rect 485 -80 486 -79
rect 611 -80 612 -79
rect 618 -80 619 -79
rect 716 -80 717 -79
rect 772 -80 773 -79
rect 849 -80 850 -79
rect 86 -82 87 -81
rect 89 -82 90 -81
rect 93 -82 94 -81
rect 275 -82 276 -81
rect 296 -82 297 -81
rect 422 -82 423 -81
rect 436 -82 437 -81
rect 457 -82 458 -81
rect 499 -82 500 -81
rect 558 -82 559 -81
rect 618 -82 619 -81
rect 674 -82 675 -81
rect 681 -82 682 -81
rect 730 -82 731 -81
rect 114 -84 115 -83
rect 275 -84 276 -83
rect 299 -84 300 -83
rect 436 -84 437 -83
rect 450 -84 451 -83
rect 597 -84 598 -83
rect 632 -84 633 -83
rect 681 -84 682 -83
rect 688 -84 689 -83
rect 744 -84 745 -83
rect 128 -86 129 -85
rect 212 -86 213 -85
rect 219 -86 220 -85
rect 331 -86 332 -85
rect 352 -86 353 -85
rect 555 -86 556 -85
rect 625 -86 626 -85
rect 632 -86 633 -85
rect 646 -86 647 -85
rect 772 -86 773 -85
rect 135 -88 136 -87
rect 317 -88 318 -87
rect 352 -88 353 -87
rect 359 -88 360 -87
rect 366 -88 367 -87
rect 387 -88 388 -87
rect 404 -88 405 -87
rect 646 -88 647 -87
rect 660 -88 661 -87
rect 674 -88 675 -87
rect 142 -90 143 -89
rect 163 -90 164 -89
rect 177 -90 178 -89
rect 341 -90 342 -89
rect 359 -90 360 -89
rect 702 -90 703 -89
rect 163 -92 164 -91
rect 327 -92 328 -91
rect 338 -92 339 -91
rect 387 -92 388 -91
rect 453 -92 454 -91
rect 688 -92 689 -91
rect 184 -94 185 -93
rect 282 -94 283 -93
rect 338 -94 339 -93
rect 394 -94 395 -93
rect 506 -94 507 -93
rect 611 -94 612 -93
rect 625 -94 626 -93
rect 653 -94 654 -93
rect 660 -94 661 -93
rect 737 -94 738 -93
rect 187 -96 188 -95
rect 226 -96 227 -95
rect 254 -96 255 -95
rect 317 -96 318 -95
rect 464 -96 465 -95
rect 506 -96 507 -95
rect 513 -96 514 -95
rect 597 -96 598 -95
rect 667 -96 668 -95
rect 719 -96 720 -95
rect 149 -98 150 -97
rect 226 -98 227 -97
rect 254 -98 255 -97
rect 261 -98 262 -97
rect 268 -98 269 -97
rect 408 -98 409 -97
rect 411 -98 412 -97
rect 513 -98 514 -97
rect 520 -98 521 -97
rect 639 -98 640 -97
rect 670 -98 671 -97
rect 807 -98 808 -97
rect 149 -100 150 -99
rect 194 -100 195 -99
rect 198 -100 199 -99
rect 233 -100 234 -99
rect 247 -100 248 -99
rect 268 -100 269 -99
rect 271 -100 272 -99
rect 310 -100 311 -99
rect 520 -100 521 -99
rect 607 -100 608 -99
rect 191 -102 192 -101
rect 240 -102 241 -101
rect 247 -102 248 -101
rect 418 -102 419 -101
rect 527 -102 528 -101
rect 765 -102 766 -101
rect 205 -104 206 -103
rect 348 -104 349 -103
rect 530 -104 531 -103
rect 793 -104 794 -103
rect 219 -106 220 -105
rect 345 -106 346 -105
rect 569 -106 570 -105
rect 653 -106 654 -105
rect 233 -108 234 -107
rect 289 -108 290 -107
rect 345 -108 346 -107
rect 590 -108 591 -107
rect 65 -110 66 -109
rect 289 -110 290 -109
rect 443 -110 444 -109
rect 569 -110 570 -109
rect 261 -112 262 -111
rect 401 -112 402 -111
rect 439 -112 440 -111
rect 443 -112 444 -111
rect 492 -112 493 -111
rect 590 -112 591 -111
rect 282 -114 283 -113
rect 537 -114 538 -113
rect 401 -116 402 -115
rect 464 -116 465 -115
rect 492 -116 493 -115
rect 583 -116 584 -115
rect 583 -118 584 -117
rect 761 -118 762 -117
rect 16 -129 17 -128
rect 439 -129 440 -128
rect 488 -129 489 -128
rect 765 -129 766 -128
rect 793 -129 794 -128
rect 828 -129 829 -128
rect 849 -129 850 -128
rect 884 -129 885 -128
rect 940 -129 941 -128
rect 968 -129 969 -128
rect 975 -129 976 -128
rect 1024 -129 1025 -128
rect 9 -131 10 -130
rect 439 -131 440 -130
rect 516 -131 517 -130
rect 597 -131 598 -130
rect 604 -131 605 -130
rect 772 -131 773 -130
rect 800 -131 801 -130
rect 912 -131 913 -130
rect 947 -131 948 -130
rect 978 -131 979 -130
rect 30 -133 31 -132
rect 54 -133 55 -132
rect 58 -133 59 -132
rect 65 -133 66 -132
rect 72 -133 73 -132
rect 75 -133 76 -132
rect 86 -133 87 -132
rect 366 -133 367 -132
rect 394 -133 395 -132
rect 985 -133 986 -132
rect 30 -135 31 -134
rect 61 -135 62 -134
rect 107 -135 108 -134
rect 114 -135 115 -134
rect 117 -135 118 -134
rect 390 -135 391 -134
rect 537 -135 538 -134
rect 835 -135 836 -134
rect 849 -135 850 -134
rect 982 -135 983 -134
rect 44 -137 45 -136
rect 271 -137 272 -136
rect 275 -137 276 -136
rect 359 -137 360 -136
rect 541 -137 542 -136
rect 597 -137 598 -136
rect 607 -137 608 -136
rect 919 -137 920 -136
rect 51 -139 52 -138
rect 401 -139 402 -138
rect 464 -139 465 -138
rect 607 -139 608 -138
rect 611 -139 612 -138
rect 842 -139 843 -138
rect 856 -139 857 -138
rect 961 -139 962 -138
rect 51 -141 52 -140
rect 142 -141 143 -140
rect 145 -141 146 -140
rect 299 -141 300 -140
rect 310 -141 311 -140
rect 401 -141 402 -140
rect 443 -141 444 -140
rect 464 -141 465 -140
rect 478 -141 479 -140
rect 611 -141 612 -140
rect 646 -141 647 -140
rect 793 -141 794 -140
rect 807 -141 808 -140
rect 891 -141 892 -140
rect 58 -143 59 -142
rect 79 -143 80 -142
rect 93 -143 94 -142
rect 275 -143 276 -142
rect 289 -143 290 -142
rect 527 -143 528 -142
rect 555 -143 556 -142
rect 996 -143 997 -142
rect 79 -145 80 -144
rect 163 -145 164 -144
rect 226 -145 227 -144
rect 296 -145 297 -144
rect 327 -145 328 -144
rect 352 -145 353 -144
rect 422 -145 423 -144
rect 478 -145 479 -144
rect 513 -145 514 -144
rect 541 -145 542 -144
rect 562 -145 563 -144
rect 772 -145 773 -144
rect 779 -145 780 -144
rect 856 -145 857 -144
rect 870 -145 871 -144
rect 926 -145 927 -144
rect 121 -147 122 -146
rect 184 -147 185 -146
rect 226 -147 227 -146
rect 362 -147 363 -146
rect 422 -147 423 -146
rect 499 -147 500 -146
rect 520 -147 521 -146
rect 527 -147 528 -146
rect 646 -147 647 -146
rect 681 -147 682 -146
rect 688 -147 689 -146
rect 758 -147 759 -146
rect 779 -147 780 -146
rect 814 -147 815 -146
rect 821 -147 822 -146
rect 954 -147 955 -146
rect 89 -149 90 -148
rect 520 -149 521 -148
rect 639 -149 640 -148
rect 821 -149 822 -148
rect 877 -149 878 -148
rect 947 -149 948 -148
rect 100 -151 101 -150
rect 121 -151 122 -150
rect 131 -151 132 -150
rect 310 -151 311 -150
rect 324 -151 325 -150
rect 352 -151 353 -150
rect 429 -151 430 -150
rect 555 -151 556 -150
rect 583 -151 584 -150
rect 639 -151 640 -150
rect 653 -151 654 -150
rect 877 -151 878 -150
rect 68 -153 69 -152
rect 100 -153 101 -152
rect 135 -153 136 -152
rect 296 -153 297 -152
rect 443 -153 444 -152
rect 709 -153 710 -152
rect 716 -153 717 -152
rect 905 -153 906 -152
rect 135 -155 136 -154
rect 170 -155 171 -154
rect 233 -155 234 -154
rect 366 -155 367 -154
rect 485 -155 486 -154
rect 583 -155 584 -154
rect 590 -155 591 -154
rect 709 -155 710 -154
rect 719 -155 720 -154
rect 800 -155 801 -154
rect 807 -155 808 -154
rect 989 -155 990 -154
rect 142 -157 143 -156
rect 191 -157 192 -156
rect 194 -157 195 -156
rect 233 -157 234 -156
rect 247 -157 248 -156
rect 324 -157 325 -156
rect 415 -157 416 -156
rect 590 -157 591 -156
rect 625 -157 626 -156
rect 653 -157 654 -156
rect 660 -157 661 -156
rect 786 -157 787 -156
rect 149 -159 150 -158
rect 187 -159 188 -158
rect 247 -159 248 -158
rect 397 -159 398 -158
rect 415 -159 416 -158
rect 471 -159 472 -158
rect 485 -159 486 -158
rect 562 -159 563 -158
rect 576 -159 577 -158
rect 625 -159 626 -158
rect 667 -159 668 -158
rect 814 -159 815 -158
rect 44 -161 45 -160
rect 149 -161 150 -160
rect 152 -161 153 -160
rect 191 -161 192 -160
rect 254 -161 255 -160
rect 320 -161 321 -160
rect 387 -161 388 -160
rect 471 -161 472 -160
rect 492 -161 493 -160
rect 576 -161 577 -160
rect 663 -161 664 -160
rect 667 -161 668 -160
rect 674 -161 675 -160
rect 765 -161 766 -160
rect 163 -163 164 -162
rect 177 -163 178 -162
rect 219 -163 220 -162
rect 254 -163 255 -162
rect 271 -163 272 -162
rect 317 -163 318 -162
rect 373 -163 374 -162
rect 387 -163 388 -162
rect 457 -163 458 -162
rect 492 -163 493 -162
rect 569 -163 570 -162
rect 674 -163 675 -162
rect 688 -163 689 -162
rect 695 -163 696 -162
rect 702 -163 703 -162
rect 898 -163 899 -162
rect 170 -165 171 -164
rect 205 -165 206 -164
rect 219 -165 220 -164
rect 306 -165 307 -164
rect 317 -165 318 -164
rect 681 -165 682 -164
rect 723 -165 724 -164
rect 933 -165 934 -164
rect 177 -167 178 -166
rect 212 -167 213 -166
rect 268 -167 269 -166
rect 702 -167 703 -166
rect 730 -167 731 -166
rect 786 -167 787 -166
rect 107 -169 108 -168
rect 268 -169 269 -168
rect 282 -169 283 -168
rect 289 -169 290 -168
rect 303 -169 304 -168
rect 373 -169 374 -168
rect 457 -169 458 -168
rect 695 -169 696 -168
rect 737 -169 738 -168
rect 870 -169 871 -168
rect 198 -171 199 -170
rect 205 -171 206 -170
rect 240 -171 241 -170
rect 282 -171 283 -170
rect 303 -171 304 -170
rect 429 -171 430 -170
rect 530 -171 531 -170
rect 737 -171 738 -170
rect 744 -171 745 -170
rect 863 -171 864 -170
rect 128 -173 129 -172
rect 240 -173 241 -172
rect 331 -173 332 -172
rect 569 -173 570 -172
rect 618 -173 619 -172
rect 723 -173 724 -172
rect 751 -173 752 -172
rect 940 -173 941 -172
rect 93 -175 94 -174
rect 331 -175 332 -174
rect 334 -175 335 -174
rect 730 -175 731 -174
rect 156 -177 157 -176
rect 198 -177 199 -176
rect 436 -177 437 -176
rect 744 -177 745 -176
rect 156 -179 157 -178
rect 212 -179 213 -178
rect 436 -179 437 -178
rect 499 -179 500 -178
rect 534 -179 535 -178
rect 618 -179 619 -178
rect 450 -181 451 -180
rect 534 -181 535 -180
rect 548 -181 549 -180
rect 751 -181 752 -180
rect 408 -183 409 -182
rect 450 -183 451 -182
rect 506 -183 507 -182
rect 548 -183 549 -182
rect 103 -185 104 -184
rect 506 -185 507 -184
rect 380 -187 381 -186
rect 408 -187 409 -186
rect 338 -189 339 -188
rect 380 -189 381 -188
rect 338 -191 339 -190
rect 345 -191 346 -190
rect 37 -193 38 -192
rect 345 -193 346 -192
rect 37 -195 38 -194
rect 261 -195 262 -194
rect 261 -197 262 -196
rect 460 -197 461 -196
rect 2 -208 3 -207
rect 30 -208 31 -207
rect 37 -208 38 -207
rect 387 -208 388 -207
rect 436 -208 437 -207
rect 590 -208 591 -207
rect 604 -208 605 -207
rect 1080 -208 1081 -207
rect 1150 -208 1151 -207
rect 1178 -208 1179 -207
rect 37 -210 38 -209
rect 387 -210 388 -209
rect 394 -210 395 -209
rect 436 -210 437 -209
rect 439 -210 440 -209
rect 842 -210 843 -209
rect 849 -210 850 -209
rect 1059 -210 1060 -209
rect 44 -212 45 -211
rect 285 -212 286 -211
rect 303 -212 304 -211
rect 313 -212 314 -211
rect 446 -212 447 -211
rect 793 -212 794 -211
rect 835 -212 836 -211
rect 1087 -212 1088 -211
rect 44 -214 45 -213
rect 65 -214 66 -213
rect 72 -214 73 -213
rect 82 -214 83 -213
rect 103 -214 104 -213
rect 240 -214 241 -213
rect 243 -214 244 -213
rect 537 -214 538 -213
rect 544 -214 545 -213
rect 821 -214 822 -213
rect 863 -214 864 -213
rect 1108 -214 1109 -213
rect 51 -216 52 -215
rect 989 -216 990 -215
rect 1024 -216 1025 -215
rect 1045 -216 1046 -215
rect 51 -218 52 -217
rect 100 -218 101 -217
rect 107 -218 108 -217
rect 303 -218 304 -217
rect 310 -218 311 -217
rect 394 -218 395 -217
rect 453 -218 454 -217
rect 877 -218 878 -217
rect 891 -218 892 -217
rect 1017 -218 1018 -217
rect 65 -220 66 -219
rect 72 -220 73 -219
rect 107 -220 108 -219
rect 443 -220 444 -219
rect 485 -220 486 -219
rect 814 -220 815 -219
rect 821 -220 822 -219
rect 828 -220 829 -219
rect 870 -220 871 -219
rect 1101 -220 1102 -219
rect 96 -222 97 -221
rect 870 -222 871 -221
rect 912 -222 913 -221
rect 1122 -222 1123 -221
rect 205 -224 206 -223
rect 271 -224 272 -223
rect 282 -224 283 -223
rect 1066 -224 1067 -223
rect 159 -226 160 -225
rect 282 -226 283 -225
rect 310 -226 311 -225
rect 331 -226 332 -225
rect 362 -226 363 -225
rect 835 -226 836 -225
rect 926 -226 927 -225
rect 1052 -226 1053 -225
rect 198 -228 199 -227
rect 205 -228 206 -227
rect 233 -228 234 -227
rect 320 -228 321 -227
rect 415 -228 416 -227
rect 443 -228 444 -227
rect 457 -228 458 -227
rect 912 -228 913 -227
rect 947 -228 948 -227
rect 1129 -228 1130 -227
rect 177 -230 178 -229
rect 198 -230 199 -229
rect 233 -230 234 -229
rect 334 -230 335 -229
rect 408 -230 409 -229
rect 415 -230 416 -229
rect 425 -230 426 -229
rect 828 -230 829 -229
rect 947 -230 948 -229
rect 975 -230 976 -229
rect 54 -232 55 -231
rect 975 -232 976 -231
rect 177 -234 178 -233
rect 317 -234 318 -233
rect 320 -234 321 -233
rect 1136 -234 1137 -233
rect 240 -236 241 -235
rect 317 -236 318 -235
rect 429 -236 430 -235
rect 457 -236 458 -235
rect 506 -236 507 -235
rect 590 -236 591 -235
rect 607 -236 608 -235
rect 1073 -236 1074 -235
rect 124 -238 125 -237
rect 429 -238 430 -237
rect 513 -238 514 -237
rect 1115 -238 1116 -237
rect 268 -240 269 -239
rect 555 -240 556 -239
rect 579 -240 580 -239
rect 1143 -240 1144 -239
rect 128 -242 129 -241
rect 268 -242 269 -241
rect 373 -242 374 -241
rect 506 -242 507 -241
rect 513 -242 514 -241
rect 548 -242 549 -241
rect 607 -242 608 -241
rect 940 -242 941 -241
rect 954 -242 955 -241
rect 1094 -242 1095 -241
rect 26 -244 27 -243
rect 954 -244 955 -243
rect 961 -244 962 -243
rect 1010 -244 1011 -243
rect 128 -246 129 -245
rect 212 -246 213 -245
rect 219 -246 220 -245
rect 373 -246 374 -245
rect 408 -246 409 -245
rect 555 -246 556 -245
rect 639 -246 640 -245
rect 877 -246 878 -245
rect 919 -246 920 -245
rect 961 -246 962 -245
rect 968 -246 969 -245
rect 982 -246 983 -245
rect 170 -248 171 -247
rect 212 -248 213 -247
rect 219 -248 220 -247
rect 226 -248 227 -247
rect 401 -248 402 -247
rect 639 -248 640 -247
rect 674 -248 675 -247
rect 793 -248 794 -247
rect 800 -248 801 -247
rect 968 -248 969 -247
rect 978 -248 979 -247
rect 982 -248 983 -247
rect 40 -250 41 -249
rect 170 -250 171 -249
rect 345 -250 346 -249
rect 401 -250 402 -249
rect 492 -250 493 -249
rect 548 -250 549 -249
rect 576 -250 577 -249
rect 674 -250 675 -249
rect 688 -250 689 -249
rect 716 -250 717 -249
rect 719 -250 720 -249
rect 1003 -250 1004 -249
rect 86 -252 87 -251
rect 492 -252 493 -251
rect 516 -252 517 -251
rect 992 -252 993 -251
rect 58 -254 59 -253
rect 86 -254 87 -253
rect 163 -254 164 -253
rect 226 -254 227 -253
rect 327 -254 328 -253
rect 688 -254 689 -253
rect 695 -254 696 -253
rect 814 -254 815 -253
rect 58 -256 59 -255
rect 289 -256 290 -255
rect 345 -256 346 -255
rect 366 -256 367 -255
rect 534 -256 535 -255
rect 933 -256 934 -255
rect 23 -258 24 -257
rect 289 -258 290 -257
rect 359 -258 360 -257
rect 366 -258 367 -257
rect 534 -258 535 -257
rect 1153 -258 1154 -257
rect 163 -260 164 -259
rect 422 -260 423 -259
rect 576 -260 577 -259
rect 905 -260 906 -259
rect 191 -262 192 -261
rect 359 -262 360 -261
rect 618 -262 619 -261
rect 716 -262 717 -261
rect 737 -262 738 -261
rect 919 -262 920 -261
rect 33 -264 34 -263
rect 191 -264 192 -263
rect 562 -264 563 -263
rect 618 -264 619 -263
rect 625 -264 626 -263
rect 737 -264 738 -263
rect 744 -264 745 -263
rect 940 -264 941 -263
rect 541 -266 542 -265
rect 562 -266 563 -265
rect 583 -266 584 -265
rect 744 -266 745 -265
rect 758 -266 759 -265
rect 1024 -266 1025 -265
rect 380 -268 381 -267
rect 583 -268 584 -267
rect 611 -268 612 -267
rect 625 -268 626 -267
rect 667 -268 668 -267
rect 800 -268 801 -267
rect 884 -268 885 -267
rect 933 -268 934 -267
rect 121 -270 122 -269
rect 380 -270 381 -269
rect 527 -270 528 -269
rect 611 -270 612 -269
rect 698 -270 699 -269
rect 842 -270 843 -269
rect 121 -272 122 -271
rect 485 -272 486 -271
rect 499 -272 500 -271
rect 527 -272 528 -271
rect 541 -272 542 -271
rect 1031 -272 1032 -271
rect 142 -274 143 -273
rect 884 -274 885 -273
rect 114 -276 115 -275
rect 142 -276 143 -275
rect 296 -276 297 -275
rect 499 -276 500 -275
rect 702 -276 703 -275
rect 926 -276 927 -275
rect 114 -278 115 -277
rect 135 -278 136 -277
rect 296 -278 297 -277
rect 604 -278 605 -277
rect 705 -278 706 -277
rect 898 -278 899 -277
rect 135 -280 136 -279
rect 422 -280 423 -279
rect 709 -280 710 -279
rect 849 -280 850 -279
rect 352 -282 353 -281
rect 667 -282 668 -281
rect 730 -282 731 -281
rect 898 -282 899 -281
rect 93 -284 94 -283
rect 352 -284 353 -283
rect 520 -284 521 -283
rect 730 -284 731 -283
rect 758 -284 759 -283
rect 1038 -284 1039 -283
rect 9 -286 10 -285
rect 93 -286 94 -285
rect 478 -286 479 -285
rect 520 -286 521 -285
rect 597 -286 598 -285
rect 709 -286 710 -285
rect 765 -286 766 -285
rect 863 -286 864 -285
rect 9 -288 10 -287
rect 79 -288 80 -287
rect 184 -288 185 -287
rect 597 -288 598 -287
rect 779 -288 780 -287
rect 891 -288 892 -287
rect 184 -290 185 -289
rect 247 -290 248 -289
rect 390 -290 391 -289
rect 765 -290 766 -289
rect 779 -290 780 -289
rect 996 -290 997 -289
rect 247 -292 248 -291
rect 275 -292 276 -291
rect 450 -292 451 -291
rect 478 -292 479 -291
rect 786 -292 787 -291
rect 905 -292 906 -291
rect 254 -294 255 -293
rect 275 -294 276 -293
rect 450 -294 451 -293
rect 751 -294 752 -293
rect 856 -294 857 -293
rect 996 -294 997 -293
rect 254 -296 255 -295
rect 324 -296 325 -295
rect 646 -296 647 -295
rect 786 -296 787 -295
rect 324 -298 325 -297
rect 338 -298 339 -297
rect 569 -298 570 -297
rect 646 -298 647 -297
rect 681 -298 682 -297
rect 856 -298 857 -297
rect 68 -300 69 -299
rect 338 -300 339 -299
rect 653 -300 654 -299
rect 681 -300 682 -299
rect 723 -300 724 -299
rect 751 -300 752 -299
rect 156 -302 157 -301
rect 569 -302 570 -301
rect 653 -302 654 -301
rect 660 -302 661 -301
rect 723 -302 724 -301
rect 807 -302 808 -301
rect 149 -304 150 -303
rect 156 -304 157 -303
rect 660 -304 661 -303
rect 695 -304 696 -303
rect 772 -304 773 -303
rect 807 -304 808 -303
rect 30 -306 31 -305
rect 772 -306 773 -305
rect 54 -308 55 -307
rect 149 -308 150 -307
rect 2 -319 3 -318
rect 40 -319 41 -318
rect 65 -319 66 -318
rect 86 -319 87 -318
rect 93 -319 94 -318
rect 226 -319 227 -318
rect 264 -319 265 -318
rect 275 -319 276 -318
rect 285 -319 286 -318
rect 1192 -319 1193 -318
rect 2 -321 3 -320
rect 44 -321 45 -320
rect 58 -321 59 -320
rect 275 -321 276 -320
rect 310 -321 311 -320
rect 450 -321 451 -320
rect 471 -321 472 -320
rect 544 -321 545 -320
rect 586 -321 587 -320
rect 1059 -321 1060 -320
rect 1101 -321 1102 -320
rect 1171 -321 1172 -320
rect 1178 -321 1179 -320
rect 1202 -321 1203 -320
rect 9 -323 10 -322
rect 30 -323 31 -322
rect 37 -323 38 -322
rect 572 -323 573 -322
rect 604 -323 605 -322
rect 618 -323 619 -322
rect 695 -323 696 -322
rect 1101 -323 1102 -322
rect 1115 -323 1116 -322
rect 1178 -323 1179 -322
rect 9 -325 10 -324
rect 233 -325 234 -324
rect 317 -325 318 -324
rect 499 -325 500 -324
rect 527 -325 528 -324
rect 541 -325 542 -324
rect 702 -325 703 -324
rect 1164 -325 1165 -324
rect 16 -327 17 -326
rect 89 -327 90 -326
rect 93 -327 94 -326
rect 177 -327 178 -326
rect 184 -327 185 -326
rect 502 -327 503 -326
rect 702 -327 703 -326
rect 709 -327 710 -326
rect 758 -327 759 -326
rect 884 -327 885 -326
rect 961 -327 962 -326
rect 1185 -327 1186 -326
rect 16 -329 17 -328
rect 313 -329 314 -328
rect 327 -329 328 -328
rect 597 -329 598 -328
rect 667 -329 668 -328
rect 758 -329 759 -328
rect 884 -329 885 -328
rect 905 -329 906 -328
rect 1031 -329 1032 -328
rect 1059 -329 1060 -328
rect 1129 -329 1130 -328
rect 1150 -329 1151 -328
rect 26 -331 27 -330
rect 191 -331 192 -330
rect 198 -331 199 -330
rect 320 -331 321 -330
rect 359 -331 360 -330
rect 667 -331 668 -330
rect 709 -331 710 -330
rect 723 -331 724 -330
rect 891 -331 892 -330
rect 905 -331 906 -330
rect 996 -331 997 -330
rect 1031 -331 1032 -330
rect 1052 -331 1053 -330
rect 1115 -331 1116 -330
rect 1136 -331 1137 -330
rect 1157 -331 1158 -330
rect 37 -333 38 -332
rect 989 -333 990 -332
rect 1087 -333 1088 -332
rect 1129 -333 1130 -332
rect 44 -335 45 -334
rect 47 -335 48 -334
rect 61 -335 62 -334
rect 233 -335 234 -334
rect 254 -335 255 -334
rect 359 -335 360 -334
rect 394 -335 395 -334
rect 411 -335 412 -334
rect 422 -335 423 -334
rect 478 -335 479 -334
rect 485 -335 486 -334
rect 618 -335 619 -334
rect 653 -335 654 -334
rect 723 -335 724 -334
rect 765 -335 766 -334
rect 996 -335 997 -334
rect 1024 -335 1025 -334
rect 1087 -335 1088 -334
rect 1094 -335 1095 -334
rect 1136 -335 1137 -334
rect 68 -337 69 -336
rect 730 -337 731 -336
rect 786 -337 787 -336
rect 891 -337 892 -336
rect 947 -337 948 -336
rect 1052 -337 1053 -336
rect 72 -339 73 -338
rect 82 -339 83 -338
rect 107 -339 108 -338
rect 110 -339 111 -338
rect 121 -339 122 -338
rect 590 -339 591 -338
rect 625 -339 626 -338
rect 765 -339 766 -338
rect 786 -339 787 -338
rect 814 -339 815 -338
rect 940 -339 941 -338
rect 947 -339 948 -338
rect 982 -339 983 -338
rect 989 -339 990 -338
rect 1045 -339 1046 -338
rect 1094 -339 1095 -338
rect 75 -341 76 -340
rect 1143 -341 1144 -340
rect 79 -343 80 -342
rect 1024 -343 1025 -342
rect 1122 -343 1123 -342
rect 1143 -343 1144 -342
rect 82 -345 83 -344
rect 1066 -345 1067 -344
rect 1073 -345 1074 -344
rect 1122 -345 1123 -344
rect 107 -347 108 -346
rect 135 -347 136 -346
rect 156 -347 157 -346
rect 453 -347 454 -346
rect 471 -347 472 -346
rect 492 -347 493 -346
rect 499 -347 500 -346
rect 562 -347 563 -346
rect 569 -347 570 -346
rect 730 -347 731 -346
rect 814 -347 815 -346
rect 821 -347 822 -346
rect 898 -347 899 -346
rect 940 -347 941 -346
rect 968 -347 969 -346
rect 982 -347 983 -346
rect 1017 -347 1018 -346
rect 1045 -347 1046 -346
rect 110 -349 111 -348
rect 135 -349 136 -348
rect 163 -349 164 -348
rect 478 -349 479 -348
rect 516 -349 517 -348
rect 898 -349 899 -348
rect 954 -349 955 -348
rect 968 -349 969 -348
rect 975 -349 976 -348
rect 1017 -349 1018 -348
rect 1038 -349 1039 -348
rect 1066 -349 1067 -348
rect 96 -351 97 -350
rect 954 -351 955 -350
rect 1003 -351 1004 -350
rect 1038 -351 1039 -350
rect 100 -353 101 -352
rect 163 -353 164 -352
rect 177 -353 178 -352
rect 282 -353 283 -352
rect 303 -353 304 -352
rect 317 -353 318 -352
rect 331 -353 332 -352
rect 422 -353 423 -352
rect 429 -353 430 -352
rect 527 -353 528 -352
rect 555 -353 556 -352
rect 597 -353 598 -352
rect 625 -353 626 -352
rect 632 -353 633 -352
rect 653 -353 654 -352
rect 674 -353 675 -352
rect 800 -353 801 -352
rect 821 -353 822 -352
rect 926 -353 927 -352
rect 975 -353 976 -352
rect 51 -355 52 -354
rect 100 -355 101 -354
rect 114 -355 115 -354
rect 121 -355 122 -354
rect 128 -355 129 -354
rect 184 -355 185 -354
rect 191 -355 192 -354
rect 212 -355 213 -354
rect 219 -355 220 -354
rect 226 -355 227 -354
rect 282 -355 283 -354
rect 373 -355 374 -354
rect 380 -355 381 -354
rect 485 -355 486 -354
rect 509 -355 510 -354
rect 632 -355 633 -354
rect 674 -355 675 -354
rect 779 -355 780 -354
rect 800 -355 801 -354
rect 1209 -355 1210 -354
rect 72 -357 73 -356
rect 114 -357 115 -356
rect 128 -357 129 -356
rect 611 -357 612 -356
rect 779 -357 780 -356
rect 807 -357 808 -356
rect 919 -357 920 -356
rect 926 -357 927 -356
rect 933 -357 934 -356
rect 1003 -357 1004 -356
rect 142 -359 143 -358
rect 219 -359 220 -358
rect 303 -359 304 -358
rect 352 -359 353 -358
rect 366 -359 367 -358
rect 380 -359 381 -358
rect 397 -359 398 -358
rect 1080 -359 1081 -358
rect 86 -361 87 -360
rect 142 -361 143 -360
rect 198 -361 199 -360
rect 205 -361 206 -360
rect 212 -361 213 -360
rect 698 -361 699 -360
rect 772 -361 773 -360
rect 807 -361 808 -360
rect 849 -361 850 -360
rect 933 -361 934 -360
rect 1010 -361 1011 -360
rect 1080 -361 1081 -360
rect 149 -363 150 -362
rect 205 -363 206 -362
rect 289 -363 290 -362
rect 352 -363 353 -362
rect 366 -363 367 -362
rect 642 -363 643 -362
rect 772 -363 773 -362
rect 793 -363 794 -362
rect 828 -363 829 -362
rect 849 -363 850 -362
rect 870 -363 871 -362
rect 919 -363 920 -362
rect 1010 -363 1011 -362
rect 1108 -363 1109 -362
rect 79 -365 80 -364
rect 828 -365 829 -364
rect 149 -367 150 -366
rect 247 -367 248 -366
rect 289 -367 290 -366
rect 551 -367 552 -366
rect 569 -367 570 -366
rect 877 -367 878 -366
rect 247 -369 248 -368
rect 268 -369 269 -368
rect 373 -369 374 -368
rect 520 -369 521 -368
rect 583 -369 584 -368
rect 793 -369 794 -368
rect 835 -369 836 -368
rect 877 -369 878 -368
rect 23 -371 24 -370
rect 835 -371 836 -370
rect 23 -373 24 -372
rect 33 -373 34 -372
rect 261 -373 262 -372
rect 268 -373 269 -372
rect 387 -373 388 -372
rect 1108 -373 1109 -372
rect 261 -375 262 -374
rect 506 -375 507 -374
rect 513 -375 514 -374
rect 555 -375 556 -374
rect 583 -375 584 -374
rect 660 -375 661 -374
rect 751 -375 752 -374
rect 870 -375 871 -374
rect 331 -377 332 -376
rect 660 -377 661 -376
rect 737 -377 738 -376
rect 751 -377 752 -376
rect 345 -379 346 -378
rect 387 -379 388 -378
rect 408 -379 409 -378
rect 961 -379 962 -378
rect 51 -381 52 -380
rect 408 -381 409 -380
rect 415 -381 416 -380
rect 429 -381 430 -380
rect 436 -381 437 -380
rect 695 -381 696 -380
rect 296 -383 297 -382
rect 345 -383 346 -382
rect 415 -383 416 -382
rect 670 -383 671 -382
rect 124 -385 125 -384
rect 296 -385 297 -384
rect 338 -385 339 -384
rect 436 -385 437 -384
rect 450 -385 451 -384
rect 457 -385 458 -384
rect 464 -385 465 -384
rect 492 -385 493 -384
rect 506 -385 507 -384
rect 744 -385 745 -384
rect 124 -387 125 -386
rect 156 -387 157 -386
rect 338 -387 339 -386
rect 576 -387 577 -386
rect 579 -387 580 -386
rect 737 -387 738 -386
rect 324 -389 325 -388
rect 576 -389 577 -388
rect 590 -389 591 -388
rect 1073 -389 1074 -388
rect 240 -391 241 -390
rect 324 -391 325 -390
rect 443 -391 444 -390
rect 457 -391 458 -390
rect 464 -391 465 -390
rect 513 -391 514 -390
rect 520 -391 521 -390
rect 534 -391 535 -390
rect 611 -391 612 -390
rect 646 -391 647 -390
rect 716 -391 717 -390
rect 744 -391 745 -390
rect 58 -393 59 -392
rect 240 -393 241 -392
rect 411 -393 412 -392
rect 716 -393 717 -392
rect 170 -395 171 -394
rect 443 -395 444 -394
rect 534 -395 535 -394
rect 548 -395 549 -394
rect 639 -395 640 -394
rect 646 -395 647 -394
rect 26 -397 27 -396
rect 170 -397 171 -396
rect 254 -397 255 -396
rect 548 -397 549 -396
rect 565 -397 566 -396
rect 639 -397 640 -396
rect 23 -408 24 -407
rect 1108 -408 1109 -407
rect 1129 -408 1130 -407
rect 1213 -408 1214 -407
rect 23 -410 24 -409
rect 264 -410 265 -409
rect 331 -410 332 -409
rect 537 -410 538 -409
rect 548 -410 549 -409
rect 1171 -410 1172 -409
rect 1209 -410 1210 -409
rect 1395 -410 1396 -409
rect 26 -412 27 -411
rect 975 -412 976 -411
rect 1017 -412 1018 -411
rect 1206 -412 1207 -411
rect 30 -414 31 -413
rect 58 -414 59 -413
rect 75 -414 76 -413
rect 121 -414 122 -413
rect 128 -414 129 -413
rect 383 -414 384 -413
rect 408 -414 409 -413
rect 429 -414 430 -413
rect 460 -414 461 -413
rect 919 -414 920 -413
rect 975 -414 976 -413
rect 1202 -414 1203 -413
rect 30 -416 31 -415
rect 940 -416 941 -415
rect 1038 -416 1039 -415
rect 1129 -416 1130 -415
rect 1136 -416 1137 -415
rect 1220 -416 1221 -415
rect 40 -418 41 -417
rect 282 -418 283 -417
rect 331 -418 332 -417
rect 653 -418 654 -417
rect 663 -418 664 -417
rect 1178 -418 1179 -417
rect 44 -420 45 -419
rect 177 -420 178 -419
rect 201 -420 202 -419
rect 205 -420 206 -419
rect 261 -420 262 -419
rect 387 -420 388 -419
rect 401 -420 402 -419
rect 429 -420 430 -419
rect 471 -420 472 -419
rect 513 -420 514 -419
rect 551 -420 552 -419
rect 807 -420 808 -419
rect 814 -420 815 -419
rect 817 -420 818 -419
rect 870 -420 871 -419
rect 940 -420 941 -419
rect 968 -420 969 -419
rect 1038 -420 1039 -419
rect 1045 -420 1046 -419
rect 1136 -420 1137 -419
rect 1143 -420 1144 -419
rect 1227 -420 1228 -419
rect 2 -422 3 -421
rect 44 -422 45 -421
rect 58 -422 59 -421
rect 65 -422 66 -421
rect 79 -422 80 -421
rect 919 -422 920 -421
rect 961 -422 962 -421
rect 1045 -422 1046 -421
rect 1059 -422 1060 -421
rect 1143 -422 1144 -421
rect 1150 -422 1151 -421
rect 1234 -422 1235 -421
rect 9 -424 10 -423
rect 79 -424 80 -423
rect 86 -424 87 -423
rect 177 -424 178 -423
rect 198 -424 199 -423
rect 205 -424 206 -423
rect 261 -424 262 -423
rect 373 -424 374 -423
rect 401 -424 402 -423
rect 611 -424 612 -423
rect 625 -424 626 -423
rect 639 -424 640 -423
rect 670 -424 671 -423
rect 1052 -424 1053 -423
rect 1066 -424 1067 -423
rect 1150 -424 1151 -423
rect 1157 -424 1158 -423
rect 1255 -424 1256 -423
rect 61 -426 62 -425
rect 1178 -426 1179 -425
rect 65 -428 66 -427
rect 555 -428 556 -427
rect 562 -428 563 -427
rect 877 -428 878 -427
rect 898 -428 899 -427
rect 961 -428 962 -427
rect 982 -428 983 -427
rect 1066 -428 1067 -427
rect 1073 -428 1074 -427
rect 1157 -428 1158 -427
rect 47 -430 48 -429
rect 877 -430 878 -429
rect 884 -430 885 -429
rect 898 -430 899 -429
rect 905 -430 906 -429
rect 968 -430 969 -429
rect 1003 -430 1004 -429
rect 1059 -430 1060 -429
rect 1080 -430 1081 -429
rect 1171 -430 1172 -429
rect 86 -432 87 -431
rect 219 -432 220 -431
rect 275 -432 276 -431
rect 387 -432 388 -431
rect 411 -432 412 -431
rect 464 -432 465 -431
rect 478 -432 479 -431
rect 516 -432 517 -431
rect 520 -432 521 -431
rect 555 -432 556 -431
rect 569 -432 570 -431
rect 933 -432 934 -431
rect 1003 -432 1004 -431
rect 1010 -432 1011 -431
rect 89 -434 90 -433
rect 1241 -434 1242 -433
rect 89 -436 90 -435
rect 821 -436 822 -435
rect 828 -436 829 -435
rect 982 -436 983 -435
rect 989 -436 990 -435
rect 1010 -436 1011 -435
rect 93 -438 94 -437
rect 124 -438 125 -437
rect 138 -438 139 -437
rect 1192 -438 1193 -437
rect 72 -440 73 -439
rect 93 -440 94 -439
rect 100 -440 101 -439
rect 408 -440 409 -439
rect 422 -440 423 -439
rect 464 -440 465 -439
rect 478 -440 479 -439
rect 758 -440 759 -439
rect 772 -440 773 -439
rect 821 -440 822 -439
rect 835 -440 836 -439
rect 905 -440 906 -439
rect 1122 -440 1123 -439
rect 1192 -440 1193 -439
rect 33 -442 34 -441
rect 772 -442 773 -441
rect 779 -442 780 -441
rect 835 -442 836 -441
rect 849 -442 850 -441
rect 870 -442 871 -441
rect 1031 -442 1032 -441
rect 1122 -442 1123 -441
rect 100 -444 101 -443
rect 142 -444 143 -443
rect 145 -444 146 -443
rect 828 -444 829 -443
rect 863 -444 864 -443
rect 933 -444 934 -443
rect 107 -446 108 -445
rect 128 -446 129 -445
rect 142 -446 143 -445
rect 184 -446 185 -445
rect 198 -446 199 -445
rect 576 -446 577 -445
rect 590 -446 591 -445
rect 663 -446 664 -445
rect 698 -446 699 -445
rect 1017 -446 1018 -445
rect 107 -448 108 -447
rect 884 -448 885 -447
rect 156 -450 157 -449
rect 548 -450 549 -449
rect 572 -450 573 -449
rect 863 -450 864 -449
rect 163 -452 164 -451
rect 282 -452 283 -451
rect 338 -452 339 -451
rect 562 -452 563 -451
rect 576 -452 577 -451
rect 618 -452 619 -451
rect 632 -452 633 -451
rect 653 -452 654 -451
rect 705 -452 706 -451
rect 1185 -452 1186 -451
rect 170 -454 171 -453
rect 569 -454 570 -453
rect 593 -454 594 -453
rect 695 -454 696 -453
rect 716 -454 717 -453
rect 779 -454 780 -453
rect 793 -454 794 -453
rect 1031 -454 1032 -453
rect 1101 -454 1102 -453
rect 1185 -454 1186 -453
rect 149 -456 150 -455
rect 170 -456 171 -455
rect 184 -456 185 -455
rect 310 -456 311 -455
rect 338 -456 339 -455
rect 492 -456 493 -455
rect 509 -456 510 -455
rect 765 -456 766 -455
rect 800 -456 801 -455
rect 849 -456 850 -455
rect 114 -458 115 -457
rect 765 -458 766 -457
rect 814 -458 815 -457
rect 926 -458 927 -457
rect 114 -460 115 -459
rect 289 -460 290 -459
rect 310 -460 311 -459
rect 317 -460 318 -459
rect 345 -460 346 -459
rect 807 -460 808 -459
rect 856 -460 857 -459
rect 926 -460 927 -459
rect 51 -462 52 -461
rect 289 -462 290 -461
rect 296 -462 297 -461
rect 345 -462 346 -461
rect 373 -462 374 -461
rect 450 -462 451 -461
rect 457 -462 458 -461
rect 471 -462 472 -461
rect 485 -462 486 -461
rect 492 -462 493 -461
rect 520 -462 521 -461
rect 583 -462 584 -461
rect 597 -462 598 -461
rect 632 -462 633 -461
rect 642 -462 643 -461
rect 989 -462 990 -461
rect 51 -464 52 -463
rect 380 -464 381 -463
rect 422 -464 423 -463
rect 793 -464 794 -463
rect 817 -464 818 -463
rect 856 -464 857 -463
rect 149 -466 150 -465
rect 240 -466 241 -465
rect 268 -466 269 -465
rect 275 -466 276 -465
rect 296 -466 297 -465
rect 397 -466 398 -465
rect 425 -466 426 -465
rect 1073 -466 1074 -465
rect 212 -468 213 -467
rect 268 -468 269 -467
rect 366 -468 367 -467
rect 450 -468 451 -467
rect 457 -468 458 -467
rect 590 -468 591 -467
rect 597 -468 598 -467
rect 1248 -468 1249 -467
rect 212 -470 213 -469
rect 233 -470 234 -469
rect 366 -470 367 -469
rect 506 -470 507 -469
rect 534 -470 535 -469
rect 583 -470 584 -469
rect 600 -470 601 -469
rect 996 -470 997 -469
rect 219 -472 220 -471
rect 324 -472 325 -471
rect 380 -472 381 -471
rect 1080 -472 1081 -471
rect 226 -474 227 -473
rect 240 -474 241 -473
rect 303 -474 304 -473
rect 324 -474 325 -473
rect 436 -474 437 -473
rect 485 -474 486 -473
rect 604 -474 605 -473
rect 625 -474 626 -473
rect 646 -474 647 -473
rect 1101 -474 1102 -473
rect 16 -476 17 -475
rect 303 -476 304 -475
rect 317 -476 318 -475
rect 534 -476 535 -475
rect 611 -476 612 -475
rect 1087 -476 1088 -475
rect 16 -478 17 -477
rect 247 -478 248 -477
rect 352 -478 353 -477
rect 436 -478 437 -477
rect 527 -478 528 -477
rect 604 -478 605 -477
rect 614 -478 615 -477
rect 1052 -478 1053 -477
rect 82 -480 83 -479
rect 646 -480 647 -479
rect 681 -480 682 -479
rect 716 -480 717 -479
rect 737 -480 738 -479
rect 758 -480 759 -479
rect 912 -480 913 -479
rect 996 -480 997 -479
rect 1024 -480 1025 -479
rect 1087 -480 1088 -479
rect 159 -482 160 -481
rect 912 -482 913 -481
rect 947 -482 948 -481
rect 1024 -482 1025 -481
rect 191 -484 192 -483
rect 226 -484 227 -483
rect 233 -484 234 -483
rect 394 -484 395 -483
rect 499 -484 500 -483
rect 681 -484 682 -483
rect 751 -484 752 -483
rect 800 -484 801 -483
rect 891 -484 892 -483
rect 947 -484 948 -483
rect 135 -486 136 -485
rect 191 -486 192 -485
rect 254 -486 255 -485
rect 394 -486 395 -485
rect 527 -486 528 -485
rect 1108 -486 1109 -485
rect 135 -488 136 -487
rect 954 -488 955 -487
rect 37 -490 38 -489
rect 954 -490 955 -489
rect 37 -492 38 -491
rect 75 -492 76 -491
rect 163 -492 164 -491
rect 499 -492 500 -491
rect 565 -492 566 -491
rect 737 -492 738 -491
rect 842 -492 843 -491
rect 891 -492 892 -491
rect 352 -494 353 -493
rect 359 -494 360 -493
rect 618 -494 619 -493
rect 674 -494 675 -493
rect 702 -494 703 -493
rect 751 -494 752 -493
rect 786 -494 787 -493
rect 842 -494 843 -493
rect 110 -496 111 -495
rect 359 -496 360 -495
rect 415 -496 416 -495
rect 702 -496 703 -495
rect 730 -496 731 -495
rect 786 -496 787 -495
rect 415 -498 416 -497
rect 1164 -498 1165 -497
rect 502 -500 503 -499
rect 674 -500 675 -499
rect 688 -500 689 -499
rect 730 -500 731 -499
rect 1094 -500 1095 -499
rect 1164 -500 1165 -499
rect 9 -502 10 -501
rect 502 -502 503 -501
rect 688 -502 689 -501
rect 723 -502 724 -501
rect 1094 -502 1095 -501
rect 1115 -502 1116 -501
rect 723 -504 724 -503
rect 744 -504 745 -503
rect 1115 -504 1116 -503
rect 1199 -504 1200 -503
rect 667 -506 668 -505
rect 1199 -506 1200 -505
rect 660 -508 661 -507
rect 667 -508 668 -507
rect 709 -508 710 -507
rect 744 -508 745 -507
rect 443 -510 444 -509
rect 709 -510 710 -509
rect 443 -512 444 -511
rect 530 -512 531 -511
rect 660 -512 661 -511
rect 1262 -512 1263 -511
rect 2 -523 3 -522
rect 1241 -523 1242 -522
rect 1248 -523 1249 -522
rect 1360 -523 1361 -522
rect 1395 -523 1396 -522
rect 1472 -523 1473 -522
rect 1500 -523 1501 -522
rect 1507 -523 1508 -522
rect 2 -525 3 -524
rect 565 -525 566 -524
rect 600 -525 601 -524
rect 1269 -525 1270 -524
rect 16 -527 17 -526
rect 254 -527 255 -526
rect 261 -527 262 -526
rect 457 -527 458 -526
rect 460 -527 461 -526
rect 919 -527 920 -526
rect 1003 -527 1004 -526
rect 1339 -527 1340 -526
rect 30 -529 31 -528
rect 583 -529 584 -528
rect 635 -529 636 -528
rect 758 -529 759 -528
rect 828 -529 829 -528
rect 919 -529 920 -528
rect 940 -529 941 -528
rect 1003 -529 1004 -528
rect 1094 -529 1095 -528
rect 1283 -529 1284 -528
rect 33 -531 34 -530
rect 72 -531 73 -530
rect 75 -531 76 -530
rect 219 -531 220 -530
rect 226 -531 227 -530
rect 380 -531 381 -530
rect 425 -531 426 -530
rect 614 -531 615 -530
rect 660 -531 661 -530
rect 814 -531 815 -530
rect 870 -531 871 -530
rect 940 -531 941 -530
rect 1024 -531 1025 -530
rect 1094 -531 1095 -530
rect 1150 -531 1151 -530
rect 1241 -531 1242 -530
rect 1255 -531 1256 -530
rect 1374 -531 1375 -530
rect 40 -533 41 -532
rect 1206 -533 1207 -532
rect 1213 -533 1214 -532
rect 1304 -533 1305 -532
rect 40 -535 41 -534
rect 1073 -535 1074 -534
rect 1080 -535 1081 -534
rect 1150 -535 1151 -534
rect 1157 -535 1158 -534
rect 1248 -535 1249 -534
rect 1262 -535 1263 -534
rect 1367 -535 1368 -534
rect 47 -537 48 -536
rect 198 -537 199 -536
rect 226 -537 227 -536
rect 275 -537 276 -536
rect 317 -537 318 -536
rect 611 -537 612 -536
rect 614 -537 615 -536
rect 821 -537 822 -536
rect 954 -537 955 -536
rect 1024 -537 1025 -536
rect 1136 -537 1137 -536
rect 1213 -537 1214 -536
rect 1220 -537 1221 -536
rect 1311 -537 1312 -536
rect 72 -539 73 -538
rect 233 -539 234 -538
rect 240 -539 241 -538
rect 261 -539 262 -538
rect 271 -539 272 -538
rect 807 -539 808 -538
rect 912 -539 913 -538
rect 954 -539 955 -538
rect 996 -539 997 -538
rect 1073 -539 1074 -538
rect 1164 -539 1165 -538
rect 1206 -539 1207 -538
rect 1227 -539 1228 -538
rect 1332 -539 1333 -538
rect 110 -541 111 -540
rect 492 -541 493 -540
rect 499 -541 500 -540
rect 1157 -541 1158 -540
rect 1171 -541 1172 -540
rect 1276 -541 1277 -540
rect 114 -543 115 -542
rect 317 -543 318 -542
rect 331 -543 332 -542
rect 509 -543 510 -542
rect 520 -543 521 -542
rect 527 -543 528 -542
rect 530 -543 531 -542
rect 751 -543 752 -542
rect 779 -543 780 -542
rect 828 -543 829 -542
rect 842 -543 843 -542
rect 912 -543 913 -542
rect 933 -543 934 -542
rect 996 -543 997 -542
rect 1017 -543 1018 -542
rect 1080 -543 1081 -542
rect 1108 -543 1109 -542
rect 1164 -543 1165 -542
rect 1178 -543 1179 -542
rect 1255 -543 1256 -542
rect 114 -545 115 -544
rect 1325 -545 1326 -544
rect 117 -547 118 -546
rect 401 -547 402 -546
rect 408 -547 409 -546
rect 499 -547 500 -546
rect 502 -547 503 -546
rect 1101 -547 1102 -546
rect 1122 -547 1123 -546
rect 1171 -547 1172 -546
rect 1185 -547 1186 -546
rect 1262 -547 1263 -546
rect 135 -549 136 -548
rect 1045 -549 1046 -548
rect 1192 -549 1193 -548
rect 1290 -549 1291 -548
rect 121 -551 122 -550
rect 135 -551 136 -550
rect 142 -551 143 -550
rect 877 -551 878 -550
rect 898 -551 899 -550
rect 1192 -551 1193 -550
rect 1199 -551 1200 -550
rect 1297 -551 1298 -550
rect 121 -553 122 -552
rect 247 -553 248 -552
rect 275 -553 276 -552
rect 383 -553 384 -552
rect 401 -553 402 -552
rect 569 -553 570 -552
rect 611 -553 612 -552
rect 1136 -553 1137 -552
rect 1234 -553 1235 -552
rect 1353 -553 1354 -552
rect 44 -555 45 -554
rect 569 -555 570 -554
rect 625 -555 626 -554
rect 751 -555 752 -554
rect 765 -555 766 -554
rect 1178 -555 1179 -554
rect 142 -557 143 -556
rect 201 -557 202 -556
rect 212 -557 213 -556
rect 331 -557 332 -556
rect 338 -557 339 -556
rect 415 -557 416 -556
rect 443 -557 444 -556
rect 492 -557 493 -556
rect 509 -557 510 -556
rect 842 -557 843 -556
rect 849 -557 850 -556
rect 898 -557 899 -556
rect 968 -557 969 -556
rect 1045 -557 1046 -556
rect 1129 -557 1130 -556
rect 1199 -557 1200 -556
rect 58 -559 59 -558
rect 415 -559 416 -558
rect 450 -559 451 -558
rect 453 -559 454 -558
rect 457 -559 458 -558
rect 562 -559 563 -558
rect 625 -559 626 -558
rect 1318 -559 1319 -558
rect 37 -561 38 -560
rect 58 -561 59 -560
rect 138 -561 139 -560
rect 212 -561 213 -560
rect 233 -561 234 -560
rect 310 -561 311 -560
rect 338 -561 339 -560
rect 373 -561 374 -560
rect 450 -561 451 -560
rect 513 -561 514 -560
rect 534 -561 535 -560
rect 1185 -561 1186 -560
rect 79 -563 80 -562
rect 534 -563 535 -562
rect 548 -563 549 -562
rect 583 -563 584 -562
rect 628 -563 629 -562
rect 1108 -563 1109 -562
rect 1143 -563 1144 -562
rect 1234 -563 1235 -562
rect 65 -565 66 -564
rect 548 -565 549 -564
rect 660 -565 661 -564
rect 905 -565 906 -564
rect 1031 -565 1032 -564
rect 1101 -565 1102 -564
rect 65 -567 66 -566
rect 163 -567 164 -566
rect 170 -567 171 -566
rect 254 -567 255 -566
rect 345 -567 346 -566
rect 422 -567 423 -566
rect 464 -567 465 -566
rect 520 -567 521 -566
rect 663 -567 664 -566
rect 779 -567 780 -566
rect 786 -567 787 -566
rect 821 -567 822 -566
rect 835 -567 836 -566
rect 905 -567 906 -566
rect 1031 -567 1032 -566
rect 1346 -567 1347 -566
rect 5 -569 6 -568
rect 422 -569 423 -568
rect 481 -569 482 -568
rect 982 -569 983 -568
rect 1052 -569 1053 -568
rect 1129 -569 1130 -568
rect 23 -571 24 -570
rect 464 -571 465 -570
rect 485 -571 486 -570
rect 513 -571 514 -570
rect 670 -571 671 -570
rect 1115 -571 1116 -570
rect 23 -573 24 -572
rect 324 -573 325 -572
rect 348 -573 349 -572
rect 968 -573 969 -572
rect 1010 -573 1011 -572
rect 1052 -573 1053 -572
rect 1059 -573 1060 -572
rect 1143 -573 1144 -572
rect 79 -575 80 -574
rect 100 -575 101 -574
rect 107 -575 108 -574
rect 982 -575 983 -574
rect 989 -575 990 -574
rect 1059 -575 1060 -574
rect 96 -577 97 -576
rect 100 -577 101 -576
rect 107 -577 108 -576
rect 159 -577 160 -576
rect 163 -577 164 -576
rect 184 -577 185 -576
rect 191 -577 192 -576
rect 198 -577 199 -576
rect 240 -577 241 -576
rect 268 -577 269 -576
rect 324 -577 325 -576
rect 471 -577 472 -576
rect 506 -577 507 -576
rect 849 -577 850 -576
rect 863 -577 864 -576
rect 933 -577 934 -576
rect 947 -577 948 -576
rect 1010 -577 1011 -576
rect 19 -579 20 -578
rect 184 -579 185 -578
rect 191 -579 192 -578
rect 205 -579 206 -578
rect 247 -579 248 -578
rect 257 -579 258 -578
rect 268 -579 269 -578
rect 705 -579 706 -578
rect 723 -579 724 -578
rect 870 -579 871 -578
rect 884 -579 885 -578
rect 947 -579 948 -578
rect 145 -581 146 -580
rect 793 -581 794 -580
rect 800 -581 801 -580
rect 877 -581 878 -580
rect 926 -581 927 -580
rect 989 -581 990 -580
rect 170 -583 171 -582
rect 219 -583 220 -582
rect 250 -583 251 -582
rect 786 -583 787 -582
rect 856 -583 857 -582
rect 926 -583 927 -582
rect 86 -585 87 -584
rect 856 -585 857 -584
rect 86 -587 87 -586
rect 555 -587 556 -586
rect 618 -587 619 -586
rect 1115 -587 1116 -586
rect 205 -589 206 -588
rect 303 -589 304 -588
rect 352 -589 353 -588
rect 446 -589 447 -588
rect 453 -589 454 -588
rect 485 -589 486 -588
rect 506 -589 507 -588
rect 975 -589 976 -588
rect 282 -591 283 -590
rect 618 -591 619 -590
rect 674 -591 675 -590
rect 1220 -591 1221 -590
rect 51 -593 52 -592
rect 282 -593 283 -592
rect 303 -593 304 -592
rect 352 -593 353 -592
rect 359 -593 360 -592
rect 408 -593 409 -592
rect 436 -593 437 -592
rect 674 -593 675 -592
rect 681 -593 682 -592
rect 758 -593 759 -592
rect 765 -593 766 -592
rect 1038 -593 1039 -592
rect 359 -595 360 -594
rect 387 -595 388 -594
rect 418 -595 419 -594
rect 436 -595 437 -594
rect 471 -595 472 -594
rect 562 -595 563 -594
rect 590 -595 591 -594
rect 681 -595 682 -594
rect 688 -595 689 -594
rect 723 -595 724 -594
rect 730 -595 731 -594
rect 800 -595 801 -594
rect 891 -595 892 -594
rect 975 -595 976 -594
rect 89 -597 90 -596
rect 891 -597 892 -596
rect 961 -597 962 -596
rect 1038 -597 1039 -596
rect 289 -599 290 -598
rect 387 -599 388 -598
rect 418 -599 419 -598
rect 1122 -599 1123 -598
rect 289 -601 290 -600
rect 394 -601 395 -600
rect 443 -601 444 -600
rect 590 -601 591 -600
rect 646 -601 647 -600
rect 730 -601 731 -600
rect 737 -601 738 -600
rect 807 -601 808 -600
rect 863 -601 864 -600
rect 961 -601 962 -600
rect 373 -603 374 -602
rect 597 -603 598 -602
rect 653 -603 654 -602
rect 737 -603 738 -602
rect 744 -603 745 -602
rect 814 -603 815 -602
rect 394 -605 395 -604
rect 429 -605 430 -604
rect 478 -605 479 -604
rect 597 -605 598 -604
rect 653 -605 654 -604
rect 709 -605 710 -604
rect 716 -605 717 -604
rect 793 -605 794 -604
rect 44 -607 45 -606
rect 709 -607 710 -606
rect 747 -607 748 -606
rect 884 -607 885 -606
rect 149 -609 150 -608
rect 429 -609 430 -608
rect 541 -609 542 -608
rect 555 -609 556 -608
rect 576 -609 577 -608
rect 646 -609 647 -608
rect 667 -609 668 -608
rect 688 -609 689 -608
rect 695 -609 696 -608
rect 1066 -609 1067 -608
rect 37 -611 38 -610
rect 576 -611 577 -610
rect 632 -611 633 -610
rect 716 -611 717 -610
rect 772 -611 773 -610
rect 835 -611 836 -610
rect 149 -613 150 -612
rect 380 -613 381 -612
rect 390 -613 391 -612
rect 1066 -613 1067 -612
rect 366 -615 367 -614
rect 541 -615 542 -614
rect 632 -615 633 -614
rect 695 -615 696 -614
rect 702 -615 703 -614
rect 1227 -615 1228 -614
rect 156 -617 157 -616
rect 702 -617 703 -616
rect 772 -617 773 -616
rect 1034 -617 1035 -616
rect 128 -619 129 -618
rect 156 -619 157 -618
rect 296 -619 297 -618
rect 366 -619 367 -618
rect 667 -619 668 -618
rect 1017 -619 1018 -618
rect 9 -621 10 -620
rect 296 -621 297 -620
rect 9 -623 10 -622
rect 604 -623 605 -622
rect 93 -625 94 -624
rect 128 -625 129 -624
rect 604 -625 605 -624
rect 698 -625 699 -624
rect 51 -627 52 -626
rect 93 -627 94 -626
rect 37 -638 38 -637
rect 324 -638 325 -637
rect 383 -638 384 -637
rect 730 -638 731 -637
rect 747 -638 748 -637
rect 996 -638 997 -637
rect 1034 -638 1035 -637
rect 1374 -638 1375 -637
rect 1472 -638 1473 -637
rect 1528 -638 1529 -637
rect 2 -640 3 -639
rect 324 -640 325 -639
rect 387 -640 388 -639
rect 450 -640 451 -639
rect 506 -640 507 -639
rect 772 -640 773 -639
rect 807 -640 808 -639
rect 1437 -640 1438 -639
rect 1507 -640 1508 -639
rect 1514 -640 1515 -639
rect 5 -642 6 -641
rect 1472 -642 1473 -641
rect 44 -644 45 -643
rect 1178 -644 1179 -643
rect 1206 -644 1207 -643
rect 1381 -644 1382 -643
rect 44 -646 45 -645
rect 233 -646 234 -645
rect 282 -646 283 -645
rect 345 -646 346 -645
rect 387 -646 388 -645
rect 541 -646 542 -645
rect 544 -646 545 -645
rect 1451 -646 1452 -645
rect 47 -648 48 -647
rect 422 -648 423 -647
rect 443 -648 444 -647
rect 548 -648 549 -647
rect 614 -648 615 -647
rect 751 -648 752 -647
rect 807 -648 808 -647
rect 926 -648 927 -647
rect 940 -648 941 -647
rect 996 -648 997 -647
rect 1101 -648 1102 -647
rect 1178 -648 1179 -647
rect 1255 -648 1256 -647
rect 1388 -648 1389 -647
rect 30 -650 31 -649
rect 422 -650 423 -649
rect 429 -650 430 -649
rect 443 -650 444 -649
rect 446 -650 447 -649
rect 1458 -650 1459 -649
rect 30 -652 31 -651
rect 352 -652 353 -651
rect 408 -652 409 -651
rect 450 -652 451 -651
rect 471 -652 472 -651
rect 772 -652 773 -651
rect 870 -652 871 -651
rect 1031 -652 1032 -651
rect 1059 -652 1060 -651
rect 1101 -652 1102 -651
rect 1150 -652 1151 -651
rect 1255 -652 1256 -651
rect 1262 -652 1263 -651
rect 1395 -652 1396 -651
rect 65 -654 66 -653
rect 93 -654 94 -653
rect 100 -654 101 -653
rect 170 -654 171 -653
rect 233 -654 234 -653
rect 390 -654 391 -653
rect 415 -654 416 -653
rect 660 -654 661 -653
rect 663 -654 664 -653
rect 1339 -654 1340 -653
rect 1346 -654 1347 -653
rect 1493 -654 1494 -653
rect 65 -656 66 -655
rect 219 -656 220 -655
rect 261 -656 262 -655
rect 282 -656 283 -655
rect 296 -656 297 -655
rect 751 -656 752 -655
rect 870 -656 871 -655
rect 1094 -656 1095 -655
rect 1150 -656 1151 -655
rect 1164 -656 1165 -655
rect 1227 -656 1228 -655
rect 1339 -656 1340 -655
rect 1353 -656 1354 -655
rect 1500 -656 1501 -655
rect 23 -658 24 -657
rect 261 -658 262 -657
rect 296 -658 297 -657
rect 394 -658 395 -657
rect 401 -658 402 -657
rect 1094 -658 1095 -657
rect 1157 -658 1158 -657
rect 1262 -658 1263 -657
rect 1283 -658 1284 -657
rect 1402 -658 1403 -657
rect 23 -660 24 -659
rect 310 -660 311 -659
rect 345 -660 346 -659
rect 464 -660 465 -659
rect 506 -660 507 -659
rect 681 -660 682 -659
rect 730 -660 731 -659
rect 737 -660 738 -659
rect 744 -660 745 -659
rect 1374 -660 1375 -659
rect 9 -662 10 -661
rect 681 -662 682 -661
rect 702 -662 703 -661
rect 737 -662 738 -661
rect 744 -662 745 -661
rect 1045 -662 1046 -661
rect 1052 -662 1053 -661
rect 1283 -662 1284 -661
rect 1290 -662 1291 -661
rect 1409 -662 1410 -661
rect 79 -664 80 -663
rect 401 -664 402 -663
rect 415 -664 416 -663
rect 621 -664 622 -663
rect 628 -664 629 -663
rect 1115 -664 1116 -663
rect 1171 -664 1172 -663
rect 1290 -664 1291 -663
rect 1304 -664 1305 -663
rect 1416 -664 1417 -663
rect 79 -666 80 -665
rect 121 -666 122 -665
rect 128 -666 129 -665
rect 170 -666 171 -665
rect 219 -666 220 -665
rect 317 -666 318 -665
rect 348 -666 349 -665
rect 408 -666 409 -665
rect 436 -666 437 -665
rect 471 -666 472 -665
rect 509 -666 510 -665
rect 534 -666 535 -665
rect 548 -666 549 -665
rect 583 -666 584 -665
rect 597 -666 598 -665
rect 926 -666 927 -665
rect 940 -666 941 -665
rect 1206 -666 1207 -665
rect 1248 -666 1249 -665
rect 1346 -666 1347 -665
rect 1360 -666 1361 -665
rect 1444 -666 1445 -665
rect 58 -668 59 -667
rect 583 -668 584 -667
rect 614 -668 615 -667
rect 1164 -668 1165 -667
rect 1171 -668 1172 -667
rect 1234 -668 1235 -667
rect 1297 -668 1298 -667
rect 1360 -668 1361 -667
rect 1367 -668 1368 -667
rect 1521 -668 1522 -667
rect 58 -670 59 -669
rect 156 -670 157 -669
rect 268 -670 269 -669
rect 1367 -670 1368 -669
rect 61 -672 62 -671
rect 1297 -672 1298 -671
rect 1311 -672 1312 -671
rect 1423 -672 1424 -671
rect 86 -674 87 -673
rect 429 -674 430 -673
rect 436 -674 437 -673
rect 604 -674 605 -673
rect 628 -674 629 -673
rect 1269 -674 1270 -673
rect 1318 -674 1319 -673
rect 1430 -674 1431 -673
rect 86 -676 87 -675
rect 331 -676 332 -675
rect 359 -676 360 -675
rect 394 -676 395 -675
rect 604 -676 605 -675
rect 695 -676 696 -675
rect 702 -676 703 -675
rect 793 -676 794 -675
rect 842 -676 843 -675
rect 1269 -676 1270 -675
rect 1325 -676 1326 -675
rect 1479 -676 1480 -675
rect 93 -678 94 -677
rect 600 -678 601 -677
rect 635 -678 636 -677
rect 1003 -678 1004 -677
rect 1010 -678 1011 -677
rect 1052 -678 1053 -677
rect 1073 -678 1074 -677
rect 1115 -678 1116 -677
rect 1129 -678 1130 -677
rect 1234 -678 1235 -677
rect 1332 -678 1333 -677
rect 1486 -678 1487 -677
rect 19 -680 20 -679
rect 1073 -680 1074 -679
rect 1080 -680 1081 -679
rect 1129 -680 1130 -679
rect 1143 -680 1144 -679
rect 1248 -680 1249 -679
rect 72 -682 73 -681
rect 1143 -682 1144 -681
rect 1199 -682 1200 -681
rect 1311 -682 1312 -681
rect 72 -684 73 -683
rect 523 -684 524 -683
rect 747 -684 748 -683
rect 1185 -684 1186 -683
rect 1199 -684 1200 -683
rect 1241 -684 1242 -683
rect 96 -686 97 -685
rect 1227 -686 1228 -685
rect 100 -688 101 -687
rect 618 -688 619 -687
rect 761 -688 762 -687
rect 1157 -688 1158 -687
rect 1213 -688 1214 -687
rect 1318 -688 1319 -687
rect 114 -690 115 -689
rect 373 -690 374 -689
rect 380 -690 381 -689
rect 464 -690 465 -689
rect 478 -690 479 -689
rect 1080 -690 1081 -689
rect 1108 -690 1109 -689
rect 1213 -690 1214 -689
rect 1220 -690 1221 -689
rect 1325 -690 1326 -689
rect 114 -692 115 -691
rect 919 -692 920 -691
rect 943 -692 944 -691
rect 1276 -692 1277 -691
rect 121 -694 122 -693
rect 481 -694 482 -693
rect 618 -694 619 -693
rect 1304 -694 1305 -693
rect 128 -696 129 -695
rect 418 -696 419 -695
rect 425 -696 426 -695
rect 695 -696 696 -695
rect 765 -696 766 -695
rect 1353 -696 1354 -695
rect 135 -698 136 -697
rect 173 -698 174 -697
rect 247 -698 248 -697
rect 331 -698 332 -697
rect 359 -698 360 -697
rect 485 -698 486 -697
rect 513 -698 514 -697
rect 765 -698 766 -697
rect 779 -698 780 -697
rect 793 -698 794 -697
rect 856 -698 857 -697
rect 1185 -698 1186 -697
rect 12 -700 13 -699
rect 856 -700 857 -699
rect 877 -700 878 -699
rect 1045 -700 1046 -699
rect 1066 -700 1067 -699
rect 1108 -700 1109 -699
rect 1136 -700 1137 -699
rect 1241 -700 1242 -699
rect 107 -702 108 -701
rect 247 -702 248 -701
rect 310 -702 311 -701
rect 527 -702 528 -701
rect 537 -702 538 -701
rect 779 -702 780 -701
rect 849 -702 850 -701
rect 877 -702 878 -701
rect 919 -702 920 -701
rect 989 -702 990 -701
rect 1017 -702 1018 -701
rect 1059 -702 1060 -701
rect 1087 -702 1088 -701
rect 1276 -702 1277 -701
rect 107 -704 108 -703
rect 240 -704 241 -703
rect 313 -704 314 -703
rect 478 -704 479 -703
rect 485 -704 486 -703
rect 492 -704 493 -703
rect 499 -704 500 -703
rect 527 -704 528 -703
rect 653 -704 654 -703
rect 1220 -704 1221 -703
rect 149 -706 150 -705
rect 156 -706 157 -705
rect 177 -706 178 -705
rect 240 -706 241 -705
rect 317 -706 318 -705
rect 716 -706 717 -705
rect 835 -706 836 -705
rect 989 -706 990 -705
rect 1024 -706 1025 -705
rect 1332 -706 1333 -705
rect 149 -708 150 -707
rect 625 -708 626 -707
rect 639 -708 640 -707
rect 653 -708 654 -707
rect 667 -708 668 -707
rect 1017 -708 1018 -707
rect 1038 -708 1039 -707
rect 1087 -708 1088 -707
rect 103 -710 104 -709
rect 639 -710 640 -709
rect 667 -710 668 -709
rect 709 -710 710 -709
rect 716 -710 717 -709
rect 800 -710 801 -709
rect 814 -710 815 -709
rect 835 -710 836 -709
rect 849 -710 850 -709
rect 891 -710 892 -709
rect 947 -710 948 -709
rect 1003 -710 1004 -709
rect 177 -712 178 -711
rect 184 -712 185 -711
rect 338 -712 339 -711
rect 513 -712 514 -711
rect 565 -712 566 -711
rect 1038 -712 1039 -711
rect 184 -714 185 -713
rect 212 -714 213 -713
rect 338 -714 339 -713
rect 674 -714 675 -713
rect 709 -714 710 -713
rect 723 -714 724 -713
rect 786 -714 787 -713
rect 800 -714 801 -713
rect 814 -714 815 -713
rect 821 -714 822 -713
rect 954 -714 955 -713
rect 1010 -714 1011 -713
rect 163 -716 164 -715
rect 212 -716 213 -715
rect 355 -716 356 -715
rect 947 -716 948 -715
rect 961 -716 962 -715
rect 1066 -716 1067 -715
rect 142 -718 143 -717
rect 163 -718 164 -717
rect 355 -718 356 -717
rect 457 -718 458 -717
rect 492 -718 493 -717
rect 660 -718 661 -717
rect 786 -718 787 -717
rect 1122 -718 1123 -717
rect 142 -720 143 -719
rect 271 -720 272 -719
rect 366 -720 367 -719
rect 723 -720 724 -719
rect 758 -720 759 -719
rect 1122 -720 1123 -719
rect 75 -722 76 -721
rect 271 -722 272 -721
rect 373 -722 374 -721
rect 520 -722 521 -721
rect 632 -722 633 -721
rect 891 -722 892 -721
rect 898 -722 899 -721
rect 954 -722 955 -721
rect 964 -722 965 -721
rect 1465 -722 1466 -721
rect 289 -724 290 -723
rect 632 -724 633 -723
rect 646 -724 647 -723
rect 674 -724 675 -723
rect 758 -724 759 -723
rect 1192 -724 1193 -723
rect 226 -726 227 -725
rect 289 -726 290 -725
rect 457 -726 458 -725
rect 576 -726 577 -725
rect 590 -726 591 -725
rect 646 -726 647 -725
rect 821 -726 822 -725
rect 887 -726 888 -725
rect 905 -726 906 -725
rect 961 -726 962 -725
rect 968 -726 969 -725
rect 1024 -726 1025 -725
rect 226 -728 227 -727
rect 254 -728 255 -727
rect 499 -728 500 -727
rect 541 -728 542 -727
rect 555 -728 556 -727
rect 590 -728 591 -727
rect 611 -728 612 -727
rect 1192 -728 1193 -727
rect 205 -730 206 -729
rect 254 -730 255 -729
rect 534 -730 535 -729
rect 555 -730 556 -729
rect 569 -730 570 -729
rect 576 -730 577 -729
rect 611 -730 612 -729
rect 1136 -730 1137 -729
rect 205 -732 206 -731
rect 275 -732 276 -731
rect 562 -732 563 -731
rect 569 -732 570 -731
rect 863 -732 864 -731
rect 898 -732 899 -731
rect 905 -732 906 -731
rect 975 -732 976 -731
rect 982 -732 983 -731
rect 1507 -732 1508 -731
rect 117 -734 118 -733
rect 982 -734 983 -733
rect 275 -736 276 -735
rect 303 -736 304 -735
rect 366 -736 367 -735
rect 975 -736 976 -735
rect 198 -738 199 -737
rect 303 -738 304 -737
rect 380 -738 381 -737
rect 562 -738 563 -737
rect 863 -738 864 -737
rect 933 -738 934 -737
rect 51 -740 52 -739
rect 198 -740 199 -739
rect 828 -740 829 -739
rect 933 -740 934 -739
rect 51 -742 52 -741
rect 75 -742 76 -741
rect 117 -742 118 -741
rect 828 -742 829 -741
rect 912 -742 913 -741
rect 968 -742 969 -741
rect 884 -744 885 -743
rect 912 -744 913 -743
rect 842 -746 843 -745
rect 884 -746 885 -745
rect 2 -757 3 -756
rect 1094 -757 1095 -756
rect 2 -759 3 -758
rect 611 -759 612 -758
rect 614 -759 615 -758
rect 1437 -759 1438 -758
rect 9 -761 10 -760
rect 338 -761 339 -760
rect 369 -761 370 -760
rect 943 -761 944 -760
rect 1066 -761 1067 -760
rect 1094 -761 1095 -760
rect 1437 -761 1438 -760
rect 1458 -761 1459 -760
rect 9 -763 10 -762
rect 642 -763 643 -762
rect 649 -763 650 -762
rect 1297 -763 1298 -762
rect 1458 -763 1459 -762
rect 1472 -763 1473 -762
rect 12 -765 13 -764
rect 968 -765 969 -764
rect 1066 -765 1067 -764
rect 1213 -765 1214 -764
rect 1472 -765 1473 -764
rect 1493 -765 1494 -764
rect 23 -767 24 -766
rect 271 -767 272 -766
rect 310 -767 311 -766
rect 712 -767 713 -766
rect 747 -767 748 -766
rect 1213 -767 1214 -766
rect 16 -769 17 -768
rect 23 -769 24 -768
rect 47 -769 48 -768
rect 632 -769 633 -768
rect 653 -769 654 -768
rect 663 -769 664 -768
rect 775 -769 776 -768
rect 1521 -769 1522 -768
rect 16 -771 17 -770
rect 184 -771 185 -770
rect 226 -771 227 -770
rect 366 -771 367 -770
rect 394 -771 395 -770
rect 397 -771 398 -770
rect 485 -771 486 -770
rect 488 -771 489 -770
rect 509 -771 510 -770
rect 1045 -771 1046 -770
rect 1164 -771 1165 -770
rect 1297 -771 1298 -770
rect 58 -773 59 -772
rect 1507 -773 1508 -772
rect 58 -775 59 -774
rect 79 -775 80 -774
rect 117 -775 118 -774
rect 723 -775 724 -774
rect 884 -775 885 -774
rect 1248 -775 1249 -774
rect 51 -777 52 -776
rect 79 -777 80 -776
rect 121 -777 122 -776
rect 310 -777 311 -776
rect 324 -777 325 -776
rect 422 -777 423 -776
rect 485 -777 486 -776
rect 527 -777 528 -776
rect 534 -777 535 -776
rect 1332 -777 1333 -776
rect 51 -779 52 -778
rect 296 -779 297 -778
rect 324 -779 325 -778
rect 439 -779 440 -778
rect 520 -779 521 -778
rect 530 -779 531 -778
rect 537 -779 538 -778
rect 751 -779 752 -778
rect 887 -779 888 -778
rect 1444 -779 1445 -778
rect 61 -781 62 -780
rect 1073 -781 1074 -780
rect 1164 -781 1165 -780
rect 1325 -781 1326 -780
rect 1332 -781 1333 -780
rect 1346 -781 1347 -780
rect 1444 -781 1445 -780
rect 1486 -781 1487 -780
rect 65 -783 66 -782
rect 460 -783 461 -782
rect 520 -783 521 -782
rect 604 -783 605 -782
rect 611 -783 612 -782
rect 898 -783 899 -782
rect 940 -783 941 -782
rect 1423 -783 1424 -782
rect 65 -785 66 -784
rect 317 -785 318 -784
rect 338 -785 339 -784
rect 352 -785 353 -784
rect 394 -785 395 -784
rect 401 -785 402 -784
rect 422 -785 423 -784
rect 576 -785 577 -784
rect 583 -785 584 -784
rect 604 -785 605 -784
rect 618 -785 619 -784
rect 702 -785 703 -784
rect 723 -785 724 -784
rect 800 -785 801 -784
rect 856 -785 857 -784
rect 898 -785 899 -784
rect 943 -785 944 -784
rect 1255 -785 1256 -784
rect 72 -787 73 -786
rect 1360 -787 1361 -786
rect 72 -789 73 -788
rect 261 -789 262 -788
rect 296 -789 297 -788
rect 768 -789 769 -788
rect 800 -789 801 -788
rect 821 -789 822 -788
rect 856 -789 857 -788
rect 947 -789 948 -788
rect 968 -789 969 -788
rect 1101 -789 1102 -788
rect 1150 -789 1151 -788
rect 1255 -789 1256 -788
rect 1360 -789 1361 -788
rect 1409 -789 1410 -788
rect 75 -791 76 -790
rect 1185 -791 1186 -790
rect 1199 -791 1200 -790
rect 1346 -791 1347 -790
rect 1409 -791 1410 -790
rect 1430 -791 1431 -790
rect 100 -793 101 -792
rect 1423 -793 1424 -792
rect 1430 -793 1431 -792
rect 1451 -793 1452 -792
rect 100 -795 101 -794
rect 359 -795 360 -794
rect 401 -795 402 -794
rect 408 -795 409 -794
rect 464 -795 465 -794
rect 576 -795 577 -794
rect 597 -795 598 -794
rect 961 -795 962 -794
rect 1017 -795 1018 -794
rect 1073 -795 1074 -794
rect 1101 -795 1102 -794
rect 1129 -795 1130 -794
rect 1199 -795 1200 -794
rect 1234 -795 1235 -794
rect 1248 -795 1249 -794
rect 1283 -795 1284 -794
rect 1451 -795 1452 -794
rect 1465 -795 1466 -794
rect 114 -797 115 -796
rect 1325 -797 1326 -796
rect 1465 -797 1466 -796
rect 1479 -797 1480 -796
rect 114 -799 115 -798
rect 282 -799 283 -798
rect 408 -799 409 -798
rect 415 -799 416 -798
rect 464 -799 465 -798
rect 1122 -799 1123 -798
rect 1129 -799 1130 -798
rect 1192 -799 1193 -798
rect 1234 -799 1235 -798
rect 1269 -799 1270 -798
rect 1283 -799 1284 -798
rect 1311 -799 1312 -798
rect 1479 -799 1480 -798
rect 1500 -799 1501 -798
rect 121 -801 122 -800
rect 177 -801 178 -800
rect 184 -801 185 -800
rect 303 -801 304 -800
rect 425 -801 426 -800
rect 1122 -801 1123 -800
rect 1171 -801 1172 -800
rect 1311 -801 1312 -800
rect 1500 -801 1501 -800
rect 1514 -801 1515 -800
rect 131 -803 132 -802
rect 170 -803 171 -802
rect 177 -803 178 -802
rect 212 -803 213 -802
rect 226 -803 227 -802
rect 380 -803 381 -802
rect 523 -803 524 -802
rect 989 -803 990 -802
rect 1017 -803 1018 -802
rect 1262 -803 1263 -802
rect 1269 -803 1270 -802
rect 1304 -803 1305 -802
rect 1514 -803 1515 -802
rect 1528 -803 1529 -802
rect 107 -805 108 -804
rect 170 -805 171 -804
rect 205 -805 206 -804
rect 317 -805 318 -804
rect 380 -805 381 -804
rect 555 -805 556 -804
rect 569 -805 570 -804
rect 884 -805 885 -804
rect 891 -805 892 -804
rect 1150 -805 1151 -804
rect 1192 -805 1193 -804
rect 1227 -805 1228 -804
rect 107 -807 108 -806
rect 219 -807 220 -806
rect 236 -807 237 -806
rect 282 -807 283 -806
rect 289 -807 290 -806
rect 303 -807 304 -806
rect 436 -807 437 -806
rect 555 -807 556 -806
rect 618 -807 619 -806
rect 926 -807 927 -806
rect 989 -807 990 -806
rect 1052 -807 1053 -806
rect 1115 -807 1116 -806
rect 1171 -807 1172 -806
rect 1227 -807 1228 -806
rect 1290 -807 1291 -806
rect 30 -809 31 -808
rect 1052 -809 1053 -808
rect 30 -811 31 -810
rect 450 -811 451 -810
rect 467 -811 468 -810
rect 1290 -811 1291 -810
rect 135 -813 136 -812
rect 691 -813 692 -812
rect 695 -813 696 -812
rect 702 -813 703 -812
rect 779 -813 780 -812
rect 1304 -813 1305 -812
rect 135 -815 136 -814
rect 163 -815 164 -814
rect 205 -815 206 -814
rect 1503 -815 1504 -814
rect 138 -817 139 -816
rect 772 -817 773 -816
rect 779 -817 780 -816
rect 793 -817 794 -816
rect 814 -817 815 -816
rect 821 -817 822 -816
rect 905 -817 906 -816
rect 926 -817 927 -816
rect 1038 -817 1039 -816
rect 1486 -817 1487 -816
rect 93 -819 94 -818
rect 814 -819 815 -818
rect 905 -819 906 -818
rect 954 -819 955 -818
rect 1038 -819 1039 -818
rect 1080 -819 1081 -818
rect 93 -821 94 -820
rect 506 -821 507 -820
rect 534 -821 535 -820
rect 597 -821 598 -820
rect 632 -821 633 -820
rect 674 -821 675 -820
rect 681 -821 682 -820
rect 695 -821 696 -820
rect 730 -821 731 -820
rect 772 -821 773 -820
rect 786 -821 787 -820
rect 1185 -821 1186 -820
rect 142 -823 143 -822
rect 359 -823 360 -822
rect 429 -823 430 -822
rect 674 -823 675 -822
rect 688 -823 689 -822
rect 730 -823 731 -822
rect 758 -823 759 -822
rect 954 -823 955 -822
rect 1045 -823 1046 -822
rect 1087 -823 1088 -822
rect 86 -825 87 -824
rect 429 -825 430 -824
rect 436 -825 437 -824
rect 891 -825 892 -824
rect 919 -825 920 -824
rect 961 -825 962 -824
rect 1080 -825 1081 -824
rect 1136 -825 1137 -824
rect 86 -827 87 -826
rect 709 -827 710 -826
rect 758 -827 759 -826
rect 807 -827 808 -826
rect 919 -827 920 -826
rect 996 -827 997 -826
rect 1087 -827 1088 -826
rect 1206 -827 1207 -826
rect 103 -829 104 -828
rect 142 -829 143 -828
rect 163 -829 164 -828
rect 1493 -829 1494 -828
rect 212 -831 213 -830
rect 366 -831 367 -830
rect 450 -831 451 -830
rect 716 -831 717 -830
rect 793 -831 794 -830
rect 835 -831 836 -830
rect 947 -831 948 -830
rect 996 -831 997 -830
rect 1136 -831 1137 -830
rect 1178 -831 1179 -830
rect 1206 -831 1207 -830
rect 1241 -831 1242 -830
rect 219 -833 220 -832
rect 268 -833 269 -832
rect 492 -833 493 -832
rect 681 -833 682 -832
rect 709 -833 710 -832
rect 1024 -833 1025 -832
rect 1241 -833 1242 -832
rect 1276 -833 1277 -832
rect 240 -835 241 -834
rect 289 -835 290 -834
rect 331 -835 332 -834
rect 492 -835 493 -834
rect 506 -835 507 -834
rect 744 -835 745 -834
rect 1024 -835 1025 -834
rect 1108 -835 1109 -834
rect 1276 -835 1277 -834
rect 1339 -835 1340 -834
rect 233 -837 234 -836
rect 240 -837 241 -836
rect 254 -837 255 -836
rect 352 -837 353 -836
rect 541 -837 542 -836
rect 1031 -837 1032 -836
rect 1108 -837 1109 -836
rect 1143 -837 1144 -836
rect 191 -839 192 -838
rect 233 -839 234 -838
rect 261 -839 262 -838
rect 663 -839 664 -838
rect 667 -839 668 -838
rect 751 -839 752 -838
rect 912 -839 913 -838
rect 1031 -839 1032 -838
rect 1143 -839 1144 -838
rect 1318 -839 1319 -838
rect 191 -841 192 -840
rect 275 -841 276 -840
rect 331 -841 332 -840
rect 373 -841 374 -840
rect 541 -841 542 -840
rect 807 -841 808 -840
rect 863 -841 864 -840
rect 912 -841 913 -840
rect 999 -841 1000 -840
rect 1339 -841 1340 -840
rect 128 -843 129 -842
rect 275 -843 276 -842
rect 373 -843 374 -842
rect 513 -843 514 -842
rect 544 -843 545 -842
rect 765 -843 766 -842
rect 1157 -843 1158 -842
rect 1318 -843 1319 -842
rect 37 -845 38 -844
rect 513 -845 514 -844
rect 548 -845 549 -844
rect 583 -845 584 -844
rect 600 -845 601 -844
rect 786 -845 787 -844
rect 838 -845 839 -844
rect 1157 -845 1158 -844
rect 128 -847 129 -846
rect 1353 -847 1354 -846
rect 198 -849 199 -848
rect 254 -849 255 -848
rect 268 -849 269 -848
rect 345 -849 346 -848
rect 530 -849 531 -848
rect 548 -849 549 -848
rect 551 -849 552 -848
rect 982 -849 983 -848
rect 1353 -849 1354 -848
rect 1367 -849 1368 -848
rect 198 -851 199 -850
rect 247 -851 248 -850
rect 345 -851 346 -850
rect 355 -851 356 -850
rect 562 -851 563 -850
rect 1178 -851 1179 -850
rect 1367 -851 1368 -850
rect 1374 -851 1375 -850
rect 44 -853 45 -852
rect 247 -853 248 -852
rect 562 -853 563 -852
rect 590 -853 591 -852
rect 639 -853 640 -852
rect 982 -853 983 -852
rect 1374 -853 1375 -852
rect 1381 -853 1382 -852
rect 44 -855 45 -854
rect 716 -855 717 -854
rect 737 -855 738 -854
rect 744 -855 745 -854
rect 765 -855 766 -854
rect 933 -855 934 -854
rect 1381 -855 1382 -854
rect 1388 -855 1389 -854
rect 166 -857 167 -856
rect 590 -857 591 -856
rect 646 -857 647 -856
rect 667 -857 668 -856
rect 737 -857 738 -856
rect 877 -857 878 -856
rect 933 -857 934 -856
rect 1003 -857 1004 -856
rect 1388 -857 1389 -856
rect 1395 -857 1396 -856
rect 457 -859 458 -858
rect 877 -859 878 -858
rect 1395 -859 1396 -858
rect 1402 -859 1403 -858
rect 457 -861 458 -860
rect 1220 -861 1221 -860
rect 1402 -861 1403 -860
rect 1416 -861 1417 -860
rect 569 -863 570 -862
rect 835 -863 836 -862
rect 625 -865 626 -864
rect 1003 -865 1004 -864
rect 40 -867 41 -866
rect 625 -867 626 -866
rect 646 -867 647 -866
rect 1262 -867 1263 -866
rect 653 -869 654 -868
rect 1115 -869 1116 -868
rect 656 -871 657 -870
rect 870 -871 871 -870
rect 660 -873 661 -872
rect 863 -873 864 -872
rect 870 -873 871 -872
rect 975 -873 976 -872
rect 149 -875 150 -874
rect 660 -875 661 -874
rect 761 -875 762 -874
rect 1220 -875 1221 -874
rect 149 -877 150 -876
rect 156 -877 157 -876
rect 828 -877 829 -876
rect 1416 -877 1417 -876
rect 156 -879 157 -878
rect 387 -879 388 -878
rect 639 -879 640 -878
rect 828 -879 829 -878
rect 975 -879 976 -878
rect 1010 -879 1011 -878
rect 369 -881 370 -880
rect 387 -881 388 -880
rect 1010 -881 1011 -880
rect 1059 -881 1060 -880
rect 842 -883 843 -882
rect 1059 -883 1060 -882
rect 842 -885 843 -884
rect 849 -885 850 -884
rect 537 -887 538 -886
rect 849 -887 850 -886
rect 40 -898 41 -897
rect 359 -898 360 -897
rect 376 -898 377 -897
rect 1178 -898 1179 -897
rect 1318 -898 1319 -897
rect 1426 -898 1427 -897
rect 1503 -898 1504 -897
rect 1514 -898 1515 -897
rect 44 -900 45 -899
rect 1101 -900 1102 -899
rect 1178 -900 1179 -899
rect 1234 -900 1235 -899
rect 51 -902 52 -901
rect 464 -902 465 -901
rect 467 -902 468 -901
rect 1073 -902 1074 -901
rect 1234 -902 1235 -901
rect 1255 -902 1256 -901
rect 51 -904 52 -903
rect 296 -904 297 -903
rect 334 -904 335 -903
rect 338 -904 339 -903
rect 352 -904 353 -903
rect 359 -904 360 -903
rect 387 -904 388 -903
rect 551 -904 552 -903
rect 646 -904 647 -903
rect 1038 -904 1039 -903
rect 1066 -904 1067 -903
rect 1069 -904 1070 -903
rect 1073 -904 1074 -903
rect 1500 -904 1501 -903
rect 30 -906 31 -905
rect 387 -906 388 -905
rect 429 -906 430 -905
rect 436 -906 437 -905
rect 443 -906 444 -905
rect 464 -906 465 -905
rect 492 -906 493 -905
rect 649 -906 650 -905
rect 656 -906 657 -905
rect 730 -906 731 -905
rect 747 -906 748 -905
rect 758 -906 759 -905
rect 761 -906 762 -905
rect 1297 -906 1298 -905
rect 30 -908 31 -907
rect 170 -908 171 -907
rect 184 -908 185 -907
rect 243 -908 244 -907
rect 296 -908 297 -907
rect 1052 -908 1053 -907
rect 1066 -908 1067 -907
rect 1108 -908 1109 -907
rect 1297 -908 1298 -907
rect 1374 -908 1375 -907
rect 16 -910 17 -909
rect 170 -910 171 -909
rect 184 -910 185 -909
rect 191 -910 192 -909
rect 198 -910 199 -909
rect 369 -910 370 -909
rect 436 -910 437 -909
rect 527 -910 528 -909
rect 534 -910 535 -909
rect 562 -910 563 -909
rect 660 -910 661 -909
rect 1045 -910 1046 -909
rect 1094 -910 1095 -909
rect 1255 -910 1256 -909
rect 1374 -910 1375 -909
rect 1437 -910 1438 -909
rect 65 -912 66 -911
rect 642 -912 643 -911
rect 691 -912 692 -911
rect 1010 -912 1011 -911
rect 1017 -912 1018 -911
rect 1318 -912 1319 -911
rect 1437 -912 1438 -911
rect 1493 -912 1494 -911
rect 65 -914 66 -913
rect 79 -914 80 -913
rect 100 -914 101 -913
rect 492 -914 493 -913
rect 495 -914 496 -913
rect 646 -914 647 -913
rect 705 -914 706 -913
rect 1164 -914 1165 -913
rect 79 -916 80 -915
rect 93 -916 94 -915
rect 100 -916 101 -915
rect 205 -916 206 -915
rect 212 -916 213 -915
rect 429 -916 430 -915
rect 450 -916 451 -915
rect 600 -916 601 -915
rect 639 -916 640 -915
rect 1094 -916 1095 -915
rect 16 -918 17 -917
rect 93 -918 94 -917
rect 114 -918 115 -917
rect 233 -918 234 -917
rect 240 -918 241 -917
rect 443 -918 444 -917
rect 509 -918 510 -917
rect 674 -918 675 -917
rect 709 -918 710 -917
rect 1409 -918 1410 -917
rect 9 -920 10 -919
rect 674 -920 675 -919
rect 712 -920 713 -919
rect 1304 -920 1305 -919
rect 9 -922 10 -921
rect 72 -922 73 -921
rect 96 -922 97 -921
rect 233 -922 234 -921
rect 338 -922 339 -921
rect 618 -922 619 -921
rect 639 -922 640 -921
rect 992 -922 993 -921
rect 1045 -922 1046 -921
rect 1122 -922 1123 -921
rect 1143 -922 1144 -921
rect 1409 -922 1410 -921
rect 72 -924 73 -923
rect 142 -924 143 -923
rect 145 -924 146 -923
rect 1052 -924 1053 -923
rect 1122 -924 1123 -923
rect 1136 -924 1137 -923
rect 1143 -924 1144 -923
rect 1199 -924 1200 -923
rect 1290 -924 1291 -923
rect 1304 -924 1305 -923
rect 114 -926 115 -925
rect 310 -926 311 -925
rect 352 -926 353 -925
rect 460 -926 461 -925
rect 513 -926 514 -925
rect 527 -926 528 -925
rect 534 -926 535 -925
rect 618 -926 619 -925
rect 667 -926 668 -925
rect 709 -926 710 -925
rect 730 -926 731 -925
rect 800 -926 801 -925
rect 807 -926 808 -925
rect 1360 -926 1361 -925
rect 142 -928 143 -927
rect 1430 -928 1431 -927
rect 163 -930 164 -929
rect 226 -930 227 -929
rect 310 -930 311 -929
rect 415 -930 416 -929
rect 513 -930 514 -929
rect 632 -930 633 -929
rect 754 -930 755 -929
rect 1227 -930 1228 -929
rect 1290 -930 1291 -929
rect 1353 -930 1354 -929
rect 1360 -930 1361 -929
rect 1423 -930 1424 -929
rect 37 -932 38 -931
rect 1227 -932 1228 -931
rect 1353 -932 1354 -931
rect 1416 -932 1417 -931
rect 37 -934 38 -933
rect 156 -934 157 -933
rect 163 -934 164 -933
rect 478 -934 479 -933
rect 520 -934 521 -933
rect 667 -934 668 -933
rect 758 -934 759 -933
rect 1276 -934 1277 -933
rect 1416 -934 1417 -933
rect 1465 -934 1466 -933
rect 2 -936 3 -935
rect 520 -936 521 -935
rect 537 -936 538 -935
rect 1325 -936 1326 -935
rect 2 -938 3 -937
rect 695 -938 696 -937
rect 768 -938 769 -937
rect 1444 -938 1445 -937
rect 131 -940 132 -939
rect 695 -940 696 -939
rect 800 -940 801 -939
rect 891 -940 892 -939
rect 908 -940 909 -939
rect 1332 -940 1333 -939
rect 1444 -940 1445 -939
rect 1472 -940 1473 -939
rect 156 -942 157 -941
rect 653 -942 654 -941
rect 807 -942 808 -941
rect 856 -942 857 -941
rect 891 -942 892 -941
rect 905 -942 906 -941
rect 940 -942 941 -941
rect 954 -942 955 -941
rect 975 -942 976 -941
rect 978 -942 979 -941
rect 989 -942 990 -941
rect 1038 -942 1039 -941
rect 1129 -942 1130 -941
rect 1136 -942 1137 -941
rect 1199 -942 1200 -941
rect 1248 -942 1249 -941
rect 1325 -942 1326 -941
rect 1381 -942 1382 -941
rect 177 -944 178 -943
rect 226 -944 227 -943
rect 380 -944 381 -943
rect 450 -944 451 -943
rect 478 -944 479 -943
rect 877 -944 878 -943
rect 943 -944 944 -943
rect 1164 -944 1165 -943
rect 1248 -944 1249 -943
rect 1283 -944 1284 -943
rect 1332 -944 1333 -943
rect 1388 -944 1389 -943
rect 128 -946 129 -945
rect 177 -946 178 -945
rect 191 -946 192 -945
rect 261 -946 262 -945
rect 275 -946 276 -945
rect 380 -946 381 -945
rect 415 -946 416 -945
rect 1185 -946 1186 -945
rect 1283 -946 1284 -945
rect 1346 -946 1347 -945
rect 1381 -946 1382 -945
rect 1451 -946 1452 -945
rect 121 -948 122 -947
rect 128 -948 129 -947
rect 198 -948 199 -947
rect 236 -948 237 -947
rect 254 -948 255 -947
rect 275 -948 276 -947
rect 373 -948 374 -947
rect 1451 -948 1452 -947
rect 121 -950 122 -949
rect 149 -950 150 -949
rect 205 -950 206 -949
rect 373 -950 374 -949
rect 537 -950 538 -949
rect 1171 -950 1172 -949
rect 1185 -950 1186 -949
rect 1241 -950 1242 -949
rect 1388 -950 1389 -949
rect 1458 -950 1459 -949
rect 149 -952 150 -951
rect 810 -952 811 -951
rect 824 -952 825 -951
rect 926 -952 927 -951
rect 975 -952 976 -951
rect 982 -952 983 -951
rect 1010 -952 1011 -951
rect 1423 -952 1424 -951
rect 212 -954 213 -953
rect 303 -954 304 -953
rect 541 -954 542 -953
rect 1220 -954 1221 -953
rect 1241 -954 1242 -953
rect 1269 -954 1270 -953
rect 254 -956 255 -955
rect 324 -956 325 -955
rect 541 -956 542 -955
rect 562 -956 563 -955
rect 576 -956 577 -955
rect 660 -956 661 -955
rect 677 -956 678 -955
rect 1220 -956 1221 -955
rect 1269 -956 1270 -955
rect 1311 -956 1312 -955
rect 261 -958 262 -957
rect 289 -958 290 -957
rect 303 -958 304 -957
rect 394 -958 395 -957
rect 544 -958 545 -957
rect 590 -958 591 -957
rect 828 -958 829 -957
rect 905 -958 906 -957
rect 926 -958 927 -957
rect 933 -958 934 -957
rect 1059 -958 1060 -957
rect 1458 -958 1459 -957
rect 44 -960 45 -959
rect 544 -960 545 -959
rect 548 -960 549 -959
rect 1430 -960 1431 -959
rect 289 -962 290 -961
rect 408 -962 409 -961
rect 551 -962 552 -961
rect 1346 -962 1347 -961
rect 324 -964 325 -963
rect 345 -964 346 -963
rect 394 -964 395 -963
rect 751 -964 752 -963
rect 828 -964 829 -963
rect 1276 -964 1277 -963
rect 1311 -964 1312 -963
rect 1339 -964 1340 -963
rect 247 -966 248 -965
rect 345 -966 346 -965
rect 401 -966 402 -965
rect 408 -966 409 -965
rect 555 -966 556 -965
rect 576 -966 577 -965
rect 590 -966 591 -965
rect 597 -966 598 -965
rect 831 -966 832 -965
rect 1031 -966 1032 -965
rect 1059 -966 1060 -965
rect 1080 -966 1081 -965
rect 1129 -966 1130 -965
rect 1192 -966 1193 -965
rect 1339 -966 1340 -965
rect 1395 -966 1396 -965
rect 86 -968 87 -967
rect 555 -968 556 -967
rect 597 -968 598 -967
rect 737 -968 738 -967
rect 838 -968 839 -967
rect 1479 -968 1480 -967
rect 86 -970 87 -969
rect 107 -970 108 -969
rect 219 -970 220 -969
rect 401 -970 402 -969
rect 723 -970 724 -969
rect 737 -970 738 -969
rect 849 -970 850 -969
rect 859 -970 860 -969
rect 877 -970 878 -969
rect 884 -970 885 -969
rect 933 -970 934 -969
rect 947 -970 948 -969
rect 996 -970 997 -969
rect 1395 -970 1396 -969
rect 107 -972 108 -971
rect 135 -972 136 -971
rect 219 -972 220 -971
rect 506 -972 507 -971
rect 625 -972 626 -971
rect 849 -972 850 -971
rect 856 -972 857 -971
rect 954 -972 955 -971
rect 968 -972 969 -971
rect 996 -972 997 -971
rect 1003 -972 1004 -971
rect 1031 -972 1032 -971
rect 1069 -972 1070 -971
rect 1108 -972 1109 -971
rect 1171 -972 1172 -971
rect 1213 -972 1214 -971
rect 135 -974 136 -973
rect 457 -974 458 -973
rect 583 -974 584 -973
rect 625 -974 626 -973
rect 884 -974 885 -973
rect 912 -974 913 -973
rect 947 -974 948 -973
rect 961 -974 962 -973
rect 1003 -974 1004 -973
rect 1115 -974 1116 -973
rect 1192 -974 1193 -973
rect 1367 -974 1368 -973
rect 247 -976 248 -975
rect 299 -976 300 -975
rect 331 -976 332 -975
rect 457 -976 458 -975
rect 611 -976 612 -975
rect 968 -976 969 -975
rect 1080 -976 1081 -975
rect 1150 -976 1151 -975
rect 1213 -976 1214 -975
rect 1262 -976 1263 -975
rect 1367 -976 1368 -975
rect 1486 -976 1487 -975
rect 282 -978 283 -977
rect 506 -978 507 -977
rect 611 -978 612 -977
rect 702 -978 703 -977
rect 716 -978 717 -977
rect 1262 -978 1263 -977
rect 282 -980 283 -979
rect 569 -980 570 -979
rect 632 -980 633 -979
rect 702 -980 703 -979
rect 863 -980 864 -979
rect 961 -980 962 -979
rect 1087 -980 1088 -979
rect 1115 -980 1116 -979
rect 1150 -980 1151 -979
rect 1206 -980 1207 -979
rect 366 -982 367 -981
rect 723 -982 724 -981
rect 835 -982 836 -981
rect 1206 -982 1207 -981
rect 268 -984 269 -983
rect 366 -984 367 -983
rect 422 -984 423 -983
rect 583 -984 584 -983
rect 688 -984 689 -983
rect 912 -984 913 -983
rect 1087 -984 1088 -983
rect 1157 -984 1158 -983
rect 268 -986 269 -985
rect 317 -986 318 -985
rect 422 -986 423 -985
rect 744 -986 745 -985
rect 751 -986 752 -985
rect 1157 -986 1158 -985
rect 317 -988 318 -987
rect 688 -988 689 -987
rect 691 -988 692 -987
rect 716 -988 717 -987
rect 744 -988 745 -987
rect 1101 -988 1102 -987
rect 569 -990 570 -989
rect 765 -990 766 -989
rect 786 -990 787 -989
rect 835 -990 836 -989
rect 863 -990 864 -989
rect 870 -990 871 -989
rect 653 -992 654 -991
rect 870 -992 871 -991
rect 765 -994 766 -993
rect 772 -994 773 -993
rect 786 -994 787 -993
rect 814 -994 815 -993
rect 548 -996 549 -995
rect 772 -996 773 -995
rect 793 -996 794 -995
rect 814 -996 815 -995
rect 779 -998 780 -997
rect 793 -998 794 -997
rect 779 -1000 780 -999
rect 842 -1000 843 -999
rect 821 -1002 822 -1001
rect 842 -1002 843 -1001
rect 821 -1004 822 -1003
rect 1017 -1004 1018 -1003
rect 72 -1015 73 -1014
rect 758 -1015 759 -1014
rect 796 -1015 797 -1014
rect 1038 -1015 1039 -1014
rect 1164 -1015 1165 -1014
rect 1591 -1015 1592 -1014
rect 72 -1017 73 -1016
rect 82 -1017 83 -1016
rect 93 -1017 94 -1016
rect 968 -1017 969 -1016
rect 989 -1017 990 -1016
rect 1234 -1017 1235 -1016
rect 1276 -1017 1277 -1016
rect 1570 -1017 1571 -1016
rect 93 -1019 94 -1018
rect 219 -1019 220 -1018
rect 226 -1019 227 -1018
rect 299 -1019 300 -1018
rect 310 -1019 311 -1018
rect 537 -1019 538 -1018
rect 541 -1019 542 -1018
rect 1311 -1019 1312 -1018
rect 1325 -1019 1326 -1018
rect 1486 -1019 1487 -1018
rect 2 -1021 3 -1020
rect 541 -1021 542 -1020
rect 548 -1021 549 -1020
rect 793 -1021 794 -1020
rect 821 -1021 822 -1020
rect 1409 -1021 1410 -1020
rect 1423 -1021 1424 -1020
rect 1444 -1021 1445 -1020
rect 1451 -1021 1452 -1020
rect 1535 -1021 1536 -1020
rect 2 -1023 3 -1022
rect 268 -1023 269 -1022
rect 310 -1023 311 -1022
rect 894 -1023 895 -1022
rect 908 -1023 909 -1022
rect 1514 -1023 1515 -1022
rect 44 -1025 45 -1024
rect 226 -1025 227 -1024
rect 240 -1025 241 -1024
rect 250 -1025 251 -1024
rect 254 -1025 255 -1024
rect 702 -1025 703 -1024
rect 705 -1025 706 -1024
rect 1451 -1025 1452 -1024
rect 23 -1027 24 -1026
rect 44 -1027 45 -1026
rect 96 -1027 97 -1026
rect 583 -1027 584 -1026
rect 590 -1027 591 -1026
rect 688 -1027 689 -1026
rect 691 -1027 692 -1026
rect 968 -1027 969 -1026
rect 992 -1027 993 -1026
rect 1059 -1027 1060 -1026
rect 1108 -1027 1109 -1026
rect 1234 -1027 1235 -1026
rect 1255 -1027 1256 -1026
rect 1409 -1027 1410 -1026
rect 1437 -1027 1438 -1026
rect 1598 -1027 1599 -1026
rect 23 -1029 24 -1028
rect 40 -1029 41 -1028
rect 107 -1029 108 -1028
rect 142 -1029 143 -1028
rect 184 -1029 185 -1028
rect 334 -1029 335 -1028
rect 376 -1029 377 -1028
rect 569 -1029 570 -1028
rect 576 -1029 577 -1028
rect 597 -1029 598 -1028
rect 600 -1029 601 -1028
rect 1255 -1029 1256 -1028
rect 1283 -1029 1284 -1028
rect 1444 -1029 1445 -1028
rect 37 -1031 38 -1030
rect 597 -1031 598 -1030
rect 607 -1031 608 -1030
rect 1052 -1031 1053 -1030
rect 1143 -1031 1144 -1030
rect 1283 -1031 1284 -1030
rect 1297 -1031 1298 -1030
rect 1479 -1031 1480 -1030
rect 37 -1033 38 -1032
rect 58 -1033 59 -1032
rect 107 -1033 108 -1032
rect 177 -1033 178 -1032
rect 184 -1033 185 -1032
rect 352 -1033 353 -1032
rect 390 -1033 391 -1032
rect 1066 -1033 1067 -1032
rect 1192 -1033 1193 -1032
rect 1472 -1033 1473 -1032
rect 33 -1035 34 -1034
rect 177 -1035 178 -1034
rect 201 -1035 202 -1034
rect 219 -1035 220 -1034
rect 240 -1035 241 -1034
rect 754 -1035 755 -1034
rect 842 -1035 843 -1034
rect 905 -1035 906 -1034
rect 940 -1035 941 -1034
rect 1059 -1035 1060 -1034
rect 1192 -1035 1193 -1034
rect 1213 -1035 1214 -1034
rect 1304 -1035 1305 -1034
rect 1423 -1035 1424 -1034
rect 58 -1037 59 -1036
rect 198 -1037 199 -1036
rect 247 -1037 248 -1036
rect 576 -1037 577 -1036
rect 593 -1037 594 -1036
rect 1318 -1037 1319 -1036
rect 1332 -1037 1333 -1036
rect 1500 -1037 1501 -1036
rect 79 -1039 80 -1038
rect 842 -1039 843 -1038
rect 856 -1039 857 -1038
rect 891 -1039 892 -1038
rect 940 -1039 941 -1038
rect 996 -1039 997 -1038
rect 1052 -1039 1053 -1038
rect 1458 -1039 1459 -1038
rect 86 -1041 87 -1040
rect 198 -1041 199 -1040
rect 247 -1041 248 -1040
rect 275 -1041 276 -1040
rect 394 -1041 395 -1040
rect 551 -1041 552 -1040
rect 569 -1041 570 -1040
rect 695 -1041 696 -1040
rect 702 -1041 703 -1040
rect 709 -1041 710 -1040
rect 716 -1041 717 -1040
rect 754 -1041 755 -1040
rect 758 -1041 759 -1040
rect 856 -1041 857 -1040
rect 859 -1041 860 -1040
rect 1416 -1041 1417 -1040
rect 114 -1043 115 -1042
rect 268 -1043 269 -1042
rect 275 -1043 276 -1042
rect 352 -1043 353 -1042
rect 415 -1043 416 -1042
rect 583 -1043 584 -1042
rect 611 -1043 612 -1042
rect 716 -1043 717 -1042
rect 719 -1043 720 -1042
rect 1325 -1043 1326 -1042
rect 1339 -1043 1340 -1042
rect 1507 -1043 1508 -1042
rect 114 -1045 115 -1044
rect 296 -1045 297 -1044
rect 331 -1045 332 -1044
rect 695 -1045 696 -1044
rect 733 -1045 734 -1044
rect 1038 -1045 1039 -1044
rect 1136 -1045 1137 -1044
rect 1213 -1045 1214 -1044
rect 1290 -1045 1291 -1044
rect 1458 -1045 1459 -1044
rect 30 -1047 31 -1046
rect 331 -1047 332 -1046
rect 408 -1047 409 -1046
rect 415 -1047 416 -1046
rect 432 -1047 433 -1046
rect 660 -1047 661 -1046
rect 663 -1047 664 -1046
rect 1577 -1047 1578 -1046
rect 30 -1049 31 -1048
rect 86 -1049 87 -1048
rect 142 -1049 143 -1048
rect 205 -1049 206 -1048
rect 254 -1049 255 -1048
rect 632 -1049 633 -1048
rect 660 -1049 661 -1048
rect 814 -1049 815 -1048
rect 859 -1049 860 -1048
rect 1437 -1049 1438 -1048
rect 156 -1051 157 -1050
rect 296 -1051 297 -1050
rect 338 -1051 339 -1050
rect 632 -1051 633 -1050
rect 667 -1051 668 -1050
rect 821 -1051 822 -1050
rect 863 -1051 864 -1050
rect 989 -1051 990 -1050
rect 996 -1051 997 -1050
rect 1024 -1051 1025 -1050
rect 1171 -1051 1172 -1050
rect 1318 -1051 1319 -1050
rect 1346 -1051 1347 -1050
rect 1521 -1051 1522 -1050
rect 135 -1053 136 -1052
rect 156 -1053 157 -1052
rect 205 -1053 206 -1052
rect 824 -1053 825 -1052
rect 870 -1053 871 -1052
rect 1402 -1053 1403 -1052
rect 121 -1055 122 -1054
rect 135 -1055 136 -1054
rect 261 -1055 262 -1054
rect 373 -1055 374 -1054
rect 408 -1055 409 -1054
rect 681 -1055 682 -1054
rect 730 -1055 731 -1054
rect 814 -1055 815 -1054
rect 936 -1055 937 -1054
rect 1290 -1055 1291 -1054
rect 1311 -1055 1312 -1054
rect 1430 -1055 1431 -1054
rect 121 -1057 122 -1056
rect 191 -1057 192 -1056
rect 212 -1057 213 -1056
rect 261 -1057 262 -1056
rect 338 -1057 339 -1056
rect 481 -1057 482 -1056
rect 485 -1057 486 -1056
rect 548 -1057 549 -1056
rect 562 -1057 563 -1056
rect 709 -1057 710 -1056
rect 747 -1057 748 -1056
rect 807 -1057 808 -1056
rect 954 -1057 955 -1056
rect 1066 -1057 1067 -1056
rect 1178 -1057 1179 -1056
rect 1332 -1057 1333 -1056
rect 1353 -1057 1354 -1056
rect 1528 -1057 1529 -1056
rect 9 -1059 10 -1058
rect 212 -1059 213 -1058
rect 359 -1059 360 -1058
rect 373 -1059 374 -1058
rect 394 -1059 395 -1058
rect 730 -1059 731 -1058
rect 793 -1059 794 -1058
rect 1402 -1059 1403 -1058
rect 145 -1061 146 -1060
rect 191 -1061 192 -1060
rect 359 -1061 360 -1060
rect 380 -1061 381 -1060
rect 446 -1061 447 -1060
rect 1024 -1061 1025 -1060
rect 1045 -1061 1046 -1060
rect 1171 -1061 1172 -1060
rect 1185 -1061 1186 -1060
rect 1339 -1061 1340 -1060
rect 1367 -1061 1368 -1060
rect 1563 -1061 1564 -1060
rect 163 -1063 164 -1062
rect 380 -1063 381 -1062
rect 460 -1063 461 -1062
rect 1276 -1063 1277 -1062
rect 1374 -1063 1375 -1062
rect 1542 -1063 1543 -1062
rect 166 -1065 167 -1064
rect 1178 -1065 1179 -1064
rect 1199 -1065 1200 -1064
rect 1353 -1065 1354 -1064
rect 1381 -1065 1382 -1064
rect 1549 -1065 1550 -1064
rect 464 -1067 465 -1066
rect 870 -1067 871 -1066
rect 933 -1067 934 -1066
rect 1045 -1067 1046 -1066
rect 1073 -1067 1074 -1066
rect 1185 -1067 1186 -1066
rect 1220 -1067 1221 -1066
rect 1374 -1067 1375 -1066
rect 1388 -1067 1389 -1066
rect 1556 -1067 1557 -1066
rect 9 -1069 10 -1068
rect 1220 -1069 1221 -1068
rect 1227 -1069 1228 -1068
rect 1381 -1069 1382 -1068
rect 1395 -1069 1396 -1068
rect 1584 -1069 1585 -1068
rect 243 -1071 244 -1070
rect 464 -1071 465 -1070
rect 478 -1071 479 -1070
rect 520 -1071 521 -1070
rect 534 -1071 535 -1070
rect 1416 -1071 1417 -1070
rect 429 -1073 430 -1072
rect 478 -1073 479 -1072
rect 485 -1073 486 -1072
rect 828 -1073 829 -1072
rect 933 -1073 934 -1072
rect 1269 -1073 1270 -1072
rect 492 -1075 493 -1074
rect 1346 -1075 1347 -1074
rect 355 -1077 356 -1076
rect 492 -1077 493 -1076
rect 495 -1077 496 -1076
rect 863 -1077 864 -1076
rect 947 -1077 948 -1076
rect 1073 -1077 1074 -1076
rect 1080 -1077 1081 -1076
rect 1367 -1077 1368 -1076
rect 499 -1079 500 -1078
rect 534 -1079 535 -1078
rect 544 -1079 545 -1078
rect 681 -1079 682 -1078
rect 828 -1079 829 -1078
rect 1136 -1079 1137 -1078
rect 1241 -1079 1242 -1078
rect 1388 -1079 1389 -1078
rect 471 -1081 472 -1080
rect 499 -1081 500 -1080
rect 555 -1081 556 -1080
rect 807 -1081 808 -1080
rect 877 -1081 878 -1080
rect 947 -1081 948 -1080
rect 954 -1081 955 -1080
rect 1493 -1081 1494 -1080
rect 443 -1083 444 -1082
rect 471 -1083 472 -1082
rect 555 -1083 556 -1082
rect 873 -1083 874 -1082
rect 957 -1083 958 -1082
rect 1157 -1083 1158 -1082
rect 1248 -1083 1249 -1082
rect 1395 -1083 1396 -1082
rect 443 -1085 444 -1084
rect 1143 -1085 1144 -1084
rect 1248 -1085 1249 -1084
rect 1360 -1085 1361 -1084
rect 562 -1087 563 -1086
rect 831 -1087 832 -1086
rect 835 -1087 836 -1086
rect 877 -1087 878 -1086
rect 975 -1087 976 -1086
rect 1108 -1087 1109 -1086
rect 1115 -1087 1116 -1086
rect 1227 -1087 1228 -1086
rect 1262 -1087 1263 -1086
rect 1430 -1087 1431 -1086
rect 79 -1089 80 -1088
rect 1262 -1089 1263 -1088
rect 611 -1091 612 -1090
rect 772 -1091 773 -1090
rect 779 -1091 780 -1090
rect 1115 -1091 1116 -1090
rect 1129 -1091 1130 -1090
rect 1269 -1091 1270 -1090
rect 250 -1093 251 -1092
rect 772 -1093 773 -1092
rect 831 -1093 832 -1092
rect 1304 -1093 1305 -1092
rect 628 -1095 629 -1094
rect 1297 -1095 1298 -1094
rect 653 -1097 654 -1096
rect 1080 -1097 1081 -1096
rect 1087 -1097 1088 -1096
rect 1241 -1097 1242 -1096
rect 604 -1099 605 -1098
rect 653 -1099 654 -1098
rect 670 -1099 671 -1098
rect 1164 -1099 1165 -1098
rect 1206 -1099 1207 -1098
rect 1360 -1099 1361 -1098
rect 674 -1101 675 -1100
rect 1465 -1101 1466 -1100
rect 674 -1103 675 -1102
rect 744 -1103 745 -1102
rect 751 -1103 752 -1102
rect 779 -1103 780 -1102
rect 835 -1103 836 -1102
rect 982 -1103 983 -1102
rect 1003 -1103 1004 -1102
rect 1157 -1103 1158 -1102
rect 513 -1105 514 -1104
rect 744 -1105 745 -1104
rect 751 -1105 752 -1104
rect 1122 -1105 1123 -1104
rect 401 -1107 402 -1106
rect 513 -1107 514 -1106
rect 639 -1107 640 -1106
rect 982 -1107 983 -1106
rect 1003 -1107 1004 -1106
rect 1017 -1107 1018 -1106
rect 1094 -1107 1095 -1106
rect 1199 -1107 1200 -1106
rect 401 -1109 402 -1108
rect 450 -1109 451 -1108
rect 457 -1109 458 -1108
rect 639 -1109 640 -1108
rect 884 -1109 885 -1108
rect 1129 -1109 1130 -1108
rect 450 -1111 451 -1110
rect 646 -1111 647 -1110
rect 737 -1111 738 -1110
rect 884 -1111 885 -1110
rect 912 -1111 913 -1110
rect 1017 -1111 1018 -1110
rect 1031 -1111 1032 -1110
rect 1094 -1111 1095 -1110
rect 1101 -1111 1102 -1110
rect 1206 -1111 1207 -1110
rect 457 -1113 458 -1112
rect 520 -1113 521 -1112
rect 604 -1113 605 -1112
rect 912 -1113 913 -1112
rect 919 -1113 920 -1112
rect 1122 -1113 1123 -1112
rect 625 -1115 626 -1114
rect 646 -1115 647 -1114
rect 723 -1115 724 -1114
rect 1031 -1115 1032 -1114
rect 282 -1117 283 -1116
rect 723 -1117 724 -1116
rect 737 -1117 738 -1116
rect 761 -1117 762 -1116
rect 849 -1117 850 -1116
rect 1101 -1117 1102 -1116
rect 282 -1119 283 -1118
rect 590 -1119 591 -1118
rect 849 -1119 850 -1118
rect 1010 -1119 1011 -1118
rect 317 -1121 318 -1120
rect 625 -1121 626 -1120
rect 898 -1121 899 -1120
rect 919 -1121 920 -1120
rect 926 -1121 927 -1120
rect 1010 -1121 1011 -1120
rect 100 -1123 101 -1122
rect 317 -1123 318 -1122
rect 436 -1123 437 -1122
rect 898 -1123 899 -1122
rect 961 -1123 962 -1122
rect 1087 -1123 1088 -1122
rect 100 -1125 101 -1124
rect 303 -1125 304 -1124
rect 387 -1125 388 -1124
rect 436 -1125 437 -1124
rect 786 -1125 787 -1124
rect 926 -1125 927 -1124
rect 975 -1125 976 -1124
rect 1426 -1125 1427 -1124
rect 65 -1127 66 -1126
rect 303 -1127 304 -1126
rect 667 -1127 668 -1126
rect 786 -1127 787 -1126
rect 800 -1127 801 -1126
rect 961 -1127 962 -1126
rect 51 -1129 52 -1128
rect 65 -1129 66 -1128
rect 765 -1129 766 -1128
rect 800 -1129 801 -1128
rect 16 -1131 17 -1130
rect 765 -1131 766 -1130
rect 16 -1133 17 -1132
rect 289 -1133 290 -1132
rect 51 -1135 52 -1134
rect 506 -1135 507 -1134
rect 233 -1137 234 -1136
rect 289 -1137 290 -1136
rect 506 -1137 507 -1136
rect 677 -1137 678 -1136
rect 149 -1139 150 -1138
rect 233 -1139 234 -1138
rect 128 -1141 129 -1140
rect 149 -1141 150 -1140
rect 128 -1143 129 -1142
rect 618 -1143 619 -1142
rect 527 -1145 528 -1144
rect 618 -1145 619 -1144
rect 366 -1147 367 -1146
rect 527 -1147 528 -1146
rect 324 -1149 325 -1148
rect 366 -1149 367 -1148
rect 324 -1151 325 -1150
rect 387 -1151 388 -1150
rect 9 -1162 10 -1161
rect 303 -1162 304 -1161
rect 341 -1162 342 -1161
rect 345 -1162 346 -1161
rect 352 -1162 353 -1161
rect 667 -1162 668 -1161
rect 670 -1162 671 -1161
rect 800 -1162 801 -1161
rect 828 -1162 829 -1161
rect 1122 -1162 1123 -1161
rect 1248 -1162 1249 -1161
rect 1251 -1162 1252 -1161
rect 9 -1164 10 -1163
rect 607 -1164 608 -1163
rect 667 -1164 668 -1163
rect 772 -1164 773 -1163
rect 782 -1164 783 -1163
rect 807 -1164 808 -1163
rect 828 -1164 829 -1163
rect 863 -1164 864 -1163
rect 894 -1164 895 -1163
rect 1367 -1164 1368 -1163
rect 12 -1166 13 -1165
rect 44 -1166 45 -1165
rect 61 -1166 62 -1165
rect 597 -1166 598 -1165
rect 719 -1166 720 -1165
rect 1129 -1166 1130 -1165
rect 1248 -1166 1249 -1165
rect 1451 -1166 1452 -1165
rect 30 -1168 31 -1167
rect 702 -1168 703 -1167
rect 719 -1168 720 -1167
rect 1458 -1168 1459 -1167
rect 33 -1170 34 -1169
rect 289 -1170 290 -1169
rect 310 -1170 311 -1169
rect 345 -1170 346 -1169
rect 408 -1170 409 -1169
rect 954 -1170 955 -1169
rect 957 -1170 958 -1169
rect 1528 -1170 1529 -1169
rect 37 -1172 38 -1171
rect 723 -1172 724 -1171
rect 730 -1172 731 -1171
rect 1472 -1172 1473 -1171
rect 1528 -1172 1529 -1171
rect 1563 -1172 1564 -1171
rect 37 -1174 38 -1173
rect 758 -1174 759 -1173
rect 772 -1174 773 -1173
rect 933 -1174 934 -1173
rect 954 -1174 955 -1173
rect 982 -1174 983 -1173
rect 989 -1174 990 -1173
rect 992 -1174 993 -1173
rect 1055 -1174 1056 -1173
rect 1563 -1174 1564 -1173
rect 40 -1176 41 -1175
rect 583 -1176 584 -1175
rect 597 -1176 598 -1175
rect 639 -1176 640 -1175
rect 702 -1176 703 -1175
rect 1269 -1176 1270 -1175
rect 1367 -1176 1368 -1175
rect 1402 -1176 1403 -1175
rect 1451 -1176 1452 -1175
rect 1500 -1176 1501 -1175
rect 44 -1178 45 -1177
rect 93 -1178 94 -1177
rect 103 -1178 104 -1177
rect 422 -1178 423 -1177
rect 457 -1178 458 -1177
rect 618 -1178 619 -1177
rect 625 -1178 626 -1177
rect 982 -1178 983 -1177
rect 989 -1178 990 -1177
rect 1031 -1178 1032 -1177
rect 1122 -1178 1123 -1177
rect 1143 -1178 1144 -1177
rect 1171 -1178 1172 -1177
rect 1472 -1178 1473 -1177
rect 51 -1180 52 -1179
rect 457 -1180 458 -1179
rect 481 -1180 482 -1179
rect 1297 -1180 1298 -1179
rect 1381 -1180 1382 -1179
rect 1458 -1180 1459 -1179
rect 51 -1182 52 -1181
rect 177 -1182 178 -1181
rect 184 -1182 185 -1181
rect 733 -1182 734 -1181
rect 754 -1182 755 -1181
rect 1059 -1182 1060 -1181
rect 1143 -1182 1144 -1181
rect 1164 -1182 1165 -1181
rect 1251 -1182 1252 -1181
rect 1500 -1182 1501 -1181
rect 79 -1184 80 -1183
rect 100 -1184 101 -1183
rect 107 -1184 108 -1183
rect 593 -1184 594 -1183
rect 618 -1184 619 -1183
rect 751 -1184 752 -1183
rect 758 -1184 759 -1183
rect 821 -1184 822 -1183
rect 831 -1184 832 -1183
rect 1108 -1184 1109 -1183
rect 1164 -1184 1165 -1183
rect 1206 -1184 1207 -1183
rect 1297 -1184 1298 -1183
rect 1325 -1184 1326 -1183
rect 1381 -1184 1382 -1183
rect 1437 -1184 1438 -1183
rect 79 -1186 80 -1185
rect 387 -1186 388 -1185
rect 408 -1186 409 -1185
rect 485 -1186 486 -1185
rect 506 -1186 507 -1185
rect 859 -1186 860 -1185
rect 863 -1186 864 -1185
rect 877 -1186 878 -1185
rect 922 -1186 923 -1185
rect 1374 -1186 1375 -1185
rect 1402 -1186 1403 -1185
rect 1423 -1186 1424 -1185
rect 82 -1188 83 -1187
rect 464 -1188 465 -1187
rect 485 -1188 486 -1187
rect 562 -1188 563 -1187
rect 569 -1188 570 -1187
rect 821 -1188 822 -1187
rect 835 -1188 836 -1187
rect 936 -1188 937 -1187
rect 996 -1188 997 -1187
rect 1108 -1188 1109 -1187
rect 1192 -1188 1193 -1187
rect 1325 -1188 1326 -1187
rect 1374 -1188 1375 -1187
rect 1430 -1188 1431 -1187
rect 86 -1190 87 -1189
rect 107 -1190 108 -1189
rect 114 -1190 115 -1189
rect 506 -1190 507 -1189
rect 509 -1190 510 -1189
rect 870 -1190 871 -1189
rect 877 -1190 878 -1189
rect 905 -1190 906 -1189
rect 1059 -1190 1060 -1189
rect 1136 -1190 1137 -1189
rect 1192 -1190 1193 -1189
rect 1388 -1190 1389 -1189
rect 1430 -1190 1431 -1189
rect 1479 -1190 1480 -1189
rect 86 -1192 87 -1191
rect 198 -1192 199 -1191
rect 205 -1192 206 -1191
rect 303 -1192 304 -1191
rect 310 -1192 311 -1191
rect 663 -1192 664 -1191
rect 723 -1192 724 -1191
rect 1017 -1192 1018 -1191
rect 1136 -1192 1137 -1191
rect 1157 -1192 1158 -1191
rect 1206 -1192 1207 -1191
rect 1227 -1192 1228 -1191
rect 1262 -1192 1263 -1191
rect 1423 -1192 1424 -1191
rect 1479 -1192 1480 -1191
rect 1549 -1192 1550 -1191
rect 93 -1194 94 -1193
rect 716 -1194 717 -1193
rect 730 -1194 731 -1193
rect 1080 -1194 1081 -1193
rect 1157 -1194 1158 -1193
rect 1174 -1194 1175 -1193
rect 1227 -1194 1228 -1193
rect 1255 -1194 1256 -1193
rect 1262 -1194 1263 -1193
rect 1486 -1194 1487 -1193
rect 100 -1196 101 -1195
rect 996 -1196 997 -1195
rect 1080 -1196 1081 -1195
rect 1094 -1196 1095 -1195
rect 1255 -1196 1256 -1195
rect 1311 -1196 1312 -1195
rect 1360 -1196 1361 -1195
rect 1486 -1196 1487 -1195
rect 114 -1198 115 -1197
rect 478 -1198 479 -1197
rect 513 -1198 514 -1197
rect 604 -1198 605 -1197
rect 611 -1198 612 -1197
rect 870 -1198 871 -1197
rect 905 -1198 906 -1197
rect 919 -1198 920 -1197
rect 940 -1198 941 -1197
rect 1017 -1198 1018 -1197
rect 1311 -1198 1312 -1197
rect 1332 -1198 1333 -1197
rect 1360 -1198 1361 -1197
rect 1395 -1198 1396 -1197
rect 2 -1200 3 -1199
rect 478 -1200 479 -1199
rect 541 -1200 542 -1199
rect 625 -1200 626 -1199
rect 639 -1200 640 -1199
rect 646 -1200 647 -1199
rect 653 -1200 654 -1199
rect 1549 -1200 1550 -1199
rect 2 -1202 3 -1201
rect 975 -1202 976 -1201
rect 1003 -1202 1004 -1201
rect 1094 -1202 1095 -1201
rect 1220 -1202 1221 -1201
rect 1332 -1202 1333 -1201
rect 1388 -1202 1389 -1201
rect 1542 -1202 1543 -1201
rect 121 -1204 122 -1203
rect 530 -1204 531 -1203
rect 541 -1204 542 -1203
rect 555 -1204 556 -1203
rect 583 -1204 584 -1203
rect 765 -1204 766 -1203
rect 786 -1204 787 -1203
rect 807 -1204 808 -1203
rect 856 -1204 857 -1203
rect 1507 -1204 1508 -1203
rect 1542 -1204 1543 -1203
rect 1598 -1204 1599 -1203
rect 121 -1206 122 -1205
rect 268 -1206 269 -1205
rect 289 -1206 290 -1205
rect 338 -1206 339 -1205
rect 366 -1206 367 -1205
rect 387 -1206 388 -1205
rect 394 -1206 395 -1205
rect 716 -1206 717 -1205
rect 751 -1206 752 -1205
rect 1129 -1206 1130 -1205
rect 1395 -1206 1396 -1205
rect 1444 -1206 1445 -1205
rect 1507 -1206 1508 -1205
rect 1570 -1206 1571 -1205
rect 131 -1208 132 -1207
rect 919 -1208 920 -1207
rect 936 -1208 937 -1207
rect 1220 -1208 1221 -1207
rect 1276 -1208 1277 -1207
rect 1444 -1208 1445 -1207
rect 166 -1210 167 -1209
rect 898 -1210 899 -1209
rect 940 -1210 941 -1209
rect 961 -1210 962 -1209
rect 975 -1210 976 -1209
rect 1073 -1210 1074 -1209
rect 1150 -1210 1151 -1209
rect 1276 -1210 1277 -1209
rect 177 -1212 178 -1211
rect 247 -1212 248 -1211
rect 254 -1212 255 -1211
rect 933 -1212 934 -1211
rect 961 -1212 962 -1211
rect 1045 -1212 1046 -1211
rect 1150 -1212 1151 -1211
rect 1178 -1212 1179 -1211
rect 16 -1214 17 -1213
rect 247 -1214 248 -1213
rect 261 -1214 262 -1213
rect 268 -1214 269 -1213
rect 362 -1214 363 -1213
rect 1045 -1214 1046 -1213
rect 1178 -1214 1179 -1213
rect 1318 -1214 1319 -1213
rect 16 -1216 17 -1215
rect 275 -1216 276 -1215
rect 366 -1216 367 -1215
rect 373 -1216 374 -1215
rect 394 -1216 395 -1215
rect 415 -1216 416 -1215
rect 422 -1216 423 -1215
rect 460 -1216 461 -1215
rect 520 -1216 521 -1215
rect 646 -1216 647 -1215
rect 653 -1216 654 -1215
rect 737 -1216 738 -1215
rect 765 -1216 766 -1215
rect 1115 -1216 1116 -1215
rect 1318 -1216 1319 -1215
rect 1346 -1216 1347 -1215
rect 65 -1218 66 -1217
rect 254 -1218 255 -1217
rect 275 -1218 276 -1217
rect 429 -1218 430 -1217
rect 436 -1218 437 -1217
rect 464 -1218 465 -1217
rect 520 -1218 521 -1217
rect 1535 -1218 1536 -1217
rect 65 -1220 66 -1219
rect 527 -1220 528 -1219
rect 548 -1220 549 -1219
rect 562 -1220 563 -1219
rect 590 -1220 591 -1219
rect 1346 -1220 1347 -1219
rect 1535 -1220 1536 -1219
rect 1584 -1220 1585 -1219
rect 170 -1222 171 -1221
rect 261 -1222 262 -1221
rect 317 -1222 318 -1221
rect 436 -1222 437 -1221
rect 527 -1222 528 -1221
rect 1269 -1222 1270 -1221
rect 170 -1224 171 -1223
rect 352 -1224 353 -1223
rect 373 -1224 374 -1223
rect 499 -1224 500 -1223
rect 548 -1224 549 -1223
rect 611 -1224 612 -1223
rect 628 -1224 629 -1223
rect 1003 -1224 1004 -1223
rect 184 -1226 185 -1225
rect 558 -1226 559 -1225
rect 590 -1226 591 -1225
rect 681 -1226 682 -1225
rect 744 -1226 745 -1225
rect 1115 -1226 1116 -1225
rect 191 -1228 192 -1227
rect 205 -1228 206 -1227
rect 212 -1228 213 -1227
rect 446 -1228 447 -1227
rect 555 -1228 556 -1227
rect 1591 -1228 1592 -1227
rect 191 -1230 192 -1229
rect 233 -1230 234 -1229
rect 240 -1230 241 -1229
rect 415 -1230 416 -1229
rect 429 -1230 430 -1229
rect 471 -1230 472 -1229
rect 604 -1230 605 -1229
rect 1283 -1230 1284 -1229
rect 58 -1232 59 -1231
rect 240 -1232 241 -1231
rect 338 -1232 339 -1231
rect 744 -1232 745 -1231
rect 786 -1232 787 -1231
rect 842 -1232 843 -1231
rect 859 -1232 860 -1231
rect 1353 -1232 1354 -1231
rect 149 -1234 150 -1233
rect 233 -1234 234 -1233
rect 380 -1234 381 -1233
rect 499 -1234 500 -1233
rect 681 -1234 682 -1233
rect 688 -1234 689 -1233
rect 796 -1234 797 -1233
rect 1010 -1234 1011 -1233
rect 1199 -1234 1200 -1233
rect 1283 -1234 1284 -1233
rect 1353 -1234 1354 -1233
rect 1493 -1234 1494 -1233
rect 128 -1236 129 -1235
rect 688 -1236 689 -1235
rect 768 -1236 769 -1235
rect 1199 -1236 1200 -1235
rect 1409 -1236 1410 -1235
rect 1493 -1236 1494 -1235
rect 149 -1238 150 -1237
rect 660 -1238 661 -1237
rect 800 -1238 801 -1237
rect 849 -1238 850 -1237
rect 898 -1238 899 -1237
rect 947 -1238 948 -1237
rect 1010 -1238 1011 -1237
rect 1066 -1238 1067 -1237
rect 1409 -1238 1410 -1237
rect 1416 -1238 1417 -1237
rect 198 -1240 199 -1239
rect 317 -1240 318 -1239
rect 401 -1240 402 -1239
rect 569 -1240 570 -1239
rect 660 -1240 661 -1239
rect 726 -1240 727 -1239
rect 814 -1240 815 -1239
rect 856 -1240 857 -1239
rect 947 -1240 948 -1239
rect 968 -1240 969 -1239
rect 1066 -1240 1067 -1239
rect 1087 -1240 1088 -1239
rect 1416 -1240 1417 -1239
rect 1465 -1240 1466 -1239
rect 212 -1242 213 -1241
rect 359 -1242 360 -1241
rect 401 -1242 402 -1241
rect 576 -1242 577 -1241
rect 632 -1242 633 -1241
rect 814 -1242 815 -1241
rect 838 -1242 839 -1241
rect 1073 -1242 1074 -1241
rect 1087 -1242 1088 -1241
rect 1101 -1242 1102 -1241
rect 1465 -1242 1466 -1241
rect 1514 -1242 1515 -1241
rect 219 -1244 220 -1243
rect 513 -1244 514 -1243
rect 576 -1244 577 -1243
rect 926 -1244 927 -1243
rect 968 -1244 969 -1243
rect 1024 -1244 1025 -1243
rect 1514 -1244 1515 -1243
rect 1577 -1244 1578 -1243
rect 142 -1246 143 -1245
rect 219 -1246 220 -1245
rect 226 -1246 227 -1245
rect 390 -1246 391 -1245
rect 450 -1246 451 -1245
rect 842 -1246 843 -1245
rect 849 -1246 850 -1245
rect 884 -1246 885 -1245
rect 912 -1246 913 -1245
rect 1101 -1246 1102 -1245
rect 58 -1248 59 -1247
rect 884 -1248 885 -1247
rect 926 -1248 927 -1247
rect 1052 -1248 1053 -1247
rect 128 -1250 129 -1249
rect 142 -1250 143 -1249
rect 226 -1250 227 -1249
rect 324 -1250 325 -1249
rect 450 -1250 451 -1249
rect 534 -1250 535 -1249
rect 632 -1250 633 -1249
rect 695 -1250 696 -1249
rect 737 -1250 738 -1249
rect 1052 -1250 1053 -1249
rect 296 -1252 297 -1251
rect 380 -1252 381 -1251
rect 471 -1252 472 -1251
rect 709 -1252 710 -1251
rect 779 -1252 780 -1251
rect 912 -1252 913 -1251
rect 1024 -1252 1025 -1251
rect 1038 -1252 1039 -1251
rect 163 -1254 164 -1253
rect 709 -1254 710 -1253
rect 779 -1254 780 -1253
rect 1437 -1254 1438 -1253
rect 156 -1256 157 -1255
rect 163 -1256 164 -1255
rect 296 -1256 297 -1255
rect 492 -1256 493 -1255
rect 534 -1256 535 -1255
rect 793 -1256 794 -1255
rect 1038 -1256 1039 -1255
rect 1185 -1256 1186 -1255
rect 135 -1258 136 -1257
rect 156 -1258 157 -1257
rect 173 -1258 174 -1257
rect 793 -1258 794 -1257
rect 1185 -1258 1186 -1257
rect 1213 -1258 1214 -1257
rect 135 -1260 136 -1259
rect 359 -1260 360 -1259
rect 492 -1260 493 -1259
rect 835 -1260 836 -1259
rect 1213 -1260 1214 -1259
rect 1234 -1260 1235 -1259
rect 320 -1262 321 -1261
rect 695 -1262 696 -1261
rect 1234 -1262 1235 -1261
rect 1241 -1262 1242 -1261
rect 324 -1264 325 -1263
rect 331 -1264 332 -1263
rect 1241 -1264 1242 -1263
rect 1290 -1264 1291 -1263
rect 331 -1266 332 -1265
rect 443 -1266 444 -1265
rect 1290 -1266 1291 -1265
rect 1304 -1266 1305 -1265
rect 443 -1268 444 -1267
rect 754 -1268 755 -1267
rect 1304 -1268 1305 -1267
rect 1339 -1268 1340 -1267
rect 1339 -1270 1340 -1269
rect 1521 -1270 1522 -1269
rect 1521 -1272 1522 -1271
rect 1556 -1272 1557 -1271
rect 891 -1274 892 -1273
rect 1556 -1274 1557 -1273
rect 355 -1276 356 -1275
rect 891 -1276 892 -1275
rect 2 -1287 3 -1286
rect 555 -1287 556 -1286
rect 562 -1287 563 -1286
rect 604 -1287 605 -1286
rect 649 -1287 650 -1286
rect 1486 -1287 1487 -1286
rect 2 -1289 3 -1288
rect 373 -1289 374 -1288
rect 478 -1289 479 -1288
rect 1290 -1289 1291 -1288
rect 1451 -1289 1452 -1288
rect 1454 -1289 1455 -1288
rect 1486 -1289 1487 -1288
rect 1514 -1289 1515 -1288
rect 30 -1291 31 -1290
rect 754 -1291 755 -1290
rect 765 -1291 766 -1290
rect 1346 -1291 1347 -1290
rect 1451 -1291 1452 -1290
rect 1465 -1291 1466 -1290
rect 1514 -1291 1515 -1290
rect 1542 -1291 1543 -1290
rect 30 -1293 31 -1292
rect 44 -1293 45 -1292
rect 61 -1293 62 -1292
rect 1472 -1293 1473 -1292
rect 37 -1295 38 -1294
rect 520 -1295 521 -1294
rect 527 -1295 528 -1294
rect 541 -1295 542 -1294
rect 548 -1295 549 -1294
rect 1549 -1295 1550 -1294
rect 37 -1297 38 -1296
rect 443 -1297 444 -1296
rect 488 -1297 489 -1296
rect 499 -1297 500 -1296
rect 509 -1297 510 -1296
rect 982 -1297 983 -1296
rect 1052 -1297 1053 -1296
rect 1458 -1297 1459 -1296
rect 1472 -1297 1473 -1296
rect 1479 -1297 1480 -1296
rect 44 -1299 45 -1298
rect 240 -1299 241 -1298
rect 338 -1299 339 -1298
rect 408 -1299 409 -1298
rect 422 -1299 423 -1298
rect 443 -1299 444 -1298
rect 467 -1299 468 -1298
rect 499 -1299 500 -1298
rect 548 -1299 549 -1298
rect 779 -1299 780 -1298
rect 782 -1299 783 -1298
rect 1521 -1299 1522 -1298
rect 68 -1301 69 -1300
rect 814 -1301 815 -1300
rect 835 -1301 836 -1300
rect 1234 -1301 1235 -1300
rect 1346 -1301 1347 -1300
rect 1367 -1301 1368 -1300
rect 1388 -1301 1389 -1300
rect 1458 -1301 1459 -1300
rect 1479 -1301 1480 -1300
rect 1507 -1301 1508 -1300
rect 100 -1303 101 -1302
rect 429 -1303 430 -1302
rect 555 -1303 556 -1302
rect 674 -1303 675 -1302
rect 719 -1303 720 -1302
rect 1521 -1303 1522 -1302
rect 100 -1305 101 -1304
rect 149 -1305 150 -1304
rect 177 -1305 178 -1304
rect 320 -1305 321 -1304
rect 345 -1305 346 -1304
rect 373 -1305 374 -1304
rect 387 -1305 388 -1304
rect 429 -1305 430 -1304
rect 562 -1305 563 -1304
rect 786 -1305 787 -1304
rect 793 -1305 794 -1304
rect 1006 -1305 1007 -1304
rect 1055 -1305 1056 -1304
rect 1528 -1305 1529 -1304
rect 79 -1307 80 -1306
rect 387 -1307 388 -1306
rect 401 -1307 402 -1306
rect 541 -1307 542 -1306
rect 674 -1307 675 -1306
rect 681 -1307 682 -1306
rect 723 -1307 724 -1306
rect 1031 -1307 1032 -1306
rect 1171 -1307 1172 -1306
rect 1402 -1307 1403 -1306
rect 1454 -1307 1455 -1306
rect 1465 -1307 1466 -1306
rect 1507 -1307 1508 -1306
rect 1535 -1307 1536 -1306
rect 79 -1309 80 -1308
rect 198 -1309 199 -1308
rect 233 -1309 234 -1308
rect 359 -1309 360 -1308
rect 418 -1309 419 -1308
rect 1367 -1309 1368 -1308
rect 1388 -1309 1389 -1308
rect 1430 -1309 1431 -1308
rect 1528 -1309 1529 -1308
rect 1556 -1309 1557 -1308
rect 82 -1311 83 -1310
rect 177 -1311 178 -1310
rect 198 -1311 199 -1310
rect 530 -1311 531 -1310
rect 632 -1311 633 -1310
rect 681 -1311 682 -1310
rect 723 -1311 724 -1310
rect 768 -1311 769 -1310
rect 779 -1311 780 -1310
rect 828 -1311 829 -1310
rect 835 -1311 836 -1310
rect 842 -1311 843 -1310
rect 880 -1311 881 -1310
rect 1500 -1311 1501 -1310
rect 86 -1313 87 -1312
rect 320 -1313 321 -1312
rect 345 -1313 346 -1312
rect 362 -1313 363 -1312
rect 422 -1313 423 -1312
rect 450 -1313 451 -1312
rect 481 -1313 482 -1312
rect 793 -1313 794 -1312
rect 828 -1313 829 -1312
rect 856 -1313 857 -1312
rect 922 -1313 923 -1312
rect 1444 -1313 1445 -1312
rect 86 -1315 87 -1314
rect 415 -1315 416 -1314
rect 450 -1315 451 -1314
rect 485 -1315 486 -1314
rect 604 -1315 605 -1314
rect 922 -1315 923 -1314
rect 933 -1315 934 -1314
rect 1493 -1315 1494 -1314
rect 9 -1317 10 -1316
rect 485 -1317 486 -1316
rect 737 -1317 738 -1316
rect 873 -1317 874 -1316
rect 933 -1317 934 -1316
rect 954 -1317 955 -1316
rect 975 -1317 976 -1316
rect 1052 -1317 1053 -1316
rect 1101 -1317 1102 -1316
rect 1535 -1317 1536 -1316
rect 9 -1319 10 -1318
rect 65 -1319 66 -1318
rect 93 -1319 94 -1318
rect 149 -1319 150 -1318
rect 212 -1319 213 -1318
rect 481 -1319 482 -1318
rect 667 -1319 668 -1318
rect 737 -1319 738 -1318
rect 744 -1319 745 -1318
rect 814 -1319 815 -1318
rect 838 -1319 839 -1318
rect 863 -1319 864 -1318
rect 898 -1319 899 -1318
rect 954 -1319 955 -1318
rect 982 -1319 983 -1318
rect 996 -1319 997 -1318
rect 1024 -1319 1025 -1318
rect 1031 -1319 1032 -1318
rect 1101 -1319 1102 -1318
rect 1213 -1319 1214 -1318
rect 1234 -1319 1235 -1318
rect 1262 -1319 1263 -1318
rect 1339 -1319 1340 -1318
rect 1493 -1319 1494 -1318
rect 93 -1321 94 -1320
rect 569 -1321 570 -1320
rect 618 -1321 619 -1320
rect 667 -1321 668 -1320
rect 688 -1321 689 -1320
rect 744 -1321 745 -1320
rect 751 -1321 752 -1320
rect 1311 -1321 1312 -1320
rect 1353 -1321 1354 -1320
rect 1430 -1321 1431 -1320
rect 103 -1323 104 -1322
rect 1423 -1323 1424 -1322
rect 110 -1325 111 -1324
rect 296 -1325 297 -1324
rect 303 -1325 304 -1324
rect 751 -1325 752 -1324
rect 765 -1325 766 -1324
rect 800 -1325 801 -1324
rect 849 -1325 850 -1324
rect 898 -1325 899 -1324
rect 961 -1325 962 -1324
rect 1024 -1325 1025 -1324
rect 1038 -1325 1039 -1324
rect 1213 -1325 1214 -1324
rect 1255 -1325 1256 -1324
rect 1500 -1325 1501 -1324
rect 128 -1327 129 -1326
rect 859 -1327 860 -1326
rect 863 -1327 864 -1326
rect 926 -1327 927 -1326
rect 940 -1327 941 -1326
rect 961 -1327 962 -1326
rect 996 -1327 997 -1326
rect 1003 -1327 1004 -1326
rect 1010 -1327 1011 -1326
rect 1038 -1327 1039 -1326
rect 1087 -1327 1088 -1326
rect 1339 -1327 1340 -1326
rect 1395 -1327 1396 -1326
rect 1402 -1327 1403 -1326
rect 1416 -1327 1417 -1326
rect 1423 -1327 1424 -1326
rect 107 -1329 108 -1328
rect 128 -1329 129 -1328
rect 131 -1329 132 -1328
rect 702 -1329 703 -1328
rect 712 -1329 713 -1328
rect 1262 -1329 1263 -1328
rect 1311 -1329 1312 -1328
rect 1360 -1329 1361 -1328
rect 1395 -1329 1396 -1328
rect 1437 -1329 1438 -1328
rect 107 -1331 108 -1330
rect 114 -1331 115 -1330
rect 215 -1331 216 -1330
rect 296 -1331 297 -1330
rect 303 -1331 304 -1330
rect 324 -1331 325 -1330
rect 352 -1331 353 -1330
rect 527 -1331 528 -1330
rect 618 -1331 619 -1330
rect 639 -1331 640 -1330
rect 730 -1331 731 -1330
rect 1087 -1331 1088 -1330
rect 1143 -1331 1144 -1330
rect 1171 -1331 1172 -1330
rect 1178 -1331 1179 -1330
rect 1290 -1331 1291 -1330
rect 1332 -1331 1333 -1330
rect 1437 -1331 1438 -1330
rect 16 -1333 17 -1332
rect 352 -1333 353 -1332
rect 436 -1333 437 -1332
rect 569 -1333 570 -1332
rect 639 -1333 640 -1332
rect 912 -1333 913 -1332
rect 926 -1333 927 -1332
rect 989 -1333 990 -1332
rect 1059 -1333 1060 -1332
rect 1143 -1333 1144 -1332
rect 1157 -1333 1158 -1332
rect 1444 -1333 1445 -1332
rect 16 -1335 17 -1334
rect 205 -1335 206 -1334
rect 233 -1335 234 -1334
rect 310 -1335 311 -1334
rect 436 -1335 437 -1334
rect 464 -1335 465 -1334
rect 471 -1335 472 -1334
rect 688 -1335 689 -1334
rect 786 -1335 787 -1334
rect 870 -1335 871 -1334
rect 940 -1335 941 -1334
rect 978 -1335 979 -1334
rect 989 -1335 990 -1334
rect 1150 -1335 1151 -1334
rect 1164 -1335 1165 -1334
rect 1178 -1335 1179 -1334
rect 1192 -1335 1193 -1334
rect 1353 -1335 1354 -1334
rect 1360 -1335 1361 -1334
rect 1374 -1335 1375 -1334
rect 51 -1337 52 -1336
rect 114 -1337 115 -1336
rect 170 -1337 171 -1336
rect 324 -1337 325 -1336
rect 457 -1337 458 -1336
rect 702 -1337 703 -1336
rect 800 -1337 801 -1336
rect 807 -1337 808 -1336
rect 842 -1337 843 -1336
rect 849 -1337 850 -1336
rect 856 -1337 857 -1336
rect 877 -1337 878 -1336
rect 947 -1337 948 -1336
rect 1010 -1337 1011 -1336
rect 1122 -1337 1123 -1336
rect 1157 -1337 1158 -1336
rect 1255 -1337 1256 -1336
rect 1276 -1337 1277 -1336
rect 1374 -1337 1375 -1336
rect 1381 -1337 1382 -1336
rect 51 -1339 52 -1338
rect 261 -1339 262 -1338
rect 275 -1339 276 -1338
rect 310 -1339 311 -1338
rect 317 -1339 318 -1338
rect 807 -1339 808 -1338
rect 877 -1339 878 -1338
rect 891 -1339 892 -1338
rect 905 -1339 906 -1338
rect 947 -1339 948 -1338
rect 1003 -1339 1004 -1338
rect 1059 -1339 1060 -1338
rect 1122 -1339 1123 -1338
rect 1227 -1339 1228 -1338
rect 1248 -1339 1249 -1338
rect 1381 -1339 1382 -1338
rect 65 -1341 66 -1340
rect 912 -1341 913 -1340
rect 1080 -1341 1081 -1340
rect 1248 -1341 1249 -1340
rect 1269 -1341 1270 -1340
rect 1276 -1341 1277 -1340
rect 142 -1343 143 -1342
rect 170 -1343 171 -1342
rect 184 -1343 185 -1342
rect 275 -1343 276 -1342
rect 317 -1343 318 -1342
rect 632 -1343 633 -1342
rect 695 -1343 696 -1342
rect 1269 -1343 1270 -1342
rect 58 -1345 59 -1344
rect 695 -1345 696 -1344
rect 884 -1345 885 -1344
rect 905 -1345 906 -1344
rect 1073 -1345 1074 -1344
rect 1080 -1345 1081 -1344
rect 1129 -1345 1130 -1344
rect 1332 -1345 1333 -1344
rect 58 -1347 59 -1346
rect 625 -1347 626 -1346
rect 884 -1347 885 -1346
rect 968 -1347 969 -1346
rect 1066 -1347 1067 -1346
rect 1073 -1347 1074 -1346
rect 1136 -1347 1137 -1346
rect 1164 -1347 1165 -1346
rect 1227 -1347 1228 -1346
rect 1318 -1347 1319 -1346
rect 135 -1349 136 -1348
rect 1129 -1349 1130 -1348
rect 1136 -1349 1137 -1348
rect 1199 -1349 1200 -1348
rect 1297 -1349 1298 -1348
rect 1318 -1349 1319 -1348
rect 72 -1351 73 -1350
rect 135 -1351 136 -1350
rect 142 -1351 143 -1350
rect 289 -1351 290 -1350
rect 457 -1351 458 -1350
rect 492 -1351 493 -1350
rect 495 -1351 496 -1350
rect 870 -1351 871 -1350
rect 891 -1351 892 -1350
rect 919 -1351 920 -1350
rect 1045 -1351 1046 -1350
rect 1066 -1351 1067 -1350
rect 1150 -1351 1151 -1350
rect 1185 -1351 1186 -1350
rect 1199 -1351 1200 -1350
rect 1206 -1351 1207 -1350
rect 1297 -1351 1298 -1350
rect 1325 -1351 1326 -1350
rect 72 -1353 73 -1352
rect 219 -1353 220 -1352
rect 226 -1353 227 -1352
rect 471 -1353 472 -1352
rect 478 -1353 479 -1352
rect 730 -1353 731 -1352
rect 1108 -1353 1109 -1352
rect 1206 -1353 1207 -1352
rect 1304 -1353 1305 -1352
rect 1325 -1353 1326 -1352
rect 121 -1355 122 -1354
rect 289 -1355 290 -1354
rect 464 -1355 465 -1354
rect 597 -1355 598 -1354
rect 625 -1355 626 -1354
rect 660 -1355 661 -1354
rect 709 -1355 710 -1354
rect 1108 -1355 1109 -1354
rect 1185 -1355 1186 -1354
rect 1563 -1355 1564 -1354
rect 121 -1357 122 -1356
rect 331 -1357 332 -1356
rect 492 -1357 493 -1356
rect 520 -1357 521 -1356
rect 523 -1357 524 -1356
rect 1045 -1357 1046 -1356
rect 163 -1359 164 -1358
rect 184 -1359 185 -1358
rect 205 -1359 206 -1358
rect 558 -1359 559 -1358
rect 597 -1359 598 -1358
rect 950 -1359 951 -1358
rect 1017 -1359 1018 -1358
rect 1304 -1359 1305 -1358
rect 163 -1361 164 -1360
rect 404 -1361 405 -1360
rect 506 -1361 507 -1360
rect 1416 -1361 1417 -1360
rect 219 -1363 220 -1362
rect 534 -1363 535 -1362
rect 611 -1363 612 -1362
rect 660 -1363 661 -1362
rect 709 -1363 710 -1362
rect 1115 -1363 1116 -1362
rect 226 -1365 227 -1364
rect 716 -1365 717 -1364
rect 845 -1365 846 -1364
rect 1115 -1365 1116 -1364
rect 240 -1367 241 -1366
rect 380 -1367 381 -1366
rect 390 -1367 391 -1366
rect 534 -1367 535 -1366
rect 551 -1367 552 -1366
rect 716 -1367 717 -1366
rect 247 -1369 248 -1368
rect 408 -1369 409 -1368
rect 506 -1369 507 -1368
rect 975 -1369 976 -1368
rect 247 -1371 248 -1370
rect 583 -1371 584 -1370
rect 590 -1371 591 -1370
rect 611 -1371 612 -1370
rect 254 -1373 255 -1372
rect 359 -1373 360 -1372
rect 380 -1373 381 -1372
rect 394 -1373 395 -1372
rect 513 -1373 514 -1372
rect 583 -1373 584 -1372
rect 590 -1373 591 -1372
rect 726 -1373 727 -1372
rect 212 -1375 213 -1374
rect 254 -1375 255 -1374
rect 261 -1375 262 -1374
rect 607 -1375 608 -1374
rect 331 -1377 332 -1376
rect 1017 -1377 1018 -1376
rect 394 -1379 395 -1378
rect 653 -1379 654 -1378
rect 513 -1381 514 -1380
rect 1283 -1381 1284 -1380
rect 516 -1383 517 -1382
rect 1283 -1383 1284 -1382
rect 523 -1385 524 -1384
rect 1192 -1385 1193 -1384
rect 576 -1387 577 -1386
rect 653 -1387 654 -1386
rect 576 -1389 577 -1388
rect 821 -1389 822 -1388
rect 758 -1391 759 -1390
rect 821 -1391 822 -1390
rect 646 -1393 647 -1392
rect 758 -1393 759 -1392
rect 646 -1395 647 -1394
rect 968 -1395 969 -1394
rect 44 -1406 45 -1405
rect 649 -1406 650 -1405
rect 684 -1406 685 -1405
rect 730 -1406 731 -1405
rect 800 -1406 801 -1405
rect 838 -1406 839 -1405
rect 842 -1406 843 -1405
rect 1353 -1406 1354 -1405
rect 44 -1408 45 -1407
rect 114 -1408 115 -1407
rect 121 -1408 122 -1407
rect 467 -1408 468 -1407
rect 471 -1408 472 -1407
rect 495 -1408 496 -1407
rect 520 -1408 521 -1407
rect 527 -1408 528 -1407
rect 646 -1408 647 -1407
rect 1269 -1408 1270 -1407
rect 1353 -1408 1354 -1407
rect 1360 -1408 1361 -1407
rect 51 -1410 52 -1409
rect 418 -1410 419 -1409
rect 478 -1410 479 -1409
rect 1192 -1410 1193 -1409
rect 1311 -1410 1312 -1409
rect 1360 -1410 1361 -1409
rect 51 -1412 52 -1411
rect 317 -1412 318 -1411
rect 320 -1412 321 -1411
rect 408 -1412 409 -1411
rect 478 -1412 479 -1411
rect 1143 -1412 1144 -1411
rect 1192 -1412 1193 -1411
rect 1297 -1412 1298 -1411
rect 65 -1414 66 -1413
rect 296 -1414 297 -1413
rect 366 -1414 367 -1413
rect 397 -1414 398 -1413
rect 408 -1414 409 -1413
rect 492 -1414 493 -1413
rect 499 -1414 500 -1413
rect 520 -1414 521 -1413
rect 646 -1414 647 -1413
rect 1115 -1414 1116 -1413
rect 1276 -1414 1277 -1413
rect 1311 -1414 1312 -1413
rect 65 -1416 66 -1415
rect 569 -1416 570 -1415
rect 712 -1416 713 -1415
rect 779 -1416 780 -1415
rect 800 -1416 801 -1415
rect 1304 -1416 1305 -1415
rect 82 -1418 83 -1417
rect 275 -1418 276 -1417
rect 296 -1418 297 -1417
rect 338 -1418 339 -1417
rect 390 -1418 391 -1417
rect 523 -1418 524 -1417
rect 562 -1418 563 -1417
rect 779 -1418 780 -1417
rect 807 -1418 808 -1417
rect 1269 -1418 1270 -1417
rect 68 -1420 69 -1419
rect 338 -1420 339 -1419
rect 394 -1420 395 -1419
rect 831 -1420 832 -1419
rect 842 -1420 843 -1419
rect 856 -1420 857 -1419
rect 873 -1420 874 -1419
rect 1234 -1420 1235 -1419
rect 1262 -1420 1263 -1419
rect 1276 -1420 1277 -1419
rect 82 -1422 83 -1421
rect 121 -1422 122 -1421
rect 184 -1422 185 -1421
rect 513 -1422 514 -1421
rect 562 -1422 563 -1421
rect 660 -1422 661 -1421
rect 723 -1422 724 -1421
rect 726 -1422 727 -1421
rect 730 -1422 731 -1421
rect 835 -1422 836 -1421
rect 856 -1422 857 -1421
rect 1206 -1422 1207 -1421
rect 1234 -1422 1235 -1421
rect 1521 -1422 1522 -1421
rect 93 -1424 94 -1423
rect 492 -1424 493 -1423
rect 513 -1424 514 -1423
rect 541 -1424 542 -1423
rect 569 -1424 570 -1423
rect 992 -1424 993 -1423
rect 1003 -1424 1004 -1423
rect 1045 -1424 1046 -1423
rect 1076 -1424 1077 -1423
rect 1318 -1424 1319 -1423
rect 1332 -1424 1333 -1423
rect 1521 -1424 1522 -1423
rect 37 -1426 38 -1425
rect 93 -1426 94 -1425
rect 100 -1426 101 -1425
rect 404 -1426 405 -1425
rect 464 -1426 465 -1425
rect 1143 -1426 1144 -1425
rect 1164 -1426 1165 -1425
rect 1262 -1426 1263 -1425
rect 37 -1428 38 -1427
rect 835 -1428 836 -1427
rect 880 -1428 881 -1427
rect 933 -1428 934 -1427
rect 950 -1428 951 -1427
rect 1465 -1428 1466 -1427
rect 100 -1430 101 -1429
rect 254 -1430 255 -1429
rect 275 -1430 276 -1429
rect 688 -1430 689 -1429
rect 723 -1430 724 -1429
rect 1213 -1430 1214 -1429
rect 1444 -1430 1445 -1429
rect 1465 -1430 1466 -1429
rect 103 -1432 104 -1431
rect 432 -1432 433 -1431
rect 436 -1432 437 -1431
rect 464 -1432 465 -1431
rect 481 -1432 482 -1431
rect 1297 -1432 1298 -1431
rect 1416 -1432 1417 -1431
rect 1444 -1432 1445 -1431
rect 114 -1434 115 -1433
rect 261 -1434 262 -1433
rect 324 -1434 325 -1433
rect 366 -1434 367 -1433
rect 436 -1434 437 -1433
rect 632 -1434 633 -1433
rect 660 -1434 661 -1433
rect 744 -1434 745 -1433
rect 768 -1434 769 -1433
rect 807 -1434 808 -1433
rect 880 -1434 881 -1433
rect 1325 -1434 1326 -1433
rect 1381 -1434 1382 -1433
rect 1416 -1434 1417 -1433
rect 135 -1436 136 -1435
rect 254 -1436 255 -1435
rect 261 -1436 262 -1435
rect 359 -1436 360 -1435
rect 541 -1436 542 -1435
rect 849 -1436 850 -1435
rect 884 -1436 885 -1435
rect 887 -1436 888 -1435
rect 919 -1436 920 -1435
rect 1507 -1436 1508 -1435
rect 79 -1438 80 -1437
rect 1507 -1438 1508 -1437
rect 135 -1440 136 -1439
rect 173 -1440 174 -1439
rect 184 -1440 185 -1439
rect 191 -1440 192 -1439
rect 205 -1440 206 -1439
rect 527 -1440 528 -1439
rect 555 -1440 556 -1439
rect 1164 -1440 1165 -1439
rect 1178 -1440 1179 -1439
rect 1332 -1440 1333 -1439
rect 1381 -1440 1382 -1439
rect 1409 -1440 1410 -1439
rect 72 -1442 73 -1441
rect 205 -1442 206 -1441
rect 219 -1442 220 -1441
rect 600 -1442 601 -1441
rect 688 -1442 689 -1441
rect 695 -1442 696 -1441
rect 744 -1442 745 -1441
rect 772 -1442 773 -1441
rect 803 -1442 804 -1441
rect 1045 -1442 1046 -1441
rect 1080 -1442 1081 -1441
rect 1206 -1442 1207 -1441
rect 1213 -1442 1214 -1441
rect 1220 -1442 1221 -1441
rect 1409 -1442 1410 -1441
rect 1458 -1442 1459 -1441
rect 72 -1444 73 -1443
rect 653 -1444 654 -1443
rect 772 -1444 773 -1443
rect 898 -1444 899 -1443
rect 905 -1444 906 -1443
rect 1080 -1444 1081 -1443
rect 1129 -1444 1130 -1443
rect 1325 -1444 1326 -1443
rect 191 -1446 192 -1445
rect 583 -1446 584 -1445
rect 653 -1446 654 -1445
rect 674 -1446 675 -1445
rect 849 -1446 850 -1445
rect 1038 -1446 1039 -1445
rect 1129 -1446 1130 -1445
rect 1255 -1446 1256 -1445
rect 219 -1448 220 -1447
rect 516 -1448 517 -1447
rect 583 -1448 584 -1447
rect 618 -1448 619 -1447
rect 859 -1448 860 -1447
rect 1458 -1448 1459 -1447
rect 233 -1450 234 -1449
rect 317 -1450 318 -1449
rect 324 -1450 325 -1449
rect 548 -1450 549 -1449
rect 884 -1450 885 -1449
rect 961 -1450 962 -1449
rect 975 -1450 976 -1449
rect 1514 -1450 1515 -1449
rect 177 -1452 178 -1451
rect 233 -1452 234 -1451
rect 240 -1452 241 -1451
rect 677 -1452 678 -1451
rect 887 -1452 888 -1451
rect 961 -1452 962 -1451
rect 978 -1452 979 -1451
rect 1248 -1452 1249 -1451
rect 1514 -1452 1515 -1451
rect 1524 -1452 1525 -1451
rect 177 -1454 178 -1453
rect 590 -1454 591 -1453
rect 674 -1454 675 -1453
rect 1248 -1454 1249 -1453
rect 1437 -1454 1438 -1453
rect 1524 -1454 1525 -1453
rect 198 -1456 199 -1455
rect 548 -1456 549 -1455
rect 898 -1456 899 -1455
rect 954 -1456 955 -1455
rect 1006 -1456 1007 -1455
rect 1423 -1456 1424 -1455
rect 16 -1458 17 -1457
rect 198 -1458 199 -1457
rect 226 -1458 227 -1457
rect 590 -1458 591 -1457
rect 905 -1458 906 -1457
rect 940 -1458 941 -1457
rect 947 -1458 948 -1457
rect 1255 -1458 1256 -1457
rect 1388 -1458 1389 -1457
rect 1423 -1458 1424 -1457
rect 16 -1460 17 -1459
rect 30 -1460 31 -1459
rect 226 -1460 227 -1459
rect 345 -1460 346 -1459
rect 359 -1460 360 -1459
rect 443 -1460 444 -1459
rect 485 -1460 486 -1459
rect 555 -1460 556 -1459
rect 919 -1460 920 -1459
rect 968 -1460 969 -1459
rect 1017 -1460 1018 -1459
rect 1087 -1460 1088 -1459
rect 1136 -1460 1137 -1459
rect 1304 -1460 1305 -1459
rect 1374 -1460 1375 -1459
rect 1388 -1460 1389 -1459
rect 30 -1462 31 -1461
rect 506 -1462 507 -1461
rect 877 -1462 878 -1461
rect 968 -1462 969 -1461
rect 989 -1462 990 -1461
rect 1136 -1462 1137 -1461
rect 1150 -1462 1151 -1461
rect 1178 -1462 1179 -1461
rect 1220 -1462 1221 -1461
rect 1227 -1462 1228 -1461
rect 107 -1464 108 -1463
rect 506 -1464 507 -1463
rect 758 -1464 759 -1463
rect 877 -1464 878 -1463
rect 926 -1464 927 -1463
rect 975 -1464 976 -1463
rect 989 -1464 990 -1463
rect 1402 -1464 1403 -1463
rect 107 -1466 108 -1465
rect 163 -1466 164 -1465
rect 240 -1466 241 -1465
rect 457 -1466 458 -1465
rect 488 -1466 489 -1465
rect 1374 -1466 1375 -1465
rect 128 -1468 129 -1467
rect 163 -1468 164 -1467
rect 247 -1468 248 -1467
rect 845 -1468 846 -1467
rect 933 -1468 934 -1467
rect 999 -1468 1000 -1467
rect 1017 -1468 1018 -1467
rect 1073 -1468 1074 -1467
rect 1087 -1468 1088 -1467
rect 1094 -1468 1095 -1467
rect 1122 -1468 1123 -1467
rect 1227 -1468 1228 -1467
rect 128 -1470 129 -1469
rect 870 -1470 871 -1469
rect 940 -1470 941 -1469
rect 982 -1470 983 -1469
rect 1020 -1470 1021 -1469
rect 1493 -1470 1494 -1469
rect 79 -1472 80 -1471
rect 870 -1472 871 -1471
rect 947 -1472 948 -1471
rect 1066 -1472 1067 -1471
rect 1094 -1472 1095 -1471
rect 1108 -1472 1109 -1471
rect 1150 -1472 1151 -1471
rect 1290 -1472 1291 -1471
rect 1486 -1472 1487 -1471
rect 1493 -1472 1494 -1471
rect 247 -1474 248 -1473
rect 289 -1474 290 -1473
rect 331 -1474 332 -1473
rect 618 -1474 619 -1473
rect 632 -1474 633 -1473
rect 1122 -1474 1123 -1473
rect 1283 -1474 1284 -1473
rect 1290 -1474 1291 -1473
rect 1479 -1474 1480 -1473
rect 1486 -1474 1487 -1473
rect 282 -1476 283 -1475
rect 289 -1476 290 -1475
rect 331 -1476 332 -1475
rect 422 -1476 423 -1475
rect 443 -1476 444 -1475
rect 579 -1476 580 -1475
rect 695 -1476 696 -1475
rect 1073 -1476 1074 -1475
rect 1283 -1476 1284 -1475
rect 1500 -1476 1501 -1475
rect 282 -1478 283 -1477
rect 303 -1478 304 -1477
rect 345 -1478 346 -1477
rect 499 -1478 500 -1477
rect 502 -1478 503 -1477
rect 926 -1478 927 -1477
rect 954 -1478 955 -1477
rect 1010 -1478 1011 -1477
rect 1024 -1478 1025 -1477
rect 1066 -1478 1067 -1477
rect 1472 -1478 1473 -1477
rect 1500 -1478 1501 -1477
rect 303 -1480 304 -1479
rect 310 -1480 311 -1479
rect 352 -1480 353 -1479
rect 457 -1480 458 -1479
rect 709 -1480 710 -1479
rect 1479 -1480 1480 -1479
rect 9 -1482 10 -1481
rect 352 -1482 353 -1481
rect 387 -1482 388 -1481
rect 422 -1482 423 -1481
rect 450 -1482 451 -1481
rect 485 -1482 486 -1481
rect 716 -1482 717 -1481
rect 1402 -1482 1403 -1481
rect 1451 -1482 1452 -1481
rect 1472 -1482 1473 -1481
rect 9 -1484 10 -1483
rect 681 -1484 682 -1483
rect 758 -1484 759 -1483
rect 765 -1484 766 -1483
rect 982 -1484 983 -1483
rect 996 -1484 997 -1483
rect 1010 -1484 1011 -1483
rect 1059 -1484 1060 -1483
rect 1430 -1484 1431 -1483
rect 1451 -1484 1452 -1483
rect 54 -1486 55 -1485
rect 709 -1486 710 -1485
rect 765 -1486 766 -1485
rect 922 -1486 923 -1485
rect 1024 -1486 1025 -1485
rect 1052 -1486 1053 -1485
rect 1059 -1486 1060 -1485
rect 1171 -1486 1172 -1485
rect 1395 -1486 1396 -1485
rect 1430 -1486 1431 -1485
rect 58 -1488 59 -1487
rect 716 -1488 717 -1487
rect 751 -1488 752 -1487
rect 1052 -1488 1053 -1487
rect 1367 -1488 1368 -1487
rect 1395 -1488 1396 -1487
rect 58 -1490 59 -1489
rect 814 -1490 815 -1489
rect 1031 -1490 1032 -1489
rect 1115 -1490 1116 -1489
rect 212 -1492 213 -1491
rect 450 -1492 451 -1491
rect 471 -1492 472 -1491
rect 1171 -1492 1172 -1491
rect 149 -1494 150 -1493
rect 212 -1494 213 -1493
rect 310 -1494 311 -1493
rect 474 -1494 475 -1493
rect 751 -1494 752 -1493
rect 821 -1494 822 -1493
rect 1031 -1494 1032 -1493
rect 1157 -1494 1158 -1493
rect 149 -1496 150 -1495
rect 170 -1496 171 -1495
rect 387 -1496 388 -1495
rect 429 -1496 430 -1495
rect 681 -1496 682 -1495
rect 1157 -1496 1158 -1495
rect 401 -1498 402 -1497
rect 1108 -1498 1109 -1497
rect 2 -1500 3 -1499
rect 401 -1500 402 -1499
rect 415 -1500 416 -1499
rect 1367 -1500 1368 -1499
rect 2 -1502 3 -1501
rect 142 -1502 143 -1501
rect 373 -1502 374 -1501
rect 415 -1502 416 -1501
rect 429 -1502 430 -1501
rect 891 -1502 892 -1501
rect 1038 -1502 1039 -1501
rect 1185 -1502 1186 -1501
rect 142 -1504 143 -1503
rect 156 -1504 157 -1503
rect 373 -1504 374 -1503
rect 380 -1504 381 -1503
rect 814 -1504 815 -1503
rect 1339 -1504 1340 -1503
rect 86 -1506 87 -1505
rect 380 -1506 381 -1505
rect 821 -1506 822 -1505
rect 863 -1506 864 -1505
rect 891 -1506 892 -1505
rect 912 -1506 913 -1505
rect 1101 -1506 1102 -1505
rect 1185 -1506 1186 -1505
rect 86 -1508 87 -1507
rect 604 -1508 605 -1507
rect 639 -1508 640 -1507
rect 863 -1508 864 -1507
rect 1101 -1508 1102 -1507
rect 1199 -1508 1200 -1507
rect 110 -1510 111 -1509
rect 1339 -1510 1340 -1509
rect 156 -1512 157 -1511
rect 576 -1512 577 -1511
rect 604 -1512 605 -1511
rect 625 -1512 626 -1511
rect 639 -1512 640 -1511
rect 667 -1512 668 -1511
rect 786 -1512 787 -1511
rect 912 -1512 913 -1511
rect 534 -1514 535 -1513
rect 667 -1514 668 -1513
rect 786 -1514 787 -1513
rect 828 -1514 829 -1513
rect 534 -1516 535 -1515
rect 597 -1516 598 -1515
rect 611 -1516 612 -1515
rect 625 -1516 626 -1515
rect 817 -1516 818 -1515
rect 1199 -1516 1200 -1515
rect 576 -1518 577 -1517
rect 1125 -1518 1126 -1517
rect 597 -1520 598 -1519
rect 1437 -1520 1438 -1519
rect 611 -1522 612 -1521
rect 702 -1522 703 -1521
rect 828 -1522 829 -1521
rect 1318 -1522 1319 -1521
rect 702 -1524 703 -1523
rect 737 -1524 738 -1523
rect 737 -1526 738 -1525
rect 793 -1526 794 -1525
rect 394 -1528 395 -1527
rect 793 -1528 794 -1527
rect 2 -1539 3 -1538
rect 131 -1539 132 -1538
rect 142 -1539 143 -1538
rect 173 -1539 174 -1538
rect 212 -1539 213 -1538
rect 432 -1539 433 -1538
rect 471 -1539 472 -1538
rect 667 -1539 668 -1538
rect 674 -1539 675 -1538
rect 1325 -1539 1326 -1538
rect 1349 -1539 1350 -1538
rect 1535 -1539 1536 -1538
rect 2 -1541 3 -1540
rect 275 -1541 276 -1540
rect 345 -1541 346 -1540
rect 856 -1541 857 -1540
rect 859 -1541 860 -1540
rect 1514 -1541 1515 -1540
rect 9 -1543 10 -1542
rect 12 -1543 13 -1542
rect 30 -1543 31 -1542
rect 446 -1543 447 -1542
rect 474 -1543 475 -1542
rect 817 -1543 818 -1542
rect 838 -1543 839 -1542
rect 1220 -1543 1221 -1542
rect 1325 -1543 1326 -1542
rect 1395 -1543 1396 -1542
rect 9 -1545 10 -1544
rect 485 -1545 486 -1544
rect 502 -1545 503 -1544
rect 625 -1545 626 -1544
rect 639 -1545 640 -1544
rect 754 -1545 755 -1544
rect 758 -1545 759 -1544
rect 768 -1545 769 -1544
rect 782 -1545 783 -1544
rect 849 -1545 850 -1544
rect 880 -1545 881 -1544
rect 1185 -1545 1186 -1544
rect 1220 -1545 1221 -1544
rect 1297 -1545 1298 -1544
rect 30 -1547 31 -1546
rect 135 -1547 136 -1546
rect 142 -1547 143 -1546
rect 632 -1547 633 -1546
rect 639 -1547 640 -1546
rect 653 -1547 654 -1546
rect 667 -1547 668 -1546
rect 807 -1547 808 -1546
rect 849 -1547 850 -1546
rect 863 -1547 864 -1546
rect 947 -1547 948 -1546
rect 950 -1547 951 -1546
rect 992 -1547 993 -1546
rect 1332 -1547 1333 -1546
rect 44 -1549 45 -1548
rect 275 -1549 276 -1548
rect 366 -1549 367 -1548
rect 632 -1549 633 -1548
rect 653 -1549 654 -1548
rect 716 -1549 717 -1548
rect 765 -1549 766 -1548
rect 1171 -1549 1172 -1548
rect 1185 -1549 1186 -1548
rect 1248 -1549 1249 -1548
rect 1297 -1549 1298 -1548
rect 1374 -1549 1375 -1548
rect 44 -1551 45 -1550
rect 611 -1551 612 -1550
rect 618 -1551 619 -1550
rect 674 -1551 675 -1550
rect 677 -1551 678 -1550
rect 1521 -1551 1522 -1550
rect 51 -1553 52 -1552
rect 107 -1553 108 -1552
rect 128 -1553 129 -1552
rect 212 -1553 213 -1552
rect 397 -1553 398 -1552
rect 1402 -1553 1403 -1552
rect 51 -1555 52 -1554
rect 562 -1555 563 -1554
rect 579 -1555 580 -1554
rect 730 -1555 731 -1554
rect 765 -1555 766 -1554
rect 957 -1555 958 -1554
rect 996 -1555 997 -1554
rect 1115 -1555 1116 -1554
rect 1122 -1555 1123 -1554
rect 1409 -1555 1410 -1554
rect 54 -1557 55 -1556
rect 772 -1557 773 -1556
rect 863 -1557 864 -1556
rect 919 -1557 920 -1556
rect 947 -1557 948 -1556
rect 1003 -1557 1004 -1556
rect 1073 -1557 1074 -1556
rect 1500 -1557 1501 -1556
rect 65 -1559 66 -1558
rect 502 -1559 503 -1558
rect 506 -1559 507 -1558
rect 807 -1559 808 -1558
rect 919 -1559 920 -1558
rect 982 -1559 983 -1558
rect 992 -1559 993 -1558
rect 1073 -1559 1074 -1558
rect 1115 -1559 1116 -1558
rect 1143 -1559 1144 -1558
rect 1150 -1559 1151 -1558
rect 1153 -1559 1154 -1558
rect 1171 -1559 1172 -1558
rect 1234 -1559 1235 -1558
rect 1374 -1559 1375 -1558
rect 1451 -1559 1452 -1558
rect 65 -1561 66 -1560
rect 72 -1561 73 -1560
rect 75 -1561 76 -1560
rect 527 -1561 528 -1560
rect 583 -1561 584 -1560
rect 649 -1561 650 -1560
rect 681 -1561 682 -1560
rect 1080 -1561 1081 -1560
rect 1101 -1561 1102 -1560
rect 1143 -1561 1144 -1560
rect 1150 -1561 1151 -1560
rect 1199 -1561 1200 -1560
rect 1234 -1561 1235 -1560
rect 1416 -1561 1417 -1560
rect 1451 -1561 1452 -1560
rect 1528 -1561 1529 -1560
rect 58 -1563 59 -1562
rect 527 -1563 528 -1562
rect 583 -1563 584 -1562
rect 590 -1563 591 -1562
rect 600 -1563 601 -1562
rect 751 -1563 752 -1562
rect 800 -1563 801 -1562
rect 1080 -1563 1081 -1562
rect 1101 -1563 1102 -1562
rect 1108 -1563 1109 -1562
rect 1192 -1563 1193 -1562
rect 1248 -1563 1249 -1562
rect 1283 -1563 1284 -1562
rect 1416 -1563 1417 -1562
rect 58 -1565 59 -1564
rect 373 -1565 374 -1564
rect 394 -1565 395 -1564
rect 1409 -1565 1410 -1564
rect 72 -1567 73 -1566
rect 254 -1567 255 -1566
rect 373 -1567 374 -1566
rect 457 -1567 458 -1566
rect 478 -1567 479 -1566
rect 831 -1567 832 -1566
rect 982 -1567 983 -1566
rect 1017 -1567 1018 -1566
rect 1059 -1567 1060 -1566
rect 1108 -1567 1109 -1566
rect 1192 -1567 1193 -1566
rect 1269 -1567 1270 -1566
rect 1283 -1567 1284 -1566
rect 1311 -1567 1312 -1566
rect 1402 -1567 1403 -1566
rect 1479 -1567 1480 -1566
rect 79 -1569 80 -1568
rect 114 -1569 115 -1568
rect 135 -1569 136 -1568
rect 723 -1569 724 -1568
rect 730 -1569 731 -1568
rect 793 -1569 794 -1568
rect 800 -1569 801 -1568
rect 842 -1569 843 -1568
rect 989 -1569 990 -1568
rect 1017 -1569 1018 -1568
rect 1024 -1569 1025 -1568
rect 1269 -1569 1270 -1568
rect 1311 -1569 1312 -1568
rect 1458 -1569 1459 -1568
rect 82 -1571 83 -1570
rect 492 -1571 493 -1570
rect 506 -1571 507 -1570
rect 870 -1571 871 -1570
rect 898 -1571 899 -1570
rect 1024 -1571 1025 -1570
rect 1059 -1571 1060 -1570
rect 1395 -1571 1396 -1570
rect 103 -1573 104 -1572
rect 226 -1573 227 -1572
rect 380 -1573 381 -1572
rect 478 -1573 479 -1572
rect 492 -1573 493 -1572
rect 520 -1573 521 -1572
rect 590 -1573 591 -1572
rect 702 -1573 703 -1572
rect 716 -1573 717 -1572
rect 737 -1573 738 -1572
rect 751 -1573 752 -1572
rect 1031 -1573 1032 -1572
rect 107 -1575 108 -1574
rect 338 -1575 339 -1574
rect 348 -1575 349 -1574
rect 380 -1575 381 -1574
rect 394 -1575 395 -1574
rect 555 -1575 556 -1574
rect 611 -1575 612 -1574
rect 660 -1575 661 -1574
rect 681 -1575 682 -1574
rect 695 -1575 696 -1574
rect 702 -1575 703 -1574
rect 786 -1575 787 -1574
rect 793 -1575 794 -1574
rect 1524 -1575 1525 -1574
rect 114 -1577 115 -1576
rect 261 -1577 262 -1576
rect 338 -1577 339 -1576
rect 726 -1577 727 -1576
rect 737 -1577 738 -1576
rect 1262 -1577 1263 -1576
rect 145 -1579 146 -1578
rect 744 -1579 745 -1578
rect 786 -1579 787 -1578
rect 814 -1579 815 -1578
rect 870 -1579 871 -1578
rect 926 -1579 927 -1578
rect 933 -1579 934 -1578
rect 1031 -1579 1032 -1578
rect 1262 -1579 1263 -1578
rect 1339 -1579 1340 -1578
rect 128 -1581 129 -1580
rect 933 -1581 934 -1580
rect 996 -1581 997 -1580
rect 1076 -1581 1077 -1580
rect 1255 -1581 1256 -1580
rect 1339 -1581 1340 -1580
rect 156 -1583 157 -1582
rect 625 -1583 626 -1582
rect 646 -1583 647 -1582
rect 831 -1583 832 -1582
rect 898 -1583 899 -1582
rect 975 -1583 976 -1582
rect 999 -1583 1000 -1582
rect 1129 -1583 1130 -1582
rect 156 -1585 157 -1584
rect 271 -1585 272 -1584
rect 408 -1585 409 -1584
rect 772 -1585 773 -1584
rect 814 -1585 815 -1584
rect 884 -1585 885 -1584
rect 975 -1585 976 -1584
rect 1038 -1585 1039 -1584
rect 1045 -1585 1046 -1584
rect 1255 -1585 1256 -1584
rect 163 -1587 164 -1586
rect 842 -1587 843 -1586
rect 884 -1587 885 -1586
rect 961 -1587 962 -1586
rect 1038 -1587 1039 -1586
rect 1087 -1587 1088 -1586
rect 1129 -1587 1130 -1586
rect 1157 -1587 1158 -1586
rect 163 -1589 164 -1588
rect 401 -1589 402 -1588
rect 429 -1589 430 -1588
rect 464 -1589 465 -1588
rect 474 -1589 475 -1588
rect 520 -1589 521 -1588
rect 555 -1589 556 -1588
rect 1367 -1589 1368 -1588
rect 170 -1591 171 -1590
rect 439 -1591 440 -1590
rect 450 -1591 451 -1590
rect 758 -1591 759 -1590
rect 817 -1591 818 -1590
rect 926 -1591 927 -1590
rect 1045 -1591 1046 -1590
rect 1094 -1591 1095 -1590
rect 1157 -1591 1158 -1590
rect 1213 -1591 1214 -1590
rect 1367 -1591 1368 -1590
rect 1444 -1591 1445 -1590
rect 170 -1593 171 -1592
rect 205 -1593 206 -1592
rect 261 -1593 262 -1592
rect 310 -1593 311 -1592
rect 352 -1593 353 -1592
rect 401 -1593 402 -1592
rect 415 -1593 416 -1592
rect 464 -1593 465 -1592
rect 499 -1593 500 -1592
rect 961 -1593 962 -1592
rect 1094 -1593 1095 -1592
rect 1276 -1593 1277 -1592
rect 100 -1595 101 -1594
rect 205 -1595 206 -1594
rect 240 -1595 241 -1594
rect 310 -1595 311 -1594
rect 331 -1595 332 -1594
rect 415 -1595 416 -1594
rect 450 -1595 451 -1594
rect 803 -1595 804 -1594
rect 1213 -1595 1214 -1594
rect 1430 -1595 1431 -1594
rect 100 -1597 101 -1596
rect 121 -1597 122 -1596
rect 177 -1597 178 -1596
rect 485 -1597 486 -1596
rect 499 -1597 500 -1596
rect 1332 -1597 1333 -1596
rect 93 -1599 94 -1598
rect 121 -1599 122 -1598
rect 177 -1599 178 -1598
rect 597 -1599 598 -1598
rect 621 -1599 622 -1598
rect 912 -1599 913 -1598
rect 1052 -1599 1053 -1598
rect 1430 -1599 1431 -1598
rect 93 -1601 94 -1600
rect 219 -1601 220 -1600
rect 240 -1601 241 -1600
rect 387 -1601 388 -1600
rect 457 -1601 458 -1600
rect 513 -1601 514 -1600
rect 646 -1601 647 -1600
rect 1136 -1601 1137 -1600
rect 1153 -1601 1154 -1600
rect 1199 -1601 1200 -1600
rect 1276 -1601 1277 -1600
rect 1346 -1601 1347 -1600
rect 86 -1603 87 -1602
rect 513 -1603 514 -1602
rect 660 -1603 661 -1602
rect 688 -1603 689 -1602
rect 695 -1603 696 -1602
rect 779 -1603 780 -1602
rect 912 -1603 913 -1602
rect 968 -1603 969 -1602
rect 989 -1603 990 -1602
rect 1346 -1603 1347 -1602
rect 86 -1605 87 -1604
rect 282 -1605 283 -1604
rect 296 -1605 297 -1604
rect 352 -1605 353 -1604
rect 369 -1605 370 -1604
rect 387 -1605 388 -1604
rect 471 -1605 472 -1604
rect 688 -1605 689 -1604
rect 723 -1605 724 -1604
rect 821 -1605 822 -1604
rect 968 -1605 969 -1604
rect 1164 -1605 1165 -1604
rect 184 -1607 185 -1606
rect 366 -1607 367 -1606
rect 684 -1607 685 -1606
rect 1507 -1607 1508 -1606
rect 184 -1609 185 -1608
rect 233 -1609 234 -1608
rect 282 -1609 283 -1608
rect 289 -1609 290 -1608
rect 331 -1609 332 -1608
rect 565 -1609 566 -1608
rect 740 -1609 741 -1608
rect 1087 -1609 1088 -1608
rect 1136 -1609 1137 -1608
rect 1178 -1609 1179 -1608
rect 191 -1611 192 -1610
rect 408 -1611 409 -1610
rect 744 -1611 745 -1610
rect 835 -1611 836 -1610
rect 1052 -1611 1053 -1610
rect 1318 -1611 1319 -1610
rect 191 -1613 192 -1612
rect 618 -1613 619 -1612
rect 709 -1613 710 -1612
rect 1318 -1613 1319 -1612
rect 198 -1615 199 -1614
rect 254 -1615 255 -1614
rect 289 -1615 290 -1614
rect 359 -1615 360 -1614
rect 548 -1615 549 -1614
rect 709 -1615 710 -1614
rect 779 -1615 780 -1614
rect 1066 -1615 1067 -1614
rect 1164 -1615 1165 -1614
rect 1227 -1615 1228 -1614
rect 198 -1617 199 -1616
rect 268 -1617 269 -1616
rect 359 -1617 360 -1616
rect 576 -1617 577 -1616
rect 821 -1617 822 -1616
rect 828 -1617 829 -1616
rect 835 -1617 836 -1616
rect 891 -1617 892 -1616
rect 905 -1617 906 -1616
rect 1066 -1617 1067 -1616
rect 1178 -1617 1179 -1616
rect 1241 -1617 1242 -1616
rect 219 -1619 220 -1618
rect 247 -1619 248 -1618
rect 541 -1619 542 -1618
rect 576 -1619 577 -1618
rect 828 -1619 829 -1618
rect 1122 -1619 1123 -1618
rect 1227 -1619 1228 -1618
rect 1353 -1619 1354 -1618
rect 226 -1621 227 -1620
rect 268 -1621 269 -1620
rect 422 -1621 423 -1620
rect 541 -1621 542 -1620
rect 548 -1621 549 -1620
rect 604 -1621 605 -1620
rect 891 -1621 892 -1620
rect 954 -1621 955 -1620
rect 1241 -1621 1242 -1620
rect 1304 -1621 1305 -1620
rect 1353 -1621 1354 -1620
rect 1381 -1621 1382 -1620
rect 233 -1623 234 -1622
rect 558 -1623 559 -1622
rect 569 -1623 570 -1622
rect 604 -1623 605 -1622
rect 905 -1623 906 -1622
rect 940 -1623 941 -1622
rect 954 -1623 955 -1622
rect 1360 -1623 1361 -1622
rect 1381 -1623 1382 -1622
rect 1465 -1623 1466 -1622
rect 247 -1625 248 -1624
rect 443 -1625 444 -1624
rect 877 -1625 878 -1624
rect 940 -1625 941 -1624
rect 1304 -1625 1305 -1624
rect 1388 -1625 1389 -1624
rect 296 -1627 297 -1626
rect 443 -1627 444 -1626
rect 877 -1627 878 -1626
rect 1206 -1627 1207 -1626
rect 1360 -1627 1361 -1626
rect 1437 -1627 1438 -1626
rect 324 -1629 325 -1628
rect 422 -1629 423 -1628
rect 436 -1629 437 -1628
rect 569 -1629 570 -1628
rect 1206 -1629 1207 -1628
rect 1290 -1629 1291 -1628
rect 1388 -1629 1389 -1628
rect 1472 -1629 1473 -1628
rect 317 -1631 318 -1630
rect 324 -1631 325 -1630
rect 1290 -1631 1291 -1630
rect 1423 -1631 1424 -1630
rect 1437 -1631 1438 -1630
rect 1486 -1631 1487 -1630
rect 37 -1633 38 -1632
rect 317 -1633 318 -1632
rect 1423 -1633 1424 -1632
rect 1493 -1633 1494 -1632
rect 37 -1635 38 -1634
rect 562 -1635 563 -1634
rect 2 -1646 3 -1645
rect 436 -1646 437 -1645
rect 446 -1646 447 -1645
rect 474 -1646 475 -1645
rect 488 -1646 489 -1645
rect 1206 -1646 1207 -1645
rect 1283 -1646 1284 -1645
rect 1346 -1646 1347 -1645
rect 1377 -1646 1378 -1645
rect 1451 -1646 1452 -1645
rect 37 -1648 38 -1647
rect 341 -1648 342 -1647
rect 429 -1648 430 -1647
rect 443 -1648 444 -1647
rect 471 -1648 472 -1647
rect 597 -1648 598 -1647
rect 621 -1648 622 -1647
rect 765 -1648 766 -1647
rect 814 -1648 815 -1647
rect 1017 -1648 1018 -1647
rect 1206 -1648 1207 -1647
rect 1297 -1648 1298 -1647
rect 37 -1650 38 -1649
rect 387 -1650 388 -1649
rect 429 -1650 430 -1649
rect 520 -1650 521 -1649
rect 555 -1650 556 -1649
rect 667 -1650 668 -1649
rect 709 -1650 710 -1649
rect 873 -1650 874 -1649
rect 877 -1650 878 -1649
rect 1003 -1650 1004 -1649
rect 1017 -1650 1018 -1649
rect 1150 -1650 1151 -1649
rect 1283 -1650 1284 -1649
rect 1367 -1650 1368 -1649
rect 65 -1652 66 -1651
rect 586 -1652 587 -1651
rect 597 -1652 598 -1651
rect 863 -1652 864 -1651
rect 877 -1652 878 -1651
rect 1297 -1652 1298 -1651
rect 1367 -1652 1368 -1651
rect 1430 -1652 1431 -1651
rect 65 -1654 66 -1653
rect 149 -1654 150 -1653
rect 163 -1654 164 -1653
rect 418 -1654 419 -1653
rect 436 -1654 437 -1653
rect 782 -1654 783 -1653
rect 828 -1654 829 -1653
rect 1094 -1654 1095 -1653
rect 1150 -1654 1151 -1653
rect 1199 -1654 1200 -1653
rect 72 -1656 73 -1655
rect 506 -1656 507 -1655
rect 513 -1656 514 -1655
rect 740 -1656 741 -1655
rect 744 -1656 745 -1655
rect 775 -1656 776 -1655
rect 817 -1656 818 -1655
rect 1199 -1656 1200 -1655
rect 82 -1658 83 -1657
rect 625 -1658 626 -1657
rect 635 -1658 636 -1657
rect 786 -1658 787 -1657
rect 828 -1658 829 -1657
rect 933 -1658 934 -1657
rect 1094 -1658 1095 -1657
rect 1304 -1658 1305 -1657
rect 128 -1660 129 -1659
rect 632 -1660 633 -1659
rect 653 -1660 654 -1659
rect 656 -1660 657 -1659
rect 667 -1660 668 -1659
rect 674 -1660 675 -1659
rect 709 -1660 710 -1659
rect 716 -1660 717 -1659
rect 719 -1660 720 -1659
rect 968 -1660 969 -1659
rect 1006 -1660 1007 -1659
rect 1304 -1660 1305 -1659
rect 128 -1662 129 -1661
rect 135 -1662 136 -1661
rect 149 -1662 150 -1661
rect 233 -1662 234 -1661
rect 240 -1662 241 -1661
rect 369 -1662 370 -1661
rect 387 -1662 388 -1661
rect 492 -1662 493 -1661
rect 513 -1662 514 -1661
rect 523 -1662 524 -1661
rect 555 -1662 556 -1661
rect 590 -1662 591 -1661
rect 604 -1662 605 -1661
rect 674 -1662 675 -1661
rect 723 -1662 724 -1661
rect 880 -1662 881 -1661
rect 933 -1662 934 -1661
rect 1080 -1662 1081 -1661
rect 9 -1664 10 -1663
rect 369 -1664 370 -1663
rect 471 -1664 472 -1663
rect 737 -1664 738 -1663
rect 751 -1664 752 -1663
rect 1346 -1664 1347 -1663
rect 9 -1666 10 -1665
rect 93 -1666 94 -1665
rect 121 -1666 122 -1665
rect 135 -1666 136 -1665
rect 142 -1666 143 -1665
rect 233 -1666 234 -1665
rect 240 -1666 241 -1665
rect 254 -1666 255 -1665
rect 303 -1666 304 -1665
rect 345 -1666 346 -1665
rect 359 -1666 360 -1665
rect 632 -1666 633 -1665
rect 653 -1666 654 -1665
rect 688 -1666 689 -1665
rect 751 -1666 752 -1665
rect 821 -1666 822 -1665
rect 863 -1666 864 -1665
rect 891 -1666 892 -1665
rect 968 -1666 969 -1665
rect 1038 -1666 1039 -1665
rect 1080 -1666 1081 -1665
rect 1185 -1666 1186 -1665
rect 93 -1668 94 -1667
rect 548 -1668 549 -1667
rect 562 -1668 563 -1667
rect 1255 -1668 1256 -1667
rect 114 -1670 115 -1669
rect 303 -1670 304 -1669
rect 310 -1670 311 -1669
rect 520 -1670 521 -1669
rect 527 -1670 528 -1669
rect 562 -1670 563 -1669
rect 565 -1670 566 -1669
rect 807 -1670 808 -1669
rect 821 -1670 822 -1669
rect 884 -1670 885 -1669
rect 891 -1670 892 -1669
rect 947 -1670 948 -1669
rect 1038 -1670 1039 -1669
rect 1143 -1670 1144 -1669
rect 1255 -1670 1256 -1669
rect 1290 -1670 1291 -1669
rect 79 -1672 80 -1671
rect 114 -1672 115 -1671
rect 121 -1672 122 -1671
rect 156 -1672 157 -1671
rect 163 -1672 164 -1671
rect 184 -1672 185 -1671
rect 198 -1672 199 -1671
rect 271 -1672 272 -1671
rect 310 -1672 311 -1671
rect 401 -1672 402 -1671
rect 408 -1672 409 -1671
rect 548 -1672 549 -1671
rect 590 -1672 591 -1671
rect 660 -1672 661 -1671
rect 758 -1672 759 -1671
rect 831 -1672 832 -1671
rect 845 -1672 846 -1671
rect 1185 -1672 1186 -1671
rect 1290 -1672 1291 -1671
rect 1374 -1672 1375 -1671
rect 58 -1674 59 -1673
rect 156 -1674 157 -1673
rect 177 -1674 178 -1673
rect 499 -1674 500 -1673
rect 604 -1674 605 -1673
rect 779 -1674 780 -1673
rect 786 -1674 787 -1673
rect 989 -1674 990 -1673
rect 58 -1676 59 -1675
rect 541 -1676 542 -1675
rect 625 -1676 626 -1675
rect 639 -1676 640 -1675
rect 656 -1676 657 -1675
rect 688 -1676 689 -1675
rect 758 -1676 759 -1675
rect 1031 -1676 1032 -1675
rect 79 -1678 80 -1677
rect 324 -1678 325 -1677
rect 345 -1678 346 -1677
rect 415 -1678 416 -1677
rect 485 -1678 486 -1677
rect 737 -1678 738 -1677
rect 765 -1678 766 -1677
rect 961 -1678 962 -1677
rect 1031 -1678 1032 -1677
rect 1157 -1678 1158 -1677
rect 110 -1680 111 -1679
rect 408 -1680 409 -1679
rect 492 -1680 493 -1679
rect 649 -1680 650 -1679
rect 660 -1680 661 -1679
rect 730 -1680 731 -1679
rect 779 -1680 780 -1679
rect 835 -1680 836 -1679
rect 880 -1680 881 -1679
rect 1010 -1680 1011 -1679
rect 1157 -1680 1158 -1679
rect 1241 -1680 1242 -1679
rect 110 -1682 111 -1681
rect 842 -1682 843 -1681
rect 884 -1682 885 -1681
rect 905 -1682 906 -1681
rect 926 -1682 927 -1681
rect 1143 -1682 1144 -1681
rect 142 -1684 143 -1683
rect 695 -1684 696 -1683
rect 730 -1684 731 -1683
rect 849 -1684 850 -1683
rect 905 -1684 906 -1683
rect 1349 -1684 1350 -1683
rect 177 -1686 178 -1685
rect 754 -1686 755 -1685
rect 835 -1686 836 -1685
rect 870 -1686 871 -1685
rect 926 -1686 927 -1685
rect 1101 -1686 1102 -1685
rect 184 -1688 185 -1687
rect 425 -1688 426 -1687
rect 506 -1688 507 -1687
rect 1241 -1688 1242 -1687
rect 198 -1690 199 -1689
rect 954 -1690 955 -1689
rect 961 -1690 962 -1689
rect 982 -1690 983 -1689
rect 1010 -1690 1011 -1689
rect 1171 -1690 1172 -1689
rect 205 -1692 206 -1691
rect 527 -1692 528 -1691
rect 576 -1692 577 -1691
rect 695 -1692 696 -1691
rect 842 -1692 843 -1691
rect 1227 -1692 1228 -1691
rect 205 -1694 206 -1693
rect 261 -1694 262 -1693
rect 268 -1694 269 -1693
rect 499 -1694 500 -1693
rect 576 -1694 577 -1693
rect 1003 -1694 1004 -1693
rect 1101 -1694 1102 -1693
rect 1220 -1694 1221 -1693
rect 1227 -1694 1228 -1693
rect 1409 -1694 1410 -1693
rect 219 -1696 220 -1695
rect 261 -1696 262 -1695
rect 268 -1696 269 -1695
rect 317 -1696 318 -1695
rect 359 -1696 360 -1695
rect 464 -1696 465 -1695
rect 611 -1696 612 -1695
rect 639 -1696 640 -1695
rect 849 -1696 850 -1695
rect 919 -1696 920 -1695
rect 947 -1696 948 -1695
rect 1045 -1696 1046 -1695
rect 1220 -1696 1221 -1695
rect 1318 -1696 1319 -1695
rect 219 -1698 220 -1697
rect 796 -1698 797 -1697
rect 870 -1698 871 -1697
rect 1234 -1698 1235 -1697
rect 1248 -1698 1249 -1697
rect 1318 -1698 1319 -1697
rect 254 -1700 255 -1699
rect 415 -1700 416 -1699
rect 464 -1700 465 -1699
rect 478 -1700 479 -1699
rect 611 -1700 612 -1699
rect 856 -1700 857 -1699
rect 901 -1700 902 -1699
rect 1248 -1700 1249 -1699
rect 289 -1702 290 -1701
rect 317 -1702 318 -1701
rect 366 -1702 367 -1701
rect 744 -1702 745 -1701
rect 856 -1702 857 -1701
rect 898 -1702 899 -1701
rect 919 -1702 920 -1701
rect 1087 -1702 1088 -1701
rect 1234 -1702 1235 -1701
rect 1388 -1702 1389 -1701
rect 212 -1704 213 -1703
rect 366 -1704 367 -1703
rect 394 -1704 395 -1703
rect 541 -1704 542 -1703
rect 898 -1704 899 -1703
rect 940 -1704 941 -1703
rect 954 -1704 955 -1703
rect 1129 -1704 1130 -1703
rect 131 -1706 132 -1705
rect 1129 -1706 1130 -1705
rect 212 -1708 213 -1707
rect 275 -1708 276 -1707
rect 282 -1708 283 -1707
rect 289 -1708 290 -1707
rect 296 -1708 297 -1707
rect 324 -1708 325 -1707
rect 394 -1708 395 -1707
rect 422 -1708 423 -1707
rect 478 -1708 479 -1707
rect 534 -1708 535 -1707
rect 940 -1708 941 -1707
rect 975 -1708 976 -1707
rect 982 -1708 983 -1707
rect 1073 -1708 1074 -1707
rect 1087 -1708 1088 -1707
rect 1192 -1708 1193 -1707
rect 75 -1710 76 -1709
rect 296 -1710 297 -1709
rect 401 -1710 402 -1709
rect 569 -1710 570 -1709
rect 975 -1710 976 -1709
rect 1122 -1710 1123 -1709
rect 1192 -1710 1193 -1709
rect 1262 -1710 1263 -1709
rect 75 -1712 76 -1711
rect 723 -1712 724 -1711
rect 996 -1712 997 -1711
rect 1171 -1712 1172 -1711
rect 1262 -1712 1263 -1711
rect 1332 -1712 1333 -1711
rect 107 -1714 108 -1713
rect 275 -1714 276 -1713
rect 282 -1714 283 -1713
rect 373 -1714 374 -1713
rect 380 -1714 381 -1713
rect 569 -1714 570 -1713
rect 996 -1714 997 -1713
rect 1108 -1714 1109 -1713
rect 1332 -1714 1333 -1713
rect 1402 -1714 1403 -1713
rect 72 -1716 73 -1715
rect 380 -1716 381 -1715
rect 422 -1716 423 -1715
rect 583 -1716 584 -1715
rect 1024 -1716 1025 -1715
rect 1409 -1716 1410 -1715
rect 107 -1718 108 -1717
rect 450 -1718 451 -1717
rect 502 -1718 503 -1717
rect 1024 -1718 1025 -1717
rect 1045 -1718 1046 -1717
rect 1164 -1718 1165 -1717
rect 1402 -1718 1403 -1717
rect 1423 -1718 1424 -1717
rect 247 -1720 248 -1719
rect 373 -1720 374 -1719
rect 534 -1720 535 -1719
rect 793 -1720 794 -1719
rect 1052 -1720 1053 -1719
rect 1122 -1720 1123 -1719
rect 1164 -1720 1165 -1719
rect 1276 -1720 1277 -1719
rect 1423 -1720 1424 -1719
rect 1437 -1720 1438 -1719
rect 145 -1722 146 -1721
rect 247 -1722 248 -1721
rect 331 -1722 332 -1721
rect 450 -1722 451 -1721
rect 793 -1722 794 -1721
rect 1311 -1722 1312 -1721
rect 331 -1724 332 -1723
rect 352 -1724 353 -1723
rect 810 -1724 811 -1723
rect 1052 -1724 1053 -1723
rect 1066 -1724 1067 -1723
rect 1388 -1724 1389 -1723
rect 338 -1726 339 -1725
rect 352 -1726 353 -1725
rect 992 -1726 993 -1725
rect 1311 -1726 1312 -1725
rect 30 -1728 31 -1727
rect 338 -1728 339 -1727
rect 992 -1728 993 -1727
rect 1339 -1728 1340 -1727
rect 16 -1730 17 -1729
rect 30 -1730 31 -1729
rect 646 -1730 647 -1729
rect 1339 -1730 1340 -1729
rect 16 -1732 17 -1731
rect 100 -1732 101 -1731
rect 646 -1732 647 -1731
rect 681 -1732 682 -1731
rect 1066 -1732 1067 -1731
rect 1115 -1732 1116 -1731
rect 1276 -1732 1277 -1731
rect 1360 -1732 1361 -1731
rect 100 -1734 101 -1733
rect 191 -1734 192 -1733
rect 530 -1734 531 -1733
rect 1115 -1734 1116 -1733
rect 191 -1736 192 -1735
rect 509 -1736 510 -1735
rect 681 -1736 682 -1735
rect 702 -1736 703 -1735
rect 716 -1736 717 -1735
rect 1360 -1736 1361 -1735
rect 702 -1738 703 -1737
rect 772 -1738 773 -1737
rect 1073 -1738 1074 -1737
rect 1178 -1738 1179 -1737
rect 772 -1740 773 -1739
rect 1269 -1740 1270 -1739
rect 1108 -1742 1109 -1741
rect 1136 -1742 1137 -1741
rect 1178 -1742 1179 -1741
rect 1381 -1742 1382 -1741
rect 1136 -1744 1137 -1743
rect 1325 -1744 1326 -1743
rect 1374 -1744 1375 -1743
rect 1381 -1744 1382 -1743
rect 618 -1746 619 -1745
rect 1325 -1746 1326 -1745
rect 44 -1748 45 -1747
rect 618 -1748 619 -1747
rect 1213 -1748 1214 -1747
rect 1269 -1748 1270 -1747
rect 44 -1750 45 -1749
rect 226 -1750 227 -1749
rect 1213 -1750 1214 -1749
rect 1395 -1750 1396 -1749
rect 86 -1752 87 -1751
rect 226 -1752 227 -1751
rect 1353 -1752 1354 -1751
rect 1395 -1752 1396 -1751
rect 86 -1754 87 -1753
rect 170 -1754 171 -1753
rect 1353 -1754 1354 -1753
rect 1416 -1754 1417 -1753
rect 170 -1756 171 -1755
rect 457 -1756 458 -1755
rect 912 -1756 913 -1755
rect 1416 -1756 1417 -1755
rect 457 -1758 458 -1757
rect 583 -1758 584 -1757
rect 912 -1758 913 -1757
rect 1059 -1758 1060 -1757
rect 1059 -1760 1060 -1759
rect 1370 -1760 1371 -1759
rect 2 -1771 3 -1770
rect 590 -1771 591 -1770
rect 667 -1771 668 -1770
rect 842 -1771 843 -1770
rect 877 -1771 878 -1770
rect 1157 -1771 1158 -1770
rect 1255 -1771 1256 -1770
rect 1258 -1771 1259 -1770
rect 1360 -1771 1361 -1770
rect 1370 -1771 1371 -1770
rect 1377 -1771 1378 -1770
rect 1395 -1771 1396 -1770
rect 19 -1773 20 -1772
rect 534 -1773 535 -1772
rect 562 -1773 563 -1772
rect 590 -1773 591 -1772
rect 667 -1773 668 -1772
rect 681 -1773 682 -1772
rect 684 -1773 685 -1772
rect 786 -1773 787 -1772
rect 793 -1773 794 -1772
rect 835 -1773 836 -1772
rect 842 -1773 843 -1772
rect 863 -1773 864 -1772
rect 887 -1773 888 -1772
rect 968 -1773 969 -1772
rect 1003 -1773 1004 -1772
rect 1066 -1773 1067 -1772
rect 1255 -1773 1256 -1772
rect 1262 -1773 1263 -1772
rect 1367 -1773 1368 -1772
rect 1402 -1773 1403 -1772
rect 61 -1775 62 -1774
rect 1227 -1775 1228 -1774
rect 1346 -1775 1347 -1774
rect 1367 -1775 1368 -1774
rect 1381 -1775 1382 -1774
rect 1430 -1775 1431 -1774
rect 72 -1777 73 -1776
rect 796 -1777 797 -1776
rect 800 -1777 801 -1776
rect 807 -1777 808 -1776
rect 814 -1777 815 -1776
rect 835 -1777 836 -1776
rect 849 -1777 850 -1776
rect 877 -1777 878 -1776
rect 898 -1777 899 -1776
rect 1192 -1777 1193 -1776
rect 1339 -1777 1340 -1776
rect 1346 -1777 1347 -1776
rect 1353 -1777 1354 -1776
rect 1381 -1777 1382 -1776
rect 30 -1779 31 -1778
rect 72 -1779 73 -1778
rect 75 -1779 76 -1778
rect 142 -1779 143 -1778
rect 247 -1779 248 -1778
rect 880 -1779 881 -1778
rect 898 -1779 899 -1778
rect 940 -1779 941 -1778
rect 968 -1779 969 -1778
rect 1059 -1779 1060 -1778
rect 1066 -1779 1067 -1778
rect 1108 -1779 1109 -1778
rect 1332 -1779 1333 -1778
rect 1339 -1779 1340 -1778
rect 1353 -1779 1354 -1778
rect 1374 -1779 1375 -1778
rect 23 -1781 24 -1780
rect 30 -1781 31 -1780
rect 89 -1781 90 -1780
rect 310 -1781 311 -1780
rect 324 -1781 325 -1780
rect 369 -1781 370 -1780
rect 373 -1781 374 -1780
rect 502 -1781 503 -1780
rect 513 -1781 514 -1780
rect 786 -1781 787 -1780
rect 793 -1781 794 -1780
rect 1395 -1781 1396 -1780
rect 23 -1783 24 -1782
rect 632 -1783 633 -1782
rect 635 -1783 636 -1782
rect 1192 -1783 1193 -1782
rect 1234 -1783 1235 -1782
rect 1332 -1783 1333 -1782
rect 51 -1785 52 -1784
rect 632 -1785 633 -1784
rect 691 -1785 692 -1784
rect 1248 -1785 1249 -1784
rect 1325 -1785 1326 -1784
rect 1374 -1785 1375 -1784
rect 51 -1787 52 -1786
rect 121 -1787 122 -1786
rect 138 -1787 139 -1786
rect 415 -1787 416 -1786
rect 436 -1787 437 -1786
rect 439 -1787 440 -1786
rect 464 -1787 465 -1786
rect 509 -1787 510 -1786
rect 513 -1787 514 -1786
rect 541 -1787 542 -1786
rect 569 -1787 570 -1786
rect 814 -1787 815 -1786
rect 849 -1787 850 -1786
rect 856 -1787 857 -1786
rect 863 -1787 864 -1786
rect 891 -1787 892 -1786
rect 908 -1787 909 -1786
rect 1150 -1787 1151 -1786
rect 1178 -1787 1179 -1786
rect 1325 -1787 1326 -1786
rect 58 -1789 59 -1788
rect 121 -1789 122 -1788
rect 191 -1789 192 -1788
rect 373 -1789 374 -1788
rect 380 -1789 381 -1788
rect 562 -1789 563 -1788
rect 569 -1789 570 -1788
rect 765 -1789 766 -1788
rect 800 -1789 801 -1788
rect 1010 -1789 1011 -1788
rect 1129 -1789 1130 -1788
rect 1150 -1789 1151 -1788
rect 1234 -1789 1235 -1788
rect 1388 -1789 1389 -1788
rect 9 -1791 10 -1790
rect 58 -1791 59 -1790
rect 82 -1791 83 -1790
rect 891 -1791 892 -1790
rect 926 -1791 927 -1790
rect 1157 -1791 1158 -1790
rect 1241 -1791 1242 -1790
rect 1248 -1791 1249 -1790
rect 9 -1793 10 -1792
rect 156 -1793 157 -1792
rect 191 -1793 192 -1792
rect 268 -1793 269 -1792
rect 275 -1793 276 -1792
rect 663 -1793 664 -1792
rect 716 -1793 717 -1792
rect 1108 -1793 1109 -1792
rect 1136 -1793 1137 -1792
rect 1241 -1793 1242 -1792
rect 37 -1795 38 -1794
rect 156 -1795 157 -1794
rect 212 -1795 213 -1794
rect 268 -1795 269 -1794
rect 289 -1795 290 -1794
rect 299 -1795 300 -1794
rect 310 -1795 311 -1794
rect 422 -1795 423 -1794
rect 436 -1795 437 -1794
rect 457 -1795 458 -1794
rect 464 -1795 465 -1794
rect 695 -1795 696 -1794
rect 719 -1795 720 -1794
rect 982 -1795 983 -1794
rect 989 -1795 990 -1794
rect 1129 -1795 1130 -1794
rect 107 -1797 108 -1796
rect 397 -1797 398 -1796
rect 415 -1797 416 -1796
rect 604 -1797 605 -1796
rect 611 -1797 612 -1796
rect 807 -1797 808 -1796
rect 810 -1797 811 -1796
rect 1388 -1797 1389 -1796
rect 100 -1799 101 -1798
rect 107 -1799 108 -1798
rect 114 -1799 115 -1798
rect 142 -1799 143 -1798
rect 212 -1799 213 -1798
rect 366 -1799 367 -1798
rect 380 -1799 381 -1798
rect 443 -1799 444 -1798
rect 527 -1799 528 -1798
rect 751 -1799 752 -1798
rect 765 -1799 766 -1798
rect 779 -1799 780 -1798
rect 803 -1799 804 -1798
rect 1227 -1799 1228 -1798
rect 1258 -1799 1259 -1798
rect 1262 -1799 1263 -1798
rect 100 -1801 101 -1800
rect 184 -1801 185 -1800
rect 226 -1801 227 -1800
rect 275 -1801 276 -1800
rect 296 -1801 297 -1800
rect 366 -1801 367 -1800
rect 387 -1801 388 -1800
rect 520 -1801 521 -1800
rect 527 -1801 528 -1800
rect 702 -1801 703 -1800
rect 719 -1801 720 -1800
rect 828 -1801 829 -1800
rect 856 -1801 857 -1800
rect 884 -1801 885 -1800
rect 926 -1801 927 -1800
rect 961 -1801 962 -1800
rect 989 -1801 990 -1800
rect 1171 -1801 1172 -1800
rect 65 -1803 66 -1802
rect 184 -1803 185 -1802
rect 247 -1803 248 -1802
rect 254 -1803 255 -1802
rect 261 -1803 262 -1802
rect 485 -1803 486 -1802
rect 534 -1803 535 -1802
rect 730 -1803 731 -1802
rect 737 -1803 738 -1802
rect 754 -1803 755 -1802
rect 779 -1803 780 -1802
rect 1220 -1803 1221 -1802
rect 65 -1805 66 -1804
rect 86 -1805 87 -1804
rect 114 -1805 115 -1804
rect 149 -1805 150 -1804
rect 163 -1805 164 -1804
rect 226 -1805 227 -1804
rect 233 -1805 234 -1804
rect 261 -1805 262 -1804
rect 296 -1805 297 -1804
rect 1062 -1805 1063 -1804
rect 1094 -1805 1095 -1804
rect 1220 -1805 1221 -1804
rect 135 -1807 136 -1806
rect 149 -1807 150 -1806
rect 163 -1807 164 -1806
rect 170 -1807 171 -1806
rect 233 -1807 234 -1806
rect 345 -1807 346 -1806
rect 352 -1807 353 -1806
rect 443 -1807 444 -1806
rect 485 -1807 486 -1806
rect 884 -1807 885 -1806
rect 919 -1807 920 -1806
rect 1171 -1807 1172 -1806
rect 37 -1809 38 -1808
rect 135 -1809 136 -1808
rect 240 -1809 241 -1808
rect 254 -1809 255 -1808
rect 324 -1809 325 -1808
rect 576 -1809 577 -1808
rect 604 -1809 605 -1808
rect 618 -1809 619 -1808
rect 695 -1809 696 -1808
rect 723 -1809 724 -1808
rect 737 -1809 738 -1808
rect 1017 -1809 1018 -1808
rect 1087 -1809 1088 -1808
rect 1094 -1809 1095 -1808
rect 1122 -1809 1123 -1808
rect 1136 -1809 1137 -1808
rect 44 -1811 45 -1810
rect 345 -1811 346 -1810
rect 352 -1811 353 -1810
rect 471 -1811 472 -1810
rect 488 -1811 489 -1810
rect 576 -1811 577 -1810
rect 611 -1811 612 -1810
rect 646 -1811 647 -1810
rect 702 -1811 703 -1810
rect 709 -1811 710 -1810
rect 723 -1811 724 -1810
rect 936 -1811 937 -1810
rect 940 -1811 941 -1810
rect 1416 -1811 1417 -1810
rect 44 -1813 45 -1812
rect 408 -1813 409 -1812
rect 492 -1813 493 -1812
rect 730 -1813 731 -1812
rect 744 -1813 745 -1812
rect 982 -1813 983 -1812
rect 996 -1813 997 -1812
rect 1003 -1813 1004 -1812
rect 1006 -1813 1007 -1812
rect 1318 -1813 1319 -1812
rect 93 -1815 94 -1814
rect 170 -1815 171 -1814
rect 240 -1815 241 -1814
rect 450 -1815 451 -1814
rect 530 -1815 531 -1814
rect 744 -1815 745 -1814
rect 751 -1815 752 -1814
rect 961 -1815 962 -1814
rect 975 -1815 976 -1814
rect 1017 -1815 1018 -1814
rect 1073 -1815 1074 -1814
rect 1087 -1815 1088 -1814
rect 1311 -1815 1312 -1814
rect 1318 -1815 1319 -1814
rect 93 -1817 94 -1816
rect 418 -1817 419 -1816
rect 450 -1817 451 -1816
rect 775 -1817 776 -1816
rect 821 -1817 822 -1816
rect 828 -1817 829 -1816
rect 870 -1817 871 -1816
rect 1416 -1817 1417 -1816
rect 128 -1819 129 -1818
rect 471 -1819 472 -1818
rect 506 -1819 507 -1818
rect 975 -1819 976 -1818
rect 996 -1819 997 -1818
rect 1143 -1819 1144 -1818
rect 1304 -1819 1305 -1818
rect 1311 -1819 1312 -1818
rect 128 -1821 129 -1820
rect 593 -1821 594 -1820
rect 597 -1821 598 -1820
rect 821 -1821 822 -1820
rect 870 -1821 871 -1820
rect 912 -1821 913 -1820
rect 919 -1821 920 -1820
rect 1080 -1821 1081 -1820
rect 1115 -1821 1116 -1820
rect 1143 -1821 1144 -1820
rect 1297 -1821 1298 -1820
rect 1304 -1821 1305 -1820
rect 317 -1823 318 -1822
rect 408 -1823 409 -1822
rect 478 -1823 479 -1822
rect 506 -1823 507 -1822
rect 541 -1823 542 -1822
rect 548 -1823 549 -1822
rect 555 -1823 556 -1822
rect 597 -1823 598 -1822
rect 618 -1823 619 -1822
rect 1024 -1823 1025 -1822
rect 1045 -1823 1046 -1822
rect 1073 -1823 1074 -1822
rect 1290 -1823 1291 -1822
rect 1297 -1823 1298 -1822
rect 282 -1825 283 -1824
rect 317 -1825 318 -1824
rect 331 -1825 332 -1824
rect 422 -1825 423 -1824
rect 432 -1825 433 -1824
rect 1045 -1825 1046 -1824
rect 1052 -1825 1053 -1824
rect 1080 -1825 1081 -1824
rect 1283 -1825 1284 -1824
rect 1290 -1825 1291 -1824
rect 282 -1827 283 -1826
rect 359 -1827 360 -1826
rect 387 -1827 388 -1826
rect 653 -1827 654 -1826
rect 681 -1827 682 -1826
rect 1115 -1827 1116 -1826
rect 219 -1829 220 -1828
rect 359 -1829 360 -1828
rect 401 -1829 402 -1828
rect 548 -1829 549 -1828
rect 555 -1829 556 -1828
rect 688 -1829 689 -1828
rect 709 -1829 710 -1828
rect 905 -1829 906 -1828
rect 933 -1829 934 -1828
rect 1024 -1829 1025 -1828
rect 1031 -1829 1032 -1828
rect 1052 -1829 1053 -1828
rect 1101 -1829 1102 -1828
rect 1283 -1829 1284 -1828
rect 79 -1831 80 -1830
rect 219 -1831 220 -1830
rect 303 -1831 304 -1830
rect 331 -1831 332 -1830
rect 338 -1831 339 -1830
rect 492 -1831 493 -1830
rect 558 -1831 559 -1830
rect 912 -1831 913 -1830
rect 1010 -1831 1011 -1830
rect 1206 -1831 1207 -1830
rect 16 -1833 17 -1832
rect 79 -1833 80 -1832
rect 303 -1833 304 -1832
rect 394 -1833 395 -1832
rect 401 -1833 402 -1832
rect 845 -1833 846 -1832
rect 873 -1833 874 -1832
rect 1122 -1833 1123 -1832
rect 1185 -1833 1186 -1832
rect 1206 -1833 1207 -1832
rect 86 -1835 87 -1834
rect 1185 -1835 1186 -1834
rect 338 -1837 339 -1836
rect 583 -1837 584 -1836
rect 586 -1837 587 -1836
rect 905 -1837 906 -1836
rect 1031 -1837 1032 -1836
rect 1038 -1837 1039 -1836
rect 1101 -1837 1102 -1836
rect 1409 -1837 1410 -1836
rect 341 -1839 342 -1838
rect 1213 -1839 1214 -1838
rect 394 -1841 395 -1840
rect 1360 -1841 1361 -1840
rect 478 -1843 479 -1842
rect 499 -1843 500 -1842
rect 583 -1843 584 -1842
rect 639 -1843 640 -1842
rect 653 -1843 654 -1842
rect 758 -1843 759 -1842
rect 901 -1843 902 -1842
rect 1409 -1843 1410 -1842
rect 289 -1845 290 -1844
rect 499 -1845 500 -1844
rect 625 -1845 626 -1844
rect 646 -1845 647 -1844
rect 688 -1845 689 -1844
rect 1178 -1845 1179 -1844
rect 1199 -1845 1200 -1844
rect 1213 -1845 1214 -1844
rect 625 -1847 626 -1846
rect 660 -1847 661 -1846
rect 716 -1847 717 -1846
rect 758 -1847 759 -1846
rect 954 -1847 955 -1846
rect 1199 -1847 1200 -1846
rect 639 -1849 640 -1848
rect 933 -1849 934 -1848
rect 947 -1849 948 -1848
rect 954 -1849 955 -1848
rect 1038 -1849 1039 -1848
rect 1276 -1849 1277 -1848
rect 572 -1851 573 -1850
rect 947 -1851 948 -1850
rect 1269 -1851 1270 -1850
rect 1276 -1851 1277 -1850
rect 660 -1853 661 -1852
rect 1402 -1853 1403 -1852
rect 772 -1855 773 -1854
rect 1269 -1855 1270 -1854
rect 429 -1857 430 -1856
rect 772 -1857 773 -1856
rect 2 -1868 3 -1867
rect 5 -1868 6 -1867
rect 9 -1868 10 -1867
rect 397 -1868 398 -1867
rect 432 -1868 433 -1867
rect 744 -1868 745 -1867
rect 751 -1868 752 -1867
rect 1283 -1868 1284 -1867
rect 1395 -1868 1396 -1867
rect 1423 -1868 1424 -1867
rect 2 -1870 3 -1869
rect 51 -1870 52 -1869
rect 100 -1870 101 -1869
rect 299 -1870 300 -1869
rect 373 -1870 374 -1869
rect 558 -1870 559 -1869
rect 565 -1870 566 -1869
rect 912 -1870 913 -1869
rect 933 -1870 934 -1869
rect 1381 -1870 1382 -1869
rect 9 -1872 10 -1871
rect 261 -1872 262 -1871
rect 282 -1872 283 -1871
rect 345 -1872 346 -1871
rect 471 -1872 472 -1871
rect 614 -1872 615 -1871
rect 618 -1872 619 -1871
rect 772 -1872 773 -1871
rect 775 -1872 776 -1871
rect 968 -1872 969 -1871
rect 1062 -1872 1063 -1871
rect 1262 -1872 1263 -1871
rect 19 -1874 20 -1873
rect 75 -1874 76 -1873
rect 100 -1874 101 -1873
rect 114 -1874 115 -1873
rect 128 -1874 129 -1873
rect 936 -1874 937 -1873
rect 968 -1874 969 -1873
rect 975 -1874 976 -1873
rect 1234 -1874 1235 -1873
rect 1395 -1874 1396 -1873
rect 26 -1876 27 -1875
rect 30 -1876 31 -1875
rect 37 -1876 38 -1875
rect 394 -1876 395 -1875
rect 401 -1876 402 -1875
rect 471 -1876 472 -1875
rect 499 -1876 500 -1875
rect 597 -1876 598 -1875
rect 618 -1876 619 -1875
rect 803 -1876 804 -1875
rect 856 -1876 857 -1875
rect 905 -1876 906 -1875
rect 912 -1876 913 -1875
rect 926 -1876 927 -1875
rect 933 -1876 934 -1875
rect 1003 -1876 1004 -1875
rect 1066 -1876 1067 -1875
rect 1234 -1876 1235 -1875
rect 30 -1878 31 -1877
rect 457 -1878 458 -1877
rect 502 -1878 503 -1877
rect 1381 -1878 1382 -1877
rect 37 -1880 38 -1879
rect 1199 -1880 1200 -1879
rect 44 -1882 45 -1881
rect 509 -1882 510 -1881
rect 523 -1882 524 -1881
rect 1206 -1882 1207 -1881
rect 44 -1884 45 -1883
rect 604 -1884 605 -1883
rect 646 -1884 647 -1883
rect 663 -1884 664 -1883
rect 681 -1884 682 -1883
rect 1398 -1884 1399 -1883
rect 51 -1886 52 -1885
rect 212 -1886 213 -1885
rect 219 -1886 220 -1885
rect 401 -1886 402 -1885
rect 527 -1886 528 -1885
rect 597 -1886 598 -1885
rect 604 -1886 605 -1885
rect 1059 -1886 1060 -1885
rect 1199 -1886 1200 -1885
rect 1241 -1886 1242 -1885
rect 58 -1888 59 -1887
rect 856 -1888 857 -1887
rect 884 -1888 885 -1887
rect 1430 -1888 1431 -1887
rect 58 -1890 59 -1889
rect 513 -1890 514 -1889
rect 555 -1890 556 -1889
rect 625 -1890 626 -1889
rect 660 -1890 661 -1889
rect 1157 -1890 1158 -1889
rect 1206 -1890 1207 -1889
rect 1297 -1890 1298 -1889
rect 40 -1892 41 -1891
rect 1157 -1892 1158 -1891
rect 1241 -1892 1242 -1891
rect 1255 -1892 1256 -1891
rect 1297 -1892 1298 -1891
rect 1332 -1892 1333 -1891
rect 61 -1894 62 -1893
rect 261 -1894 262 -1893
rect 282 -1894 283 -1893
rect 408 -1894 409 -1893
rect 513 -1894 514 -1893
rect 723 -1894 724 -1893
rect 726 -1894 727 -1893
rect 1262 -1894 1263 -1893
rect 1332 -1894 1333 -1893
rect 1367 -1894 1368 -1893
rect 79 -1896 80 -1895
rect 212 -1896 213 -1895
rect 219 -1896 220 -1895
rect 352 -1896 353 -1895
rect 355 -1896 356 -1895
rect 975 -1896 976 -1895
rect 996 -1896 997 -1895
rect 1066 -1896 1067 -1895
rect 1122 -1896 1123 -1895
rect 1367 -1896 1368 -1895
rect 79 -1898 80 -1897
rect 142 -1898 143 -1897
rect 170 -1898 171 -1897
rect 642 -1898 643 -1897
rect 688 -1898 689 -1897
rect 1171 -1898 1172 -1897
rect 1255 -1898 1256 -1897
rect 1311 -1898 1312 -1897
rect 89 -1900 90 -1899
rect 646 -1900 647 -1899
rect 660 -1900 661 -1899
rect 688 -1900 689 -1899
rect 691 -1900 692 -1899
rect 1171 -1900 1172 -1899
rect 1311 -1900 1312 -1899
rect 1339 -1900 1340 -1899
rect 121 -1902 122 -1901
rect 499 -1902 500 -1901
rect 625 -1902 626 -1901
rect 709 -1902 710 -1901
rect 737 -1902 738 -1901
rect 996 -1902 997 -1901
rect 1003 -1902 1004 -1901
rect 1073 -1902 1074 -1901
rect 1122 -1902 1123 -1901
rect 1220 -1902 1221 -1901
rect 1339 -1902 1340 -1901
rect 1388 -1902 1389 -1901
rect 121 -1904 122 -1903
rect 506 -1904 507 -1903
rect 702 -1904 703 -1903
rect 719 -1904 720 -1903
rect 737 -1904 738 -1903
rect 807 -1904 808 -1903
rect 870 -1904 871 -1903
rect 884 -1904 885 -1903
rect 926 -1904 927 -1903
rect 1017 -1904 1018 -1903
rect 1038 -1904 1039 -1903
rect 1220 -1904 1221 -1903
rect 1388 -1904 1389 -1903
rect 1416 -1904 1417 -1903
rect 128 -1906 129 -1905
rect 443 -1906 444 -1905
rect 506 -1906 507 -1905
rect 1248 -1906 1249 -1905
rect 135 -1908 136 -1907
rect 1143 -1908 1144 -1907
rect 1248 -1908 1249 -1907
rect 1304 -1908 1305 -1907
rect 135 -1910 136 -1909
rect 149 -1910 150 -1909
rect 170 -1910 171 -1909
rect 1374 -1910 1375 -1909
rect 142 -1912 143 -1911
rect 296 -1912 297 -1911
rect 338 -1912 339 -1911
rect 1017 -1912 1018 -1911
rect 1038 -1912 1039 -1911
rect 1108 -1912 1109 -1911
rect 1143 -1912 1144 -1911
rect 1192 -1912 1193 -1911
rect 1374 -1912 1375 -1911
rect 1409 -1912 1410 -1911
rect 149 -1914 150 -1913
rect 667 -1914 668 -1913
rect 716 -1914 717 -1913
rect 1304 -1914 1305 -1913
rect 205 -1916 206 -1915
rect 569 -1916 570 -1915
rect 611 -1916 612 -1915
rect 702 -1916 703 -1915
rect 716 -1916 717 -1915
rect 758 -1916 759 -1915
rect 772 -1916 773 -1915
rect 828 -1916 829 -1915
rect 870 -1916 871 -1915
rect 891 -1916 892 -1915
rect 1059 -1916 1060 -1915
rect 1129 -1916 1130 -1915
rect 1192 -1916 1193 -1915
rect 1276 -1916 1277 -1915
rect 205 -1918 206 -1917
rect 331 -1918 332 -1917
rect 338 -1918 339 -1917
rect 366 -1918 367 -1917
rect 387 -1918 388 -1917
rect 663 -1918 664 -1917
rect 744 -1918 745 -1917
rect 821 -1918 822 -1917
rect 828 -1918 829 -1917
rect 863 -1918 864 -1917
rect 891 -1918 892 -1917
rect 947 -1918 948 -1917
rect 1108 -1918 1109 -1917
rect 1402 -1918 1403 -1917
rect 93 -1920 94 -1919
rect 863 -1920 864 -1919
rect 898 -1920 899 -1919
rect 947 -1920 948 -1919
rect 1024 -1920 1025 -1919
rect 1402 -1920 1403 -1919
rect 93 -1922 94 -1921
rect 198 -1922 199 -1921
rect 233 -1922 234 -1921
rect 429 -1922 430 -1921
rect 492 -1922 493 -1921
rect 667 -1922 668 -1921
rect 751 -1922 752 -1921
rect 1073 -1922 1074 -1921
rect 1129 -1922 1130 -1921
rect 1325 -1922 1326 -1921
rect 198 -1924 199 -1923
rect 786 -1924 787 -1923
rect 800 -1924 801 -1923
rect 954 -1924 955 -1923
rect 1024 -1924 1025 -1923
rect 1087 -1924 1088 -1923
rect 1276 -1924 1277 -1923
rect 1318 -1924 1319 -1923
rect 1325 -1924 1326 -1923
rect 1353 -1924 1354 -1923
rect 86 -1926 87 -1925
rect 1353 -1926 1354 -1925
rect 86 -1928 87 -1927
rect 348 -1928 349 -1927
rect 352 -1928 353 -1927
rect 387 -1928 388 -1927
rect 408 -1928 409 -1927
rect 527 -1928 528 -1927
rect 569 -1928 570 -1927
rect 576 -1928 577 -1927
rect 611 -1928 612 -1927
rect 709 -1928 710 -1927
rect 723 -1928 724 -1927
rect 786 -1928 787 -1927
rect 800 -1928 801 -1927
rect 940 -1928 941 -1927
rect 954 -1928 955 -1927
rect 1045 -1928 1046 -1927
rect 1087 -1928 1088 -1927
rect 1269 -1928 1270 -1927
rect 1318 -1928 1319 -1927
rect 1346 -1928 1347 -1927
rect 138 -1930 139 -1929
rect 1045 -1930 1046 -1929
rect 1346 -1930 1347 -1929
rect 1360 -1930 1361 -1929
rect 233 -1932 234 -1931
rect 632 -1932 633 -1931
rect 653 -1932 654 -1931
rect 898 -1932 899 -1931
rect 940 -1932 941 -1931
rect 1115 -1932 1116 -1931
rect 240 -1934 241 -1933
rect 684 -1934 685 -1933
rect 754 -1934 755 -1933
rect 877 -1934 878 -1933
rect 989 -1934 990 -1933
rect 1360 -1934 1361 -1933
rect 240 -1936 241 -1935
rect 422 -1936 423 -1935
rect 429 -1936 430 -1935
rect 908 -1936 909 -1935
rect 989 -1936 990 -1935
rect 1052 -1936 1053 -1935
rect 1115 -1936 1116 -1935
rect 1185 -1936 1186 -1935
rect 191 -1938 192 -1937
rect 422 -1938 423 -1937
rect 464 -1938 465 -1937
rect 492 -1938 493 -1937
rect 520 -1938 521 -1937
rect 576 -1938 577 -1937
rect 674 -1938 675 -1937
rect 754 -1938 755 -1937
rect 758 -1938 759 -1937
rect 765 -1938 766 -1937
rect 782 -1938 783 -1937
rect 1101 -1938 1102 -1937
rect 1150 -1938 1151 -1937
rect 1185 -1938 1186 -1937
rect 72 -1940 73 -1939
rect 191 -1940 192 -1939
rect 247 -1940 248 -1939
rect 394 -1940 395 -1939
rect 464 -1940 465 -1939
rect 793 -1940 794 -1939
rect 807 -1940 808 -1939
rect 1283 -1940 1284 -1939
rect 72 -1942 73 -1941
rect 173 -1942 174 -1941
rect 268 -1942 269 -1941
rect 443 -1942 444 -1941
rect 485 -1942 486 -1941
rect 793 -1942 794 -1941
rect 821 -1942 822 -1941
rect 849 -1942 850 -1941
rect 1010 -1942 1011 -1941
rect 1150 -1942 1151 -1941
rect 107 -1944 108 -1943
rect 247 -1944 248 -1943
rect 268 -1944 269 -1943
rect 275 -1944 276 -1943
rect 289 -1944 290 -1943
rect 632 -1944 633 -1943
rect 765 -1944 766 -1943
rect 814 -1944 815 -1943
rect 835 -1944 836 -1943
rect 877 -1944 878 -1943
rect 1010 -1944 1011 -1943
rect 1080 -1944 1081 -1943
rect 1101 -1944 1102 -1943
rect 1178 -1944 1179 -1943
rect 16 -1946 17 -1945
rect 107 -1946 108 -1945
rect 163 -1946 164 -1945
rect 289 -1946 290 -1945
rect 296 -1946 297 -1945
rect 541 -1946 542 -1945
rect 572 -1946 573 -1945
rect 814 -1946 815 -1945
rect 835 -1946 836 -1945
rect 842 -1946 843 -1945
rect 1052 -1946 1053 -1945
rect 1094 -1946 1095 -1945
rect 1178 -1946 1179 -1945
rect 1227 -1946 1228 -1945
rect 16 -1948 17 -1947
rect 23 -1948 24 -1947
rect 163 -1948 164 -1947
rect 593 -1948 594 -1947
rect 842 -1948 843 -1947
rect 961 -1948 962 -1947
rect 1080 -1948 1081 -1947
rect 1136 -1948 1137 -1947
rect 23 -1950 24 -1949
rect 1213 -1950 1214 -1949
rect 229 -1952 230 -1951
rect 275 -1952 276 -1951
rect 310 -1952 311 -1951
rect 485 -1952 486 -1951
rect 579 -1952 580 -1951
rect 674 -1952 675 -1951
rect 705 -1952 706 -1951
rect 1136 -1952 1137 -1951
rect 1213 -1952 1214 -1951
rect 1290 -1952 1291 -1951
rect 310 -1954 311 -1953
rect 324 -1954 325 -1953
rect 331 -1954 332 -1953
rect 548 -1954 549 -1953
rect 887 -1954 888 -1953
rect 1290 -1954 1291 -1953
rect 65 -1956 66 -1955
rect 324 -1956 325 -1955
rect 345 -1956 346 -1955
rect 516 -1956 517 -1955
rect 548 -1956 549 -1955
rect 562 -1956 563 -1955
rect 961 -1956 962 -1955
rect 982 -1956 983 -1955
rect 1094 -1956 1095 -1955
rect 1164 -1956 1165 -1955
rect 65 -1958 66 -1957
rect 114 -1958 115 -1957
rect 317 -1958 318 -1957
rect 562 -1958 563 -1957
rect 779 -1958 780 -1957
rect 1164 -1958 1165 -1957
rect 317 -1960 318 -1959
rect 436 -1960 437 -1959
rect 478 -1960 479 -1959
rect 541 -1960 542 -1959
rect 681 -1960 682 -1959
rect 779 -1960 780 -1959
rect 982 -1960 983 -1959
rect 1031 -1960 1032 -1959
rect 359 -1962 360 -1961
rect 457 -1962 458 -1961
rect 919 -1962 920 -1961
rect 1031 -1962 1032 -1961
rect 359 -1964 360 -1963
rect 450 -1964 451 -1963
rect 590 -1964 591 -1963
rect 919 -1964 920 -1963
rect 177 -1966 178 -1965
rect 450 -1966 451 -1965
rect 583 -1966 584 -1965
rect 590 -1966 591 -1965
rect 177 -1968 178 -1967
rect 226 -1968 227 -1967
rect 366 -1968 367 -1967
rect 639 -1968 640 -1967
rect 184 -1970 185 -1969
rect 226 -1970 227 -1969
rect 373 -1970 374 -1969
rect 1269 -1970 1270 -1969
rect 68 -1972 69 -1971
rect 184 -1972 185 -1971
rect 380 -1972 381 -1971
rect 520 -1972 521 -1971
rect 583 -1972 584 -1971
rect 1227 -1972 1228 -1971
rect 156 -1974 157 -1973
rect 380 -1974 381 -1973
rect 415 -1974 416 -1973
rect 478 -1974 479 -1973
rect 639 -1974 640 -1973
rect 653 -1974 654 -1973
rect 5 -1976 6 -1975
rect 415 -1976 416 -1975
rect 436 -1976 437 -1975
rect 852 -1976 853 -1975
rect 156 -1978 157 -1977
rect 695 -1978 696 -1977
rect 695 -1980 696 -1979
rect 730 -1980 731 -1979
rect 534 -1982 535 -1981
rect 730 -1982 731 -1981
rect 411 -1984 412 -1983
rect 534 -1984 535 -1983
rect 2 -1995 3 -1994
rect 37 -1995 38 -1994
rect 51 -1995 52 -1994
rect 660 -1995 661 -1994
rect 663 -1995 664 -1994
rect 996 -1995 997 -1994
rect 1139 -1995 1140 -1994
rect 1367 -1995 1368 -1994
rect 5 -1997 6 -1996
rect 191 -1997 192 -1996
rect 205 -1997 206 -1996
rect 320 -1997 321 -1996
rect 324 -1997 325 -1996
rect 376 -1997 377 -1996
rect 408 -1997 409 -1996
rect 1262 -1997 1263 -1996
rect 37 -1999 38 -1998
rect 338 -1999 339 -1998
rect 408 -1999 409 -1998
rect 541 -1999 542 -1998
rect 579 -1999 580 -1998
rect 1185 -1999 1186 -1998
rect 1262 -1999 1263 -1998
rect 1283 -1999 1284 -1998
rect 51 -2001 52 -2000
rect 261 -2001 262 -2000
rect 268 -2001 269 -2000
rect 355 -2001 356 -2000
rect 373 -2001 374 -2000
rect 1185 -2001 1186 -2000
rect 1283 -2001 1284 -2000
rect 1325 -2001 1326 -2000
rect 58 -2003 59 -2002
rect 488 -2003 489 -2002
rect 502 -2003 503 -2002
rect 1304 -2003 1305 -2002
rect 1325 -2003 1326 -2002
rect 1388 -2003 1389 -2002
rect 58 -2005 59 -2004
rect 247 -2005 248 -2004
rect 261 -2005 262 -2004
rect 387 -2005 388 -2004
rect 411 -2005 412 -2004
rect 1234 -2005 1235 -2004
rect 65 -2007 66 -2006
rect 289 -2007 290 -2006
rect 334 -2007 335 -2006
rect 1276 -2007 1277 -2006
rect 65 -2009 66 -2008
rect 303 -2009 304 -2008
rect 338 -2009 339 -2008
rect 394 -2009 395 -2008
rect 415 -2009 416 -2008
rect 541 -2009 542 -2008
rect 614 -2009 615 -2008
rect 1241 -2009 1242 -2008
rect 68 -2011 69 -2010
rect 324 -2011 325 -2010
rect 373 -2011 374 -2010
rect 478 -2011 479 -2010
rect 513 -2011 514 -2010
rect 1290 -2011 1291 -2010
rect 72 -2013 73 -2012
rect 1227 -2013 1228 -2012
rect 1290 -2013 1291 -2012
rect 1332 -2013 1333 -2012
rect 72 -2015 73 -2014
rect 331 -2015 332 -2014
rect 387 -2015 388 -2014
rect 485 -2015 486 -2014
rect 513 -2015 514 -2014
rect 625 -2015 626 -2014
rect 639 -2015 640 -2014
rect 1080 -2015 1081 -2014
rect 1108 -2015 1109 -2014
rect 1304 -2015 1305 -2014
rect 93 -2017 94 -2016
rect 205 -2017 206 -2016
rect 268 -2017 269 -2016
rect 429 -2017 430 -2016
rect 453 -2017 454 -2016
rect 1241 -2017 1242 -2016
rect 93 -2019 94 -2018
rect 639 -2019 640 -2018
rect 646 -2019 647 -2018
rect 660 -2019 661 -2018
rect 691 -2019 692 -2018
rect 1360 -2019 1361 -2018
rect 96 -2021 97 -2020
rect 100 -2021 101 -2020
rect 107 -2021 108 -2020
rect 247 -2021 248 -2020
rect 289 -2021 290 -2020
rect 436 -2021 437 -2020
rect 478 -2021 479 -2020
rect 527 -2021 528 -2020
rect 604 -2021 605 -2020
rect 625 -2021 626 -2020
rect 646 -2021 647 -2020
rect 681 -2021 682 -2020
rect 705 -2021 706 -2020
rect 772 -2021 773 -2020
rect 782 -2021 783 -2020
rect 821 -2021 822 -2020
rect 849 -2021 850 -2020
rect 933 -2021 934 -2020
rect 947 -2021 948 -2020
rect 1143 -2021 1144 -2020
rect 1213 -2021 1214 -2020
rect 1276 -2021 1277 -2020
rect 100 -2023 101 -2022
rect 173 -2023 174 -2022
rect 177 -2023 178 -2022
rect 331 -2023 332 -2022
rect 415 -2023 416 -2022
rect 492 -2023 493 -2022
rect 516 -2023 517 -2022
rect 765 -2023 766 -2022
rect 807 -2023 808 -2022
rect 1045 -2023 1046 -2022
rect 1059 -2023 1060 -2022
rect 1080 -2023 1081 -2022
rect 1129 -2023 1130 -2022
rect 1234 -2023 1235 -2022
rect 121 -2025 122 -2024
rect 492 -2025 493 -2024
rect 499 -2025 500 -2024
rect 807 -2025 808 -2024
rect 821 -2025 822 -2024
rect 1199 -2025 1200 -2024
rect 1206 -2025 1207 -2024
rect 1213 -2025 1214 -2024
rect 1227 -2025 1228 -2024
rect 1255 -2025 1256 -2024
rect 23 -2027 24 -2026
rect 121 -2027 122 -2026
rect 128 -2027 129 -2026
rect 681 -2027 682 -2026
rect 726 -2027 727 -2026
rect 1402 -2027 1403 -2026
rect 16 -2029 17 -2028
rect 128 -2029 129 -2028
rect 131 -2029 132 -2028
rect 394 -2029 395 -2028
rect 422 -2029 423 -2028
rect 509 -2029 510 -2028
rect 520 -2029 521 -2028
rect 590 -2029 591 -2028
rect 621 -2029 622 -2028
rect 1353 -2029 1354 -2028
rect 16 -2031 17 -2030
rect 240 -2031 241 -2030
rect 296 -2031 297 -2030
rect 499 -2031 500 -2030
rect 520 -2031 521 -2030
rect 817 -2031 818 -2030
rect 849 -2031 850 -2030
rect 856 -2031 857 -2030
rect 912 -2031 913 -2030
rect 1108 -2031 1109 -2030
rect 1129 -2031 1130 -2030
rect 1136 -2031 1137 -2030
rect 1143 -2031 1144 -2030
rect 1164 -2031 1165 -2030
rect 1199 -2031 1200 -2030
rect 1220 -2031 1221 -2030
rect 23 -2033 24 -2032
rect 156 -2033 157 -2032
rect 163 -2033 164 -2032
rect 226 -2033 227 -2032
rect 296 -2033 297 -2032
rect 611 -2033 612 -2032
rect 730 -2033 731 -2032
rect 733 -2033 734 -2032
rect 737 -2033 738 -2032
rect 772 -2033 773 -2032
rect 779 -2033 780 -2032
rect 1164 -2033 1165 -2032
rect 1206 -2033 1207 -2032
rect 1318 -2033 1319 -2032
rect 9 -2035 10 -2034
rect 163 -2035 164 -2034
rect 166 -2035 167 -2034
rect 1017 -2035 1018 -2034
rect 1059 -2035 1060 -2034
rect 1094 -2035 1095 -2034
rect 1220 -2035 1221 -2034
rect 1248 -2035 1249 -2034
rect 1318 -2035 1319 -2034
rect 1381 -2035 1382 -2034
rect 9 -2037 10 -2036
rect 1255 -2037 1256 -2036
rect 135 -2039 136 -2038
rect 156 -2039 157 -2038
rect 173 -2039 174 -2038
rect 212 -2039 213 -2038
rect 219 -2039 220 -2038
rect 240 -2039 241 -2038
rect 303 -2039 304 -2038
rect 310 -2039 311 -2038
rect 422 -2039 423 -2038
rect 450 -2039 451 -2038
rect 527 -2039 528 -2038
rect 548 -2039 549 -2038
rect 555 -2039 556 -2038
rect 604 -2039 605 -2038
rect 716 -2039 717 -2038
rect 737 -2039 738 -2038
rect 754 -2039 755 -2038
rect 898 -2039 899 -2038
rect 933 -2039 934 -2038
rect 992 -2039 993 -2038
rect 996 -2039 997 -2038
rect 1122 -2039 1123 -2038
rect 1248 -2039 1249 -2038
rect 1269 -2039 1270 -2038
rect 110 -2041 111 -2040
rect 212 -2041 213 -2040
rect 219 -2041 220 -2040
rect 534 -2041 535 -2040
rect 548 -2041 549 -2040
rect 782 -2041 783 -2040
rect 842 -2041 843 -2040
rect 912 -2041 913 -2040
rect 968 -2041 969 -2040
rect 1045 -2041 1046 -2040
rect 1094 -2041 1095 -2040
rect 1192 -2041 1193 -2040
rect 1269 -2041 1270 -2040
rect 1311 -2041 1312 -2040
rect 135 -2043 136 -2042
rect 670 -2043 671 -2042
rect 730 -2043 731 -2042
rect 800 -2043 801 -2042
rect 828 -2043 829 -2042
rect 842 -2043 843 -2042
rect 852 -2043 853 -2042
rect 905 -2043 906 -2042
rect 971 -2043 972 -2042
rect 1297 -2043 1298 -2042
rect 1311 -2043 1312 -2042
rect 1374 -2043 1375 -2042
rect 142 -2045 143 -2044
rect 310 -2045 311 -2044
rect 429 -2045 430 -2044
rect 824 -2045 825 -2044
rect 856 -2045 857 -2044
rect 954 -2045 955 -2044
rect 1017 -2045 1018 -2044
rect 1087 -2045 1088 -2044
rect 1101 -2045 1102 -2044
rect 1192 -2045 1193 -2044
rect 1297 -2045 1298 -2044
rect 1339 -2045 1340 -2044
rect 142 -2047 143 -2046
rect 359 -2047 360 -2046
rect 436 -2047 437 -2046
rect 471 -2047 472 -2046
rect 485 -2047 486 -2046
rect 716 -2047 717 -2046
rect 765 -2047 766 -2046
rect 863 -2047 864 -2046
rect 870 -2047 871 -2046
rect 898 -2047 899 -2046
rect 954 -2047 955 -2046
rect 989 -2047 990 -2046
rect 1073 -2047 1074 -2046
rect 1087 -2047 1088 -2046
rect 1101 -2047 1102 -2046
rect 1115 -2047 1116 -2046
rect 30 -2049 31 -2048
rect 359 -2049 360 -2048
rect 443 -2049 444 -2048
rect 450 -2049 451 -2048
rect 457 -2049 458 -2048
rect 471 -2049 472 -2048
rect 555 -2049 556 -2048
rect 586 -2049 587 -2048
rect 590 -2049 591 -2048
rect 632 -2049 633 -2048
rect 779 -2049 780 -2048
rect 1346 -2049 1347 -2048
rect 30 -2051 31 -2050
rect 40 -2051 41 -2050
rect 170 -2051 171 -2050
rect 443 -2051 444 -2050
rect 457 -2051 458 -2050
rect 464 -2051 465 -2050
rect 569 -2051 570 -2050
rect 611 -2051 612 -2050
rect 786 -2051 787 -2050
rect 800 -2051 801 -2050
rect 863 -2051 864 -2050
rect 894 -2051 895 -2050
rect 1066 -2051 1067 -2050
rect 1073 -2051 1074 -2050
rect 75 -2053 76 -2052
rect 170 -2053 171 -2052
rect 177 -2053 178 -2052
rect 723 -2053 724 -2052
rect 744 -2053 745 -2052
rect 786 -2053 787 -2052
rect 870 -2053 871 -2052
rect 1115 -2053 1116 -2052
rect 191 -2055 192 -2054
rect 618 -2055 619 -2054
rect 674 -2055 675 -2054
rect 723 -2055 724 -2054
rect 733 -2055 734 -2054
rect 744 -2055 745 -2054
rect 891 -2055 892 -2054
rect 905 -2055 906 -2054
rect 149 -2057 150 -2056
rect 618 -2057 619 -2056
rect 674 -2057 675 -2056
rect 695 -2057 696 -2056
rect 149 -2059 150 -2058
rect 1157 -2059 1158 -2058
rect 198 -2061 199 -2060
rect 464 -2061 465 -2060
rect 506 -2061 507 -2060
rect 1066 -2061 1067 -2060
rect 184 -2063 185 -2062
rect 198 -2063 199 -2062
rect 226 -2063 227 -2062
rect 751 -2063 752 -2062
rect 184 -2065 185 -2064
rect 254 -2065 255 -2064
rect 562 -2065 563 -2064
rect 1157 -2065 1158 -2064
rect 229 -2067 230 -2066
rect 506 -2067 507 -2066
rect 562 -2067 563 -2066
rect 975 -2067 976 -2066
rect 233 -2069 234 -2068
rect 534 -2069 535 -2068
rect 569 -2069 570 -2068
rect 667 -2069 668 -2068
rect 695 -2069 696 -2068
rect 793 -2069 794 -2068
rect 975 -2069 976 -2068
rect 982 -2069 983 -2068
rect 86 -2071 87 -2070
rect 233 -2071 234 -2070
rect 254 -2071 255 -2070
rect 282 -2071 283 -2070
rect 576 -2071 577 -2070
rect 632 -2071 633 -2070
rect 667 -2071 668 -2070
rect 1150 -2071 1151 -2070
rect 86 -2073 87 -2072
rect 107 -2073 108 -2072
rect 282 -2073 283 -2072
rect 345 -2073 346 -2072
rect 576 -2073 577 -2072
rect 961 -2073 962 -2072
rect 982 -2073 983 -2072
rect 1395 -2073 1396 -2072
rect 345 -2075 346 -2074
rect 401 -2075 402 -2074
rect 579 -2075 580 -2074
rect 947 -2075 948 -2074
rect 1150 -2075 1151 -2074
rect 1171 -2075 1172 -2074
rect 401 -2077 402 -2076
rect 642 -2077 643 -2076
rect 751 -2077 752 -2076
rect 758 -2077 759 -2076
rect 793 -2077 794 -2076
rect 1003 -2077 1004 -2076
rect 1171 -2077 1172 -2076
rect 1178 -2077 1179 -2076
rect 597 -2079 598 -2078
rect 828 -2079 829 -2078
rect 835 -2079 836 -2078
rect 1003 -2079 1004 -2078
rect 523 -2081 524 -2080
rect 597 -2081 598 -2080
rect 688 -2081 689 -2080
rect 758 -2081 759 -2080
rect 814 -2081 815 -2080
rect 835 -2081 836 -2080
rect 926 -2081 927 -2080
rect 961 -2081 962 -2080
rect 583 -2083 584 -2082
rect 688 -2083 689 -2082
rect 709 -2083 710 -2082
rect 1178 -2083 1179 -2082
rect 380 -2085 381 -2084
rect 709 -2085 710 -2084
rect 814 -2085 815 -2084
rect 1052 -2085 1053 -2084
rect 44 -2087 45 -2086
rect 380 -2087 381 -2086
rect 583 -2087 584 -2086
rect 653 -2087 654 -2086
rect 919 -2087 920 -2086
rect 926 -2087 927 -2086
rect 940 -2087 941 -2086
rect 1052 -2087 1053 -2086
rect 2 -2089 3 -2088
rect 653 -2089 654 -2088
rect 940 -2089 941 -2088
rect 1038 -2089 1039 -2088
rect 44 -2091 45 -2090
rect 79 -2091 80 -2090
rect 352 -2091 353 -2090
rect 919 -2091 920 -2090
rect 968 -2091 969 -2090
rect 1038 -2091 1039 -2090
rect 79 -2093 80 -2092
rect 317 -2093 318 -2092
rect 275 -2095 276 -2094
rect 352 -2095 353 -2094
rect 275 -2097 276 -2096
rect 366 -2097 367 -2096
rect 317 -2099 318 -2098
rect 1122 -2099 1123 -2098
rect 366 -2101 367 -2100
rect 702 -2101 703 -2100
rect 702 -2103 703 -2102
rect 810 -2103 811 -2102
rect 9 -2114 10 -2113
rect 44 -2114 45 -2113
rect 51 -2114 52 -2113
rect 667 -2114 668 -2113
rect 765 -2114 766 -2113
rect 768 -2114 769 -2113
rect 793 -2114 794 -2113
rect 891 -2114 892 -2113
rect 936 -2114 937 -2113
rect 975 -2114 976 -2113
rect 989 -2114 990 -2113
rect 1045 -2114 1046 -2113
rect 1115 -2114 1116 -2113
rect 1262 -2114 1263 -2113
rect 9 -2116 10 -2115
rect 471 -2116 472 -2115
rect 478 -2116 479 -2115
rect 691 -2116 692 -2115
rect 695 -2116 696 -2115
rect 793 -2116 794 -2115
rect 814 -2116 815 -2115
rect 905 -2116 906 -2115
rect 968 -2116 969 -2115
rect 1115 -2116 1116 -2115
rect 1118 -2116 1119 -2115
rect 1213 -2116 1214 -2115
rect 1262 -2116 1263 -2115
rect 1283 -2116 1284 -2115
rect 30 -2118 31 -2117
rect 44 -2118 45 -2117
rect 51 -2118 52 -2117
rect 660 -2118 661 -2117
rect 667 -2118 668 -2117
rect 737 -2118 738 -2117
rect 765 -2118 766 -2117
rect 835 -2118 836 -2117
rect 891 -2118 892 -2117
rect 1052 -2118 1053 -2117
rect 1139 -2118 1140 -2117
rect 1276 -2118 1277 -2117
rect 75 -2120 76 -2119
rect 709 -2120 710 -2119
rect 814 -2120 815 -2119
rect 898 -2120 899 -2119
rect 905 -2120 906 -2119
rect 954 -2120 955 -2119
rect 985 -2120 986 -2119
rect 1283 -2120 1284 -2119
rect 107 -2122 108 -2121
rect 1192 -2122 1193 -2121
rect 1213 -2122 1214 -2121
rect 1241 -2122 1242 -2121
rect 1276 -2122 1277 -2121
rect 1290 -2122 1291 -2121
rect 107 -2124 108 -2123
rect 411 -2124 412 -2123
rect 450 -2124 451 -2123
rect 1080 -2124 1081 -2123
rect 1192 -2124 1193 -2123
rect 1220 -2124 1221 -2123
rect 1241 -2124 1242 -2123
rect 1255 -2124 1256 -2123
rect 1290 -2124 1291 -2123
rect 1297 -2124 1298 -2123
rect 40 -2126 41 -2125
rect 1220 -2126 1221 -2125
rect 1297 -2126 1298 -2125
rect 1318 -2126 1319 -2125
rect 110 -2128 111 -2127
rect 268 -2128 269 -2127
rect 320 -2128 321 -2127
rect 485 -2128 486 -2127
rect 488 -2128 489 -2127
rect 898 -2128 899 -2127
rect 989 -2128 990 -2127
rect 1010 -2128 1011 -2127
rect 1045 -2128 1046 -2127
rect 1087 -2128 1088 -2127
rect 1206 -2128 1207 -2127
rect 1255 -2128 1256 -2127
rect 131 -2130 132 -2129
rect 156 -2130 157 -2129
rect 170 -2130 171 -2129
rect 177 -2130 178 -2129
rect 184 -2130 185 -2129
rect 334 -2130 335 -2129
rect 345 -2130 346 -2129
rect 555 -2130 556 -2129
rect 579 -2130 580 -2129
rect 681 -2130 682 -2129
rect 695 -2130 696 -2129
rect 982 -2130 983 -2129
rect 992 -2130 993 -2129
rect 1311 -2130 1312 -2129
rect 37 -2132 38 -2131
rect 184 -2132 185 -2131
rect 191 -2132 192 -2131
rect 677 -2132 678 -2131
rect 821 -2132 822 -2131
rect 849 -2132 850 -2131
rect 856 -2132 857 -2131
rect 954 -2132 955 -2131
rect 996 -2132 997 -2131
rect 1087 -2132 1088 -2131
rect 1206 -2132 1207 -2131
rect 1234 -2132 1235 -2131
rect 79 -2134 80 -2133
rect 177 -2134 178 -2133
rect 191 -2134 192 -2133
rect 317 -2134 318 -2133
rect 331 -2134 332 -2133
rect 975 -2134 976 -2133
rect 996 -2134 997 -2133
rect 1031 -2134 1032 -2133
rect 1080 -2134 1081 -2133
rect 1122 -2134 1123 -2133
rect 79 -2136 80 -2135
rect 541 -2136 542 -2135
rect 555 -2136 556 -2135
rect 653 -2136 654 -2135
rect 660 -2136 661 -2135
rect 730 -2136 731 -2135
rect 849 -2136 850 -2135
rect 884 -2136 885 -2135
rect 940 -2136 941 -2135
rect 1010 -2136 1011 -2135
rect 1031 -2136 1032 -2135
rect 1038 -2136 1039 -2135
rect 138 -2138 139 -2137
rect 156 -2138 157 -2137
rect 163 -2138 164 -2137
rect 982 -2138 983 -2137
rect 1003 -2138 1004 -2137
rect 1311 -2138 1312 -2137
rect 170 -2140 171 -2139
rect 621 -2140 622 -2139
rect 628 -2140 629 -2139
rect 1234 -2140 1235 -2139
rect 205 -2142 206 -2141
rect 208 -2142 209 -2141
rect 219 -2142 220 -2141
rect 971 -2142 972 -2141
rect 1003 -2142 1004 -2141
rect 1024 -2142 1025 -2141
rect 1038 -2142 1039 -2141
rect 1094 -2142 1095 -2141
rect 205 -2144 206 -2143
rect 233 -2144 234 -2143
rect 247 -2144 248 -2143
rect 471 -2144 472 -2143
rect 478 -2144 479 -2143
rect 639 -2144 640 -2143
rect 649 -2144 650 -2143
rect 744 -2144 745 -2143
rect 884 -2144 885 -2143
rect 919 -2144 920 -2143
rect 1094 -2144 1095 -2143
rect 1129 -2144 1130 -2143
rect 247 -2146 248 -2145
rect 299 -2146 300 -2145
rect 317 -2146 318 -2145
rect 338 -2146 339 -2145
rect 352 -2146 353 -2145
rect 425 -2146 426 -2145
rect 450 -2146 451 -2145
rect 782 -2146 783 -2145
rect 1129 -2146 1130 -2145
rect 1164 -2146 1165 -2145
rect 5 -2148 6 -2147
rect 352 -2148 353 -2147
rect 373 -2148 374 -2147
rect 681 -2148 682 -2147
rect 702 -2148 703 -2147
rect 856 -2148 857 -2147
rect 1164 -2148 1165 -2147
rect 1185 -2148 1186 -2147
rect 72 -2150 73 -2149
rect 338 -2150 339 -2149
rect 394 -2150 395 -2149
rect 968 -2150 969 -2149
rect 1185 -2150 1186 -2149
rect 1199 -2150 1200 -2149
rect 72 -2152 73 -2151
rect 149 -2152 150 -2151
rect 254 -2152 255 -2151
rect 348 -2152 349 -2151
rect 394 -2152 395 -2151
rect 422 -2152 423 -2151
rect 464 -2152 465 -2151
rect 709 -2152 710 -2151
rect 730 -2152 731 -2151
rect 824 -2152 825 -2151
rect 1199 -2152 1200 -2151
rect 1227 -2152 1228 -2151
rect 2 -2154 3 -2153
rect 149 -2154 150 -2153
rect 261 -2154 262 -2153
rect 268 -2154 269 -2153
rect 310 -2154 311 -2153
rect 373 -2154 374 -2153
rect 397 -2154 398 -2153
rect 453 -2154 454 -2153
rect 464 -2154 465 -2153
rect 530 -2154 531 -2153
rect 541 -2154 542 -2153
rect 590 -2154 591 -2153
rect 597 -2154 598 -2153
rect 737 -2154 738 -2153
rect 744 -2154 745 -2153
rect 947 -2154 948 -2153
rect 1227 -2154 1228 -2153
rect 1248 -2154 1249 -2153
rect 65 -2156 66 -2155
rect 254 -2156 255 -2155
rect 261 -2156 262 -2155
rect 275 -2156 276 -2155
rect 296 -2156 297 -2155
rect 310 -2156 311 -2155
rect 404 -2156 405 -2155
rect 688 -2156 689 -2155
rect 702 -2156 703 -2155
rect 723 -2156 724 -2155
rect 768 -2156 769 -2155
rect 835 -2156 836 -2155
rect 1248 -2156 1249 -2155
rect 1269 -2156 1270 -2155
rect 65 -2158 66 -2157
rect 86 -2158 87 -2157
rect 275 -2158 276 -2157
rect 303 -2158 304 -2157
rect 453 -2158 454 -2157
rect 807 -2158 808 -2157
rect 1269 -2158 1270 -2157
rect 1304 -2158 1305 -2157
rect 86 -2160 87 -2159
rect 226 -2160 227 -2159
rect 240 -2160 241 -2159
rect 303 -2160 304 -2159
rect 485 -2160 486 -2159
rect 527 -2160 528 -2159
rect 548 -2160 549 -2159
rect 947 -2160 948 -2159
rect 1304 -2160 1305 -2159
rect 1325 -2160 1326 -2159
rect 198 -2162 199 -2161
rect 226 -2162 227 -2161
rect 240 -2162 241 -2161
rect 359 -2162 360 -2161
rect 443 -2162 444 -2161
rect 548 -2162 549 -2161
rect 590 -2162 591 -2161
rect 716 -2162 717 -2161
rect 723 -2162 724 -2161
rect 758 -2162 759 -2161
rect 772 -2162 773 -2161
rect 919 -2162 920 -2161
rect 198 -2164 199 -2163
rect 387 -2164 388 -2163
rect 436 -2164 437 -2163
rect 443 -2164 444 -2163
rect 499 -2164 500 -2163
rect 1178 -2164 1179 -2163
rect 128 -2166 129 -2165
rect 1178 -2166 1179 -2165
rect 114 -2168 115 -2167
rect 128 -2168 129 -2167
rect 219 -2168 220 -2167
rect 527 -2168 528 -2167
rect 576 -2168 577 -2167
rect 772 -2168 773 -2167
rect 807 -2168 808 -2167
rect 1122 -2168 1123 -2167
rect 296 -2170 297 -2169
rect 331 -2170 332 -2169
rect 359 -2170 360 -2169
rect 894 -2170 895 -2169
rect 324 -2172 325 -2171
rect 387 -2172 388 -2171
rect 415 -2172 416 -2171
rect 436 -2172 437 -2171
rect 499 -2172 500 -2171
rect 810 -2172 811 -2171
rect 212 -2174 213 -2173
rect 415 -2174 416 -2173
rect 502 -2174 503 -2173
rect 779 -2174 780 -2173
rect 212 -2176 213 -2175
rect 492 -2176 493 -2175
rect 520 -2176 521 -2175
rect 639 -2176 640 -2175
rect 653 -2176 654 -2175
rect 817 -2176 818 -2175
rect 324 -2178 325 -2177
rect 401 -2178 402 -2177
rect 492 -2178 493 -2177
rect 926 -2178 927 -2177
rect 401 -2180 402 -2179
rect 1024 -2180 1025 -2179
rect 523 -2182 524 -2181
rect 940 -2182 941 -2181
rect 576 -2184 577 -2183
rect 674 -2184 675 -2183
rect 716 -2184 717 -2183
rect 751 -2184 752 -2183
rect 758 -2184 759 -2183
rect 786 -2184 787 -2183
rect 597 -2186 598 -2185
rect 618 -2186 619 -2185
rect 621 -2186 622 -2185
rect 828 -2186 829 -2185
rect 506 -2188 507 -2187
rect 618 -2188 619 -2187
rect 632 -2188 633 -2187
rect 926 -2188 927 -2187
rect 93 -2190 94 -2189
rect 506 -2190 507 -2189
rect 611 -2190 612 -2189
rect 688 -2190 689 -2189
rect 751 -2190 752 -2189
rect 800 -2190 801 -2189
rect 828 -2190 829 -2189
rect 863 -2190 864 -2189
rect 93 -2192 94 -2191
rect 282 -2192 283 -2191
rect 583 -2192 584 -2191
rect 611 -2192 612 -2191
rect 786 -2192 787 -2191
rect 1136 -2192 1137 -2191
rect 117 -2194 118 -2193
rect 632 -2194 633 -2193
rect 800 -2194 801 -2193
rect 842 -2194 843 -2193
rect 863 -2194 864 -2193
rect 912 -2194 913 -2193
rect 1136 -2194 1137 -2193
rect 1157 -2194 1158 -2193
rect 282 -2196 283 -2195
rect 513 -2196 514 -2195
rect 534 -2196 535 -2195
rect 583 -2196 584 -2195
rect 842 -2196 843 -2195
rect 877 -2196 878 -2195
rect 912 -2196 913 -2195
rect 933 -2196 934 -2195
rect 1017 -2196 1018 -2195
rect 1157 -2196 1158 -2195
rect 37 -2198 38 -2197
rect 877 -2198 878 -2197
rect 933 -2198 934 -2197
rect 1108 -2198 1109 -2197
rect 380 -2200 381 -2199
rect 513 -2200 514 -2199
rect 534 -2200 535 -2199
rect 569 -2200 570 -2199
rect 1017 -2200 1018 -2199
rect 1059 -2200 1060 -2199
rect 1108 -2200 1109 -2199
rect 1150 -2200 1151 -2199
rect 135 -2202 136 -2201
rect 380 -2202 381 -2201
rect 520 -2202 521 -2201
rect 1059 -2202 1060 -2201
rect 135 -2204 136 -2203
rect 366 -2204 367 -2203
rect 569 -2204 570 -2203
rect 625 -2204 626 -2203
rect 16 -2206 17 -2205
rect 366 -2206 367 -2205
rect 562 -2206 563 -2205
rect 625 -2206 626 -2205
rect 16 -2208 17 -2207
rect 457 -2208 458 -2207
rect 562 -2208 563 -2207
rect 604 -2208 605 -2207
rect 58 -2210 59 -2209
rect 457 -2210 458 -2209
rect 604 -2210 605 -2209
rect 646 -2210 647 -2209
rect 58 -2212 59 -2211
rect 142 -2212 143 -2211
rect 152 -2212 153 -2211
rect 1150 -2212 1151 -2211
rect 100 -2214 101 -2213
rect 646 -2214 647 -2213
rect 100 -2216 101 -2215
rect 289 -2216 290 -2215
rect 121 -2218 122 -2217
rect 142 -2218 143 -2217
rect 289 -2218 290 -2217
rect 429 -2218 430 -2217
rect 23 -2220 24 -2219
rect 429 -2220 430 -2219
rect 23 -2222 24 -2221
rect 26 -2222 27 -2221
rect 121 -2222 122 -2221
rect 408 -2222 409 -2221
rect 408 -2224 409 -2223
rect 1066 -2224 1067 -2223
rect 1066 -2226 1067 -2225
rect 1101 -2226 1102 -2225
rect 1101 -2228 1102 -2227
rect 1143 -2228 1144 -2227
rect 1143 -2230 1144 -2229
rect 1171 -2230 1172 -2229
rect 1073 -2232 1074 -2231
rect 1171 -2232 1172 -2231
rect 870 -2234 871 -2233
rect 1073 -2234 1074 -2233
rect 870 -2236 871 -2235
rect 1052 -2236 1053 -2235
rect 5 -2247 6 -2246
rect 44 -2247 45 -2246
rect 61 -2247 62 -2246
rect 492 -2247 493 -2246
rect 516 -2247 517 -2246
rect 726 -2247 727 -2246
rect 747 -2247 748 -2246
rect 1087 -2247 1088 -2246
rect 23 -2249 24 -2248
rect 1024 -2249 1025 -2248
rect 1034 -2249 1035 -2248
rect 1290 -2249 1291 -2248
rect 23 -2251 24 -2250
rect 401 -2251 402 -2250
rect 408 -2251 409 -2250
rect 415 -2251 416 -2250
rect 425 -2251 426 -2250
rect 688 -2251 689 -2250
rect 761 -2251 762 -2250
rect 856 -2251 857 -2250
rect 870 -2251 871 -2250
rect 1234 -2251 1235 -2250
rect 33 -2253 34 -2252
rect 198 -2253 199 -2252
rect 205 -2253 206 -2252
rect 338 -2253 339 -2252
rect 387 -2253 388 -2252
rect 523 -2253 524 -2252
rect 527 -2253 528 -2252
rect 737 -2253 738 -2252
rect 810 -2253 811 -2252
rect 961 -2253 962 -2252
rect 982 -2253 983 -2252
rect 1276 -2253 1277 -2252
rect 9 -2255 10 -2254
rect 198 -2255 199 -2254
rect 205 -2255 206 -2254
rect 373 -2255 374 -2254
rect 387 -2255 388 -2254
rect 422 -2255 423 -2254
rect 520 -2255 521 -2254
rect 562 -2255 563 -2254
rect 579 -2255 580 -2254
rect 968 -2255 969 -2254
rect 982 -2255 983 -2254
rect 985 -2255 986 -2254
rect 1024 -2255 1025 -2254
rect 1094 -2255 1095 -2254
rect 9 -2257 10 -2256
rect 359 -2257 360 -2256
rect 411 -2257 412 -2256
rect 464 -2257 465 -2256
rect 527 -2257 528 -2256
rect 933 -2257 934 -2256
rect 961 -2257 962 -2256
rect 1017 -2257 1018 -2256
rect 1094 -2257 1095 -2256
rect 1150 -2257 1151 -2256
rect 37 -2259 38 -2258
rect 975 -2259 976 -2258
rect 1017 -2259 1018 -2258
rect 1080 -2259 1081 -2258
rect 1150 -2259 1151 -2258
rect 1220 -2259 1221 -2258
rect 37 -2261 38 -2260
rect 341 -2261 342 -2260
rect 359 -2261 360 -2260
rect 485 -2261 486 -2260
rect 530 -2261 531 -2260
rect 926 -2261 927 -2260
rect 933 -2261 934 -2260
rect 1059 -2261 1060 -2260
rect 1080 -2261 1081 -2260
rect 1297 -2261 1298 -2260
rect 40 -2263 41 -2262
rect 352 -2263 353 -2262
rect 464 -2263 465 -2262
rect 849 -2263 850 -2262
rect 856 -2263 857 -2262
rect 1010 -2263 1011 -2262
rect 1059 -2263 1060 -2262
rect 1122 -2263 1123 -2262
rect 40 -2265 41 -2264
rect 926 -2265 927 -2264
rect 975 -2265 976 -2264
rect 1269 -2265 1270 -2264
rect 44 -2267 45 -2266
rect 380 -2267 381 -2266
rect 485 -2267 486 -2266
rect 513 -2267 514 -2266
rect 548 -2267 549 -2266
rect 688 -2267 689 -2266
rect 695 -2267 696 -2266
rect 849 -2267 850 -2266
rect 870 -2267 871 -2266
rect 940 -2267 941 -2266
rect 1122 -2267 1123 -2266
rect 1192 -2267 1193 -2266
rect 79 -2269 80 -2268
rect 415 -2269 416 -2268
rect 548 -2269 549 -2268
rect 604 -2269 605 -2268
rect 625 -2269 626 -2268
rect 639 -2269 640 -2268
rect 674 -2269 675 -2268
rect 772 -2269 773 -2268
rect 873 -2269 874 -2268
rect 1031 -2269 1032 -2268
rect 1192 -2269 1193 -2268
rect 1241 -2269 1242 -2268
rect 16 -2271 17 -2270
rect 79 -2271 80 -2270
rect 86 -2271 87 -2270
rect 296 -2271 297 -2270
rect 306 -2271 307 -2270
rect 408 -2271 409 -2270
rect 492 -2271 493 -2270
rect 1031 -2271 1032 -2270
rect 1129 -2271 1130 -2270
rect 1241 -2271 1242 -2270
rect 16 -2273 17 -2272
rect 317 -2273 318 -2272
rect 320 -2273 321 -2272
rect 1234 -2273 1235 -2272
rect 86 -2275 87 -2274
rect 723 -2275 724 -2274
rect 737 -2275 738 -2274
rect 744 -2275 745 -2274
rect 772 -2275 773 -2274
rect 800 -2275 801 -2274
rect 96 -2277 97 -2276
rect 618 -2277 619 -2276
rect 628 -2277 629 -2276
rect 968 -2277 969 -2276
rect 100 -2279 101 -2278
rect 114 -2279 115 -2278
rect 117 -2279 118 -2278
rect 1178 -2279 1179 -2278
rect 100 -2281 101 -2280
rect 345 -2281 346 -2280
rect 352 -2281 353 -2280
rect 478 -2281 479 -2280
rect 513 -2281 514 -2280
rect 1129 -2281 1130 -2280
rect 1178 -2281 1179 -2280
rect 1255 -2281 1256 -2280
rect 114 -2283 115 -2282
rect 191 -2283 192 -2282
rect 240 -2283 241 -2282
rect 520 -2283 521 -2282
rect 558 -2283 559 -2282
rect 681 -2283 682 -2282
rect 695 -2283 696 -2282
rect 793 -2283 794 -2282
rect 800 -2283 801 -2282
rect 814 -2283 815 -2282
rect 121 -2285 122 -2284
rect 744 -2285 745 -2284
rect 793 -2285 794 -2284
rect 810 -2285 811 -2284
rect 814 -2285 815 -2284
rect 877 -2285 878 -2284
rect 121 -2287 122 -2286
rect 450 -2287 451 -2286
rect 555 -2287 556 -2286
rect 681 -2287 682 -2286
rect 877 -2287 878 -2286
rect 947 -2287 948 -2286
rect 149 -2289 150 -2288
rect 919 -2289 920 -2288
rect 947 -2289 948 -2288
rect 1045 -2289 1046 -2288
rect 149 -2291 150 -2290
rect 436 -2291 437 -2290
rect 450 -2291 451 -2290
rect 583 -2291 584 -2290
rect 593 -2291 594 -2290
rect 835 -2291 836 -2290
rect 919 -2291 920 -2290
rect 989 -2291 990 -2290
rect 1045 -2291 1046 -2290
rect 1304 -2291 1305 -2290
rect 152 -2293 153 -2292
rect 807 -2293 808 -2292
rect 989 -2293 990 -2292
rect 1066 -2293 1067 -2292
rect 156 -2295 157 -2294
rect 296 -2295 297 -2294
rect 331 -2295 332 -2294
rect 940 -2295 941 -2294
rect 1066 -2295 1067 -2294
rect 1164 -2295 1165 -2294
rect 2 -2297 3 -2296
rect 331 -2297 332 -2296
rect 341 -2297 342 -2296
rect 457 -2297 458 -2296
rect 562 -2297 563 -2296
rect 660 -2297 661 -2296
rect 677 -2297 678 -2296
rect 1136 -2297 1137 -2296
rect 2 -2299 3 -2298
rect 478 -2299 479 -2298
rect 569 -2299 570 -2298
rect 583 -2299 584 -2298
rect 604 -2299 605 -2298
rect 702 -2299 703 -2298
rect 786 -2299 787 -2298
rect 835 -2299 836 -2298
rect 107 -2301 108 -2300
rect 457 -2301 458 -2300
rect 471 -2301 472 -2300
rect 569 -2301 570 -2300
rect 611 -2301 612 -2300
rect 618 -2301 619 -2300
rect 635 -2301 636 -2300
rect 758 -2301 759 -2300
rect 807 -2301 808 -2300
rect 1003 -2301 1004 -2300
rect 107 -2303 108 -2302
rect 128 -2303 129 -2302
rect 156 -2303 157 -2302
rect 184 -2303 185 -2302
rect 191 -2303 192 -2302
rect 289 -2303 290 -2302
rect 380 -2303 381 -2302
rect 576 -2303 577 -2302
rect 611 -2303 612 -2302
rect 632 -2303 633 -2302
rect 639 -2303 640 -2302
rect 709 -2303 710 -2302
rect 758 -2303 759 -2302
rect 1171 -2303 1172 -2302
rect 75 -2305 76 -2304
rect 632 -2305 633 -2304
rect 646 -2305 647 -2304
rect 1164 -2305 1165 -2304
rect 128 -2307 129 -2306
rect 394 -2307 395 -2306
rect 471 -2307 472 -2306
rect 506 -2307 507 -2306
rect 576 -2307 577 -2306
rect 1220 -2307 1221 -2306
rect 51 -2309 52 -2308
rect 394 -2309 395 -2308
rect 499 -2309 500 -2308
rect 506 -2309 507 -2308
rect 597 -2309 598 -2308
rect 646 -2309 647 -2308
rect 660 -2309 661 -2308
rect 1283 -2309 1284 -2308
rect 51 -2311 52 -2310
rect 138 -2311 139 -2310
rect 163 -2311 164 -2310
rect 289 -2311 290 -2310
rect 338 -2311 339 -2310
rect 1171 -2311 1172 -2310
rect 138 -2313 139 -2312
rect 1087 -2313 1088 -2312
rect 163 -2315 164 -2314
rect 404 -2315 405 -2314
rect 499 -2315 500 -2314
rect 534 -2315 535 -2314
rect 590 -2315 591 -2314
rect 597 -2315 598 -2314
rect 702 -2315 703 -2314
rect 751 -2315 752 -2314
rect 1003 -2315 1004 -2314
rect 1206 -2315 1207 -2314
rect 177 -2317 178 -2316
rect 345 -2317 346 -2316
rect 534 -2317 535 -2316
rect 863 -2317 864 -2316
rect 1206 -2317 1207 -2316
rect 1248 -2317 1249 -2316
rect 170 -2319 171 -2318
rect 177 -2319 178 -2318
rect 184 -2319 185 -2318
rect 233 -2319 234 -2318
rect 254 -2319 255 -2318
rect 373 -2319 374 -2318
rect 590 -2319 591 -2318
rect 1136 -2319 1137 -2318
rect 1248 -2319 1249 -2318
rect 1311 -2319 1312 -2318
rect 93 -2321 94 -2320
rect 254 -2321 255 -2320
rect 261 -2321 262 -2320
rect 401 -2321 402 -2320
rect 709 -2321 710 -2320
rect 716 -2321 717 -2320
rect 751 -2321 752 -2320
rect 842 -2321 843 -2320
rect 863 -2321 864 -2320
rect 954 -2321 955 -2320
rect 65 -2323 66 -2322
rect 93 -2323 94 -2322
rect 170 -2323 171 -2322
rect 317 -2323 318 -2322
rect 397 -2323 398 -2322
rect 842 -2323 843 -2322
rect 954 -2323 955 -2322
rect 1108 -2323 1109 -2322
rect 30 -2325 31 -2324
rect 65 -2325 66 -2324
rect 219 -2325 220 -2324
rect 240 -2325 241 -2324
rect 261 -2325 262 -2324
rect 555 -2325 556 -2324
rect 716 -2325 717 -2324
rect 765 -2325 766 -2324
rect 1108 -2325 1109 -2324
rect 1185 -2325 1186 -2324
rect 30 -2327 31 -2326
rect 425 -2327 426 -2326
rect 1185 -2327 1186 -2326
rect 1227 -2327 1228 -2326
rect 135 -2329 136 -2328
rect 765 -2329 766 -2328
rect 891 -2329 892 -2328
rect 1227 -2329 1228 -2328
rect 135 -2331 136 -2330
rect 366 -2331 367 -2330
rect 397 -2331 398 -2330
rect 730 -2331 731 -2330
rect 891 -2331 892 -2330
rect 996 -2331 997 -2330
rect 219 -2333 220 -2332
rect 324 -2333 325 -2332
rect 366 -2333 367 -2332
rect 541 -2333 542 -2332
rect 730 -2333 731 -2332
rect 821 -2333 822 -2332
rect 996 -2333 997 -2332
rect 1073 -2333 1074 -2332
rect 226 -2335 227 -2334
rect 786 -2335 787 -2334
rect 821 -2335 822 -2334
rect 884 -2335 885 -2334
rect 1073 -2335 1074 -2334
rect 1143 -2335 1144 -2334
rect 142 -2337 143 -2336
rect 226 -2337 227 -2336
rect 233 -2337 234 -2336
rect 268 -2337 269 -2336
rect 282 -2337 283 -2336
rect 663 -2337 664 -2336
rect 779 -2337 780 -2336
rect 884 -2337 885 -2336
rect 1143 -2337 1144 -2336
rect 1199 -2337 1200 -2336
rect 142 -2339 143 -2338
rect 828 -2339 829 -2338
rect 268 -2341 269 -2340
rect 310 -2341 311 -2340
rect 324 -2341 325 -2340
rect 443 -2341 444 -2340
rect 541 -2341 542 -2340
rect 653 -2341 654 -2340
rect 779 -2341 780 -2340
rect 912 -2341 913 -2340
rect 275 -2343 276 -2342
rect 310 -2343 311 -2342
rect 443 -2343 444 -2342
rect 453 -2343 454 -2342
rect 621 -2343 622 -2342
rect 1199 -2343 1200 -2342
rect 275 -2345 276 -2344
rect 429 -2345 430 -2344
rect 653 -2345 654 -2344
rect 667 -2345 668 -2344
rect 828 -2345 829 -2344
rect 898 -2345 899 -2344
rect 912 -2345 913 -2344
rect 1052 -2345 1053 -2344
rect 72 -2347 73 -2346
rect 667 -2347 668 -2346
rect 898 -2347 899 -2346
rect 905 -2347 906 -2346
rect 72 -2349 73 -2348
rect 247 -2349 248 -2348
rect 282 -2349 283 -2348
rect 299 -2349 300 -2348
rect 436 -2349 437 -2348
rect 1052 -2349 1053 -2348
rect 58 -2351 59 -2350
rect 247 -2351 248 -2350
rect 905 -2351 906 -2350
rect 1115 -2351 1116 -2350
rect 58 -2353 59 -2352
rect 1010 -2353 1011 -2352
rect 1038 -2353 1039 -2352
rect 1115 -2353 1116 -2352
rect 212 -2355 213 -2354
rect 429 -2355 430 -2354
rect 1038 -2355 1039 -2354
rect 1101 -2355 1102 -2354
rect 212 -2357 213 -2356
rect 303 -2357 304 -2356
rect 1101 -2357 1102 -2356
rect 1157 -2357 1158 -2356
rect 1157 -2359 1158 -2358
rect 1213 -2359 1214 -2358
rect 1213 -2361 1214 -2360
rect 1262 -2361 1263 -2360
rect 9 -2372 10 -2371
rect 376 -2372 377 -2371
rect 394 -2372 395 -2371
rect 1234 -2372 1235 -2371
rect 23 -2374 24 -2373
rect 341 -2374 342 -2373
rect 352 -2374 353 -2373
rect 436 -2374 437 -2373
rect 446 -2374 447 -2373
rect 779 -2374 780 -2373
rect 796 -2374 797 -2373
rect 954 -2374 955 -2373
rect 1031 -2374 1032 -2373
rect 1073 -2374 1074 -2373
rect 1104 -2374 1105 -2373
rect 1115 -2374 1116 -2373
rect 30 -2376 31 -2375
rect 201 -2376 202 -2375
rect 303 -2376 304 -2375
rect 842 -2376 843 -2375
rect 849 -2376 850 -2375
rect 919 -2376 920 -2375
rect 954 -2376 955 -2375
rect 1045 -2376 1046 -2375
rect 1073 -2376 1074 -2375
rect 1199 -2376 1200 -2375
rect 37 -2378 38 -2377
rect 296 -2378 297 -2377
rect 303 -2378 304 -2377
rect 425 -2378 426 -2377
rect 464 -2378 465 -2377
rect 758 -2378 759 -2377
rect 779 -2378 780 -2377
rect 1010 -2378 1011 -2377
rect 1034 -2378 1035 -2377
rect 1178 -2378 1179 -2377
rect 40 -2380 41 -2379
rect 940 -2380 941 -2379
rect 1010 -2380 1011 -2379
rect 1059 -2380 1060 -2379
rect 54 -2382 55 -2381
rect 254 -2382 255 -2381
rect 320 -2382 321 -2381
rect 786 -2382 787 -2381
rect 807 -2382 808 -2381
rect 1143 -2382 1144 -2381
rect 61 -2384 62 -2383
rect 569 -2384 570 -2383
rect 576 -2384 577 -2383
rect 905 -2384 906 -2383
rect 908 -2384 909 -2383
rect 1220 -2384 1221 -2383
rect 72 -2386 73 -2385
rect 513 -2386 514 -2385
rect 520 -2386 521 -2385
rect 810 -2386 811 -2385
rect 842 -2386 843 -2385
rect 1108 -2386 1109 -2385
rect 72 -2388 73 -2387
rect 170 -2388 171 -2387
rect 184 -2388 185 -2387
rect 306 -2388 307 -2387
rect 338 -2388 339 -2387
rect 443 -2388 444 -2387
rect 485 -2388 486 -2387
rect 849 -2388 850 -2387
rect 898 -2388 899 -2387
rect 1013 -2388 1014 -2387
rect 1059 -2388 1060 -2387
rect 1080 -2388 1081 -2387
rect 79 -2390 80 -2389
rect 149 -2390 150 -2389
rect 163 -2390 164 -2389
rect 296 -2390 297 -2389
rect 359 -2390 360 -2389
rect 362 -2390 363 -2389
rect 366 -2390 367 -2389
rect 516 -2390 517 -2389
rect 520 -2390 521 -2389
rect 593 -2390 594 -2389
rect 614 -2390 615 -2389
rect 863 -2390 864 -2389
rect 898 -2390 899 -2389
rect 1157 -2390 1158 -2389
rect 44 -2392 45 -2391
rect 79 -2392 80 -2391
rect 86 -2392 87 -2391
rect 366 -2392 367 -2391
rect 394 -2392 395 -2391
rect 471 -2392 472 -2391
rect 516 -2392 517 -2391
rect 1164 -2392 1165 -2391
rect 86 -2394 87 -2393
rect 282 -2394 283 -2393
rect 359 -2394 360 -2393
rect 408 -2394 409 -2393
rect 422 -2394 423 -2393
rect 688 -2394 689 -2393
rect 723 -2394 724 -2393
rect 772 -2394 773 -2393
rect 786 -2394 787 -2393
rect 852 -2394 853 -2393
rect 905 -2394 906 -2393
rect 1241 -2394 1242 -2393
rect 93 -2396 94 -2395
rect 422 -2396 423 -2395
rect 450 -2396 451 -2395
rect 863 -2396 864 -2395
rect 919 -2396 920 -2395
rect 996 -2396 997 -2395
rect 1080 -2396 1081 -2395
rect 1136 -2396 1137 -2395
rect 93 -2398 94 -2397
rect 397 -2398 398 -2397
rect 450 -2398 451 -2397
rect 870 -2398 871 -2397
rect 884 -2398 885 -2397
rect 996 -2398 997 -2397
rect 100 -2400 101 -2399
rect 744 -2400 745 -2399
rect 751 -2400 752 -2399
rect 758 -2400 759 -2399
rect 765 -2400 766 -2399
rect 807 -2400 808 -2399
rect 870 -2400 871 -2399
rect 912 -2400 913 -2399
rect 940 -2400 941 -2399
rect 1122 -2400 1123 -2399
rect 100 -2402 101 -2401
rect 142 -2402 143 -2401
rect 184 -2402 185 -2401
rect 562 -2402 563 -2401
rect 569 -2402 570 -2401
rect 625 -2402 626 -2401
rect 635 -2402 636 -2401
rect 702 -2402 703 -2401
rect 709 -2402 710 -2401
rect 884 -2402 885 -2401
rect 912 -2402 913 -2401
rect 1171 -2402 1172 -2401
rect 107 -2404 108 -2403
rect 170 -2404 171 -2403
rect 198 -2404 199 -2403
rect 439 -2404 440 -2403
rect 457 -2404 458 -2403
rect 485 -2404 486 -2403
rect 548 -2404 549 -2403
rect 576 -2404 577 -2403
rect 590 -2404 591 -2403
rect 653 -2404 654 -2403
rect 660 -2404 661 -2403
rect 1227 -2404 1228 -2403
rect 107 -2406 108 -2405
rect 597 -2406 598 -2405
rect 611 -2406 612 -2405
rect 653 -2406 654 -2405
rect 663 -2406 664 -2405
rect 1066 -2406 1067 -2405
rect 58 -2408 59 -2407
rect 597 -2408 598 -2407
rect 646 -2408 647 -2407
rect 744 -2408 745 -2407
rect 751 -2408 752 -2407
rect 891 -2408 892 -2407
rect 961 -2408 962 -2407
rect 1108 -2408 1109 -2407
rect 58 -2410 59 -2409
rect 247 -2410 248 -2409
rect 261 -2410 262 -2409
rect 590 -2410 591 -2409
rect 646 -2410 647 -2409
rect 933 -2410 934 -2409
rect 1066 -2410 1067 -2409
rect 1129 -2410 1130 -2409
rect 121 -2412 122 -2411
rect 254 -2412 255 -2411
rect 261 -2412 262 -2411
rect 506 -2412 507 -2411
rect 555 -2412 556 -2411
rect 730 -2412 731 -2411
rect 765 -2412 766 -2411
rect 975 -2412 976 -2411
rect 1129 -2412 1130 -2411
rect 1248 -2412 1249 -2411
rect 124 -2414 125 -2413
rect 968 -2414 969 -2413
rect 128 -2416 129 -2415
rect 163 -2416 164 -2415
rect 198 -2416 199 -2415
rect 226 -2416 227 -2415
rect 247 -2416 248 -2415
rect 324 -2416 325 -2415
rect 362 -2416 363 -2415
rect 408 -2416 409 -2415
rect 415 -2416 416 -2415
rect 660 -2416 661 -2415
rect 667 -2416 668 -2415
rect 702 -2416 703 -2415
rect 709 -2416 710 -2415
rect 989 -2416 990 -2415
rect 128 -2418 129 -2417
rect 138 -2418 139 -2417
rect 142 -2418 143 -2417
rect 317 -2418 318 -2417
rect 387 -2418 388 -2417
rect 625 -2418 626 -2417
rect 667 -2418 668 -2417
rect 828 -2418 829 -2417
rect 877 -2418 878 -2417
rect 933 -2418 934 -2417
rect 989 -2418 990 -2417
rect 1192 -2418 1193 -2417
rect 131 -2420 132 -2419
rect 548 -2420 549 -2419
rect 558 -2420 559 -2419
rect 639 -2420 640 -2419
rect 674 -2420 675 -2419
rect 975 -2420 976 -2419
rect 1192 -2420 1193 -2419
rect 1206 -2420 1207 -2419
rect 226 -2422 227 -2421
rect 331 -2422 332 -2421
rect 380 -2422 381 -2421
rect 674 -2422 675 -2421
rect 681 -2422 682 -2421
rect 723 -2422 724 -2421
rect 726 -2422 727 -2421
rect 961 -2422 962 -2421
rect 51 -2424 52 -2423
rect 380 -2424 381 -2423
rect 387 -2424 388 -2423
rect 429 -2424 430 -2423
rect 439 -2424 440 -2423
rect 761 -2424 762 -2423
rect 772 -2424 773 -2423
rect 856 -2424 857 -2423
rect 877 -2424 878 -2423
rect 1017 -2424 1018 -2423
rect 275 -2426 276 -2425
rect 726 -2426 727 -2425
rect 814 -2426 815 -2425
rect 891 -2426 892 -2425
rect 1017 -2426 1018 -2425
rect 1213 -2426 1214 -2425
rect 212 -2428 213 -2427
rect 275 -2428 276 -2427
rect 282 -2428 283 -2427
rect 401 -2428 402 -2427
rect 415 -2428 416 -2427
rect 464 -2428 465 -2427
rect 471 -2428 472 -2427
rect 604 -2428 605 -2427
rect 611 -2428 612 -2427
rect 968 -2428 969 -2427
rect 212 -2430 213 -2429
rect 240 -2430 241 -2429
rect 289 -2430 290 -2429
rect 324 -2430 325 -2429
rect 331 -2430 332 -2429
rect 373 -2430 374 -2429
rect 401 -2430 402 -2429
rect 513 -2430 514 -2429
rect 579 -2430 580 -2429
rect 730 -2430 731 -2429
rect 814 -2430 815 -2429
rect 1094 -2430 1095 -2429
rect 177 -2432 178 -2431
rect 240 -2432 241 -2431
rect 289 -2432 290 -2431
rect 352 -2432 353 -2431
rect 373 -2432 374 -2431
rect 828 -2432 829 -2431
rect 856 -2432 857 -2431
rect 1038 -2432 1039 -2431
rect 156 -2434 157 -2433
rect 177 -2434 178 -2433
rect 317 -2434 318 -2433
rect 345 -2434 346 -2433
rect 429 -2434 430 -2433
rect 534 -2434 535 -2433
rect 604 -2434 605 -2433
rect 1087 -2434 1088 -2433
rect 156 -2436 157 -2435
rect 233 -2436 234 -2435
rect 345 -2436 346 -2435
rect 467 -2436 468 -2435
rect 478 -2436 479 -2435
rect 562 -2436 563 -2435
rect 618 -2436 619 -2435
rect 681 -2436 682 -2435
rect 688 -2436 689 -2435
rect 926 -2436 927 -2435
rect 982 -2436 983 -2435
rect 1087 -2436 1088 -2435
rect 233 -2438 234 -2437
rect 527 -2438 528 -2437
rect 534 -2438 535 -2437
rect 632 -2438 633 -2437
rect 639 -2438 640 -2437
rect 737 -2438 738 -2437
rect 926 -2438 927 -2437
rect 1003 -2438 1004 -2437
rect 457 -2440 458 -2439
rect 492 -2440 493 -2439
rect 499 -2440 500 -2439
rect 506 -2440 507 -2439
rect 527 -2440 528 -2439
rect 695 -2440 696 -2439
rect 737 -2440 738 -2439
rect 943 -2440 944 -2439
rect 982 -2440 983 -2439
rect 1101 -2440 1102 -2439
rect 478 -2442 479 -2441
rect 583 -2442 584 -2441
rect 618 -2442 619 -2441
rect 716 -2442 717 -2441
rect 821 -2442 822 -2441
rect 1003 -2442 1004 -2441
rect 1094 -2442 1095 -2441
rect 1101 -2442 1102 -2441
rect 268 -2444 269 -2443
rect 583 -2444 584 -2443
rect 632 -2444 633 -2443
rect 800 -2444 801 -2443
rect 821 -2444 822 -2443
rect 1052 -2444 1053 -2443
rect 205 -2446 206 -2445
rect 268 -2446 269 -2445
rect 492 -2446 493 -2445
rect 793 -2446 794 -2445
rect 205 -2448 206 -2447
rect 219 -2448 220 -2447
rect 499 -2448 500 -2447
rect 572 -2448 573 -2447
rect 695 -2448 696 -2447
rect 1150 -2448 1151 -2447
rect 191 -2450 192 -2449
rect 219 -2450 220 -2449
rect 541 -2450 542 -2449
rect 800 -2450 801 -2449
rect 16 -2452 17 -2451
rect 191 -2452 192 -2451
rect 443 -2452 444 -2451
rect 541 -2452 542 -2451
rect 716 -2452 717 -2451
rect 835 -2452 836 -2451
rect 835 -2454 836 -2453
rect 1024 -2454 1025 -2453
rect 947 -2456 948 -2455
rect 1024 -2456 1025 -2455
rect 947 -2458 948 -2457
rect 1185 -2458 1186 -2457
rect 58 -2469 59 -2468
rect 460 -2469 461 -2468
rect 471 -2469 472 -2468
rect 523 -2469 524 -2468
rect 530 -2469 531 -2468
rect 583 -2469 584 -2468
rect 625 -2469 626 -2468
rect 866 -2469 867 -2468
rect 961 -2469 962 -2468
rect 1101 -2469 1102 -2468
rect 1108 -2469 1109 -2468
rect 1143 -2469 1144 -2468
rect 1185 -2469 1186 -2468
rect 1192 -2469 1193 -2468
rect 65 -2471 66 -2470
rect 352 -2471 353 -2470
rect 366 -2471 367 -2470
rect 586 -2471 587 -2470
rect 625 -2471 626 -2470
rect 821 -2471 822 -2470
rect 828 -2471 829 -2470
rect 870 -2471 871 -2470
rect 1013 -2471 1014 -2470
rect 1129 -2471 1130 -2470
rect 72 -2473 73 -2472
rect 131 -2473 132 -2472
rect 149 -2473 150 -2472
rect 352 -2473 353 -2472
rect 366 -2473 367 -2472
rect 604 -2473 605 -2472
rect 639 -2473 640 -2472
rect 642 -2473 643 -2472
rect 674 -2473 675 -2472
rect 758 -2473 759 -2472
rect 793 -2473 794 -2472
rect 807 -2473 808 -2472
rect 828 -2473 829 -2472
rect 856 -2473 857 -2472
rect 863 -2473 864 -2472
rect 870 -2473 871 -2472
rect 1024 -2473 1025 -2472
rect 1104 -2473 1105 -2472
rect 79 -2475 80 -2474
rect 471 -2475 472 -2474
rect 478 -2475 479 -2474
rect 695 -2475 696 -2474
rect 723 -2475 724 -2474
rect 947 -2475 948 -2474
rect 1038 -2475 1039 -2474
rect 1073 -2475 1074 -2474
rect 1087 -2475 1088 -2474
rect 1178 -2475 1179 -2474
rect 86 -2477 87 -2476
rect 166 -2477 167 -2476
rect 191 -2477 192 -2476
rect 691 -2477 692 -2476
rect 740 -2477 741 -2476
rect 877 -2477 878 -2476
rect 926 -2477 927 -2476
rect 947 -2477 948 -2476
rect 1052 -2477 1053 -2476
rect 1059 -2477 1060 -2476
rect 107 -2479 108 -2478
rect 467 -2479 468 -2478
rect 492 -2479 493 -2478
rect 604 -2479 605 -2478
rect 618 -2479 619 -2478
rect 723 -2479 724 -2478
rect 758 -2479 759 -2478
rect 842 -2479 843 -2478
rect 863 -2479 864 -2478
rect 982 -2479 983 -2478
rect 124 -2481 125 -2480
rect 226 -2481 227 -2480
rect 247 -2481 248 -2480
rect 492 -2481 493 -2480
rect 499 -2481 500 -2480
rect 583 -2481 584 -2480
rect 639 -2481 640 -2480
rect 786 -2481 787 -2480
rect 800 -2481 801 -2480
rect 810 -2481 811 -2480
rect 926 -2481 927 -2480
rect 996 -2481 997 -2480
rect 173 -2483 174 -2482
rect 247 -2483 248 -2482
rect 278 -2483 279 -2482
rect 359 -2483 360 -2482
rect 373 -2483 374 -2482
rect 443 -2483 444 -2482
rect 446 -2483 447 -2482
rect 849 -2483 850 -2482
rect 201 -2485 202 -2484
rect 226 -2485 227 -2484
rect 282 -2485 283 -2484
rect 478 -2485 479 -2484
rect 499 -2485 500 -2484
rect 744 -2485 745 -2484
rect 772 -2485 773 -2484
rect 793 -2485 794 -2484
rect 800 -2485 801 -2484
rect 912 -2485 913 -2484
rect 212 -2487 213 -2486
rect 551 -2487 552 -2486
rect 565 -2487 566 -2486
rect 975 -2487 976 -2486
rect 219 -2489 220 -2488
rect 355 -2489 356 -2488
rect 359 -2489 360 -2488
rect 376 -2489 377 -2488
rect 380 -2489 381 -2488
rect 684 -2489 685 -2488
rect 730 -2489 731 -2488
rect 786 -2489 787 -2488
rect 807 -2489 808 -2488
rect 989 -2489 990 -2488
rect 205 -2491 206 -2490
rect 380 -2491 381 -2490
rect 390 -2491 391 -2490
rect 513 -2491 514 -2490
rect 520 -2491 521 -2490
rect 695 -2491 696 -2490
rect 730 -2491 731 -2490
rect 751 -2491 752 -2490
rect 772 -2491 773 -2490
rect 835 -2491 836 -2490
rect 912 -2491 913 -2490
rect 954 -2491 955 -2490
rect 975 -2491 976 -2490
rect 1003 -2491 1004 -2490
rect 93 -2493 94 -2492
rect 520 -2493 521 -2492
rect 544 -2493 545 -2492
rect 572 -2493 573 -2492
rect 597 -2493 598 -2492
rect 744 -2493 745 -2492
rect 954 -2493 955 -2492
rect 1017 -2493 1018 -2492
rect 114 -2495 115 -2494
rect 572 -2495 573 -2494
rect 597 -2495 598 -2494
rect 737 -2495 738 -2494
rect 1017 -2495 1018 -2494
rect 1031 -2495 1032 -2494
rect 282 -2497 283 -2496
rect 345 -2497 346 -2496
rect 373 -2497 374 -2496
rect 534 -2497 535 -2496
rect 548 -2497 549 -2496
rect 943 -2497 944 -2496
rect 1031 -2497 1032 -2496
rect 1066 -2497 1067 -2496
rect 289 -2499 290 -2498
rect 611 -2499 612 -2498
rect 646 -2499 647 -2498
rect 751 -2499 752 -2498
rect 1066 -2499 1067 -2498
rect 1080 -2499 1081 -2498
rect 233 -2501 234 -2500
rect 289 -2501 290 -2500
rect 296 -2501 297 -2500
rect 677 -2501 678 -2500
rect 170 -2503 171 -2502
rect 233 -2503 234 -2502
rect 296 -2503 297 -2502
rect 303 -2503 304 -2502
rect 317 -2503 318 -2502
rect 439 -2503 440 -2502
rect 443 -2503 444 -2502
rect 555 -2503 556 -2502
rect 569 -2503 570 -2502
rect 779 -2503 780 -2502
rect 100 -2505 101 -2504
rect 303 -2505 304 -2504
rect 327 -2505 328 -2504
rect 401 -2505 402 -2504
rect 415 -2505 416 -2504
rect 534 -2505 535 -2504
rect 541 -2505 542 -2504
rect 611 -2505 612 -2504
rect 642 -2505 643 -2504
rect 646 -2505 647 -2504
rect 653 -2505 654 -2504
rect 737 -2505 738 -2504
rect 240 -2507 241 -2506
rect 415 -2507 416 -2506
rect 422 -2507 423 -2506
rect 618 -2507 619 -2506
rect 653 -2507 654 -2506
rect 702 -2507 703 -2506
rect 275 -2509 276 -2508
rect 317 -2509 318 -2508
rect 331 -2509 332 -2508
rect 464 -2509 465 -2508
rect 509 -2509 510 -2508
rect 968 -2509 969 -2508
rect 128 -2511 129 -2510
rect 331 -2511 332 -2510
rect 345 -2511 346 -2510
rect 485 -2511 486 -2510
rect 513 -2511 514 -2510
rect 709 -2511 710 -2510
rect 121 -2513 122 -2512
rect 128 -2513 129 -2512
rect 310 -2513 311 -2512
rect 401 -2513 402 -2512
rect 429 -2513 430 -2512
rect 660 -2513 661 -2512
rect 667 -2513 668 -2512
rect 674 -2513 675 -2512
rect 702 -2513 703 -2512
rect 716 -2513 717 -2512
rect 184 -2515 185 -2514
rect 310 -2515 311 -2514
rect 408 -2515 409 -2514
rect 429 -2515 430 -2514
rect 436 -2515 437 -2514
rect 905 -2515 906 -2514
rect 268 -2517 269 -2516
rect 408 -2517 409 -2516
rect 450 -2517 451 -2516
rect 474 -2517 475 -2516
rect 485 -2517 486 -2516
rect 814 -2517 815 -2516
rect 142 -2519 143 -2518
rect 268 -2519 269 -2518
rect 387 -2519 388 -2518
rect 436 -2519 437 -2518
rect 527 -2519 528 -2518
rect 709 -2519 710 -2518
rect 177 -2521 178 -2520
rect 450 -2521 451 -2520
rect 548 -2521 549 -2520
rect 919 -2521 920 -2520
rect 387 -2523 388 -2522
rect 394 -2523 395 -2522
rect 555 -2523 556 -2522
rect 688 -2523 689 -2522
rect 324 -2525 325 -2524
rect 394 -2525 395 -2524
rect 569 -2525 570 -2524
rect 681 -2525 682 -2524
rect 576 -2527 577 -2526
rect 667 -2527 668 -2526
rect 681 -2527 682 -2526
rect 933 -2527 934 -2526
rect 457 -2529 458 -2528
rect 576 -2529 577 -2528
rect 590 -2529 591 -2528
rect 779 -2529 780 -2528
rect 884 -2529 885 -2528
rect 933 -2529 934 -2528
rect 422 -2531 423 -2530
rect 457 -2531 458 -2530
rect 590 -2531 591 -2530
rect 891 -2531 892 -2530
rect 632 -2533 633 -2532
rect 716 -2533 717 -2532
rect 562 -2535 563 -2534
rect 632 -2535 633 -2534
rect 660 -2535 661 -2534
rect 765 -2535 766 -2534
rect 506 -2537 507 -2536
rect 562 -2537 563 -2536
rect 765 -2537 766 -2536
rect 898 -2537 899 -2536
rect 261 -2539 262 -2538
rect 506 -2539 507 -2538
rect 156 -2541 157 -2540
rect 261 -2541 262 -2540
rect 131 -2552 132 -2551
rect 135 -2552 136 -2551
rect 226 -2552 227 -2551
rect 257 -2552 258 -2551
rect 261 -2552 262 -2551
rect 366 -2552 367 -2551
rect 380 -2552 381 -2551
rect 527 -2552 528 -2551
rect 530 -2552 531 -2551
rect 702 -2552 703 -2551
rect 716 -2552 717 -2551
rect 807 -2552 808 -2551
rect 814 -2552 815 -2551
rect 828 -2552 829 -2551
rect 866 -2552 867 -2551
rect 926 -2552 927 -2551
rect 933 -2552 934 -2551
rect 964 -2552 965 -2551
rect 968 -2552 969 -2551
rect 975 -2552 976 -2551
rect 1013 -2552 1014 -2551
rect 1038 -2552 1039 -2551
rect 1045 -2552 1046 -2551
rect 1052 -2552 1053 -2551
rect 1059 -2552 1060 -2551
rect 1066 -2552 1067 -2551
rect 1143 -2552 1144 -2551
rect 1178 -2552 1179 -2551
rect 1181 -2552 1182 -2551
rect 1185 -2552 1186 -2551
rect 128 -2554 129 -2553
rect 135 -2554 136 -2553
rect 233 -2554 234 -2553
rect 275 -2554 276 -2553
rect 282 -2554 283 -2553
rect 387 -2554 388 -2553
rect 394 -2554 395 -2553
rect 471 -2554 472 -2553
rect 478 -2554 479 -2553
rect 677 -2554 678 -2553
rect 681 -2554 682 -2553
rect 772 -2554 773 -2553
rect 870 -2554 871 -2553
rect 887 -2554 888 -2553
rect 898 -2554 899 -2553
rect 912 -2554 913 -2553
rect 1024 -2554 1025 -2553
rect 1031 -2554 1032 -2553
rect 247 -2556 248 -2555
rect 324 -2556 325 -2555
rect 331 -2556 332 -2555
rect 485 -2556 486 -2555
rect 492 -2556 493 -2555
rect 684 -2556 685 -2555
rect 688 -2556 689 -2555
rect 730 -2556 731 -2555
rect 744 -2556 745 -2555
rect 793 -2556 794 -2555
rect 884 -2556 885 -2555
rect 954 -2556 955 -2555
rect 268 -2558 269 -2557
rect 324 -2558 325 -2557
rect 345 -2558 346 -2557
rect 366 -2558 367 -2557
rect 401 -2558 402 -2557
rect 548 -2558 549 -2557
rect 551 -2558 552 -2557
rect 653 -2558 654 -2557
rect 663 -2558 664 -2557
rect 667 -2558 668 -2557
rect 681 -2558 682 -2557
rect 779 -2558 780 -2557
rect 947 -2558 948 -2557
rect 954 -2558 955 -2557
rect 289 -2560 290 -2559
rect 383 -2560 384 -2559
rect 415 -2560 416 -2559
rect 492 -2560 493 -2559
rect 506 -2560 507 -2559
rect 611 -2560 612 -2559
rect 621 -2560 622 -2559
rect 800 -2560 801 -2559
rect 303 -2562 304 -2561
rect 593 -2562 594 -2561
rect 600 -2562 601 -2561
rect 646 -2562 647 -2561
rect 660 -2562 661 -2561
rect 667 -2562 668 -2561
rect 716 -2562 717 -2561
rect 758 -2562 759 -2561
rect 310 -2564 311 -2563
rect 649 -2564 650 -2563
rect 723 -2564 724 -2563
rect 810 -2564 811 -2563
rect 317 -2566 318 -2565
rect 331 -2566 332 -2565
rect 359 -2566 360 -2565
rect 506 -2566 507 -2565
rect 523 -2566 524 -2565
rect 541 -2566 542 -2565
rect 565 -2566 566 -2565
rect 639 -2566 640 -2565
rect 723 -2566 724 -2565
rect 765 -2566 766 -2565
rect 429 -2568 430 -2567
rect 488 -2568 489 -2567
rect 527 -2568 528 -2567
rect 555 -2568 556 -2567
rect 569 -2568 570 -2567
rect 674 -2568 675 -2567
rect 730 -2568 731 -2567
rect 751 -2568 752 -2567
rect 436 -2570 437 -2569
rect 544 -2570 545 -2569
rect 576 -2570 577 -2569
rect 590 -2570 591 -2569
rect 632 -2570 633 -2569
rect 712 -2570 713 -2569
rect 747 -2570 748 -2569
rect 786 -2570 787 -2569
rect 443 -2572 444 -2571
rect 460 -2572 461 -2571
rect 513 -2572 514 -2571
rect 555 -2572 556 -2571
rect 576 -2572 577 -2571
rect 597 -2572 598 -2571
rect 695 -2572 696 -2571
rect 751 -2572 752 -2571
rect 338 -2574 339 -2573
rect 513 -2574 514 -2573
rect 530 -2574 531 -2573
rect 562 -2574 563 -2573
rect 296 -2576 297 -2575
rect 338 -2576 339 -2575
rect 373 -2576 374 -2575
rect 443 -2576 444 -2575
rect 450 -2576 451 -2575
rect 569 -2576 570 -2575
rect 352 -2578 353 -2577
rect 450 -2578 451 -2577
rect 464 -2578 465 -2577
rect 597 -2578 598 -2577
rect 373 -2580 374 -2579
rect 422 -2580 423 -2579
rect 534 -2580 535 -2579
rect 646 -2580 647 -2579
rect 408 -2582 409 -2581
rect 534 -2582 535 -2581
rect 541 -2582 542 -2581
rect 709 -2582 710 -2581
rect 562 -2584 563 -2583
rect 625 -2584 626 -2583
rect 604 -2586 605 -2585
rect 709 -2586 710 -2585
rect 131 -2597 132 -2596
rect 135 -2597 136 -2596
rect 324 -2597 325 -2596
rect 383 -2597 384 -2596
rect 443 -2597 444 -2596
rect 516 -2597 517 -2596
rect 534 -2597 535 -2596
rect 663 -2597 664 -2596
rect 674 -2597 675 -2596
rect 723 -2597 724 -2596
rect 751 -2597 752 -2596
rect 807 -2597 808 -2596
rect 810 -2597 811 -2596
rect 814 -2597 815 -2596
rect 884 -2597 885 -2596
rect 898 -2597 899 -2596
rect 954 -2597 955 -2596
rect 964 -2597 965 -2596
rect 1010 -2597 1011 -2596
rect 1017 -2597 1018 -2596
rect 1045 -2597 1046 -2596
rect 1052 -2597 1053 -2596
rect 1055 -2597 1056 -2596
rect 1059 -2597 1060 -2596
rect 331 -2599 332 -2598
rect 348 -2599 349 -2598
rect 366 -2599 367 -2598
rect 380 -2599 381 -2598
rect 450 -2599 451 -2598
rect 544 -2599 545 -2598
rect 548 -2599 549 -2598
rect 576 -2599 577 -2598
rect 660 -2599 661 -2598
rect 667 -2599 668 -2598
rect 684 -2599 685 -2598
rect 716 -2599 717 -2598
rect 961 -2599 962 -2598
rect 968 -2599 969 -2598
rect 1013 -2599 1014 -2598
rect 1024 -2599 1025 -2598
rect 338 -2601 339 -2600
rect 373 -2601 374 -2600
rect 471 -2601 472 -2600
rect 551 -2601 552 -2600
rect 555 -2601 556 -2600
rect 600 -2601 601 -2600
rect 709 -2601 710 -2600
rect 730 -2601 731 -2600
rect 492 -2603 493 -2602
rect 565 -2603 566 -2602
rect 569 -2603 570 -2602
rect 681 -2603 682 -2602
rect 499 -2605 500 -2604
rect 513 -2605 514 -2604
rect 506 -2607 507 -2606
rect 649 -2607 650 -2606
<< metal2 >>
rect 215 -15 216 1
rect 240 -15 241 1
rect 247 -15 248 1
rect 478 -15 479 1
rect 562 -15 563 1
rect 639 -15 640 1
rect 667 -15 668 1
rect 702 -15 703 1
rect 800 -15 801 1
rect 828 -15 829 1
rect 261 -15 262 -1
rect 268 -15 269 -1
rect 275 -15 276 -1
rect 408 -15 409 -1
rect 411 -15 412 -1
rect 506 -15 507 -1
rect 576 -15 577 -1
rect 607 -15 608 -1
rect 681 -15 682 -1
rect 803 -15 804 -1
rect 338 -15 339 -3
rect 380 -15 381 -3
rect 387 -15 388 -3
rect 583 -15 584 -3
rect 586 -15 587 -3
rect 709 -15 710 -3
rect 373 -15 374 -5
rect 401 -15 402 -5
rect 415 -15 416 -5
rect 457 -15 458 -5
rect 464 -15 465 -5
rect 527 -15 528 -5
rect 604 -15 605 -5
rect 765 -15 766 -5
rect 397 -15 398 -7
rect 485 -15 486 -7
rect 425 -15 426 -9
rect 569 -15 570 -9
rect 429 -15 430 -11
rect 516 -15 517 -11
rect 467 -15 468 -13
rect 499 -15 500 -13
rect 156 -25 157 -23
rect 156 -58 157 -24
rect 156 -25 157 -23
rect 156 -58 157 -24
rect 163 -58 164 -24
rect 285 -25 286 -23
rect 292 -58 293 -24
rect 338 -25 339 -23
rect 359 -58 360 -24
rect 467 -25 468 -23
rect 478 -25 479 -23
rect 604 -58 605 -24
rect 621 -58 622 -24
rect 723 -58 724 -24
rect 800 -25 801 -23
rect 905 -58 906 -24
rect 191 -58 192 -26
rect 247 -27 248 -23
rect 254 -58 255 -26
rect 401 -27 402 -23
rect 404 -27 405 -23
rect 443 -58 444 -26
rect 464 -58 465 -26
rect 607 -27 608 -23
rect 639 -27 640 -23
rect 688 -58 689 -26
rect 702 -27 703 -23
rect 751 -58 752 -26
rect 828 -27 829 -23
rect 849 -58 850 -26
rect 215 -29 216 -23
rect 219 -58 220 -28
rect 226 -58 227 -28
rect 275 -29 276 -23
rect 282 -29 283 -23
rect 394 -58 395 -28
rect 401 -58 402 -28
rect 411 -58 412 -28
rect 436 -58 437 -28
rect 460 -29 461 -23
rect 481 -29 482 -23
rect 660 -58 661 -28
rect 667 -29 668 -23
rect 674 -58 675 -28
rect 709 -29 710 -23
rect 758 -58 759 -28
rect 765 -29 766 -23
rect 828 -58 829 -28
rect 233 -58 234 -30
rect 240 -31 241 -23
rect 247 -58 248 -30
rect 261 -31 262 -23
rect 268 -58 269 -30
rect 383 -31 384 -23
rect 408 -31 409 -23
rect 471 -58 472 -30
rect 485 -31 486 -23
rect 520 -58 521 -30
rect 527 -31 528 -23
rect 541 -58 542 -30
rect 551 -31 552 -23
rect 597 -58 598 -30
rect 639 -58 640 -30
rect 681 -31 682 -23
rect 719 -58 720 -30
rect 877 -58 878 -30
rect 261 -58 262 -32
rect 387 -33 388 -23
rect 492 -58 493 -32
rect 548 -33 549 -23
rect 555 -58 556 -32
rect 681 -58 682 -32
rect 275 -58 276 -34
rect 355 -58 356 -34
rect 366 -58 367 -34
rect 513 -35 514 -23
rect 516 -35 517 -23
rect 632 -58 633 -34
rect 653 -58 654 -34
rect 716 -58 717 -34
rect 282 -58 283 -36
rect 425 -37 426 -23
rect 499 -37 500 -23
rect 513 -58 514 -36
rect 534 -58 535 -36
rect 702 -58 703 -36
rect 296 -58 297 -38
rect 429 -39 430 -23
rect 502 -58 503 -38
rect 527 -58 528 -38
rect 548 -58 549 -38
rect 618 -58 619 -38
rect 303 -58 304 -40
rect 397 -41 398 -23
rect 429 -58 430 -40
rect 537 -58 538 -40
rect 569 -41 570 -23
rect 625 -58 626 -40
rect 310 -58 311 -42
rect 422 -58 423 -42
rect 457 -43 458 -23
rect 569 -58 570 -42
rect 576 -43 577 -23
rect 611 -58 612 -42
rect 317 -58 318 -44
rect 579 -58 580 -44
rect 583 -45 584 -23
rect 646 -58 647 -44
rect 324 -58 325 -46
rect 373 -47 374 -23
rect 380 -47 381 -23
rect 485 -58 486 -46
rect 506 -47 507 -23
rect 583 -58 584 -46
rect 593 -58 594 -46
rect 772 -58 773 -46
rect 331 -58 332 -48
rect 418 -58 419 -48
rect 457 -58 458 -48
rect 478 -58 479 -48
rect 506 -58 507 -48
rect 562 -49 563 -23
rect 345 -58 346 -50
rect 667 -58 668 -50
rect 373 -58 374 -52
rect 415 -53 416 -23
rect 380 -58 381 -54
rect 562 -58 563 -54
rect 387 -58 388 -56
rect 499 -58 500 -56
rect 23 -119 24 -67
rect 355 -68 356 -66
rect 415 -68 416 -66
rect 548 -68 549 -66
rect 562 -68 563 -66
rect 709 -119 710 -67
rect 723 -68 724 -66
rect 779 -119 780 -67
rect 828 -68 829 -66
rect 870 -119 871 -67
rect 877 -68 878 -66
rect 940 -119 941 -67
rect 1500 -119 1501 -67
rect 1507 -119 1508 -67
rect 30 -119 31 -69
rect 152 -70 153 -66
rect 156 -119 157 -69
rect 292 -70 293 -66
rect 303 -70 304 -66
rect 303 -119 304 -69
rect 303 -70 304 -66
rect 303 -119 304 -69
rect 313 -119 314 -69
rect 397 -119 398 -69
rect 422 -70 423 -66
rect 548 -119 549 -69
rect 562 -119 563 -69
rect 639 -70 640 -66
rect 663 -119 664 -69
rect 856 -119 857 -69
rect 905 -70 906 -66
rect 947 -119 948 -69
rect 37 -119 38 -71
rect 331 -72 332 -66
rect 373 -72 374 -66
rect 415 -119 416 -71
rect 478 -72 479 -66
rect 695 -119 696 -71
rect 702 -72 703 -66
rect 800 -119 801 -71
rect 849 -72 850 -66
rect 877 -119 878 -71
rect 44 -119 45 -73
rect 159 -74 160 -66
rect 170 -119 171 -73
rect 310 -74 311 -66
rect 324 -74 325 -66
rect 380 -119 381 -73
rect 394 -74 395 -66
rect 478 -119 479 -73
rect 481 -74 482 -66
rect 485 -74 486 -66
rect 499 -74 500 -66
rect 534 -119 535 -73
rect 541 -74 542 -66
rect 579 -74 580 -66
rect 604 -74 605 -66
rect 723 -119 724 -73
rect 751 -74 752 -66
rect 814 -119 815 -73
rect 51 -119 52 -75
rect 366 -76 367 -66
rect 373 -119 374 -75
rect 429 -76 430 -66
rect 471 -76 472 -66
rect 541 -119 542 -75
rect 576 -76 577 -66
rect 821 -119 822 -75
rect 75 -119 76 -77
rect 100 -119 101 -77
rect 107 -119 108 -77
rect 117 -119 118 -77
rect 121 -119 122 -77
rect 450 -78 451 -66
rect 471 -119 472 -77
rect 555 -78 556 -66
rect 576 -119 577 -77
rect 593 -78 594 -66
rect 604 -119 605 -77
rect 751 -119 752 -77
rect 758 -78 759 -66
rect 786 -119 787 -77
rect 79 -119 80 -79
rect 383 -80 384 -66
rect 429 -119 430 -79
rect 457 -80 458 -66
rect 485 -119 486 -79
rect 611 -80 612 -66
rect 618 -80 619 -66
rect 716 -119 717 -79
rect 772 -80 773 -66
rect 849 -119 850 -79
rect 86 -119 87 -81
rect 89 -119 90 -81
rect 93 -119 94 -81
rect 275 -82 276 -66
rect 296 -82 297 -66
rect 422 -119 423 -81
rect 436 -82 437 -66
rect 457 -119 458 -81
rect 499 -119 500 -81
rect 558 -82 559 -66
rect 618 -119 619 -81
rect 674 -82 675 -66
rect 681 -82 682 -66
rect 730 -119 731 -81
rect 114 -119 115 -83
rect 275 -119 276 -83
rect 299 -119 300 -83
rect 436 -119 437 -83
rect 450 -119 451 -83
rect 597 -84 598 -66
rect 632 -84 633 -66
rect 681 -119 682 -83
rect 688 -84 689 -66
rect 744 -119 745 -83
rect 128 -119 129 -85
rect 212 -119 213 -85
rect 219 -86 220 -66
rect 331 -119 332 -85
rect 352 -86 353 -66
rect 555 -119 556 -85
rect 625 -86 626 -66
rect 632 -119 633 -85
rect 646 -86 647 -66
rect 772 -119 773 -85
rect 135 -119 136 -87
rect 317 -88 318 -66
rect 352 -119 353 -87
rect 359 -88 360 -66
rect 366 -119 367 -87
rect 387 -88 388 -66
rect 404 -119 405 -87
rect 646 -119 647 -87
rect 660 -88 661 -66
rect 674 -119 675 -87
rect 142 -119 143 -89
rect 163 -90 164 -66
rect 177 -119 178 -89
rect 341 -90 342 -66
rect 359 -119 360 -89
rect 702 -119 703 -89
rect 163 -119 164 -91
rect 327 -119 328 -91
rect 338 -92 339 -66
rect 387 -119 388 -91
rect 453 -92 454 -66
rect 688 -119 689 -91
rect 184 -119 185 -93
rect 282 -94 283 -66
rect 338 -119 339 -93
rect 394 -119 395 -93
rect 506 -94 507 -66
rect 611 -119 612 -93
rect 625 -119 626 -93
rect 653 -94 654 -66
rect 660 -119 661 -93
rect 737 -119 738 -93
rect 187 -119 188 -95
rect 226 -96 227 -66
rect 254 -96 255 -66
rect 317 -119 318 -95
rect 464 -96 465 -66
rect 506 -119 507 -95
rect 513 -96 514 -66
rect 597 -119 598 -95
rect 667 -119 668 -95
rect 719 -96 720 -66
rect 149 -98 150 -66
rect 226 -119 227 -97
rect 254 -119 255 -97
rect 261 -98 262 -66
rect 268 -98 269 -66
rect 408 -119 409 -97
rect 411 -98 412 -66
rect 513 -119 514 -97
rect 520 -98 521 -66
rect 639 -119 640 -97
rect 670 -98 671 -66
rect 807 -119 808 -97
rect 149 -119 150 -99
rect 194 -119 195 -99
rect 198 -119 199 -99
rect 233 -100 234 -66
rect 247 -100 248 -66
rect 268 -119 269 -99
rect 271 -119 272 -99
rect 310 -119 311 -99
rect 520 -119 521 -99
rect 607 -119 608 -99
rect 191 -102 192 -66
rect 240 -119 241 -101
rect 247 -119 248 -101
rect 418 -102 419 -66
rect 527 -102 528 -66
rect 765 -119 766 -101
rect 205 -119 206 -103
rect 348 -104 349 -66
rect 530 -119 531 -103
rect 793 -119 794 -103
rect 219 -119 220 -105
rect 345 -106 346 -66
rect 569 -106 570 -66
rect 653 -119 654 -105
rect 233 -119 234 -107
rect 289 -108 290 -66
rect 345 -119 346 -107
rect 590 -108 591 -66
rect 65 -119 66 -109
rect 289 -119 290 -109
rect 443 -110 444 -66
rect 569 -119 570 -109
rect 261 -119 262 -111
rect 401 -112 402 -66
rect 439 -119 440 -111
rect 443 -119 444 -111
rect 492 -112 493 -66
rect 590 -119 591 -111
rect 282 -119 283 -113
rect 537 -114 538 -66
rect 401 -119 402 -115
rect 464 -119 465 -115
rect 492 -119 493 -115
rect 583 -116 584 -66
rect 583 -119 584 -117
rect 761 -119 762 -117
rect 16 -198 17 -128
rect 439 -129 440 -127
rect 488 -198 489 -128
rect 765 -129 766 -127
rect 793 -129 794 -127
rect 828 -198 829 -128
rect 849 -129 850 -127
rect 884 -198 885 -128
rect 940 -129 941 -127
rect 968 -198 969 -128
rect 975 -198 976 -128
rect 1024 -198 1025 -128
rect 1500 -129 1501 -127
rect 1500 -198 1501 -128
rect 1500 -129 1501 -127
rect 1500 -198 1501 -128
rect 9 -198 10 -130
rect 439 -198 440 -130
rect 516 -198 517 -130
rect 597 -131 598 -127
rect 604 -198 605 -130
rect 772 -131 773 -127
rect 800 -131 801 -127
rect 912 -198 913 -130
rect 947 -131 948 -127
rect 978 -198 979 -130
rect 23 -133 24 -127
rect 23 -198 24 -132
rect 23 -133 24 -127
rect 23 -198 24 -132
rect 30 -133 31 -127
rect 54 -198 55 -132
rect 58 -133 59 -127
rect 65 -198 66 -132
rect 72 -198 73 -132
rect 75 -133 76 -127
rect 86 -198 87 -132
rect 366 -133 367 -127
rect 394 -198 395 -132
rect 985 -198 986 -132
rect 30 -198 31 -134
rect 61 -135 62 -127
rect 107 -135 108 -127
rect 114 -198 115 -134
rect 117 -135 118 -127
rect 390 -198 391 -134
rect 537 -198 538 -134
rect 835 -198 836 -134
rect 849 -198 850 -134
rect 982 -198 983 -134
rect 44 -137 45 -127
rect 271 -137 272 -127
rect 275 -137 276 -127
rect 359 -198 360 -136
rect 541 -137 542 -127
rect 597 -198 598 -136
rect 607 -137 608 -127
rect 919 -198 920 -136
rect 51 -139 52 -127
rect 401 -139 402 -127
rect 464 -139 465 -127
rect 607 -198 608 -138
rect 611 -139 612 -127
rect 842 -198 843 -138
rect 856 -139 857 -127
rect 961 -198 962 -138
rect 51 -198 52 -140
rect 142 -141 143 -127
rect 145 -198 146 -140
rect 299 -141 300 -127
rect 310 -141 311 -127
rect 401 -198 402 -140
rect 443 -141 444 -127
rect 464 -198 465 -140
rect 478 -141 479 -127
rect 611 -198 612 -140
rect 632 -141 633 -127
rect 632 -198 633 -140
rect 632 -141 633 -127
rect 632 -198 633 -140
rect 646 -141 647 -127
rect 793 -198 794 -140
rect 807 -141 808 -127
rect 891 -198 892 -140
rect 58 -198 59 -142
rect 79 -143 80 -127
rect 93 -143 94 -127
rect 275 -198 276 -142
rect 289 -143 290 -127
rect 527 -143 528 -127
rect 555 -143 556 -127
rect 996 -198 997 -142
rect 79 -198 80 -144
rect 163 -145 164 -127
rect 226 -145 227 -127
rect 296 -145 297 -127
rect 327 -145 328 -127
rect 352 -145 353 -127
rect 422 -145 423 -127
rect 478 -198 479 -144
rect 513 -145 514 -127
rect 541 -198 542 -144
rect 562 -145 563 -127
rect 772 -198 773 -144
rect 779 -145 780 -127
rect 856 -198 857 -144
rect 870 -145 871 -127
rect 926 -198 927 -144
rect 121 -147 122 -127
rect 184 -198 185 -146
rect 226 -198 227 -146
rect 362 -147 363 -127
rect 422 -198 423 -146
rect 499 -147 500 -127
rect 520 -147 521 -127
rect 527 -198 528 -146
rect 646 -198 647 -146
rect 681 -147 682 -127
rect 688 -147 689 -127
rect 758 -198 759 -146
rect 779 -198 780 -146
rect 814 -147 815 -127
rect 821 -147 822 -127
rect 954 -198 955 -146
rect 89 -149 90 -127
rect 520 -198 521 -148
rect 639 -149 640 -127
rect 821 -198 822 -148
rect 877 -149 878 -127
rect 947 -198 948 -148
rect 100 -151 101 -127
rect 121 -198 122 -150
rect 131 -151 132 -127
rect 310 -198 311 -150
rect 324 -151 325 -127
rect 352 -198 353 -150
rect 429 -151 430 -127
rect 555 -198 556 -150
rect 583 -151 584 -127
rect 639 -198 640 -150
rect 653 -151 654 -127
rect 877 -198 878 -150
rect 68 -153 69 -127
rect 100 -198 101 -152
rect 135 -153 136 -127
rect 296 -198 297 -152
rect 443 -198 444 -152
rect 709 -153 710 -127
rect 716 -153 717 -127
rect 905 -198 906 -152
rect 135 -198 136 -154
rect 170 -155 171 -127
rect 233 -155 234 -127
rect 366 -198 367 -154
rect 485 -155 486 -127
rect 583 -198 584 -154
rect 590 -155 591 -127
rect 709 -198 710 -154
rect 719 -198 720 -154
rect 800 -198 801 -154
rect 807 -198 808 -154
rect 989 -198 990 -154
rect 142 -198 143 -156
rect 191 -157 192 -127
rect 194 -157 195 -127
rect 233 -198 234 -156
rect 247 -157 248 -127
rect 324 -198 325 -156
rect 415 -157 416 -127
rect 590 -198 591 -156
rect 625 -157 626 -127
rect 653 -198 654 -156
rect 660 -198 661 -156
rect 786 -157 787 -127
rect 149 -159 150 -127
rect 187 -159 188 -127
rect 247 -198 248 -158
rect 397 -159 398 -127
rect 415 -198 416 -158
rect 471 -159 472 -127
rect 485 -198 486 -158
rect 562 -198 563 -158
rect 576 -159 577 -127
rect 625 -198 626 -158
rect 667 -159 668 -127
rect 814 -198 815 -158
rect 44 -198 45 -160
rect 149 -198 150 -160
rect 152 -198 153 -160
rect 191 -198 192 -160
rect 254 -161 255 -127
rect 320 -198 321 -160
rect 387 -161 388 -127
rect 471 -198 472 -160
rect 492 -161 493 -127
rect 576 -198 577 -160
rect 663 -161 664 -127
rect 667 -198 668 -160
rect 674 -161 675 -127
rect 765 -198 766 -160
rect 163 -198 164 -162
rect 177 -163 178 -127
rect 219 -163 220 -127
rect 254 -198 255 -162
rect 271 -198 272 -162
rect 317 -163 318 -127
rect 373 -163 374 -127
rect 387 -198 388 -162
rect 457 -163 458 -127
rect 492 -198 493 -162
rect 569 -163 570 -127
rect 674 -198 675 -162
rect 688 -198 689 -162
rect 695 -163 696 -127
rect 702 -163 703 -127
rect 898 -198 899 -162
rect 170 -198 171 -164
rect 205 -165 206 -127
rect 219 -198 220 -164
rect 306 -198 307 -164
rect 317 -198 318 -164
rect 681 -198 682 -164
rect 723 -165 724 -127
rect 933 -198 934 -164
rect 177 -198 178 -166
rect 212 -167 213 -127
rect 268 -167 269 -127
rect 702 -198 703 -166
rect 730 -167 731 -127
rect 786 -198 787 -166
rect 107 -198 108 -168
rect 268 -198 269 -168
rect 282 -169 283 -127
rect 289 -198 290 -168
rect 303 -169 304 -127
rect 373 -198 374 -168
rect 457 -198 458 -168
rect 695 -198 696 -168
rect 737 -169 738 -127
rect 870 -198 871 -168
rect 198 -171 199 -127
rect 205 -198 206 -170
rect 240 -171 241 -127
rect 282 -198 283 -170
rect 303 -198 304 -170
rect 429 -198 430 -170
rect 530 -171 531 -127
rect 737 -198 738 -170
rect 744 -171 745 -127
rect 863 -198 864 -170
rect 128 -198 129 -172
rect 240 -198 241 -172
rect 331 -173 332 -127
rect 569 -198 570 -172
rect 618 -173 619 -127
rect 723 -198 724 -172
rect 751 -173 752 -127
rect 940 -198 941 -172
rect 93 -198 94 -174
rect 331 -198 332 -174
rect 334 -198 335 -174
rect 730 -198 731 -174
rect 156 -177 157 -127
rect 198 -198 199 -176
rect 436 -177 437 -127
rect 744 -198 745 -176
rect 156 -198 157 -178
rect 212 -198 213 -178
rect 436 -198 437 -178
rect 499 -198 500 -178
rect 534 -179 535 -127
rect 618 -198 619 -178
rect 450 -181 451 -127
rect 534 -198 535 -180
rect 548 -181 549 -127
rect 751 -198 752 -180
rect 408 -183 409 -127
rect 450 -198 451 -182
rect 506 -183 507 -127
rect 548 -198 549 -182
rect 103 -198 104 -184
rect 506 -198 507 -184
rect 380 -187 381 -127
rect 408 -198 409 -186
rect 338 -189 339 -127
rect 380 -198 381 -188
rect 338 -198 339 -190
rect 345 -191 346 -127
rect 37 -193 38 -127
rect 345 -198 346 -192
rect 37 -198 38 -194
rect 261 -195 262 -127
rect 261 -198 262 -196
rect 460 -198 461 -196
rect 2 -309 3 -207
rect 30 -208 31 -206
rect 37 -208 38 -206
rect 387 -208 388 -206
rect 436 -208 437 -206
rect 590 -208 591 -206
rect 604 -208 605 -206
rect 1080 -309 1081 -207
rect 1150 -309 1151 -207
rect 1178 -309 1179 -207
rect 1500 -208 1501 -206
rect 1500 -309 1501 -207
rect 1500 -208 1501 -206
rect 1500 -309 1501 -207
rect 16 -210 17 -206
rect 16 -309 17 -209
rect 16 -210 17 -206
rect 16 -309 17 -209
rect 37 -309 38 -209
rect 387 -309 388 -209
rect 394 -210 395 -206
rect 436 -309 437 -209
rect 439 -210 440 -206
rect 842 -210 843 -206
rect 849 -210 850 -206
rect 1059 -309 1060 -209
rect 44 -212 45 -206
rect 285 -309 286 -211
rect 303 -212 304 -206
rect 313 -309 314 -211
rect 446 -212 447 -206
rect 793 -212 794 -206
rect 835 -212 836 -206
rect 1087 -309 1088 -211
rect 44 -309 45 -213
rect 65 -214 66 -206
rect 72 -214 73 -206
rect 82 -309 83 -213
rect 103 -214 104 -206
rect 240 -214 241 -206
rect 243 -214 244 -206
rect 537 -214 538 -206
rect 544 -309 545 -213
rect 821 -214 822 -206
rect 863 -214 864 -206
rect 1108 -309 1109 -213
rect 51 -216 52 -206
rect 989 -309 990 -215
rect 1024 -216 1025 -206
rect 1045 -309 1046 -215
rect 51 -309 52 -217
rect 100 -309 101 -217
rect 107 -218 108 -206
rect 303 -309 304 -217
rect 310 -218 311 -206
rect 394 -309 395 -217
rect 453 -309 454 -217
rect 877 -218 878 -206
rect 891 -218 892 -206
rect 1017 -309 1018 -217
rect 65 -309 66 -219
rect 72 -309 73 -219
rect 107 -309 108 -219
rect 443 -220 444 -206
rect 464 -220 465 -206
rect 464 -309 465 -219
rect 464 -220 465 -206
rect 464 -309 465 -219
rect 471 -220 472 -206
rect 471 -309 472 -219
rect 471 -220 472 -206
rect 471 -309 472 -219
rect 485 -220 486 -206
rect 814 -220 815 -206
rect 821 -309 822 -219
rect 828 -220 829 -206
rect 870 -220 871 -206
rect 1101 -309 1102 -219
rect 96 -309 97 -221
rect 870 -309 871 -221
rect 912 -222 913 -206
rect 1122 -309 1123 -221
rect 205 -224 206 -206
rect 271 -224 272 -206
rect 282 -224 283 -206
rect 1066 -309 1067 -223
rect 159 -226 160 -206
rect 282 -309 283 -225
rect 310 -309 311 -225
rect 331 -309 332 -225
rect 362 -309 363 -225
rect 835 -309 836 -225
rect 926 -226 927 -206
rect 1052 -309 1053 -225
rect 198 -228 199 -206
rect 205 -309 206 -227
rect 233 -228 234 -206
rect 320 -228 321 -206
rect 415 -228 416 -206
rect 443 -309 444 -227
rect 457 -228 458 -206
rect 912 -309 913 -227
rect 947 -228 948 -206
rect 1129 -309 1130 -227
rect 177 -230 178 -206
rect 198 -309 199 -229
rect 233 -309 234 -229
rect 334 -230 335 -206
rect 408 -230 409 -206
rect 415 -309 416 -229
rect 425 -309 426 -229
rect 828 -309 829 -229
rect 947 -309 948 -229
rect 975 -230 976 -206
rect 54 -232 55 -206
rect 975 -309 976 -231
rect 177 -309 178 -233
rect 317 -234 318 -206
rect 320 -309 321 -233
rect 1136 -309 1137 -233
rect 240 -309 241 -235
rect 317 -309 318 -235
rect 429 -236 430 -206
rect 457 -309 458 -235
rect 506 -236 507 -206
rect 590 -309 591 -235
rect 607 -236 608 -206
rect 1073 -309 1074 -235
rect 124 -309 125 -237
rect 429 -309 430 -237
rect 513 -238 514 -206
rect 1115 -309 1116 -237
rect 261 -240 262 -206
rect 261 -309 262 -239
rect 261 -240 262 -206
rect 261 -309 262 -239
rect 268 -240 269 -206
rect 555 -240 556 -206
rect 579 -309 580 -239
rect 1143 -309 1144 -239
rect 128 -242 129 -206
rect 268 -309 269 -241
rect 373 -242 374 -206
rect 506 -309 507 -241
rect 513 -309 514 -241
rect 548 -242 549 -206
rect 607 -309 608 -241
rect 940 -242 941 -206
rect 954 -242 955 -206
rect 1094 -309 1095 -241
rect 26 -309 27 -243
rect 954 -309 955 -243
rect 961 -244 962 -206
rect 1010 -309 1011 -243
rect 128 -309 129 -245
rect 212 -246 213 -206
rect 219 -246 220 -206
rect 373 -309 374 -245
rect 408 -309 409 -245
rect 555 -309 556 -245
rect 632 -246 633 -206
rect 632 -309 633 -245
rect 632 -246 633 -206
rect 632 -309 633 -245
rect 639 -246 640 -206
rect 877 -309 878 -245
rect 919 -246 920 -206
rect 961 -309 962 -245
rect 968 -246 969 -206
rect 982 -246 983 -206
rect 170 -248 171 -206
rect 212 -309 213 -247
rect 219 -309 220 -247
rect 226 -248 227 -206
rect 401 -248 402 -206
rect 639 -309 640 -247
rect 674 -248 675 -206
rect 793 -309 794 -247
rect 800 -248 801 -206
rect 968 -309 969 -247
rect 978 -248 979 -206
rect 982 -309 983 -247
rect 40 -309 41 -249
rect 170 -309 171 -249
rect 345 -250 346 -206
rect 401 -309 402 -249
rect 492 -250 493 -206
rect 548 -309 549 -249
rect 576 -250 577 -206
rect 674 -309 675 -249
rect 688 -250 689 -206
rect 716 -250 717 -206
rect 719 -250 720 -206
rect 1003 -309 1004 -249
rect 86 -252 87 -206
rect 492 -309 493 -251
rect 516 -252 517 -206
rect 992 -252 993 -206
rect 58 -254 59 -206
rect 86 -309 87 -253
rect 163 -254 164 -206
rect 226 -309 227 -253
rect 327 -309 328 -253
rect 688 -309 689 -253
rect 695 -254 696 -206
rect 814 -309 815 -253
rect 58 -309 59 -255
rect 289 -256 290 -206
rect 345 -309 346 -255
rect 366 -256 367 -206
rect 534 -256 535 -206
rect 933 -256 934 -206
rect 23 -258 24 -206
rect 289 -309 290 -257
rect 359 -258 360 -206
rect 366 -309 367 -257
rect 534 -309 535 -257
rect 1153 -309 1154 -257
rect 163 -309 164 -259
rect 422 -260 423 -206
rect 576 -309 577 -259
rect 905 -260 906 -206
rect 191 -262 192 -206
rect 359 -309 360 -261
rect 618 -262 619 -206
rect 716 -309 717 -261
rect 737 -262 738 -206
rect 919 -309 920 -261
rect 33 -309 34 -263
rect 191 -309 192 -263
rect 562 -264 563 -206
rect 618 -309 619 -263
rect 625 -264 626 -206
rect 737 -309 738 -263
rect 744 -264 745 -206
rect 940 -309 941 -263
rect 541 -266 542 -206
rect 562 -309 563 -265
rect 583 -266 584 -206
rect 744 -309 745 -265
rect 758 -266 759 -206
rect 1024 -309 1025 -265
rect 380 -268 381 -206
rect 583 -309 584 -267
rect 611 -268 612 -206
rect 625 -309 626 -267
rect 667 -268 668 -206
rect 800 -309 801 -267
rect 884 -268 885 -206
rect 933 -309 934 -267
rect 121 -270 122 -206
rect 380 -309 381 -269
rect 527 -270 528 -206
rect 611 -309 612 -269
rect 698 -309 699 -269
rect 842 -309 843 -269
rect 121 -309 122 -271
rect 485 -309 486 -271
rect 499 -272 500 -206
rect 527 -309 528 -271
rect 541 -309 542 -271
rect 1031 -309 1032 -271
rect 142 -274 143 -206
rect 884 -309 885 -273
rect 114 -276 115 -206
rect 142 -309 143 -275
rect 296 -276 297 -206
rect 499 -309 500 -275
rect 702 -276 703 -206
rect 926 -309 927 -275
rect 114 -309 115 -277
rect 135 -278 136 -206
rect 296 -309 297 -277
rect 604 -309 605 -277
rect 705 -309 706 -277
rect 898 -278 899 -206
rect 135 -309 136 -279
rect 422 -309 423 -279
rect 709 -280 710 -206
rect 849 -309 850 -279
rect 352 -282 353 -206
rect 667 -309 668 -281
rect 730 -282 731 -206
rect 898 -309 899 -281
rect 93 -284 94 -206
rect 352 -309 353 -283
rect 520 -284 521 -206
rect 730 -309 731 -283
rect 758 -309 759 -283
rect 1038 -309 1039 -283
rect 9 -286 10 -206
rect 93 -309 94 -285
rect 478 -286 479 -206
rect 520 -309 521 -285
rect 597 -286 598 -206
rect 709 -309 710 -285
rect 765 -286 766 -206
rect 863 -309 864 -285
rect 9 -309 10 -287
rect 79 -288 80 -206
rect 184 -288 185 -206
rect 597 -309 598 -287
rect 779 -288 780 -206
rect 891 -309 892 -287
rect 184 -309 185 -289
rect 247 -290 248 -206
rect 390 -290 391 -206
rect 765 -309 766 -289
rect 779 -309 780 -289
rect 996 -290 997 -206
rect 247 -309 248 -291
rect 275 -292 276 -206
rect 450 -292 451 -206
rect 478 -309 479 -291
rect 786 -292 787 -206
rect 905 -309 906 -291
rect 254 -294 255 -206
rect 275 -309 276 -293
rect 450 -309 451 -293
rect 751 -294 752 -206
rect 856 -294 857 -206
rect 996 -309 997 -293
rect 254 -309 255 -295
rect 324 -296 325 -206
rect 646 -296 647 -206
rect 786 -309 787 -295
rect 324 -309 325 -297
rect 338 -298 339 -206
rect 569 -298 570 -206
rect 646 -309 647 -297
rect 681 -298 682 -206
rect 856 -309 857 -297
rect 68 -309 69 -299
rect 338 -309 339 -299
rect 653 -300 654 -206
rect 681 -309 682 -299
rect 723 -300 724 -206
rect 751 -309 752 -299
rect 156 -302 157 -206
rect 569 -309 570 -301
rect 653 -309 654 -301
rect 660 -302 661 -206
rect 723 -309 724 -301
rect 807 -302 808 -206
rect 149 -304 150 -206
rect 156 -309 157 -303
rect 660 -309 661 -303
rect 695 -309 696 -303
rect 772 -304 773 -206
rect 807 -309 808 -303
rect 30 -309 31 -305
rect 772 -309 773 -305
rect 54 -309 55 -307
rect 149 -309 150 -307
rect 2 -319 3 -317
rect 40 -398 41 -318
rect 65 -398 66 -318
rect 86 -319 87 -317
rect 93 -319 94 -317
rect 226 -319 227 -317
rect 264 -398 265 -318
rect 275 -319 276 -317
rect 285 -319 286 -317
rect 1192 -398 1193 -318
rect 1500 -319 1501 -317
rect 1500 -398 1501 -318
rect 1500 -319 1501 -317
rect 1500 -398 1501 -318
rect 2 -398 3 -320
rect 44 -321 45 -317
rect 58 -321 59 -317
rect 275 -398 276 -320
rect 310 -398 311 -320
rect 450 -321 451 -317
rect 471 -321 472 -317
rect 544 -321 545 -317
rect 586 -321 587 -317
rect 1059 -321 1060 -317
rect 1101 -321 1102 -317
rect 1171 -398 1172 -320
rect 1178 -321 1179 -317
rect 1202 -398 1203 -320
rect 9 -323 10 -317
rect 30 -398 31 -322
rect 37 -323 38 -317
rect 572 -398 573 -322
rect 604 -398 605 -322
rect 618 -323 619 -317
rect 681 -323 682 -317
rect 681 -398 682 -322
rect 681 -323 682 -317
rect 681 -398 682 -322
rect 688 -323 689 -317
rect 688 -398 689 -322
rect 688 -323 689 -317
rect 688 -398 689 -322
rect 695 -323 696 -317
rect 1101 -398 1102 -322
rect 1115 -323 1116 -317
rect 1178 -398 1179 -322
rect 9 -398 10 -324
rect 233 -325 234 -317
rect 317 -325 318 -317
rect 499 -325 500 -317
rect 527 -325 528 -317
rect 541 -398 542 -324
rect 702 -325 703 -317
rect 1164 -398 1165 -324
rect 16 -327 17 -317
rect 89 -398 90 -326
rect 93 -398 94 -326
rect 177 -327 178 -317
rect 184 -327 185 -317
rect 502 -398 503 -326
rect 702 -398 703 -326
rect 709 -327 710 -317
rect 758 -327 759 -317
rect 884 -327 885 -317
rect 912 -327 913 -317
rect 912 -398 913 -326
rect 912 -327 913 -317
rect 912 -398 913 -326
rect 961 -327 962 -317
rect 1185 -398 1186 -326
rect 16 -398 17 -328
rect 313 -329 314 -317
rect 327 -329 328 -317
rect 597 -329 598 -317
rect 667 -329 668 -317
rect 758 -398 759 -328
rect 842 -329 843 -317
rect 842 -398 843 -328
rect 842 -329 843 -317
rect 842 -398 843 -328
rect 856 -329 857 -317
rect 856 -398 857 -328
rect 856 -329 857 -317
rect 856 -398 857 -328
rect 863 -329 864 -317
rect 863 -398 864 -328
rect 863 -329 864 -317
rect 863 -398 864 -328
rect 884 -398 885 -328
rect 905 -329 906 -317
rect 1031 -329 1032 -317
rect 1059 -398 1060 -328
rect 1129 -329 1130 -317
rect 1150 -398 1151 -328
rect 26 -331 27 -317
rect 191 -331 192 -317
rect 198 -331 199 -317
rect 320 -331 321 -317
rect 359 -331 360 -317
rect 667 -398 668 -330
rect 709 -398 710 -330
rect 723 -331 724 -317
rect 891 -331 892 -317
rect 905 -398 906 -330
rect 996 -331 997 -317
rect 1031 -398 1032 -330
rect 1052 -331 1053 -317
rect 1115 -398 1116 -330
rect 1136 -331 1137 -317
rect 1157 -398 1158 -330
rect 37 -398 38 -332
rect 989 -333 990 -317
rect 1087 -333 1088 -317
rect 1129 -398 1130 -332
rect 44 -398 45 -334
rect 47 -398 48 -334
rect 61 -398 62 -334
rect 233 -398 234 -334
rect 254 -335 255 -317
rect 359 -398 360 -334
rect 394 -335 395 -317
rect 411 -335 412 -317
rect 422 -335 423 -317
rect 478 -335 479 -317
rect 485 -335 486 -317
rect 618 -398 619 -334
rect 653 -335 654 -317
rect 723 -398 724 -334
rect 765 -335 766 -317
rect 996 -398 997 -334
rect 1024 -335 1025 -317
rect 1087 -398 1088 -334
rect 1094 -335 1095 -317
rect 1136 -398 1137 -334
rect 68 -337 69 -317
rect 730 -337 731 -317
rect 786 -337 787 -317
rect 891 -398 892 -336
rect 947 -337 948 -317
rect 1052 -398 1053 -336
rect 72 -339 73 -317
rect 82 -339 83 -317
rect 107 -339 108 -317
rect 110 -349 111 -338
rect 121 -339 122 -317
rect 590 -339 591 -317
rect 625 -339 626 -317
rect 765 -398 766 -338
rect 786 -398 787 -338
rect 814 -339 815 -317
rect 940 -339 941 -317
rect 947 -398 948 -338
rect 982 -339 983 -317
rect 989 -398 990 -338
rect 1045 -339 1046 -317
rect 1094 -398 1095 -338
rect 75 -398 76 -340
rect 1143 -341 1144 -317
rect 79 -343 80 -317
rect 1024 -398 1025 -342
rect 1122 -343 1123 -317
rect 1143 -398 1144 -342
rect 82 -398 83 -344
rect 1066 -345 1067 -317
rect 1073 -345 1074 -317
rect 1122 -398 1123 -344
rect 107 -398 108 -346
rect 135 -347 136 -317
rect 156 -347 157 -317
rect 453 -347 454 -317
rect 471 -398 472 -346
rect 492 -347 493 -317
rect 499 -398 500 -346
rect 562 -347 563 -317
rect 569 -347 570 -317
rect 730 -398 731 -346
rect 814 -398 815 -346
rect 821 -347 822 -317
rect 898 -347 899 -317
rect 940 -398 941 -346
rect 968 -347 969 -317
rect 982 -398 983 -346
rect 1017 -347 1018 -317
rect 1045 -398 1046 -346
rect 135 -398 136 -348
rect 163 -349 164 -317
rect 478 -398 479 -348
rect 516 -398 517 -348
rect 898 -398 899 -348
rect 954 -349 955 -317
rect 968 -398 969 -348
rect 975 -349 976 -317
rect 1017 -398 1018 -348
rect 1038 -349 1039 -317
rect 1066 -398 1067 -348
rect 96 -351 97 -317
rect 954 -398 955 -350
rect 1003 -351 1004 -317
rect 1038 -398 1039 -350
rect 100 -353 101 -317
rect 163 -398 164 -352
rect 177 -398 178 -352
rect 282 -353 283 -317
rect 303 -353 304 -317
rect 317 -398 318 -352
rect 331 -353 332 -317
rect 422 -398 423 -352
rect 429 -353 430 -317
rect 527 -398 528 -352
rect 555 -353 556 -317
rect 597 -398 598 -352
rect 625 -398 626 -352
rect 632 -353 633 -317
rect 653 -398 654 -352
rect 674 -353 675 -317
rect 800 -353 801 -317
rect 821 -398 822 -352
rect 926 -353 927 -317
rect 975 -398 976 -352
rect 51 -355 52 -317
rect 100 -398 101 -354
rect 114 -355 115 -317
rect 121 -398 122 -354
rect 128 -355 129 -317
rect 184 -398 185 -354
rect 191 -398 192 -354
rect 212 -355 213 -317
rect 219 -355 220 -317
rect 226 -398 227 -354
rect 282 -398 283 -354
rect 373 -355 374 -317
rect 380 -355 381 -317
rect 485 -398 486 -354
rect 509 -398 510 -354
rect 632 -398 633 -354
rect 674 -398 675 -354
rect 779 -355 780 -317
rect 800 -398 801 -354
rect 1209 -398 1210 -354
rect 72 -398 73 -356
rect 114 -398 115 -356
rect 128 -398 129 -356
rect 611 -357 612 -317
rect 779 -398 780 -356
rect 807 -357 808 -317
rect 919 -357 920 -317
rect 926 -398 927 -356
rect 933 -357 934 -317
rect 1003 -398 1004 -356
rect 142 -359 143 -317
rect 219 -398 220 -358
rect 303 -398 304 -358
rect 352 -359 353 -317
rect 366 -359 367 -317
rect 380 -398 381 -358
rect 397 -398 398 -358
rect 1080 -359 1081 -317
rect 86 -398 87 -360
rect 142 -398 143 -360
rect 198 -398 199 -360
rect 205 -361 206 -317
rect 212 -398 213 -360
rect 698 -361 699 -317
rect 772 -361 773 -317
rect 807 -398 808 -360
rect 849 -361 850 -317
rect 933 -398 934 -360
rect 1010 -361 1011 -317
rect 1080 -398 1081 -360
rect 149 -363 150 -317
rect 205 -398 206 -362
rect 289 -363 290 -317
rect 352 -398 353 -362
rect 366 -398 367 -362
rect 642 -398 643 -362
rect 772 -398 773 -362
rect 793 -363 794 -317
rect 828 -363 829 -317
rect 849 -398 850 -362
rect 870 -363 871 -317
rect 919 -398 920 -362
rect 1010 -398 1011 -362
rect 1108 -363 1109 -317
rect 79 -398 80 -364
rect 828 -398 829 -364
rect 149 -398 150 -366
rect 247 -367 248 -317
rect 289 -398 290 -366
rect 551 -398 552 -366
rect 569 -398 570 -366
rect 877 -367 878 -317
rect 247 -398 248 -368
rect 268 -369 269 -317
rect 373 -398 374 -368
rect 520 -369 521 -317
rect 583 -369 584 -317
rect 793 -398 794 -368
rect 835 -369 836 -317
rect 877 -398 878 -368
rect 23 -371 24 -317
rect 835 -398 836 -370
rect 23 -398 24 -372
rect 33 -373 34 -317
rect 261 -373 262 -317
rect 268 -398 269 -372
rect 387 -373 388 -317
rect 1108 -398 1109 -372
rect 261 -398 262 -374
rect 506 -375 507 -317
rect 513 -375 514 -317
rect 555 -398 556 -374
rect 583 -398 584 -374
rect 660 -375 661 -317
rect 751 -375 752 -317
rect 870 -398 871 -374
rect 331 -398 332 -376
rect 660 -398 661 -376
rect 737 -377 738 -317
rect 751 -398 752 -376
rect 345 -379 346 -317
rect 387 -398 388 -378
rect 401 -379 402 -317
rect 401 -398 402 -378
rect 401 -379 402 -317
rect 401 -398 402 -378
rect 408 -379 409 -317
rect 961 -398 962 -378
rect 51 -398 52 -380
rect 408 -398 409 -380
rect 415 -381 416 -317
rect 429 -398 430 -380
rect 436 -381 437 -317
rect 695 -398 696 -380
rect 296 -383 297 -317
rect 345 -398 346 -382
rect 415 -398 416 -382
rect 670 -398 671 -382
rect 124 -385 125 -317
rect 296 -398 297 -384
rect 338 -385 339 -317
rect 436 -398 437 -384
rect 450 -398 451 -384
rect 457 -385 458 -317
rect 464 -385 465 -317
rect 492 -398 493 -384
rect 506 -398 507 -384
rect 744 -385 745 -317
rect 124 -398 125 -386
rect 156 -398 157 -386
rect 338 -398 339 -386
rect 576 -387 577 -317
rect 579 -387 580 -317
rect 737 -398 738 -386
rect 324 -389 325 -317
rect 576 -398 577 -388
rect 590 -398 591 -388
rect 1073 -398 1074 -388
rect 240 -391 241 -317
rect 324 -398 325 -390
rect 443 -391 444 -317
rect 457 -398 458 -390
rect 464 -398 465 -390
rect 513 -398 514 -390
rect 520 -398 521 -390
rect 534 -391 535 -317
rect 611 -398 612 -390
rect 646 -391 647 -317
rect 716 -391 717 -317
rect 744 -398 745 -390
rect 58 -398 59 -392
rect 240 -398 241 -392
rect 411 -398 412 -392
rect 716 -398 717 -392
rect 170 -395 171 -317
rect 443 -398 444 -394
rect 534 -398 535 -394
rect 548 -395 549 -317
rect 639 -395 640 -317
rect 646 -398 647 -394
rect 26 -398 27 -396
rect 170 -398 171 -396
rect 254 -398 255 -396
rect 548 -398 549 -396
rect 565 -398 566 -396
rect 639 -398 640 -396
rect 23 -408 24 -406
rect 1108 -408 1109 -406
rect 1129 -408 1130 -406
rect 1213 -513 1214 -407
rect 1500 -408 1501 -406
rect 1500 -513 1501 -407
rect 1500 -408 1501 -406
rect 1500 -513 1501 -407
rect 23 -513 24 -409
rect 264 -410 265 -406
rect 331 -410 332 -406
rect 537 -513 538 -409
rect 541 -410 542 -406
rect 541 -513 542 -409
rect 541 -410 542 -406
rect 541 -513 542 -409
rect 548 -410 549 -406
rect 1171 -410 1172 -406
rect 1209 -410 1210 -406
rect 1395 -513 1396 -409
rect 26 -412 27 -406
rect 975 -412 976 -406
rect 1017 -412 1018 -406
rect 1206 -513 1207 -411
rect 30 -414 31 -406
rect 58 -414 59 -406
rect 75 -414 76 -406
rect 121 -513 122 -413
rect 128 -414 129 -406
rect 383 -513 384 -413
rect 408 -414 409 -406
rect 429 -414 430 -406
rect 460 -513 461 -413
rect 919 -414 920 -406
rect 975 -513 976 -413
rect 1202 -414 1203 -406
rect 30 -513 31 -415
rect 940 -416 941 -406
rect 1038 -416 1039 -406
rect 1129 -513 1130 -415
rect 1136 -416 1137 -406
rect 1220 -513 1221 -415
rect 40 -513 41 -417
rect 282 -418 283 -406
rect 331 -513 332 -417
rect 653 -418 654 -406
rect 663 -418 664 -406
rect 1178 -418 1179 -406
rect 44 -420 45 -406
rect 177 -420 178 -406
rect 201 -513 202 -419
rect 205 -420 206 -406
rect 261 -420 262 -406
rect 387 -420 388 -406
rect 401 -420 402 -406
rect 429 -513 430 -419
rect 471 -420 472 -406
rect 513 -513 514 -419
rect 551 -420 552 -406
rect 807 -420 808 -406
rect 814 -420 815 -406
rect 817 -464 818 -419
rect 870 -420 871 -406
rect 940 -513 941 -419
rect 968 -420 969 -406
rect 1038 -513 1039 -419
rect 1045 -420 1046 -406
rect 1136 -513 1137 -419
rect 1143 -420 1144 -406
rect 1227 -513 1228 -419
rect 2 -422 3 -406
rect 44 -513 45 -421
rect 58 -513 59 -421
rect 65 -422 66 -406
rect 79 -422 80 -406
rect 919 -513 920 -421
rect 961 -422 962 -406
rect 1045 -513 1046 -421
rect 1059 -422 1060 -406
rect 1143 -513 1144 -421
rect 1150 -422 1151 -406
rect 1234 -513 1235 -421
rect 9 -424 10 -406
rect 79 -513 80 -423
rect 86 -424 87 -406
rect 177 -513 178 -423
rect 198 -424 199 -406
rect 205 -513 206 -423
rect 261 -513 262 -423
rect 373 -424 374 -406
rect 401 -513 402 -423
rect 611 -424 612 -406
rect 625 -424 626 -406
rect 639 -513 640 -423
rect 670 -424 671 -406
rect 1052 -424 1053 -406
rect 1066 -424 1067 -406
rect 1150 -513 1151 -423
rect 1157 -424 1158 -406
rect 1255 -513 1256 -423
rect 61 -426 62 -406
rect 1178 -513 1179 -425
rect 65 -513 66 -427
rect 555 -428 556 -406
rect 562 -428 563 -406
rect 877 -428 878 -406
rect 898 -428 899 -406
rect 961 -513 962 -427
rect 982 -428 983 -406
rect 1066 -513 1067 -427
rect 1073 -428 1074 -406
rect 1157 -513 1158 -427
rect 47 -430 48 -406
rect 877 -513 878 -429
rect 884 -430 885 -406
rect 898 -513 899 -429
rect 905 -430 906 -406
rect 968 -513 969 -429
rect 1003 -430 1004 -406
rect 1059 -513 1060 -429
rect 1080 -430 1081 -406
rect 1171 -513 1172 -429
rect 86 -513 87 -431
rect 219 -432 220 -406
rect 275 -432 276 -406
rect 387 -513 388 -431
rect 411 -432 412 -406
rect 464 -432 465 -406
rect 478 -432 479 -406
rect 516 -432 517 -406
rect 520 -432 521 -406
rect 555 -513 556 -431
rect 569 -432 570 -406
rect 933 -432 934 -406
rect 1003 -513 1004 -431
rect 1010 -432 1011 -406
rect 89 -434 90 -406
rect 1241 -513 1242 -433
rect 89 -513 90 -435
rect 821 -436 822 -406
rect 828 -436 829 -406
rect 982 -513 983 -435
rect 989 -436 990 -406
rect 1010 -513 1011 -435
rect 93 -438 94 -406
rect 124 -438 125 -406
rect 138 -513 139 -437
rect 1192 -438 1193 -406
rect 72 -513 73 -439
rect 93 -513 94 -439
rect 100 -440 101 -406
rect 408 -513 409 -439
rect 422 -440 423 -406
rect 464 -513 465 -439
rect 478 -513 479 -439
rect 758 -440 759 -406
rect 772 -440 773 -406
rect 821 -513 822 -439
rect 835 -440 836 -406
rect 905 -513 906 -439
rect 1122 -440 1123 -406
rect 1192 -513 1193 -439
rect 33 -513 34 -441
rect 772 -513 773 -441
rect 779 -442 780 -406
rect 835 -513 836 -441
rect 849 -442 850 -406
rect 870 -513 871 -441
rect 1031 -442 1032 -406
rect 1122 -513 1123 -441
rect 100 -513 101 -443
rect 142 -444 143 -406
rect 145 -513 146 -443
rect 828 -513 829 -443
rect 863 -444 864 -406
rect 933 -513 934 -443
rect 107 -446 108 -406
rect 128 -513 129 -445
rect 142 -513 143 -445
rect 184 -446 185 -406
rect 198 -513 199 -445
rect 576 -446 577 -406
rect 590 -446 591 -406
rect 663 -513 664 -445
rect 698 -513 699 -445
rect 1017 -513 1018 -445
rect 107 -513 108 -447
rect 884 -513 885 -447
rect 156 -450 157 -406
rect 548 -513 549 -449
rect 572 -450 573 -406
rect 863 -513 864 -449
rect 163 -452 164 -406
rect 282 -513 283 -451
rect 338 -452 339 -406
rect 562 -513 563 -451
rect 576 -513 577 -451
rect 618 -452 619 -406
rect 632 -452 633 -406
rect 653 -513 654 -451
rect 705 -513 706 -451
rect 1185 -452 1186 -406
rect 170 -454 171 -406
rect 569 -513 570 -453
rect 593 -454 594 -406
rect 695 -454 696 -406
rect 716 -454 717 -406
rect 779 -513 780 -453
rect 793 -454 794 -406
rect 1031 -513 1032 -453
rect 1101 -454 1102 -406
rect 1185 -513 1186 -453
rect 149 -456 150 -406
rect 170 -513 171 -455
rect 184 -513 185 -455
rect 310 -456 311 -406
rect 338 -513 339 -455
rect 492 -456 493 -406
rect 509 -513 510 -455
rect 765 -456 766 -406
rect 800 -456 801 -406
rect 849 -513 850 -455
rect 114 -458 115 -406
rect 765 -513 766 -457
rect 814 -513 815 -457
rect 926 -458 927 -406
rect 114 -513 115 -459
rect 289 -460 290 -406
rect 310 -513 311 -459
rect 317 -460 318 -406
rect 345 -460 346 -406
rect 807 -513 808 -459
rect 856 -460 857 -406
rect 926 -513 927 -459
rect 51 -462 52 -406
rect 289 -513 290 -461
rect 296 -462 297 -406
rect 345 -513 346 -461
rect 373 -513 374 -461
rect 450 -462 451 -406
rect 457 -462 458 -406
rect 471 -513 472 -461
rect 485 -462 486 -406
rect 492 -513 493 -461
rect 520 -513 521 -461
rect 583 -462 584 -406
rect 597 -462 598 -406
rect 632 -513 633 -461
rect 642 -462 643 -406
rect 989 -513 990 -461
rect 51 -513 52 -463
rect 380 -464 381 -406
rect 422 -513 423 -463
rect 793 -513 794 -463
rect 856 -513 857 -463
rect 149 -513 150 -465
rect 240 -466 241 -406
rect 268 -466 269 -406
rect 275 -513 276 -465
rect 296 -513 297 -465
rect 397 -466 398 -406
rect 425 -513 426 -465
rect 1073 -513 1074 -465
rect 212 -468 213 -406
rect 268 -513 269 -467
rect 366 -468 367 -406
rect 450 -513 451 -467
rect 457 -513 458 -467
rect 590 -513 591 -467
rect 597 -513 598 -467
rect 1248 -513 1249 -467
rect 212 -513 213 -469
rect 233 -470 234 -406
rect 366 -513 367 -469
rect 506 -513 507 -469
rect 534 -470 535 -406
rect 583 -513 584 -469
rect 600 -513 601 -469
rect 996 -470 997 -406
rect 219 -513 220 -471
rect 324 -472 325 -406
rect 380 -513 381 -471
rect 1080 -513 1081 -471
rect 226 -474 227 -406
rect 240 -513 241 -473
rect 303 -474 304 -406
rect 324 -513 325 -473
rect 436 -474 437 -406
rect 485 -513 486 -473
rect 604 -474 605 -406
rect 625 -513 626 -473
rect 646 -474 647 -406
rect 1101 -513 1102 -473
rect 16 -476 17 -406
rect 303 -513 304 -475
rect 317 -513 318 -475
rect 534 -513 535 -475
rect 611 -513 612 -475
rect 1087 -476 1088 -406
rect 16 -513 17 -477
rect 247 -478 248 -406
rect 352 -478 353 -406
rect 436 -513 437 -477
rect 527 -478 528 -406
rect 604 -513 605 -477
rect 614 -513 615 -477
rect 1052 -513 1053 -477
rect 82 -480 83 -406
rect 646 -513 647 -479
rect 681 -480 682 -406
rect 716 -513 717 -479
rect 737 -480 738 -406
rect 758 -513 759 -479
rect 912 -480 913 -406
rect 996 -513 997 -479
rect 1024 -480 1025 -406
rect 1087 -513 1088 -479
rect 159 -513 160 -481
rect 912 -513 913 -481
rect 947 -482 948 -406
rect 1024 -513 1025 -481
rect 191 -484 192 -406
rect 226 -513 227 -483
rect 233 -513 234 -483
rect 394 -484 395 -406
rect 499 -484 500 -406
rect 681 -513 682 -483
rect 751 -484 752 -406
rect 800 -513 801 -483
rect 891 -484 892 -406
rect 947 -513 948 -483
rect 135 -486 136 -406
rect 191 -513 192 -485
rect 254 -486 255 -406
rect 394 -513 395 -485
rect 527 -513 528 -485
rect 1108 -513 1109 -485
rect 135 -513 136 -487
rect 954 -488 955 -406
rect 37 -490 38 -406
rect 954 -513 955 -489
rect 37 -513 38 -491
rect 75 -513 76 -491
rect 163 -513 164 -491
rect 499 -513 500 -491
rect 565 -492 566 -406
rect 737 -513 738 -491
rect 842 -492 843 -406
rect 891 -513 892 -491
rect 352 -513 353 -493
rect 359 -494 360 -406
rect 618 -513 619 -493
rect 674 -494 675 -406
rect 702 -494 703 -406
rect 751 -513 752 -493
rect 786 -494 787 -406
rect 842 -513 843 -493
rect 110 -513 111 -495
rect 359 -513 360 -495
rect 415 -496 416 -406
rect 702 -513 703 -495
rect 730 -496 731 -406
rect 786 -513 787 -495
rect 415 -513 416 -497
rect 1164 -498 1165 -406
rect 502 -500 503 -406
rect 674 -513 675 -499
rect 688 -500 689 -406
rect 730 -513 731 -499
rect 1094 -500 1095 -406
rect 1164 -513 1165 -499
rect 9 -513 10 -501
rect 502 -513 503 -501
rect 688 -513 689 -501
rect 723 -502 724 -406
rect 1094 -513 1095 -501
rect 1115 -502 1116 -406
rect 723 -513 724 -503
rect 744 -504 745 -406
rect 1115 -513 1116 -503
rect 1199 -504 1200 -406
rect 667 -506 668 -406
rect 1199 -513 1200 -505
rect 660 -508 661 -406
rect 667 -513 668 -507
rect 709 -508 710 -406
rect 744 -513 745 -507
rect 443 -510 444 -406
rect 709 -513 710 -509
rect 443 -513 444 -511
rect 530 -513 531 -511
rect 660 -513 661 -511
rect 1262 -513 1263 -511
rect 2 -523 3 -521
rect 1241 -523 1242 -521
rect 1248 -523 1249 -521
rect 1360 -628 1361 -522
rect 1395 -523 1396 -521
rect 1472 -628 1473 -522
rect 1500 -523 1501 -521
rect 1507 -628 1508 -522
rect 2 -628 3 -524
rect 565 -628 566 -524
rect 600 -525 601 -521
rect 1269 -628 1270 -524
rect 16 -527 17 -521
rect 254 -527 255 -521
rect 261 -527 262 -521
rect 457 -527 458 -521
rect 460 -527 461 -521
rect 919 -527 920 -521
rect 1003 -527 1004 -521
rect 1339 -628 1340 -526
rect 30 -628 31 -528
rect 583 -529 584 -521
rect 635 -628 636 -528
rect 758 -529 759 -521
rect 828 -529 829 -521
rect 919 -628 920 -528
rect 940 -529 941 -521
rect 1003 -628 1004 -528
rect 1087 -529 1088 -521
rect 1087 -628 1088 -528
rect 1087 -529 1088 -521
rect 1087 -628 1088 -528
rect 1094 -529 1095 -521
rect 1283 -628 1284 -528
rect 33 -531 34 -521
rect 72 -531 73 -521
rect 75 -628 76 -530
rect 219 -531 220 -521
rect 226 -531 227 -521
rect 380 -531 381 -521
rect 425 -531 426 -521
rect 614 -531 615 -521
rect 639 -531 640 -521
rect 639 -628 640 -530
rect 639 -531 640 -521
rect 639 -628 640 -530
rect 660 -531 661 -521
rect 814 -531 815 -521
rect 870 -531 871 -521
rect 940 -628 941 -530
rect 1024 -531 1025 -521
rect 1094 -628 1095 -530
rect 1150 -531 1151 -521
rect 1241 -628 1242 -530
rect 1255 -531 1256 -521
rect 1374 -628 1375 -530
rect 40 -533 41 -521
rect 1206 -533 1207 -521
rect 1213 -533 1214 -521
rect 1304 -628 1305 -532
rect 40 -628 41 -534
rect 1073 -535 1074 -521
rect 1080 -535 1081 -521
rect 1150 -628 1151 -534
rect 1157 -535 1158 -521
rect 1248 -628 1249 -534
rect 1262 -535 1263 -521
rect 1367 -628 1368 -534
rect 47 -628 48 -536
rect 198 -537 199 -521
rect 226 -628 227 -536
rect 275 -537 276 -521
rect 317 -537 318 -521
rect 611 -537 612 -521
rect 614 -628 615 -536
rect 821 -537 822 -521
rect 954 -537 955 -521
rect 1024 -628 1025 -536
rect 1136 -537 1137 -521
rect 1213 -628 1214 -536
rect 1220 -537 1221 -521
rect 1311 -628 1312 -536
rect 72 -628 73 -538
rect 233 -539 234 -521
rect 240 -539 241 -521
rect 261 -628 262 -538
rect 271 -628 272 -538
rect 807 -539 808 -521
rect 912 -539 913 -521
rect 954 -628 955 -538
rect 996 -539 997 -521
rect 1073 -628 1074 -538
rect 1164 -539 1165 -521
rect 1206 -628 1207 -538
rect 1227 -539 1228 -521
rect 1332 -628 1333 -538
rect 110 -541 111 -521
rect 492 -541 493 -521
rect 499 -541 500 -521
rect 1157 -628 1158 -540
rect 1171 -541 1172 -521
rect 1276 -628 1277 -540
rect 114 -543 115 -521
rect 317 -628 318 -542
rect 331 -543 332 -521
rect 509 -543 510 -521
rect 520 -543 521 -521
rect 527 -628 528 -542
rect 530 -543 531 -521
rect 751 -543 752 -521
rect 779 -543 780 -521
rect 828 -628 829 -542
rect 842 -543 843 -521
rect 912 -628 913 -542
rect 933 -543 934 -521
rect 996 -628 997 -542
rect 1017 -543 1018 -521
rect 1080 -628 1081 -542
rect 1108 -543 1109 -521
rect 1164 -628 1165 -542
rect 1178 -543 1179 -521
rect 1255 -628 1256 -542
rect 114 -628 115 -544
rect 1325 -628 1326 -544
rect 117 -628 118 -546
rect 401 -547 402 -521
rect 408 -547 409 -521
rect 499 -628 500 -546
rect 502 -547 503 -521
rect 1101 -547 1102 -521
rect 1122 -547 1123 -521
rect 1171 -628 1172 -546
rect 1185 -547 1186 -521
rect 1262 -628 1263 -546
rect 135 -549 136 -521
rect 1045 -549 1046 -521
rect 1192 -549 1193 -521
rect 1290 -628 1291 -548
rect 121 -551 122 -521
rect 135 -628 136 -550
rect 142 -551 143 -521
rect 877 -551 878 -521
rect 898 -551 899 -521
rect 1192 -628 1193 -550
rect 1199 -551 1200 -521
rect 1297 -628 1298 -550
rect 121 -628 122 -552
rect 247 -553 248 -521
rect 275 -628 276 -552
rect 383 -553 384 -521
rect 401 -628 402 -552
rect 569 -553 570 -521
rect 611 -628 612 -552
rect 1136 -628 1137 -552
rect 1234 -553 1235 -521
rect 1353 -628 1354 -552
rect 44 -555 45 -521
rect 569 -628 570 -554
rect 625 -555 626 -521
rect 751 -628 752 -554
rect 765 -555 766 -521
rect 1178 -628 1179 -554
rect 142 -628 143 -556
rect 201 -557 202 -521
rect 212 -557 213 -521
rect 331 -628 332 -556
rect 338 -557 339 -521
rect 415 -557 416 -521
rect 443 -557 444 -521
rect 492 -628 493 -556
rect 509 -628 510 -556
rect 842 -628 843 -556
rect 849 -557 850 -521
rect 898 -628 899 -556
rect 968 -557 969 -521
rect 1045 -628 1046 -556
rect 1129 -557 1130 -521
rect 1199 -628 1200 -556
rect 58 -559 59 -521
rect 415 -628 416 -558
rect 450 -559 451 -521
rect 453 -589 454 -558
rect 457 -628 458 -558
rect 562 -559 563 -521
rect 625 -628 626 -558
rect 1318 -628 1319 -558
rect 37 -561 38 -521
rect 58 -628 59 -560
rect 138 -561 139 -521
rect 212 -628 213 -560
rect 233 -628 234 -560
rect 310 -561 311 -521
rect 338 -628 339 -560
rect 373 -561 374 -521
rect 450 -628 451 -560
rect 513 -561 514 -521
rect 534 -561 535 -521
rect 1185 -628 1186 -560
rect 79 -563 80 -521
rect 534 -628 535 -562
rect 548 -563 549 -521
rect 583 -628 584 -562
rect 628 -628 629 -562
rect 1108 -628 1109 -562
rect 1143 -563 1144 -521
rect 1234 -628 1235 -562
rect 65 -565 66 -521
rect 548 -628 549 -564
rect 660 -628 661 -564
rect 905 -565 906 -521
rect 1031 -565 1032 -521
rect 1101 -628 1102 -564
rect 65 -628 66 -566
rect 163 -567 164 -521
rect 170 -567 171 -521
rect 254 -628 255 -566
rect 345 -567 346 -521
rect 422 -567 423 -521
rect 464 -567 465 -521
rect 520 -628 521 -566
rect 663 -567 664 -521
rect 779 -628 780 -566
rect 786 -567 787 -521
rect 821 -628 822 -566
rect 835 -567 836 -521
rect 905 -628 906 -566
rect 1031 -628 1032 -566
rect 1346 -628 1347 -566
rect 5 -569 6 -521
rect 422 -628 423 -568
rect 481 -628 482 -568
rect 982 -569 983 -521
rect 1052 -569 1053 -521
rect 1129 -628 1130 -568
rect 23 -571 24 -521
rect 464 -628 465 -570
rect 485 -571 486 -521
rect 513 -628 514 -570
rect 670 -628 671 -570
rect 1115 -571 1116 -521
rect 23 -628 24 -572
rect 324 -573 325 -521
rect 348 -628 349 -572
rect 968 -628 969 -572
rect 1010 -573 1011 -521
rect 1052 -628 1053 -572
rect 1059 -573 1060 -521
rect 1143 -628 1144 -572
rect 79 -628 80 -574
rect 100 -575 101 -521
rect 107 -575 108 -521
rect 982 -628 983 -574
rect 989 -575 990 -521
rect 1059 -628 1060 -574
rect 96 -628 97 -576
rect 100 -628 101 -576
rect 107 -628 108 -576
rect 159 -577 160 -521
rect 163 -628 164 -576
rect 184 -577 185 -521
rect 191 -577 192 -521
rect 198 -628 199 -576
rect 240 -628 241 -576
rect 268 -577 269 -521
rect 324 -628 325 -576
rect 471 -577 472 -521
rect 506 -577 507 -521
rect 849 -628 850 -576
rect 863 -577 864 -521
rect 933 -628 934 -576
rect 947 -577 948 -521
rect 1010 -628 1011 -576
rect 19 -628 20 -578
rect 184 -628 185 -578
rect 191 -628 192 -578
rect 205 -579 206 -521
rect 247 -628 248 -578
rect 257 -579 258 -521
rect 268 -628 269 -578
rect 705 -579 706 -521
rect 723 -579 724 -521
rect 870 -628 871 -578
rect 884 -579 885 -521
rect 947 -628 948 -578
rect 145 -581 146 -521
rect 793 -581 794 -521
rect 800 -581 801 -521
rect 877 -628 878 -580
rect 926 -581 927 -521
rect 989 -628 990 -580
rect 170 -628 171 -582
rect 219 -628 220 -582
rect 250 -583 251 -521
rect 786 -628 787 -582
rect 856 -583 857 -521
rect 926 -628 927 -582
rect 86 -585 87 -521
rect 856 -628 857 -584
rect 86 -628 87 -586
rect 555 -587 556 -521
rect 618 -587 619 -521
rect 1115 -628 1116 -586
rect 177 -589 178 -521
rect 177 -628 178 -588
rect 177 -589 178 -521
rect 177 -628 178 -588
rect 205 -628 206 -588
rect 303 -589 304 -521
rect 352 -589 353 -521
rect 446 -628 447 -588
rect 485 -628 486 -588
rect 506 -628 507 -588
rect 975 -589 976 -521
rect 282 -591 283 -521
rect 618 -628 619 -590
rect 674 -591 675 -521
rect 1220 -628 1221 -590
rect 51 -593 52 -521
rect 282 -628 283 -592
rect 303 -628 304 -592
rect 352 -628 353 -592
rect 359 -593 360 -521
rect 408 -628 409 -592
rect 436 -593 437 -521
rect 674 -628 675 -592
rect 681 -593 682 -521
rect 758 -628 759 -592
rect 765 -628 766 -592
rect 1038 -593 1039 -521
rect 359 -628 360 -594
rect 387 -595 388 -521
rect 418 -595 419 -521
rect 436 -628 437 -594
rect 471 -628 472 -594
rect 562 -628 563 -594
rect 590 -595 591 -521
rect 681 -628 682 -594
rect 688 -595 689 -521
rect 723 -628 724 -594
rect 730 -595 731 -521
rect 800 -628 801 -594
rect 891 -595 892 -521
rect 975 -628 976 -594
rect 89 -597 90 -521
rect 891 -628 892 -596
rect 961 -597 962 -521
rect 1038 -628 1039 -596
rect 289 -599 290 -521
rect 387 -628 388 -598
rect 418 -628 419 -598
rect 1122 -628 1123 -598
rect 289 -628 290 -600
rect 394 -601 395 -521
rect 443 -628 444 -600
rect 590 -628 591 -600
rect 646 -601 647 -521
rect 730 -628 731 -600
rect 737 -601 738 -521
rect 807 -628 808 -600
rect 863 -628 864 -600
rect 961 -628 962 -600
rect 373 -628 374 -602
rect 597 -603 598 -521
rect 653 -603 654 -521
rect 737 -628 738 -602
rect 744 -603 745 -521
rect 814 -628 815 -602
rect 394 -628 395 -604
rect 429 -605 430 -521
rect 478 -605 479 -521
rect 597 -628 598 -604
rect 653 -628 654 -604
rect 709 -605 710 -521
rect 716 -605 717 -521
rect 793 -628 794 -604
rect 44 -628 45 -606
rect 709 -628 710 -606
rect 747 -628 748 -606
rect 884 -628 885 -606
rect 149 -609 150 -521
rect 429 -628 430 -608
rect 541 -609 542 -521
rect 555 -628 556 -608
rect 576 -609 577 -521
rect 646 -628 647 -608
rect 667 -609 668 -521
rect 688 -628 689 -608
rect 695 -609 696 -521
rect 1066 -609 1067 -521
rect 37 -628 38 -610
rect 576 -628 577 -610
rect 632 -611 633 -521
rect 716 -628 717 -610
rect 772 -611 773 -521
rect 835 -628 836 -610
rect 149 -628 150 -612
rect 380 -628 381 -612
rect 390 -628 391 -612
rect 1066 -628 1067 -612
rect 366 -615 367 -521
rect 541 -628 542 -614
rect 632 -628 633 -614
rect 695 -628 696 -614
rect 702 -615 703 -521
rect 1227 -628 1228 -614
rect 156 -617 157 -521
rect 702 -628 703 -616
rect 772 -628 773 -616
rect 1034 -628 1035 -616
rect 128 -619 129 -521
rect 156 -628 157 -618
rect 296 -619 297 -521
rect 366 -628 367 -618
rect 667 -628 668 -618
rect 1017 -628 1018 -618
rect 9 -621 10 -521
rect 296 -628 297 -620
rect 9 -628 10 -622
rect 604 -623 605 -521
rect 93 -625 94 -521
rect 128 -628 129 -624
rect 604 -628 605 -624
rect 698 -625 699 -521
rect 51 -628 52 -626
rect 93 -628 94 -626
rect 16 -638 17 -636
rect 16 -747 17 -637
rect 16 -638 17 -636
rect 16 -747 17 -637
rect 37 -747 38 -637
rect 324 -638 325 -636
rect 383 -638 384 -636
rect 730 -638 731 -636
rect 747 -638 748 -636
rect 996 -638 997 -636
rect 1034 -638 1035 -636
rect 1374 -638 1375 -636
rect 1472 -638 1473 -636
rect 1528 -747 1529 -637
rect 2 -640 3 -636
rect 324 -747 325 -639
rect 387 -640 388 -636
rect 450 -640 451 -636
rect 506 -640 507 -636
rect 772 -640 773 -636
rect 807 -640 808 -636
rect 1437 -747 1438 -639
rect 1507 -640 1508 -636
rect 1514 -747 1515 -639
rect 5 -747 6 -641
rect 1472 -747 1473 -641
rect 44 -644 45 -636
rect 1178 -644 1179 -636
rect 1206 -644 1207 -636
rect 1381 -747 1382 -643
rect 44 -747 45 -645
rect 233 -646 234 -636
rect 282 -646 283 -636
rect 345 -646 346 -636
rect 387 -747 388 -645
rect 541 -646 542 -636
rect 544 -747 545 -645
rect 1451 -747 1452 -645
rect 47 -648 48 -636
rect 422 -648 423 -636
rect 443 -648 444 -636
rect 548 -648 549 -636
rect 614 -648 615 -636
rect 751 -648 752 -636
rect 807 -747 808 -647
rect 926 -648 927 -636
rect 940 -648 941 -636
rect 996 -747 997 -647
rect 1101 -648 1102 -636
rect 1178 -747 1179 -647
rect 1255 -648 1256 -636
rect 1388 -747 1389 -647
rect 30 -650 31 -636
rect 422 -747 423 -649
rect 429 -650 430 -636
rect 443 -747 444 -649
rect 446 -650 447 -636
rect 1458 -747 1459 -649
rect 30 -747 31 -651
rect 352 -747 353 -651
rect 408 -652 409 -636
rect 450 -747 451 -651
rect 471 -652 472 -636
rect 772 -747 773 -651
rect 870 -652 871 -636
rect 1031 -747 1032 -651
rect 1059 -652 1060 -636
rect 1101 -747 1102 -651
rect 1150 -652 1151 -636
rect 1255 -747 1256 -651
rect 1262 -652 1263 -636
rect 1395 -747 1396 -651
rect 65 -654 66 -636
rect 93 -654 94 -636
rect 100 -654 101 -636
rect 170 -654 171 -636
rect 191 -654 192 -636
rect 191 -747 192 -653
rect 191 -654 192 -636
rect 191 -747 192 -653
rect 233 -747 234 -653
rect 390 -654 391 -636
rect 415 -654 416 -636
rect 660 -654 661 -636
rect 663 -747 664 -653
rect 1339 -654 1340 -636
rect 1346 -654 1347 -636
rect 1493 -747 1494 -653
rect 65 -747 66 -655
rect 219 -656 220 -636
rect 261 -656 262 -636
rect 282 -747 283 -655
rect 296 -656 297 -636
rect 751 -747 752 -655
rect 870 -747 871 -655
rect 1094 -656 1095 -636
rect 1150 -747 1151 -655
rect 1164 -656 1165 -636
rect 1227 -656 1228 -636
rect 1339 -747 1340 -655
rect 1353 -656 1354 -636
rect 1500 -747 1501 -655
rect 23 -658 24 -636
rect 261 -747 262 -657
rect 296 -747 297 -657
rect 394 -658 395 -636
rect 401 -658 402 -636
rect 1094 -747 1095 -657
rect 1157 -658 1158 -636
rect 1262 -747 1263 -657
rect 1283 -658 1284 -636
rect 1402 -747 1403 -657
rect 23 -747 24 -659
rect 310 -660 311 -636
rect 345 -747 346 -659
rect 464 -660 465 -636
rect 506 -747 507 -659
rect 681 -660 682 -636
rect 688 -660 689 -636
rect 688 -747 689 -659
rect 688 -660 689 -636
rect 688 -747 689 -659
rect 730 -747 731 -659
rect 737 -660 738 -636
rect 744 -660 745 -636
rect 1374 -747 1375 -659
rect 9 -662 10 -636
rect 681 -747 682 -661
rect 702 -662 703 -636
rect 737 -747 738 -661
rect 744 -747 745 -661
rect 1045 -662 1046 -636
rect 1052 -662 1053 -636
rect 1283 -747 1284 -661
rect 1290 -662 1291 -636
rect 1409 -747 1410 -661
rect 79 -664 80 -636
rect 401 -747 402 -663
rect 415 -747 416 -663
rect 621 -747 622 -663
rect 628 -664 629 -636
rect 1115 -664 1116 -636
rect 1171 -664 1172 -636
rect 1290 -747 1291 -663
rect 1304 -664 1305 -636
rect 1416 -747 1417 -663
rect 79 -747 80 -665
rect 121 -666 122 -636
rect 128 -666 129 -636
rect 170 -747 171 -665
rect 219 -747 220 -665
rect 317 -666 318 -636
rect 348 -666 349 -636
rect 408 -747 409 -665
rect 436 -666 437 -636
rect 471 -747 472 -665
rect 509 -666 510 -636
rect 534 -666 535 -636
rect 548 -747 549 -665
rect 583 -666 584 -636
rect 597 -666 598 -636
rect 926 -747 927 -665
rect 940 -747 941 -665
rect 1206 -747 1207 -665
rect 1248 -666 1249 -636
rect 1346 -747 1347 -665
rect 1360 -666 1361 -636
rect 1444 -747 1445 -665
rect 58 -668 59 -636
rect 583 -747 584 -667
rect 614 -747 615 -667
rect 1164 -747 1165 -667
rect 1171 -747 1172 -667
rect 1234 -668 1235 -636
rect 1297 -668 1298 -636
rect 1360 -747 1361 -667
rect 1367 -668 1368 -636
rect 1521 -747 1522 -667
rect 58 -747 59 -669
rect 156 -670 157 -636
rect 268 -747 269 -669
rect 1367 -747 1368 -669
rect 61 -747 62 -671
rect 1297 -747 1298 -671
rect 1311 -672 1312 -636
rect 1423 -747 1424 -671
rect 86 -674 87 -636
rect 429 -747 430 -673
rect 436 -747 437 -673
rect 604 -674 605 -636
rect 628 -747 629 -673
rect 1269 -674 1270 -636
rect 1318 -674 1319 -636
rect 1430 -747 1431 -673
rect 86 -747 87 -675
rect 331 -676 332 -636
rect 359 -676 360 -636
rect 394 -747 395 -675
rect 604 -747 605 -675
rect 695 -676 696 -636
rect 702 -747 703 -675
rect 793 -676 794 -636
rect 842 -676 843 -636
rect 1269 -747 1270 -675
rect 1325 -676 1326 -636
rect 1479 -747 1480 -675
rect 93 -747 94 -677
rect 600 -747 601 -677
rect 635 -678 636 -636
rect 1003 -678 1004 -636
rect 1010 -678 1011 -636
rect 1052 -747 1053 -677
rect 1073 -678 1074 -636
rect 1115 -747 1116 -677
rect 1129 -678 1130 -636
rect 1234 -747 1235 -677
rect 1332 -678 1333 -636
rect 1486 -747 1487 -677
rect 19 -680 20 -636
rect 1073 -747 1074 -679
rect 1080 -680 1081 -636
rect 1129 -747 1130 -679
rect 1143 -680 1144 -636
rect 1248 -747 1249 -679
rect 72 -682 73 -636
rect 1143 -747 1144 -681
rect 1199 -682 1200 -636
rect 1311 -747 1312 -681
rect 72 -747 73 -683
rect 523 -747 524 -683
rect 747 -747 748 -683
rect 1185 -684 1186 -636
rect 1199 -747 1200 -683
rect 1241 -684 1242 -636
rect 96 -686 97 -636
rect 1227 -747 1228 -685
rect 100 -747 101 -687
rect 618 -688 619 -636
rect 761 -747 762 -687
rect 1157 -747 1158 -687
rect 1213 -688 1214 -636
rect 1318 -747 1319 -687
rect 114 -690 115 -636
rect 373 -690 374 -636
rect 380 -690 381 -636
rect 464 -747 465 -689
rect 478 -690 479 -636
rect 1080 -747 1081 -689
rect 1108 -690 1109 -636
rect 1213 -747 1214 -689
rect 1220 -690 1221 -636
rect 1325 -747 1326 -689
rect 114 -747 115 -691
rect 919 -692 920 -636
rect 943 -747 944 -691
rect 1276 -692 1277 -636
rect 121 -747 122 -693
rect 481 -694 482 -636
rect 618 -747 619 -693
rect 1304 -747 1305 -693
rect 128 -747 129 -695
rect 418 -696 419 -636
rect 425 -747 426 -695
rect 695 -747 696 -695
rect 765 -696 766 -636
rect 1353 -747 1354 -695
rect 135 -698 136 -636
rect 173 -698 174 -636
rect 247 -698 248 -636
rect 331 -747 332 -697
rect 359 -747 360 -697
rect 485 -698 486 -636
rect 513 -698 514 -636
rect 765 -747 766 -697
rect 779 -698 780 -636
rect 793 -747 794 -697
rect 856 -698 857 -636
rect 1185 -747 1186 -697
rect 12 -747 13 -699
rect 856 -747 857 -699
rect 877 -700 878 -636
rect 1045 -747 1046 -699
rect 1066 -700 1067 -636
rect 1108 -747 1109 -699
rect 1136 -700 1137 -636
rect 1241 -747 1242 -699
rect 107 -702 108 -636
rect 247 -747 248 -701
rect 310 -747 311 -701
rect 527 -702 528 -636
rect 537 -747 538 -701
rect 779 -747 780 -701
rect 849 -702 850 -636
rect 877 -747 878 -701
rect 919 -747 920 -701
rect 989 -702 990 -636
rect 1017 -702 1018 -636
rect 1059 -747 1060 -701
rect 1087 -702 1088 -636
rect 1276 -747 1277 -701
rect 107 -747 108 -703
rect 240 -704 241 -636
rect 313 -704 314 -636
rect 478 -747 479 -703
rect 485 -747 486 -703
rect 492 -704 493 -636
rect 499 -704 500 -636
rect 527 -747 528 -703
rect 653 -704 654 -636
rect 1220 -747 1221 -703
rect 149 -706 150 -636
rect 156 -747 157 -705
rect 177 -706 178 -636
rect 240 -747 241 -705
rect 317 -747 318 -705
rect 716 -706 717 -636
rect 835 -706 836 -636
rect 989 -747 990 -705
rect 1024 -706 1025 -636
rect 1332 -747 1333 -705
rect 149 -747 150 -707
rect 625 -708 626 -636
rect 639 -708 640 -636
rect 653 -747 654 -707
rect 667 -708 668 -636
rect 1017 -747 1018 -707
rect 1038 -708 1039 -636
rect 1087 -747 1088 -707
rect 103 -747 104 -709
rect 639 -747 640 -709
rect 667 -747 668 -709
rect 709 -710 710 -636
rect 716 -747 717 -709
rect 800 -710 801 -636
rect 814 -710 815 -636
rect 835 -747 836 -709
rect 849 -747 850 -709
rect 891 -710 892 -636
rect 947 -710 948 -636
rect 1003 -747 1004 -709
rect 177 -747 178 -711
rect 184 -712 185 -636
rect 338 -712 339 -636
rect 513 -747 514 -711
rect 565 -747 566 -711
rect 1038 -747 1039 -711
rect 184 -747 185 -713
rect 212 -714 213 -636
rect 338 -747 339 -713
rect 674 -714 675 -636
rect 709 -747 710 -713
rect 723 -714 724 -636
rect 786 -714 787 -636
rect 800 -747 801 -713
rect 814 -747 815 -713
rect 821 -714 822 -636
rect 954 -714 955 -636
rect 1010 -747 1011 -713
rect 163 -716 164 -636
rect 212 -747 213 -715
rect 355 -716 356 -636
rect 947 -747 948 -715
rect 961 -716 962 -636
rect 1066 -747 1067 -715
rect 142 -718 143 -636
rect 163 -747 164 -717
rect 355 -747 356 -717
rect 457 -718 458 -636
rect 492 -747 493 -717
rect 660 -747 661 -717
rect 786 -747 787 -717
rect 1122 -718 1123 -636
rect 142 -747 143 -719
rect 271 -720 272 -636
rect 366 -720 367 -636
rect 723 -747 724 -719
rect 758 -720 759 -636
rect 1122 -747 1123 -719
rect 75 -722 76 -636
rect 271 -747 272 -721
rect 373 -747 374 -721
rect 520 -722 521 -636
rect 632 -722 633 -636
rect 891 -747 892 -721
rect 898 -722 899 -636
rect 954 -747 955 -721
rect 964 -722 965 -636
rect 1465 -747 1466 -721
rect 289 -724 290 -636
rect 632 -747 633 -723
rect 646 -724 647 -636
rect 674 -747 675 -723
rect 758 -747 759 -723
rect 1192 -724 1193 -636
rect 226 -726 227 -636
rect 289 -747 290 -725
rect 457 -747 458 -725
rect 576 -726 577 -636
rect 590 -726 591 -636
rect 646 -747 647 -725
rect 821 -747 822 -725
rect 887 -747 888 -725
rect 905 -726 906 -636
rect 961 -747 962 -725
rect 968 -726 969 -636
rect 1024 -747 1025 -725
rect 226 -747 227 -727
rect 254 -728 255 -636
rect 499 -747 500 -727
rect 541 -747 542 -727
rect 555 -728 556 -636
rect 590 -747 591 -727
rect 611 -728 612 -636
rect 1192 -747 1193 -727
rect 205 -730 206 -636
rect 254 -747 255 -729
rect 534 -747 535 -729
rect 555 -747 556 -729
rect 569 -730 570 -636
rect 576 -747 577 -729
rect 611 -747 612 -729
rect 1136 -747 1137 -729
rect 205 -747 206 -731
rect 275 -732 276 -636
rect 562 -732 563 -636
rect 569 -747 570 -731
rect 863 -732 864 -636
rect 898 -747 899 -731
rect 905 -747 906 -731
rect 975 -732 976 -636
rect 982 -732 983 -636
rect 1507 -747 1508 -731
rect 117 -734 118 -636
rect 982 -747 983 -733
rect 275 -747 276 -735
rect 303 -736 304 -636
rect 366 -747 367 -735
rect 975 -747 976 -735
rect 198 -738 199 -636
rect 303 -747 304 -737
rect 380 -747 381 -737
rect 562 -747 563 -737
rect 863 -747 864 -737
rect 933 -738 934 -636
rect 51 -740 52 -636
rect 198 -747 199 -739
rect 828 -740 829 -636
rect 933 -747 934 -739
rect 51 -747 52 -741
rect 75 -747 76 -741
rect 117 -747 118 -741
rect 828 -747 829 -741
rect 912 -742 913 -636
rect 968 -747 969 -741
rect 884 -744 885 -636
rect 912 -747 913 -743
rect 842 -747 843 -745
rect 884 -747 885 -745
rect 2 -757 3 -755
rect 1094 -757 1095 -755
rect 2 -888 3 -758
rect 611 -759 612 -755
rect 614 -759 615 -755
rect 1437 -759 1438 -755
rect 9 -761 10 -755
rect 338 -761 339 -755
rect 369 -761 370 -755
rect 943 -761 944 -755
rect 1066 -761 1067 -755
rect 1094 -888 1095 -760
rect 1437 -888 1438 -760
rect 1458 -761 1459 -755
rect 9 -888 10 -762
rect 642 -888 643 -762
rect 649 -888 650 -762
rect 1297 -763 1298 -755
rect 1458 -888 1459 -762
rect 1472 -763 1473 -755
rect 12 -765 13 -755
rect 968 -765 969 -755
rect 1066 -888 1067 -764
rect 1213 -765 1214 -755
rect 1472 -888 1473 -764
rect 1493 -765 1494 -755
rect 23 -767 24 -755
rect 271 -767 272 -755
rect 310 -767 311 -755
rect 712 -888 713 -766
rect 747 -767 748 -755
rect 1213 -888 1214 -766
rect 16 -769 17 -755
rect 23 -888 24 -768
rect 47 -888 48 -768
rect 632 -769 633 -755
rect 653 -769 654 -755
rect 663 -769 664 -755
rect 775 -769 776 -755
rect 1521 -769 1522 -755
rect 16 -888 17 -770
rect 184 -771 185 -755
rect 226 -771 227 -755
rect 366 -771 367 -755
rect 394 -771 395 -755
rect 397 -849 398 -770
rect 443 -771 444 -755
rect 443 -888 444 -770
rect 443 -771 444 -755
rect 443 -888 444 -770
rect 471 -771 472 -755
rect 471 -888 472 -770
rect 471 -771 472 -755
rect 471 -888 472 -770
rect 478 -771 479 -755
rect 478 -888 479 -770
rect 478 -771 479 -755
rect 478 -888 479 -770
rect 485 -771 486 -755
rect 488 -849 489 -770
rect 499 -771 500 -755
rect 499 -888 500 -770
rect 499 -771 500 -755
rect 499 -888 500 -770
rect 509 -888 510 -770
rect 1045 -771 1046 -755
rect 1164 -771 1165 -755
rect 1297 -888 1298 -770
rect 58 -773 59 -755
rect 1507 -773 1508 -755
rect 58 -888 59 -774
rect 79 -775 80 -755
rect 117 -775 118 -755
rect 723 -775 724 -755
rect 884 -775 885 -755
rect 1248 -775 1249 -755
rect 51 -777 52 -755
rect 79 -888 80 -776
rect 121 -777 122 -755
rect 310 -888 311 -776
rect 324 -777 325 -755
rect 422 -777 423 -755
rect 485 -888 486 -776
rect 527 -777 528 -755
rect 534 -777 535 -755
rect 1332 -777 1333 -755
rect 51 -888 52 -778
rect 296 -779 297 -755
rect 324 -888 325 -778
rect 439 -888 440 -778
rect 520 -779 521 -755
rect 530 -779 531 -755
rect 537 -779 538 -755
rect 751 -779 752 -755
rect 887 -779 888 -755
rect 1444 -779 1445 -755
rect 61 -781 62 -755
rect 1073 -781 1074 -755
rect 1164 -888 1165 -780
rect 1325 -781 1326 -755
rect 1332 -888 1333 -780
rect 1346 -781 1347 -755
rect 1444 -888 1445 -780
rect 1486 -781 1487 -755
rect 65 -783 66 -755
rect 460 -888 461 -782
rect 520 -888 521 -782
rect 604 -783 605 -755
rect 611 -888 612 -782
rect 898 -783 899 -755
rect 940 -783 941 -755
rect 1423 -783 1424 -755
rect 65 -888 66 -784
rect 317 -785 318 -755
rect 338 -888 339 -784
rect 352 -785 353 -755
rect 394 -888 395 -784
rect 401 -785 402 -755
rect 422 -888 423 -784
rect 576 -785 577 -755
rect 583 -785 584 -755
rect 604 -888 605 -784
rect 618 -785 619 -755
rect 702 -785 703 -755
rect 723 -888 724 -784
rect 800 -785 801 -755
rect 856 -785 857 -755
rect 898 -888 899 -784
rect 943 -888 944 -784
rect 1255 -785 1256 -755
rect 72 -787 73 -755
rect 1360 -787 1361 -755
rect 72 -888 73 -788
rect 261 -789 262 -755
rect 296 -888 297 -788
rect 768 -888 769 -788
rect 800 -888 801 -788
rect 821 -789 822 -755
rect 856 -888 857 -788
rect 947 -789 948 -755
rect 968 -888 969 -788
rect 1101 -789 1102 -755
rect 1150 -789 1151 -755
rect 1255 -888 1256 -788
rect 1360 -888 1361 -788
rect 1409 -789 1410 -755
rect 75 -791 76 -755
rect 1185 -791 1186 -755
rect 1199 -791 1200 -755
rect 1346 -888 1347 -790
rect 1409 -888 1410 -790
rect 1430 -791 1431 -755
rect 100 -793 101 -755
rect 1423 -888 1424 -792
rect 1430 -888 1431 -792
rect 1451 -793 1452 -755
rect 100 -888 101 -794
rect 359 -795 360 -755
rect 401 -888 402 -794
rect 408 -795 409 -755
rect 464 -795 465 -755
rect 576 -888 577 -794
rect 597 -795 598 -755
rect 961 -795 962 -755
rect 1017 -795 1018 -755
rect 1073 -888 1074 -794
rect 1101 -888 1102 -794
rect 1129 -795 1130 -755
rect 1199 -888 1200 -794
rect 1234 -795 1235 -755
rect 1248 -888 1249 -794
rect 1283 -795 1284 -755
rect 1451 -888 1452 -794
rect 1465 -795 1466 -755
rect 114 -797 115 -755
rect 1325 -888 1326 -796
rect 1465 -888 1466 -796
rect 1479 -797 1480 -755
rect 114 -888 115 -798
rect 282 -799 283 -755
rect 408 -888 409 -798
rect 464 -888 465 -798
rect 1122 -799 1123 -755
rect 1129 -888 1130 -798
rect 1192 -799 1193 -755
rect 1234 -888 1235 -798
rect 1269 -799 1270 -755
rect 1283 -888 1284 -798
rect 1311 -799 1312 -755
rect 1479 -888 1480 -798
rect 1500 -799 1501 -755
rect 121 -888 122 -800
rect 177 -801 178 -755
rect 184 -888 185 -800
rect 303 -801 304 -755
rect 425 -801 426 -755
rect 1122 -888 1123 -800
rect 1171 -801 1172 -755
rect 1311 -888 1312 -800
rect 1500 -888 1501 -800
rect 1514 -801 1515 -755
rect 131 -888 132 -802
rect 170 -803 171 -755
rect 177 -888 178 -802
rect 212 -803 213 -755
rect 226 -888 227 -802
rect 380 -803 381 -755
rect 523 -803 524 -755
rect 989 -803 990 -755
rect 1017 -888 1018 -802
rect 1262 -803 1263 -755
rect 1269 -888 1270 -802
rect 1304 -803 1305 -755
rect 1514 -888 1515 -802
rect 1528 -803 1529 -755
rect 107 -805 108 -755
rect 170 -888 171 -804
rect 205 -805 206 -755
rect 317 -888 318 -804
rect 380 -888 381 -804
rect 555 -805 556 -755
rect 569 -805 570 -755
rect 884 -888 885 -804
rect 891 -805 892 -755
rect 1150 -888 1151 -804
rect 1192 -888 1193 -804
rect 1227 -805 1228 -755
rect 107 -888 108 -806
rect 219 -807 220 -755
rect 236 -888 237 -806
rect 282 -888 283 -806
rect 289 -807 290 -755
rect 303 -888 304 -806
rect 436 -807 437 -755
rect 555 -888 556 -806
rect 618 -888 619 -806
rect 926 -807 927 -755
rect 989 -888 990 -806
rect 1052 -807 1053 -755
rect 1115 -807 1116 -755
rect 1171 -888 1172 -806
rect 1227 -888 1228 -806
rect 1290 -807 1291 -755
rect 30 -809 31 -755
rect 1052 -888 1053 -808
rect 30 -888 31 -810
rect 450 -811 451 -755
rect 467 -888 468 -810
rect 1290 -888 1291 -810
rect 135 -813 136 -755
rect 691 -888 692 -812
rect 695 -813 696 -755
rect 702 -888 703 -812
rect 779 -813 780 -755
rect 1304 -888 1305 -812
rect 135 -888 136 -814
rect 163 -815 164 -755
rect 205 -888 206 -814
rect 1503 -888 1504 -814
rect 138 -817 139 -755
rect 772 -817 773 -755
rect 779 -888 780 -816
rect 793 -817 794 -755
rect 814 -817 815 -755
rect 821 -888 822 -816
rect 905 -817 906 -755
rect 926 -888 927 -816
rect 1038 -817 1039 -755
rect 1486 -888 1487 -816
rect 93 -819 94 -755
rect 814 -888 815 -818
rect 905 -888 906 -818
rect 954 -819 955 -755
rect 1038 -888 1039 -818
rect 1080 -819 1081 -755
rect 93 -888 94 -820
rect 506 -821 507 -755
rect 534 -888 535 -820
rect 597 -888 598 -820
rect 632 -888 633 -820
rect 674 -821 675 -755
rect 681 -821 682 -755
rect 695 -888 696 -820
rect 730 -821 731 -755
rect 772 -888 773 -820
rect 786 -821 787 -755
rect 1185 -888 1186 -820
rect 142 -823 143 -755
rect 359 -888 360 -822
rect 429 -823 430 -755
rect 674 -888 675 -822
rect 688 -823 689 -755
rect 730 -888 731 -822
rect 758 -823 759 -755
rect 954 -888 955 -822
rect 1045 -888 1046 -822
rect 1087 -823 1088 -755
rect 86 -825 87 -755
rect 429 -888 430 -824
rect 436 -888 437 -824
rect 891 -888 892 -824
rect 919 -825 920 -755
rect 961 -888 962 -824
rect 1080 -888 1081 -824
rect 1136 -825 1137 -755
rect 86 -888 87 -826
rect 709 -827 710 -755
rect 758 -888 759 -826
rect 807 -827 808 -755
rect 919 -888 920 -826
rect 996 -827 997 -755
rect 1087 -888 1088 -826
rect 1206 -827 1207 -755
rect 103 -829 104 -755
rect 142 -888 143 -828
rect 163 -888 164 -828
rect 1493 -888 1494 -828
rect 212 -888 213 -830
rect 366 -888 367 -830
rect 450 -888 451 -830
rect 716 -831 717 -755
rect 793 -888 794 -830
rect 835 -831 836 -755
rect 947 -888 948 -830
rect 996 -888 997 -830
rect 1136 -888 1137 -830
rect 1178 -831 1179 -755
rect 1206 -888 1207 -830
rect 1241 -831 1242 -755
rect 219 -888 220 -832
rect 268 -833 269 -755
rect 492 -833 493 -755
rect 681 -888 682 -832
rect 709 -888 710 -832
rect 1024 -833 1025 -755
rect 1241 -888 1242 -832
rect 1276 -833 1277 -755
rect 240 -835 241 -755
rect 289 -888 290 -834
rect 331 -835 332 -755
rect 492 -888 493 -834
rect 506 -888 507 -834
rect 744 -835 745 -755
rect 1024 -888 1025 -834
rect 1108 -835 1109 -755
rect 1276 -888 1277 -834
rect 1339 -835 1340 -755
rect 233 -837 234 -755
rect 240 -888 241 -836
rect 254 -837 255 -755
rect 352 -888 353 -836
rect 541 -837 542 -755
rect 1031 -837 1032 -755
rect 1108 -888 1109 -836
rect 1143 -837 1144 -755
rect 191 -839 192 -755
rect 233 -888 234 -838
rect 261 -888 262 -838
rect 663 -888 664 -838
rect 667 -839 668 -755
rect 751 -888 752 -838
rect 912 -839 913 -755
rect 1031 -888 1032 -838
rect 1143 -888 1144 -838
rect 1318 -839 1319 -755
rect 191 -888 192 -840
rect 275 -841 276 -755
rect 331 -888 332 -840
rect 373 -841 374 -755
rect 541 -888 542 -840
rect 807 -888 808 -840
rect 863 -841 864 -755
rect 912 -888 913 -840
rect 999 -888 1000 -840
rect 1339 -888 1340 -840
rect 128 -843 129 -755
rect 275 -888 276 -842
rect 373 -888 374 -842
rect 513 -843 514 -755
rect 544 -843 545 -755
rect 765 -843 766 -755
rect 1157 -843 1158 -755
rect 1318 -888 1319 -842
rect 37 -845 38 -755
rect 513 -888 514 -844
rect 548 -845 549 -755
rect 583 -888 584 -844
rect 600 -845 601 -755
rect 786 -888 787 -844
rect 838 -888 839 -844
rect 1157 -888 1158 -844
rect 128 -888 129 -846
rect 1353 -847 1354 -755
rect 198 -849 199 -755
rect 254 -888 255 -848
rect 268 -888 269 -848
rect 345 -849 346 -755
rect 530 -888 531 -848
rect 548 -888 549 -848
rect 551 -888 552 -848
rect 982 -849 983 -755
rect 1353 -888 1354 -848
rect 1367 -849 1368 -755
rect 198 -888 199 -850
rect 247 -851 248 -755
rect 345 -888 346 -850
rect 355 -851 356 -755
rect 562 -851 563 -755
rect 1178 -888 1179 -850
rect 1367 -888 1368 -850
rect 1374 -851 1375 -755
rect 44 -853 45 -755
rect 247 -888 248 -852
rect 562 -888 563 -852
rect 590 -853 591 -755
rect 639 -853 640 -755
rect 982 -888 983 -852
rect 1374 -888 1375 -852
rect 1381 -853 1382 -755
rect 44 -888 45 -854
rect 716 -888 717 -854
rect 737 -855 738 -755
rect 744 -888 745 -854
rect 765 -888 766 -854
rect 933 -855 934 -755
rect 1381 -888 1382 -854
rect 1388 -855 1389 -755
rect 166 -888 167 -856
rect 590 -888 591 -856
rect 646 -857 647 -755
rect 667 -888 668 -856
rect 737 -888 738 -856
rect 877 -857 878 -755
rect 933 -888 934 -856
rect 1003 -857 1004 -755
rect 1388 -888 1389 -856
rect 1395 -857 1396 -755
rect 457 -859 458 -755
rect 877 -888 878 -858
rect 1395 -888 1396 -858
rect 1402 -859 1403 -755
rect 457 -888 458 -860
rect 1220 -861 1221 -755
rect 1402 -888 1403 -860
rect 1416 -861 1417 -755
rect 569 -888 570 -862
rect 835 -888 836 -862
rect 625 -865 626 -755
rect 1003 -888 1004 -864
rect 40 -888 41 -866
rect 625 -888 626 -866
rect 646 -888 647 -866
rect 1262 -888 1263 -866
rect 653 -888 654 -868
rect 1115 -888 1116 -868
rect 656 -888 657 -870
rect 870 -871 871 -755
rect 660 -873 661 -755
rect 863 -888 864 -872
rect 870 -888 871 -872
rect 975 -873 976 -755
rect 149 -875 150 -755
rect 660 -888 661 -874
rect 761 -875 762 -755
rect 1220 -888 1221 -874
rect 149 -888 150 -876
rect 156 -877 157 -755
rect 828 -877 829 -755
rect 1416 -888 1417 -876
rect 156 -888 157 -878
rect 387 -879 388 -755
rect 639 -888 640 -878
rect 828 -888 829 -878
rect 975 -888 976 -878
rect 1010 -879 1011 -755
rect 369 -888 370 -880
rect 387 -888 388 -880
rect 1010 -888 1011 -880
rect 1059 -881 1060 -755
rect 842 -883 843 -755
rect 1059 -888 1060 -882
rect 842 -888 843 -884
rect 849 -885 850 -755
rect 537 -888 538 -886
rect 849 -888 850 -886
rect 23 -898 24 -896
rect 23 -1005 24 -897
rect 23 -898 24 -896
rect 23 -1005 24 -897
rect 40 -898 41 -896
rect 359 -898 360 -896
rect 376 -1005 377 -897
rect 1178 -898 1179 -896
rect 1318 -898 1319 -896
rect 1426 -1005 1427 -897
rect 1503 -898 1504 -896
rect 1514 -898 1515 -896
rect 44 -900 45 -896
rect 1101 -900 1102 -896
rect 1178 -1005 1179 -899
rect 1234 -900 1235 -896
rect 1402 -900 1403 -896
rect 1402 -1005 1403 -899
rect 1402 -900 1403 -896
rect 1402 -1005 1403 -899
rect 51 -902 52 -896
rect 464 -902 465 -896
rect 467 -902 468 -896
rect 1073 -902 1074 -896
rect 1234 -1005 1235 -901
rect 1255 -902 1256 -896
rect 51 -1005 52 -903
rect 296 -904 297 -896
rect 334 -1005 335 -903
rect 338 -904 339 -896
rect 352 -904 353 -896
rect 359 -1005 360 -903
rect 387 -904 388 -896
rect 551 -904 552 -896
rect 604 -904 605 -896
rect 604 -1005 605 -903
rect 604 -904 605 -896
rect 604 -1005 605 -903
rect 646 -904 647 -896
rect 1038 -904 1039 -896
rect 1066 -904 1067 -896
rect 1069 -904 1070 -896
rect 1073 -1005 1074 -903
rect 1500 -904 1501 -896
rect 30 -906 31 -896
rect 387 -1005 388 -905
rect 429 -906 430 -896
rect 436 -906 437 -896
rect 443 -906 444 -896
rect 464 -1005 465 -905
rect 471 -906 472 -896
rect 471 -1005 472 -905
rect 471 -906 472 -896
rect 471 -1005 472 -905
rect 485 -906 486 -896
rect 485 -1005 486 -905
rect 485 -906 486 -896
rect 485 -1005 486 -905
rect 492 -906 493 -896
rect 649 -906 650 -896
rect 656 -906 657 -896
rect 730 -906 731 -896
rect 747 -1005 748 -905
rect 758 -906 759 -896
rect 761 -1005 762 -905
rect 1297 -906 1298 -896
rect 30 -1005 31 -907
rect 170 -908 171 -896
rect 184 -908 185 -896
rect 243 -1005 244 -907
rect 296 -1005 297 -907
rect 1052 -908 1053 -896
rect 1066 -1005 1067 -907
rect 1108 -908 1109 -896
rect 1297 -1005 1298 -907
rect 1374 -908 1375 -896
rect 16 -910 17 -896
rect 170 -1005 171 -909
rect 184 -1005 185 -909
rect 191 -910 192 -896
rect 198 -910 199 -896
rect 369 -910 370 -896
rect 436 -1005 437 -909
rect 527 -910 528 -896
rect 534 -910 535 -896
rect 562 -910 563 -896
rect 660 -910 661 -896
rect 1045 -910 1046 -896
rect 1094 -910 1095 -896
rect 1255 -1005 1256 -909
rect 1374 -1005 1375 -909
rect 1437 -910 1438 -896
rect 58 -912 59 -896
rect 58 -1005 59 -911
rect 58 -912 59 -896
rect 58 -1005 59 -911
rect 65 -912 66 -896
rect 642 -912 643 -896
rect 681 -912 682 -896
rect 681 -1005 682 -911
rect 681 -912 682 -896
rect 681 -1005 682 -911
rect 691 -912 692 -896
rect 1010 -912 1011 -896
rect 1017 -912 1018 -896
rect 1318 -1005 1319 -911
rect 1437 -1005 1438 -911
rect 1493 -912 1494 -896
rect 65 -1005 66 -913
rect 79 -914 80 -896
rect 100 -914 101 -896
rect 492 -1005 493 -913
rect 495 -1005 496 -913
rect 646 -1005 647 -913
rect 705 -1005 706 -913
rect 1164 -914 1165 -896
rect 79 -1005 80 -915
rect 93 -916 94 -896
rect 100 -1005 101 -915
rect 205 -916 206 -896
rect 212 -916 213 -896
rect 429 -1005 430 -915
rect 450 -916 451 -896
rect 600 -1005 601 -915
rect 639 -916 640 -896
rect 1094 -1005 1095 -915
rect 16 -1005 17 -917
rect 93 -1005 94 -917
rect 114 -918 115 -896
rect 233 -918 234 -896
rect 240 -918 241 -896
rect 443 -1005 444 -917
rect 499 -918 500 -896
rect 499 -1005 500 -917
rect 499 -918 500 -896
rect 499 -1005 500 -917
rect 509 -918 510 -896
rect 674 -918 675 -896
rect 709 -918 710 -896
rect 1409 -918 1410 -896
rect 9 -920 10 -896
rect 674 -1005 675 -919
rect 712 -920 713 -896
rect 1304 -920 1305 -896
rect 9 -1005 10 -921
rect 72 -922 73 -896
rect 96 -1005 97 -921
rect 233 -1005 234 -921
rect 338 -1005 339 -921
rect 618 -922 619 -896
rect 639 -1005 640 -921
rect 992 -1005 993 -921
rect 1024 -922 1025 -896
rect 1024 -1005 1025 -921
rect 1024 -922 1025 -896
rect 1024 -1005 1025 -921
rect 1045 -1005 1046 -921
rect 1122 -922 1123 -896
rect 1143 -922 1144 -896
rect 1409 -1005 1410 -921
rect 72 -1005 73 -923
rect 142 -924 143 -896
rect 145 -1005 146 -923
rect 1052 -1005 1053 -923
rect 1122 -1005 1123 -923
rect 1136 -924 1137 -896
rect 1143 -1005 1144 -923
rect 1199 -924 1200 -896
rect 1290 -924 1291 -896
rect 1304 -1005 1305 -923
rect 114 -1005 115 -925
rect 310 -926 311 -896
rect 352 -1005 353 -925
rect 460 -926 461 -896
rect 513 -926 514 -896
rect 527 -1005 528 -925
rect 534 -1005 535 -925
rect 618 -1005 619 -925
rect 667 -926 668 -896
rect 709 -1005 710 -925
rect 730 -1005 731 -925
rect 800 -926 801 -896
rect 807 -926 808 -896
rect 1360 -926 1361 -896
rect 142 -1005 143 -927
rect 1430 -928 1431 -896
rect 163 -930 164 -896
rect 226 -930 227 -896
rect 310 -1005 311 -929
rect 415 -930 416 -896
rect 513 -1005 514 -929
rect 632 -930 633 -896
rect 754 -1005 755 -929
rect 1227 -930 1228 -896
rect 1290 -1005 1291 -929
rect 1353 -930 1354 -896
rect 1360 -1005 1361 -929
rect 1423 -930 1424 -896
rect 37 -932 38 -896
rect 1227 -1005 1228 -931
rect 1353 -1005 1354 -931
rect 1416 -932 1417 -896
rect 37 -1005 38 -933
rect 156 -934 157 -896
rect 163 -1005 164 -933
rect 478 -934 479 -896
rect 520 -934 521 -896
rect 667 -1005 668 -933
rect 758 -1005 759 -933
rect 1276 -934 1277 -896
rect 1416 -1005 1417 -933
rect 1465 -934 1466 -896
rect 2 -936 3 -896
rect 520 -1005 521 -935
rect 537 -936 538 -896
rect 1325 -936 1326 -896
rect 2 -1005 3 -937
rect 695 -938 696 -896
rect 768 -938 769 -896
rect 1444 -938 1445 -896
rect 131 -940 132 -896
rect 695 -1005 696 -939
rect 800 -1005 801 -939
rect 891 -940 892 -896
rect 898 -940 899 -896
rect 898 -1005 899 -939
rect 898 -940 899 -896
rect 898 -1005 899 -939
rect 908 -1005 909 -939
rect 1332 -940 1333 -896
rect 1444 -1005 1445 -939
rect 1472 -940 1473 -896
rect 156 -1005 157 -941
rect 653 -942 654 -896
rect 807 -1005 808 -941
rect 856 -942 857 -896
rect 891 -1005 892 -941
rect 905 -942 906 -896
rect 919 -942 920 -896
rect 919 -1005 920 -941
rect 919 -942 920 -896
rect 919 -1005 920 -941
rect 940 -1005 941 -941
rect 954 -942 955 -896
rect 975 -942 976 -896
rect 978 -972 979 -941
rect 989 -942 990 -896
rect 1038 -1005 1039 -941
rect 1129 -942 1130 -896
rect 1136 -1005 1137 -941
rect 1199 -1005 1200 -941
rect 1248 -942 1249 -896
rect 1325 -1005 1326 -941
rect 1381 -942 1382 -896
rect 177 -944 178 -896
rect 226 -1005 227 -943
rect 380 -944 381 -896
rect 450 -1005 451 -943
rect 478 -1005 479 -943
rect 877 -944 878 -896
rect 943 -944 944 -896
rect 1164 -1005 1165 -943
rect 1248 -1005 1249 -943
rect 1283 -944 1284 -896
rect 1332 -1005 1333 -943
rect 1388 -944 1389 -896
rect 128 -946 129 -896
rect 177 -1005 178 -945
rect 191 -1005 192 -945
rect 261 -946 262 -896
rect 275 -946 276 -896
rect 380 -1005 381 -945
rect 415 -1005 416 -945
rect 1185 -946 1186 -896
rect 1283 -1005 1284 -945
rect 1346 -946 1347 -896
rect 1381 -1005 1382 -945
rect 1451 -946 1452 -896
rect 121 -948 122 -896
rect 128 -1005 129 -947
rect 198 -1005 199 -947
rect 236 -948 237 -896
rect 254 -948 255 -896
rect 275 -1005 276 -947
rect 373 -948 374 -896
rect 1451 -1005 1452 -947
rect 121 -1005 122 -949
rect 149 -950 150 -896
rect 205 -1005 206 -949
rect 373 -1005 374 -949
rect 537 -1005 538 -949
rect 1171 -950 1172 -896
rect 1185 -1005 1186 -949
rect 1241 -950 1242 -896
rect 1388 -1005 1389 -949
rect 1458 -950 1459 -896
rect 149 -1005 150 -951
rect 810 -952 811 -896
rect 824 -1005 825 -951
rect 926 -952 927 -896
rect 975 -1005 976 -951
rect 1010 -1005 1011 -951
rect 1423 -1005 1424 -951
rect 212 -1005 213 -953
rect 303 -954 304 -896
rect 541 -954 542 -896
rect 1220 -954 1221 -896
rect 1241 -1005 1242 -953
rect 1269 -954 1270 -896
rect 254 -1005 255 -955
rect 324 -956 325 -896
rect 541 -1005 542 -955
rect 562 -1005 563 -955
rect 576 -956 577 -896
rect 660 -1005 661 -955
rect 677 -1005 678 -955
rect 1220 -1005 1221 -955
rect 1269 -1005 1270 -955
rect 1311 -956 1312 -896
rect 261 -1005 262 -957
rect 289 -958 290 -896
rect 303 -1005 304 -957
rect 394 -958 395 -896
rect 544 -958 545 -896
rect 590 -958 591 -896
rect 828 -958 829 -896
rect 905 -1005 906 -957
rect 926 -1005 927 -957
rect 933 -958 934 -896
rect 1059 -958 1060 -896
rect 1458 -1005 1459 -957
rect 44 -1005 45 -959
rect 544 -1005 545 -959
rect 548 -960 549 -896
rect 1430 -1005 1431 -959
rect 289 -1005 290 -961
rect 408 -962 409 -896
rect 551 -1005 552 -961
rect 1346 -1005 1347 -961
rect 324 -1005 325 -963
rect 345 -964 346 -896
rect 394 -1005 395 -963
rect 751 -964 752 -896
rect 828 -1005 829 -963
rect 1276 -1005 1277 -963
rect 1311 -1005 1312 -963
rect 1339 -964 1340 -896
rect 247 -966 248 -896
rect 345 -1005 346 -965
rect 401 -966 402 -896
rect 408 -1005 409 -965
rect 555 -966 556 -896
rect 576 -1005 577 -965
rect 590 -1005 591 -965
rect 597 -966 598 -896
rect 831 -1005 832 -965
rect 1031 -966 1032 -896
rect 1059 -1005 1060 -965
rect 1080 -966 1081 -896
rect 1129 -1005 1130 -965
rect 1192 -966 1193 -896
rect 1339 -1005 1340 -965
rect 1395 -966 1396 -896
rect 86 -968 87 -896
rect 555 -1005 556 -967
rect 597 -1005 598 -967
rect 737 -968 738 -896
rect 838 -968 839 -896
rect 1479 -968 1480 -896
rect 86 -1005 87 -969
rect 107 -970 108 -896
rect 219 -970 220 -896
rect 401 -1005 402 -969
rect 723 -970 724 -896
rect 737 -1005 738 -969
rect 849 -970 850 -896
rect 859 -1005 860 -969
rect 877 -1005 878 -969
rect 884 -970 885 -896
rect 933 -1005 934 -969
rect 947 -970 948 -896
rect 996 -970 997 -896
rect 1395 -1005 1396 -969
rect 107 -1005 108 -971
rect 135 -972 136 -896
rect 219 -1005 220 -971
rect 506 -972 507 -896
rect 625 -972 626 -896
rect 849 -1005 850 -971
rect 856 -1005 857 -971
rect 954 -1005 955 -971
rect 968 -972 969 -896
rect 996 -1005 997 -971
rect 1003 -972 1004 -896
rect 1031 -1005 1032 -971
rect 1069 -1005 1070 -971
rect 1108 -1005 1109 -971
rect 1171 -1005 1172 -971
rect 1213 -972 1214 -896
rect 135 -1005 136 -973
rect 457 -974 458 -896
rect 583 -974 584 -896
rect 625 -1005 626 -973
rect 884 -1005 885 -973
rect 912 -974 913 -896
rect 947 -1005 948 -973
rect 961 -974 962 -896
rect 1003 -1005 1004 -973
rect 1115 -974 1116 -896
rect 1192 -1005 1193 -973
rect 1367 -974 1368 -896
rect 247 -1005 248 -975
rect 299 -1005 300 -975
rect 331 -976 332 -896
rect 457 -1005 458 -975
rect 611 -976 612 -896
rect 968 -1005 969 -975
rect 1080 -1005 1081 -975
rect 1150 -976 1151 -896
rect 1213 -1005 1214 -975
rect 1262 -976 1263 -896
rect 1367 -1005 1368 -975
rect 1486 -976 1487 -896
rect 282 -978 283 -896
rect 506 -1005 507 -977
rect 611 -1005 612 -977
rect 702 -978 703 -896
rect 716 -978 717 -896
rect 1262 -1005 1263 -977
rect 282 -1005 283 -979
rect 569 -980 570 -896
rect 632 -1005 633 -979
rect 702 -1005 703 -979
rect 863 -980 864 -896
rect 961 -1005 962 -979
rect 1087 -980 1088 -896
rect 1115 -1005 1116 -979
rect 1150 -1005 1151 -979
rect 1206 -980 1207 -896
rect 366 -982 367 -896
rect 723 -1005 724 -981
rect 835 -982 836 -896
rect 1206 -1005 1207 -981
rect 268 -984 269 -896
rect 366 -1005 367 -983
rect 422 -984 423 -896
rect 583 -1005 584 -983
rect 688 -984 689 -896
rect 912 -1005 913 -983
rect 1087 -1005 1088 -983
rect 1157 -984 1158 -896
rect 268 -1005 269 -985
rect 317 -986 318 -896
rect 422 -1005 423 -985
rect 744 -986 745 -896
rect 751 -1005 752 -985
rect 1157 -1005 1158 -985
rect 317 -1005 318 -987
rect 688 -1005 689 -987
rect 691 -1005 692 -987
rect 716 -1005 717 -987
rect 744 -1005 745 -987
rect 1101 -1005 1102 -987
rect 569 -1005 570 -989
rect 765 -990 766 -896
rect 786 -990 787 -896
rect 835 -1005 836 -989
rect 863 -1005 864 -989
rect 870 -990 871 -896
rect 653 -1005 654 -991
rect 870 -1005 871 -991
rect 765 -1005 766 -993
rect 772 -994 773 -896
rect 786 -1005 787 -993
rect 814 -994 815 -896
rect 548 -1005 549 -995
rect 772 -1005 773 -995
rect 793 -996 794 -896
rect 814 -1005 815 -995
rect 779 -998 780 -896
rect 793 -1005 794 -997
rect 779 -1005 780 -999
rect 842 -1000 843 -896
rect 821 -1002 822 -896
rect 842 -1005 843 -1001
rect 821 -1005 822 -1003
rect 1017 -1005 1018 -1003
rect 72 -1015 73 -1013
rect 758 -1015 759 -1013
rect 796 -1152 797 -1014
rect 1038 -1015 1039 -1013
rect 1150 -1015 1151 -1013
rect 1150 -1152 1151 -1014
rect 1150 -1015 1151 -1013
rect 1150 -1152 1151 -1014
rect 1164 -1015 1165 -1013
rect 1591 -1152 1592 -1014
rect 72 -1152 73 -1016
rect 82 -1152 83 -1016
rect 93 -1017 94 -1013
rect 968 -1017 969 -1013
rect 989 -1017 990 -1013
rect 1234 -1017 1235 -1013
rect 1276 -1017 1277 -1013
rect 1570 -1152 1571 -1016
rect 93 -1152 94 -1018
rect 219 -1019 220 -1013
rect 226 -1019 227 -1013
rect 299 -1019 300 -1013
rect 310 -1019 311 -1013
rect 537 -1019 538 -1013
rect 541 -1019 542 -1013
rect 1311 -1019 1312 -1013
rect 1325 -1019 1326 -1013
rect 1486 -1152 1487 -1018
rect 2 -1021 3 -1013
rect 541 -1152 542 -1020
rect 548 -1021 549 -1013
rect 793 -1021 794 -1013
rect 821 -1021 822 -1013
rect 1409 -1021 1410 -1013
rect 1423 -1021 1424 -1013
rect 1444 -1021 1445 -1013
rect 1451 -1021 1452 -1013
rect 1535 -1152 1536 -1020
rect 2 -1152 3 -1022
rect 268 -1023 269 -1013
rect 310 -1152 311 -1022
rect 894 -1152 895 -1022
rect 908 -1023 909 -1013
rect 1514 -1152 1515 -1022
rect 44 -1025 45 -1013
rect 226 -1152 227 -1024
rect 240 -1025 241 -1013
rect 250 -1093 251 -1024
rect 254 -1025 255 -1013
rect 702 -1025 703 -1013
rect 705 -1025 706 -1013
rect 1451 -1152 1452 -1024
rect 23 -1027 24 -1013
rect 44 -1152 45 -1026
rect 96 -1027 97 -1013
rect 583 -1027 584 -1013
rect 590 -1027 591 -1013
rect 688 -1152 689 -1026
rect 691 -1027 692 -1013
rect 968 -1152 969 -1026
rect 992 -1027 993 -1013
rect 1059 -1027 1060 -1013
rect 1108 -1027 1109 -1013
rect 1234 -1152 1235 -1026
rect 1255 -1027 1256 -1013
rect 1409 -1152 1410 -1026
rect 1437 -1027 1438 -1013
rect 1598 -1152 1599 -1026
rect 23 -1152 24 -1028
rect 40 -1152 41 -1028
rect 107 -1029 108 -1013
rect 142 -1029 143 -1013
rect 170 -1029 171 -1013
rect 170 -1152 171 -1028
rect 170 -1029 171 -1013
rect 170 -1152 171 -1028
rect 184 -1029 185 -1013
rect 334 -1029 335 -1013
rect 345 -1029 346 -1013
rect 345 -1152 346 -1028
rect 345 -1029 346 -1013
rect 345 -1152 346 -1028
rect 376 -1029 377 -1013
rect 569 -1029 570 -1013
rect 576 -1029 577 -1013
rect 597 -1029 598 -1013
rect 600 -1029 601 -1013
rect 1255 -1152 1256 -1028
rect 1283 -1029 1284 -1013
rect 1444 -1152 1445 -1028
rect 37 -1031 38 -1013
rect 597 -1152 598 -1030
rect 607 -1152 608 -1030
rect 1052 -1031 1053 -1013
rect 1143 -1031 1144 -1013
rect 1283 -1152 1284 -1030
rect 1297 -1031 1298 -1013
rect 1479 -1152 1480 -1030
rect 37 -1152 38 -1032
rect 58 -1033 59 -1013
rect 107 -1152 108 -1032
rect 177 -1033 178 -1013
rect 184 -1152 185 -1032
rect 352 -1033 353 -1013
rect 390 -1152 391 -1032
rect 1066 -1033 1067 -1013
rect 1192 -1033 1193 -1013
rect 1472 -1152 1473 -1032
rect 33 -1152 34 -1034
rect 177 -1152 178 -1034
rect 201 -1152 202 -1034
rect 219 -1152 220 -1034
rect 240 -1152 241 -1034
rect 754 -1035 755 -1013
rect 842 -1035 843 -1013
rect 905 -1152 906 -1034
rect 940 -1035 941 -1013
rect 1059 -1152 1060 -1034
rect 1192 -1152 1193 -1034
rect 1213 -1035 1214 -1013
rect 1304 -1035 1305 -1013
rect 1423 -1152 1424 -1034
rect 58 -1152 59 -1036
rect 198 -1037 199 -1013
rect 247 -1037 248 -1013
rect 576 -1152 577 -1036
rect 593 -1152 594 -1036
rect 1318 -1037 1319 -1013
rect 1332 -1037 1333 -1013
rect 1500 -1152 1501 -1036
rect 79 -1039 80 -1013
rect 842 -1152 843 -1038
rect 856 -1039 857 -1013
rect 891 -1039 892 -1013
rect 940 -1152 941 -1038
rect 996 -1039 997 -1013
rect 1052 -1152 1053 -1038
rect 1458 -1039 1459 -1013
rect 86 -1041 87 -1013
rect 198 -1152 199 -1040
rect 247 -1152 248 -1040
rect 275 -1041 276 -1013
rect 394 -1041 395 -1013
rect 551 -1041 552 -1013
rect 569 -1152 570 -1040
rect 695 -1041 696 -1013
rect 702 -1152 703 -1040
rect 709 -1041 710 -1013
rect 716 -1041 717 -1013
rect 754 -1152 755 -1040
rect 758 -1152 759 -1040
rect 856 -1152 857 -1040
rect 859 -1041 860 -1013
rect 1416 -1041 1417 -1013
rect 114 -1043 115 -1013
rect 268 -1152 269 -1042
rect 275 -1152 276 -1042
rect 352 -1152 353 -1042
rect 415 -1043 416 -1013
rect 583 -1152 584 -1042
rect 611 -1043 612 -1013
rect 716 -1152 717 -1042
rect 719 -1152 720 -1042
rect 1325 -1152 1326 -1042
rect 1339 -1043 1340 -1013
rect 1507 -1152 1508 -1042
rect 114 -1152 115 -1044
rect 296 -1045 297 -1013
rect 331 -1045 332 -1013
rect 695 -1152 696 -1044
rect 733 -1152 734 -1044
rect 1038 -1152 1039 -1044
rect 1136 -1045 1137 -1013
rect 1213 -1152 1214 -1044
rect 1290 -1045 1291 -1013
rect 1458 -1152 1459 -1044
rect 30 -1047 31 -1013
rect 331 -1152 332 -1046
rect 408 -1047 409 -1013
rect 415 -1152 416 -1046
rect 422 -1047 423 -1013
rect 422 -1152 423 -1046
rect 422 -1047 423 -1013
rect 422 -1152 423 -1046
rect 432 -1152 433 -1046
rect 660 -1047 661 -1013
rect 663 -1152 664 -1046
rect 1577 -1152 1578 -1046
rect 30 -1152 31 -1048
rect 86 -1152 87 -1048
rect 142 -1152 143 -1048
rect 205 -1049 206 -1013
rect 254 -1152 255 -1048
rect 632 -1049 633 -1013
rect 660 -1152 661 -1048
rect 814 -1049 815 -1013
rect 859 -1152 860 -1048
rect 1437 -1152 1438 -1048
rect 156 -1051 157 -1013
rect 296 -1152 297 -1050
rect 338 -1051 339 -1013
rect 632 -1152 633 -1050
rect 667 -1051 668 -1013
rect 821 -1152 822 -1050
rect 863 -1051 864 -1013
rect 989 -1152 990 -1050
rect 996 -1152 997 -1050
rect 1024 -1051 1025 -1013
rect 1171 -1051 1172 -1013
rect 1318 -1152 1319 -1050
rect 1346 -1051 1347 -1013
rect 1521 -1152 1522 -1050
rect 135 -1053 136 -1013
rect 156 -1152 157 -1052
rect 205 -1152 206 -1052
rect 824 -1053 825 -1013
rect 870 -1053 871 -1013
rect 1402 -1053 1403 -1013
rect 121 -1055 122 -1013
rect 135 -1152 136 -1054
rect 261 -1055 262 -1013
rect 373 -1055 374 -1013
rect 408 -1152 409 -1054
rect 681 -1055 682 -1013
rect 730 -1055 731 -1013
rect 814 -1152 815 -1054
rect 936 -1152 937 -1054
rect 1290 -1152 1291 -1054
rect 1311 -1152 1312 -1054
rect 1430 -1055 1431 -1013
rect 121 -1152 122 -1056
rect 191 -1057 192 -1013
rect 212 -1057 213 -1013
rect 261 -1152 262 -1056
rect 338 -1152 339 -1056
rect 481 -1057 482 -1013
rect 485 -1057 486 -1013
rect 548 -1152 549 -1056
rect 562 -1057 563 -1013
rect 709 -1152 710 -1056
rect 747 -1057 748 -1013
rect 807 -1057 808 -1013
rect 954 -1057 955 -1013
rect 1066 -1152 1067 -1056
rect 1178 -1057 1179 -1013
rect 1332 -1152 1333 -1056
rect 1353 -1057 1354 -1013
rect 1528 -1152 1529 -1056
rect 9 -1059 10 -1013
rect 212 -1152 213 -1058
rect 359 -1059 360 -1013
rect 373 -1152 374 -1058
rect 394 -1152 395 -1058
rect 730 -1152 731 -1058
rect 793 -1152 794 -1058
rect 1402 -1152 1403 -1058
rect 145 -1061 146 -1013
rect 191 -1152 192 -1060
rect 359 -1152 360 -1060
rect 380 -1061 381 -1013
rect 446 -1152 447 -1060
rect 1024 -1152 1025 -1060
rect 1045 -1061 1046 -1013
rect 1171 -1152 1172 -1060
rect 1185 -1061 1186 -1013
rect 1339 -1152 1340 -1060
rect 1367 -1061 1368 -1013
rect 1563 -1152 1564 -1060
rect 163 -1063 164 -1013
rect 380 -1152 381 -1062
rect 460 -1152 461 -1062
rect 1276 -1152 1277 -1062
rect 1374 -1063 1375 -1013
rect 1542 -1152 1543 -1062
rect 166 -1152 167 -1064
rect 1178 -1152 1179 -1064
rect 1199 -1065 1200 -1013
rect 1353 -1152 1354 -1064
rect 1381 -1065 1382 -1013
rect 1549 -1152 1550 -1064
rect 464 -1067 465 -1013
rect 870 -1152 871 -1066
rect 933 -1067 934 -1013
rect 1045 -1152 1046 -1066
rect 1073 -1067 1074 -1013
rect 1185 -1152 1186 -1066
rect 1220 -1067 1221 -1013
rect 1374 -1152 1375 -1066
rect 1388 -1067 1389 -1013
rect 1556 -1152 1557 -1066
rect 9 -1152 10 -1068
rect 1220 -1152 1221 -1068
rect 1227 -1069 1228 -1013
rect 1381 -1152 1382 -1068
rect 1395 -1069 1396 -1013
rect 1584 -1152 1585 -1068
rect 243 -1071 244 -1013
rect 464 -1152 465 -1070
rect 478 -1071 479 -1013
rect 520 -1071 521 -1013
rect 534 -1071 535 -1013
rect 1416 -1152 1417 -1070
rect 429 -1073 430 -1013
rect 478 -1152 479 -1072
rect 485 -1152 486 -1072
rect 828 -1073 829 -1013
rect 933 -1152 934 -1072
rect 1269 -1073 1270 -1013
rect 492 -1075 493 -1013
rect 1346 -1152 1347 -1074
rect 355 -1152 356 -1076
rect 492 -1152 493 -1076
rect 495 -1077 496 -1013
rect 863 -1152 864 -1076
rect 947 -1077 948 -1013
rect 1073 -1152 1074 -1076
rect 1080 -1077 1081 -1013
rect 1367 -1152 1368 -1076
rect 499 -1079 500 -1013
rect 534 -1152 535 -1078
rect 544 -1079 545 -1013
rect 681 -1152 682 -1078
rect 828 -1152 829 -1078
rect 1136 -1152 1137 -1078
rect 1241 -1079 1242 -1013
rect 1388 -1152 1389 -1078
rect 471 -1081 472 -1013
rect 499 -1152 500 -1080
rect 555 -1081 556 -1013
rect 807 -1152 808 -1080
rect 877 -1081 878 -1013
rect 947 -1152 948 -1080
rect 954 -1152 955 -1080
rect 1493 -1152 1494 -1080
rect 443 -1083 444 -1013
rect 471 -1152 472 -1082
rect 555 -1152 556 -1082
rect 873 -1083 874 -1013
rect 957 -1152 958 -1082
rect 1157 -1083 1158 -1013
rect 1248 -1083 1249 -1013
rect 1395 -1152 1396 -1082
rect 443 -1152 444 -1084
rect 1143 -1152 1144 -1084
rect 1248 -1152 1249 -1084
rect 1360 -1085 1361 -1013
rect 562 -1152 563 -1086
rect 831 -1087 832 -1013
rect 835 -1087 836 -1013
rect 877 -1152 878 -1086
rect 975 -1087 976 -1013
rect 1108 -1152 1109 -1086
rect 1115 -1087 1116 -1013
rect 1227 -1152 1228 -1086
rect 1262 -1087 1263 -1013
rect 1430 -1152 1431 -1086
rect 79 -1152 80 -1088
rect 1262 -1152 1263 -1088
rect 611 -1152 612 -1090
rect 772 -1091 773 -1013
rect 779 -1091 780 -1013
rect 1115 -1152 1116 -1090
rect 1129 -1091 1130 -1013
rect 1269 -1152 1270 -1090
rect 772 -1152 773 -1092
rect 831 -1152 832 -1092
rect 1304 -1152 1305 -1092
rect 628 -1152 629 -1094
rect 1297 -1152 1298 -1094
rect 653 -1097 654 -1013
rect 1080 -1152 1081 -1096
rect 1087 -1097 1088 -1013
rect 1241 -1152 1242 -1096
rect 604 -1099 605 -1013
rect 653 -1152 654 -1098
rect 670 -1152 671 -1098
rect 1164 -1152 1165 -1098
rect 1206 -1099 1207 -1013
rect 1360 -1152 1361 -1098
rect 674 -1101 675 -1013
rect 1465 -1152 1466 -1100
rect 674 -1152 675 -1102
rect 744 -1103 745 -1013
rect 751 -1103 752 -1013
rect 779 -1152 780 -1102
rect 835 -1152 836 -1102
rect 982 -1103 983 -1013
rect 1003 -1103 1004 -1013
rect 1157 -1152 1158 -1102
rect 513 -1105 514 -1013
rect 744 -1152 745 -1104
rect 751 -1152 752 -1104
rect 1122 -1105 1123 -1013
rect 401 -1107 402 -1013
rect 513 -1152 514 -1106
rect 639 -1107 640 -1013
rect 982 -1152 983 -1106
rect 1003 -1152 1004 -1106
rect 1017 -1107 1018 -1013
rect 1094 -1107 1095 -1013
rect 1199 -1152 1200 -1106
rect 401 -1152 402 -1108
rect 450 -1109 451 -1013
rect 457 -1109 458 -1013
rect 639 -1152 640 -1108
rect 884 -1109 885 -1013
rect 1129 -1152 1130 -1108
rect 450 -1152 451 -1110
rect 646 -1111 647 -1013
rect 737 -1111 738 -1013
rect 884 -1152 885 -1110
rect 912 -1111 913 -1013
rect 1017 -1152 1018 -1110
rect 1031 -1111 1032 -1013
rect 1094 -1152 1095 -1110
rect 1101 -1111 1102 -1013
rect 1206 -1152 1207 -1110
rect 457 -1152 458 -1112
rect 520 -1152 521 -1112
rect 604 -1152 605 -1112
rect 912 -1152 913 -1112
rect 919 -1113 920 -1013
rect 1122 -1152 1123 -1112
rect 625 -1115 626 -1013
rect 646 -1152 647 -1114
rect 723 -1115 724 -1013
rect 1031 -1152 1032 -1114
rect 282 -1117 283 -1013
rect 723 -1152 724 -1116
rect 737 -1152 738 -1116
rect 761 -1117 762 -1013
rect 849 -1117 850 -1013
rect 1101 -1152 1102 -1116
rect 282 -1152 283 -1118
rect 590 -1152 591 -1118
rect 849 -1152 850 -1118
rect 1010 -1119 1011 -1013
rect 317 -1121 318 -1013
rect 625 -1152 626 -1120
rect 898 -1121 899 -1013
rect 919 -1152 920 -1120
rect 926 -1121 927 -1013
rect 1010 -1152 1011 -1120
rect 100 -1123 101 -1013
rect 317 -1152 318 -1122
rect 436 -1123 437 -1013
rect 898 -1152 899 -1122
rect 961 -1123 962 -1013
rect 1087 -1152 1088 -1122
rect 100 -1152 101 -1124
rect 303 -1125 304 -1013
rect 387 -1125 388 -1013
rect 436 -1152 437 -1124
rect 786 -1125 787 -1013
rect 926 -1152 927 -1124
rect 975 -1152 976 -1124
rect 1426 -1125 1427 -1013
rect 65 -1127 66 -1013
rect 303 -1152 304 -1126
rect 667 -1152 668 -1126
rect 786 -1152 787 -1126
rect 800 -1127 801 -1013
rect 961 -1152 962 -1126
rect 51 -1129 52 -1013
rect 65 -1152 66 -1128
rect 765 -1129 766 -1013
rect 800 -1152 801 -1128
rect 16 -1131 17 -1013
rect 765 -1152 766 -1130
rect 16 -1152 17 -1132
rect 289 -1133 290 -1013
rect 51 -1152 52 -1134
rect 506 -1135 507 -1013
rect 233 -1137 234 -1013
rect 289 -1152 290 -1136
rect 506 -1152 507 -1136
rect 677 -1137 678 -1013
rect 149 -1139 150 -1013
rect 233 -1152 234 -1138
rect 128 -1141 129 -1013
rect 149 -1152 150 -1140
rect 128 -1152 129 -1142
rect 618 -1143 619 -1013
rect 527 -1145 528 -1013
rect 618 -1152 619 -1144
rect 366 -1147 367 -1013
rect 527 -1152 528 -1146
rect 324 -1149 325 -1013
rect 366 -1152 367 -1148
rect 324 -1152 325 -1150
rect 387 -1152 388 -1150
rect 9 -1162 10 -1160
rect 303 -1162 304 -1160
rect 341 -1277 342 -1161
rect 345 -1162 346 -1160
rect 352 -1162 353 -1160
rect 667 -1162 668 -1160
rect 670 -1162 671 -1160
rect 800 -1162 801 -1160
rect 828 -1162 829 -1160
rect 1122 -1162 1123 -1160
rect 1248 -1162 1249 -1160
rect 1251 -1162 1252 -1160
rect 9 -1277 10 -1163
rect 607 -1277 608 -1163
rect 667 -1277 668 -1163
rect 772 -1164 773 -1160
rect 782 -1277 783 -1163
rect 807 -1164 808 -1160
rect 828 -1277 829 -1163
rect 863 -1164 864 -1160
rect 894 -1164 895 -1160
rect 1367 -1164 1368 -1160
rect 12 -1166 13 -1160
rect 44 -1166 45 -1160
rect 61 -1277 62 -1165
rect 597 -1166 598 -1160
rect 674 -1166 675 -1160
rect 674 -1277 675 -1165
rect 674 -1166 675 -1160
rect 674 -1277 675 -1165
rect 719 -1166 720 -1160
rect 1129 -1166 1130 -1160
rect 1248 -1277 1249 -1165
rect 1451 -1166 1452 -1160
rect 23 -1168 24 -1160
rect 23 -1277 24 -1167
rect 23 -1168 24 -1160
rect 23 -1277 24 -1167
rect 30 -1277 31 -1167
rect 702 -1168 703 -1160
rect 719 -1277 720 -1167
rect 1458 -1168 1459 -1160
rect 33 -1170 34 -1160
rect 289 -1170 290 -1160
rect 310 -1170 311 -1160
rect 345 -1277 346 -1169
rect 408 -1170 409 -1160
rect 954 -1170 955 -1160
rect 957 -1170 958 -1160
rect 1528 -1170 1529 -1160
rect 37 -1172 38 -1160
rect 723 -1172 724 -1160
rect 730 -1172 731 -1160
rect 1472 -1172 1473 -1160
rect 1528 -1277 1529 -1171
rect 1563 -1172 1564 -1160
rect 37 -1277 38 -1173
rect 758 -1174 759 -1160
rect 772 -1277 773 -1173
rect 933 -1174 934 -1160
rect 954 -1277 955 -1173
rect 982 -1174 983 -1160
rect 989 -1174 990 -1160
rect 992 -1182 993 -1173
rect 1055 -1277 1056 -1173
rect 1563 -1277 1564 -1173
rect 40 -1176 41 -1160
rect 583 -1176 584 -1160
rect 597 -1277 598 -1175
rect 639 -1176 640 -1160
rect 702 -1277 703 -1175
rect 1269 -1176 1270 -1160
rect 1367 -1277 1368 -1175
rect 1402 -1176 1403 -1160
rect 1451 -1277 1452 -1175
rect 1500 -1176 1501 -1160
rect 44 -1277 45 -1177
rect 93 -1178 94 -1160
rect 103 -1277 104 -1177
rect 422 -1178 423 -1160
rect 457 -1178 458 -1160
rect 618 -1178 619 -1160
rect 625 -1178 626 -1160
rect 982 -1277 983 -1177
rect 989 -1277 990 -1177
rect 1122 -1277 1123 -1177
rect 1143 -1178 1144 -1160
rect 1171 -1178 1172 -1160
rect 1472 -1277 1473 -1177
rect 51 -1180 52 -1160
rect 457 -1277 458 -1179
rect 481 -1277 482 -1179
rect 1297 -1180 1298 -1160
rect 1381 -1180 1382 -1160
rect 1458 -1277 1459 -1179
rect 51 -1277 52 -1181
rect 177 -1182 178 -1160
rect 184 -1182 185 -1160
rect 733 -1182 734 -1160
rect 754 -1182 755 -1160
rect 1059 -1182 1060 -1160
rect 1143 -1277 1144 -1181
rect 1164 -1182 1165 -1160
rect 1251 -1277 1252 -1181
rect 1500 -1277 1501 -1181
rect 72 -1184 73 -1160
rect 72 -1277 73 -1183
rect 72 -1184 73 -1160
rect 72 -1277 73 -1183
rect 79 -1184 80 -1160
rect 100 -1184 101 -1160
rect 107 -1184 108 -1160
rect 593 -1184 594 -1160
rect 618 -1277 619 -1183
rect 751 -1184 752 -1160
rect 758 -1277 759 -1183
rect 821 -1184 822 -1160
rect 831 -1184 832 -1160
rect 1108 -1184 1109 -1160
rect 1164 -1277 1165 -1183
rect 1206 -1184 1207 -1160
rect 1297 -1277 1298 -1183
rect 1325 -1184 1326 -1160
rect 1381 -1277 1382 -1183
rect 1437 -1184 1438 -1160
rect 79 -1277 80 -1185
rect 387 -1186 388 -1160
rect 408 -1277 409 -1185
rect 485 -1186 486 -1160
rect 506 -1186 507 -1160
rect 859 -1186 860 -1160
rect 863 -1277 864 -1185
rect 877 -1186 878 -1160
rect 922 -1277 923 -1185
rect 1374 -1186 1375 -1160
rect 1402 -1277 1403 -1185
rect 1423 -1186 1424 -1160
rect 82 -1188 83 -1160
rect 464 -1188 465 -1160
rect 485 -1277 486 -1187
rect 562 -1188 563 -1160
rect 569 -1188 570 -1160
rect 821 -1277 822 -1187
rect 835 -1188 836 -1160
rect 936 -1188 937 -1160
rect 996 -1188 997 -1160
rect 1108 -1277 1109 -1187
rect 1192 -1188 1193 -1160
rect 1325 -1277 1326 -1187
rect 1374 -1277 1375 -1187
rect 1430 -1188 1431 -1160
rect 86 -1190 87 -1160
rect 107 -1277 108 -1189
rect 114 -1190 115 -1160
rect 506 -1277 507 -1189
rect 509 -1277 510 -1189
rect 870 -1190 871 -1160
rect 877 -1277 878 -1189
rect 905 -1190 906 -1160
rect 1059 -1277 1060 -1189
rect 1136 -1190 1137 -1160
rect 1192 -1277 1193 -1189
rect 1388 -1190 1389 -1160
rect 1430 -1277 1431 -1189
rect 1479 -1190 1480 -1160
rect 86 -1277 87 -1191
rect 198 -1192 199 -1160
rect 205 -1192 206 -1160
rect 303 -1277 304 -1191
rect 310 -1277 311 -1191
rect 663 -1192 664 -1160
rect 723 -1277 724 -1191
rect 1017 -1192 1018 -1160
rect 1136 -1277 1137 -1191
rect 1157 -1192 1158 -1160
rect 1206 -1277 1207 -1191
rect 1227 -1192 1228 -1160
rect 1262 -1192 1263 -1160
rect 1423 -1277 1424 -1191
rect 1479 -1277 1480 -1191
rect 1549 -1192 1550 -1160
rect 93 -1277 94 -1193
rect 716 -1194 717 -1160
rect 730 -1277 731 -1193
rect 1080 -1194 1081 -1160
rect 1157 -1277 1158 -1193
rect 1174 -1277 1175 -1193
rect 1227 -1277 1228 -1193
rect 1255 -1194 1256 -1160
rect 1262 -1277 1263 -1193
rect 1486 -1194 1487 -1160
rect 100 -1277 101 -1195
rect 996 -1277 997 -1195
rect 1080 -1277 1081 -1195
rect 1094 -1196 1095 -1160
rect 1255 -1277 1256 -1195
rect 1311 -1196 1312 -1160
rect 1360 -1196 1361 -1160
rect 1486 -1277 1487 -1195
rect 114 -1277 115 -1197
rect 478 -1198 479 -1160
rect 513 -1198 514 -1160
rect 604 -1198 605 -1160
rect 611 -1198 612 -1160
rect 870 -1277 871 -1197
rect 905 -1277 906 -1197
rect 919 -1198 920 -1160
rect 940 -1198 941 -1160
rect 1017 -1277 1018 -1197
rect 1311 -1277 1312 -1197
rect 1332 -1198 1333 -1160
rect 1360 -1277 1361 -1197
rect 1395 -1198 1396 -1160
rect 2 -1200 3 -1160
rect 478 -1277 479 -1199
rect 541 -1200 542 -1160
rect 625 -1277 626 -1199
rect 639 -1277 640 -1199
rect 646 -1200 647 -1160
rect 653 -1200 654 -1160
rect 1549 -1277 1550 -1199
rect 2 -1277 3 -1201
rect 975 -1202 976 -1160
rect 1003 -1202 1004 -1160
rect 1094 -1277 1095 -1201
rect 1220 -1202 1221 -1160
rect 1332 -1277 1333 -1201
rect 1388 -1277 1389 -1201
rect 1542 -1202 1543 -1160
rect 121 -1204 122 -1160
rect 530 -1277 531 -1203
rect 541 -1277 542 -1203
rect 555 -1204 556 -1160
rect 583 -1277 584 -1203
rect 765 -1204 766 -1160
rect 786 -1204 787 -1160
rect 807 -1277 808 -1203
rect 856 -1204 857 -1160
rect 1507 -1204 1508 -1160
rect 1542 -1277 1543 -1203
rect 1598 -1204 1599 -1160
rect 121 -1277 122 -1205
rect 268 -1206 269 -1160
rect 282 -1206 283 -1160
rect 282 -1277 283 -1205
rect 282 -1206 283 -1160
rect 282 -1277 283 -1205
rect 289 -1277 290 -1205
rect 338 -1206 339 -1160
rect 366 -1206 367 -1160
rect 387 -1277 388 -1205
rect 394 -1206 395 -1160
rect 716 -1277 717 -1205
rect 751 -1277 752 -1205
rect 1129 -1277 1130 -1205
rect 1395 -1277 1396 -1205
rect 1444 -1206 1445 -1160
rect 1507 -1277 1508 -1205
rect 1570 -1206 1571 -1160
rect 131 -1277 132 -1207
rect 919 -1277 920 -1207
rect 936 -1277 937 -1207
rect 1220 -1277 1221 -1207
rect 1276 -1208 1277 -1160
rect 1444 -1277 1445 -1207
rect 166 -1210 167 -1160
rect 898 -1210 899 -1160
rect 940 -1277 941 -1209
rect 961 -1210 962 -1160
rect 975 -1277 976 -1209
rect 1073 -1210 1074 -1160
rect 1150 -1210 1151 -1160
rect 1276 -1277 1277 -1209
rect 177 -1277 178 -1211
rect 247 -1212 248 -1160
rect 254 -1212 255 -1160
rect 933 -1277 934 -1211
rect 961 -1277 962 -1211
rect 1045 -1212 1046 -1160
rect 1150 -1277 1151 -1211
rect 1178 -1212 1179 -1160
rect 16 -1214 17 -1160
rect 247 -1277 248 -1213
rect 261 -1214 262 -1160
rect 268 -1277 269 -1213
rect 362 -1277 363 -1213
rect 1045 -1277 1046 -1213
rect 1178 -1277 1179 -1213
rect 1318 -1214 1319 -1160
rect 16 -1277 17 -1215
rect 275 -1216 276 -1160
rect 366 -1277 367 -1215
rect 373 -1216 374 -1160
rect 394 -1277 395 -1215
rect 415 -1216 416 -1160
rect 422 -1277 423 -1215
rect 460 -1216 461 -1160
rect 520 -1216 521 -1160
rect 646 -1277 647 -1215
rect 653 -1277 654 -1215
rect 737 -1216 738 -1160
rect 765 -1277 766 -1215
rect 1115 -1216 1116 -1160
rect 1318 -1277 1319 -1215
rect 1346 -1216 1347 -1160
rect 65 -1218 66 -1160
rect 254 -1277 255 -1217
rect 275 -1277 276 -1217
rect 429 -1218 430 -1160
rect 436 -1218 437 -1160
rect 464 -1277 465 -1217
rect 520 -1277 521 -1217
rect 1535 -1218 1536 -1160
rect 65 -1277 66 -1219
rect 527 -1220 528 -1160
rect 548 -1220 549 -1160
rect 562 -1277 563 -1219
rect 590 -1220 591 -1160
rect 1346 -1277 1347 -1219
rect 1535 -1277 1536 -1219
rect 1584 -1220 1585 -1160
rect 170 -1222 171 -1160
rect 261 -1277 262 -1221
rect 317 -1222 318 -1160
rect 436 -1277 437 -1221
rect 527 -1277 528 -1221
rect 1269 -1277 1270 -1221
rect 170 -1277 171 -1223
rect 352 -1277 353 -1223
rect 373 -1277 374 -1223
rect 499 -1224 500 -1160
rect 548 -1277 549 -1223
rect 611 -1277 612 -1223
rect 628 -1224 629 -1160
rect 1003 -1277 1004 -1223
rect 184 -1277 185 -1225
rect 558 -1277 559 -1225
rect 590 -1277 591 -1225
rect 681 -1226 682 -1160
rect 744 -1226 745 -1160
rect 1115 -1277 1116 -1225
rect 191 -1228 192 -1160
rect 205 -1277 206 -1227
rect 212 -1228 213 -1160
rect 446 -1228 447 -1160
rect 555 -1277 556 -1227
rect 1591 -1228 1592 -1160
rect 191 -1277 192 -1229
rect 233 -1230 234 -1160
rect 240 -1230 241 -1160
rect 415 -1277 416 -1229
rect 429 -1277 430 -1229
rect 471 -1230 472 -1160
rect 604 -1277 605 -1229
rect 1283 -1230 1284 -1160
rect 58 -1232 59 -1160
rect 240 -1277 241 -1231
rect 338 -1277 339 -1231
rect 744 -1277 745 -1231
rect 786 -1277 787 -1231
rect 842 -1232 843 -1160
rect 859 -1277 860 -1231
rect 1353 -1232 1354 -1160
rect 149 -1234 150 -1160
rect 233 -1277 234 -1233
rect 380 -1234 381 -1160
rect 499 -1277 500 -1233
rect 681 -1277 682 -1233
rect 688 -1234 689 -1160
rect 796 -1234 797 -1160
rect 1010 -1234 1011 -1160
rect 1199 -1234 1200 -1160
rect 1283 -1277 1284 -1233
rect 1353 -1277 1354 -1233
rect 1493 -1234 1494 -1160
rect 128 -1236 129 -1160
rect 688 -1277 689 -1235
rect 768 -1277 769 -1235
rect 1199 -1277 1200 -1235
rect 1409 -1236 1410 -1160
rect 1493 -1277 1494 -1235
rect 149 -1277 150 -1237
rect 660 -1238 661 -1160
rect 800 -1277 801 -1237
rect 849 -1238 850 -1160
rect 898 -1277 899 -1237
rect 947 -1238 948 -1160
rect 1010 -1277 1011 -1237
rect 1066 -1238 1067 -1160
rect 1409 -1277 1410 -1237
rect 1416 -1238 1417 -1160
rect 198 -1277 199 -1239
rect 317 -1277 318 -1239
rect 401 -1240 402 -1160
rect 569 -1277 570 -1239
rect 660 -1277 661 -1239
rect 726 -1277 727 -1239
rect 814 -1240 815 -1160
rect 856 -1277 857 -1239
rect 947 -1277 948 -1239
rect 968 -1240 969 -1160
rect 1066 -1277 1067 -1239
rect 1087 -1240 1088 -1160
rect 1416 -1277 1417 -1239
rect 1465 -1240 1466 -1160
rect 212 -1277 213 -1241
rect 359 -1242 360 -1160
rect 401 -1277 402 -1241
rect 576 -1242 577 -1160
rect 632 -1242 633 -1160
rect 814 -1277 815 -1241
rect 838 -1277 839 -1241
rect 1073 -1277 1074 -1241
rect 1087 -1277 1088 -1241
rect 1101 -1242 1102 -1160
rect 1465 -1277 1466 -1241
rect 1514 -1242 1515 -1160
rect 219 -1244 220 -1160
rect 513 -1277 514 -1243
rect 576 -1277 577 -1243
rect 926 -1244 927 -1160
rect 968 -1277 969 -1243
rect 1024 -1244 1025 -1160
rect 1514 -1277 1515 -1243
rect 1577 -1244 1578 -1160
rect 142 -1246 143 -1160
rect 219 -1277 220 -1245
rect 226 -1246 227 -1160
rect 390 -1246 391 -1160
rect 450 -1246 451 -1160
rect 842 -1277 843 -1245
rect 849 -1277 850 -1245
rect 884 -1246 885 -1160
rect 912 -1246 913 -1160
rect 1101 -1277 1102 -1245
rect 58 -1277 59 -1247
rect 884 -1277 885 -1247
rect 926 -1277 927 -1247
rect 1052 -1248 1053 -1160
rect 128 -1277 129 -1249
rect 142 -1277 143 -1249
rect 226 -1277 227 -1249
rect 324 -1250 325 -1160
rect 450 -1277 451 -1249
rect 534 -1250 535 -1160
rect 632 -1277 633 -1249
rect 695 -1250 696 -1160
rect 737 -1277 738 -1249
rect 1052 -1277 1053 -1249
rect 296 -1252 297 -1160
rect 380 -1277 381 -1251
rect 471 -1277 472 -1251
rect 709 -1252 710 -1160
rect 779 -1252 780 -1160
rect 912 -1277 913 -1251
rect 1024 -1277 1025 -1251
rect 1038 -1252 1039 -1160
rect 163 -1254 164 -1160
rect 709 -1277 710 -1253
rect 779 -1277 780 -1253
rect 1437 -1277 1438 -1253
rect 156 -1256 157 -1160
rect 163 -1277 164 -1255
rect 296 -1277 297 -1255
rect 492 -1256 493 -1160
rect 534 -1277 535 -1255
rect 793 -1256 794 -1160
rect 1038 -1277 1039 -1255
rect 1185 -1256 1186 -1160
rect 135 -1258 136 -1160
rect 156 -1277 157 -1257
rect 173 -1277 174 -1257
rect 793 -1277 794 -1257
rect 1185 -1277 1186 -1257
rect 1213 -1258 1214 -1160
rect 135 -1277 136 -1259
rect 359 -1277 360 -1259
rect 492 -1277 493 -1259
rect 835 -1277 836 -1259
rect 1213 -1277 1214 -1259
rect 1234 -1260 1235 -1160
rect 320 -1277 321 -1261
rect 695 -1277 696 -1261
rect 1234 -1277 1235 -1261
rect 1241 -1262 1242 -1160
rect 324 -1277 325 -1263
rect 331 -1264 332 -1160
rect 1241 -1277 1242 -1263
rect 1290 -1264 1291 -1160
rect 331 -1277 332 -1265
rect 443 -1266 444 -1160
rect 1290 -1277 1291 -1265
rect 1304 -1266 1305 -1160
rect 443 -1277 444 -1267
rect 754 -1277 755 -1267
rect 1304 -1277 1305 -1267
rect 1339 -1268 1340 -1160
rect 1339 -1277 1340 -1269
rect 1521 -1270 1522 -1160
rect 1521 -1277 1522 -1271
rect 1556 -1272 1557 -1160
rect 891 -1274 892 -1160
rect 1556 -1277 1557 -1273
rect 355 -1276 356 -1160
rect 891 -1277 892 -1275
rect 2 -1287 3 -1285
rect 555 -1287 556 -1285
rect 562 -1287 563 -1285
rect 604 -1287 605 -1285
rect 649 -1396 650 -1286
rect 1486 -1287 1487 -1285
rect 2 -1396 3 -1288
rect 373 -1289 374 -1285
rect 478 -1289 479 -1285
rect 1290 -1289 1291 -1285
rect 1409 -1289 1410 -1285
rect 1409 -1396 1410 -1288
rect 1409 -1289 1410 -1285
rect 1409 -1396 1410 -1288
rect 1451 -1289 1452 -1285
rect 1454 -1307 1455 -1288
rect 1486 -1396 1487 -1288
rect 1514 -1289 1515 -1285
rect 23 -1291 24 -1285
rect 23 -1396 24 -1290
rect 23 -1291 24 -1285
rect 23 -1396 24 -1290
rect 30 -1291 31 -1285
rect 754 -1291 755 -1285
rect 765 -1291 766 -1285
rect 1346 -1291 1347 -1285
rect 1451 -1396 1452 -1290
rect 1465 -1291 1466 -1285
rect 1514 -1396 1515 -1290
rect 1542 -1291 1543 -1285
rect 30 -1396 31 -1292
rect 44 -1293 45 -1285
rect 61 -1293 62 -1285
rect 1472 -1293 1473 -1285
rect 37 -1295 38 -1285
rect 520 -1295 521 -1285
rect 527 -1295 528 -1285
rect 541 -1295 542 -1285
rect 548 -1295 549 -1285
rect 1549 -1295 1550 -1285
rect 37 -1396 38 -1296
rect 443 -1297 444 -1285
rect 488 -1396 489 -1296
rect 499 -1297 500 -1285
rect 509 -1297 510 -1285
rect 982 -1297 983 -1285
rect 1052 -1297 1053 -1285
rect 1458 -1297 1459 -1285
rect 1472 -1396 1473 -1296
rect 1479 -1297 1480 -1285
rect 44 -1396 45 -1298
rect 240 -1299 241 -1285
rect 268 -1299 269 -1285
rect 268 -1396 269 -1298
rect 268 -1299 269 -1285
rect 268 -1396 269 -1298
rect 282 -1299 283 -1285
rect 282 -1396 283 -1298
rect 282 -1299 283 -1285
rect 282 -1396 283 -1298
rect 338 -1396 339 -1298
rect 408 -1299 409 -1285
rect 422 -1299 423 -1285
rect 443 -1396 444 -1298
rect 467 -1396 468 -1298
rect 499 -1396 500 -1298
rect 548 -1396 549 -1298
rect 779 -1299 780 -1285
rect 782 -1299 783 -1285
rect 1521 -1299 1522 -1285
rect 68 -1396 69 -1300
rect 814 -1301 815 -1285
rect 835 -1301 836 -1285
rect 1234 -1301 1235 -1285
rect 1241 -1301 1242 -1285
rect 1241 -1396 1242 -1300
rect 1241 -1301 1242 -1285
rect 1241 -1396 1242 -1300
rect 1346 -1396 1347 -1300
rect 1367 -1301 1368 -1285
rect 1388 -1301 1389 -1285
rect 1458 -1396 1459 -1300
rect 1479 -1396 1480 -1300
rect 1507 -1301 1508 -1285
rect 100 -1303 101 -1285
rect 429 -1303 430 -1285
rect 555 -1396 556 -1302
rect 674 -1303 675 -1285
rect 719 -1303 720 -1285
rect 1521 -1396 1522 -1302
rect 100 -1396 101 -1304
rect 149 -1305 150 -1285
rect 156 -1305 157 -1285
rect 156 -1396 157 -1304
rect 156 -1305 157 -1285
rect 156 -1396 157 -1304
rect 177 -1305 178 -1285
rect 320 -1305 321 -1285
rect 345 -1305 346 -1285
rect 373 -1396 374 -1304
rect 387 -1305 388 -1285
rect 429 -1396 430 -1304
rect 562 -1396 563 -1304
rect 786 -1305 787 -1285
rect 793 -1305 794 -1285
rect 1006 -1396 1007 -1304
rect 1055 -1305 1056 -1285
rect 1528 -1305 1529 -1285
rect 79 -1307 80 -1285
rect 387 -1396 388 -1306
rect 401 -1307 402 -1285
rect 541 -1396 542 -1306
rect 674 -1396 675 -1306
rect 681 -1307 682 -1285
rect 723 -1307 724 -1285
rect 1031 -1307 1032 -1285
rect 1094 -1307 1095 -1285
rect 1094 -1396 1095 -1306
rect 1094 -1307 1095 -1285
rect 1094 -1396 1095 -1306
rect 1171 -1307 1172 -1285
rect 1402 -1307 1403 -1285
rect 1465 -1396 1466 -1306
rect 1507 -1396 1508 -1306
rect 1535 -1307 1536 -1285
rect 79 -1396 80 -1308
rect 198 -1309 199 -1285
rect 233 -1309 234 -1285
rect 359 -1309 360 -1285
rect 366 -1309 367 -1285
rect 366 -1396 367 -1308
rect 366 -1309 367 -1285
rect 366 -1396 367 -1308
rect 418 -1396 419 -1308
rect 1367 -1396 1368 -1308
rect 1388 -1396 1389 -1308
rect 1430 -1309 1431 -1285
rect 1528 -1396 1529 -1308
rect 1556 -1309 1557 -1285
rect 82 -1396 83 -1310
rect 177 -1396 178 -1310
rect 191 -1311 192 -1285
rect 191 -1396 192 -1310
rect 191 -1311 192 -1285
rect 191 -1396 192 -1310
rect 198 -1396 199 -1310
rect 530 -1311 531 -1285
rect 632 -1311 633 -1285
rect 681 -1396 682 -1310
rect 723 -1396 724 -1310
rect 768 -1311 769 -1285
rect 772 -1311 773 -1285
rect 772 -1396 773 -1310
rect 772 -1311 773 -1285
rect 772 -1396 773 -1310
rect 779 -1396 780 -1310
rect 828 -1311 829 -1285
rect 835 -1396 836 -1310
rect 842 -1311 843 -1285
rect 880 -1396 881 -1310
rect 1500 -1311 1501 -1285
rect 86 -1313 87 -1285
rect 320 -1396 321 -1312
rect 345 -1396 346 -1312
rect 362 -1313 363 -1285
rect 422 -1396 423 -1312
rect 450 -1313 451 -1285
rect 481 -1313 482 -1285
rect 793 -1396 794 -1312
rect 828 -1396 829 -1312
rect 856 -1313 857 -1285
rect 922 -1313 923 -1285
rect 1444 -1313 1445 -1285
rect 86 -1396 87 -1314
rect 415 -1315 416 -1285
rect 450 -1396 451 -1314
rect 485 -1315 486 -1285
rect 604 -1396 605 -1314
rect 922 -1396 923 -1314
rect 933 -1315 934 -1285
rect 1493 -1315 1494 -1285
rect 9 -1317 10 -1285
rect 485 -1396 486 -1316
rect 737 -1317 738 -1285
rect 873 -1396 874 -1316
rect 933 -1396 934 -1316
rect 954 -1317 955 -1285
rect 975 -1317 976 -1285
rect 1052 -1396 1053 -1316
rect 1101 -1317 1102 -1285
rect 1535 -1396 1536 -1316
rect 9 -1396 10 -1318
rect 65 -1319 66 -1285
rect 93 -1319 94 -1285
rect 149 -1396 150 -1318
rect 212 -1319 213 -1285
rect 481 -1396 482 -1318
rect 667 -1319 668 -1285
rect 737 -1396 738 -1318
rect 744 -1319 745 -1285
rect 814 -1396 815 -1318
rect 838 -1319 839 -1285
rect 863 -1319 864 -1285
rect 898 -1319 899 -1285
rect 954 -1396 955 -1318
rect 982 -1396 983 -1318
rect 996 -1319 997 -1285
rect 1024 -1319 1025 -1285
rect 1031 -1396 1032 -1318
rect 1101 -1396 1102 -1318
rect 1213 -1319 1214 -1285
rect 1220 -1319 1221 -1285
rect 1220 -1396 1221 -1318
rect 1220 -1319 1221 -1285
rect 1220 -1396 1221 -1318
rect 1234 -1396 1235 -1318
rect 1262 -1319 1263 -1285
rect 1339 -1319 1340 -1285
rect 1493 -1396 1494 -1318
rect 93 -1396 94 -1320
rect 569 -1321 570 -1285
rect 618 -1321 619 -1285
rect 667 -1396 668 -1320
rect 688 -1321 689 -1285
rect 744 -1396 745 -1320
rect 751 -1321 752 -1285
rect 1311 -1321 1312 -1285
rect 1353 -1321 1354 -1285
rect 1430 -1396 1431 -1320
rect 103 -1323 104 -1285
rect 1423 -1323 1424 -1285
rect 110 -1396 111 -1324
rect 296 -1325 297 -1285
rect 303 -1325 304 -1285
rect 751 -1396 752 -1324
rect 765 -1396 766 -1324
rect 800 -1325 801 -1285
rect 849 -1325 850 -1285
rect 898 -1396 899 -1324
rect 961 -1325 962 -1285
rect 1024 -1396 1025 -1324
rect 1038 -1325 1039 -1285
rect 1213 -1396 1214 -1324
rect 1255 -1325 1256 -1285
rect 1500 -1396 1501 -1324
rect 128 -1327 129 -1285
rect 859 -1327 860 -1285
rect 863 -1396 864 -1326
rect 926 -1327 927 -1285
rect 940 -1327 941 -1285
rect 961 -1396 962 -1326
rect 996 -1396 997 -1326
rect 1003 -1327 1004 -1285
rect 1010 -1327 1011 -1285
rect 1038 -1396 1039 -1326
rect 1087 -1327 1088 -1285
rect 1339 -1396 1340 -1326
rect 1395 -1327 1396 -1285
rect 1402 -1396 1403 -1326
rect 1416 -1327 1417 -1285
rect 1423 -1396 1424 -1326
rect 107 -1329 108 -1285
rect 128 -1396 129 -1328
rect 131 -1329 132 -1285
rect 702 -1329 703 -1285
rect 712 -1396 713 -1328
rect 1262 -1396 1263 -1328
rect 1311 -1396 1312 -1328
rect 1360 -1329 1361 -1285
rect 1395 -1396 1396 -1328
rect 1437 -1329 1438 -1285
rect 107 -1396 108 -1330
rect 114 -1331 115 -1285
rect 215 -1396 216 -1330
rect 296 -1396 297 -1330
rect 303 -1396 304 -1330
rect 324 -1331 325 -1285
rect 352 -1331 353 -1285
rect 527 -1396 528 -1330
rect 618 -1396 619 -1330
rect 639 -1331 640 -1285
rect 730 -1331 731 -1285
rect 1087 -1396 1088 -1330
rect 1143 -1331 1144 -1285
rect 1171 -1396 1172 -1330
rect 1178 -1331 1179 -1285
rect 1290 -1396 1291 -1330
rect 1332 -1331 1333 -1285
rect 1437 -1396 1438 -1330
rect 16 -1333 17 -1285
rect 352 -1396 353 -1332
rect 436 -1333 437 -1285
rect 569 -1396 570 -1332
rect 639 -1396 640 -1332
rect 912 -1333 913 -1285
rect 926 -1396 927 -1332
rect 989 -1333 990 -1285
rect 1059 -1333 1060 -1285
rect 1143 -1396 1144 -1332
rect 1157 -1333 1158 -1285
rect 1444 -1396 1445 -1332
rect 16 -1396 17 -1334
rect 205 -1335 206 -1285
rect 233 -1396 234 -1334
rect 310 -1335 311 -1285
rect 436 -1396 437 -1334
rect 464 -1335 465 -1285
rect 471 -1335 472 -1285
rect 688 -1396 689 -1334
rect 786 -1396 787 -1334
rect 870 -1335 871 -1285
rect 940 -1396 941 -1334
rect 978 -1396 979 -1334
rect 989 -1396 990 -1334
rect 1150 -1335 1151 -1285
rect 1164 -1335 1165 -1285
rect 1178 -1396 1179 -1334
rect 1192 -1335 1193 -1285
rect 1353 -1396 1354 -1334
rect 1360 -1396 1361 -1334
rect 1374 -1335 1375 -1285
rect 51 -1337 52 -1285
rect 114 -1396 115 -1336
rect 170 -1337 171 -1285
rect 324 -1396 325 -1336
rect 457 -1337 458 -1285
rect 702 -1396 703 -1336
rect 800 -1396 801 -1336
rect 807 -1337 808 -1285
rect 842 -1396 843 -1336
rect 849 -1396 850 -1336
rect 856 -1396 857 -1336
rect 877 -1337 878 -1285
rect 947 -1337 948 -1285
rect 1010 -1396 1011 -1336
rect 1122 -1337 1123 -1285
rect 1157 -1396 1158 -1336
rect 1255 -1396 1256 -1336
rect 1276 -1337 1277 -1285
rect 1374 -1396 1375 -1336
rect 1381 -1337 1382 -1285
rect 51 -1396 52 -1338
rect 261 -1339 262 -1285
rect 275 -1339 276 -1285
rect 310 -1396 311 -1338
rect 317 -1339 318 -1285
rect 807 -1396 808 -1338
rect 877 -1396 878 -1338
rect 891 -1339 892 -1285
rect 905 -1339 906 -1285
rect 947 -1396 948 -1338
rect 1003 -1396 1004 -1338
rect 1059 -1396 1060 -1338
rect 1122 -1396 1123 -1338
rect 1227 -1339 1228 -1285
rect 1248 -1339 1249 -1285
rect 1381 -1396 1382 -1338
rect 65 -1396 66 -1340
rect 912 -1396 913 -1340
rect 1080 -1341 1081 -1285
rect 1248 -1396 1249 -1340
rect 1269 -1341 1270 -1285
rect 1276 -1396 1277 -1340
rect 142 -1343 143 -1285
rect 170 -1396 171 -1342
rect 184 -1343 185 -1285
rect 275 -1396 276 -1342
rect 317 -1396 318 -1342
rect 632 -1396 633 -1342
rect 695 -1343 696 -1285
rect 1269 -1396 1270 -1342
rect 58 -1345 59 -1285
rect 695 -1396 696 -1344
rect 884 -1345 885 -1285
rect 905 -1396 906 -1344
rect 1073 -1345 1074 -1285
rect 1080 -1396 1081 -1344
rect 1129 -1345 1130 -1285
rect 1332 -1396 1333 -1344
rect 58 -1396 59 -1346
rect 625 -1347 626 -1285
rect 884 -1396 885 -1346
rect 968 -1347 969 -1285
rect 1066 -1347 1067 -1285
rect 1073 -1396 1074 -1346
rect 1136 -1347 1137 -1285
rect 1164 -1396 1165 -1346
rect 1227 -1396 1228 -1346
rect 1318 -1347 1319 -1285
rect 135 -1349 136 -1285
rect 1129 -1396 1130 -1348
rect 1136 -1396 1137 -1348
rect 1199 -1349 1200 -1285
rect 1297 -1349 1298 -1285
rect 1318 -1396 1319 -1348
rect 72 -1351 73 -1285
rect 135 -1396 136 -1350
rect 142 -1396 143 -1350
rect 289 -1351 290 -1285
rect 457 -1396 458 -1350
rect 492 -1351 493 -1285
rect 495 -1396 496 -1350
rect 870 -1396 871 -1350
rect 891 -1396 892 -1350
rect 919 -1396 920 -1350
rect 1045 -1351 1046 -1285
rect 1066 -1396 1067 -1350
rect 1150 -1396 1151 -1350
rect 1185 -1351 1186 -1285
rect 1199 -1396 1200 -1350
rect 1206 -1351 1207 -1285
rect 1297 -1396 1298 -1350
rect 1325 -1351 1326 -1285
rect 72 -1396 73 -1352
rect 219 -1353 220 -1285
rect 226 -1353 227 -1285
rect 471 -1396 472 -1352
rect 478 -1396 479 -1352
rect 730 -1396 731 -1352
rect 1108 -1353 1109 -1285
rect 1206 -1396 1207 -1352
rect 1304 -1353 1305 -1285
rect 1325 -1396 1326 -1352
rect 121 -1355 122 -1285
rect 289 -1396 290 -1354
rect 464 -1396 465 -1354
rect 597 -1355 598 -1285
rect 625 -1396 626 -1354
rect 660 -1355 661 -1285
rect 709 -1355 710 -1285
rect 1108 -1396 1109 -1354
rect 1185 -1396 1186 -1354
rect 1563 -1355 1564 -1285
rect 121 -1396 122 -1356
rect 331 -1357 332 -1285
rect 492 -1396 493 -1356
rect 520 -1396 521 -1356
rect 523 -1357 524 -1285
rect 1045 -1396 1046 -1356
rect 163 -1359 164 -1285
rect 184 -1396 185 -1358
rect 205 -1396 206 -1358
rect 558 -1359 559 -1285
rect 597 -1396 598 -1358
rect 950 -1396 951 -1358
rect 1017 -1359 1018 -1285
rect 1304 -1396 1305 -1358
rect 163 -1396 164 -1360
rect 404 -1396 405 -1360
rect 506 -1361 507 -1285
rect 1416 -1396 1417 -1360
rect 219 -1396 220 -1362
rect 534 -1363 535 -1285
rect 611 -1363 612 -1285
rect 660 -1396 661 -1362
rect 709 -1396 710 -1362
rect 1115 -1363 1116 -1285
rect 226 -1396 227 -1364
rect 716 -1365 717 -1285
rect 845 -1396 846 -1364
rect 1115 -1396 1116 -1364
rect 240 -1396 241 -1366
rect 380 -1367 381 -1285
rect 390 -1396 391 -1366
rect 534 -1396 535 -1366
rect 551 -1367 552 -1285
rect 716 -1396 717 -1366
rect 247 -1369 248 -1285
rect 408 -1396 409 -1368
rect 506 -1396 507 -1368
rect 975 -1396 976 -1368
rect 247 -1396 248 -1370
rect 583 -1371 584 -1285
rect 590 -1371 591 -1285
rect 611 -1396 612 -1370
rect 254 -1373 255 -1285
rect 359 -1396 360 -1372
rect 380 -1396 381 -1372
rect 394 -1373 395 -1285
rect 513 -1373 514 -1285
rect 583 -1396 584 -1372
rect 590 -1396 591 -1372
rect 726 -1373 727 -1285
rect 212 -1396 213 -1374
rect 254 -1396 255 -1374
rect 261 -1396 262 -1374
rect 607 -1375 608 -1285
rect 331 -1396 332 -1376
rect 1017 -1396 1018 -1376
rect 394 -1396 395 -1378
rect 653 -1379 654 -1285
rect 513 -1396 514 -1380
rect 1283 -1381 1284 -1285
rect 516 -1396 517 -1382
rect 1283 -1396 1284 -1382
rect 523 -1396 524 -1384
rect 1192 -1396 1193 -1384
rect 576 -1387 577 -1285
rect 653 -1396 654 -1386
rect 576 -1396 577 -1388
rect 821 -1389 822 -1285
rect 758 -1391 759 -1285
rect 821 -1396 822 -1390
rect 646 -1393 647 -1285
rect 758 -1396 759 -1392
rect 646 -1396 647 -1394
rect 968 -1396 969 -1394
rect 23 -1406 24 -1404
rect 23 -1529 24 -1405
rect 23 -1406 24 -1404
rect 23 -1529 24 -1405
rect 44 -1406 45 -1404
rect 649 -1406 650 -1404
rect 684 -1529 685 -1405
rect 730 -1406 731 -1404
rect 800 -1406 801 -1404
rect 838 -1529 839 -1405
rect 842 -1406 843 -1404
rect 1353 -1406 1354 -1404
rect 1528 -1406 1529 -1404
rect 1528 -1529 1529 -1405
rect 1528 -1406 1529 -1404
rect 1528 -1529 1529 -1405
rect 1535 -1406 1536 -1404
rect 1535 -1529 1536 -1405
rect 1535 -1406 1536 -1404
rect 1535 -1529 1536 -1405
rect 44 -1529 45 -1407
rect 114 -1408 115 -1404
rect 121 -1408 122 -1404
rect 467 -1408 468 -1404
rect 471 -1408 472 -1404
rect 495 -1408 496 -1404
rect 520 -1408 521 -1404
rect 527 -1408 528 -1404
rect 646 -1408 647 -1404
rect 1269 -1408 1270 -1404
rect 1346 -1408 1347 -1404
rect 1346 -1529 1347 -1407
rect 1346 -1408 1347 -1404
rect 1346 -1529 1347 -1407
rect 1353 -1529 1354 -1407
rect 1360 -1408 1361 -1404
rect 51 -1410 52 -1404
rect 418 -1410 419 -1404
rect 478 -1410 479 -1404
rect 1192 -1410 1193 -1404
rect 1241 -1410 1242 -1404
rect 1241 -1529 1242 -1409
rect 1241 -1410 1242 -1404
rect 1241 -1529 1242 -1409
rect 1311 -1410 1312 -1404
rect 1360 -1529 1361 -1409
rect 51 -1529 52 -1411
rect 317 -1412 318 -1404
rect 320 -1412 321 -1404
rect 408 -1412 409 -1404
rect 478 -1529 479 -1411
rect 1143 -1412 1144 -1404
rect 1192 -1529 1193 -1411
rect 1297 -1412 1298 -1404
rect 65 -1414 66 -1404
rect 296 -1414 297 -1404
rect 366 -1414 367 -1404
rect 397 -1529 398 -1413
rect 408 -1529 409 -1413
rect 492 -1414 493 -1404
rect 499 -1414 500 -1404
rect 520 -1529 521 -1413
rect 646 -1529 647 -1413
rect 1115 -1414 1116 -1404
rect 1276 -1414 1277 -1404
rect 1311 -1529 1312 -1413
rect 65 -1529 66 -1415
rect 569 -1416 570 -1404
rect 712 -1416 713 -1404
rect 779 -1416 780 -1404
rect 800 -1529 801 -1415
rect 1304 -1416 1305 -1404
rect 82 -1418 83 -1404
rect 275 -1418 276 -1404
rect 296 -1529 297 -1417
rect 338 -1418 339 -1404
rect 390 -1418 391 -1404
rect 523 -1418 524 -1404
rect 562 -1418 563 -1404
rect 779 -1529 780 -1417
rect 807 -1418 808 -1404
rect 1269 -1529 1270 -1417
rect 68 -1420 69 -1404
rect 338 -1529 339 -1419
rect 394 -1420 395 -1404
rect 831 -1529 832 -1419
rect 842 -1529 843 -1419
rect 856 -1420 857 -1404
rect 873 -1420 874 -1404
rect 1234 -1420 1235 -1404
rect 1262 -1420 1263 -1404
rect 1276 -1529 1277 -1419
rect 82 -1529 83 -1421
rect 121 -1529 122 -1421
rect 184 -1422 185 -1404
rect 513 -1422 514 -1404
rect 562 -1529 563 -1421
rect 660 -1422 661 -1404
rect 723 -1422 724 -1404
rect 726 -1529 727 -1421
rect 730 -1529 731 -1421
rect 835 -1422 836 -1404
rect 856 -1529 857 -1421
rect 1206 -1422 1207 -1404
rect 1234 -1529 1235 -1421
rect 1521 -1422 1522 -1404
rect 93 -1424 94 -1404
rect 492 -1529 493 -1423
rect 513 -1529 514 -1423
rect 541 -1424 542 -1404
rect 569 -1529 570 -1423
rect 992 -1529 993 -1423
rect 1003 -1529 1004 -1423
rect 1045 -1424 1046 -1404
rect 1076 -1529 1077 -1423
rect 1318 -1424 1319 -1404
rect 1332 -1424 1333 -1404
rect 1521 -1529 1522 -1423
rect 37 -1426 38 -1404
rect 93 -1529 94 -1425
rect 100 -1426 101 -1404
rect 404 -1426 405 -1404
rect 464 -1426 465 -1404
rect 1143 -1529 1144 -1425
rect 1164 -1426 1165 -1404
rect 1262 -1529 1263 -1425
rect 37 -1529 38 -1427
rect 835 -1529 836 -1427
rect 880 -1428 881 -1404
rect 933 -1428 934 -1404
rect 950 -1428 951 -1404
rect 1465 -1428 1466 -1404
rect 100 -1529 101 -1429
rect 254 -1430 255 -1404
rect 268 -1430 269 -1404
rect 268 -1529 269 -1429
rect 268 -1430 269 -1404
rect 268 -1529 269 -1429
rect 275 -1529 276 -1429
rect 688 -1430 689 -1404
rect 723 -1529 724 -1429
rect 1213 -1430 1214 -1404
rect 1444 -1430 1445 -1404
rect 1465 -1529 1466 -1429
rect 103 -1529 104 -1431
rect 432 -1529 433 -1431
rect 436 -1432 437 -1404
rect 464 -1529 465 -1431
rect 481 -1432 482 -1404
rect 1297 -1529 1298 -1431
rect 1416 -1432 1417 -1404
rect 1444 -1529 1445 -1431
rect 114 -1529 115 -1433
rect 261 -1434 262 -1404
rect 324 -1434 325 -1404
rect 366 -1529 367 -1433
rect 436 -1529 437 -1433
rect 632 -1434 633 -1404
rect 660 -1529 661 -1433
rect 744 -1434 745 -1404
rect 768 -1529 769 -1433
rect 807 -1529 808 -1433
rect 880 -1529 881 -1433
rect 1325 -1434 1326 -1404
rect 1381 -1434 1382 -1404
rect 1416 -1529 1417 -1433
rect 135 -1436 136 -1404
rect 254 -1529 255 -1435
rect 261 -1529 262 -1435
rect 359 -1436 360 -1404
rect 541 -1529 542 -1435
rect 849 -1436 850 -1404
rect 884 -1436 885 -1404
rect 887 -1452 888 -1435
rect 919 -1436 920 -1404
rect 1507 -1436 1508 -1404
rect 79 -1438 80 -1404
rect 1507 -1529 1508 -1437
rect 135 -1529 136 -1439
rect 173 -1529 174 -1439
rect 184 -1529 185 -1439
rect 191 -1440 192 -1404
rect 205 -1440 206 -1404
rect 527 -1529 528 -1439
rect 555 -1440 556 -1404
rect 1164 -1529 1165 -1439
rect 1178 -1440 1179 -1404
rect 1332 -1529 1333 -1439
rect 1381 -1529 1382 -1439
rect 1409 -1440 1410 -1404
rect 72 -1442 73 -1404
rect 205 -1529 206 -1441
rect 219 -1442 220 -1404
rect 600 -1529 601 -1441
rect 688 -1529 689 -1441
rect 695 -1442 696 -1404
rect 744 -1529 745 -1441
rect 772 -1442 773 -1404
rect 803 -1529 804 -1441
rect 1045 -1529 1046 -1441
rect 1080 -1442 1081 -1404
rect 1206 -1529 1207 -1441
rect 1213 -1529 1214 -1441
rect 1220 -1442 1221 -1404
rect 1409 -1529 1410 -1441
rect 1458 -1442 1459 -1404
rect 72 -1529 73 -1443
rect 653 -1444 654 -1404
rect 772 -1529 773 -1443
rect 898 -1444 899 -1404
rect 905 -1444 906 -1404
rect 1080 -1529 1081 -1443
rect 1129 -1444 1130 -1404
rect 1325 -1529 1326 -1443
rect 191 -1529 192 -1445
rect 583 -1446 584 -1404
rect 653 -1529 654 -1445
rect 674 -1446 675 -1404
rect 849 -1529 850 -1445
rect 1038 -1446 1039 -1404
rect 1129 -1529 1130 -1445
rect 1255 -1446 1256 -1404
rect 219 -1529 220 -1447
rect 516 -1448 517 -1404
rect 583 -1529 584 -1447
rect 618 -1448 619 -1404
rect 859 -1529 860 -1447
rect 1458 -1529 1459 -1447
rect 233 -1450 234 -1404
rect 317 -1529 318 -1449
rect 324 -1529 325 -1449
rect 548 -1450 549 -1404
rect 884 -1529 885 -1449
rect 961 -1450 962 -1404
rect 975 -1450 976 -1404
rect 1514 -1450 1515 -1404
rect 177 -1452 178 -1404
rect 233 -1529 234 -1451
rect 240 -1452 241 -1404
rect 677 -1529 678 -1451
rect 961 -1529 962 -1451
rect 978 -1452 979 -1404
rect 1248 -1452 1249 -1404
rect 1514 -1529 1515 -1451
rect 1524 -1452 1525 -1404
rect 177 -1529 178 -1453
rect 590 -1454 591 -1404
rect 674 -1529 675 -1453
rect 1248 -1529 1249 -1453
rect 1437 -1454 1438 -1404
rect 1524 -1529 1525 -1453
rect 198 -1456 199 -1404
rect 548 -1529 549 -1455
rect 898 -1529 899 -1455
rect 954 -1456 955 -1404
rect 1006 -1456 1007 -1404
rect 1423 -1456 1424 -1404
rect 16 -1458 17 -1404
rect 198 -1529 199 -1457
rect 226 -1458 227 -1404
rect 590 -1529 591 -1457
rect 905 -1529 906 -1457
rect 940 -1458 941 -1404
rect 947 -1458 948 -1404
rect 1255 -1529 1256 -1457
rect 1388 -1458 1389 -1404
rect 1423 -1529 1424 -1457
rect 16 -1529 17 -1459
rect 30 -1460 31 -1404
rect 226 -1529 227 -1459
rect 345 -1460 346 -1404
rect 359 -1529 360 -1459
rect 443 -1460 444 -1404
rect 485 -1460 486 -1404
rect 555 -1529 556 -1459
rect 919 -1529 920 -1459
rect 968 -1460 969 -1404
rect 1017 -1460 1018 -1404
rect 1087 -1460 1088 -1404
rect 1136 -1460 1137 -1404
rect 1304 -1529 1305 -1459
rect 1374 -1460 1375 -1404
rect 1388 -1529 1389 -1459
rect 30 -1529 31 -1461
rect 506 -1462 507 -1404
rect 877 -1462 878 -1404
rect 968 -1529 969 -1461
rect 989 -1462 990 -1404
rect 1136 -1529 1137 -1461
rect 1150 -1462 1151 -1404
rect 1178 -1529 1179 -1461
rect 1220 -1529 1221 -1461
rect 1227 -1462 1228 -1404
rect 107 -1464 108 -1404
rect 506 -1529 507 -1463
rect 758 -1464 759 -1404
rect 877 -1529 878 -1463
rect 926 -1464 927 -1404
rect 975 -1529 976 -1463
rect 989 -1529 990 -1463
rect 1402 -1464 1403 -1404
rect 107 -1529 108 -1465
rect 163 -1466 164 -1404
rect 240 -1529 241 -1465
rect 457 -1466 458 -1404
rect 488 -1466 489 -1404
rect 1374 -1529 1375 -1465
rect 128 -1468 129 -1404
rect 163 -1529 164 -1467
rect 247 -1468 248 -1404
rect 845 -1468 846 -1404
rect 933 -1529 934 -1467
rect 999 -1529 1000 -1467
rect 1017 -1529 1018 -1467
rect 1073 -1468 1074 -1404
rect 1087 -1529 1088 -1467
rect 1094 -1468 1095 -1404
rect 1122 -1468 1123 -1404
rect 1227 -1529 1228 -1467
rect 128 -1529 129 -1469
rect 870 -1470 871 -1404
rect 940 -1529 941 -1469
rect 982 -1470 983 -1404
rect 1020 -1470 1021 -1404
rect 1493 -1470 1494 -1404
rect 79 -1529 80 -1471
rect 870 -1529 871 -1471
rect 947 -1529 948 -1471
rect 1066 -1472 1067 -1404
rect 1094 -1529 1095 -1471
rect 1108 -1472 1109 -1404
rect 1150 -1529 1151 -1471
rect 1290 -1472 1291 -1404
rect 1486 -1472 1487 -1404
rect 1493 -1529 1494 -1471
rect 247 -1529 248 -1473
rect 289 -1474 290 -1404
rect 331 -1474 332 -1404
rect 618 -1529 619 -1473
rect 632 -1529 633 -1473
rect 1122 -1529 1123 -1473
rect 1283 -1474 1284 -1404
rect 1290 -1529 1291 -1473
rect 1479 -1474 1480 -1404
rect 1486 -1529 1487 -1473
rect 282 -1476 283 -1404
rect 289 -1529 290 -1475
rect 331 -1529 332 -1475
rect 422 -1476 423 -1404
rect 443 -1529 444 -1475
rect 579 -1529 580 -1475
rect 695 -1529 696 -1475
rect 1073 -1529 1074 -1475
rect 1283 -1529 1284 -1475
rect 1500 -1476 1501 -1404
rect 282 -1529 283 -1477
rect 303 -1478 304 -1404
rect 345 -1529 346 -1477
rect 499 -1529 500 -1477
rect 502 -1529 503 -1477
rect 926 -1529 927 -1477
rect 954 -1529 955 -1477
rect 1010 -1478 1011 -1404
rect 1024 -1478 1025 -1404
rect 1066 -1529 1067 -1477
rect 1472 -1478 1473 -1404
rect 1500 -1529 1501 -1477
rect 303 -1529 304 -1479
rect 310 -1480 311 -1404
rect 352 -1480 353 -1404
rect 457 -1529 458 -1479
rect 709 -1480 710 -1404
rect 1479 -1529 1480 -1479
rect 9 -1482 10 -1404
rect 352 -1529 353 -1481
rect 387 -1482 388 -1404
rect 422 -1529 423 -1481
rect 450 -1482 451 -1404
rect 485 -1529 486 -1481
rect 716 -1482 717 -1404
rect 1402 -1529 1403 -1481
rect 1451 -1482 1452 -1404
rect 1472 -1529 1473 -1481
rect 9 -1529 10 -1483
rect 681 -1484 682 -1404
rect 758 -1529 759 -1483
rect 765 -1484 766 -1404
rect 982 -1529 983 -1483
rect 996 -1484 997 -1404
rect 1010 -1529 1011 -1483
rect 1059 -1484 1060 -1404
rect 1430 -1484 1431 -1404
rect 1451 -1529 1452 -1483
rect 54 -1529 55 -1485
rect 709 -1529 710 -1485
rect 765 -1529 766 -1485
rect 922 -1486 923 -1404
rect 1024 -1529 1025 -1485
rect 1052 -1486 1053 -1404
rect 1059 -1529 1060 -1485
rect 1171 -1486 1172 -1404
rect 1395 -1486 1396 -1404
rect 1430 -1529 1431 -1485
rect 58 -1488 59 -1404
rect 716 -1529 717 -1487
rect 751 -1488 752 -1404
rect 1052 -1529 1053 -1487
rect 1367 -1488 1368 -1404
rect 1395 -1529 1396 -1487
rect 58 -1529 59 -1489
rect 814 -1490 815 -1404
rect 1031 -1490 1032 -1404
rect 1115 -1529 1116 -1489
rect 212 -1492 213 -1404
rect 450 -1529 451 -1491
rect 471 -1529 472 -1491
rect 1171 -1529 1172 -1491
rect 149 -1494 150 -1404
rect 212 -1529 213 -1493
rect 310 -1529 311 -1493
rect 474 -1529 475 -1493
rect 751 -1529 752 -1493
rect 821 -1494 822 -1404
rect 1031 -1529 1032 -1493
rect 1157 -1494 1158 -1404
rect 149 -1529 150 -1495
rect 170 -1496 171 -1404
rect 387 -1529 388 -1495
rect 429 -1496 430 -1404
rect 681 -1529 682 -1495
rect 1157 -1529 1158 -1495
rect 401 -1498 402 -1404
rect 1108 -1529 1109 -1497
rect 2 -1500 3 -1404
rect 401 -1529 402 -1499
rect 415 -1500 416 -1404
rect 1367 -1529 1368 -1499
rect 2 -1529 3 -1501
rect 142 -1502 143 -1404
rect 373 -1502 374 -1404
rect 415 -1529 416 -1501
rect 429 -1529 430 -1501
rect 891 -1502 892 -1404
rect 1038 -1529 1039 -1501
rect 1185 -1502 1186 -1404
rect 142 -1529 143 -1503
rect 156 -1504 157 -1404
rect 373 -1529 374 -1503
rect 380 -1504 381 -1404
rect 814 -1529 815 -1503
rect 1339 -1504 1340 -1404
rect 86 -1506 87 -1404
rect 380 -1529 381 -1505
rect 821 -1529 822 -1505
rect 863 -1506 864 -1404
rect 891 -1529 892 -1505
rect 912 -1506 913 -1404
rect 1101 -1506 1102 -1404
rect 1185 -1529 1186 -1505
rect 86 -1529 87 -1507
rect 604 -1508 605 -1404
rect 639 -1508 640 -1404
rect 863 -1529 864 -1507
rect 1101 -1529 1102 -1507
rect 1199 -1508 1200 -1404
rect 110 -1510 111 -1404
rect 1339 -1529 1340 -1509
rect 156 -1529 157 -1511
rect 576 -1512 577 -1404
rect 604 -1529 605 -1511
rect 625 -1512 626 -1404
rect 639 -1529 640 -1511
rect 667 -1512 668 -1404
rect 786 -1512 787 -1404
rect 912 -1529 913 -1511
rect 534 -1514 535 -1404
rect 667 -1529 668 -1513
rect 786 -1529 787 -1513
rect 828 -1514 829 -1404
rect 534 -1529 535 -1515
rect 597 -1516 598 -1404
rect 611 -1516 612 -1404
rect 625 -1529 626 -1515
rect 817 -1529 818 -1515
rect 1199 -1529 1200 -1515
rect 576 -1529 577 -1517
rect 1125 -1529 1126 -1517
rect 597 -1529 598 -1519
rect 1437 -1529 1438 -1519
rect 611 -1529 612 -1521
rect 702 -1522 703 -1404
rect 828 -1529 829 -1521
rect 1318 -1529 1319 -1521
rect 702 -1529 703 -1523
rect 737 -1524 738 -1404
rect 737 -1529 738 -1525
rect 793 -1526 794 -1404
rect 394 -1529 395 -1527
rect 793 -1529 794 -1527
rect 2 -1539 3 -1537
rect 131 -1636 132 -1538
rect 142 -1539 143 -1537
rect 173 -1539 174 -1537
rect 212 -1539 213 -1537
rect 432 -1539 433 -1537
rect 471 -1539 472 -1537
rect 667 -1539 668 -1537
rect 674 -1539 675 -1537
rect 1325 -1539 1326 -1537
rect 1349 -1636 1350 -1538
rect 1535 -1539 1536 -1537
rect 2 -1636 3 -1540
rect 275 -1541 276 -1537
rect 303 -1541 304 -1537
rect 303 -1636 304 -1540
rect 303 -1541 304 -1537
rect 303 -1636 304 -1540
rect 345 -1541 346 -1537
rect 856 -1636 857 -1540
rect 859 -1541 860 -1537
rect 1514 -1541 1515 -1537
rect 9 -1543 10 -1537
rect 12 -1601 13 -1542
rect 16 -1543 17 -1537
rect 16 -1636 17 -1542
rect 16 -1543 17 -1537
rect 16 -1636 17 -1542
rect 23 -1543 24 -1537
rect 23 -1636 24 -1542
rect 23 -1543 24 -1537
rect 23 -1636 24 -1542
rect 30 -1543 31 -1537
rect 446 -1636 447 -1542
rect 474 -1543 475 -1537
rect 817 -1543 818 -1537
rect 838 -1543 839 -1537
rect 1220 -1543 1221 -1537
rect 1325 -1636 1326 -1542
rect 1395 -1543 1396 -1537
rect 9 -1636 10 -1544
rect 485 -1545 486 -1537
rect 502 -1545 503 -1537
rect 625 -1545 626 -1537
rect 639 -1545 640 -1537
rect 754 -1636 755 -1544
rect 758 -1545 759 -1537
rect 768 -1545 769 -1537
rect 782 -1636 783 -1544
rect 849 -1545 850 -1537
rect 880 -1636 881 -1544
rect 1185 -1545 1186 -1537
rect 1220 -1636 1221 -1544
rect 1297 -1545 1298 -1537
rect 30 -1636 31 -1546
rect 135 -1547 136 -1537
rect 142 -1636 143 -1546
rect 632 -1547 633 -1537
rect 639 -1636 640 -1546
rect 653 -1547 654 -1537
rect 667 -1636 668 -1546
rect 807 -1547 808 -1537
rect 849 -1636 850 -1546
rect 863 -1547 864 -1537
rect 947 -1547 948 -1537
rect 950 -1601 951 -1546
rect 992 -1547 993 -1537
rect 1332 -1547 1333 -1537
rect 44 -1549 45 -1537
rect 275 -1636 276 -1548
rect 366 -1549 367 -1537
rect 632 -1636 633 -1548
rect 653 -1636 654 -1548
rect 716 -1549 717 -1537
rect 765 -1549 766 -1537
rect 1171 -1549 1172 -1537
rect 1185 -1636 1186 -1548
rect 1248 -1549 1249 -1537
rect 1297 -1636 1298 -1548
rect 1374 -1549 1375 -1537
rect 44 -1636 45 -1550
rect 611 -1551 612 -1537
rect 618 -1551 619 -1537
rect 674 -1636 675 -1550
rect 677 -1551 678 -1537
rect 1521 -1551 1522 -1537
rect 51 -1553 52 -1537
rect 107 -1553 108 -1537
rect 128 -1553 129 -1537
rect 212 -1636 213 -1552
rect 397 -1553 398 -1537
rect 1402 -1553 1403 -1537
rect 51 -1636 52 -1554
rect 562 -1555 563 -1537
rect 579 -1555 580 -1537
rect 730 -1555 731 -1537
rect 765 -1636 766 -1554
rect 957 -1636 958 -1554
rect 996 -1555 997 -1537
rect 1115 -1555 1116 -1537
rect 1122 -1555 1123 -1537
rect 1409 -1555 1410 -1537
rect 54 -1557 55 -1537
rect 772 -1557 773 -1537
rect 863 -1636 864 -1556
rect 919 -1557 920 -1537
rect 947 -1636 948 -1556
rect 1003 -1557 1004 -1537
rect 1010 -1557 1011 -1537
rect 1010 -1636 1011 -1556
rect 1010 -1557 1011 -1537
rect 1010 -1636 1011 -1556
rect 1073 -1557 1074 -1537
rect 1500 -1557 1501 -1537
rect 65 -1559 66 -1537
rect 502 -1636 503 -1558
rect 506 -1559 507 -1537
rect 807 -1636 808 -1558
rect 919 -1636 920 -1558
rect 982 -1559 983 -1537
rect 992 -1636 993 -1558
rect 1073 -1636 1074 -1558
rect 1115 -1636 1116 -1558
rect 1143 -1559 1144 -1537
rect 1150 -1559 1151 -1537
rect 1153 -1559 1154 -1537
rect 1171 -1636 1172 -1558
rect 1234 -1559 1235 -1537
rect 1374 -1636 1375 -1558
rect 1451 -1559 1452 -1537
rect 65 -1636 66 -1560
rect 72 -1561 73 -1537
rect 75 -1636 76 -1560
rect 527 -1561 528 -1537
rect 534 -1561 535 -1537
rect 534 -1636 535 -1560
rect 534 -1561 535 -1537
rect 534 -1636 535 -1560
rect 583 -1561 584 -1537
rect 649 -1636 650 -1560
rect 681 -1561 682 -1537
rect 1080 -1561 1081 -1537
rect 1101 -1561 1102 -1537
rect 1143 -1636 1144 -1560
rect 1150 -1636 1151 -1560
rect 1199 -1561 1200 -1537
rect 1234 -1636 1235 -1560
rect 1416 -1561 1417 -1537
rect 1451 -1636 1452 -1560
rect 1528 -1561 1529 -1537
rect 58 -1563 59 -1537
rect 527 -1636 528 -1562
rect 583 -1636 584 -1562
rect 590 -1563 591 -1537
rect 600 -1563 601 -1537
rect 751 -1563 752 -1537
rect 800 -1563 801 -1537
rect 1080 -1636 1081 -1562
rect 1101 -1636 1102 -1562
rect 1108 -1563 1109 -1537
rect 1192 -1563 1193 -1537
rect 1248 -1636 1249 -1562
rect 1283 -1563 1284 -1537
rect 1416 -1636 1417 -1562
rect 58 -1636 59 -1564
rect 373 -1565 374 -1537
rect 394 -1565 395 -1537
rect 1409 -1636 1410 -1564
rect 72 -1636 73 -1566
rect 254 -1567 255 -1537
rect 373 -1636 374 -1566
rect 457 -1567 458 -1537
rect 478 -1567 479 -1537
rect 831 -1567 832 -1537
rect 982 -1636 983 -1566
rect 1017 -1567 1018 -1537
rect 1059 -1567 1060 -1537
rect 1108 -1636 1109 -1566
rect 1192 -1636 1193 -1566
rect 1269 -1567 1270 -1537
rect 1283 -1636 1284 -1566
rect 1311 -1567 1312 -1537
rect 1402 -1636 1403 -1566
rect 1479 -1567 1480 -1537
rect 79 -1636 80 -1568
rect 114 -1569 115 -1537
rect 135 -1636 136 -1568
rect 723 -1569 724 -1537
rect 730 -1636 731 -1568
rect 793 -1569 794 -1537
rect 800 -1636 801 -1568
rect 842 -1569 843 -1537
rect 989 -1569 990 -1537
rect 1017 -1636 1018 -1568
rect 1024 -1569 1025 -1537
rect 1269 -1636 1270 -1568
rect 1311 -1636 1312 -1568
rect 1458 -1569 1459 -1537
rect 82 -1571 83 -1537
rect 492 -1571 493 -1537
rect 506 -1636 507 -1570
rect 870 -1571 871 -1537
rect 898 -1571 899 -1537
rect 1024 -1636 1025 -1570
rect 1059 -1636 1060 -1570
rect 1395 -1636 1396 -1570
rect 103 -1573 104 -1537
rect 226 -1573 227 -1537
rect 380 -1573 381 -1537
rect 478 -1636 479 -1572
rect 492 -1636 493 -1572
rect 520 -1573 521 -1537
rect 590 -1636 591 -1572
rect 702 -1573 703 -1537
rect 716 -1636 717 -1572
rect 737 -1573 738 -1537
rect 751 -1636 752 -1572
rect 1031 -1573 1032 -1537
rect 107 -1636 108 -1574
rect 338 -1575 339 -1537
rect 348 -1636 349 -1574
rect 380 -1636 381 -1574
rect 394 -1636 395 -1574
rect 555 -1575 556 -1537
rect 611 -1636 612 -1574
rect 660 -1575 661 -1537
rect 681 -1636 682 -1574
rect 695 -1575 696 -1537
rect 702 -1636 703 -1574
rect 786 -1575 787 -1537
rect 793 -1636 794 -1574
rect 1524 -1575 1525 -1537
rect 114 -1636 115 -1576
rect 261 -1577 262 -1537
rect 338 -1636 339 -1576
rect 726 -1577 727 -1537
rect 737 -1636 738 -1576
rect 1262 -1577 1263 -1537
rect 145 -1636 146 -1578
rect 744 -1579 745 -1537
rect 786 -1636 787 -1578
rect 814 -1579 815 -1537
rect 870 -1636 871 -1578
rect 926 -1579 927 -1537
rect 933 -1579 934 -1537
rect 1031 -1636 1032 -1578
rect 1262 -1636 1263 -1578
rect 1339 -1579 1340 -1537
rect 128 -1636 129 -1580
rect 933 -1636 934 -1580
rect 996 -1636 997 -1580
rect 1076 -1581 1077 -1537
rect 1255 -1581 1256 -1537
rect 1339 -1636 1340 -1580
rect 149 -1583 150 -1537
rect 149 -1636 150 -1582
rect 149 -1583 150 -1537
rect 149 -1636 150 -1582
rect 156 -1583 157 -1537
rect 625 -1636 626 -1582
rect 646 -1583 647 -1537
rect 831 -1636 832 -1582
rect 898 -1636 899 -1582
rect 975 -1583 976 -1537
rect 999 -1583 1000 -1537
rect 1129 -1583 1130 -1537
rect 156 -1636 157 -1584
rect 271 -1636 272 -1584
rect 408 -1585 409 -1537
rect 772 -1636 773 -1584
rect 814 -1636 815 -1584
rect 884 -1585 885 -1537
rect 975 -1636 976 -1584
rect 1038 -1585 1039 -1537
rect 1045 -1585 1046 -1537
rect 1255 -1636 1256 -1584
rect 163 -1587 164 -1537
rect 842 -1636 843 -1586
rect 884 -1636 885 -1586
rect 961 -1587 962 -1537
rect 1038 -1636 1039 -1586
rect 1087 -1587 1088 -1537
rect 1129 -1636 1130 -1586
rect 1157 -1587 1158 -1537
rect 163 -1636 164 -1588
rect 401 -1589 402 -1537
rect 429 -1636 430 -1588
rect 464 -1589 465 -1537
rect 474 -1636 475 -1588
rect 520 -1636 521 -1588
rect 555 -1636 556 -1588
rect 1367 -1589 1368 -1537
rect 170 -1591 171 -1537
rect 439 -1636 440 -1590
rect 450 -1591 451 -1537
rect 758 -1636 759 -1590
rect 817 -1636 818 -1590
rect 926 -1636 927 -1590
rect 1045 -1636 1046 -1590
rect 1094 -1591 1095 -1537
rect 1157 -1636 1158 -1590
rect 1213 -1591 1214 -1537
rect 1367 -1636 1368 -1590
rect 1444 -1591 1445 -1537
rect 170 -1636 171 -1592
rect 205 -1593 206 -1537
rect 261 -1636 262 -1592
rect 310 -1593 311 -1537
rect 352 -1593 353 -1537
rect 401 -1636 402 -1592
rect 415 -1593 416 -1537
rect 464 -1636 465 -1592
rect 499 -1593 500 -1537
rect 961 -1636 962 -1592
rect 1094 -1636 1095 -1592
rect 1276 -1593 1277 -1537
rect 100 -1595 101 -1537
rect 205 -1636 206 -1594
rect 240 -1595 241 -1537
rect 310 -1636 311 -1594
rect 331 -1595 332 -1537
rect 415 -1636 416 -1594
rect 450 -1636 451 -1594
rect 803 -1595 804 -1537
rect 1213 -1636 1214 -1594
rect 1430 -1595 1431 -1537
rect 100 -1636 101 -1596
rect 121 -1597 122 -1537
rect 177 -1597 178 -1537
rect 485 -1636 486 -1596
rect 499 -1636 500 -1596
rect 1332 -1636 1333 -1596
rect 93 -1599 94 -1537
rect 121 -1636 122 -1598
rect 177 -1636 178 -1598
rect 621 -1636 622 -1598
rect 912 -1599 913 -1537
rect 1052 -1599 1053 -1537
rect 1430 -1636 1431 -1598
rect 93 -1636 94 -1600
rect 219 -1601 220 -1537
rect 240 -1636 241 -1600
rect 387 -1601 388 -1537
rect 457 -1636 458 -1600
rect 513 -1601 514 -1537
rect 646 -1636 647 -1600
rect 1136 -1601 1137 -1537
rect 1153 -1636 1154 -1600
rect 1199 -1636 1200 -1600
rect 1276 -1636 1277 -1600
rect 1346 -1601 1347 -1537
rect 86 -1603 87 -1537
rect 513 -1636 514 -1602
rect 660 -1636 661 -1602
rect 688 -1603 689 -1537
rect 695 -1636 696 -1602
rect 779 -1603 780 -1537
rect 912 -1636 913 -1602
rect 968 -1603 969 -1537
rect 989 -1636 990 -1602
rect 1346 -1636 1347 -1602
rect 86 -1636 87 -1604
rect 282 -1605 283 -1537
rect 296 -1605 297 -1537
rect 352 -1636 353 -1604
rect 369 -1636 370 -1604
rect 387 -1636 388 -1604
rect 471 -1636 472 -1604
rect 688 -1636 689 -1604
rect 723 -1636 724 -1604
rect 821 -1605 822 -1537
rect 968 -1636 969 -1604
rect 1164 -1605 1165 -1537
rect 184 -1607 185 -1537
rect 366 -1636 367 -1606
rect 684 -1607 685 -1537
rect 1507 -1607 1508 -1537
rect 184 -1636 185 -1608
rect 233 -1609 234 -1537
rect 282 -1636 283 -1608
rect 289 -1609 290 -1537
rect 331 -1636 332 -1608
rect 565 -1636 566 -1608
rect 740 -1636 741 -1608
rect 1087 -1636 1088 -1608
rect 1136 -1636 1137 -1608
rect 1178 -1609 1179 -1537
rect 191 -1611 192 -1537
rect 408 -1636 409 -1610
rect 744 -1636 745 -1610
rect 835 -1611 836 -1537
rect 1052 -1636 1053 -1610
rect 1318 -1611 1319 -1537
rect 191 -1636 192 -1612
rect 618 -1636 619 -1612
rect 709 -1613 710 -1537
rect 1318 -1636 1319 -1612
rect 198 -1615 199 -1537
rect 254 -1636 255 -1614
rect 289 -1636 290 -1614
rect 359 -1615 360 -1537
rect 548 -1615 549 -1537
rect 709 -1636 710 -1614
rect 779 -1636 780 -1614
rect 1066 -1615 1067 -1537
rect 1164 -1636 1165 -1614
rect 1227 -1615 1228 -1537
rect 198 -1636 199 -1616
rect 268 -1617 269 -1537
rect 359 -1636 360 -1616
rect 576 -1617 577 -1537
rect 821 -1636 822 -1616
rect 828 -1617 829 -1537
rect 835 -1636 836 -1616
rect 891 -1617 892 -1537
rect 905 -1617 906 -1537
rect 1066 -1636 1067 -1616
rect 1178 -1636 1179 -1616
rect 1241 -1617 1242 -1537
rect 219 -1636 220 -1618
rect 247 -1619 248 -1537
rect 541 -1619 542 -1537
rect 576 -1636 577 -1618
rect 828 -1636 829 -1618
rect 1122 -1636 1123 -1618
rect 1227 -1636 1228 -1618
rect 1353 -1619 1354 -1537
rect 226 -1636 227 -1620
rect 268 -1636 269 -1620
rect 422 -1621 423 -1537
rect 541 -1636 542 -1620
rect 548 -1636 549 -1620
rect 604 -1621 605 -1537
rect 891 -1636 892 -1620
rect 954 -1621 955 -1537
rect 1241 -1636 1242 -1620
rect 1304 -1621 1305 -1537
rect 1353 -1636 1354 -1620
rect 1381 -1621 1382 -1537
rect 233 -1636 234 -1622
rect 558 -1636 559 -1622
rect 569 -1623 570 -1537
rect 604 -1636 605 -1622
rect 905 -1636 906 -1622
rect 940 -1623 941 -1537
rect 954 -1636 955 -1622
rect 1360 -1623 1361 -1537
rect 1381 -1636 1382 -1622
rect 1465 -1623 1466 -1537
rect 247 -1636 248 -1624
rect 443 -1625 444 -1537
rect 877 -1625 878 -1537
rect 940 -1636 941 -1624
rect 1304 -1636 1305 -1624
rect 1388 -1625 1389 -1537
rect 296 -1636 297 -1626
rect 443 -1636 444 -1626
rect 877 -1636 878 -1626
rect 1206 -1627 1207 -1537
rect 1360 -1636 1361 -1626
rect 1437 -1627 1438 -1537
rect 324 -1629 325 -1537
rect 422 -1636 423 -1628
rect 436 -1629 437 -1537
rect 569 -1636 570 -1628
rect 1206 -1636 1207 -1628
rect 1290 -1629 1291 -1537
rect 1388 -1636 1389 -1628
rect 1472 -1629 1473 -1537
rect 317 -1631 318 -1537
rect 324 -1636 325 -1630
rect 1290 -1636 1291 -1630
rect 1423 -1631 1424 -1537
rect 1437 -1636 1438 -1630
rect 1486 -1631 1487 -1537
rect 37 -1633 38 -1537
rect 317 -1636 318 -1632
rect 1423 -1636 1424 -1632
rect 1493 -1633 1494 -1537
rect 37 -1636 38 -1634
rect 562 -1636 563 -1634
rect 2 -1646 3 -1644
rect 436 -1646 437 -1644
rect 446 -1646 447 -1644
rect 474 -1646 475 -1644
rect 488 -1761 489 -1645
rect 1206 -1646 1207 -1644
rect 1283 -1646 1284 -1644
rect 1346 -1646 1347 -1644
rect 1377 -1761 1378 -1645
rect 1451 -1646 1452 -1644
rect 23 -1648 24 -1644
rect 23 -1761 24 -1647
rect 23 -1648 24 -1644
rect 23 -1761 24 -1647
rect 37 -1648 38 -1644
rect 341 -1761 342 -1647
rect 429 -1648 430 -1644
rect 443 -1761 444 -1647
rect 471 -1648 472 -1644
rect 597 -1648 598 -1644
rect 621 -1648 622 -1644
rect 765 -1648 766 -1644
rect 800 -1648 801 -1644
rect 800 -1761 801 -1647
rect 800 -1648 801 -1644
rect 800 -1761 801 -1647
rect 814 -1761 815 -1647
rect 1017 -1648 1018 -1644
rect 1206 -1761 1207 -1647
rect 1297 -1648 1298 -1644
rect 37 -1761 38 -1649
rect 387 -1650 388 -1644
rect 429 -1761 430 -1649
rect 520 -1650 521 -1644
rect 555 -1650 556 -1644
rect 667 -1650 668 -1644
rect 709 -1650 710 -1644
rect 873 -1761 874 -1649
rect 877 -1650 878 -1644
rect 1003 -1650 1004 -1644
rect 1017 -1761 1018 -1649
rect 1150 -1650 1151 -1644
rect 1283 -1761 1284 -1649
rect 1367 -1650 1368 -1644
rect 51 -1652 52 -1644
rect 51 -1761 52 -1651
rect 51 -1652 52 -1644
rect 51 -1761 52 -1651
rect 65 -1652 66 -1644
rect 586 -1761 587 -1651
rect 597 -1761 598 -1651
rect 863 -1652 864 -1644
rect 877 -1761 878 -1651
rect 1297 -1761 1298 -1651
rect 1367 -1761 1368 -1651
rect 1430 -1652 1431 -1644
rect 65 -1761 66 -1653
rect 149 -1654 150 -1644
rect 163 -1654 164 -1644
rect 418 -1761 419 -1653
rect 436 -1761 437 -1653
rect 782 -1654 783 -1644
rect 828 -1654 829 -1644
rect 1094 -1654 1095 -1644
rect 1150 -1761 1151 -1653
rect 1199 -1654 1200 -1644
rect 72 -1656 73 -1644
rect 506 -1656 507 -1644
rect 513 -1656 514 -1644
rect 740 -1656 741 -1644
rect 744 -1656 745 -1644
rect 775 -1761 776 -1655
rect 817 -1656 818 -1644
rect 1199 -1761 1200 -1655
rect 82 -1761 83 -1657
rect 625 -1658 626 -1644
rect 635 -1761 636 -1657
rect 786 -1658 787 -1644
rect 828 -1761 829 -1657
rect 933 -1658 934 -1644
rect 1094 -1761 1095 -1657
rect 1304 -1658 1305 -1644
rect 128 -1660 129 -1644
rect 632 -1660 633 -1644
rect 653 -1660 654 -1644
rect 656 -1676 657 -1659
rect 667 -1761 668 -1659
rect 674 -1660 675 -1644
rect 709 -1761 710 -1659
rect 716 -1660 717 -1644
rect 719 -1761 720 -1659
rect 968 -1660 969 -1644
rect 1006 -1761 1007 -1659
rect 1304 -1761 1305 -1659
rect 128 -1761 129 -1661
rect 135 -1662 136 -1644
rect 149 -1761 150 -1661
rect 233 -1662 234 -1644
rect 240 -1662 241 -1644
rect 369 -1662 370 -1644
rect 387 -1761 388 -1661
rect 492 -1662 493 -1644
rect 513 -1761 514 -1661
rect 523 -1761 524 -1661
rect 555 -1761 556 -1661
rect 590 -1662 591 -1644
rect 604 -1662 605 -1644
rect 674 -1761 675 -1661
rect 723 -1662 724 -1644
rect 880 -1662 881 -1644
rect 933 -1761 934 -1661
rect 1080 -1662 1081 -1644
rect 9 -1664 10 -1644
rect 369 -1761 370 -1663
rect 471 -1761 472 -1663
rect 737 -1664 738 -1644
rect 751 -1664 752 -1644
rect 1346 -1761 1347 -1663
rect 9 -1761 10 -1665
rect 93 -1666 94 -1644
rect 121 -1666 122 -1644
rect 135 -1761 136 -1665
rect 142 -1666 143 -1644
rect 233 -1761 234 -1665
rect 240 -1761 241 -1665
rect 254 -1666 255 -1644
rect 303 -1666 304 -1644
rect 345 -1666 346 -1644
rect 359 -1666 360 -1644
rect 632 -1761 633 -1665
rect 653 -1761 654 -1665
rect 688 -1666 689 -1644
rect 751 -1761 752 -1665
rect 821 -1666 822 -1644
rect 863 -1761 864 -1665
rect 891 -1666 892 -1644
rect 968 -1761 969 -1665
rect 1038 -1666 1039 -1644
rect 1080 -1761 1081 -1665
rect 1185 -1666 1186 -1644
rect 93 -1761 94 -1667
rect 548 -1668 549 -1644
rect 562 -1668 563 -1644
rect 1255 -1668 1256 -1644
rect 114 -1670 115 -1644
rect 303 -1761 304 -1669
rect 310 -1670 311 -1644
rect 520 -1761 521 -1669
rect 527 -1670 528 -1644
rect 562 -1761 563 -1669
rect 565 -1670 566 -1644
rect 807 -1670 808 -1644
rect 821 -1761 822 -1669
rect 884 -1670 885 -1644
rect 891 -1761 892 -1669
rect 947 -1670 948 -1644
rect 1038 -1761 1039 -1669
rect 1143 -1670 1144 -1644
rect 1255 -1761 1256 -1669
rect 1290 -1670 1291 -1644
rect 79 -1672 80 -1644
rect 114 -1761 115 -1671
rect 121 -1761 122 -1671
rect 156 -1672 157 -1644
rect 163 -1761 164 -1671
rect 184 -1672 185 -1644
rect 198 -1672 199 -1644
rect 271 -1672 272 -1644
rect 310 -1761 311 -1671
rect 401 -1672 402 -1644
rect 408 -1672 409 -1644
rect 548 -1761 549 -1671
rect 590 -1761 591 -1671
rect 660 -1672 661 -1644
rect 758 -1672 759 -1644
rect 831 -1672 832 -1644
rect 845 -1761 846 -1671
rect 1185 -1761 1186 -1671
rect 1290 -1761 1291 -1671
rect 1374 -1672 1375 -1644
rect 58 -1674 59 -1644
rect 156 -1761 157 -1673
rect 177 -1674 178 -1644
rect 499 -1674 500 -1644
rect 604 -1761 605 -1673
rect 779 -1674 780 -1644
rect 786 -1761 787 -1673
rect 989 -1761 990 -1673
rect 58 -1761 59 -1675
rect 541 -1676 542 -1644
rect 625 -1761 626 -1675
rect 639 -1676 640 -1644
rect 688 -1761 689 -1675
rect 758 -1761 759 -1675
rect 1031 -1676 1032 -1644
rect 79 -1761 80 -1677
rect 324 -1678 325 -1644
rect 345 -1761 346 -1677
rect 415 -1678 416 -1644
rect 485 -1678 486 -1644
rect 737 -1761 738 -1677
rect 765 -1761 766 -1677
rect 961 -1678 962 -1644
rect 1031 -1761 1032 -1677
rect 1157 -1678 1158 -1644
rect 110 -1680 111 -1644
rect 408 -1761 409 -1679
rect 492 -1761 493 -1679
rect 649 -1680 650 -1644
rect 660 -1761 661 -1679
rect 730 -1680 731 -1644
rect 779 -1761 780 -1679
rect 835 -1680 836 -1644
rect 880 -1761 881 -1679
rect 1010 -1680 1011 -1644
rect 1157 -1761 1158 -1679
rect 1241 -1680 1242 -1644
rect 110 -1761 111 -1681
rect 842 -1682 843 -1644
rect 884 -1761 885 -1681
rect 905 -1682 906 -1644
rect 926 -1682 927 -1644
rect 1143 -1761 1144 -1681
rect 142 -1761 143 -1683
rect 695 -1684 696 -1644
rect 730 -1761 731 -1683
rect 849 -1684 850 -1644
rect 905 -1761 906 -1683
rect 1349 -1684 1350 -1644
rect 177 -1761 178 -1685
rect 754 -1686 755 -1644
rect 835 -1761 836 -1685
rect 870 -1686 871 -1644
rect 926 -1761 927 -1685
rect 1101 -1686 1102 -1644
rect 184 -1761 185 -1687
rect 425 -1761 426 -1687
rect 506 -1761 507 -1687
rect 1241 -1761 1242 -1687
rect 198 -1761 199 -1689
rect 954 -1690 955 -1644
rect 961 -1761 962 -1689
rect 982 -1690 983 -1644
rect 1010 -1761 1011 -1689
rect 1171 -1690 1172 -1644
rect 205 -1692 206 -1644
rect 527 -1761 528 -1691
rect 576 -1692 577 -1644
rect 695 -1761 696 -1691
rect 842 -1761 843 -1691
rect 1227 -1692 1228 -1644
rect 205 -1761 206 -1693
rect 261 -1694 262 -1644
rect 268 -1694 269 -1644
rect 499 -1761 500 -1693
rect 576 -1761 577 -1693
rect 1003 -1761 1004 -1693
rect 1101 -1761 1102 -1693
rect 1220 -1694 1221 -1644
rect 1227 -1761 1228 -1693
rect 1409 -1694 1410 -1644
rect 219 -1696 220 -1644
rect 261 -1761 262 -1695
rect 268 -1761 269 -1695
rect 317 -1696 318 -1644
rect 359 -1761 360 -1695
rect 464 -1696 465 -1644
rect 611 -1696 612 -1644
rect 639 -1761 640 -1695
rect 849 -1761 850 -1695
rect 919 -1696 920 -1644
rect 947 -1761 948 -1695
rect 1045 -1696 1046 -1644
rect 1220 -1761 1221 -1695
rect 1318 -1696 1319 -1644
rect 219 -1761 220 -1697
rect 796 -1761 797 -1697
rect 870 -1761 871 -1697
rect 1234 -1698 1235 -1644
rect 1248 -1698 1249 -1644
rect 1318 -1761 1319 -1697
rect 254 -1761 255 -1699
rect 415 -1761 416 -1699
rect 464 -1761 465 -1699
rect 478 -1700 479 -1644
rect 611 -1761 612 -1699
rect 856 -1700 857 -1644
rect 901 -1761 902 -1699
rect 1248 -1761 1249 -1699
rect 289 -1702 290 -1644
rect 317 -1761 318 -1701
rect 366 -1702 367 -1644
rect 744 -1761 745 -1701
rect 856 -1761 857 -1701
rect 898 -1702 899 -1644
rect 919 -1761 920 -1701
rect 1087 -1702 1088 -1644
rect 1234 -1761 1235 -1701
rect 1388 -1702 1389 -1644
rect 212 -1704 213 -1644
rect 366 -1761 367 -1703
rect 394 -1704 395 -1644
rect 541 -1761 542 -1703
rect 898 -1761 899 -1703
rect 940 -1704 941 -1644
rect 954 -1761 955 -1703
rect 1129 -1704 1130 -1644
rect 131 -1706 132 -1644
rect 1129 -1761 1130 -1705
rect 212 -1761 213 -1707
rect 275 -1708 276 -1644
rect 282 -1708 283 -1644
rect 289 -1761 290 -1707
rect 296 -1708 297 -1644
rect 324 -1761 325 -1707
rect 394 -1761 395 -1707
rect 422 -1708 423 -1644
rect 478 -1761 479 -1707
rect 534 -1708 535 -1644
rect 940 -1761 941 -1707
rect 975 -1708 976 -1644
rect 982 -1761 983 -1707
rect 1073 -1708 1074 -1644
rect 1087 -1761 1088 -1707
rect 1192 -1708 1193 -1644
rect 75 -1710 76 -1644
rect 296 -1761 297 -1709
rect 401 -1761 402 -1709
rect 569 -1710 570 -1644
rect 975 -1761 976 -1709
rect 1122 -1710 1123 -1644
rect 1192 -1761 1193 -1709
rect 1262 -1710 1263 -1644
rect 75 -1761 76 -1711
rect 723 -1761 724 -1711
rect 996 -1712 997 -1644
rect 1171 -1761 1172 -1711
rect 1262 -1761 1263 -1711
rect 1332 -1712 1333 -1644
rect 107 -1714 108 -1644
rect 275 -1761 276 -1713
rect 282 -1761 283 -1713
rect 373 -1714 374 -1644
rect 380 -1714 381 -1644
rect 569 -1761 570 -1713
rect 996 -1761 997 -1713
rect 1108 -1714 1109 -1644
rect 1332 -1761 1333 -1713
rect 1402 -1714 1403 -1644
rect 72 -1761 73 -1715
rect 380 -1761 381 -1715
rect 422 -1761 423 -1715
rect 583 -1716 584 -1644
rect 1024 -1716 1025 -1644
rect 1409 -1761 1410 -1715
rect 107 -1761 108 -1717
rect 450 -1718 451 -1644
rect 502 -1718 503 -1644
rect 1024 -1761 1025 -1717
rect 1045 -1761 1046 -1717
rect 1164 -1718 1165 -1644
rect 1402 -1761 1403 -1717
rect 1423 -1718 1424 -1644
rect 247 -1720 248 -1644
rect 373 -1761 374 -1719
rect 534 -1761 535 -1719
rect 793 -1720 794 -1644
rect 1052 -1720 1053 -1644
rect 1122 -1761 1123 -1719
rect 1164 -1761 1165 -1719
rect 1276 -1720 1277 -1644
rect 1423 -1761 1424 -1719
rect 1437 -1720 1438 -1644
rect 145 -1722 146 -1644
rect 247 -1761 248 -1721
rect 331 -1722 332 -1644
rect 450 -1761 451 -1721
rect 793 -1761 794 -1721
rect 1311 -1722 1312 -1644
rect 331 -1761 332 -1723
rect 352 -1724 353 -1644
rect 810 -1761 811 -1723
rect 1052 -1761 1053 -1723
rect 1066 -1724 1067 -1644
rect 1388 -1761 1389 -1723
rect 338 -1726 339 -1644
rect 352 -1761 353 -1725
rect 992 -1726 993 -1644
rect 1311 -1761 1312 -1725
rect 30 -1728 31 -1644
rect 338 -1761 339 -1727
rect 992 -1761 993 -1727
rect 1339 -1728 1340 -1644
rect 16 -1730 17 -1644
rect 30 -1761 31 -1729
rect 646 -1730 647 -1644
rect 1339 -1761 1340 -1729
rect 16 -1761 17 -1731
rect 100 -1732 101 -1644
rect 646 -1761 647 -1731
rect 681 -1732 682 -1644
rect 1066 -1761 1067 -1731
rect 1115 -1732 1116 -1644
rect 1276 -1761 1277 -1731
rect 1360 -1732 1361 -1644
rect 100 -1761 101 -1733
rect 191 -1734 192 -1644
rect 530 -1761 531 -1733
rect 1115 -1761 1116 -1733
rect 191 -1761 192 -1735
rect 509 -1761 510 -1735
rect 681 -1761 682 -1735
rect 702 -1736 703 -1644
rect 716 -1761 717 -1735
rect 1360 -1761 1361 -1735
rect 702 -1761 703 -1737
rect 772 -1738 773 -1644
rect 1073 -1761 1074 -1737
rect 1178 -1738 1179 -1644
rect 772 -1761 773 -1739
rect 1269 -1740 1270 -1644
rect 1108 -1761 1109 -1741
rect 1136 -1742 1137 -1644
rect 1178 -1761 1179 -1741
rect 1381 -1742 1382 -1644
rect 1136 -1761 1137 -1743
rect 1325 -1744 1326 -1644
rect 1374 -1761 1375 -1743
rect 1381 -1761 1382 -1743
rect 618 -1746 619 -1644
rect 1325 -1761 1326 -1745
rect 44 -1748 45 -1644
rect 618 -1761 619 -1747
rect 1213 -1748 1214 -1644
rect 1269 -1761 1270 -1747
rect 44 -1761 45 -1749
rect 226 -1750 227 -1644
rect 1213 -1761 1214 -1749
rect 1395 -1750 1396 -1644
rect 86 -1752 87 -1644
rect 226 -1761 227 -1751
rect 1353 -1752 1354 -1644
rect 1395 -1761 1396 -1751
rect 86 -1761 87 -1753
rect 170 -1754 171 -1644
rect 1353 -1761 1354 -1753
rect 1416 -1754 1417 -1644
rect 170 -1761 171 -1755
rect 457 -1756 458 -1644
rect 912 -1756 913 -1644
rect 1416 -1761 1417 -1755
rect 457 -1761 458 -1757
rect 583 -1761 584 -1757
rect 912 -1761 913 -1757
rect 1059 -1758 1060 -1644
rect 1059 -1761 1060 -1759
rect 1370 -1761 1371 -1759
rect 2 -1858 3 -1770
rect 590 -1771 591 -1769
rect 667 -1771 668 -1769
rect 842 -1771 843 -1769
rect 877 -1771 878 -1769
rect 1157 -1771 1158 -1769
rect 1164 -1771 1165 -1769
rect 1164 -1858 1165 -1770
rect 1164 -1771 1165 -1769
rect 1164 -1858 1165 -1770
rect 1255 -1771 1256 -1769
rect 1258 -1771 1259 -1769
rect 1360 -1771 1361 -1769
rect 1370 -1771 1371 -1769
rect 1377 -1771 1378 -1769
rect 1395 -1771 1396 -1769
rect 1423 -1771 1424 -1769
rect 1423 -1858 1424 -1770
rect 1423 -1771 1424 -1769
rect 1423 -1858 1424 -1770
rect 19 -1858 20 -1772
rect 534 -1773 535 -1769
rect 562 -1773 563 -1769
rect 590 -1858 591 -1772
rect 667 -1858 668 -1772
rect 681 -1773 682 -1769
rect 684 -1858 685 -1772
rect 786 -1773 787 -1769
rect 793 -1773 794 -1769
rect 835 -1773 836 -1769
rect 842 -1858 843 -1772
rect 863 -1773 864 -1769
rect 887 -1858 888 -1772
rect 968 -1773 969 -1769
rect 1003 -1773 1004 -1769
rect 1066 -1773 1067 -1769
rect 1255 -1858 1256 -1772
rect 1262 -1773 1263 -1769
rect 1367 -1773 1368 -1769
rect 1402 -1773 1403 -1769
rect 61 -1858 62 -1774
rect 1227 -1775 1228 -1769
rect 1346 -1775 1347 -1769
rect 1367 -1858 1368 -1774
rect 1381 -1775 1382 -1769
rect 1430 -1858 1431 -1774
rect 72 -1777 73 -1769
rect 796 -1777 797 -1769
rect 800 -1777 801 -1769
rect 807 -1777 808 -1769
rect 814 -1777 815 -1769
rect 835 -1858 836 -1776
rect 849 -1777 850 -1769
rect 877 -1858 878 -1776
rect 898 -1777 899 -1769
rect 1192 -1777 1193 -1769
rect 1339 -1777 1340 -1769
rect 1346 -1858 1347 -1776
rect 1353 -1777 1354 -1769
rect 1381 -1858 1382 -1776
rect 30 -1779 31 -1769
rect 72 -1858 73 -1778
rect 75 -1779 76 -1769
rect 142 -1779 143 -1769
rect 177 -1779 178 -1769
rect 177 -1858 178 -1778
rect 177 -1779 178 -1769
rect 177 -1858 178 -1778
rect 198 -1779 199 -1769
rect 198 -1858 199 -1778
rect 198 -1779 199 -1769
rect 198 -1858 199 -1778
rect 205 -1779 206 -1769
rect 205 -1858 206 -1778
rect 205 -1779 206 -1769
rect 205 -1858 206 -1778
rect 247 -1779 248 -1769
rect 880 -1779 881 -1769
rect 898 -1858 899 -1778
rect 940 -1779 941 -1769
rect 968 -1858 969 -1778
rect 1059 -1779 1060 -1769
rect 1066 -1858 1067 -1778
rect 1108 -1779 1109 -1769
rect 1332 -1779 1333 -1769
rect 1339 -1858 1340 -1778
rect 1353 -1858 1354 -1778
rect 1374 -1779 1375 -1769
rect 23 -1781 24 -1769
rect 30 -1858 31 -1780
rect 89 -1858 90 -1780
rect 310 -1781 311 -1769
rect 324 -1781 325 -1769
rect 369 -1781 370 -1769
rect 373 -1781 374 -1769
rect 502 -1858 503 -1780
rect 513 -1781 514 -1769
rect 786 -1858 787 -1780
rect 793 -1858 794 -1780
rect 1395 -1858 1396 -1780
rect 23 -1858 24 -1782
rect 632 -1783 633 -1769
rect 635 -1783 636 -1769
rect 1192 -1858 1193 -1782
rect 1234 -1783 1235 -1769
rect 1332 -1858 1333 -1782
rect 51 -1785 52 -1769
rect 632 -1858 633 -1784
rect 674 -1785 675 -1769
rect 674 -1858 675 -1784
rect 674 -1785 675 -1769
rect 674 -1858 675 -1784
rect 691 -1858 692 -1784
rect 1248 -1785 1249 -1769
rect 1325 -1785 1326 -1769
rect 1374 -1858 1375 -1784
rect 51 -1858 52 -1786
rect 121 -1787 122 -1769
rect 138 -1858 139 -1786
rect 415 -1787 416 -1769
rect 436 -1787 437 -1769
rect 439 -1799 440 -1786
rect 464 -1787 465 -1769
rect 509 -1787 510 -1769
rect 513 -1858 514 -1786
rect 541 -1787 542 -1769
rect 569 -1787 570 -1769
rect 814 -1858 815 -1786
rect 849 -1858 850 -1786
rect 856 -1787 857 -1769
rect 863 -1858 864 -1786
rect 891 -1787 892 -1769
rect 908 -1858 909 -1786
rect 1150 -1787 1151 -1769
rect 1178 -1787 1179 -1769
rect 1325 -1858 1326 -1786
rect 58 -1789 59 -1769
rect 121 -1858 122 -1788
rect 191 -1789 192 -1769
rect 373 -1858 374 -1788
rect 380 -1789 381 -1769
rect 562 -1858 563 -1788
rect 569 -1858 570 -1788
rect 765 -1789 766 -1769
rect 800 -1858 801 -1788
rect 1010 -1789 1011 -1769
rect 1129 -1789 1130 -1769
rect 1150 -1858 1151 -1788
rect 1234 -1858 1235 -1788
rect 1388 -1789 1389 -1769
rect 9 -1791 10 -1769
rect 58 -1858 59 -1790
rect 82 -1791 83 -1769
rect 891 -1858 892 -1790
rect 926 -1791 927 -1769
rect 1157 -1858 1158 -1790
rect 1241 -1791 1242 -1769
rect 1248 -1858 1249 -1790
rect 9 -1858 10 -1792
rect 156 -1793 157 -1769
rect 191 -1858 192 -1792
rect 268 -1793 269 -1769
rect 275 -1793 276 -1769
rect 663 -1858 664 -1792
rect 716 -1793 717 -1769
rect 1108 -1858 1109 -1792
rect 1136 -1793 1137 -1769
rect 1241 -1858 1242 -1792
rect 37 -1795 38 -1769
rect 156 -1858 157 -1794
rect 212 -1795 213 -1769
rect 268 -1858 269 -1794
rect 289 -1795 290 -1769
rect 299 -1858 300 -1794
rect 310 -1858 311 -1794
rect 422 -1795 423 -1769
rect 436 -1858 437 -1794
rect 464 -1858 465 -1794
rect 695 -1795 696 -1769
rect 719 -1795 720 -1769
rect 982 -1795 983 -1769
rect 989 -1795 990 -1769
rect 1129 -1858 1130 -1794
rect 107 -1797 108 -1769
rect 397 -1858 398 -1796
rect 415 -1858 416 -1796
rect 604 -1797 605 -1769
rect 611 -1797 612 -1769
rect 807 -1858 808 -1796
rect 810 -1797 811 -1769
rect 1388 -1858 1389 -1796
rect 100 -1799 101 -1769
rect 107 -1858 108 -1798
rect 114 -1799 115 -1769
rect 142 -1858 143 -1798
rect 212 -1858 213 -1798
rect 366 -1799 367 -1769
rect 380 -1858 381 -1798
rect 443 -1799 444 -1769
rect 527 -1799 528 -1769
rect 751 -1799 752 -1769
rect 765 -1858 766 -1798
rect 779 -1799 780 -1769
rect 803 -1858 804 -1798
rect 1227 -1858 1228 -1798
rect 1258 -1858 1259 -1798
rect 1262 -1858 1263 -1798
rect 100 -1858 101 -1800
rect 184 -1801 185 -1769
rect 226 -1801 227 -1769
rect 275 -1858 276 -1800
rect 296 -1801 297 -1769
rect 366 -1858 367 -1800
rect 387 -1801 388 -1769
rect 520 -1858 521 -1800
rect 527 -1858 528 -1800
rect 702 -1801 703 -1769
rect 719 -1858 720 -1800
rect 828 -1801 829 -1769
rect 856 -1858 857 -1800
rect 884 -1801 885 -1769
rect 926 -1858 927 -1800
rect 961 -1801 962 -1769
rect 989 -1858 990 -1800
rect 1171 -1801 1172 -1769
rect 65 -1803 66 -1769
rect 184 -1858 185 -1802
rect 247 -1858 248 -1802
rect 254 -1803 255 -1769
rect 261 -1803 262 -1769
rect 485 -1803 486 -1769
rect 534 -1858 535 -1802
rect 730 -1803 731 -1769
rect 737 -1803 738 -1769
rect 754 -1858 755 -1802
rect 779 -1858 780 -1802
rect 1220 -1803 1221 -1769
rect 65 -1858 66 -1804
rect 86 -1805 87 -1769
rect 114 -1858 115 -1804
rect 149 -1805 150 -1769
rect 163 -1805 164 -1769
rect 226 -1858 227 -1804
rect 233 -1805 234 -1769
rect 261 -1858 262 -1804
rect 296 -1858 297 -1804
rect 1062 -1858 1063 -1804
rect 1094 -1805 1095 -1769
rect 1220 -1858 1221 -1804
rect 135 -1807 136 -1769
rect 149 -1858 150 -1806
rect 163 -1858 164 -1806
rect 170 -1807 171 -1769
rect 233 -1858 234 -1806
rect 345 -1807 346 -1769
rect 352 -1807 353 -1769
rect 443 -1858 444 -1806
rect 485 -1858 486 -1806
rect 884 -1858 885 -1806
rect 919 -1807 920 -1769
rect 1171 -1858 1172 -1806
rect 37 -1858 38 -1808
rect 135 -1858 136 -1808
rect 240 -1809 241 -1769
rect 254 -1858 255 -1808
rect 324 -1858 325 -1808
rect 576 -1809 577 -1769
rect 604 -1858 605 -1808
rect 618 -1809 619 -1769
rect 695 -1858 696 -1808
rect 723 -1809 724 -1769
rect 737 -1858 738 -1808
rect 1017 -1809 1018 -1769
rect 1087 -1809 1088 -1769
rect 1094 -1858 1095 -1808
rect 1122 -1809 1123 -1769
rect 1136 -1858 1137 -1808
rect 44 -1811 45 -1769
rect 345 -1858 346 -1810
rect 352 -1858 353 -1810
rect 471 -1811 472 -1769
rect 488 -1811 489 -1769
rect 576 -1858 577 -1810
rect 611 -1858 612 -1810
rect 646 -1811 647 -1769
rect 702 -1858 703 -1810
rect 709 -1811 710 -1769
rect 723 -1858 724 -1810
rect 936 -1858 937 -1810
rect 940 -1858 941 -1810
rect 1416 -1811 1417 -1769
rect 44 -1858 45 -1812
rect 408 -1813 409 -1769
rect 492 -1813 493 -1769
rect 730 -1858 731 -1812
rect 744 -1813 745 -1769
rect 982 -1858 983 -1812
rect 996 -1813 997 -1769
rect 1003 -1858 1004 -1812
rect 1006 -1813 1007 -1769
rect 1318 -1813 1319 -1769
rect 93 -1815 94 -1769
rect 170 -1858 171 -1814
rect 240 -1858 241 -1814
rect 450 -1815 451 -1769
rect 530 -1815 531 -1769
rect 744 -1858 745 -1814
rect 751 -1858 752 -1814
rect 961 -1858 962 -1814
rect 975 -1815 976 -1769
rect 1017 -1858 1018 -1814
rect 1073 -1815 1074 -1769
rect 1087 -1858 1088 -1814
rect 1311 -1815 1312 -1769
rect 1318 -1858 1319 -1814
rect 93 -1858 94 -1816
rect 418 -1817 419 -1769
rect 450 -1858 451 -1816
rect 775 -1817 776 -1769
rect 821 -1817 822 -1769
rect 828 -1858 829 -1816
rect 870 -1817 871 -1769
rect 1416 -1858 1417 -1816
rect 128 -1819 129 -1769
rect 471 -1858 472 -1818
rect 506 -1819 507 -1769
rect 975 -1858 976 -1818
rect 996 -1858 997 -1818
rect 1143 -1819 1144 -1769
rect 1304 -1819 1305 -1769
rect 1311 -1858 1312 -1818
rect 128 -1858 129 -1820
rect 593 -1858 594 -1820
rect 597 -1821 598 -1769
rect 821 -1858 822 -1820
rect 870 -1858 871 -1820
rect 912 -1821 913 -1769
rect 919 -1858 920 -1820
rect 1080 -1821 1081 -1769
rect 1115 -1821 1116 -1769
rect 1143 -1858 1144 -1820
rect 1297 -1821 1298 -1769
rect 1304 -1858 1305 -1820
rect 317 -1823 318 -1769
rect 408 -1858 409 -1822
rect 478 -1823 479 -1769
rect 506 -1858 507 -1822
rect 541 -1858 542 -1822
rect 548 -1823 549 -1769
rect 555 -1823 556 -1769
rect 597 -1858 598 -1822
rect 618 -1858 619 -1822
rect 1024 -1823 1025 -1769
rect 1045 -1823 1046 -1769
rect 1073 -1858 1074 -1822
rect 1290 -1823 1291 -1769
rect 1297 -1858 1298 -1822
rect 282 -1825 283 -1769
rect 317 -1858 318 -1824
rect 331 -1825 332 -1769
rect 422 -1858 423 -1824
rect 432 -1858 433 -1824
rect 1045 -1858 1046 -1824
rect 1052 -1825 1053 -1769
rect 1080 -1858 1081 -1824
rect 1283 -1825 1284 -1769
rect 1290 -1858 1291 -1824
rect 282 -1858 283 -1826
rect 359 -1827 360 -1769
rect 387 -1858 388 -1826
rect 653 -1827 654 -1769
rect 681 -1858 682 -1826
rect 1115 -1858 1116 -1826
rect 219 -1829 220 -1769
rect 359 -1858 360 -1828
rect 401 -1829 402 -1769
rect 548 -1858 549 -1828
rect 555 -1858 556 -1828
rect 688 -1829 689 -1769
rect 709 -1858 710 -1828
rect 905 -1829 906 -1769
rect 933 -1829 934 -1769
rect 1024 -1858 1025 -1828
rect 1031 -1829 1032 -1769
rect 1052 -1858 1053 -1828
rect 1101 -1829 1102 -1769
rect 1283 -1858 1284 -1828
rect 79 -1831 80 -1769
rect 219 -1858 220 -1830
rect 303 -1831 304 -1769
rect 331 -1858 332 -1830
rect 338 -1831 339 -1769
rect 492 -1858 493 -1830
rect 558 -1858 559 -1830
rect 912 -1858 913 -1830
rect 1010 -1858 1011 -1830
rect 1206 -1831 1207 -1769
rect 16 -1833 17 -1769
rect 79 -1858 80 -1832
rect 303 -1858 304 -1832
rect 394 -1833 395 -1769
rect 401 -1858 402 -1832
rect 845 -1833 846 -1769
rect 873 -1833 874 -1769
rect 1122 -1858 1123 -1832
rect 1185 -1833 1186 -1769
rect 1206 -1858 1207 -1832
rect 86 -1858 87 -1834
rect 1185 -1858 1186 -1834
rect 338 -1858 339 -1836
rect 583 -1837 584 -1769
rect 586 -1837 587 -1769
rect 905 -1858 906 -1836
rect 1031 -1858 1032 -1836
rect 1038 -1837 1039 -1769
rect 1101 -1858 1102 -1836
rect 1409 -1837 1410 -1769
rect 341 -1839 342 -1769
rect 1213 -1839 1214 -1769
rect 394 -1858 395 -1840
rect 1360 -1858 1361 -1840
rect 478 -1858 479 -1842
rect 499 -1843 500 -1769
rect 583 -1858 584 -1842
rect 639 -1843 640 -1769
rect 653 -1858 654 -1842
rect 758 -1843 759 -1769
rect 901 -1843 902 -1769
rect 1409 -1858 1410 -1842
rect 289 -1858 290 -1844
rect 499 -1858 500 -1844
rect 625 -1845 626 -1769
rect 646 -1858 647 -1844
rect 688 -1858 689 -1844
rect 1178 -1858 1179 -1844
rect 1199 -1845 1200 -1769
rect 1213 -1858 1214 -1844
rect 625 -1858 626 -1846
rect 660 -1847 661 -1769
rect 716 -1858 717 -1846
rect 758 -1858 759 -1846
rect 954 -1847 955 -1769
rect 1199 -1858 1200 -1846
rect 639 -1858 640 -1848
rect 933 -1858 934 -1848
rect 947 -1849 948 -1769
rect 954 -1858 955 -1848
rect 1038 -1858 1039 -1848
rect 1276 -1849 1277 -1769
rect 572 -1858 573 -1850
rect 947 -1858 948 -1850
rect 1269 -1851 1270 -1769
rect 1276 -1858 1277 -1850
rect 660 -1858 661 -1852
rect 1402 -1858 1403 -1852
rect 772 -1855 773 -1769
rect 1269 -1858 1270 -1854
rect 429 -1857 430 -1769
rect 772 -1858 773 -1856
rect 2 -1868 3 -1866
rect 5 -1976 6 -1867
rect 9 -1868 10 -1866
rect 397 -1868 398 -1866
rect 432 -1868 433 -1866
rect 744 -1868 745 -1866
rect 751 -1868 752 -1866
rect 1283 -1868 1284 -1866
rect 1395 -1868 1396 -1866
rect 1423 -1868 1424 -1866
rect 2 -1985 3 -1869
rect 51 -1870 52 -1866
rect 100 -1870 101 -1866
rect 299 -1870 300 -1866
rect 303 -1870 304 -1866
rect 303 -1985 304 -1869
rect 303 -1870 304 -1866
rect 303 -1985 304 -1869
rect 373 -1870 374 -1866
rect 558 -1870 559 -1866
rect 565 -1985 566 -1869
rect 912 -1870 913 -1866
rect 933 -1870 934 -1866
rect 1381 -1870 1382 -1866
rect 9 -1985 10 -1871
rect 261 -1872 262 -1866
rect 282 -1872 283 -1866
rect 345 -1872 346 -1866
rect 471 -1872 472 -1866
rect 614 -1985 615 -1871
rect 618 -1872 619 -1866
rect 772 -1872 773 -1866
rect 775 -1872 776 -1866
rect 968 -1872 969 -1866
rect 1062 -1872 1063 -1866
rect 1262 -1872 1263 -1866
rect 19 -1874 20 -1866
rect 75 -1985 76 -1873
rect 100 -1985 101 -1873
rect 114 -1874 115 -1866
rect 128 -1874 129 -1866
rect 936 -1874 937 -1866
rect 968 -1985 969 -1873
rect 975 -1874 976 -1866
rect 1234 -1874 1235 -1866
rect 1395 -1985 1396 -1873
rect 26 -1985 27 -1875
rect 30 -1876 31 -1866
rect 37 -1876 38 -1866
rect 394 -1876 395 -1866
rect 401 -1876 402 -1866
rect 471 -1985 472 -1875
rect 499 -1876 500 -1866
rect 597 -1876 598 -1866
rect 618 -1985 619 -1875
rect 803 -1876 804 -1866
rect 856 -1876 857 -1866
rect 905 -1985 906 -1875
rect 912 -1985 913 -1875
rect 926 -1876 927 -1866
rect 933 -1985 934 -1875
rect 1003 -1876 1004 -1866
rect 1066 -1876 1067 -1866
rect 1234 -1985 1235 -1875
rect 30 -1985 31 -1877
rect 457 -1878 458 -1866
rect 502 -1878 503 -1866
rect 1381 -1985 1382 -1877
rect 37 -1985 38 -1879
rect 1199 -1880 1200 -1866
rect 44 -1882 45 -1866
rect 509 -1985 510 -1881
rect 523 -1985 524 -1881
rect 1206 -1882 1207 -1866
rect 44 -1985 45 -1883
rect 604 -1884 605 -1866
rect 646 -1884 647 -1866
rect 663 -1884 664 -1866
rect 681 -1884 682 -1866
rect 1398 -1884 1399 -1866
rect 51 -1985 52 -1885
rect 212 -1886 213 -1866
rect 219 -1886 220 -1866
rect 401 -1985 402 -1885
rect 527 -1886 528 -1866
rect 597 -1985 598 -1885
rect 604 -1985 605 -1885
rect 1059 -1886 1060 -1866
rect 1199 -1985 1200 -1885
rect 1241 -1886 1242 -1866
rect 58 -1888 59 -1866
rect 856 -1985 857 -1887
rect 884 -1888 885 -1866
rect 1430 -1888 1431 -1866
rect 58 -1985 59 -1889
rect 513 -1890 514 -1866
rect 555 -1985 556 -1889
rect 625 -1890 626 -1866
rect 660 -1890 661 -1866
rect 1157 -1890 1158 -1866
rect 1206 -1985 1207 -1889
rect 1297 -1890 1298 -1866
rect 40 -1985 41 -1891
rect 1157 -1985 1158 -1891
rect 1241 -1985 1242 -1891
rect 1255 -1892 1256 -1866
rect 1297 -1985 1298 -1891
rect 1332 -1892 1333 -1866
rect 61 -1894 62 -1866
rect 261 -1985 262 -1893
rect 282 -1985 283 -1893
rect 408 -1894 409 -1866
rect 513 -1985 514 -1893
rect 723 -1894 724 -1866
rect 726 -1985 727 -1893
rect 1262 -1985 1263 -1893
rect 1332 -1985 1333 -1893
rect 1367 -1894 1368 -1866
rect 79 -1896 80 -1866
rect 212 -1985 213 -1895
rect 219 -1985 220 -1895
rect 352 -1896 353 -1866
rect 355 -1985 356 -1895
rect 975 -1985 976 -1895
rect 996 -1896 997 -1866
rect 1066 -1985 1067 -1895
rect 1122 -1896 1123 -1866
rect 1367 -1985 1368 -1895
rect 79 -1985 80 -1897
rect 142 -1898 143 -1866
rect 170 -1898 171 -1866
rect 642 -1985 643 -1897
rect 688 -1898 689 -1866
rect 1171 -1898 1172 -1866
rect 1255 -1985 1256 -1897
rect 1311 -1898 1312 -1866
rect 89 -1900 90 -1866
rect 646 -1985 647 -1899
rect 660 -1985 661 -1899
rect 688 -1985 689 -1899
rect 691 -1900 692 -1866
rect 1171 -1985 1172 -1899
rect 1311 -1985 1312 -1899
rect 1339 -1900 1340 -1866
rect 121 -1902 122 -1866
rect 499 -1985 500 -1901
rect 625 -1985 626 -1901
rect 709 -1902 710 -1866
rect 737 -1902 738 -1866
rect 996 -1985 997 -1901
rect 1003 -1985 1004 -1901
rect 1073 -1902 1074 -1866
rect 1122 -1985 1123 -1901
rect 1220 -1902 1221 -1866
rect 1339 -1985 1340 -1901
rect 1388 -1902 1389 -1866
rect 121 -1985 122 -1903
rect 506 -1904 507 -1866
rect 702 -1904 703 -1866
rect 719 -1904 720 -1866
rect 737 -1985 738 -1903
rect 807 -1904 808 -1866
rect 870 -1904 871 -1866
rect 884 -1985 885 -1903
rect 926 -1985 927 -1903
rect 1017 -1904 1018 -1866
rect 1038 -1904 1039 -1866
rect 1220 -1985 1221 -1903
rect 1388 -1985 1389 -1903
rect 1416 -1904 1417 -1866
rect 128 -1985 129 -1905
rect 443 -1906 444 -1866
rect 506 -1985 507 -1905
rect 1248 -1906 1249 -1866
rect 135 -1908 136 -1866
rect 1143 -1908 1144 -1866
rect 1248 -1985 1249 -1907
rect 1304 -1908 1305 -1866
rect 135 -1985 136 -1909
rect 149 -1910 150 -1866
rect 170 -1985 171 -1909
rect 1374 -1910 1375 -1866
rect 142 -1985 143 -1911
rect 296 -1912 297 -1866
rect 338 -1912 339 -1866
rect 1017 -1985 1018 -1911
rect 1038 -1985 1039 -1911
rect 1108 -1912 1109 -1866
rect 1143 -1985 1144 -1911
rect 1192 -1912 1193 -1866
rect 1374 -1985 1375 -1911
rect 1409 -1912 1410 -1866
rect 149 -1985 150 -1913
rect 667 -1914 668 -1866
rect 716 -1914 717 -1866
rect 1304 -1985 1305 -1913
rect 205 -1916 206 -1866
rect 569 -1916 570 -1866
rect 611 -1916 612 -1866
rect 702 -1985 703 -1915
rect 716 -1985 717 -1915
rect 758 -1916 759 -1866
rect 772 -1985 773 -1915
rect 828 -1916 829 -1866
rect 870 -1985 871 -1915
rect 891 -1916 892 -1866
rect 1059 -1985 1060 -1915
rect 1129 -1916 1130 -1866
rect 1192 -1985 1193 -1915
rect 1276 -1916 1277 -1866
rect 205 -1985 206 -1917
rect 331 -1918 332 -1866
rect 338 -1985 339 -1917
rect 366 -1918 367 -1866
rect 387 -1918 388 -1866
rect 663 -1985 664 -1917
rect 744 -1985 745 -1917
rect 821 -1918 822 -1866
rect 828 -1985 829 -1917
rect 863 -1918 864 -1866
rect 891 -1985 892 -1917
rect 947 -1918 948 -1866
rect 1108 -1985 1109 -1917
rect 1402 -1918 1403 -1866
rect 93 -1920 94 -1866
rect 863 -1985 864 -1919
rect 898 -1920 899 -1866
rect 947 -1985 948 -1919
rect 1024 -1920 1025 -1866
rect 1402 -1985 1403 -1919
rect 93 -1985 94 -1921
rect 198 -1922 199 -1866
rect 233 -1922 234 -1866
rect 429 -1922 430 -1866
rect 492 -1922 493 -1866
rect 667 -1985 668 -1921
rect 751 -1985 752 -1921
rect 1073 -1985 1074 -1921
rect 1129 -1985 1130 -1921
rect 1325 -1922 1326 -1866
rect 198 -1985 199 -1923
rect 786 -1924 787 -1866
rect 800 -1924 801 -1866
rect 954 -1924 955 -1866
rect 1024 -1985 1025 -1923
rect 1087 -1924 1088 -1866
rect 1276 -1985 1277 -1923
rect 1318 -1924 1319 -1866
rect 1325 -1985 1326 -1923
rect 1353 -1924 1354 -1866
rect 86 -1926 87 -1866
rect 1353 -1985 1354 -1925
rect 86 -1985 87 -1927
rect 348 -1928 349 -1866
rect 352 -1985 353 -1927
rect 387 -1985 388 -1927
rect 408 -1985 409 -1927
rect 527 -1985 528 -1927
rect 569 -1985 570 -1927
rect 576 -1928 577 -1866
rect 611 -1985 612 -1927
rect 709 -1985 710 -1927
rect 723 -1985 724 -1927
rect 786 -1985 787 -1927
rect 800 -1985 801 -1927
rect 940 -1928 941 -1866
rect 954 -1985 955 -1927
rect 1045 -1928 1046 -1866
rect 1087 -1985 1088 -1927
rect 1269 -1928 1270 -1866
rect 1318 -1985 1319 -1927
rect 1346 -1928 1347 -1866
rect 138 -1930 139 -1866
rect 1045 -1985 1046 -1929
rect 1346 -1985 1347 -1929
rect 1360 -1930 1361 -1866
rect 233 -1985 234 -1931
rect 632 -1932 633 -1866
rect 653 -1932 654 -1866
rect 898 -1985 899 -1931
rect 940 -1985 941 -1931
rect 1115 -1932 1116 -1866
rect 240 -1934 241 -1866
rect 684 -1934 685 -1866
rect 754 -1934 755 -1866
rect 877 -1934 878 -1866
rect 989 -1934 990 -1866
rect 1360 -1985 1361 -1933
rect 240 -1985 241 -1935
rect 422 -1936 423 -1866
rect 429 -1985 430 -1935
rect 908 -1936 909 -1866
rect 989 -1985 990 -1935
rect 1052 -1936 1053 -1866
rect 1115 -1985 1116 -1935
rect 1185 -1936 1186 -1866
rect 191 -1938 192 -1866
rect 422 -1985 423 -1937
rect 464 -1938 465 -1866
rect 492 -1985 493 -1937
rect 520 -1938 521 -1866
rect 576 -1985 577 -1937
rect 674 -1938 675 -1866
rect 754 -1985 755 -1937
rect 758 -1985 759 -1937
rect 765 -1938 766 -1866
rect 782 -1985 783 -1937
rect 1101 -1938 1102 -1866
rect 1150 -1938 1151 -1866
rect 1185 -1985 1186 -1937
rect 72 -1940 73 -1866
rect 191 -1985 192 -1939
rect 247 -1940 248 -1866
rect 394 -1985 395 -1939
rect 464 -1985 465 -1939
rect 793 -1940 794 -1866
rect 807 -1985 808 -1939
rect 1283 -1985 1284 -1939
rect 72 -1985 73 -1941
rect 173 -1985 174 -1941
rect 254 -1942 255 -1866
rect 254 -1985 255 -1941
rect 254 -1942 255 -1866
rect 254 -1985 255 -1941
rect 268 -1942 269 -1866
rect 443 -1985 444 -1941
rect 485 -1942 486 -1866
rect 793 -1985 794 -1941
rect 821 -1985 822 -1941
rect 849 -1942 850 -1866
rect 1010 -1942 1011 -1866
rect 1150 -1985 1151 -1941
rect 107 -1944 108 -1866
rect 247 -1985 248 -1943
rect 268 -1985 269 -1943
rect 275 -1944 276 -1866
rect 289 -1944 290 -1866
rect 632 -1985 633 -1943
rect 765 -1985 766 -1943
rect 814 -1944 815 -1866
rect 835 -1944 836 -1866
rect 877 -1985 878 -1943
rect 1010 -1985 1011 -1943
rect 1080 -1944 1081 -1866
rect 1101 -1985 1102 -1943
rect 1178 -1944 1179 -1866
rect 16 -1946 17 -1866
rect 107 -1985 108 -1945
rect 163 -1946 164 -1866
rect 289 -1985 290 -1945
rect 296 -1985 297 -1945
rect 541 -1946 542 -1866
rect 572 -1946 573 -1866
rect 814 -1985 815 -1945
rect 835 -1985 836 -1945
rect 842 -1946 843 -1866
rect 1052 -1985 1053 -1945
rect 1094 -1946 1095 -1866
rect 1178 -1985 1179 -1945
rect 1227 -1946 1228 -1866
rect 16 -1985 17 -1947
rect 23 -1948 24 -1866
rect 163 -1985 164 -1947
rect 593 -1948 594 -1866
rect 842 -1985 843 -1947
rect 961 -1948 962 -1866
rect 1080 -1985 1081 -1947
rect 1136 -1948 1137 -1866
rect 23 -1985 24 -1949
rect 1213 -1950 1214 -1866
rect 229 -1985 230 -1951
rect 275 -1985 276 -1951
rect 310 -1952 311 -1866
rect 485 -1985 486 -1951
rect 579 -1985 580 -1951
rect 674 -1985 675 -1951
rect 705 -1985 706 -1951
rect 1136 -1985 1137 -1951
rect 1213 -1985 1214 -1951
rect 1290 -1952 1291 -1866
rect 310 -1985 311 -1953
rect 324 -1954 325 -1866
rect 331 -1985 332 -1953
rect 548 -1954 549 -1866
rect 887 -1954 888 -1866
rect 1290 -1985 1291 -1953
rect 65 -1956 66 -1866
rect 324 -1985 325 -1955
rect 345 -1985 346 -1955
rect 516 -1985 517 -1955
rect 548 -1985 549 -1955
rect 562 -1956 563 -1866
rect 961 -1985 962 -1955
rect 982 -1956 983 -1866
rect 1094 -1985 1095 -1955
rect 1164 -1956 1165 -1866
rect 65 -1985 66 -1957
rect 114 -1985 115 -1957
rect 317 -1958 318 -1866
rect 562 -1985 563 -1957
rect 779 -1958 780 -1866
rect 1164 -1985 1165 -1957
rect 317 -1985 318 -1959
rect 436 -1960 437 -1866
rect 478 -1960 479 -1866
rect 541 -1985 542 -1959
rect 681 -1985 682 -1959
rect 779 -1985 780 -1959
rect 982 -1985 983 -1959
rect 1031 -1960 1032 -1866
rect 359 -1962 360 -1866
rect 457 -1985 458 -1961
rect 919 -1962 920 -1866
rect 1031 -1985 1032 -1961
rect 359 -1985 360 -1963
rect 450 -1964 451 -1866
rect 590 -1964 591 -1866
rect 919 -1985 920 -1963
rect 177 -1966 178 -1866
rect 450 -1985 451 -1965
rect 583 -1966 584 -1866
rect 590 -1985 591 -1965
rect 177 -1985 178 -1967
rect 226 -1968 227 -1866
rect 366 -1985 367 -1967
rect 639 -1968 640 -1866
rect 184 -1970 185 -1866
rect 226 -1985 227 -1969
rect 373 -1985 374 -1969
rect 1269 -1985 1270 -1969
rect 68 -1985 69 -1971
rect 184 -1985 185 -1971
rect 380 -1972 381 -1866
rect 520 -1985 521 -1971
rect 583 -1985 584 -1971
rect 1227 -1985 1228 -1971
rect 156 -1974 157 -1866
rect 380 -1985 381 -1973
rect 415 -1974 416 -1866
rect 478 -1985 479 -1973
rect 639 -1985 640 -1973
rect 653 -1985 654 -1973
rect 415 -1985 416 -1975
rect 436 -1985 437 -1975
rect 852 -1985 853 -1975
rect 156 -1985 157 -1977
rect 695 -1978 696 -1866
rect 695 -1985 696 -1979
rect 730 -1980 731 -1866
rect 534 -1982 535 -1866
rect 730 -1985 731 -1981
rect 411 -1985 412 -1983
rect 534 -1985 535 -1983
rect 2 -1995 3 -1993
rect 37 -1995 38 -1993
rect 51 -1995 52 -1993
rect 660 -1995 661 -1993
rect 663 -1995 664 -1993
rect 996 -1995 997 -1993
rect 1010 -1995 1011 -1993
rect 1010 -2104 1011 -1994
rect 1010 -1995 1011 -1993
rect 1010 -2104 1011 -1994
rect 1024 -1995 1025 -1993
rect 1024 -2104 1025 -1994
rect 1024 -1995 1025 -1993
rect 1024 -2104 1025 -1994
rect 1031 -1995 1032 -1993
rect 1031 -2104 1032 -1994
rect 1031 -1995 1032 -1993
rect 1031 -2104 1032 -1994
rect 1139 -2104 1140 -1994
rect 1367 -1995 1368 -1993
rect 5 -2104 6 -1996
rect 191 -1997 192 -1993
rect 205 -1997 206 -1993
rect 320 -2104 321 -1996
rect 324 -1997 325 -1993
rect 376 -1997 377 -1993
rect 408 -1997 409 -1993
rect 1262 -1997 1263 -1993
rect 37 -2104 38 -1998
rect 338 -1999 339 -1993
rect 408 -2104 409 -1998
rect 541 -1999 542 -1993
rect 579 -1999 580 -1993
rect 1185 -1999 1186 -1993
rect 1262 -2104 1263 -1998
rect 1283 -1999 1284 -1993
rect 51 -2104 52 -2000
rect 261 -2001 262 -1993
rect 268 -2001 269 -1993
rect 355 -2001 356 -1993
rect 373 -2001 374 -1993
rect 1185 -2104 1186 -2000
rect 1283 -2104 1284 -2000
rect 1325 -2001 1326 -1993
rect 58 -2003 59 -1993
rect 488 -2104 489 -2002
rect 502 -2104 503 -2002
rect 1304 -2003 1305 -1993
rect 1325 -2104 1326 -2002
rect 1388 -2003 1389 -1993
rect 58 -2104 59 -2004
rect 247 -2005 248 -1993
rect 261 -2104 262 -2004
rect 387 -2005 388 -1993
rect 411 -2005 412 -1993
rect 1234 -2005 1235 -1993
rect 65 -2007 66 -1993
rect 289 -2007 290 -1993
rect 334 -2104 335 -2006
rect 1276 -2007 1277 -1993
rect 65 -2104 66 -2008
rect 303 -2009 304 -1993
rect 338 -2104 339 -2008
rect 394 -2009 395 -1993
rect 415 -2009 416 -1993
rect 541 -2104 542 -2008
rect 614 -2009 615 -1993
rect 1241 -2009 1242 -1993
rect 68 -2011 69 -1993
rect 324 -2104 325 -2010
rect 373 -2104 374 -2010
rect 478 -2011 479 -1993
rect 513 -2011 514 -1993
rect 1290 -2011 1291 -1993
rect 72 -2013 73 -1993
rect 1227 -2013 1228 -1993
rect 1290 -2104 1291 -2012
rect 1332 -2013 1333 -1993
rect 72 -2104 73 -2014
rect 331 -2015 332 -1993
rect 387 -2104 388 -2014
rect 485 -2015 486 -1993
rect 513 -2104 514 -2014
rect 625 -2015 626 -1993
rect 639 -2015 640 -1993
rect 1080 -2015 1081 -1993
rect 1108 -2015 1109 -1993
rect 1304 -2104 1305 -2014
rect 93 -2017 94 -1993
rect 205 -2104 206 -2016
rect 268 -2104 269 -2016
rect 429 -2017 430 -1993
rect 453 -2104 454 -2016
rect 1241 -2104 1242 -2016
rect 93 -2104 94 -2018
rect 639 -2104 640 -2018
rect 646 -2019 647 -1993
rect 660 -2104 661 -2018
rect 691 -2104 692 -2018
rect 1360 -2019 1361 -1993
rect 96 -2104 97 -2020
rect 100 -2021 101 -1993
rect 107 -2021 108 -1993
rect 247 -2104 248 -2020
rect 289 -2104 290 -2020
rect 436 -2021 437 -1993
rect 478 -2104 479 -2020
rect 527 -2021 528 -1993
rect 604 -2021 605 -1993
rect 625 -2104 626 -2020
rect 646 -2104 647 -2020
rect 681 -2021 682 -1993
rect 705 -2021 706 -1993
rect 772 -2021 773 -1993
rect 782 -2021 783 -1993
rect 821 -2021 822 -1993
rect 849 -2021 850 -1993
rect 933 -2021 934 -1993
rect 947 -2021 948 -1993
rect 1143 -2021 1144 -1993
rect 1213 -2021 1214 -1993
rect 1276 -2104 1277 -2020
rect 100 -2104 101 -2022
rect 173 -2023 174 -1993
rect 177 -2023 178 -1993
rect 331 -2104 332 -2022
rect 415 -2104 416 -2022
rect 492 -2023 493 -1993
rect 516 -2023 517 -1993
rect 765 -2023 766 -1993
rect 807 -2023 808 -1993
rect 1045 -2023 1046 -1993
rect 1059 -2023 1060 -1993
rect 1080 -2104 1081 -2022
rect 1129 -2023 1130 -1993
rect 1234 -2104 1235 -2022
rect 114 -2025 115 -1993
rect 114 -2104 115 -2024
rect 114 -2025 115 -1993
rect 114 -2104 115 -2024
rect 121 -2025 122 -1993
rect 492 -2104 493 -2024
rect 499 -2025 500 -1993
rect 807 -2104 808 -2024
rect 821 -2104 822 -2024
rect 1199 -2025 1200 -1993
rect 1206 -2025 1207 -1993
rect 1213 -2104 1214 -2024
rect 1227 -2104 1228 -2024
rect 1255 -2025 1256 -1993
rect 23 -2027 24 -1993
rect 121 -2104 122 -2026
rect 128 -2027 129 -1993
rect 681 -2104 682 -2026
rect 726 -2027 727 -1993
rect 1402 -2027 1403 -1993
rect 16 -2029 17 -1993
rect 128 -2104 129 -2028
rect 131 -2104 132 -2028
rect 394 -2104 395 -2028
rect 422 -2029 423 -1993
rect 509 -2029 510 -1993
rect 520 -2029 521 -1993
rect 590 -2029 591 -1993
rect 621 -2104 622 -2028
rect 1353 -2029 1354 -1993
rect 16 -2104 17 -2030
rect 240 -2031 241 -1993
rect 296 -2031 297 -1993
rect 499 -2104 500 -2030
rect 520 -2104 521 -2030
rect 817 -2104 818 -2030
rect 849 -2104 850 -2030
rect 856 -2031 857 -1993
rect 877 -2031 878 -1993
rect 877 -2104 878 -2030
rect 877 -2031 878 -1993
rect 877 -2104 878 -2030
rect 884 -2031 885 -1993
rect 884 -2104 885 -2030
rect 884 -2031 885 -1993
rect 884 -2104 885 -2030
rect 912 -2031 913 -1993
rect 1108 -2104 1109 -2030
rect 1129 -2104 1130 -2030
rect 1136 -2031 1137 -1993
rect 1143 -2104 1144 -2030
rect 1164 -2031 1165 -1993
rect 1199 -2104 1200 -2030
rect 1220 -2031 1221 -1993
rect 23 -2104 24 -2032
rect 156 -2033 157 -1993
rect 163 -2033 164 -1993
rect 226 -2033 227 -1993
rect 296 -2104 297 -2032
rect 611 -2033 612 -1993
rect 730 -2033 731 -1993
rect 733 -2055 734 -2032
rect 737 -2033 738 -1993
rect 772 -2104 773 -2032
rect 779 -2033 780 -1993
rect 1164 -2104 1165 -2032
rect 1206 -2104 1207 -2032
rect 1318 -2033 1319 -1993
rect 9 -2035 10 -1993
rect 163 -2104 164 -2034
rect 166 -2104 167 -2034
rect 1017 -2035 1018 -1993
rect 1059 -2104 1060 -2034
rect 1094 -2035 1095 -1993
rect 1220 -2104 1221 -2034
rect 1248 -2035 1249 -1993
rect 1318 -2104 1319 -2034
rect 1381 -2035 1382 -1993
rect 9 -2104 10 -2036
rect 1255 -2104 1256 -2036
rect 135 -2039 136 -1993
rect 156 -2104 157 -2038
rect 173 -2104 174 -2038
rect 212 -2039 213 -1993
rect 219 -2039 220 -1993
rect 240 -2104 241 -2038
rect 303 -2104 304 -2038
rect 310 -2039 311 -1993
rect 422 -2104 423 -2038
rect 450 -2039 451 -1993
rect 527 -2104 528 -2038
rect 548 -2039 549 -1993
rect 555 -2039 556 -1993
rect 604 -2104 605 -2038
rect 716 -2039 717 -1993
rect 737 -2104 738 -2038
rect 754 -2039 755 -1993
rect 898 -2039 899 -1993
rect 933 -2104 934 -2038
rect 992 -2104 993 -2038
rect 996 -2104 997 -2038
rect 1122 -2039 1123 -1993
rect 1248 -2104 1249 -2038
rect 1269 -2039 1270 -1993
rect 110 -2104 111 -2040
rect 212 -2104 213 -2040
rect 219 -2104 220 -2040
rect 534 -2041 535 -1993
rect 548 -2104 549 -2040
rect 782 -2104 783 -2040
rect 842 -2041 843 -1993
rect 912 -2104 913 -2040
rect 968 -2041 969 -1993
rect 1045 -2104 1046 -2040
rect 1094 -2104 1095 -2040
rect 1192 -2041 1193 -1993
rect 1269 -2104 1270 -2040
rect 1311 -2041 1312 -1993
rect 135 -2104 136 -2042
rect 670 -2104 671 -2042
rect 730 -2104 731 -2042
rect 800 -2043 801 -1993
rect 828 -2043 829 -1993
rect 842 -2104 843 -2042
rect 852 -2043 853 -1993
rect 905 -2043 906 -1993
rect 971 -2104 972 -2042
rect 1297 -2043 1298 -1993
rect 1311 -2104 1312 -2042
rect 1374 -2043 1375 -1993
rect 142 -2045 143 -1993
rect 310 -2104 311 -2044
rect 429 -2104 430 -2044
rect 824 -2104 825 -2044
rect 856 -2104 857 -2044
rect 954 -2045 955 -1993
rect 1017 -2104 1018 -2044
rect 1087 -2045 1088 -1993
rect 1101 -2045 1102 -1993
rect 1192 -2104 1193 -2044
rect 1297 -2104 1298 -2044
rect 1339 -2045 1340 -1993
rect 142 -2104 143 -2046
rect 359 -2047 360 -1993
rect 436 -2104 437 -2046
rect 471 -2047 472 -1993
rect 485 -2104 486 -2046
rect 716 -2104 717 -2046
rect 765 -2104 766 -2046
rect 863 -2047 864 -1993
rect 870 -2047 871 -1993
rect 898 -2104 899 -2046
rect 954 -2104 955 -2046
rect 989 -2047 990 -1993
rect 1073 -2047 1074 -1993
rect 1087 -2104 1088 -2046
rect 1101 -2104 1102 -2046
rect 1115 -2047 1116 -1993
rect 30 -2049 31 -1993
rect 359 -2104 360 -2048
rect 443 -2049 444 -1993
rect 450 -2104 451 -2048
rect 457 -2049 458 -1993
rect 471 -2104 472 -2048
rect 555 -2104 556 -2048
rect 586 -2049 587 -1993
rect 590 -2104 591 -2048
rect 632 -2049 633 -1993
rect 779 -2104 780 -2048
rect 1346 -2049 1347 -1993
rect 30 -2104 31 -2050
rect 40 -2051 41 -1993
rect 170 -2051 171 -1993
rect 443 -2104 444 -2050
rect 457 -2104 458 -2050
rect 464 -2051 465 -1993
rect 569 -2051 570 -1993
rect 611 -2104 612 -2050
rect 786 -2051 787 -1993
rect 800 -2104 801 -2050
rect 863 -2104 864 -2050
rect 894 -2104 895 -2050
rect 1066 -2051 1067 -1993
rect 1073 -2104 1074 -2050
rect 75 -2053 76 -1993
rect 170 -2104 171 -2052
rect 177 -2104 178 -2052
rect 723 -2053 724 -1993
rect 744 -2053 745 -1993
rect 786 -2104 787 -2052
rect 870 -2104 871 -2052
rect 1115 -2104 1116 -2052
rect 191 -2104 192 -2054
rect 618 -2055 619 -1993
rect 674 -2055 675 -1993
rect 723 -2104 724 -2054
rect 744 -2104 745 -2054
rect 891 -2055 892 -1993
rect 905 -2104 906 -2054
rect 149 -2057 150 -1993
rect 618 -2104 619 -2056
rect 674 -2104 675 -2056
rect 695 -2057 696 -1993
rect 149 -2104 150 -2058
rect 1157 -2059 1158 -1993
rect 198 -2061 199 -1993
rect 464 -2104 465 -2060
rect 506 -2061 507 -1993
rect 1066 -2104 1067 -2060
rect 184 -2063 185 -1993
rect 198 -2104 199 -2062
rect 226 -2104 227 -2062
rect 751 -2063 752 -1993
rect 184 -2104 185 -2064
rect 254 -2065 255 -1993
rect 562 -2065 563 -1993
rect 1157 -2104 1158 -2064
rect 229 -2067 230 -1993
rect 506 -2104 507 -2066
rect 562 -2104 563 -2066
rect 975 -2067 976 -1993
rect 233 -2069 234 -1993
rect 534 -2104 535 -2068
rect 569 -2104 570 -2068
rect 667 -2069 668 -1993
rect 695 -2104 696 -2068
rect 793 -2069 794 -1993
rect 975 -2104 976 -2068
rect 982 -2069 983 -1993
rect 86 -2071 87 -1993
rect 233 -2104 234 -2070
rect 254 -2104 255 -2070
rect 282 -2071 283 -1993
rect 576 -2071 577 -1993
rect 632 -2104 633 -2070
rect 667 -2104 668 -2070
rect 1150 -2071 1151 -1993
rect 86 -2104 87 -2072
rect 107 -2104 108 -2072
rect 282 -2104 283 -2072
rect 345 -2073 346 -1993
rect 576 -2104 577 -2072
rect 961 -2073 962 -1993
rect 982 -2104 983 -2072
rect 1395 -2073 1396 -1993
rect 345 -2104 346 -2074
rect 401 -2075 402 -1993
rect 579 -2104 580 -2074
rect 947 -2104 948 -2074
rect 1150 -2104 1151 -2074
rect 1171 -2075 1172 -1993
rect 401 -2104 402 -2076
rect 642 -2077 643 -1993
rect 751 -2104 752 -2076
rect 758 -2077 759 -1993
rect 793 -2104 794 -2076
rect 1003 -2077 1004 -1993
rect 1171 -2104 1172 -2076
rect 1178 -2077 1179 -1993
rect 597 -2079 598 -1993
rect 828 -2104 829 -2078
rect 835 -2079 836 -1993
rect 1003 -2104 1004 -2078
rect 523 -2081 524 -1993
rect 597 -2104 598 -2080
rect 688 -2081 689 -1993
rect 758 -2104 759 -2080
rect 814 -2081 815 -1993
rect 835 -2104 836 -2080
rect 926 -2081 927 -1993
rect 961 -2104 962 -2080
rect 583 -2083 584 -1993
rect 688 -2104 689 -2082
rect 709 -2083 710 -1993
rect 1178 -2104 1179 -2082
rect 380 -2085 381 -1993
rect 709 -2104 710 -2084
rect 814 -2104 815 -2084
rect 1052 -2085 1053 -1993
rect 44 -2087 45 -1993
rect 380 -2104 381 -2086
rect 583 -2104 584 -2086
rect 653 -2087 654 -1993
rect 919 -2087 920 -1993
rect 926 -2104 927 -2086
rect 940 -2087 941 -1993
rect 1052 -2104 1053 -2086
rect 2 -2104 3 -2088
rect 653 -2104 654 -2088
rect 940 -2104 941 -2088
rect 1038 -2089 1039 -1993
rect 44 -2104 45 -2090
rect 79 -2091 80 -1993
rect 352 -2091 353 -1993
rect 919 -2104 920 -2090
rect 968 -2104 969 -2090
rect 1038 -2104 1039 -2090
rect 79 -2104 80 -2092
rect 317 -2093 318 -1993
rect 275 -2095 276 -1993
rect 352 -2104 353 -2094
rect 275 -2104 276 -2096
rect 366 -2097 367 -1993
rect 317 -2104 318 -2098
rect 1122 -2104 1123 -2098
rect 366 -2104 367 -2100
rect 702 -2101 703 -1993
rect 702 -2104 703 -2102
rect 810 -2103 811 -1993
rect 9 -2114 10 -2112
rect 44 -2114 45 -2112
rect 51 -2114 52 -2112
rect 667 -2114 668 -2112
rect 765 -2114 766 -2112
rect 768 -2114 769 -2112
rect 793 -2114 794 -2112
rect 891 -2114 892 -2112
rect 936 -2237 937 -2113
rect 975 -2114 976 -2112
rect 989 -2114 990 -2112
rect 1045 -2114 1046 -2112
rect 1115 -2114 1116 -2112
rect 1262 -2114 1263 -2112
rect 9 -2237 10 -2115
rect 471 -2116 472 -2112
rect 478 -2116 479 -2112
rect 691 -2116 692 -2112
rect 695 -2116 696 -2112
rect 793 -2237 794 -2115
rect 814 -2116 815 -2112
rect 905 -2116 906 -2112
rect 961 -2116 962 -2112
rect 961 -2237 962 -2115
rect 961 -2116 962 -2112
rect 961 -2237 962 -2115
rect 968 -2116 969 -2112
rect 1115 -2237 1116 -2115
rect 1118 -2116 1119 -2112
rect 1213 -2116 1214 -2112
rect 1262 -2237 1263 -2115
rect 1283 -2116 1284 -2112
rect 30 -2118 31 -2112
rect 44 -2237 45 -2117
rect 51 -2237 52 -2117
rect 660 -2118 661 -2112
rect 667 -2237 668 -2117
rect 737 -2118 738 -2112
rect 765 -2237 766 -2117
rect 835 -2118 836 -2112
rect 891 -2237 892 -2117
rect 1052 -2118 1053 -2112
rect 1139 -2118 1140 -2112
rect 1276 -2118 1277 -2112
rect 75 -2237 76 -2119
rect 709 -2120 710 -2112
rect 814 -2237 815 -2119
rect 898 -2120 899 -2112
rect 905 -2237 906 -2119
rect 954 -2120 955 -2112
rect 985 -2237 986 -2119
rect 1283 -2237 1284 -2119
rect 107 -2122 108 -2112
rect 1192 -2122 1193 -2112
rect 1213 -2237 1214 -2121
rect 1241 -2122 1242 -2112
rect 1276 -2237 1277 -2121
rect 1290 -2122 1291 -2112
rect 107 -2237 108 -2123
rect 411 -2237 412 -2123
rect 450 -2124 451 -2112
rect 1080 -2124 1081 -2112
rect 1192 -2237 1193 -2123
rect 1220 -2124 1221 -2112
rect 1241 -2237 1242 -2123
rect 1255 -2124 1256 -2112
rect 1290 -2237 1291 -2123
rect 1297 -2124 1298 -2112
rect 40 -2237 41 -2125
rect 1220 -2237 1221 -2125
rect 1297 -2237 1298 -2125
rect 1318 -2126 1319 -2112
rect 110 -2128 111 -2112
rect 268 -2128 269 -2112
rect 320 -2128 321 -2112
rect 485 -2128 486 -2112
rect 488 -2128 489 -2112
rect 898 -2237 899 -2127
rect 989 -2237 990 -2127
rect 1010 -2128 1011 -2112
rect 1045 -2237 1046 -2127
rect 1087 -2128 1088 -2112
rect 1206 -2128 1207 -2112
rect 1255 -2237 1256 -2127
rect 131 -2130 132 -2112
rect 156 -2130 157 -2112
rect 170 -2130 171 -2112
rect 177 -2130 178 -2112
rect 184 -2130 185 -2112
rect 334 -2130 335 -2112
rect 345 -2237 346 -2129
rect 555 -2130 556 -2112
rect 579 -2130 580 -2112
rect 681 -2130 682 -2112
rect 695 -2237 696 -2129
rect 982 -2130 983 -2112
rect 992 -2130 993 -2112
rect 1311 -2130 1312 -2112
rect 37 -2132 38 -2112
rect 184 -2237 185 -2131
rect 191 -2132 192 -2112
rect 677 -2237 678 -2131
rect 821 -2237 822 -2131
rect 849 -2132 850 -2112
rect 856 -2132 857 -2112
rect 954 -2237 955 -2131
rect 996 -2132 997 -2112
rect 1087 -2237 1088 -2131
rect 1206 -2237 1207 -2131
rect 1234 -2132 1235 -2112
rect 79 -2134 80 -2112
rect 177 -2237 178 -2133
rect 191 -2237 192 -2133
rect 317 -2134 318 -2112
rect 331 -2134 332 -2112
rect 975 -2237 976 -2133
rect 996 -2237 997 -2133
rect 1031 -2134 1032 -2112
rect 1080 -2237 1081 -2133
rect 1122 -2134 1123 -2112
rect 79 -2237 80 -2135
rect 541 -2136 542 -2112
rect 555 -2237 556 -2135
rect 653 -2136 654 -2112
rect 660 -2237 661 -2135
rect 730 -2136 731 -2112
rect 849 -2237 850 -2135
rect 884 -2136 885 -2112
rect 940 -2136 941 -2112
rect 1010 -2237 1011 -2135
rect 1031 -2237 1032 -2135
rect 1038 -2136 1039 -2112
rect 138 -2237 139 -2137
rect 156 -2237 157 -2137
rect 163 -2237 164 -2137
rect 982 -2237 983 -2137
rect 1003 -2138 1004 -2112
rect 1311 -2237 1312 -2137
rect 170 -2237 171 -2139
rect 621 -2140 622 -2112
rect 628 -2237 629 -2139
rect 1234 -2237 1235 -2139
rect 205 -2142 206 -2112
rect 208 -2156 209 -2141
rect 219 -2142 220 -2112
rect 971 -2142 972 -2112
rect 1003 -2237 1004 -2141
rect 1024 -2142 1025 -2112
rect 1038 -2237 1039 -2141
rect 1094 -2142 1095 -2112
rect 205 -2237 206 -2143
rect 247 -2144 248 -2112
rect 471 -2237 472 -2143
rect 478 -2237 479 -2143
rect 639 -2144 640 -2112
rect 649 -2237 650 -2143
rect 744 -2144 745 -2112
rect 884 -2237 885 -2143
rect 919 -2144 920 -2112
rect 1094 -2237 1095 -2143
rect 1129 -2144 1130 -2112
rect 247 -2237 248 -2145
rect 299 -2237 300 -2145
rect 317 -2237 318 -2145
rect 338 -2146 339 -2112
rect 352 -2146 353 -2112
rect 425 -2237 426 -2145
rect 450 -2237 451 -2145
rect 782 -2146 783 -2112
rect 1129 -2237 1130 -2145
rect 1164 -2146 1165 -2112
rect 5 -2148 6 -2112
rect 352 -2237 353 -2147
rect 373 -2148 374 -2112
rect 681 -2237 682 -2147
rect 702 -2148 703 -2112
rect 856 -2237 857 -2147
rect 1164 -2237 1165 -2147
rect 1185 -2148 1186 -2112
rect 72 -2150 73 -2112
rect 338 -2237 339 -2149
rect 394 -2150 395 -2112
rect 968 -2237 969 -2149
rect 1185 -2237 1186 -2149
rect 1199 -2150 1200 -2112
rect 72 -2237 73 -2151
rect 149 -2152 150 -2112
rect 254 -2152 255 -2112
rect 348 -2152 349 -2112
rect 394 -2237 395 -2151
rect 422 -2152 423 -2112
rect 464 -2152 465 -2112
rect 709 -2237 710 -2151
rect 730 -2237 731 -2151
rect 824 -2152 825 -2112
rect 1199 -2237 1200 -2151
rect 1227 -2152 1228 -2112
rect 2 -2237 3 -2153
rect 149 -2237 150 -2153
rect 261 -2154 262 -2112
rect 268 -2237 269 -2153
rect 310 -2154 311 -2112
rect 373 -2237 374 -2153
rect 397 -2237 398 -2153
rect 453 -2154 454 -2112
rect 464 -2237 465 -2153
rect 530 -2237 531 -2153
rect 541 -2237 542 -2153
rect 590 -2154 591 -2112
rect 597 -2154 598 -2112
rect 737 -2237 738 -2153
rect 744 -2237 745 -2153
rect 947 -2154 948 -2112
rect 1227 -2237 1228 -2153
rect 1248 -2154 1249 -2112
rect 65 -2156 66 -2112
rect 254 -2237 255 -2155
rect 261 -2237 262 -2155
rect 275 -2156 276 -2112
rect 296 -2156 297 -2112
rect 310 -2237 311 -2155
rect 404 -2237 405 -2155
rect 688 -2156 689 -2112
rect 702 -2237 703 -2155
rect 723 -2156 724 -2112
rect 768 -2237 769 -2155
rect 835 -2237 836 -2155
rect 1248 -2237 1249 -2155
rect 1269 -2156 1270 -2112
rect 65 -2237 66 -2157
rect 86 -2158 87 -2112
rect 275 -2237 276 -2157
rect 303 -2158 304 -2112
rect 453 -2237 454 -2157
rect 807 -2158 808 -2112
rect 1269 -2237 1270 -2157
rect 1304 -2158 1305 -2112
rect 86 -2237 87 -2159
rect 226 -2160 227 -2112
rect 240 -2160 241 -2112
rect 303 -2237 304 -2159
rect 485 -2237 486 -2159
rect 527 -2160 528 -2112
rect 548 -2160 549 -2112
rect 947 -2237 948 -2159
rect 1304 -2237 1305 -2159
rect 1325 -2160 1326 -2112
rect 198 -2162 199 -2112
rect 226 -2237 227 -2161
rect 240 -2237 241 -2161
rect 359 -2162 360 -2112
rect 443 -2162 444 -2112
rect 548 -2237 549 -2161
rect 590 -2237 591 -2161
rect 716 -2162 717 -2112
rect 723 -2237 724 -2161
rect 758 -2162 759 -2112
rect 772 -2162 773 -2112
rect 919 -2237 920 -2161
rect 198 -2237 199 -2163
rect 387 -2164 388 -2112
rect 436 -2164 437 -2112
rect 443 -2237 444 -2163
rect 499 -2164 500 -2112
rect 1178 -2164 1179 -2112
rect 128 -2166 129 -2112
rect 1178 -2237 1179 -2165
rect 114 -2168 115 -2112
rect 128 -2237 129 -2167
rect 219 -2237 220 -2167
rect 527 -2237 528 -2167
rect 576 -2168 577 -2112
rect 772 -2237 773 -2167
rect 807 -2237 808 -2167
rect 1122 -2237 1123 -2167
rect 296 -2237 297 -2169
rect 331 -2237 332 -2169
rect 359 -2237 360 -2169
rect 894 -2170 895 -2112
rect 324 -2172 325 -2112
rect 387 -2237 388 -2171
rect 415 -2172 416 -2112
rect 436 -2237 437 -2171
rect 499 -2237 500 -2171
rect 810 -2237 811 -2171
rect 212 -2174 213 -2112
rect 415 -2237 416 -2173
rect 502 -2174 503 -2112
rect 779 -2237 780 -2173
rect 212 -2237 213 -2175
rect 492 -2176 493 -2112
rect 520 -2176 521 -2112
rect 639 -2237 640 -2175
rect 653 -2237 654 -2175
rect 817 -2176 818 -2112
rect 324 -2237 325 -2177
rect 401 -2178 402 -2112
rect 492 -2237 493 -2177
rect 926 -2178 927 -2112
rect 401 -2237 402 -2179
rect 1024 -2237 1025 -2179
rect 523 -2237 524 -2181
rect 940 -2237 941 -2181
rect 576 -2237 577 -2183
rect 674 -2184 675 -2112
rect 716 -2237 717 -2183
rect 751 -2184 752 -2112
rect 758 -2237 759 -2183
rect 786 -2184 787 -2112
rect 597 -2237 598 -2185
rect 618 -2186 619 -2112
rect 621 -2237 622 -2185
rect 828 -2186 829 -2112
rect 506 -2188 507 -2112
rect 618 -2237 619 -2187
rect 632 -2188 633 -2112
rect 926 -2237 927 -2187
rect 93 -2190 94 -2112
rect 506 -2237 507 -2189
rect 611 -2190 612 -2112
rect 688 -2237 689 -2189
rect 751 -2237 752 -2189
rect 800 -2190 801 -2112
rect 828 -2237 829 -2189
rect 863 -2190 864 -2112
rect 93 -2237 94 -2191
rect 282 -2192 283 -2112
rect 583 -2192 584 -2112
rect 611 -2237 612 -2191
rect 786 -2237 787 -2191
rect 1136 -2192 1137 -2112
rect 117 -2237 118 -2193
rect 632 -2237 633 -2193
rect 800 -2237 801 -2193
rect 842 -2194 843 -2112
rect 863 -2237 864 -2193
rect 912 -2194 913 -2112
rect 1136 -2237 1137 -2193
rect 1157 -2194 1158 -2112
rect 282 -2237 283 -2195
rect 513 -2196 514 -2112
rect 534 -2196 535 -2112
rect 583 -2237 584 -2195
rect 842 -2237 843 -2195
rect 877 -2196 878 -2112
rect 912 -2237 913 -2195
rect 933 -2196 934 -2112
rect 1017 -2196 1018 -2112
rect 1157 -2237 1158 -2195
rect 37 -2237 38 -2197
rect 877 -2237 878 -2197
rect 933 -2237 934 -2197
rect 1108 -2198 1109 -2112
rect 380 -2200 381 -2112
rect 513 -2237 514 -2199
rect 534 -2237 535 -2199
rect 569 -2200 570 -2112
rect 1017 -2237 1018 -2199
rect 1059 -2200 1060 -2112
rect 1108 -2237 1109 -2199
rect 1150 -2200 1151 -2112
rect 135 -2202 136 -2112
rect 380 -2237 381 -2201
rect 520 -2237 521 -2201
rect 1059 -2237 1060 -2201
rect 135 -2237 136 -2203
rect 366 -2204 367 -2112
rect 569 -2237 570 -2203
rect 625 -2204 626 -2112
rect 16 -2206 17 -2112
rect 366 -2237 367 -2205
rect 562 -2206 563 -2112
rect 625 -2237 626 -2205
rect 16 -2237 17 -2207
rect 457 -2208 458 -2112
rect 562 -2237 563 -2207
rect 604 -2208 605 -2112
rect 58 -2210 59 -2112
rect 457 -2237 458 -2209
rect 604 -2237 605 -2209
rect 646 -2210 647 -2112
rect 58 -2237 59 -2211
rect 142 -2212 143 -2112
rect 152 -2237 153 -2211
rect 1150 -2237 1151 -2211
rect 100 -2214 101 -2112
rect 646 -2237 647 -2213
rect 100 -2237 101 -2215
rect 289 -2216 290 -2112
rect 121 -2218 122 -2112
rect 142 -2237 143 -2217
rect 289 -2237 290 -2217
rect 429 -2218 430 -2112
rect 23 -2220 24 -2112
rect 429 -2237 430 -2219
rect 23 -2237 24 -2221
rect 26 -2237 27 -2221
rect 121 -2237 122 -2221
rect 408 -2222 409 -2112
rect 408 -2237 409 -2223
rect 1066 -2224 1067 -2112
rect 1066 -2237 1067 -2225
rect 1101 -2226 1102 -2112
rect 1101 -2237 1102 -2227
rect 1143 -2228 1144 -2112
rect 1143 -2237 1144 -2229
rect 1171 -2230 1172 -2112
rect 1073 -2232 1074 -2112
rect 1171 -2237 1172 -2231
rect 870 -2234 871 -2112
rect 1073 -2237 1074 -2233
rect 870 -2237 871 -2235
rect 1052 -2237 1053 -2235
rect 5 -2362 6 -2246
rect 44 -2247 45 -2245
rect 61 -2362 62 -2246
rect 492 -2247 493 -2245
rect 516 -2362 517 -2246
rect 726 -2362 727 -2246
rect 747 -2362 748 -2246
rect 1087 -2247 1088 -2245
rect 23 -2249 24 -2245
rect 1024 -2249 1025 -2245
rect 1034 -2362 1035 -2248
rect 1290 -2249 1291 -2245
rect 23 -2362 24 -2250
rect 401 -2251 402 -2245
rect 408 -2251 409 -2245
rect 415 -2251 416 -2245
rect 425 -2251 426 -2245
rect 688 -2251 689 -2245
rect 761 -2362 762 -2250
rect 856 -2251 857 -2245
rect 870 -2251 871 -2245
rect 1234 -2251 1235 -2245
rect 33 -2253 34 -2245
rect 198 -2253 199 -2245
rect 205 -2253 206 -2245
rect 338 -2253 339 -2245
rect 387 -2253 388 -2245
rect 523 -2253 524 -2245
rect 527 -2253 528 -2245
rect 737 -2253 738 -2245
rect 810 -2253 811 -2245
rect 961 -2253 962 -2245
rect 982 -2253 983 -2245
rect 1276 -2253 1277 -2245
rect 9 -2255 10 -2245
rect 198 -2362 199 -2254
rect 205 -2362 206 -2254
rect 373 -2255 374 -2245
rect 387 -2362 388 -2254
rect 422 -2255 423 -2245
rect 520 -2255 521 -2245
rect 562 -2255 563 -2245
rect 579 -2362 580 -2254
rect 968 -2255 969 -2245
rect 982 -2362 983 -2254
rect 985 -2255 986 -2245
rect 1024 -2362 1025 -2254
rect 1094 -2255 1095 -2245
rect 9 -2362 10 -2256
rect 359 -2257 360 -2245
rect 411 -2257 412 -2245
rect 464 -2257 465 -2245
rect 527 -2362 528 -2256
rect 933 -2257 934 -2245
rect 961 -2362 962 -2256
rect 1017 -2257 1018 -2245
rect 1094 -2362 1095 -2256
rect 1150 -2257 1151 -2245
rect 37 -2259 38 -2245
rect 975 -2259 976 -2245
rect 1017 -2362 1018 -2258
rect 1080 -2259 1081 -2245
rect 1150 -2362 1151 -2258
rect 1220 -2259 1221 -2245
rect 37 -2362 38 -2260
rect 341 -2261 342 -2245
rect 359 -2362 360 -2260
rect 485 -2261 486 -2245
rect 530 -2261 531 -2245
rect 926 -2261 927 -2245
rect 933 -2362 934 -2260
rect 1059 -2261 1060 -2245
rect 1080 -2362 1081 -2260
rect 1297 -2261 1298 -2245
rect 40 -2263 41 -2245
rect 352 -2263 353 -2245
rect 464 -2362 465 -2262
rect 849 -2263 850 -2245
rect 856 -2362 857 -2262
rect 1010 -2263 1011 -2245
rect 1059 -2362 1060 -2262
rect 1122 -2263 1123 -2245
rect 40 -2362 41 -2264
rect 926 -2362 927 -2264
rect 975 -2362 976 -2264
rect 1269 -2265 1270 -2245
rect 44 -2362 45 -2266
rect 380 -2267 381 -2245
rect 485 -2362 486 -2266
rect 513 -2267 514 -2245
rect 548 -2267 549 -2245
rect 688 -2362 689 -2266
rect 695 -2267 696 -2245
rect 849 -2362 850 -2266
rect 870 -2362 871 -2266
rect 940 -2267 941 -2245
rect 1122 -2362 1123 -2266
rect 1192 -2267 1193 -2245
rect 79 -2269 80 -2245
rect 415 -2362 416 -2268
rect 548 -2362 549 -2268
rect 604 -2269 605 -2245
rect 625 -2362 626 -2268
rect 639 -2269 640 -2245
rect 674 -2362 675 -2268
rect 772 -2269 773 -2245
rect 873 -2269 874 -2245
rect 1031 -2269 1032 -2245
rect 1192 -2362 1193 -2268
rect 1241 -2269 1242 -2245
rect 16 -2271 17 -2245
rect 79 -2362 80 -2270
rect 86 -2271 87 -2245
rect 296 -2271 297 -2245
rect 306 -2362 307 -2270
rect 408 -2362 409 -2270
rect 492 -2362 493 -2270
rect 1031 -2362 1032 -2270
rect 1129 -2271 1130 -2245
rect 1241 -2362 1242 -2270
rect 16 -2362 17 -2272
rect 317 -2273 318 -2245
rect 320 -2362 321 -2272
rect 1234 -2362 1235 -2272
rect 86 -2362 87 -2274
rect 723 -2275 724 -2245
rect 737 -2362 738 -2274
rect 744 -2275 745 -2245
rect 772 -2362 773 -2274
rect 800 -2275 801 -2245
rect 96 -2362 97 -2276
rect 618 -2277 619 -2245
rect 628 -2277 629 -2245
rect 968 -2362 969 -2276
rect 100 -2279 101 -2245
rect 114 -2279 115 -2245
rect 117 -2279 118 -2245
rect 1178 -2279 1179 -2245
rect 100 -2362 101 -2280
rect 345 -2281 346 -2245
rect 352 -2362 353 -2280
rect 478 -2281 479 -2245
rect 513 -2362 514 -2280
rect 1129 -2362 1130 -2280
rect 1178 -2362 1179 -2280
rect 1255 -2281 1256 -2245
rect 114 -2362 115 -2282
rect 191 -2283 192 -2245
rect 240 -2283 241 -2245
rect 520 -2362 521 -2282
rect 558 -2283 559 -2245
rect 681 -2283 682 -2245
rect 695 -2362 696 -2282
rect 793 -2283 794 -2245
rect 800 -2362 801 -2282
rect 814 -2283 815 -2245
rect 121 -2285 122 -2245
rect 744 -2362 745 -2284
rect 793 -2362 794 -2284
rect 810 -2362 811 -2284
rect 814 -2362 815 -2284
rect 877 -2285 878 -2245
rect 121 -2362 122 -2286
rect 450 -2287 451 -2245
rect 555 -2287 556 -2245
rect 681 -2362 682 -2286
rect 877 -2362 878 -2286
rect 947 -2287 948 -2245
rect 149 -2289 150 -2245
rect 919 -2289 920 -2245
rect 947 -2362 948 -2288
rect 1045 -2289 1046 -2245
rect 149 -2362 150 -2290
rect 436 -2291 437 -2245
rect 450 -2362 451 -2290
rect 583 -2291 584 -2245
rect 593 -2362 594 -2290
rect 835 -2291 836 -2245
rect 919 -2362 920 -2290
rect 989 -2291 990 -2245
rect 1045 -2362 1046 -2290
rect 1304 -2291 1305 -2245
rect 152 -2362 153 -2292
rect 807 -2293 808 -2245
rect 989 -2362 990 -2292
rect 1066 -2293 1067 -2245
rect 156 -2295 157 -2245
rect 296 -2362 297 -2294
rect 331 -2295 332 -2245
rect 940 -2362 941 -2294
rect 1066 -2362 1067 -2294
rect 1164 -2295 1165 -2245
rect 2 -2297 3 -2245
rect 331 -2362 332 -2296
rect 341 -2362 342 -2296
rect 457 -2297 458 -2245
rect 562 -2362 563 -2296
rect 660 -2297 661 -2245
rect 677 -2297 678 -2245
rect 1136 -2297 1137 -2245
rect 2 -2362 3 -2298
rect 478 -2362 479 -2298
rect 569 -2299 570 -2245
rect 583 -2362 584 -2298
rect 604 -2362 605 -2298
rect 702 -2299 703 -2245
rect 786 -2299 787 -2245
rect 835 -2362 836 -2298
rect 107 -2301 108 -2245
rect 457 -2362 458 -2300
rect 471 -2301 472 -2245
rect 569 -2362 570 -2300
rect 611 -2301 612 -2245
rect 618 -2362 619 -2300
rect 635 -2362 636 -2300
rect 758 -2301 759 -2245
rect 807 -2362 808 -2300
rect 1003 -2301 1004 -2245
rect 107 -2362 108 -2302
rect 128 -2303 129 -2245
rect 156 -2362 157 -2302
rect 184 -2303 185 -2245
rect 191 -2362 192 -2302
rect 289 -2303 290 -2245
rect 380 -2362 381 -2302
rect 576 -2303 577 -2245
rect 611 -2362 612 -2302
rect 632 -2303 633 -2245
rect 639 -2362 640 -2302
rect 709 -2303 710 -2245
rect 758 -2362 759 -2302
rect 1171 -2303 1172 -2245
rect 75 -2305 76 -2245
rect 632 -2362 633 -2304
rect 646 -2305 647 -2245
rect 1164 -2362 1165 -2304
rect 128 -2362 129 -2306
rect 394 -2307 395 -2245
rect 471 -2362 472 -2306
rect 506 -2307 507 -2245
rect 576 -2362 577 -2306
rect 1220 -2362 1221 -2306
rect 51 -2309 52 -2245
rect 394 -2362 395 -2308
rect 499 -2309 500 -2245
rect 506 -2362 507 -2308
rect 597 -2309 598 -2245
rect 646 -2362 647 -2308
rect 660 -2362 661 -2308
rect 1283 -2309 1284 -2245
rect 51 -2362 52 -2310
rect 138 -2311 139 -2245
rect 163 -2311 164 -2245
rect 289 -2362 290 -2310
rect 338 -2362 339 -2310
rect 1171 -2362 1172 -2310
rect 138 -2362 139 -2312
rect 1087 -2362 1088 -2312
rect 163 -2362 164 -2314
rect 404 -2315 405 -2245
rect 499 -2362 500 -2314
rect 534 -2315 535 -2245
rect 590 -2315 591 -2245
rect 597 -2362 598 -2314
rect 702 -2362 703 -2314
rect 751 -2315 752 -2245
rect 1003 -2362 1004 -2314
rect 1206 -2315 1207 -2245
rect 177 -2317 178 -2245
rect 345 -2362 346 -2316
rect 534 -2362 535 -2316
rect 863 -2317 864 -2245
rect 1206 -2362 1207 -2316
rect 1248 -2317 1249 -2245
rect 170 -2319 171 -2245
rect 177 -2362 178 -2318
rect 184 -2362 185 -2318
rect 233 -2319 234 -2245
rect 254 -2319 255 -2245
rect 373 -2362 374 -2318
rect 590 -2362 591 -2318
rect 1136 -2362 1137 -2318
rect 1248 -2362 1249 -2318
rect 1311 -2319 1312 -2245
rect 93 -2321 94 -2245
rect 254 -2362 255 -2320
rect 261 -2321 262 -2245
rect 401 -2362 402 -2320
rect 709 -2362 710 -2320
rect 716 -2321 717 -2245
rect 751 -2362 752 -2320
rect 842 -2321 843 -2245
rect 863 -2362 864 -2320
rect 954 -2321 955 -2245
rect 65 -2323 66 -2245
rect 93 -2362 94 -2322
rect 170 -2362 171 -2322
rect 317 -2362 318 -2322
rect 397 -2323 398 -2245
rect 842 -2362 843 -2322
rect 954 -2362 955 -2322
rect 1108 -2323 1109 -2245
rect 30 -2325 31 -2245
rect 65 -2362 66 -2324
rect 219 -2325 220 -2245
rect 240 -2362 241 -2324
rect 261 -2362 262 -2324
rect 555 -2362 556 -2324
rect 716 -2362 717 -2324
rect 765 -2325 766 -2245
rect 1108 -2362 1109 -2324
rect 1185 -2325 1186 -2245
rect 30 -2362 31 -2326
rect 425 -2362 426 -2326
rect 1185 -2362 1186 -2326
rect 1227 -2327 1228 -2245
rect 135 -2329 136 -2245
rect 765 -2362 766 -2328
rect 891 -2329 892 -2245
rect 1227 -2362 1228 -2328
rect 135 -2362 136 -2330
rect 366 -2331 367 -2245
rect 397 -2362 398 -2330
rect 730 -2331 731 -2245
rect 891 -2362 892 -2330
rect 996 -2331 997 -2245
rect 219 -2362 220 -2332
rect 324 -2333 325 -2245
rect 366 -2362 367 -2332
rect 541 -2333 542 -2245
rect 730 -2362 731 -2332
rect 821 -2333 822 -2245
rect 996 -2362 997 -2332
rect 1073 -2333 1074 -2245
rect 226 -2335 227 -2245
rect 786 -2362 787 -2334
rect 821 -2362 822 -2334
rect 884 -2335 885 -2245
rect 1073 -2362 1074 -2334
rect 1143 -2335 1144 -2245
rect 142 -2337 143 -2245
rect 226 -2362 227 -2336
rect 233 -2362 234 -2336
rect 268 -2337 269 -2245
rect 282 -2337 283 -2245
rect 663 -2362 664 -2336
rect 779 -2337 780 -2245
rect 884 -2362 885 -2336
rect 1143 -2362 1144 -2336
rect 1199 -2337 1200 -2245
rect 142 -2362 143 -2338
rect 828 -2339 829 -2245
rect 268 -2362 269 -2340
rect 310 -2341 311 -2245
rect 324 -2362 325 -2340
rect 443 -2341 444 -2245
rect 541 -2362 542 -2340
rect 653 -2341 654 -2245
rect 779 -2362 780 -2340
rect 912 -2341 913 -2245
rect 275 -2343 276 -2245
rect 310 -2362 311 -2342
rect 443 -2362 444 -2342
rect 453 -2343 454 -2245
rect 621 -2343 622 -2245
rect 1199 -2362 1200 -2342
rect 275 -2362 276 -2344
rect 429 -2345 430 -2245
rect 653 -2362 654 -2344
rect 667 -2345 668 -2245
rect 828 -2362 829 -2344
rect 898 -2345 899 -2245
rect 912 -2362 913 -2344
rect 1052 -2345 1053 -2245
rect 72 -2347 73 -2245
rect 667 -2362 668 -2346
rect 898 -2362 899 -2346
rect 905 -2347 906 -2245
rect 72 -2362 73 -2348
rect 247 -2349 248 -2245
rect 282 -2362 283 -2348
rect 299 -2349 300 -2245
rect 436 -2362 437 -2348
rect 1052 -2362 1053 -2348
rect 58 -2351 59 -2245
rect 247 -2362 248 -2350
rect 905 -2362 906 -2350
rect 1115 -2351 1116 -2245
rect 58 -2362 59 -2352
rect 1010 -2362 1011 -2352
rect 1038 -2353 1039 -2245
rect 1115 -2362 1116 -2352
rect 212 -2355 213 -2245
rect 429 -2362 430 -2354
rect 1038 -2362 1039 -2354
rect 1101 -2355 1102 -2245
rect 212 -2362 213 -2356
rect 303 -2357 304 -2245
rect 1101 -2362 1102 -2356
rect 1157 -2357 1158 -2245
rect 1157 -2362 1158 -2358
rect 1213 -2359 1214 -2245
rect 1213 -2362 1214 -2360
rect 1262 -2361 1263 -2245
rect 9 -2372 10 -2370
rect 376 -2459 377 -2371
rect 394 -2372 395 -2370
rect 1234 -2372 1235 -2370
rect 23 -2374 24 -2370
rect 341 -2374 342 -2370
rect 352 -2374 353 -2370
rect 436 -2374 437 -2370
rect 446 -2459 447 -2373
rect 779 -2374 780 -2370
rect 796 -2459 797 -2373
rect 954 -2374 955 -2370
rect 1031 -2459 1032 -2373
rect 1073 -2374 1074 -2370
rect 1104 -2459 1105 -2373
rect 1115 -2374 1116 -2370
rect 30 -2376 31 -2370
rect 201 -2459 202 -2375
rect 303 -2376 304 -2370
rect 842 -2376 843 -2370
rect 849 -2376 850 -2370
rect 919 -2376 920 -2370
rect 954 -2459 955 -2375
rect 1045 -2376 1046 -2370
rect 1073 -2459 1074 -2375
rect 1199 -2376 1200 -2370
rect 37 -2378 38 -2370
rect 296 -2378 297 -2370
rect 303 -2459 304 -2377
rect 425 -2378 426 -2370
rect 464 -2378 465 -2370
rect 758 -2378 759 -2370
rect 779 -2459 780 -2377
rect 1010 -2378 1011 -2370
rect 1034 -2378 1035 -2370
rect 1178 -2378 1179 -2370
rect 40 -2380 41 -2370
rect 940 -2380 941 -2370
rect 1010 -2459 1011 -2379
rect 1059 -2380 1060 -2370
rect 54 -2382 55 -2370
rect 254 -2382 255 -2370
rect 310 -2382 311 -2370
rect 310 -2459 311 -2381
rect 310 -2382 311 -2370
rect 310 -2459 311 -2381
rect 320 -2382 321 -2370
rect 786 -2382 787 -2370
rect 807 -2382 808 -2370
rect 1143 -2382 1144 -2370
rect 61 -2384 62 -2370
rect 569 -2384 570 -2370
rect 576 -2384 577 -2370
rect 905 -2384 906 -2370
rect 908 -2459 909 -2383
rect 1220 -2384 1221 -2370
rect 65 -2386 66 -2370
rect 65 -2459 66 -2385
rect 65 -2386 66 -2370
rect 65 -2459 66 -2385
rect 72 -2386 73 -2370
rect 513 -2386 514 -2370
rect 520 -2386 521 -2370
rect 810 -2386 811 -2370
rect 842 -2459 843 -2385
rect 1108 -2386 1109 -2370
rect 72 -2459 73 -2387
rect 170 -2388 171 -2370
rect 184 -2388 185 -2370
rect 306 -2388 307 -2370
rect 338 -2459 339 -2387
rect 443 -2388 444 -2370
rect 485 -2388 486 -2370
rect 849 -2459 850 -2387
rect 898 -2388 899 -2370
rect 1013 -2459 1014 -2387
rect 1059 -2459 1060 -2387
rect 1080 -2388 1081 -2370
rect 79 -2390 80 -2370
rect 149 -2459 150 -2389
rect 163 -2390 164 -2370
rect 296 -2459 297 -2389
rect 359 -2390 360 -2370
rect 362 -2416 363 -2389
rect 366 -2390 367 -2370
rect 516 -2390 517 -2370
rect 520 -2459 521 -2389
rect 593 -2390 594 -2370
rect 614 -2459 615 -2389
rect 863 -2390 864 -2370
rect 898 -2459 899 -2389
rect 1157 -2390 1158 -2370
rect 44 -2392 45 -2370
rect 79 -2459 80 -2391
rect 86 -2392 87 -2370
rect 366 -2459 367 -2391
rect 394 -2459 395 -2391
rect 471 -2392 472 -2370
rect 516 -2459 517 -2391
rect 1164 -2392 1165 -2370
rect 86 -2459 87 -2393
rect 282 -2394 283 -2370
rect 359 -2459 360 -2393
rect 408 -2394 409 -2370
rect 422 -2394 423 -2370
rect 688 -2394 689 -2370
rect 723 -2394 724 -2370
rect 772 -2394 773 -2370
rect 786 -2459 787 -2393
rect 852 -2394 853 -2370
rect 905 -2459 906 -2393
rect 1241 -2394 1242 -2370
rect 93 -2396 94 -2370
rect 422 -2459 423 -2395
rect 450 -2396 451 -2370
rect 863 -2459 864 -2395
rect 919 -2459 920 -2395
rect 996 -2396 997 -2370
rect 1080 -2459 1081 -2395
rect 1136 -2396 1137 -2370
rect 93 -2459 94 -2397
rect 397 -2398 398 -2370
rect 450 -2459 451 -2397
rect 870 -2398 871 -2370
rect 884 -2398 885 -2370
rect 996 -2459 997 -2397
rect 100 -2400 101 -2370
rect 744 -2400 745 -2370
rect 751 -2400 752 -2370
rect 758 -2459 759 -2399
rect 765 -2400 766 -2370
rect 807 -2459 808 -2399
rect 870 -2459 871 -2399
rect 912 -2400 913 -2370
rect 940 -2459 941 -2399
rect 1122 -2400 1123 -2370
rect 100 -2459 101 -2401
rect 142 -2402 143 -2370
rect 184 -2459 185 -2401
rect 562 -2402 563 -2370
rect 569 -2459 570 -2401
rect 625 -2402 626 -2370
rect 635 -2402 636 -2370
rect 702 -2402 703 -2370
rect 709 -2402 710 -2370
rect 884 -2459 885 -2401
rect 912 -2459 913 -2401
rect 1171 -2402 1172 -2370
rect 107 -2404 108 -2370
rect 170 -2459 171 -2403
rect 198 -2404 199 -2370
rect 439 -2404 440 -2370
rect 457 -2404 458 -2370
rect 485 -2459 486 -2403
rect 548 -2404 549 -2370
rect 576 -2459 577 -2403
rect 590 -2404 591 -2370
rect 653 -2404 654 -2370
rect 660 -2404 661 -2370
rect 1227 -2404 1228 -2370
rect 107 -2459 108 -2405
rect 597 -2406 598 -2370
rect 611 -2406 612 -2370
rect 653 -2459 654 -2405
rect 663 -2459 664 -2405
rect 1066 -2406 1067 -2370
rect 58 -2408 59 -2370
rect 597 -2459 598 -2407
rect 646 -2408 647 -2370
rect 744 -2459 745 -2407
rect 751 -2459 752 -2407
rect 891 -2408 892 -2370
rect 961 -2408 962 -2370
rect 1108 -2459 1109 -2407
rect 58 -2459 59 -2409
rect 247 -2410 248 -2370
rect 261 -2410 262 -2370
rect 590 -2459 591 -2409
rect 646 -2459 647 -2409
rect 933 -2410 934 -2370
rect 1066 -2459 1067 -2409
rect 1129 -2410 1130 -2370
rect 114 -2412 115 -2370
rect 114 -2459 115 -2411
rect 114 -2412 115 -2370
rect 114 -2459 115 -2411
rect 121 -2412 122 -2370
rect 254 -2459 255 -2411
rect 261 -2459 262 -2411
rect 506 -2412 507 -2370
rect 555 -2459 556 -2411
rect 730 -2412 731 -2370
rect 765 -2459 766 -2411
rect 975 -2412 976 -2370
rect 1129 -2459 1130 -2411
rect 1248 -2412 1249 -2370
rect 124 -2459 125 -2413
rect 968 -2414 969 -2370
rect 128 -2416 129 -2370
rect 163 -2459 164 -2415
rect 198 -2459 199 -2415
rect 226 -2416 227 -2370
rect 247 -2459 248 -2415
rect 324 -2416 325 -2370
rect 408 -2459 409 -2415
rect 415 -2416 416 -2370
rect 660 -2459 661 -2415
rect 667 -2416 668 -2370
rect 702 -2459 703 -2415
rect 709 -2459 710 -2415
rect 989 -2416 990 -2370
rect 128 -2459 129 -2417
rect 138 -2418 139 -2370
rect 142 -2459 143 -2417
rect 317 -2418 318 -2370
rect 387 -2418 388 -2370
rect 625 -2459 626 -2417
rect 667 -2459 668 -2417
rect 828 -2418 829 -2370
rect 877 -2418 878 -2370
rect 933 -2459 934 -2417
rect 989 -2459 990 -2417
rect 1192 -2418 1193 -2370
rect 131 -2459 132 -2419
rect 548 -2459 549 -2419
rect 558 -2420 559 -2370
rect 639 -2420 640 -2370
rect 674 -2420 675 -2370
rect 975 -2459 976 -2419
rect 1192 -2459 1193 -2419
rect 1206 -2420 1207 -2370
rect 135 -2422 136 -2370
rect 135 -2459 136 -2421
rect 135 -2422 136 -2370
rect 135 -2459 136 -2421
rect 226 -2459 227 -2421
rect 331 -2422 332 -2370
rect 380 -2422 381 -2370
rect 674 -2459 675 -2421
rect 681 -2422 682 -2370
rect 723 -2459 724 -2421
rect 726 -2422 727 -2370
rect 961 -2459 962 -2421
rect 51 -2424 52 -2370
rect 380 -2459 381 -2423
rect 387 -2459 388 -2423
rect 429 -2424 430 -2370
rect 439 -2459 440 -2423
rect 761 -2424 762 -2370
rect 772 -2459 773 -2423
rect 856 -2424 857 -2370
rect 877 -2459 878 -2423
rect 1017 -2424 1018 -2370
rect 275 -2426 276 -2370
rect 726 -2459 727 -2425
rect 814 -2426 815 -2370
rect 891 -2459 892 -2425
rect 1017 -2459 1018 -2425
rect 1213 -2426 1214 -2370
rect 212 -2428 213 -2370
rect 275 -2459 276 -2427
rect 282 -2459 283 -2427
rect 401 -2428 402 -2370
rect 415 -2459 416 -2427
rect 464 -2459 465 -2427
rect 471 -2459 472 -2427
rect 604 -2428 605 -2370
rect 611 -2459 612 -2427
rect 968 -2459 969 -2427
rect 212 -2459 213 -2429
rect 240 -2430 241 -2370
rect 289 -2430 290 -2370
rect 324 -2459 325 -2429
rect 331 -2459 332 -2429
rect 373 -2430 374 -2370
rect 401 -2459 402 -2429
rect 513 -2459 514 -2429
rect 579 -2430 580 -2370
rect 730 -2459 731 -2429
rect 814 -2459 815 -2429
rect 1094 -2430 1095 -2370
rect 177 -2432 178 -2370
rect 240 -2459 241 -2431
rect 289 -2459 290 -2431
rect 352 -2459 353 -2431
rect 373 -2459 374 -2431
rect 828 -2459 829 -2431
rect 856 -2459 857 -2431
rect 1038 -2432 1039 -2370
rect 156 -2434 157 -2370
rect 177 -2459 178 -2433
rect 317 -2459 318 -2433
rect 345 -2434 346 -2370
rect 429 -2459 430 -2433
rect 534 -2434 535 -2370
rect 604 -2459 605 -2433
rect 1087 -2434 1088 -2370
rect 156 -2459 157 -2435
rect 233 -2436 234 -2370
rect 345 -2459 346 -2435
rect 467 -2459 468 -2435
rect 478 -2436 479 -2370
rect 562 -2459 563 -2435
rect 618 -2436 619 -2370
rect 681 -2459 682 -2435
rect 688 -2459 689 -2435
rect 926 -2436 927 -2370
rect 982 -2436 983 -2370
rect 1087 -2459 1088 -2435
rect 233 -2459 234 -2437
rect 527 -2438 528 -2370
rect 534 -2459 535 -2437
rect 632 -2438 633 -2370
rect 639 -2459 640 -2437
rect 737 -2438 738 -2370
rect 926 -2459 927 -2437
rect 1003 -2438 1004 -2370
rect 457 -2459 458 -2439
rect 492 -2440 493 -2370
rect 499 -2440 500 -2370
rect 506 -2459 507 -2439
rect 527 -2459 528 -2439
rect 695 -2440 696 -2370
rect 737 -2459 738 -2439
rect 943 -2459 944 -2439
rect 982 -2459 983 -2439
rect 1101 -2440 1102 -2370
rect 478 -2459 479 -2441
rect 583 -2442 584 -2370
rect 618 -2459 619 -2441
rect 716 -2442 717 -2370
rect 821 -2442 822 -2370
rect 1003 -2459 1004 -2441
rect 1094 -2459 1095 -2441
rect 1101 -2459 1102 -2441
rect 268 -2444 269 -2370
rect 583 -2459 584 -2443
rect 632 -2459 633 -2443
rect 800 -2444 801 -2370
rect 821 -2459 822 -2443
rect 1052 -2444 1053 -2370
rect 205 -2446 206 -2370
rect 268 -2459 269 -2445
rect 492 -2459 493 -2445
rect 793 -2446 794 -2370
rect 205 -2459 206 -2447
rect 219 -2448 220 -2370
rect 499 -2459 500 -2447
rect 572 -2459 573 -2447
rect 695 -2459 696 -2447
rect 1150 -2448 1151 -2370
rect 191 -2450 192 -2370
rect 219 -2459 220 -2449
rect 541 -2450 542 -2370
rect 800 -2459 801 -2449
rect 16 -2452 17 -2370
rect 191 -2459 192 -2451
rect 443 -2459 444 -2451
rect 541 -2459 542 -2451
rect 716 -2459 717 -2451
rect 835 -2452 836 -2370
rect 835 -2459 836 -2453
rect 1024 -2454 1025 -2370
rect 947 -2456 948 -2370
rect 1024 -2459 1025 -2455
rect 947 -2459 948 -2457
rect 1185 -2458 1186 -2370
rect 58 -2469 59 -2467
rect 460 -2542 461 -2468
rect 471 -2469 472 -2467
rect 523 -2542 524 -2468
rect 530 -2542 531 -2468
rect 583 -2469 584 -2467
rect 625 -2469 626 -2467
rect 866 -2542 867 -2468
rect 961 -2469 962 -2467
rect 1101 -2469 1102 -2467
rect 1108 -2469 1109 -2467
rect 1143 -2542 1144 -2468
rect 1185 -2542 1186 -2468
rect 1192 -2469 1193 -2467
rect 65 -2471 66 -2467
rect 352 -2471 353 -2467
rect 366 -2471 367 -2467
rect 586 -2542 587 -2470
rect 625 -2542 626 -2470
rect 821 -2471 822 -2467
rect 828 -2471 829 -2467
rect 870 -2471 871 -2467
rect 1013 -2471 1014 -2467
rect 1129 -2471 1130 -2467
rect 72 -2473 73 -2467
rect 131 -2473 132 -2467
rect 135 -2473 136 -2467
rect 135 -2542 136 -2472
rect 135 -2473 136 -2467
rect 135 -2542 136 -2472
rect 149 -2473 150 -2467
rect 352 -2542 353 -2472
rect 366 -2542 367 -2472
rect 604 -2473 605 -2467
rect 639 -2473 640 -2467
rect 642 -2505 643 -2472
rect 674 -2473 675 -2467
rect 758 -2473 759 -2467
rect 793 -2473 794 -2467
rect 807 -2473 808 -2467
rect 828 -2542 829 -2472
rect 856 -2473 857 -2467
rect 863 -2473 864 -2467
rect 870 -2542 871 -2472
rect 1024 -2473 1025 -2467
rect 1104 -2473 1105 -2467
rect 79 -2475 80 -2467
rect 471 -2542 472 -2474
rect 478 -2475 479 -2467
rect 695 -2475 696 -2467
rect 723 -2475 724 -2467
rect 947 -2475 948 -2467
rect 1038 -2542 1039 -2474
rect 1073 -2475 1074 -2467
rect 1087 -2475 1088 -2467
rect 1178 -2542 1179 -2474
rect 86 -2477 87 -2467
rect 166 -2477 167 -2467
rect 191 -2477 192 -2467
rect 691 -2542 692 -2476
rect 740 -2542 741 -2476
rect 877 -2477 878 -2467
rect 926 -2477 927 -2467
rect 947 -2542 948 -2476
rect 1052 -2542 1053 -2476
rect 1059 -2477 1060 -2467
rect 1094 -2477 1095 -2467
rect 1094 -2542 1095 -2476
rect 1094 -2477 1095 -2467
rect 1094 -2542 1095 -2476
rect 107 -2479 108 -2467
rect 467 -2479 468 -2467
rect 492 -2479 493 -2467
rect 604 -2542 605 -2478
rect 618 -2479 619 -2467
rect 723 -2542 724 -2478
rect 758 -2542 759 -2478
rect 842 -2479 843 -2467
rect 863 -2542 864 -2478
rect 982 -2479 983 -2467
rect 124 -2481 125 -2467
rect 226 -2481 227 -2467
rect 247 -2481 248 -2467
rect 492 -2542 493 -2480
rect 499 -2481 500 -2467
rect 583 -2542 584 -2480
rect 639 -2542 640 -2480
rect 786 -2481 787 -2467
rect 800 -2481 801 -2467
rect 810 -2542 811 -2480
rect 926 -2542 927 -2480
rect 996 -2481 997 -2467
rect 173 -2483 174 -2467
rect 247 -2542 248 -2482
rect 254 -2483 255 -2467
rect 254 -2542 255 -2482
rect 254 -2483 255 -2467
rect 254 -2542 255 -2482
rect 278 -2542 279 -2482
rect 359 -2483 360 -2467
rect 373 -2483 374 -2467
rect 443 -2483 444 -2467
rect 446 -2483 447 -2467
rect 849 -2483 850 -2467
rect 201 -2485 202 -2467
rect 226 -2542 227 -2484
rect 282 -2485 283 -2467
rect 478 -2542 479 -2484
rect 499 -2542 500 -2484
rect 744 -2485 745 -2467
rect 772 -2485 773 -2467
rect 793 -2542 794 -2484
rect 800 -2542 801 -2484
rect 912 -2485 913 -2467
rect 212 -2487 213 -2467
rect 551 -2542 552 -2486
rect 565 -2487 566 -2467
rect 975 -2487 976 -2467
rect 219 -2489 220 -2467
rect 355 -2489 356 -2467
rect 359 -2542 360 -2488
rect 376 -2489 377 -2467
rect 380 -2489 381 -2467
rect 684 -2542 685 -2488
rect 730 -2489 731 -2467
rect 786 -2542 787 -2488
rect 807 -2542 808 -2488
rect 989 -2489 990 -2467
rect 205 -2491 206 -2467
rect 380 -2542 381 -2490
rect 390 -2542 391 -2490
rect 513 -2491 514 -2467
rect 520 -2491 521 -2467
rect 695 -2542 696 -2490
rect 730 -2542 731 -2490
rect 751 -2491 752 -2467
rect 772 -2542 773 -2490
rect 835 -2491 836 -2467
rect 912 -2542 913 -2490
rect 954 -2491 955 -2467
rect 975 -2542 976 -2490
rect 1003 -2491 1004 -2467
rect 93 -2493 94 -2467
rect 520 -2542 521 -2492
rect 544 -2542 545 -2492
rect 572 -2493 573 -2467
rect 597 -2493 598 -2467
rect 744 -2542 745 -2492
rect 954 -2542 955 -2492
rect 1017 -2493 1018 -2467
rect 114 -2495 115 -2467
rect 572 -2542 573 -2494
rect 597 -2542 598 -2494
rect 737 -2495 738 -2467
rect 1017 -2542 1018 -2494
rect 1031 -2495 1032 -2467
rect 282 -2542 283 -2496
rect 345 -2497 346 -2467
rect 373 -2542 374 -2496
rect 534 -2497 535 -2467
rect 548 -2497 549 -2467
rect 943 -2497 944 -2467
rect 1031 -2542 1032 -2496
rect 1066 -2497 1067 -2467
rect 289 -2499 290 -2467
rect 611 -2499 612 -2467
rect 646 -2499 647 -2467
rect 751 -2542 752 -2498
rect 1066 -2542 1067 -2498
rect 1080 -2499 1081 -2467
rect 233 -2501 234 -2467
rect 289 -2542 290 -2500
rect 296 -2501 297 -2467
rect 677 -2501 678 -2467
rect 170 -2503 171 -2467
rect 233 -2542 234 -2502
rect 296 -2542 297 -2502
rect 303 -2503 304 -2467
rect 317 -2503 318 -2467
rect 439 -2503 440 -2467
rect 443 -2542 444 -2502
rect 555 -2503 556 -2467
rect 569 -2503 570 -2467
rect 779 -2503 780 -2467
rect 100 -2505 101 -2467
rect 303 -2542 304 -2504
rect 327 -2542 328 -2504
rect 401 -2505 402 -2467
rect 415 -2505 416 -2467
rect 534 -2542 535 -2504
rect 541 -2505 542 -2467
rect 611 -2542 612 -2504
rect 646 -2542 647 -2504
rect 653 -2505 654 -2467
rect 737 -2542 738 -2504
rect 240 -2507 241 -2467
rect 415 -2542 416 -2506
rect 422 -2507 423 -2467
rect 618 -2542 619 -2506
rect 653 -2542 654 -2506
rect 702 -2507 703 -2467
rect 275 -2509 276 -2467
rect 317 -2542 318 -2508
rect 331 -2509 332 -2467
rect 464 -2542 465 -2508
rect 509 -2542 510 -2508
rect 968 -2509 969 -2467
rect 128 -2511 129 -2467
rect 331 -2542 332 -2510
rect 338 -2511 339 -2467
rect 338 -2542 339 -2510
rect 338 -2511 339 -2467
rect 338 -2542 339 -2510
rect 345 -2542 346 -2510
rect 485 -2511 486 -2467
rect 513 -2542 514 -2510
rect 709 -2511 710 -2467
rect 121 -2513 122 -2467
rect 128 -2542 129 -2512
rect 310 -2513 311 -2467
rect 401 -2542 402 -2512
rect 429 -2513 430 -2467
rect 660 -2513 661 -2467
rect 667 -2513 668 -2467
rect 674 -2542 675 -2512
rect 702 -2542 703 -2512
rect 716 -2513 717 -2467
rect 184 -2515 185 -2467
rect 310 -2542 311 -2514
rect 408 -2515 409 -2467
rect 429 -2542 430 -2514
rect 436 -2515 437 -2467
rect 905 -2515 906 -2467
rect 268 -2517 269 -2467
rect 408 -2542 409 -2516
rect 450 -2517 451 -2467
rect 474 -2542 475 -2516
rect 485 -2542 486 -2516
rect 814 -2517 815 -2467
rect 142 -2519 143 -2467
rect 268 -2542 269 -2518
rect 387 -2519 388 -2467
rect 436 -2542 437 -2518
rect 527 -2519 528 -2467
rect 709 -2542 710 -2518
rect 177 -2521 178 -2467
rect 450 -2542 451 -2520
rect 548 -2542 549 -2520
rect 919 -2521 920 -2467
rect 387 -2542 388 -2522
rect 394 -2523 395 -2467
rect 555 -2542 556 -2522
rect 688 -2523 689 -2467
rect 324 -2525 325 -2467
rect 394 -2542 395 -2524
rect 569 -2542 570 -2524
rect 681 -2525 682 -2467
rect 576 -2527 577 -2467
rect 667 -2542 668 -2526
rect 681 -2542 682 -2526
rect 933 -2527 934 -2467
rect 457 -2529 458 -2467
rect 576 -2542 577 -2528
rect 590 -2529 591 -2467
rect 779 -2542 780 -2528
rect 884 -2529 885 -2467
rect 933 -2542 934 -2528
rect 422 -2542 423 -2530
rect 457 -2542 458 -2530
rect 590 -2542 591 -2530
rect 891 -2531 892 -2467
rect 632 -2533 633 -2467
rect 716 -2542 717 -2532
rect 562 -2535 563 -2467
rect 632 -2542 633 -2534
rect 660 -2542 661 -2534
rect 765 -2535 766 -2467
rect 506 -2537 507 -2467
rect 562 -2542 563 -2536
rect 765 -2542 766 -2536
rect 898 -2537 899 -2467
rect 261 -2539 262 -2467
rect 506 -2542 507 -2538
rect 156 -2541 157 -2467
rect 261 -2542 262 -2540
rect 131 -2587 132 -2551
rect 135 -2552 136 -2550
rect 226 -2552 227 -2550
rect 257 -2587 258 -2551
rect 261 -2552 262 -2550
rect 366 -2552 367 -2550
rect 380 -2552 381 -2550
rect 527 -2552 528 -2550
rect 530 -2552 531 -2550
rect 702 -2552 703 -2550
rect 716 -2552 717 -2550
rect 807 -2552 808 -2550
rect 814 -2587 815 -2551
rect 828 -2552 829 -2550
rect 866 -2552 867 -2550
rect 926 -2552 927 -2550
rect 933 -2552 934 -2550
rect 964 -2587 965 -2551
rect 968 -2587 969 -2551
rect 975 -2552 976 -2550
rect 1013 -2587 1014 -2551
rect 1038 -2552 1039 -2550
rect 1045 -2587 1046 -2551
rect 1052 -2552 1053 -2550
rect 1059 -2587 1060 -2551
rect 1066 -2552 1067 -2550
rect 1143 -2552 1144 -2550
rect 1178 -2552 1179 -2550
rect 1181 -2552 1182 -2550
rect 1185 -2552 1186 -2550
rect 128 -2554 129 -2550
rect 135 -2587 136 -2553
rect 233 -2554 234 -2550
rect 275 -2554 276 -2550
rect 282 -2554 283 -2550
rect 387 -2554 388 -2550
rect 394 -2554 395 -2550
rect 471 -2587 472 -2553
rect 478 -2554 479 -2550
rect 677 -2587 678 -2553
rect 681 -2554 682 -2550
rect 772 -2554 773 -2550
rect 870 -2554 871 -2550
rect 887 -2587 888 -2553
rect 898 -2587 899 -2553
rect 912 -2554 913 -2550
rect 1017 -2554 1018 -2550
rect 1017 -2587 1018 -2553
rect 1017 -2554 1018 -2550
rect 1017 -2587 1018 -2553
rect 1024 -2587 1025 -2553
rect 1031 -2554 1032 -2550
rect 247 -2556 248 -2550
rect 324 -2556 325 -2550
rect 331 -2556 332 -2550
rect 485 -2556 486 -2550
rect 492 -2556 493 -2550
rect 684 -2556 685 -2550
rect 688 -2556 689 -2550
rect 730 -2556 731 -2550
rect 744 -2556 745 -2550
rect 793 -2556 794 -2550
rect 884 -2587 885 -2555
rect 954 -2556 955 -2550
rect 254 -2558 255 -2550
rect 254 -2587 255 -2557
rect 254 -2558 255 -2550
rect 254 -2587 255 -2557
rect 268 -2558 269 -2550
rect 324 -2587 325 -2557
rect 345 -2558 346 -2550
rect 366 -2587 367 -2557
rect 401 -2558 402 -2550
rect 548 -2558 549 -2550
rect 551 -2587 552 -2557
rect 653 -2558 654 -2550
rect 663 -2587 664 -2557
rect 667 -2558 668 -2550
rect 681 -2587 682 -2557
rect 779 -2558 780 -2550
rect 947 -2558 948 -2550
rect 954 -2587 955 -2557
rect 289 -2560 290 -2550
rect 383 -2587 384 -2559
rect 415 -2560 416 -2550
rect 492 -2587 493 -2559
rect 499 -2560 500 -2550
rect 499 -2587 500 -2559
rect 499 -2560 500 -2550
rect 499 -2587 500 -2559
rect 506 -2560 507 -2550
rect 611 -2560 612 -2550
rect 621 -2560 622 -2550
rect 800 -2560 801 -2550
rect 303 -2562 304 -2550
rect 593 -2562 594 -2550
rect 600 -2587 601 -2561
rect 646 -2562 647 -2550
rect 660 -2562 661 -2550
rect 667 -2587 668 -2561
rect 691 -2562 692 -2550
rect 691 -2587 692 -2561
rect 691 -2562 692 -2550
rect 691 -2587 692 -2561
rect 716 -2587 717 -2561
rect 758 -2562 759 -2550
rect 310 -2564 311 -2550
rect 649 -2587 650 -2563
rect 723 -2564 724 -2550
rect 810 -2587 811 -2563
rect 317 -2566 318 -2550
rect 331 -2587 332 -2565
rect 359 -2566 360 -2550
rect 506 -2587 507 -2565
rect 523 -2566 524 -2550
rect 541 -2566 542 -2550
rect 565 -2587 566 -2565
rect 639 -2566 640 -2550
rect 723 -2587 724 -2565
rect 765 -2566 766 -2550
rect 429 -2568 430 -2550
rect 488 -2568 489 -2550
rect 527 -2587 528 -2567
rect 555 -2568 556 -2550
rect 569 -2568 570 -2550
rect 674 -2568 675 -2550
rect 730 -2587 731 -2567
rect 751 -2568 752 -2550
rect 436 -2570 437 -2550
rect 544 -2587 545 -2569
rect 576 -2570 577 -2550
rect 590 -2570 591 -2550
rect 632 -2570 633 -2550
rect 712 -2587 713 -2569
rect 747 -2570 748 -2550
rect 786 -2570 787 -2550
rect 443 -2572 444 -2550
rect 460 -2572 461 -2550
rect 513 -2572 514 -2550
rect 555 -2587 556 -2571
rect 576 -2587 577 -2571
rect 597 -2572 598 -2550
rect 695 -2572 696 -2550
rect 751 -2587 752 -2571
rect 338 -2574 339 -2550
rect 513 -2587 514 -2573
rect 530 -2587 531 -2573
rect 562 -2574 563 -2550
rect 296 -2576 297 -2550
rect 338 -2587 339 -2575
rect 373 -2576 374 -2550
rect 443 -2587 444 -2575
rect 450 -2576 451 -2550
rect 569 -2587 570 -2575
rect 352 -2578 353 -2550
rect 450 -2587 451 -2577
rect 464 -2578 465 -2550
rect 597 -2587 598 -2577
rect 373 -2587 374 -2579
rect 422 -2580 423 -2550
rect 534 -2580 535 -2550
rect 646 -2587 647 -2579
rect 408 -2582 409 -2550
rect 534 -2587 535 -2581
rect 541 -2587 542 -2581
rect 709 -2582 710 -2550
rect 562 -2587 563 -2583
rect 625 -2584 626 -2550
rect 604 -2586 605 -2550
rect 709 -2587 710 -2585
rect 131 -2597 132 -2595
rect 135 -2597 136 -2595
rect 324 -2597 325 -2595
rect 383 -2597 384 -2595
rect 443 -2597 444 -2595
rect 516 -2597 517 -2595
rect 534 -2597 535 -2595
rect 663 -2597 664 -2595
rect 674 -2597 675 -2595
rect 723 -2597 724 -2595
rect 751 -2597 752 -2595
rect 807 -2597 808 -2595
rect 810 -2597 811 -2595
rect 814 -2597 815 -2595
rect 884 -2597 885 -2595
rect 898 -2597 899 -2595
rect 954 -2597 955 -2595
rect 964 -2597 965 -2595
rect 1010 -2597 1011 -2595
rect 1017 -2597 1018 -2595
rect 1045 -2597 1046 -2595
rect 1052 -2597 1053 -2595
rect 1055 -2597 1056 -2595
rect 1059 -2597 1060 -2595
rect 331 -2599 332 -2595
rect 348 -2599 349 -2595
rect 366 -2599 367 -2595
rect 380 -2599 381 -2595
rect 450 -2599 451 -2595
rect 544 -2599 545 -2595
rect 548 -2599 549 -2595
rect 576 -2599 577 -2595
rect 660 -2599 661 -2595
rect 667 -2599 668 -2595
rect 684 -2599 685 -2595
rect 716 -2599 717 -2595
rect 961 -2599 962 -2595
rect 968 -2599 969 -2595
rect 1013 -2599 1014 -2595
rect 1024 -2599 1025 -2595
rect 338 -2601 339 -2595
rect 373 -2601 374 -2595
rect 471 -2601 472 -2595
rect 551 -2601 552 -2595
rect 555 -2601 556 -2595
rect 600 -2601 601 -2595
rect 709 -2601 710 -2595
rect 730 -2601 731 -2595
rect 492 -2603 493 -2595
rect 565 -2603 566 -2595
rect 569 -2603 570 -2595
rect 681 -2603 682 -2595
rect 499 -2605 500 -2595
rect 513 -2605 514 -2595
rect 506 -2607 507 -2595
rect 649 -2607 650 -2595
<< labels >>
rlabel pdiffusion 157 -20 157 -20 0 cellNo=95
rlabel pdiffusion 213 -20 213 -20 0 cellNo=341
rlabel pdiffusion 241 -20 241 -20 0 feedthrough
rlabel pdiffusion 248 -20 248 -20 0 feedthrough
rlabel pdiffusion 262 -20 262 -20 0 feedthrough
rlabel pdiffusion 269 -20 269 -20 0 cellNo=486
rlabel pdiffusion 276 -20 276 -20 0 feedthrough
rlabel pdiffusion 283 -20 283 -20 0 cellNo=262
rlabel pdiffusion 339 -20 339 -20 0 feedthrough
rlabel pdiffusion 374 -20 374 -20 0 feedthrough
rlabel pdiffusion 381 -20 381 -20 0 cellNo=510
rlabel pdiffusion 388 -20 388 -20 0 feedthrough
rlabel pdiffusion 395 -20 395 -20 0 cellNo=19
rlabel pdiffusion 402 -20 402 -20 0 cellNo=449
rlabel pdiffusion 409 -20 409 -20 0 cellNo=394
rlabel pdiffusion 416 -20 416 -20 0 feedthrough
rlabel pdiffusion 423 -20 423 -20 0 cellNo=465
rlabel pdiffusion 430 -20 430 -20 0 feedthrough
rlabel pdiffusion 458 -20 458 -20 0 cellNo=565
rlabel pdiffusion 465 -20 465 -20 0 cellNo=508
rlabel pdiffusion 479 -20 479 -20 0 cellNo=566
rlabel pdiffusion 486 -20 486 -20 0 feedthrough
rlabel pdiffusion 500 -20 500 -20 0 feedthrough
rlabel pdiffusion 507 -20 507 -20 0 feedthrough
rlabel pdiffusion 514 -20 514 -20 0 cellNo=451
rlabel pdiffusion 528 -20 528 -20 0 feedthrough
rlabel pdiffusion 549 -20 549 -20 0 cellNo=201
rlabel pdiffusion 563 -20 563 -20 0 cellNo=109
rlabel pdiffusion 570 -20 570 -20 0 feedthrough
rlabel pdiffusion 577 -20 577 -20 0 feedthrough
rlabel pdiffusion 584 -20 584 -20 0 cellNo=214
rlabel pdiffusion 605 -20 605 -20 0 cellNo=110
rlabel pdiffusion 640 -20 640 -20 0 feedthrough
rlabel pdiffusion 668 -20 668 -20 0 feedthrough
rlabel pdiffusion 682 -20 682 -20 0 feedthrough
rlabel pdiffusion 703 -20 703 -20 0 cellNo=49
rlabel pdiffusion 710 -20 710 -20 0 feedthrough
rlabel pdiffusion 766 -20 766 -20 0 feedthrough
rlabel pdiffusion 801 -20 801 -20 0 cellNo=230
rlabel pdiffusion 829 -20 829 -20 0 feedthrough
rlabel pdiffusion 150 -63 150 -63 0 cellNo=363
rlabel pdiffusion 157 -63 157 -63 0 cellNo=435
rlabel pdiffusion 164 -63 164 -63 0 feedthrough
rlabel pdiffusion 192 -63 192 -63 0 feedthrough
rlabel pdiffusion 220 -63 220 -63 0 feedthrough
rlabel pdiffusion 227 -63 227 -63 0 feedthrough
rlabel pdiffusion 234 -63 234 -63 0 feedthrough
rlabel pdiffusion 248 -63 248 -63 0 feedthrough
rlabel pdiffusion 255 -63 255 -63 0 feedthrough
rlabel pdiffusion 262 -63 262 -63 0 feedthrough
rlabel pdiffusion 269 -63 269 -63 0 feedthrough
rlabel pdiffusion 276 -63 276 -63 0 feedthrough
rlabel pdiffusion 283 -63 283 -63 0 feedthrough
rlabel pdiffusion 290 -63 290 -63 0 cellNo=468
rlabel pdiffusion 297 -63 297 -63 0 feedthrough
rlabel pdiffusion 304 -63 304 -63 0 feedthrough
rlabel pdiffusion 311 -63 311 -63 0 cellNo=175
rlabel pdiffusion 318 -63 318 -63 0 feedthrough
rlabel pdiffusion 325 -63 325 -63 0 feedthrough
rlabel pdiffusion 332 -63 332 -63 0 feedthrough
rlabel pdiffusion 339 -63 339 -63 0 cellNo=82
rlabel pdiffusion 346 -63 346 -63 0 cellNo=483
rlabel pdiffusion 353 -63 353 -63 0 cellNo=477
rlabel pdiffusion 360 -63 360 -63 0 feedthrough
rlabel pdiffusion 367 -63 367 -63 0 feedthrough
rlabel pdiffusion 374 -63 374 -63 0 feedthrough
rlabel pdiffusion 381 -63 381 -63 0 cellNo=282
rlabel pdiffusion 388 -63 388 -63 0 feedthrough
rlabel pdiffusion 395 -63 395 -63 0 feedthrough
rlabel pdiffusion 402 -63 402 -63 0 feedthrough
rlabel pdiffusion 409 -63 409 -63 0 cellNo=165
rlabel pdiffusion 416 -63 416 -63 0 cellNo=234
rlabel pdiffusion 423 -63 423 -63 0 feedthrough
rlabel pdiffusion 430 -63 430 -63 0 feedthrough
rlabel pdiffusion 437 -63 437 -63 0 feedthrough
rlabel pdiffusion 444 -63 444 -63 0 feedthrough
rlabel pdiffusion 451 -63 451 -63 0 cellNo=103
rlabel pdiffusion 458 -63 458 -63 0 feedthrough
rlabel pdiffusion 465 -63 465 -63 0 feedthrough
rlabel pdiffusion 472 -63 472 -63 0 feedthrough
rlabel pdiffusion 479 -63 479 -63 0 cellNo=357
rlabel pdiffusion 486 -63 486 -63 0 feedthrough
rlabel pdiffusion 493 -63 493 -63 0 feedthrough
rlabel pdiffusion 500 -63 500 -63 0 cellNo=554
rlabel pdiffusion 507 -63 507 -63 0 feedthrough
rlabel pdiffusion 514 -63 514 -63 0 feedthrough
rlabel pdiffusion 521 -63 521 -63 0 feedthrough
rlabel pdiffusion 528 -63 528 -63 0 feedthrough
rlabel pdiffusion 535 -63 535 -63 0 cellNo=511
rlabel pdiffusion 542 -63 542 -63 0 feedthrough
rlabel pdiffusion 549 -63 549 -63 0 feedthrough
rlabel pdiffusion 556 -63 556 -63 0 cellNo=548
rlabel pdiffusion 563 -63 563 -63 0 feedthrough
rlabel pdiffusion 570 -63 570 -63 0 feedthrough
rlabel pdiffusion 577 -63 577 -63 0 cellNo=399
rlabel pdiffusion 584 -63 584 -63 0 feedthrough
rlabel pdiffusion 591 -63 591 -63 0 cellNo=176
rlabel pdiffusion 598 -63 598 -63 0 feedthrough
rlabel pdiffusion 605 -63 605 -63 0 feedthrough
rlabel pdiffusion 612 -63 612 -63 0 feedthrough
rlabel pdiffusion 619 -63 619 -63 0 cellNo=164
rlabel pdiffusion 626 -63 626 -63 0 feedthrough
rlabel pdiffusion 633 -63 633 -63 0 feedthrough
rlabel pdiffusion 640 -63 640 -63 0 feedthrough
rlabel pdiffusion 647 -63 647 -63 0 feedthrough
rlabel pdiffusion 654 -63 654 -63 0 feedthrough
rlabel pdiffusion 661 -63 661 -63 0 feedthrough
rlabel pdiffusion 668 -63 668 -63 0 cellNo=326
rlabel pdiffusion 675 -63 675 -63 0 feedthrough
rlabel pdiffusion 682 -63 682 -63 0 feedthrough
rlabel pdiffusion 689 -63 689 -63 0 feedthrough
rlabel pdiffusion 703 -63 703 -63 0 feedthrough
rlabel pdiffusion 717 -63 717 -63 0 cellNo=11
rlabel pdiffusion 724 -63 724 -63 0 feedthrough
rlabel pdiffusion 752 -63 752 -63 0 feedthrough
rlabel pdiffusion 759 -63 759 -63 0 feedthrough
rlabel pdiffusion 773 -63 773 -63 0 feedthrough
rlabel pdiffusion 829 -63 829 -63 0 feedthrough
rlabel pdiffusion 850 -63 850 -63 0 feedthrough
rlabel pdiffusion 878 -63 878 -63 0 feedthrough
rlabel pdiffusion 906 -63 906 -63 0 feedthrough
rlabel pdiffusion 24 -124 24 -124 0 feedthrough
rlabel pdiffusion 31 -124 31 -124 0 feedthrough
rlabel pdiffusion 38 -124 38 -124 0 feedthrough
rlabel pdiffusion 45 -124 45 -124 0 feedthrough
rlabel pdiffusion 52 -124 52 -124 0 feedthrough
rlabel pdiffusion 59 -124 59 -124 0 cellNo=302
rlabel pdiffusion 66 -124 66 -124 0 cellNo=144
rlabel pdiffusion 73 -124 73 -124 0 cellNo=338
rlabel pdiffusion 80 -124 80 -124 0 feedthrough
rlabel pdiffusion 87 -124 87 -124 0 cellNo=182
rlabel pdiffusion 94 -124 94 -124 0 feedthrough
rlabel pdiffusion 101 -124 101 -124 0 feedthrough
rlabel pdiffusion 108 -124 108 -124 0 feedthrough
rlabel pdiffusion 115 -124 115 -124 0 cellNo=140
rlabel pdiffusion 122 -124 122 -124 0 feedthrough
rlabel pdiffusion 129 -124 129 -124 0 cellNo=52
rlabel pdiffusion 136 -124 136 -124 0 feedthrough
rlabel pdiffusion 143 -124 143 -124 0 feedthrough
rlabel pdiffusion 150 -124 150 -124 0 feedthrough
rlabel pdiffusion 157 -124 157 -124 0 feedthrough
rlabel pdiffusion 164 -124 164 -124 0 feedthrough
rlabel pdiffusion 171 -124 171 -124 0 feedthrough
rlabel pdiffusion 178 -124 178 -124 0 feedthrough
rlabel pdiffusion 185 -124 185 -124 0 cellNo=192
rlabel pdiffusion 192 -124 192 -124 0 cellNo=87
rlabel pdiffusion 199 -124 199 -124 0 feedthrough
rlabel pdiffusion 206 -124 206 -124 0 feedthrough
rlabel pdiffusion 213 -124 213 -124 0 feedthrough
rlabel pdiffusion 220 -124 220 -124 0 feedthrough
rlabel pdiffusion 227 -124 227 -124 0 feedthrough
rlabel pdiffusion 234 -124 234 -124 0 feedthrough
rlabel pdiffusion 241 -124 241 -124 0 feedthrough
rlabel pdiffusion 248 -124 248 -124 0 feedthrough
rlabel pdiffusion 255 -124 255 -124 0 feedthrough
rlabel pdiffusion 262 -124 262 -124 0 feedthrough
rlabel pdiffusion 269 -124 269 -124 0 cellNo=429
rlabel pdiffusion 276 -124 276 -124 0 feedthrough
rlabel pdiffusion 283 -124 283 -124 0 feedthrough
rlabel pdiffusion 290 -124 290 -124 0 feedthrough
rlabel pdiffusion 297 -124 297 -124 0 cellNo=276
rlabel pdiffusion 304 -124 304 -124 0 feedthrough
rlabel pdiffusion 311 -124 311 -124 0 cellNo=450
rlabel pdiffusion 318 -124 318 -124 0 feedthrough
rlabel pdiffusion 325 -124 325 -124 0 cellNo=312
rlabel pdiffusion 332 -124 332 -124 0 feedthrough
rlabel pdiffusion 339 -124 339 -124 0 feedthrough
rlabel pdiffusion 346 -124 346 -124 0 feedthrough
rlabel pdiffusion 353 -124 353 -124 0 feedthrough
rlabel pdiffusion 360 -124 360 -124 0 cellNo=151
rlabel pdiffusion 367 -124 367 -124 0 feedthrough
rlabel pdiffusion 374 -124 374 -124 0 feedthrough
rlabel pdiffusion 381 -124 381 -124 0 feedthrough
rlabel pdiffusion 388 -124 388 -124 0 feedthrough
rlabel pdiffusion 395 -124 395 -124 0 cellNo=298
rlabel pdiffusion 402 -124 402 -124 0 cellNo=63
rlabel pdiffusion 409 -124 409 -124 0 feedthrough
rlabel pdiffusion 416 -124 416 -124 0 feedthrough
rlabel pdiffusion 423 -124 423 -124 0 feedthrough
rlabel pdiffusion 430 -124 430 -124 0 feedthrough
rlabel pdiffusion 437 -124 437 -124 0 cellNo=393
rlabel pdiffusion 444 -124 444 -124 0 feedthrough
rlabel pdiffusion 451 -124 451 -124 0 feedthrough
rlabel pdiffusion 458 -124 458 -124 0 feedthrough
rlabel pdiffusion 465 -124 465 -124 0 feedthrough
rlabel pdiffusion 472 -124 472 -124 0 feedthrough
rlabel pdiffusion 479 -124 479 -124 0 feedthrough
rlabel pdiffusion 486 -124 486 -124 0 feedthrough
rlabel pdiffusion 493 -124 493 -124 0 feedthrough
rlabel pdiffusion 500 -124 500 -124 0 feedthrough
rlabel pdiffusion 507 -124 507 -124 0 feedthrough
rlabel pdiffusion 514 -124 514 -124 0 feedthrough
rlabel pdiffusion 521 -124 521 -124 0 feedthrough
rlabel pdiffusion 528 -124 528 -124 0 cellNo=166
rlabel pdiffusion 535 -124 535 -124 0 feedthrough
rlabel pdiffusion 542 -124 542 -124 0 feedthrough
rlabel pdiffusion 549 -124 549 -124 0 feedthrough
rlabel pdiffusion 556 -124 556 -124 0 feedthrough
rlabel pdiffusion 563 -124 563 -124 0 feedthrough
rlabel pdiffusion 570 -124 570 -124 0 feedthrough
rlabel pdiffusion 577 -124 577 -124 0 feedthrough
rlabel pdiffusion 584 -124 584 -124 0 feedthrough
rlabel pdiffusion 591 -124 591 -124 0 feedthrough
rlabel pdiffusion 598 -124 598 -124 0 feedthrough
rlabel pdiffusion 605 -124 605 -124 0 cellNo=497
rlabel pdiffusion 612 -124 612 -124 0 feedthrough
rlabel pdiffusion 619 -124 619 -124 0 feedthrough
rlabel pdiffusion 626 -124 626 -124 0 feedthrough
rlabel pdiffusion 633 -124 633 -124 0 feedthrough
rlabel pdiffusion 640 -124 640 -124 0 feedthrough
rlabel pdiffusion 647 -124 647 -124 0 feedthrough
rlabel pdiffusion 654 -124 654 -124 0 feedthrough
rlabel pdiffusion 661 -124 661 -124 0 cellNo=377
rlabel pdiffusion 668 -124 668 -124 0 feedthrough
rlabel pdiffusion 675 -124 675 -124 0 feedthrough
rlabel pdiffusion 682 -124 682 -124 0 feedthrough
rlabel pdiffusion 689 -124 689 -124 0 feedthrough
rlabel pdiffusion 696 -124 696 -124 0 feedthrough
rlabel pdiffusion 703 -124 703 -124 0 feedthrough
rlabel pdiffusion 710 -124 710 -124 0 feedthrough
rlabel pdiffusion 717 -124 717 -124 0 feedthrough
rlabel pdiffusion 724 -124 724 -124 0 feedthrough
rlabel pdiffusion 731 -124 731 -124 0 feedthrough
rlabel pdiffusion 738 -124 738 -124 0 feedthrough
rlabel pdiffusion 745 -124 745 -124 0 feedthrough
rlabel pdiffusion 752 -124 752 -124 0 feedthrough
rlabel pdiffusion 759 -124 759 -124 0 cellNo=25
rlabel pdiffusion 766 -124 766 -124 0 feedthrough
rlabel pdiffusion 773 -124 773 -124 0 feedthrough
rlabel pdiffusion 780 -124 780 -124 0 feedthrough
rlabel pdiffusion 787 -124 787 -124 0 feedthrough
rlabel pdiffusion 794 -124 794 -124 0 feedthrough
rlabel pdiffusion 801 -124 801 -124 0 feedthrough
rlabel pdiffusion 808 -124 808 -124 0 feedthrough
rlabel pdiffusion 815 -124 815 -124 0 feedthrough
rlabel pdiffusion 822 -124 822 -124 0 feedthrough
rlabel pdiffusion 850 -124 850 -124 0 feedthrough
rlabel pdiffusion 857 -124 857 -124 0 feedthrough
rlabel pdiffusion 871 -124 871 -124 0 feedthrough
rlabel pdiffusion 878 -124 878 -124 0 feedthrough
rlabel pdiffusion 941 -124 941 -124 0 feedthrough
rlabel pdiffusion 948 -124 948 -124 0 feedthrough
rlabel pdiffusion 1501 -124 1501 -124 0 feedthrough
rlabel pdiffusion 1508 -124 1508 -124 0 cellNo=174
rlabel pdiffusion 10 -203 10 -203 0 feedthrough
rlabel pdiffusion 17 -203 17 -203 0 feedthrough
rlabel pdiffusion 24 -203 24 -203 0 feedthrough
rlabel pdiffusion 31 -203 31 -203 0 feedthrough
rlabel pdiffusion 38 -203 38 -203 0 feedthrough
rlabel pdiffusion 45 -203 45 -203 0 feedthrough
rlabel pdiffusion 52 -203 52 -203 0 cellNo=415
rlabel pdiffusion 59 -203 59 -203 0 feedthrough
rlabel pdiffusion 66 -203 66 -203 0 feedthrough
rlabel pdiffusion 73 -203 73 -203 0 feedthrough
rlabel pdiffusion 80 -203 80 -203 0 feedthrough
rlabel pdiffusion 87 -203 87 -203 0 feedthrough
rlabel pdiffusion 94 -203 94 -203 0 feedthrough
rlabel pdiffusion 101 -203 101 -203 0 cellNo=421
rlabel pdiffusion 108 -203 108 -203 0 feedthrough
rlabel pdiffusion 115 -203 115 -203 0 feedthrough
rlabel pdiffusion 122 -203 122 -203 0 feedthrough
rlabel pdiffusion 129 -203 129 -203 0 feedthrough
rlabel pdiffusion 136 -203 136 -203 0 feedthrough
rlabel pdiffusion 143 -203 143 -203 0 cellNo=241
rlabel pdiffusion 150 -203 150 -203 0 cellNo=271
rlabel pdiffusion 157 -203 157 -203 0 cellNo=539
rlabel pdiffusion 164 -203 164 -203 0 feedthrough
rlabel pdiffusion 171 -203 171 -203 0 feedthrough
rlabel pdiffusion 178 -203 178 -203 0 feedthrough
rlabel pdiffusion 185 -203 185 -203 0 feedthrough
rlabel pdiffusion 192 -203 192 -203 0 feedthrough
rlabel pdiffusion 199 -203 199 -203 0 feedthrough
rlabel pdiffusion 206 -203 206 -203 0 feedthrough
rlabel pdiffusion 213 -203 213 -203 0 feedthrough
rlabel pdiffusion 220 -203 220 -203 0 feedthrough
rlabel pdiffusion 227 -203 227 -203 0 feedthrough
rlabel pdiffusion 234 -203 234 -203 0 feedthrough
rlabel pdiffusion 241 -203 241 -203 0 cellNo=78
rlabel pdiffusion 248 -203 248 -203 0 feedthrough
rlabel pdiffusion 255 -203 255 -203 0 feedthrough
rlabel pdiffusion 262 -203 262 -203 0 feedthrough
rlabel pdiffusion 269 -203 269 -203 0 cellNo=401
rlabel pdiffusion 276 -203 276 -203 0 feedthrough
rlabel pdiffusion 283 -203 283 -203 0 feedthrough
rlabel pdiffusion 290 -203 290 -203 0 feedthrough
rlabel pdiffusion 297 -203 297 -203 0 feedthrough
rlabel pdiffusion 304 -203 304 -203 0 cellNo=122
rlabel pdiffusion 311 -203 311 -203 0 feedthrough
rlabel pdiffusion 318 -203 318 -203 0 cellNo=414
rlabel pdiffusion 325 -203 325 -203 0 feedthrough
rlabel pdiffusion 332 -203 332 -203 0 cellNo=319
rlabel pdiffusion 339 -203 339 -203 0 feedthrough
rlabel pdiffusion 346 -203 346 -203 0 feedthrough
rlabel pdiffusion 353 -203 353 -203 0 feedthrough
rlabel pdiffusion 360 -203 360 -203 0 feedthrough
rlabel pdiffusion 367 -203 367 -203 0 feedthrough
rlabel pdiffusion 374 -203 374 -203 0 feedthrough
rlabel pdiffusion 381 -203 381 -203 0 feedthrough
rlabel pdiffusion 388 -203 388 -203 0 cellNo=40
rlabel pdiffusion 395 -203 395 -203 0 feedthrough
rlabel pdiffusion 402 -203 402 -203 0 feedthrough
rlabel pdiffusion 409 -203 409 -203 0 feedthrough
rlabel pdiffusion 416 -203 416 -203 0 feedthrough
rlabel pdiffusion 423 -203 423 -203 0 feedthrough
rlabel pdiffusion 430 -203 430 -203 0 feedthrough
rlabel pdiffusion 437 -203 437 -203 0 cellNo=184
rlabel pdiffusion 444 -203 444 -203 0 cellNo=286
rlabel pdiffusion 451 -203 451 -203 0 feedthrough
rlabel pdiffusion 458 -203 458 -203 0 cellNo=461
rlabel pdiffusion 465 -203 465 -203 0 feedthrough
rlabel pdiffusion 472 -203 472 -203 0 feedthrough
rlabel pdiffusion 479 -203 479 -203 0 feedthrough
rlabel pdiffusion 486 -203 486 -203 0 cellNo=124
rlabel pdiffusion 493 -203 493 -203 0 feedthrough
rlabel pdiffusion 500 -203 500 -203 0 feedthrough
rlabel pdiffusion 507 -203 507 -203 0 feedthrough
rlabel pdiffusion 514 -203 514 -203 0 cellNo=368
rlabel pdiffusion 521 -203 521 -203 0 feedthrough
rlabel pdiffusion 528 -203 528 -203 0 feedthrough
rlabel pdiffusion 535 -203 535 -203 0 cellNo=154
rlabel pdiffusion 542 -203 542 -203 0 feedthrough
rlabel pdiffusion 549 -203 549 -203 0 feedthrough
rlabel pdiffusion 556 -203 556 -203 0 feedthrough
rlabel pdiffusion 563 -203 563 -203 0 feedthrough
rlabel pdiffusion 570 -203 570 -203 0 feedthrough
rlabel pdiffusion 577 -203 577 -203 0 feedthrough
rlabel pdiffusion 584 -203 584 -203 0 feedthrough
rlabel pdiffusion 591 -203 591 -203 0 feedthrough
rlabel pdiffusion 598 -203 598 -203 0 feedthrough
rlabel pdiffusion 605 -203 605 -203 0 cellNo=595
rlabel pdiffusion 612 -203 612 -203 0 feedthrough
rlabel pdiffusion 619 -203 619 -203 0 feedthrough
rlabel pdiffusion 626 -203 626 -203 0 feedthrough
rlabel pdiffusion 633 -203 633 -203 0 feedthrough
rlabel pdiffusion 640 -203 640 -203 0 feedthrough
rlabel pdiffusion 647 -203 647 -203 0 feedthrough
rlabel pdiffusion 654 -203 654 -203 0 feedthrough
rlabel pdiffusion 661 -203 661 -203 0 feedthrough
rlabel pdiffusion 668 -203 668 -203 0 feedthrough
rlabel pdiffusion 675 -203 675 -203 0 feedthrough
rlabel pdiffusion 682 -203 682 -203 0 feedthrough
rlabel pdiffusion 689 -203 689 -203 0 feedthrough
rlabel pdiffusion 696 -203 696 -203 0 feedthrough
rlabel pdiffusion 703 -203 703 -203 0 feedthrough
rlabel pdiffusion 710 -203 710 -203 0 feedthrough
rlabel pdiffusion 717 -203 717 -203 0 cellNo=141
rlabel pdiffusion 724 -203 724 -203 0 feedthrough
rlabel pdiffusion 731 -203 731 -203 0 feedthrough
rlabel pdiffusion 738 -203 738 -203 0 feedthrough
rlabel pdiffusion 745 -203 745 -203 0 feedthrough
rlabel pdiffusion 752 -203 752 -203 0 feedthrough
rlabel pdiffusion 759 -203 759 -203 0 feedthrough
rlabel pdiffusion 766 -203 766 -203 0 feedthrough
rlabel pdiffusion 773 -203 773 -203 0 feedthrough
rlabel pdiffusion 780 -203 780 -203 0 feedthrough
rlabel pdiffusion 787 -203 787 -203 0 feedthrough
rlabel pdiffusion 794 -203 794 -203 0 feedthrough
rlabel pdiffusion 801 -203 801 -203 0 feedthrough
rlabel pdiffusion 808 -203 808 -203 0 feedthrough
rlabel pdiffusion 815 -203 815 -203 0 feedthrough
rlabel pdiffusion 822 -203 822 -203 0 feedthrough
rlabel pdiffusion 829 -203 829 -203 0 feedthrough
rlabel pdiffusion 836 -203 836 -203 0 feedthrough
rlabel pdiffusion 843 -203 843 -203 0 feedthrough
rlabel pdiffusion 850 -203 850 -203 0 feedthrough
rlabel pdiffusion 857 -203 857 -203 0 feedthrough
rlabel pdiffusion 864 -203 864 -203 0 feedthrough
rlabel pdiffusion 871 -203 871 -203 0 feedthrough
rlabel pdiffusion 878 -203 878 -203 0 feedthrough
rlabel pdiffusion 885 -203 885 -203 0 feedthrough
rlabel pdiffusion 892 -203 892 -203 0 feedthrough
rlabel pdiffusion 899 -203 899 -203 0 feedthrough
rlabel pdiffusion 906 -203 906 -203 0 feedthrough
rlabel pdiffusion 913 -203 913 -203 0 feedthrough
rlabel pdiffusion 920 -203 920 -203 0 feedthrough
rlabel pdiffusion 927 -203 927 -203 0 feedthrough
rlabel pdiffusion 934 -203 934 -203 0 feedthrough
rlabel pdiffusion 941 -203 941 -203 0 feedthrough
rlabel pdiffusion 948 -203 948 -203 0 feedthrough
rlabel pdiffusion 955 -203 955 -203 0 feedthrough
rlabel pdiffusion 962 -203 962 -203 0 feedthrough
rlabel pdiffusion 969 -203 969 -203 0 feedthrough
rlabel pdiffusion 976 -203 976 -203 0 cellNo=405
rlabel pdiffusion 983 -203 983 -203 0 cellNo=503
rlabel pdiffusion 990 -203 990 -203 0 cellNo=599
rlabel pdiffusion 997 -203 997 -203 0 feedthrough
rlabel pdiffusion 1025 -203 1025 -203 0 feedthrough
rlabel pdiffusion 1501 -203 1501 -203 0 feedthrough
rlabel pdiffusion 3 -314 3 -314 0 feedthrough
rlabel pdiffusion 10 -314 10 -314 0 feedthrough
rlabel pdiffusion 17 -314 17 -314 0 feedthrough
rlabel pdiffusion 24 -314 24 -314 0 cellNo=222
rlabel pdiffusion 31 -314 31 -314 0 cellNo=28
rlabel pdiffusion 38 -314 38 -314 0 cellNo=310
rlabel pdiffusion 45 -314 45 -314 0 feedthrough
rlabel pdiffusion 52 -314 52 -314 0 cellNo=137
rlabel pdiffusion 59 -314 59 -314 0 feedthrough
rlabel pdiffusion 66 -314 66 -314 0 cellNo=29
rlabel pdiffusion 73 -314 73 -314 0 feedthrough
rlabel pdiffusion 80 -314 80 -314 0 cellNo=170
rlabel pdiffusion 87 -314 87 -314 0 feedthrough
rlabel pdiffusion 94 -314 94 -314 0 cellNo=518
rlabel pdiffusion 101 -314 101 -314 0 feedthrough
rlabel pdiffusion 108 -314 108 -314 0 feedthrough
rlabel pdiffusion 115 -314 115 -314 0 feedthrough
rlabel pdiffusion 122 -314 122 -314 0 cellNo=515
rlabel pdiffusion 129 -314 129 -314 0 feedthrough
rlabel pdiffusion 136 -314 136 -314 0 feedthrough
rlabel pdiffusion 143 -314 143 -314 0 feedthrough
rlabel pdiffusion 150 -314 150 -314 0 feedthrough
rlabel pdiffusion 157 -314 157 -314 0 feedthrough
rlabel pdiffusion 164 -314 164 -314 0 feedthrough
rlabel pdiffusion 171 -314 171 -314 0 feedthrough
rlabel pdiffusion 178 -314 178 -314 0 feedthrough
rlabel pdiffusion 185 -314 185 -314 0 feedthrough
rlabel pdiffusion 192 -314 192 -314 0 feedthrough
rlabel pdiffusion 199 -314 199 -314 0 feedthrough
rlabel pdiffusion 206 -314 206 -314 0 feedthrough
rlabel pdiffusion 213 -314 213 -314 0 feedthrough
rlabel pdiffusion 220 -314 220 -314 0 feedthrough
rlabel pdiffusion 227 -314 227 -314 0 feedthrough
rlabel pdiffusion 234 -314 234 -314 0 feedthrough
rlabel pdiffusion 241 -314 241 -314 0 feedthrough
rlabel pdiffusion 248 -314 248 -314 0 feedthrough
rlabel pdiffusion 255 -314 255 -314 0 feedthrough
rlabel pdiffusion 262 -314 262 -314 0 feedthrough
rlabel pdiffusion 269 -314 269 -314 0 feedthrough
rlabel pdiffusion 276 -314 276 -314 0 feedthrough
rlabel pdiffusion 283 -314 283 -314 0 cellNo=179
rlabel pdiffusion 290 -314 290 -314 0 feedthrough
rlabel pdiffusion 297 -314 297 -314 0 feedthrough
rlabel pdiffusion 304 -314 304 -314 0 feedthrough
rlabel pdiffusion 311 -314 311 -314 0 cellNo=309
rlabel pdiffusion 318 -314 318 -314 0 cellNo=1
rlabel pdiffusion 325 -314 325 -314 0 cellNo=383
rlabel pdiffusion 332 -314 332 -314 0 feedthrough
rlabel pdiffusion 339 -314 339 -314 0 feedthrough
rlabel pdiffusion 346 -314 346 -314 0 feedthrough
rlabel pdiffusion 353 -314 353 -314 0 feedthrough
rlabel pdiffusion 360 -314 360 -314 0 cellNo=297
rlabel pdiffusion 367 -314 367 -314 0 feedthrough
rlabel pdiffusion 374 -314 374 -314 0 feedthrough
rlabel pdiffusion 381 -314 381 -314 0 feedthrough
rlabel pdiffusion 388 -314 388 -314 0 feedthrough
rlabel pdiffusion 395 -314 395 -314 0 feedthrough
rlabel pdiffusion 402 -314 402 -314 0 feedthrough
rlabel pdiffusion 409 -314 409 -314 0 cellNo=346
rlabel pdiffusion 416 -314 416 -314 0 feedthrough
rlabel pdiffusion 423 -314 423 -314 0 cellNo=22
rlabel pdiffusion 430 -314 430 -314 0 feedthrough
rlabel pdiffusion 437 -314 437 -314 0 feedthrough
rlabel pdiffusion 444 -314 444 -314 0 feedthrough
rlabel pdiffusion 451 -314 451 -314 0 cellNo=315
rlabel pdiffusion 458 -314 458 -314 0 feedthrough
rlabel pdiffusion 465 -314 465 -314 0 feedthrough
rlabel pdiffusion 472 -314 472 -314 0 feedthrough
rlabel pdiffusion 479 -314 479 -314 0 feedthrough
rlabel pdiffusion 486 -314 486 -314 0 feedthrough
rlabel pdiffusion 493 -314 493 -314 0 feedthrough
rlabel pdiffusion 500 -314 500 -314 0 feedthrough
rlabel pdiffusion 507 -314 507 -314 0 feedthrough
rlabel pdiffusion 514 -314 514 -314 0 feedthrough
rlabel pdiffusion 521 -314 521 -314 0 feedthrough
rlabel pdiffusion 528 -314 528 -314 0 feedthrough
rlabel pdiffusion 535 -314 535 -314 0 feedthrough
rlabel pdiffusion 542 -314 542 -314 0 cellNo=156
rlabel pdiffusion 549 -314 549 -314 0 feedthrough
rlabel pdiffusion 556 -314 556 -314 0 feedthrough
rlabel pdiffusion 563 -314 563 -314 0 feedthrough
rlabel pdiffusion 570 -314 570 -314 0 feedthrough
rlabel pdiffusion 577 -314 577 -314 0 cellNo=359
rlabel pdiffusion 584 -314 584 -314 0 cellNo=592
rlabel pdiffusion 591 -314 591 -314 0 feedthrough
rlabel pdiffusion 598 -314 598 -314 0 feedthrough
rlabel pdiffusion 605 -314 605 -314 0 cellNo=390
rlabel pdiffusion 612 -314 612 -314 0 feedthrough
rlabel pdiffusion 619 -314 619 -314 0 feedthrough
rlabel pdiffusion 626 -314 626 -314 0 feedthrough
rlabel pdiffusion 633 -314 633 -314 0 feedthrough
rlabel pdiffusion 640 -314 640 -314 0 feedthrough
rlabel pdiffusion 647 -314 647 -314 0 feedthrough
rlabel pdiffusion 654 -314 654 -314 0 feedthrough
rlabel pdiffusion 661 -314 661 -314 0 feedthrough
rlabel pdiffusion 668 -314 668 -314 0 feedthrough
rlabel pdiffusion 675 -314 675 -314 0 feedthrough
rlabel pdiffusion 682 -314 682 -314 0 feedthrough
rlabel pdiffusion 689 -314 689 -314 0 feedthrough
rlabel pdiffusion 696 -314 696 -314 0 cellNo=553
rlabel pdiffusion 703 -314 703 -314 0 cellNo=295
rlabel pdiffusion 710 -314 710 -314 0 feedthrough
rlabel pdiffusion 717 -314 717 -314 0 feedthrough
rlabel pdiffusion 724 -314 724 -314 0 feedthrough
rlabel pdiffusion 731 -314 731 -314 0 feedthrough
rlabel pdiffusion 738 -314 738 -314 0 feedthrough
rlabel pdiffusion 745 -314 745 -314 0 feedthrough
rlabel pdiffusion 752 -314 752 -314 0 feedthrough
rlabel pdiffusion 759 -314 759 -314 0 cellNo=153
rlabel pdiffusion 766 -314 766 -314 0 feedthrough
rlabel pdiffusion 773 -314 773 -314 0 feedthrough
rlabel pdiffusion 780 -314 780 -314 0 feedthrough
rlabel pdiffusion 787 -314 787 -314 0 feedthrough
rlabel pdiffusion 794 -314 794 -314 0 feedthrough
rlabel pdiffusion 801 -314 801 -314 0 feedthrough
rlabel pdiffusion 808 -314 808 -314 0 feedthrough
rlabel pdiffusion 815 -314 815 -314 0 feedthrough
rlabel pdiffusion 822 -314 822 -314 0 feedthrough
rlabel pdiffusion 829 -314 829 -314 0 feedthrough
rlabel pdiffusion 836 -314 836 -314 0 feedthrough
rlabel pdiffusion 843 -314 843 -314 0 feedthrough
rlabel pdiffusion 850 -314 850 -314 0 feedthrough
rlabel pdiffusion 857 -314 857 -314 0 feedthrough
rlabel pdiffusion 864 -314 864 -314 0 feedthrough
rlabel pdiffusion 871 -314 871 -314 0 feedthrough
rlabel pdiffusion 878 -314 878 -314 0 feedthrough
rlabel pdiffusion 885 -314 885 -314 0 feedthrough
rlabel pdiffusion 892 -314 892 -314 0 feedthrough
rlabel pdiffusion 899 -314 899 -314 0 feedthrough
rlabel pdiffusion 906 -314 906 -314 0 feedthrough
rlabel pdiffusion 913 -314 913 -314 0 feedthrough
rlabel pdiffusion 920 -314 920 -314 0 feedthrough
rlabel pdiffusion 927 -314 927 -314 0 feedthrough
rlabel pdiffusion 934 -314 934 -314 0 feedthrough
rlabel pdiffusion 941 -314 941 -314 0 feedthrough
rlabel pdiffusion 948 -314 948 -314 0 feedthrough
rlabel pdiffusion 955 -314 955 -314 0 feedthrough
rlabel pdiffusion 962 -314 962 -314 0 feedthrough
rlabel pdiffusion 969 -314 969 -314 0 feedthrough
rlabel pdiffusion 976 -314 976 -314 0 feedthrough
rlabel pdiffusion 983 -314 983 -314 0 feedthrough
rlabel pdiffusion 990 -314 990 -314 0 feedthrough
rlabel pdiffusion 997 -314 997 -314 0 feedthrough
rlabel pdiffusion 1004 -314 1004 -314 0 feedthrough
rlabel pdiffusion 1011 -314 1011 -314 0 feedthrough
rlabel pdiffusion 1018 -314 1018 -314 0 feedthrough
rlabel pdiffusion 1025 -314 1025 -314 0 feedthrough
rlabel pdiffusion 1032 -314 1032 -314 0 feedthrough
rlabel pdiffusion 1039 -314 1039 -314 0 feedthrough
rlabel pdiffusion 1046 -314 1046 -314 0 feedthrough
rlabel pdiffusion 1053 -314 1053 -314 0 feedthrough
rlabel pdiffusion 1060 -314 1060 -314 0 feedthrough
rlabel pdiffusion 1067 -314 1067 -314 0 feedthrough
rlabel pdiffusion 1074 -314 1074 -314 0 feedthrough
rlabel pdiffusion 1081 -314 1081 -314 0 feedthrough
rlabel pdiffusion 1088 -314 1088 -314 0 feedthrough
rlabel pdiffusion 1095 -314 1095 -314 0 feedthrough
rlabel pdiffusion 1102 -314 1102 -314 0 feedthrough
rlabel pdiffusion 1109 -314 1109 -314 0 feedthrough
rlabel pdiffusion 1116 -314 1116 -314 0 feedthrough
rlabel pdiffusion 1123 -314 1123 -314 0 feedthrough
rlabel pdiffusion 1130 -314 1130 -314 0 feedthrough
rlabel pdiffusion 1137 -314 1137 -314 0 feedthrough
rlabel pdiffusion 1144 -314 1144 -314 0 feedthrough
rlabel pdiffusion 1151 -314 1151 -314 0 cellNo=516
rlabel pdiffusion 1179 -314 1179 -314 0 feedthrough
rlabel pdiffusion 1501 -314 1501 -314 0 feedthrough
rlabel pdiffusion 3 -403 3 -403 0 feedthrough
rlabel pdiffusion 10 -403 10 -403 0 feedthrough
rlabel pdiffusion 17 -403 17 -403 0 feedthrough
rlabel pdiffusion 24 -403 24 -403 0 cellNo=261
rlabel pdiffusion 31 -403 31 -403 0 feedthrough
rlabel pdiffusion 38 -403 38 -403 0 cellNo=9
rlabel pdiffusion 45 -403 45 -403 0 cellNo=26
rlabel pdiffusion 52 -403 52 -403 0 feedthrough
rlabel pdiffusion 59 -403 59 -403 0 cellNo=506
rlabel pdiffusion 66 -403 66 -403 0 feedthrough
rlabel pdiffusion 73 -403 73 -403 0 cellNo=35
rlabel pdiffusion 80 -403 80 -403 0 cellNo=356
rlabel pdiffusion 87 -403 87 -403 0 cellNo=466
rlabel pdiffusion 94 -403 94 -403 0 feedthrough
rlabel pdiffusion 101 -403 101 -403 0 feedthrough
rlabel pdiffusion 108 -403 108 -403 0 feedthrough
rlabel pdiffusion 115 -403 115 -403 0 feedthrough
rlabel pdiffusion 122 -403 122 -403 0 cellNo=65
rlabel pdiffusion 129 -403 129 -403 0 feedthrough
rlabel pdiffusion 136 -403 136 -403 0 feedthrough
rlabel pdiffusion 143 -403 143 -403 0 feedthrough
rlabel pdiffusion 150 -403 150 -403 0 feedthrough
rlabel pdiffusion 157 -403 157 -403 0 feedthrough
rlabel pdiffusion 164 -403 164 -403 0 feedthrough
rlabel pdiffusion 171 -403 171 -403 0 feedthrough
rlabel pdiffusion 178 -403 178 -403 0 feedthrough
rlabel pdiffusion 185 -403 185 -403 0 feedthrough
rlabel pdiffusion 192 -403 192 -403 0 feedthrough
rlabel pdiffusion 199 -403 199 -403 0 feedthrough
rlabel pdiffusion 206 -403 206 -403 0 feedthrough
rlabel pdiffusion 213 -403 213 -403 0 feedthrough
rlabel pdiffusion 220 -403 220 -403 0 feedthrough
rlabel pdiffusion 227 -403 227 -403 0 feedthrough
rlabel pdiffusion 234 -403 234 -403 0 feedthrough
rlabel pdiffusion 241 -403 241 -403 0 feedthrough
rlabel pdiffusion 248 -403 248 -403 0 feedthrough
rlabel pdiffusion 255 -403 255 -403 0 feedthrough
rlabel pdiffusion 262 -403 262 -403 0 cellNo=314
rlabel pdiffusion 269 -403 269 -403 0 feedthrough
rlabel pdiffusion 276 -403 276 -403 0 feedthrough
rlabel pdiffusion 283 -403 283 -403 0 feedthrough
rlabel pdiffusion 290 -403 290 -403 0 cellNo=533
rlabel pdiffusion 297 -403 297 -403 0 feedthrough
rlabel pdiffusion 304 -403 304 -403 0 feedthrough
rlabel pdiffusion 311 -403 311 -403 0 feedthrough
rlabel pdiffusion 318 -403 318 -403 0 feedthrough
rlabel pdiffusion 325 -403 325 -403 0 feedthrough
rlabel pdiffusion 332 -403 332 -403 0 feedthrough
rlabel pdiffusion 339 -403 339 -403 0 feedthrough
rlabel pdiffusion 346 -403 346 -403 0 feedthrough
rlabel pdiffusion 353 -403 353 -403 0 feedthrough
rlabel pdiffusion 360 -403 360 -403 0 feedthrough
rlabel pdiffusion 367 -403 367 -403 0 feedthrough
rlabel pdiffusion 374 -403 374 -403 0 feedthrough
rlabel pdiffusion 381 -403 381 -403 0 feedthrough
rlabel pdiffusion 388 -403 388 -403 0 feedthrough
rlabel pdiffusion 395 -403 395 -403 0 cellNo=54
rlabel pdiffusion 402 -403 402 -403 0 feedthrough
rlabel pdiffusion 409 -403 409 -403 0 cellNo=327
rlabel pdiffusion 416 -403 416 -403 0 feedthrough
rlabel pdiffusion 423 -403 423 -403 0 feedthrough
rlabel pdiffusion 430 -403 430 -403 0 feedthrough
rlabel pdiffusion 437 -403 437 -403 0 feedthrough
rlabel pdiffusion 444 -403 444 -403 0 feedthrough
rlabel pdiffusion 451 -403 451 -403 0 feedthrough
rlabel pdiffusion 458 -403 458 -403 0 feedthrough
rlabel pdiffusion 465 -403 465 -403 0 feedthrough
rlabel pdiffusion 472 -403 472 -403 0 feedthrough
rlabel pdiffusion 479 -403 479 -403 0 feedthrough
rlabel pdiffusion 486 -403 486 -403 0 feedthrough
rlabel pdiffusion 493 -403 493 -403 0 feedthrough
rlabel pdiffusion 500 -403 500 -403 0 cellNo=227
rlabel pdiffusion 507 -403 507 -403 0 cellNo=237
rlabel pdiffusion 514 -403 514 -403 0 cellNo=69
rlabel pdiffusion 521 -403 521 -403 0 feedthrough
rlabel pdiffusion 528 -403 528 -403 0 feedthrough
rlabel pdiffusion 535 -403 535 -403 0 feedthrough
rlabel pdiffusion 542 -403 542 -403 0 feedthrough
rlabel pdiffusion 549 -403 549 -403 0 cellNo=134
rlabel pdiffusion 556 -403 556 -403 0 feedthrough
rlabel pdiffusion 563 -403 563 -403 0 cellNo=249
rlabel pdiffusion 570 -403 570 -403 0 cellNo=70
rlabel pdiffusion 577 -403 577 -403 0 feedthrough
rlabel pdiffusion 584 -403 584 -403 0 feedthrough
rlabel pdiffusion 591 -403 591 -403 0 cellNo=102
rlabel pdiffusion 598 -403 598 -403 0 feedthrough
rlabel pdiffusion 605 -403 605 -403 0 feedthrough
rlabel pdiffusion 612 -403 612 -403 0 feedthrough
rlabel pdiffusion 619 -403 619 -403 0 feedthrough
rlabel pdiffusion 626 -403 626 -403 0 feedthrough
rlabel pdiffusion 633 -403 633 -403 0 feedthrough
rlabel pdiffusion 640 -403 640 -403 0 cellNo=591
rlabel pdiffusion 647 -403 647 -403 0 feedthrough
rlabel pdiffusion 654 -403 654 -403 0 feedthrough
rlabel pdiffusion 661 -403 661 -403 0 cellNo=7
rlabel pdiffusion 668 -403 668 -403 0 cellNo=77
rlabel pdiffusion 675 -403 675 -403 0 feedthrough
rlabel pdiffusion 682 -403 682 -403 0 feedthrough
rlabel pdiffusion 689 -403 689 -403 0 feedthrough
rlabel pdiffusion 696 -403 696 -403 0 feedthrough
rlabel pdiffusion 703 -403 703 -403 0 feedthrough
rlabel pdiffusion 710 -403 710 -403 0 feedthrough
rlabel pdiffusion 717 -403 717 -403 0 feedthrough
rlabel pdiffusion 724 -403 724 -403 0 feedthrough
rlabel pdiffusion 731 -403 731 -403 0 feedthrough
rlabel pdiffusion 738 -403 738 -403 0 feedthrough
rlabel pdiffusion 745 -403 745 -403 0 feedthrough
rlabel pdiffusion 752 -403 752 -403 0 feedthrough
rlabel pdiffusion 759 -403 759 -403 0 feedthrough
rlabel pdiffusion 766 -403 766 -403 0 feedthrough
rlabel pdiffusion 773 -403 773 -403 0 feedthrough
rlabel pdiffusion 780 -403 780 -403 0 feedthrough
rlabel pdiffusion 787 -403 787 -403 0 feedthrough
rlabel pdiffusion 794 -403 794 -403 0 feedthrough
rlabel pdiffusion 801 -403 801 -403 0 feedthrough
rlabel pdiffusion 808 -403 808 -403 0 feedthrough
rlabel pdiffusion 815 -403 815 -403 0 feedthrough
rlabel pdiffusion 822 -403 822 -403 0 feedthrough
rlabel pdiffusion 829 -403 829 -403 0 feedthrough
rlabel pdiffusion 836 -403 836 -403 0 feedthrough
rlabel pdiffusion 843 -403 843 -403 0 feedthrough
rlabel pdiffusion 850 -403 850 -403 0 feedthrough
rlabel pdiffusion 857 -403 857 -403 0 feedthrough
rlabel pdiffusion 864 -403 864 -403 0 feedthrough
rlabel pdiffusion 871 -403 871 -403 0 feedthrough
rlabel pdiffusion 878 -403 878 -403 0 feedthrough
rlabel pdiffusion 885 -403 885 -403 0 feedthrough
rlabel pdiffusion 892 -403 892 -403 0 feedthrough
rlabel pdiffusion 899 -403 899 -403 0 feedthrough
rlabel pdiffusion 906 -403 906 -403 0 feedthrough
rlabel pdiffusion 913 -403 913 -403 0 feedthrough
rlabel pdiffusion 920 -403 920 -403 0 feedthrough
rlabel pdiffusion 927 -403 927 -403 0 feedthrough
rlabel pdiffusion 934 -403 934 -403 0 feedthrough
rlabel pdiffusion 941 -403 941 -403 0 feedthrough
rlabel pdiffusion 948 -403 948 -403 0 feedthrough
rlabel pdiffusion 955 -403 955 -403 0 feedthrough
rlabel pdiffusion 962 -403 962 -403 0 feedthrough
rlabel pdiffusion 969 -403 969 -403 0 feedthrough
rlabel pdiffusion 976 -403 976 -403 0 feedthrough
rlabel pdiffusion 983 -403 983 -403 0 feedthrough
rlabel pdiffusion 990 -403 990 -403 0 feedthrough
rlabel pdiffusion 997 -403 997 -403 0 feedthrough
rlabel pdiffusion 1004 -403 1004 -403 0 feedthrough
rlabel pdiffusion 1011 -403 1011 -403 0 feedthrough
rlabel pdiffusion 1018 -403 1018 -403 0 feedthrough
rlabel pdiffusion 1025 -403 1025 -403 0 feedthrough
rlabel pdiffusion 1032 -403 1032 -403 0 feedthrough
rlabel pdiffusion 1039 -403 1039 -403 0 feedthrough
rlabel pdiffusion 1046 -403 1046 -403 0 feedthrough
rlabel pdiffusion 1053 -403 1053 -403 0 feedthrough
rlabel pdiffusion 1060 -403 1060 -403 0 feedthrough
rlabel pdiffusion 1067 -403 1067 -403 0 feedthrough
rlabel pdiffusion 1074 -403 1074 -403 0 feedthrough
rlabel pdiffusion 1081 -403 1081 -403 0 feedthrough
rlabel pdiffusion 1088 -403 1088 -403 0 feedthrough
rlabel pdiffusion 1095 -403 1095 -403 0 feedthrough
rlabel pdiffusion 1102 -403 1102 -403 0 feedthrough
rlabel pdiffusion 1109 -403 1109 -403 0 feedthrough
rlabel pdiffusion 1116 -403 1116 -403 0 feedthrough
rlabel pdiffusion 1123 -403 1123 -403 0 feedthrough
rlabel pdiffusion 1130 -403 1130 -403 0 feedthrough
rlabel pdiffusion 1137 -403 1137 -403 0 feedthrough
rlabel pdiffusion 1144 -403 1144 -403 0 feedthrough
rlabel pdiffusion 1151 -403 1151 -403 0 feedthrough
rlabel pdiffusion 1158 -403 1158 -403 0 feedthrough
rlabel pdiffusion 1165 -403 1165 -403 0 feedthrough
rlabel pdiffusion 1172 -403 1172 -403 0 feedthrough
rlabel pdiffusion 1179 -403 1179 -403 0 feedthrough
rlabel pdiffusion 1186 -403 1186 -403 0 feedthrough
rlabel pdiffusion 1193 -403 1193 -403 0 feedthrough
rlabel pdiffusion 1200 -403 1200 -403 0 cellNo=457
rlabel pdiffusion 1207 -403 1207 -403 0 cellNo=14
rlabel pdiffusion 1501 -403 1501 -403 0 feedthrough
rlabel pdiffusion 3 -518 3 -518 0 cellNo=233
rlabel pdiffusion 10 -518 10 -518 0 feedthrough
rlabel pdiffusion 17 -518 17 -518 0 feedthrough
rlabel pdiffusion 24 -518 24 -518 0 feedthrough
rlabel pdiffusion 31 -518 31 -518 0 cellNo=4
rlabel pdiffusion 38 -518 38 -518 0 cellNo=481
rlabel pdiffusion 45 -518 45 -518 0 feedthrough
rlabel pdiffusion 52 -518 52 -518 0 feedthrough
rlabel pdiffusion 59 -518 59 -518 0 feedthrough
rlabel pdiffusion 66 -518 66 -518 0 feedthrough
rlabel pdiffusion 73 -518 73 -518 0 cellNo=322
rlabel pdiffusion 80 -518 80 -518 0 feedthrough
rlabel pdiffusion 87 -518 87 -518 0 cellNo=333
rlabel pdiffusion 94 -518 94 -518 0 feedthrough
rlabel pdiffusion 101 -518 101 -518 0 feedthrough
rlabel pdiffusion 108 -518 108 -518 0 cellNo=206
rlabel pdiffusion 115 -518 115 -518 0 feedthrough
rlabel pdiffusion 122 -518 122 -518 0 feedthrough
rlabel pdiffusion 129 -518 129 -518 0 feedthrough
rlabel pdiffusion 136 -518 136 -518 0 cellNo=59
rlabel pdiffusion 143 -518 143 -518 0 cellNo=446
rlabel pdiffusion 150 -518 150 -518 0 feedthrough
rlabel pdiffusion 157 -518 157 -518 0 cellNo=267
rlabel pdiffusion 164 -518 164 -518 0 feedthrough
rlabel pdiffusion 171 -518 171 -518 0 feedthrough
rlabel pdiffusion 178 -518 178 -518 0 feedthrough
rlabel pdiffusion 185 -518 185 -518 0 feedthrough
rlabel pdiffusion 192 -518 192 -518 0 feedthrough
rlabel pdiffusion 199 -518 199 -518 0 cellNo=55
rlabel pdiffusion 206 -518 206 -518 0 feedthrough
rlabel pdiffusion 213 -518 213 -518 0 feedthrough
rlabel pdiffusion 220 -518 220 -518 0 feedthrough
rlabel pdiffusion 227 -518 227 -518 0 feedthrough
rlabel pdiffusion 234 -518 234 -518 0 feedthrough
rlabel pdiffusion 241 -518 241 -518 0 feedthrough
rlabel pdiffusion 248 -518 248 -518 0 cellNo=329
rlabel pdiffusion 255 -518 255 -518 0 cellNo=107
rlabel pdiffusion 262 -518 262 -518 0 feedthrough
rlabel pdiffusion 269 -518 269 -518 0 feedthrough
rlabel pdiffusion 276 -518 276 -518 0 feedthrough
rlabel pdiffusion 283 -518 283 -518 0 feedthrough
rlabel pdiffusion 290 -518 290 -518 0 feedthrough
rlabel pdiffusion 297 -518 297 -518 0 feedthrough
rlabel pdiffusion 304 -518 304 -518 0 feedthrough
rlabel pdiffusion 311 -518 311 -518 0 feedthrough
rlabel pdiffusion 318 -518 318 -518 0 feedthrough
rlabel pdiffusion 325 -518 325 -518 0 feedthrough
rlabel pdiffusion 332 -518 332 -518 0 feedthrough
rlabel pdiffusion 339 -518 339 -518 0 feedthrough
rlabel pdiffusion 346 -518 346 -518 0 feedthrough
rlabel pdiffusion 353 -518 353 -518 0 feedthrough
rlabel pdiffusion 360 -518 360 -518 0 feedthrough
rlabel pdiffusion 367 -518 367 -518 0 feedthrough
rlabel pdiffusion 374 -518 374 -518 0 feedthrough
rlabel pdiffusion 381 -518 381 -518 0 cellNo=238
rlabel pdiffusion 388 -518 388 -518 0 feedthrough
rlabel pdiffusion 395 -518 395 -518 0 feedthrough
rlabel pdiffusion 402 -518 402 -518 0 feedthrough
rlabel pdiffusion 409 -518 409 -518 0 feedthrough
rlabel pdiffusion 416 -518 416 -518 0 cellNo=469
rlabel pdiffusion 423 -518 423 -518 0 cellNo=51
rlabel pdiffusion 430 -518 430 -518 0 feedthrough
rlabel pdiffusion 437 -518 437 -518 0 feedthrough
rlabel pdiffusion 444 -518 444 -518 0 feedthrough
rlabel pdiffusion 451 -518 451 -518 0 feedthrough
rlabel pdiffusion 458 -518 458 -518 0 cellNo=374
rlabel pdiffusion 465 -518 465 -518 0 feedthrough
rlabel pdiffusion 472 -518 472 -518 0 feedthrough
rlabel pdiffusion 479 -518 479 -518 0 feedthrough
rlabel pdiffusion 486 -518 486 -518 0 feedthrough
rlabel pdiffusion 493 -518 493 -518 0 feedthrough
rlabel pdiffusion 500 -518 500 -518 0 cellNo=579
rlabel pdiffusion 507 -518 507 -518 0 cellNo=416
rlabel pdiffusion 514 -518 514 -518 0 feedthrough
rlabel pdiffusion 521 -518 521 -518 0 feedthrough
rlabel pdiffusion 528 -518 528 -518 0 cellNo=536
rlabel pdiffusion 535 -518 535 -518 0 cellNo=56
rlabel pdiffusion 542 -518 542 -518 0 feedthrough
rlabel pdiffusion 549 -518 549 -518 0 feedthrough
rlabel pdiffusion 556 -518 556 -518 0 feedthrough
rlabel pdiffusion 563 -518 563 -518 0 feedthrough
rlabel pdiffusion 570 -518 570 -518 0 feedthrough
rlabel pdiffusion 577 -518 577 -518 0 feedthrough
rlabel pdiffusion 584 -518 584 -518 0 feedthrough
rlabel pdiffusion 591 -518 591 -518 0 feedthrough
rlabel pdiffusion 598 -518 598 -518 0 cellNo=219
rlabel pdiffusion 605 -518 605 -518 0 feedthrough
rlabel pdiffusion 612 -518 612 -518 0 cellNo=104
rlabel pdiffusion 619 -518 619 -518 0 feedthrough
rlabel pdiffusion 626 -518 626 -518 0 feedthrough
rlabel pdiffusion 633 -518 633 -518 0 feedthrough
rlabel pdiffusion 640 -518 640 -518 0 feedthrough
rlabel pdiffusion 647 -518 647 -518 0 feedthrough
rlabel pdiffusion 654 -518 654 -518 0 feedthrough
rlabel pdiffusion 661 -518 661 -518 0 cellNo=160
rlabel pdiffusion 668 -518 668 -518 0 feedthrough
rlabel pdiffusion 675 -518 675 -518 0 feedthrough
rlabel pdiffusion 682 -518 682 -518 0 feedthrough
rlabel pdiffusion 689 -518 689 -518 0 feedthrough
rlabel pdiffusion 696 -518 696 -518 0 cellNo=400
rlabel pdiffusion 703 -518 703 -518 0 cellNo=283
rlabel pdiffusion 710 -518 710 -518 0 feedthrough
rlabel pdiffusion 717 -518 717 -518 0 feedthrough
rlabel pdiffusion 724 -518 724 -518 0 feedthrough
rlabel pdiffusion 731 -518 731 -518 0 feedthrough
rlabel pdiffusion 738 -518 738 -518 0 feedthrough
rlabel pdiffusion 745 -518 745 -518 0 feedthrough
rlabel pdiffusion 752 -518 752 -518 0 feedthrough
rlabel pdiffusion 759 -518 759 -518 0 feedthrough
rlabel pdiffusion 766 -518 766 -518 0 feedthrough
rlabel pdiffusion 773 -518 773 -518 0 feedthrough
rlabel pdiffusion 780 -518 780 -518 0 feedthrough
rlabel pdiffusion 787 -518 787 -518 0 feedthrough
rlabel pdiffusion 794 -518 794 -518 0 feedthrough
rlabel pdiffusion 801 -518 801 -518 0 feedthrough
rlabel pdiffusion 808 -518 808 -518 0 feedthrough
rlabel pdiffusion 815 -518 815 -518 0 feedthrough
rlabel pdiffusion 822 -518 822 -518 0 feedthrough
rlabel pdiffusion 829 -518 829 -518 0 feedthrough
rlabel pdiffusion 836 -518 836 -518 0 feedthrough
rlabel pdiffusion 843 -518 843 -518 0 feedthrough
rlabel pdiffusion 850 -518 850 -518 0 feedthrough
rlabel pdiffusion 857 -518 857 -518 0 feedthrough
rlabel pdiffusion 864 -518 864 -518 0 feedthrough
rlabel pdiffusion 871 -518 871 -518 0 feedthrough
rlabel pdiffusion 878 -518 878 -518 0 feedthrough
rlabel pdiffusion 885 -518 885 -518 0 feedthrough
rlabel pdiffusion 892 -518 892 -518 0 feedthrough
rlabel pdiffusion 899 -518 899 -518 0 feedthrough
rlabel pdiffusion 906 -518 906 -518 0 feedthrough
rlabel pdiffusion 913 -518 913 -518 0 feedthrough
rlabel pdiffusion 920 -518 920 -518 0 feedthrough
rlabel pdiffusion 927 -518 927 -518 0 feedthrough
rlabel pdiffusion 934 -518 934 -518 0 feedthrough
rlabel pdiffusion 941 -518 941 -518 0 feedthrough
rlabel pdiffusion 948 -518 948 -518 0 feedthrough
rlabel pdiffusion 955 -518 955 -518 0 feedthrough
rlabel pdiffusion 962 -518 962 -518 0 feedthrough
rlabel pdiffusion 969 -518 969 -518 0 feedthrough
rlabel pdiffusion 976 -518 976 -518 0 feedthrough
rlabel pdiffusion 983 -518 983 -518 0 feedthrough
rlabel pdiffusion 990 -518 990 -518 0 feedthrough
rlabel pdiffusion 997 -518 997 -518 0 feedthrough
rlabel pdiffusion 1004 -518 1004 -518 0 feedthrough
rlabel pdiffusion 1011 -518 1011 -518 0 feedthrough
rlabel pdiffusion 1018 -518 1018 -518 0 feedthrough
rlabel pdiffusion 1025 -518 1025 -518 0 feedthrough
rlabel pdiffusion 1032 -518 1032 -518 0 feedthrough
rlabel pdiffusion 1039 -518 1039 -518 0 feedthrough
rlabel pdiffusion 1046 -518 1046 -518 0 feedthrough
rlabel pdiffusion 1053 -518 1053 -518 0 feedthrough
rlabel pdiffusion 1060 -518 1060 -518 0 feedthrough
rlabel pdiffusion 1067 -518 1067 -518 0 feedthrough
rlabel pdiffusion 1074 -518 1074 -518 0 feedthrough
rlabel pdiffusion 1081 -518 1081 -518 0 feedthrough
rlabel pdiffusion 1088 -518 1088 -518 0 feedthrough
rlabel pdiffusion 1095 -518 1095 -518 0 feedthrough
rlabel pdiffusion 1102 -518 1102 -518 0 feedthrough
rlabel pdiffusion 1109 -518 1109 -518 0 feedthrough
rlabel pdiffusion 1116 -518 1116 -518 0 feedthrough
rlabel pdiffusion 1123 -518 1123 -518 0 feedthrough
rlabel pdiffusion 1130 -518 1130 -518 0 feedthrough
rlabel pdiffusion 1137 -518 1137 -518 0 feedthrough
rlabel pdiffusion 1144 -518 1144 -518 0 feedthrough
rlabel pdiffusion 1151 -518 1151 -518 0 feedthrough
rlabel pdiffusion 1158 -518 1158 -518 0 feedthrough
rlabel pdiffusion 1165 -518 1165 -518 0 feedthrough
rlabel pdiffusion 1172 -518 1172 -518 0 feedthrough
rlabel pdiffusion 1179 -518 1179 -518 0 feedthrough
rlabel pdiffusion 1186 -518 1186 -518 0 feedthrough
rlabel pdiffusion 1193 -518 1193 -518 0 feedthrough
rlabel pdiffusion 1200 -518 1200 -518 0 feedthrough
rlabel pdiffusion 1207 -518 1207 -518 0 feedthrough
rlabel pdiffusion 1214 -518 1214 -518 0 feedthrough
rlabel pdiffusion 1221 -518 1221 -518 0 feedthrough
rlabel pdiffusion 1228 -518 1228 -518 0 feedthrough
rlabel pdiffusion 1235 -518 1235 -518 0 feedthrough
rlabel pdiffusion 1242 -518 1242 -518 0 feedthrough
rlabel pdiffusion 1249 -518 1249 -518 0 feedthrough
rlabel pdiffusion 1256 -518 1256 -518 0 feedthrough
rlabel pdiffusion 1263 -518 1263 -518 0 feedthrough
rlabel pdiffusion 1396 -518 1396 -518 0 feedthrough
rlabel pdiffusion 1501 -518 1501 -518 0 feedthrough
rlabel pdiffusion 3 -633 3 -633 0 feedthrough
rlabel pdiffusion 10 -633 10 -633 0 feedthrough
rlabel pdiffusion 17 -633 17 -633 0 cellNo=258
rlabel pdiffusion 24 -633 24 -633 0 feedthrough
rlabel pdiffusion 31 -633 31 -633 0 feedthrough
rlabel pdiffusion 38 -633 38 -633 0 cellNo=116
rlabel pdiffusion 45 -633 45 -633 0 cellNo=422
rlabel pdiffusion 52 -633 52 -633 0 feedthrough
rlabel pdiffusion 59 -633 59 -633 0 feedthrough
rlabel pdiffusion 66 -633 66 -633 0 feedthrough
rlabel pdiffusion 73 -633 73 -633 0 cellNo=263
rlabel pdiffusion 80 -633 80 -633 0 feedthrough
rlabel pdiffusion 87 -633 87 -633 0 feedthrough
rlabel pdiffusion 94 -633 94 -633 0 cellNo=437
rlabel pdiffusion 101 -633 101 -633 0 feedthrough
rlabel pdiffusion 108 -633 108 -633 0 feedthrough
rlabel pdiffusion 115 -633 115 -633 0 cellNo=419
rlabel pdiffusion 122 -633 122 -633 0 feedthrough
rlabel pdiffusion 129 -633 129 -633 0 feedthrough
rlabel pdiffusion 136 -633 136 -633 0 feedthrough
rlabel pdiffusion 143 -633 143 -633 0 feedthrough
rlabel pdiffusion 150 -633 150 -633 0 feedthrough
rlabel pdiffusion 157 -633 157 -633 0 feedthrough
rlabel pdiffusion 164 -633 164 -633 0 feedthrough
rlabel pdiffusion 171 -633 171 -633 0 cellNo=126
rlabel pdiffusion 178 -633 178 -633 0 feedthrough
rlabel pdiffusion 185 -633 185 -633 0 feedthrough
rlabel pdiffusion 192 -633 192 -633 0 feedthrough
rlabel pdiffusion 199 -633 199 -633 0 feedthrough
rlabel pdiffusion 206 -633 206 -633 0 feedthrough
rlabel pdiffusion 213 -633 213 -633 0 feedthrough
rlabel pdiffusion 220 -633 220 -633 0 feedthrough
rlabel pdiffusion 227 -633 227 -633 0 feedthrough
rlabel pdiffusion 234 -633 234 -633 0 feedthrough
rlabel pdiffusion 241 -633 241 -633 0 feedthrough
rlabel pdiffusion 248 -633 248 -633 0 feedthrough
rlabel pdiffusion 255 -633 255 -633 0 feedthrough
rlabel pdiffusion 262 -633 262 -633 0 feedthrough
rlabel pdiffusion 269 -633 269 -633 0 cellNo=18
rlabel pdiffusion 276 -633 276 -633 0 feedthrough
rlabel pdiffusion 283 -633 283 -633 0 feedthrough
rlabel pdiffusion 290 -633 290 -633 0 feedthrough
rlabel pdiffusion 297 -633 297 -633 0 feedthrough
rlabel pdiffusion 304 -633 304 -633 0 feedthrough
rlabel pdiffusion 311 -633 311 -633 0 cellNo=496
rlabel pdiffusion 318 -633 318 -633 0 feedthrough
rlabel pdiffusion 325 -633 325 -633 0 feedthrough
rlabel pdiffusion 332 -633 332 -633 0 feedthrough
rlabel pdiffusion 339 -633 339 -633 0 feedthrough
rlabel pdiffusion 346 -633 346 -633 0 cellNo=386
rlabel pdiffusion 353 -633 353 -633 0 cellNo=247
rlabel pdiffusion 360 -633 360 -633 0 feedthrough
rlabel pdiffusion 367 -633 367 -633 0 feedthrough
rlabel pdiffusion 374 -633 374 -633 0 feedthrough
rlabel pdiffusion 381 -633 381 -633 0 cellNo=491
rlabel pdiffusion 388 -633 388 -633 0 cellNo=145
rlabel pdiffusion 395 -633 395 -633 0 feedthrough
rlabel pdiffusion 402 -633 402 -633 0 feedthrough
rlabel pdiffusion 409 -633 409 -633 0 feedthrough
rlabel pdiffusion 416 -633 416 -633 0 cellNo=410
rlabel pdiffusion 423 -633 423 -633 0 feedthrough
rlabel pdiffusion 430 -633 430 -633 0 feedthrough
rlabel pdiffusion 437 -633 437 -633 0 feedthrough
rlabel pdiffusion 444 -633 444 -633 0 cellNo=132
rlabel pdiffusion 451 -633 451 -633 0 feedthrough
rlabel pdiffusion 458 -633 458 -633 0 feedthrough
rlabel pdiffusion 465 -633 465 -633 0 feedthrough
rlabel pdiffusion 472 -633 472 -633 0 feedthrough
rlabel pdiffusion 479 -633 479 -633 0 cellNo=53
rlabel pdiffusion 486 -633 486 -633 0 feedthrough
rlabel pdiffusion 493 -633 493 -633 0 feedthrough
rlabel pdiffusion 500 -633 500 -633 0 feedthrough
rlabel pdiffusion 507 -633 507 -633 0 cellNo=423
rlabel pdiffusion 514 -633 514 -633 0 feedthrough
rlabel pdiffusion 521 -633 521 -633 0 feedthrough
rlabel pdiffusion 528 -633 528 -633 0 feedthrough
rlabel pdiffusion 535 -633 535 -633 0 feedthrough
rlabel pdiffusion 542 -633 542 -633 0 feedthrough
rlabel pdiffusion 549 -633 549 -633 0 feedthrough
rlabel pdiffusion 556 -633 556 -633 0 feedthrough
rlabel pdiffusion 563 -633 563 -633 0 cellNo=112
rlabel pdiffusion 570 -633 570 -633 0 feedthrough
rlabel pdiffusion 577 -633 577 -633 0 feedthrough
rlabel pdiffusion 584 -633 584 -633 0 feedthrough
rlabel pdiffusion 591 -633 591 -633 0 feedthrough
rlabel pdiffusion 598 -633 598 -633 0 feedthrough
rlabel pdiffusion 605 -633 605 -633 0 feedthrough
rlabel pdiffusion 612 -633 612 -633 0 cellNo=191
rlabel pdiffusion 619 -633 619 -633 0 feedthrough
rlabel pdiffusion 626 -633 626 -633 0 cellNo=337
rlabel pdiffusion 633 -633 633 -633 0 cellNo=348
rlabel pdiffusion 640 -633 640 -633 0 feedthrough
rlabel pdiffusion 647 -633 647 -633 0 feedthrough
rlabel pdiffusion 654 -633 654 -633 0 feedthrough
rlabel pdiffusion 661 -633 661 -633 0 feedthrough
rlabel pdiffusion 668 -633 668 -633 0 cellNo=113
rlabel pdiffusion 675 -633 675 -633 0 feedthrough
rlabel pdiffusion 682 -633 682 -633 0 feedthrough
rlabel pdiffusion 689 -633 689 -633 0 feedthrough
rlabel pdiffusion 696 -633 696 -633 0 feedthrough
rlabel pdiffusion 703 -633 703 -633 0 feedthrough
rlabel pdiffusion 710 -633 710 -633 0 feedthrough
rlabel pdiffusion 717 -633 717 -633 0 feedthrough
rlabel pdiffusion 724 -633 724 -633 0 feedthrough
rlabel pdiffusion 731 -633 731 -633 0 feedthrough
rlabel pdiffusion 738 -633 738 -633 0 feedthrough
rlabel pdiffusion 745 -633 745 -633 0 cellNo=148
rlabel pdiffusion 752 -633 752 -633 0 feedthrough
rlabel pdiffusion 759 -633 759 -633 0 feedthrough
rlabel pdiffusion 766 -633 766 -633 0 feedthrough
rlabel pdiffusion 773 -633 773 -633 0 feedthrough
rlabel pdiffusion 780 -633 780 -633 0 feedthrough
rlabel pdiffusion 787 -633 787 -633 0 feedthrough
rlabel pdiffusion 794 -633 794 -633 0 feedthrough
rlabel pdiffusion 801 -633 801 -633 0 feedthrough
rlabel pdiffusion 808 -633 808 -633 0 feedthrough
rlabel pdiffusion 815 -633 815 -633 0 feedthrough
rlabel pdiffusion 822 -633 822 -633 0 feedthrough
rlabel pdiffusion 829 -633 829 -633 0 feedthrough
rlabel pdiffusion 836 -633 836 -633 0 feedthrough
rlabel pdiffusion 843 -633 843 -633 0 feedthrough
rlabel pdiffusion 850 -633 850 -633 0 feedthrough
rlabel pdiffusion 857 -633 857 -633 0 feedthrough
rlabel pdiffusion 864 -633 864 -633 0 feedthrough
rlabel pdiffusion 871 -633 871 -633 0 feedthrough
rlabel pdiffusion 878 -633 878 -633 0 feedthrough
rlabel pdiffusion 885 -633 885 -633 0 feedthrough
rlabel pdiffusion 892 -633 892 -633 0 feedthrough
rlabel pdiffusion 899 -633 899 -633 0 feedthrough
rlabel pdiffusion 906 -633 906 -633 0 feedthrough
rlabel pdiffusion 913 -633 913 -633 0 feedthrough
rlabel pdiffusion 920 -633 920 -633 0 feedthrough
rlabel pdiffusion 927 -633 927 -633 0 feedthrough
rlabel pdiffusion 934 -633 934 -633 0 feedthrough
rlabel pdiffusion 941 -633 941 -633 0 feedthrough
rlabel pdiffusion 948 -633 948 -633 0 feedthrough
rlabel pdiffusion 955 -633 955 -633 0 feedthrough
rlabel pdiffusion 962 -633 962 -633 0 cellNo=340
rlabel pdiffusion 969 -633 969 -633 0 feedthrough
rlabel pdiffusion 976 -633 976 -633 0 feedthrough
rlabel pdiffusion 983 -633 983 -633 0 feedthrough
rlabel pdiffusion 990 -633 990 -633 0 feedthrough
rlabel pdiffusion 997 -633 997 -633 0 feedthrough
rlabel pdiffusion 1004 -633 1004 -633 0 feedthrough
rlabel pdiffusion 1011 -633 1011 -633 0 feedthrough
rlabel pdiffusion 1018 -633 1018 -633 0 feedthrough
rlabel pdiffusion 1025 -633 1025 -633 0 feedthrough
rlabel pdiffusion 1032 -633 1032 -633 0 cellNo=60
rlabel pdiffusion 1039 -633 1039 -633 0 feedthrough
rlabel pdiffusion 1046 -633 1046 -633 0 feedthrough
rlabel pdiffusion 1053 -633 1053 -633 0 feedthrough
rlabel pdiffusion 1060 -633 1060 -633 0 feedthrough
rlabel pdiffusion 1067 -633 1067 -633 0 feedthrough
rlabel pdiffusion 1074 -633 1074 -633 0 feedthrough
rlabel pdiffusion 1081 -633 1081 -633 0 feedthrough
rlabel pdiffusion 1088 -633 1088 -633 0 feedthrough
rlabel pdiffusion 1095 -633 1095 -633 0 feedthrough
rlabel pdiffusion 1102 -633 1102 -633 0 feedthrough
rlabel pdiffusion 1109 -633 1109 -633 0 feedthrough
rlabel pdiffusion 1116 -633 1116 -633 0 feedthrough
rlabel pdiffusion 1123 -633 1123 -633 0 feedthrough
rlabel pdiffusion 1130 -633 1130 -633 0 feedthrough
rlabel pdiffusion 1137 -633 1137 -633 0 feedthrough
rlabel pdiffusion 1144 -633 1144 -633 0 feedthrough
rlabel pdiffusion 1151 -633 1151 -633 0 feedthrough
rlabel pdiffusion 1158 -633 1158 -633 0 feedthrough
rlabel pdiffusion 1165 -633 1165 -633 0 feedthrough
rlabel pdiffusion 1172 -633 1172 -633 0 feedthrough
rlabel pdiffusion 1179 -633 1179 -633 0 feedthrough
rlabel pdiffusion 1186 -633 1186 -633 0 feedthrough
rlabel pdiffusion 1193 -633 1193 -633 0 feedthrough
rlabel pdiffusion 1200 -633 1200 -633 0 feedthrough
rlabel pdiffusion 1207 -633 1207 -633 0 feedthrough
rlabel pdiffusion 1214 -633 1214 -633 0 feedthrough
rlabel pdiffusion 1221 -633 1221 -633 0 feedthrough
rlabel pdiffusion 1228 -633 1228 -633 0 feedthrough
rlabel pdiffusion 1235 -633 1235 -633 0 feedthrough
rlabel pdiffusion 1242 -633 1242 -633 0 feedthrough
rlabel pdiffusion 1249 -633 1249 -633 0 feedthrough
rlabel pdiffusion 1256 -633 1256 -633 0 feedthrough
rlabel pdiffusion 1263 -633 1263 -633 0 feedthrough
rlabel pdiffusion 1270 -633 1270 -633 0 feedthrough
rlabel pdiffusion 1277 -633 1277 -633 0 feedthrough
rlabel pdiffusion 1284 -633 1284 -633 0 feedthrough
rlabel pdiffusion 1291 -633 1291 -633 0 feedthrough
rlabel pdiffusion 1298 -633 1298 -633 0 feedthrough
rlabel pdiffusion 1305 -633 1305 -633 0 feedthrough
rlabel pdiffusion 1312 -633 1312 -633 0 feedthrough
rlabel pdiffusion 1319 -633 1319 -633 0 feedthrough
rlabel pdiffusion 1326 -633 1326 -633 0 feedthrough
rlabel pdiffusion 1333 -633 1333 -633 0 feedthrough
rlabel pdiffusion 1340 -633 1340 -633 0 feedthrough
rlabel pdiffusion 1347 -633 1347 -633 0 feedthrough
rlabel pdiffusion 1354 -633 1354 -633 0 feedthrough
rlabel pdiffusion 1361 -633 1361 -633 0 feedthrough
rlabel pdiffusion 1368 -633 1368 -633 0 feedthrough
rlabel pdiffusion 1375 -633 1375 -633 0 feedthrough
rlabel pdiffusion 1473 -633 1473 -633 0 feedthrough
rlabel pdiffusion 1508 -633 1508 -633 0 feedthrough
rlabel pdiffusion 3 -752 3 -752 0 cellNo=169
rlabel pdiffusion 10 -752 10 -752 0 cellNo=334
rlabel pdiffusion 17 -752 17 -752 0 feedthrough
rlabel pdiffusion 24 -752 24 -752 0 feedthrough
rlabel pdiffusion 31 -752 31 -752 0 feedthrough
rlabel pdiffusion 38 -752 38 -752 0 feedthrough
rlabel pdiffusion 45 -752 45 -752 0 feedthrough
rlabel pdiffusion 52 -752 52 -752 0 feedthrough
rlabel pdiffusion 59 -752 59 -752 0 cellNo=88
rlabel pdiffusion 66 -752 66 -752 0 feedthrough
rlabel pdiffusion 73 -752 73 -752 0 cellNo=125
rlabel pdiffusion 80 -752 80 -752 0 feedthrough
rlabel pdiffusion 87 -752 87 -752 0 feedthrough
rlabel pdiffusion 94 -752 94 -752 0 feedthrough
rlabel pdiffusion 101 -752 101 -752 0 cellNo=480
rlabel pdiffusion 108 -752 108 -752 0 feedthrough
rlabel pdiffusion 115 -752 115 -752 0 cellNo=385
rlabel pdiffusion 122 -752 122 -752 0 feedthrough
rlabel pdiffusion 129 -752 129 -752 0 feedthrough
rlabel pdiffusion 136 -752 136 -752 0 cellNo=99
rlabel pdiffusion 143 -752 143 -752 0 feedthrough
rlabel pdiffusion 150 -752 150 -752 0 feedthrough
rlabel pdiffusion 157 -752 157 -752 0 feedthrough
rlabel pdiffusion 164 -752 164 -752 0 feedthrough
rlabel pdiffusion 171 -752 171 -752 0 feedthrough
rlabel pdiffusion 178 -752 178 -752 0 feedthrough
rlabel pdiffusion 185 -752 185 -752 0 feedthrough
rlabel pdiffusion 192 -752 192 -752 0 feedthrough
rlabel pdiffusion 199 -752 199 -752 0 feedthrough
rlabel pdiffusion 206 -752 206 -752 0 feedthrough
rlabel pdiffusion 213 -752 213 -752 0 feedthrough
rlabel pdiffusion 220 -752 220 -752 0 feedthrough
rlabel pdiffusion 227 -752 227 -752 0 feedthrough
rlabel pdiffusion 234 -752 234 -752 0 feedthrough
rlabel pdiffusion 241 -752 241 -752 0 feedthrough
rlabel pdiffusion 248 -752 248 -752 0 feedthrough
rlabel pdiffusion 255 -752 255 -752 0 feedthrough
rlabel pdiffusion 262 -752 262 -752 0 feedthrough
rlabel pdiffusion 269 -752 269 -752 0 cellNo=157
rlabel pdiffusion 276 -752 276 -752 0 feedthrough
rlabel pdiffusion 283 -752 283 -752 0 feedthrough
rlabel pdiffusion 290 -752 290 -752 0 feedthrough
rlabel pdiffusion 297 -752 297 -752 0 feedthrough
rlabel pdiffusion 304 -752 304 -752 0 feedthrough
rlabel pdiffusion 311 -752 311 -752 0 feedthrough
rlabel pdiffusion 318 -752 318 -752 0 feedthrough
rlabel pdiffusion 325 -752 325 -752 0 feedthrough
rlabel pdiffusion 332 -752 332 -752 0 feedthrough
rlabel pdiffusion 339 -752 339 -752 0 feedthrough
rlabel pdiffusion 346 -752 346 -752 0 feedthrough
rlabel pdiffusion 353 -752 353 -752 0 cellNo=114
rlabel pdiffusion 360 -752 360 -752 0 feedthrough
rlabel pdiffusion 367 -752 367 -752 0 cellNo=20
rlabel pdiffusion 374 -752 374 -752 0 feedthrough
rlabel pdiffusion 381 -752 381 -752 0 feedthrough
rlabel pdiffusion 388 -752 388 -752 0 feedthrough
rlabel pdiffusion 395 -752 395 -752 0 feedthrough
rlabel pdiffusion 402 -752 402 -752 0 feedthrough
rlabel pdiffusion 409 -752 409 -752 0 feedthrough
rlabel pdiffusion 416 -752 416 -752 0 feedthrough
rlabel pdiffusion 423 -752 423 -752 0 cellNo=274
rlabel pdiffusion 430 -752 430 -752 0 feedthrough
rlabel pdiffusion 437 -752 437 -752 0 feedthrough
rlabel pdiffusion 444 -752 444 -752 0 feedthrough
rlabel pdiffusion 451 -752 451 -752 0 feedthrough
rlabel pdiffusion 458 -752 458 -752 0 feedthrough
rlabel pdiffusion 465 -752 465 -752 0 feedthrough
rlabel pdiffusion 472 -752 472 -752 0 feedthrough
rlabel pdiffusion 479 -752 479 -752 0 feedthrough
rlabel pdiffusion 486 -752 486 -752 0 feedthrough
rlabel pdiffusion 493 -752 493 -752 0 feedthrough
rlabel pdiffusion 500 -752 500 -752 0 feedthrough
rlabel pdiffusion 507 -752 507 -752 0 feedthrough
rlabel pdiffusion 514 -752 514 -752 0 feedthrough
rlabel pdiffusion 521 -752 521 -752 0 cellNo=66
rlabel pdiffusion 528 -752 528 -752 0 feedthrough
rlabel pdiffusion 535 -752 535 -752 0 cellNo=139
rlabel pdiffusion 542 -752 542 -752 0 cellNo=96
rlabel pdiffusion 549 -752 549 -752 0 feedthrough
rlabel pdiffusion 556 -752 556 -752 0 feedthrough
rlabel pdiffusion 563 -752 563 -752 0 cellNo=597
rlabel pdiffusion 570 -752 570 -752 0 feedthrough
rlabel pdiffusion 577 -752 577 -752 0 feedthrough
rlabel pdiffusion 584 -752 584 -752 0 feedthrough
rlabel pdiffusion 591 -752 591 -752 0 feedthrough
rlabel pdiffusion 598 -752 598 -752 0 cellNo=576
rlabel pdiffusion 605 -752 605 -752 0 feedthrough
rlabel pdiffusion 612 -752 612 -752 0 cellNo=202
rlabel pdiffusion 619 -752 619 -752 0 cellNo=24
rlabel pdiffusion 626 -752 626 -752 0 cellNo=207
rlabel pdiffusion 633 -752 633 -752 0 feedthrough
rlabel pdiffusion 640 -752 640 -752 0 feedthrough
rlabel pdiffusion 647 -752 647 -752 0 feedthrough
rlabel pdiffusion 654 -752 654 -752 0 feedthrough
rlabel pdiffusion 661 -752 661 -752 0 cellNo=354
rlabel pdiffusion 668 -752 668 -752 0 feedthrough
rlabel pdiffusion 675 -752 675 -752 0 feedthrough
rlabel pdiffusion 682 -752 682 -752 0 feedthrough
rlabel pdiffusion 689 -752 689 -752 0 feedthrough
rlabel pdiffusion 696 -752 696 -752 0 feedthrough
rlabel pdiffusion 703 -752 703 -752 0 feedthrough
rlabel pdiffusion 710 -752 710 -752 0 feedthrough
rlabel pdiffusion 717 -752 717 -752 0 feedthrough
rlabel pdiffusion 724 -752 724 -752 0 feedthrough
rlabel pdiffusion 731 -752 731 -752 0 feedthrough
rlabel pdiffusion 738 -752 738 -752 0 feedthrough
rlabel pdiffusion 745 -752 745 -752 0 cellNo=92
rlabel pdiffusion 752 -752 752 -752 0 feedthrough
rlabel pdiffusion 759 -752 759 -752 0 cellNo=6
rlabel pdiffusion 766 -752 766 -752 0 feedthrough
rlabel pdiffusion 773 -752 773 -752 0 cellNo=90
rlabel pdiffusion 780 -752 780 -752 0 feedthrough
rlabel pdiffusion 787 -752 787 -752 0 feedthrough
rlabel pdiffusion 794 -752 794 -752 0 feedthrough
rlabel pdiffusion 801 -752 801 -752 0 feedthrough
rlabel pdiffusion 808 -752 808 -752 0 feedthrough
rlabel pdiffusion 815 -752 815 -752 0 feedthrough
rlabel pdiffusion 822 -752 822 -752 0 feedthrough
rlabel pdiffusion 829 -752 829 -752 0 feedthrough
rlabel pdiffusion 836 -752 836 -752 0 feedthrough
rlabel pdiffusion 843 -752 843 -752 0 feedthrough
rlabel pdiffusion 850 -752 850 -752 0 feedthrough
rlabel pdiffusion 857 -752 857 -752 0 feedthrough
rlabel pdiffusion 864 -752 864 -752 0 feedthrough
rlabel pdiffusion 871 -752 871 -752 0 feedthrough
rlabel pdiffusion 878 -752 878 -752 0 feedthrough
rlabel pdiffusion 885 -752 885 -752 0 cellNo=254
rlabel pdiffusion 892 -752 892 -752 0 feedthrough
rlabel pdiffusion 899 -752 899 -752 0 feedthrough
rlabel pdiffusion 906 -752 906 -752 0 feedthrough
rlabel pdiffusion 913 -752 913 -752 0 feedthrough
rlabel pdiffusion 920 -752 920 -752 0 feedthrough
rlabel pdiffusion 927 -752 927 -752 0 feedthrough
rlabel pdiffusion 934 -752 934 -752 0 feedthrough
rlabel pdiffusion 941 -752 941 -752 0 cellNo=397
rlabel pdiffusion 948 -752 948 -752 0 feedthrough
rlabel pdiffusion 955 -752 955 -752 0 feedthrough
rlabel pdiffusion 962 -752 962 -752 0 feedthrough
rlabel pdiffusion 969 -752 969 -752 0 feedthrough
rlabel pdiffusion 976 -752 976 -752 0 feedthrough
rlabel pdiffusion 983 -752 983 -752 0 feedthrough
rlabel pdiffusion 990 -752 990 -752 0 feedthrough
rlabel pdiffusion 997 -752 997 -752 0 feedthrough
rlabel pdiffusion 1004 -752 1004 -752 0 feedthrough
rlabel pdiffusion 1011 -752 1011 -752 0 feedthrough
rlabel pdiffusion 1018 -752 1018 -752 0 feedthrough
rlabel pdiffusion 1025 -752 1025 -752 0 feedthrough
rlabel pdiffusion 1032 -752 1032 -752 0 feedthrough
rlabel pdiffusion 1039 -752 1039 -752 0 feedthrough
rlabel pdiffusion 1046 -752 1046 -752 0 feedthrough
rlabel pdiffusion 1053 -752 1053 -752 0 feedthrough
rlabel pdiffusion 1060 -752 1060 -752 0 feedthrough
rlabel pdiffusion 1067 -752 1067 -752 0 feedthrough
rlabel pdiffusion 1074 -752 1074 -752 0 feedthrough
rlabel pdiffusion 1081 -752 1081 -752 0 feedthrough
rlabel pdiffusion 1088 -752 1088 -752 0 feedthrough
rlabel pdiffusion 1095 -752 1095 -752 0 feedthrough
rlabel pdiffusion 1102 -752 1102 -752 0 feedthrough
rlabel pdiffusion 1109 -752 1109 -752 0 feedthrough
rlabel pdiffusion 1116 -752 1116 -752 0 feedthrough
rlabel pdiffusion 1123 -752 1123 -752 0 feedthrough
rlabel pdiffusion 1130 -752 1130 -752 0 feedthrough
rlabel pdiffusion 1137 -752 1137 -752 0 feedthrough
rlabel pdiffusion 1144 -752 1144 -752 0 feedthrough
rlabel pdiffusion 1151 -752 1151 -752 0 feedthrough
rlabel pdiffusion 1158 -752 1158 -752 0 feedthrough
rlabel pdiffusion 1165 -752 1165 -752 0 feedthrough
rlabel pdiffusion 1172 -752 1172 -752 0 feedthrough
rlabel pdiffusion 1179 -752 1179 -752 0 feedthrough
rlabel pdiffusion 1186 -752 1186 -752 0 feedthrough
rlabel pdiffusion 1193 -752 1193 -752 0 feedthrough
rlabel pdiffusion 1200 -752 1200 -752 0 feedthrough
rlabel pdiffusion 1207 -752 1207 -752 0 feedthrough
rlabel pdiffusion 1214 -752 1214 -752 0 feedthrough
rlabel pdiffusion 1221 -752 1221 -752 0 feedthrough
rlabel pdiffusion 1228 -752 1228 -752 0 feedthrough
rlabel pdiffusion 1235 -752 1235 -752 0 feedthrough
rlabel pdiffusion 1242 -752 1242 -752 0 feedthrough
rlabel pdiffusion 1249 -752 1249 -752 0 feedthrough
rlabel pdiffusion 1256 -752 1256 -752 0 feedthrough
rlabel pdiffusion 1263 -752 1263 -752 0 feedthrough
rlabel pdiffusion 1270 -752 1270 -752 0 feedthrough
rlabel pdiffusion 1277 -752 1277 -752 0 feedthrough
rlabel pdiffusion 1284 -752 1284 -752 0 feedthrough
rlabel pdiffusion 1291 -752 1291 -752 0 feedthrough
rlabel pdiffusion 1298 -752 1298 -752 0 feedthrough
rlabel pdiffusion 1305 -752 1305 -752 0 feedthrough
rlabel pdiffusion 1312 -752 1312 -752 0 feedthrough
rlabel pdiffusion 1319 -752 1319 -752 0 feedthrough
rlabel pdiffusion 1326 -752 1326 -752 0 feedthrough
rlabel pdiffusion 1333 -752 1333 -752 0 feedthrough
rlabel pdiffusion 1340 -752 1340 -752 0 feedthrough
rlabel pdiffusion 1347 -752 1347 -752 0 feedthrough
rlabel pdiffusion 1354 -752 1354 -752 0 feedthrough
rlabel pdiffusion 1361 -752 1361 -752 0 feedthrough
rlabel pdiffusion 1368 -752 1368 -752 0 feedthrough
rlabel pdiffusion 1375 -752 1375 -752 0 feedthrough
rlabel pdiffusion 1382 -752 1382 -752 0 feedthrough
rlabel pdiffusion 1389 -752 1389 -752 0 feedthrough
rlabel pdiffusion 1396 -752 1396 -752 0 feedthrough
rlabel pdiffusion 1403 -752 1403 -752 0 feedthrough
rlabel pdiffusion 1410 -752 1410 -752 0 feedthrough
rlabel pdiffusion 1417 -752 1417 -752 0 feedthrough
rlabel pdiffusion 1424 -752 1424 -752 0 feedthrough
rlabel pdiffusion 1431 -752 1431 -752 0 feedthrough
rlabel pdiffusion 1438 -752 1438 -752 0 feedthrough
rlabel pdiffusion 1445 -752 1445 -752 0 feedthrough
rlabel pdiffusion 1452 -752 1452 -752 0 feedthrough
rlabel pdiffusion 1459 -752 1459 -752 0 feedthrough
rlabel pdiffusion 1466 -752 1466 -752 0 feedthrough
rlabel pdiffusion 1473 -752 1473 -752 0 feedthrough
rlabel pdiffusion 1480 -752 1480 -752 0 feedthrough
rlabel pdiffusion 1487 -752 1487 -752 0 feedthrough
rlabel pdiffusion 1494 -752 1494 -752 0 feedthrough
rlabel pdiffusion 1501 -752 1501 -752 0 feedthrough
rlabel pdiffusion 1508 -752 1508 -752 0 feedthrough
rlabel pdiffusion 1515 -752 1515 -752 0 feedthrough
rlabel pdiffusion 1522 -752 1522 -752 0 feedthrough
rlabel pdiffusion 1529 -752 1529 -752 0 feedthrough
rlabel pdiffusion 3 -893 3 -893 0 feedthrough
rlabel pdiffusion 10 -893 10 -893 0 feedthrough
rlabel pdiffusion 17 -893 17 -893 0 feedthrough
rlabel pdiffusion 24 -893 24 -893 0 feedthrough
rlabel pdiffusion 31 -893 31 -893 0 feedthrough
rlabel pdiffusion 38 -893 38 -893 0 cellNo=5
rlabel pdiffusion 45 -893 45 -893 0 cellNo=485
rlabel pdiffusion 52 -893 52 -893 0 feedthrough
rlabel pdiffusion 59 -893 59 -893 0 feedthrough
rlabel pdiffusion 66 -893 66 -893 0 feedthrough
rlabel pdiffusion 73 -893 73 -893 0 feedthrough
rlabel pdiffusion 80 -893 80 -893 0 feedthrough
rlabel pdiffusion 87 -893 87 -893 0 feedthrough
rlabel pdiffusion 94 -893 94 -893 0 feedthrough
rlabel pdiffusion 101 -893 101 -893 0 feedthrough
rlabel pdiffusion 108 -893 108 -893 0 feedthrough
rlabel pdiffusion 115 -893 115 -893 0 feedthrough
rlabel pdiffusion 122 -893 122 -893 0 feedthrough
rlabel pdiffusion 129 -893 129 -893 0 cellNo=181
rlabel pdiffusion 136 -893 136 -893 0 feedthrough
rlabel pdiffusion 143 -893 143 -893 0 feedthrough
rlabel pdiffusion 150 -893 150 -893 0 feedthrough
rlabel pdiffusion 157 -893 157 -893 0 feedthrough
rlabel pdiffusion 164 -893 164 -893 0 cellNo=412
rlabel pdiffusion 171 -893 171 -893 0 feedthrough
rlabel pdiffusion 178 -893 178 -893 0 feedthrough
rlabel pdiffusion 185 -893 185 -893 0 feedthrough
rlabel pdiffusion 192 -893 192 -893 0 feedthrough
rlabel pdiffusion 199 -893 199 -893 0 feedthrough
rlabel pdiffusion 206 -893 206 -893 0 feedthrough
rlabel pdiffusion 213 -893 213 -893 0 feedthrough
rlabel pdiffusion 220 -893 220 -893 0 feedthrough
rlabel pdiffusion 227 -893 227 -893 0 feedthrough
rlabel pdiffusion 234 -893 234 -893 0 cellNo=240
rlabel pdiffusion 241 -893 241 -893 0 feedthrough
rlabel pdiffusion 248 -893 248 -893 0 feedthrough
rlabel pdiffusion 255 -893 255 -893 0 feedthrough
rlabel pdiffusion 262 -893 262 -893 0 feedthrough
rlabel pdiffusion 269 -893 269 -893 0 feedthrough
rlabel pdiffusion 276 -893 276 -893 0 feedthrough
rlabel pdiffusion 283 -893 283 -893 0 feedthrough
rlabel pdiffusion 290 -893 290 -893 0 feedthrough
rlabel pdiffusion 297 -893 297 -893 0 feedthrough
rlabel pdiffusion 304 -893 304 -893 0 feedthrough
rlabel pdiffusion 311 -893 311 -893 0 feedthrough
rlabel pdiffusion 318 -893 318 -893 0 feedthrough
rlabel pdiffusion 325 -893 325 -893 0 feedthrough
rlabel pdiffusion 332 -893 332 -893 0 feedthrough
rlabel pdiffusion 339 -893 339 -893 0 feedthrough
rlabel pdiffusion 346 -893 346 -893 0 feedthrough
rlabel pdiffusion 353 -893 353 -893 0 feedthrough
rlabel pdiffusion 360 -893 360 -893 0 feedthrough
rlabel pdiffusion 367 -893 367 -893 0 cellNo=200
rlabel pdiffusion 374 -893 374 -893 0 feedthrough
rlabel pdiffusion 381 -893 381 -893 0 feedthrough
rlabel pdiffusion 388 -893 388 -893 0 feedthrough
rlabel pdiffusion 395 -893 395 -893 0 feedthrough
rlabel pdiffusion 402 -893 402 -893 0 feedthrough
rlabel pdiffusion 409 -893 409 -893 0 feedthrough
rlabel pdiffusion 416 -893 416 -893 0 feedthrough
rlabel pdiffusion 423 -893 423 -893 0 feedthrough
rlabel pdiffusion 430 -893 430 -893 0 feedthrough
rlabel pdiffusion 437 -893 437 -893 0 cellNo=101
rlabel pdiffusion 444 -893 444 -893 0 feedthrough
rlabel pdiffusion 451 -893 451 -893 0 feedthrough
rlabel pdiffusion 458 -893 458 -893 0 cellNo=304
rlabel pdiffusion 465 -893 465 -893 0 cellNo=551
rlabel pdiffusion 472 -893 472 -893 0 feedthrough
rlabel pdiffusion 479 -893 479 -893 0 feedthrough
rlabel pdiffusion 486 -893 486 -893 0 feedthrough
rlabel pdiffusion 493 -893 493 -893 0 feedthrough
rlabel pdiffusion 500 -893 500 -893 0 feedthrough
rlabel pdiffusion 507 -893 507 -893 0 cellNo=198
rlabel pdiffusion 514 -893 514 -893 0 feedthrough
rlabel pdiffusion 521 -893 521 -893 0 feedthrough
rlabel pdiffusion 528 -893 528 -893 0 feedthrough
rlabel pdiffusion 535 -893 535 -893 0 cellNo=10
rlabel pdiffusion 542 -893 542 -893 0 cellNo=245
rlabel pdiffusion 549 -893 549 -893 0 cellNo=225
rlabel pdiffusion 556 -893 556 -893 0 feedthrough
rlabel pdiffusion 563 -893 563 -893 0 feedthrough
rlabel pdiffusion 570 -893 570 -893 0 feedthrough
rlabel pdiffusion 577 -893 577 -893 0 feedthrough
rlabel pdiffusion 584 -893 584 -893 0 feedthrough
rlabel pdiffusion 591 -893 591 -893 0 feedthrough
rlabel pdiffusion 598 -893 598 -893 0 feedthrough
rlabel pdiffusion 605 -893 605 -893 0 feedthrough
rlabel pdiffusion 612 -893 612 -893 0 feedthrough
rlabel pdiffusion 619 -893 619 -893 0 feedthrough
rlabel pdiffusion 626 -893 626 -893 0 feedthrough
rlabel pdiffusion 633 -893 633 -893 0 feedthrough
rlabel pdiffusion 640 -893 640 -893 0 cellNo=369
rlabel pdiffusion 647 -893 647 -893 0 cellNo=128
rlabel pdiffusion 654 -893 654 -893 0 cellNo=172
rlabel pdiffusion 661 -893 661 -893 0 cellNo=64
rlabel pdiffusion 668 -893 668 -893 0 feedthrough
rlabel pdiffusion 675 -893 675 -893 0 feedthrough
rlabel pdiffusion 682 -893 682 -893 0 feedthrough
rlabel pdiffusion 689 -893 689 -893 0 cellNo=453
rlabel pdiffusion 696 -893 696 -893 0 feedthrough
rlabel pdiffusion 703 -893 703 -893 0 feedthrough
rlabel pdiffusion 710 -893 710 -893 0 cellNo=522
rlabel pdiffusion 717 -893 717 -893 0 feedthrough
rlabel pdiffusion 724 -893 724 -893 0 feedthrough
rlabel pdiffusion 731 -893 731 -893 0 feedthrough
rlabel pdiffusion 738 -893 738 -893 0 feedthrough
rlabel pdiffusion 745 -893 745 -893 0 feedthrough
rlabel pdiffusion 752 -893 752 -893 0 feedthrough
rlabel pdiffusion 759 -893 759 -893 0 feedthrough
rlabel pdiffusion 766 -893 766 -893 0 cellNo=89
rlabel pdiffusion 773 -893 773 -893 0 feedthrough
rlabel pdiffusion 780 -893 780 -893 0 feedthrough
rlabel pdiffusion 787 -893 787 -893 0 feedthrough
rlabel pdiffusion 794 -893 794 -893 0 feedthrough
rlabel pdiffusion 801 -893 801 -893 0 feedthrough
rlabel pdiffusion 808 -893 808 -893 0 cellNo=342
rlabel pdiffusion 815 -893 815 -893 0 feedthrough
rlabel pdiffusion 822 -893 822 -893 0 feedthrough
rlabel pdiffusion 829 -893 829 -893 0 feedthrough
rlabel pdiffusion 836 -893 836 -893 0 cellNo=281
rlabel pdiffusion 843 -893 843 -893 0 feedthrough
rlabel pdiffusion 850 -893 850 -893 0 feedthrough
rlabel pdiffusion 857 -893 857 -893 0 feedthrough
rlabel pdiffusion 864 -893 864 -893 0 feedthrough
rlabel pdiffusion 871 -893 871 -893 0 feedthrough
rlabel pdiffusion 878 -893 878 -893 0 feedthrough
rlabel pdiffusion 885 -893 885 -893 0 feedthrough
rlabel pdiffusion 892 -893 892 -893 0 feedthrough
rlabel pdiffusion 899 -893 899 -893 0 feedthrough
rlabel pdiffusion 906 -893 906 -893 0 feedthrough
rlabel pdiffusion 913 -893 913 -893 0 feedthrough
rlabel pdiffusion 920 -893 920 -893 0 feedthrough
rlabel pdiffusion 927 -893 927 -893 0 feedthrough
rlabel pdiffusion 934 -893 934 -893 0 feedthrough
rlabel pdiffusion 941 -893 941 -893 0 cellNo=244
rlabel pdiffusion 948 -893 948 -893 0 feedthrough
rlabel pdiffusion 955 -893 955 -893 0 feedthrough
rlabel pdiffusion 962 -893 962 -893 0 feedthrough
rlabel pdiffusion 969 -893 969 -893 0 feedthrough
rlabel pdiffusion 976 -893 976 -893 0 feedthrough
rlabel pdiffusion 983 -893 983 -893 0 feedthrough
rlabel pdiffusion 990 -893 990 -893 0 feedthrough
rlabel pdiffusion 997 -893 997 -893 0 cellNo=195
rlabel pdiffusion 1004 -893 1004 -893 0 feedthrough
rlabel pdiffusion 1011 -893 1011 -893 0 feedthrough
rlabel pdiffusion 1018 -893 1018 -893 0 feedthrough
rlabel pdiffusion 1025 -893 1025 -893 0 feedthrough
rlabel pdiffusion 1032 -893 1032 -893 0 feedthrough
rlabel pdiffusion 1039 -893 1039 -893 0 feedthrough
rlabel pdiffusion 1046 -893 1046 -893 0 feedthrough
rlabel pdiffusion 1053 -893 1053 -893 0 feedthrough
rlabel pdiffusion 1060 -893 1060 -893 0 feedthrough
rlabel pdiffusion 1067 -893 1067 -893 0 feedthrough
rlabel pdiffusion 1074 -893 1074 -893 0 feedthrough
rlabel pdiffusion 1081 -893 1081 -893 0 feedthrough
rlabel pdiffusion 1088 -893 1088 -893 0 feedthrough
rlabel pdiffusion 1095 -893 1095 -893 0 feedthrough
rlabel pdiffusion 1102 -893 1102 -893 0 feedthrough
rlabel pdiffusion 1109 -893 1109 -893 0 feedthrough
rlabel pdiffusion 1116 -893 1116 -893 0 feedthrough
rlabel pdiffusion 1123 -893 1123 -893 0 feedthrough
rlabel pdiffusion 1130 -893 1130 -893 0 feedthrough
rlabel pdiffusion 1137 -893 1137 -893 0 feedthrough
rlabel pdiffusion 1144 -893 1144 -893 0 feedthrough
rlabel pdiffusion 1151 -893 1151 -893 0 feedthrough
rlabel pdiffusion 1158 -893 1158 -893 0 feedthrough
rlabel pdiffusion 1165 -893 1165 -893 0 feedthrough
rlabel pdiffusion 1172 -893 1172 -893 0 feedthrough
rlabel pdiffusion 1179 -893 1179 -893 0 feedthrough
rlabel pdiffusion 1186 -893 1186 -893 0 feedthrough
rlabel pdiffusion 1193 -893 1193 -893 0 feedthrough
rlabel pdiffusion 1200 -893 1200 -893 0 feedthrough
rlabel pdiffusion 1207 -893 1207 -893 0 feedthrough
rlabel pdiffusion 1214 -893 1214 -893 0 feedthrough
rlabel pdiffusion 1221 -893 1221 -893 0 feedthrough
rlabel pdiffusion 1228 -893 1228 -893 0 feedthrough
rlabel pdiffusion 1235 -893 1235 -893 0 feedthrough
rlabel pdiffusion 1242 -893 1242 -893 0 feedthrough
rlabel pdiffusion 1249 -893 1249 -893 0 feedthrough
rlabel pdiffusion 1256 -893 1256 -893 0 feedthrough
rlabel pdiffusion 1263 -893 1263 -893 0 feedthrough
rlabel pdiffusion 1270 -893 1270 -893 0 feedthrough
rlabel pdiffusion 1277 -893 1277 -893 0 feedthrough
rlabel pdiffusion 1284 -893 1284 -893 0 feedthrough
rlabel pdiffusion 1291 -893 1291 -893 0 feedthrough
rlabel pdiffusion 1298 -893 1298 -893 0 feedthrough
rlabel pdiffusion 1305 -893 1305 -893 0 feedthrough
rlabel pdiffusion 1312 -893 1312 -893 0 feedthrough
rlabel pdiffusion 1319 -893 1319 -893 0 feedthrough
rlabel pdiffusion 1326 -893 1326 -893 0 feedthrough
rlabel pdiffusion 1333 -893 1333 -893 0 feedthrough
rlabel pdiffusion 1340 -893 1340 -893 0 feedthrough
rlabel pdiffusion 1347 -893 1347 -893 0 feedthrough
rlabel pdiffusion 1354 -893 1354 -893 0 feedthrough
rlabel pdiffusion 1361 -893 1361 -893 0 feedthrough
rlabel pdiffusion 1368 -893 1368 -893 0 feedthrough
rlabel pdiffusion 1375 -893 1375 -893 0 feedthrough
rlabel pdiffusion 1382 -893 1382 -893 0 feedthrough
rlabel pdiffusion 1389 -893 1389 -893 0 feedthrough
rlabel pdiffusion 1396 -893 1396 -893 0 feedthrough
rlabel pdiffusion 1403 -893 1403 -893 0 feedthrough
rlabel pdiffusion 1410 -893 1410 -893 0 feedthrough
rlabel pdiffusion 1417 -893 1417 -893 0 feedthrough
rlabel pdiffusion 1424 -893 1424 -893 0 feedthrough
rlabel pdiffusion 1431 -893 1431 -893 0 feedthrough
rlabel pdiffusion 1438 -893 1438 -893 0 feedthrough
rlabel pdiffusion 1445 -893 1445 -893 0 feedthrough
rlabel pdiffusion 1452 -893 1452 -893 0 feedthrough
rlabel pdiffusion 1459 -893 1459 -893 0 feedthrough
rlabel pdiffusion 1466 -893 1466 -893 0 feedthrough
rlabel pdiffusion 1473 -893 1473 -893 0 feedthrough
rlabel pdiffusion 1480 -893 1480 -893 0 feedthrough
rlabel pdiffusion 1487 -893 1487 -893 0 feedthrough
rlabel pdiffusion 1494 -893 1494 -893 0 feedthrough
rlabel pdiffusion 1501 -893 1501 -893 0 cellNo=72
rlabel pdiffusion 1515 -893 1515 -893 0 feedthrough
rlabel pdiffusion 3 -1010 3 -1010 0 feedthrough
rlabel pdiffusion 10 -1010 10 -1010 0 feedthrough
rlabel pdiffusion 17 -1010 17 -1010 0 feedthrough
rlabel pdiffusion 24 -1010 24 -1010 0 feedthrough
rlabel pdiffusion 31 -1010 31 -1010 0 feedthrough
rlabel pdiffusion 38 -1010 38 -1010 0 feedthrough
rlabel pdiffusion 45 -1010 45 -1010 0 feedthrough
rlabel pdiffusion 52 -1010 52 -1010 0 feedthrough
rlabel pdiffusion 59 -1010 59 -1010 0 feedthrough
rlabel pdiffusion 66 -1010 66 -1010 0 feedthrough
rlabel pdiffusion 73 -1010 73 -1010 0 feedthrough
rlabel pdiffusion 80 -1010 80 -1010 0 feedthrough
rlabel pdiffusion 87 -1010 87 -1010 0 feedthrough
rlabel pdiffusion 94 -1010 94 -1010 0 cellNo=589
rlabel pdiffusion 101 -1010 101 -1010 0 feedthrough
rlabel pdiffusion 108 -1010 108 -1010 0 feedthrough
rlabel pdiffusion 115 -1010 115 -1010 0 feedthrough
rlabel pdiffusion 122 -1010 122 -1010 0 feedthrough
rlabel pdiffusion 129 -1010 129 -1010 0 feedthrough
rlabel pdiffusion 136 -1010 136 -1010 0 feedthrough
rlabel pdiffusion 143 -1010 143 -1010 0 cellNo=243
rlabel pdiffusion 150 -1010 150 -1010 0 feedthrough
rlabel pdiffusion 157 -1010 157 -1010 0 feedthrough
rlabel pdiffusion 164 -1010 164 -1010 0 feedthrough
rlabel pdiffusion 171 -1010 171 -1010 0 feedthrough
rlabel pdiffusion 178 -1010 178 -1010 0 feedthrough
rlabel pdiffusion 185 -1010 185 -1010 0 feedthrough
rlabel pdiffusion 192 -1010 192 -1010 0 feedthrough
rlabel pdiffusion 199 -1010 199 -1010 0 feedthrough
rlabel pdiffusion 206 -1010 206 -1010 0 feedthrough
rlabel pdiffusion 213 -1010 213 -1010 0 feedthrough
rlabel pdiffusion 220 -1010 220 -1010 0 feedthrough
rlabel pdiffusion 227 -1010 227 -1010 0 feedthrough
rlabel pdiffusion 234 -1010 234 -1010 0 feedthrough
rlabel pdiffusion 241 -1010 241 -1010 0 cellNo=210
rlabel pdiffusion 248 -1010 248 -1010 0 feedthrough
rlabel pdiffusion 255 -1010 255 -1010 0 feedthrough
rlabel pdiffusion 262 -1010 262 -1010 0 feedthrough
rlabel pdiffusion 269 -1010 269 -1010 0 feedthrough
rlabel pdiffusion 276 -1010 276 -1010 0 feedthrough
rlabel pdiffusion 283 -1010 283 -1010 0 feedthrough
rlabel pdiffusion 290 -1010 290 -1010 0 feedthrough
rlabel pdiffusion 297 -1010 297 -1010 0 cellNo=15
rlabel pdiffusion 304 -1010 304 -1010 0 feedthrough
rlabel pdiffusion 311 -1010 311 -1010 0 feedthrough
rlabel pdiffusion 318 -1010 318 -1010 0 feedthrough
rlabel pdiffusion 325 -1010 325 -1010 0 feedthrough
rlabel pdiffusion 332 -1010 332 -1010 0 cellNo=253
rlabel pdiffusion 339 -1010 339 -1010 0 feedthrough
rlabel pdiffusion 346 -1010 346 -1010 0 feedthrough
rlabel pdiffusion 353 -1010 353 -1010 0 feedthrough
rlabel pdiffusion 360 -1010 360 -1010 0 feedthrough
rlabel pdiffusion 367 -1010 367 -1010 0 feedthrough
rlabel pdiffusion 374 -1010 374 -1010 0 cellNo=239
rlabel pdiffusion 381 -1010 381 -1010 0 feedthrough
rlabel pdiffusion 388 -1010 388 -1010 0 feedthrough
rlabel pdiffusion 395 -1010 395 -1010 0 feedthrough
rlabel pdiffusion 402 -1010 402 -1010 0 feedthrough
rlabel pdiffusion 409 -1010 409 -1010 0 feedthrough
rlabel pdiffusion 416 -1010 416 -1010 0 feedthrough
rlabel pdiffusion 423 -1010 423 -1010 0 feedthrough
rlabel pdiffusion 430 -1010 430 -1010 0 feedthrough
rlabel pdiffusion 437 -1010 437 -1010 0 feedthrough
rlabel pdiffusion 444 -1010 444 -1010 0 feedthrough
rlabel pdiffusion 451 -1010 451 -1010 0 feedthrough
rlabel pdiffusion 458 -1010 458 -1010 0 feedthrough
rlabel pdiffusion 465 -1010 465 -1010 0 feedthrough
rlabel pdiffusion 472 -1010 472 -1010 0 feedthrough
rlabel pdiffusion 479 -1010 479 -1010 0 cellNo=344
rlabel pdiffusion 486 -1010 486 -1010 0 feedthrough
rlabel pdiffusion 493 -1010 493 -1010 0 cellNo=504
rlabel pdiffusion 500 -1010 500 -1010 0 feedthrough
rlabel pdiffusion 507 -1010 507 -1010 0 feedthrough
rlabel pdiffusion 514 -1010 514 -1010 0 feedthrough
rlabel pdiffusion 521 -1010 521 -1010 0 feedthrough
rlabel pdiffusion 528 -1010 528 -1010 0 feedthrough
rlabel pdiffusion 535 -1010 535 -1010 0 cellNo=117
rlabel pdiffusion 542 -1010 542 -1010 0 cellNo=552
rlabel pdiffusion 549 -1010 549 -1010 0 cellNo=252
rlabel pdiffusion 556 -1010 556 -1010 0 feedthrough
rlabel pdiffusion 563 -1010 563 -1010 0 feedthrough
rlabel pdiffusion 570 -1010 570 -1010 0 feedthrough
rlabel pdiffusion 577 -1010 577 -1010 0 feedthrough
rlabel pdiffusion 584 -1010 584 -1010 0 feedthrough
rlabel pdiffusion 591 -1010 591 -1010 0 feedthrough
rlabel pdiffusion 598 -1010 598 -1010 0 cellNo=331
rlabel pdiffusion 605 -1010 605 -1010 0 feedthrough
rlabel pdiffusion 612 -1010 612 -1010 0 feedthrough
rlabel pdiffusion 619 -1010 619 -1010 0 feedthrough
rlabel pdiffusion 626 -1010 626 -1010 0 feedthrough
rlabel pdiffusion 633 -1010 633 -1010 0 feedthrough
rlabel pdiffusion 640 -1010 640 -1010 0 feedthrough
rlabel pdiffusion 647 -1010 647 -1010 0 feedthrough
rlabel pdiffusion 654 -1010 654 -1010 0 feedthrough
rlabel pdiffusion 661 -1010 661 -1010 0 feedthrough
rlabel pdiffusion 668 -1010 668 -1010 0 feedthrough
rlabel pdiffusion 675 -1010 675 -1010 0 cellNo=149
rlabel pdiffusion 682 -1010 682 -1010 0 feedthrough
rlabel pdiffusion 689 -1010 689 -1010 0 cellNo=189
rlabel pdiffusion 696 -1010 696 -1010 0 feedthrough
rlabel pdiffusion 703 -1010 703 -1010 0 cellNo=404
rlabel pdiffusion 710 -1010 710 -1010 0 feedthrough
rlabel pdiffusion 717 -1010 717 -1010 0 feedthrough
rlabel pdiffusion 724 -1010 724 -1010 0 feedthrough
rlabel pdiffusion 731 -1010 731 -1010 0 feedthrough
rlabel pdiffusion 738 -1010 738 -1010 0 feedthrough
rlabel pdiffusion 745 -1010 745 -1010 0 cellNo=91
rlabel pdiffusion 752 -1010 752 -1010 0 cellNo=562
rlabel pdiffusion 759 -1010 759 -1010 0 cellNo=402
rlabel pdiffusion 766 -1010 766 -1010 0 feedthrough
rlabel pdiffusion 773 -1010 773 -1010 0 feedthrough
rlabel pdiffusion 780 -1010 780 -1010 0 feedthrough
rlabel pdiffusion 787 -1010 787 -1010 0 feedthrough
rlabel pdiffusion 794 -1010 794 -1010 0 feedthrough
rlabel pdiffusion 801 -1010 801 -1010 0 feedthrough
rlabel pdiffusion 808 -1010 808 -1010 0 feedthrough
rlabel pdiffusion 815 -1010 815 -1010 0 feedthrough
rlabel pdiffusion 822 -1010 822 -1010 0 cellNo=259
rlabel pdiffusion 829 -1010 829 -1010 0 cellNo=307
rlabel pdiffusion 836 -1010 836 -1010 0 feedthrough
rlabel pdiffusion 843 -1010 843 -1010 0 feedthrough
rlabel pdiffusion 850 -1010 850 -1010 0 feedthrough
rlabel pdiffusion 857 -1010 857 -1010 0 cellNo=220
rlabel pdiffusion 864 -1010 864 -1010 0 feedthrough
rlabel pdiffusion 871 -1010 871 -1010 0 cellNo=373
rlabel pdiffusion 878 -1010 878 -1010 0 feedthrough
rlabel pdiffusion 885 -1010 885 -1010 0 feedthrough
rlabel pdiffusion 892 -1010 892 -1010 0 feedthrough
rlabel pdiffusion 899 -1010 899 -1010 0 feedthrough
rlabel pdiffusion 906 -1010 906 -1010 0 cellNo=292
rlabel pdiffusion 913 -1010 913 -1010 0 feedthrough
rlabel pdiffusion 920 -1010 920 -1010 0 feedthrough
rlabel pdiffusion 927 -1010 927 -1010 0 feedthrough
rlabel pdiffusion 934 -1010 934 -1010 0 feedthrough
rlabel pdiffusion 941 -1010 941 -1010 0 feedthrough
rlabel pdiffusion 948 -1010 948 -1010 0 feedthrough
rlabel pdiffusion 955 -1010 955 -1010 0 feedthrough
rlabel pdiffusion 962 -1010 962 -1010 0 feedthrough
rlabel pdiffusion 969 -1010 969 -1010 0 feedthrough
rlabel pdiffusion 976 -1010 976 -1010 0 feedthrough
rlabel pdiffusion 983 -1010 983 -1010 0 feedthrough
rlabel pdiffusion 990 -1010 990 -1010 0 cellNo=98
rlabel pdiffusion 997 -1010 997 -1010 0 feedthrough
rlabel pdiffusion 1004 -1010 1004 -1010 0 feedthrough
rlabel pdiffusion 1011 -1010 1011 -1010 0 feedthrough
rlabel pdiffusion 1018 -1010 1018 -1010 0 feedthrough
rlabel pdiffusion 1025 -1010 1025 -1010 0 feedthrough
rlabel pdiffusion 1032 -1010 1032 -1010 0 feedthrough
rlabel pdiffusion 1039 -1010 1039 -1010 0 feedthrough
rlabel pdiffusion 1046 -1010 1046 -1010 0 feedthrough
rlabel pdiffusion 1053 -1010 1053 -1010 0 feedthrough
rlabel pdiffusion 1060 -1010 1060 -1010 0 feedthrough
rlabel pdiffusion 1067 -1010 1067 -1010 0 feedthrough
rlabel pdiffusion 1074 -1010 1074 -1010 0 feedthrough
rlabel pdiffusion 1081 -1010 1081 -1010 0 feedthrough
rlabel pdiffusion 1088 -1010 1088 -1010 0 feedthrough
rlabel pdiffusion 1095 -1010 1095 -1010 0 feedthrough
rlabel pdiffusion 1102 -1010 1102 -1010 0 feedthrough
rlabel pdiffusion 1109 -1010 1109 -1010 0 feedthrough
rlabel pdiffusion 1116 -1010 1116 -1010 0 feedthrough
rlabel pdiffusion 1123 -1010 1123 -1010 0 feedthrough
rlabel pdiffusion 1130 -1010 1130 -1010 0 feedthrough
rlabel pdiffusion 1137 -1010 1137 -1010 0 feedthrough
rlabel pdiffusion 1144 -1010 1144 -1010 0 feedthrough
rlabel pdiffusion 1151 -1010 1151 -1010 0 feedthrough
rlabel pdiffusion 1158 -1010 1158 -1010 0 feedthrough
rlabel pdiffusion 1165 -1010 1165 -1010 0 feedthrough
rlabel pdiffusion 1172 -1010 1172 -1010 0 feedthrough
rlabel pdiffusion 1179 -1010 1179 -1010 0 feedthrough
rlabel pdiffusion 1186 -1010 1186 -1010 0 feedthrough
rlabel pdiffusion 1193 -1010 1193 -1010 0 feedthrough
rlabel pdiffusion 1200 -1010 1200 -1010 0 feedthrough
rlabel pdiffusion 1207 -1010 1207 -1010 0 feedthrough
rlabel pdiffusion 1214 -1010 1214 -1010 0 feedthrough
rlabel pdiffusion 1221 -1010 1221 -1010 0 feedthrough
rlabel pdiffusion 1228 -1010 1228 -1010 0 feedthrough
rlabel pdiffusion 1235 -1010 1235 -1010 0 feedthrough
rlabel pdiffusion 1242 -1010 1242 -1010 0 feedthrough
rlabel pdiffusion 1249 -1010 1249 -1010 0 feedthrough
rlabel pdiffusion 1256 -1010 1256 -1010 0 feedthrough
rlabel pdiffusion 1263 -1010 1263 -1010 0 feedthrough
rlabel pdiffusion 1270 -1010 1270 -1010 0 feedthrough
rlabel pdiffusion 1277 -1010 1277 -1010 0 feedthrough
rlabel pdiffusion 1284 -1010 1284 -1010 0 feedthrough
rlabel pdiffusion 1291 -1010 1291 -1010 0 feedthrough
rlabel pdiffusion 1298 -1010 1298 -1010 0 feedthrough
rlabel pdiffusion 1305 -1010 1305 -1010 0 feedthrough
rlabel pdiffusion 1312 -1010 1312 -1010 0 feedthrough
rlabel pdiffusion 1319 -1010 1319 -1010 0 feedthrough
rlabel pdiffusion 1326 -1010 1326 -1010 0 feedthrough
rlabel pdiffusion 1333 -1010 1333 -1010 0 feedthrough
rlabel pdiffusion 1340 -1010 1340 -1010 0 feedthrough
rlabel pdiffusion 1347 -1010 1347 -1010 0 feedthrough
rlabel pdiffusion 1354 -1010 1354 -1010 0 feedthrough
rlabel pdiffusion 1361 -1010 1361 -1010 0 feedthrough
rlabel pdiffusion 1368 -1010 1368 -1010 0 feedthrough
rlabel pdiffusion 1375 -1010 1375 -1010 0 feedthrough
rlabel pdiffusion 1382 -1010 1382 -1010 0 feedthrough
rlabel pdiffusion 1389 -1010 1389 -1010 0 feedthrough
rlabel pdiffusion 1396 -1010 1396 -1010 0 feedthrough
rlabel pdiffusion 1403 -1010 1403 -1010 0 feedthrough
rlabel pdiffusion 1410 -1010 1410 -1010 0 feedthrough
rlabel pdiffusion 1417 -1010 1417 -1010 0 feedthrough
rlabel pdiffusion 1424 -1010 1424 -1010 0 cellNo=108
rlabel pdiffusion 1431 -1010 1431 -1010 0 feedthrough
rlabel pdiffusion 1438 -1010 1438 -1010 0 feedthrough
rlabel pdiffusion 1445 -1010 1445 -1010 0 feedthrough
rlabel pdiffusion 1452 -1010 1452 -1010 0 feedthrough
rlabel pdiffusion 1459 -1010 1459 -1010 0 feedthrough
rlabel pdiffusion 3 -1157 3 -1157 0 feedthrough
rlabel pdiffusion 10 -1157 10 -1157 0 cellNo=563
rlabel pdiffusion 17 -1157 17 -1157 0 feedthrough
rlabel pdiffusion 24 -1157 24 -1157 0 feedthrough
rlabel pdiffusion 31 -1157 31 -1157 0 cellNo=50
rlabel pdiffusion 38 -1157 38 -1157 0 cellNo=432
rlabel pdiffusion 45 -1157 45 -1157 0 feedthrough
rlabel pdiffusion 52 -1157 52 -1157 0 feedthrough
rlabel pdiffusion 59 -1157 59 -1157 0 feedthrough
rlabel pdiffusion 66 -1157 66 -1157 0 feedthrough
rlabel pdiffusion 73 -1157 73 -1157 0 feedthrough
rlabel pdiffusion 80 -1157 80 -1157 0 cellNo=376
rlabel pdiffusion 87 -1157 87 -1157 0 feedthrough
rlabel pdiffusion 94 -1157 94 -1157 0 feedthrough
rlabel pdiffusion 101 -1157 101 -1157 0 feedthrough
rlabel pdiffusion 108 -1157 108 -1157 0 feedthrough
rlabel pdiffusion 115 -1157 115 -1157 0 feedthrough
rlabel pdiffusion 122 -1157 122 -1157 0 feedthrough
rlabel pdiffusion 129 -1157 129 -1157 0 feedthrough
rlabel pdiffusion 136 -1157 136 -1157 0 feedthrough
rlabel pdiffusion 143 -1157 143 -1157 0 feedthrough
rlabel pdiffusion 150 -1157 150 -1157 0 feedthrough
rlabel pdiffusion 157 -1157 157 -1157 0 feedthrough
rlabel pdiffusion 164 -1157 164 -1157 0 cellNo=320
rlabel pdiffusion 171 -1157 171 -1157 0 feedthrough
rlabel pdiffusion 178 -1157 178 -1157 0 feedthrough
rlabel pdiffusion 185 -1157 185 -1157 0 feedthrough
rlabel pdiffusion 192 -1157 192 -1157 0 feedthrough
rlabel pdiffusion 199 -1157 199 -1157 0 cellNo=285
rlabel pdiffusion 206 -1157 206 -1157 0 feedthrough
rlabel pdiffusion 213 -1157 213 -1157 0 feedthrough
rlabel pdiffusion 220 -1157 220 -1157 0 feedthrough
rlabel pdiffusion 227 -1157 227 -1157 0 feedthrough
rlabel pdiffusion 234 -1157 234 -1157 0 feedthrough
rlabel pdiffusion 241 -1157 241 -1157 0 feedthrough
rlabel pdiffusion 248 -1157 248 -1157 0 feedthrough
rlabel pdiffusion 255 -1157 255 -1157 0 feedthrough
rlabel pdiffusion 262 -1157 262 -1157 0 feedthrough
rlabel pdiffusion 269 -1157 269 -1157 0 feedthrough
rlabel pdiffusion 276 -1157 276 -1157 0 feedthrough
rlabel pdiffusion 283 -1157 283 -1157 0 feedthrough
rlabel pdiffusion 290 -1157 290 -1157 0 feedthrough
rlabel pdiffusion 297 -1157 297 -1157 0 feedthrough
rlabel pdiffusion 304 -1157 304 -1157 0 feedthrough
rlabel pdiffusion 311 -1157 311 -1157 0 feedthrough
rlabel pdiffusion 318 -1157 318 -1157 0 feedthrough
rlabel pdiffusion 325 -1157 325 -1157 0 feedthrough
rlabel pdiffusion 332 -1157 332 -1157 0 feedthrough
rlabel pdiffusion 339 -1157 339 -1157 0 feedthrough
rlabel pdiffusion 346 -1157 346 -1157 0 feedthrough
rlabel pdiffusion 353 -1157 353 -1157 0 cellNo=411
rlabel pdiffusion 360 -1157 360 -1157 0 feedthrough
rlabel pdiffusion 367 -1157 367 -1157 0 feedthrough
rlabel pdiffusion 374 -1157 374 -1157 0 feedthrough
rlabel pdiffusion 381 -1157 381 -1157 0 feedthrough
rlabel pdiffusion 388 -1157 388 -1157 0 cellNo=444
rlabel pdiffusion 395 -1157 395 -1157 0 feedthrough
rlabel pdiffusion 402 -1157 402 -1157 0 feedthrough
rlabel pdiffusion 409 -1157 409 -1157 0 feedthrough
rlabel pdiffusion 416 -1157 416 -1157 0 feedthrough
rlabel pdiffusion 423 -1157 423 -1157 0 feedthrough
rlabel pdiffusion 430 -1157 430 -1157 0 cellNo=159
rlabel pdiffusion 437 -1157 437 -1157 0 feedthrough
rlabel pdiffusion 444 -1157 444 -1157 0 cellNo=458
rlabel pdiffusion 451 -1157 451 -1157 0 feedthrough
rlabel pdiffusion 458 -1157 458 -1157 0 cellNo=596
rlabel pdiffusion 465 -1157 465 -1157 0 feedthrough
rlabel pdiffusion 472 -1157 472 -1157 0 feedthrough
rlabel pdiffusion 479 -1157 479 -1157 0 feedthrough
rlabel pdiffusion 486 -1157 486 -1157 0 feedthrough
rlabel pdiffusion 493 -1157 493 -1157 0 feedthrough
rlabel pdiffusion 500 -1157 500 -1157 0 feedthrough
rlabel pdiffusion 507 -1157 507 -1157 0 feedthrough
rlabel pdiffusion 514 -1157 514 -1157 0 feedthrough
rlabel pdiffusion 521 -1157 521 -1157 0 feedthrough
rlabel pdiffusion 528 -1157 528 -1157 0 feedthrough
rlabel pdiffusion 535 -1157 535 -1157 0 feedthrough
rlabel pdiffusion 542 -1157 542 -1157 0 feedthrough
rlabel pdiffusion 549 -1157 549 -1157 0 feedthrough
rlabel pdiffusion 556 -1157 556 -1157 0 feedthrough
rlabel pdiffusion 563 -1157 563 -1157 0 feedthrough
rlabel pdiffusion 570 -1157 570 -1157 0 feedthrough
rlabel pdiffusion 577 -1157 577 -1157 0 feedthrough
rlabel pdiffusion 584 -1157 584 -1157 0 feedthrough
rlabel pdiffusion 591 -1157 591 -1157 0 cellNo=265
rlabel pdiffusion 598 -1157 598 -1157 0 feedthrough
rlabel pdiffusion 605 -1157 605 -1157 0 cellNo=513
rlabel pdiffusion 612 -1157 612 -1157 0 feedthrough
rlabel pdiffusion 619 -1157 619 -1157 0 feedthrough
rlabel pdiffusion 626 -1157 626 -1157 0 cellNo=583
rlabel pdiffusion 633 -1157 633 -1157 0 feedthrough
rlabel pdiffusion 640 -1157 640 -1157 0 feedthrough
rlabel pdiffusion 647 -1157 647 -1157 0 feedthrough
rlabel pdiffusion 654 -1157 654 -1157 0 feedthrough
rlabel pdiffusion 661 -1157 661 -1157 0 cellNo=277
rlabel pdiffusion 668 -1157 668 -1157 0 cellNo=224
rlabel pdiffusion 675 -1157 675 -1157 0 feedthrough
rlabel pdiffusion 682 -1157 682 -1157 0 feedthrough
rlabel pdiffusion 689 -1157 689 -1157 0 feedthrough
rlabel pdiffusion 696 -1157 696 -1157 0 feedthrough
rlabel pdiffusion 703 -1157 703 -1157 0 feedthrough
rlabel pdiffusion 710 -1157 710 -1157 0 feedthrough
rlabel pdiffusion 717 -1157 717 -1157 0 cellNo=426
rlabel pdiffusion 724 -1157 724 -1157 0 feedthrough
rlabel pdiffusion 731 -1157 731 -1157 0 cellNo=39
rlabel pdiffusion 738 -1157 738 -1157 0 feedthrough
rlabel pdiffusion 745 -1157 745 -1157 0 feedthrough
rlabel pdiffusion 752 -1157 752 -1157 0 cellNo=428
rlabel pdiffusion 759 -1157 759 -1157 0 feedthrough
rlabel pdiffusion 766 -1157 766 -1157 0 feedthrough
rlabel pdiffusion 773 -1157 773 -1157 0 feedthrough
rlabel pdiffusion 780 -1157 780 -1157 0 feedthrough
rlabel pdiffusion 787 -1157 787 -1157 0 feedthrough
rlabel pdiffusion 794 -1157 794 -1157 0 cellNo=355
rlabel pdiffusion 801 -1157 801 -1157 0 feedthrough
rlabel pdiffusion 808 -1157 808 -1157 0 feedthrough
rlabel pdiffusion 815 -1157 815 -1157 0 feedthrough
rlabel pdiffusion 822 -1157 822 -1157 0 feedthrough
rlabel pdiffusion 829 -1157 829 -1157 0 cellNo=75
rlabel pdiffusion 836 -1157 836 -1157 0 feedthrough
rlabel pdiffusion 843 -1157 843 -1157 0 feedthrough
rlabel pdiffusion 850 -1157 850 -1157 0 feedthrough
rlabel pdiffusion 857 -1157 857 -1157 0 cellNo=367
rlabel pdiffusion 864 -1157 864 -1157 0 feedthrough
rlabel pdiffusion 871 -1157 871 -1157 0 feedthrough
rlabel pdiffusion 878 -1157 878 -1157 0 feedthrough
rlabel pdiffusion 885 -1157 885 -1157 0 feedthrough
rlabel pdiffusion 892 -1157 892 -1157 0 cellNo=362
rlabel pdiffusion 899 -1157 899 -1157 0 feedthrough
rlabel pdiffusion 906 -1157 906 -1157 0 feedthrough
rlabel pdiffusion 913 -1157 913 -1157 0 feedthrough
rlabel pdiffusion 920 -1157 920 -1157 0 feedthrough
rlabel pdiffusion 927 -1157 927 -1157 0 feedthrough
rlabel pdiffusion 934 -1157 934 -1157 0 cellNo=535
rlabel pdiffusion 941 -1157 941 -1157 0 feedthrough
rlabel pdiffusion 948 -1157 948 -1157 0 feedthrough
rlabel pdiffusion 955 -1157 955 -1157 0 cellNo=218
rlabel pdiffusion 962 -1157 962 -1157 0 feedthrough
rlabel pdiffusion 969 -1157 969 -1157 0 feedthrough
rlabel pdiffusion 976 -1157 976 -1157 0 feedthrough
rlabel pdiffusion 983 -1157 983 -1157 0 feedthrough
rlabel pdiffusion 990 -1157 990 -1157 0 feedthrough
rlabel pdiffusion 997 -1157 997 -1157 0 feedthrough
rlabel pdiffusion 1004 -1157 1004 -1157 0 feedthrough
rlabel pdiffusion 1011 -1157 1011 -1157 0 feedthrough
rlabel pdiffusion 1018 -1157 1018 -1157 0 feedthrough
rlabel pdiffusion 1025 -1157 1025 -1157 0 feedthrough
rlabel pdiffusion 1032 -1157 1032 -1157 0 feedthrough
rlabel pdiffusion 1039 -1157 1039 -1157 0 feedthrough
rlabel pdiffusion 1046 -1157 1046 -1157 0 feedthrough
rlabel pdiffusion 1053 -1157 1053 -1157 0 feedthrough
rlabel pdiffusion 1060 -1157 1060 -1157 0 feedthrough
rlabel pdiffusion 1067 -1157 1067 -1157 0 feedthrough
rlabel pdiffusion 1074 -1157 1074 -1157 0 feedthrough
rlabel pdiffusion 1081 -1157 1081 -1157 0 feedthrough
rlabel pdiffusion 1088 -1157 1088 -1157 0 feedthrough
rlabel pdiffusion 1095 -1157 1095 -1157 0 feedthrough
rlabel pdiffusion 1102 -1157 1102 -1157 0 feedthrough
rlabel pdiffusion 1109 -1157 1109 -1157 0 feedthrough
rlabel pdiffusion 1116 -1157 1116 -1157 0 feedthrough
rlabel pdiffusion 1123 -1157 1123 -1157 0 feedthrough
rlabel pdiffusion 1130 -1157 1130 -1157 0 feedthrough
rlabel pdiffusion 1137 -1157 1137 -1157 0 feedthrough
rlabel pdiffusion 1144 -1157 1144 -1157 0 feedthrough
rlabel pdiffusion 1151 -1157 1151 -1157 0 feedthrough
rlabel pdiffusion 1158 -1157 1158 -1157 0 feedthrough
rlabel pdiffusion 1165 -1157 1165 -1157 0 feedthrough
rlabel pdiffusion 1172 -1157 1172 -1157 0 feedthrough
rlabel pdiffusion 1179 -1157 1179 -1157 0 feedthrough
rlabel pdiffusion 1186 -1157 1186 -1157 0 feedthrough
rlabel pdiffusion 1193 -1157 1193 -1157 0 feedthrough
rlabel pdiffusion 1200 -1157 1200 -1157 0 feedthrough
rlabel pdiffusion 1207 -1157 1207 -1157 0 feedthrough
rlabel pdiffusion 1214 -1157 1214 -1157 0 feedthrough
rlabel pdiffusion 1221 -1157 1221 -1157 0 feedthrough
rlabel pdiffusion 1228 -1157 1228 -1157 0 feedthrough
rlabel pdiffusion 1235 -1157 1235 -1157 0 feedthrough
rlabel pdiffusion 1242 -1157 1242 -1157 0 feedthrough
rlabel pdiffusion 1249 -1157 1249 -1157 0 feedthrough
rlabel pdiffusion 1256 -1157 1256 -1157 0 feedthrough
rlabel pdiffusion 1263 -1157 1263 -1157 0 feedthrough
rlabel pdiffusion 1270 -1157 1270 -1157 0 feedthrough
rlabel pdiffusion 1277 -1157 1277 -1157 0 feedthrough
rlabel pdiffusion 1284 -1157 1284 -1157 0 feedthrough
rlabel pdiffusion 1291 -1157 1291 -1157 0 feedthrough
rlabel pdiffusion 1298 -1157 1298 -1157 0 feedthrough
rlabel pdiffusion 1305 -1157 1305 -1157 0 feedthrough
rlabel pdiffusion 1312 -1157 1312 -1157 0 feedthrough
rlabel pdiffusion 1319 -1157 1319 -1157 0 feedthrough
rlabel pdiffusion 1326 -1157 1326 -1157 0 feedthrough
rlabel pdiffusion 1333 -1157 1333 -1157 0 feedthrough
rlabel pdiffusion 1340 -1157 1340 -1157 0 feedthrough
rlabel pdiffusion 1347 -1157 1347 -1157 0 feedthrough
rlabel pdiffusion 1354 -1157 1354 -1157 0 feedthrough
rlabel pdiffusion 1361 -1157 1361 -1157 0 feedthrough
rlabel pdiffusion 1368 -1157 1368 -1157 0 feedthrough
rlabel pdiffusion 1375 -1157 1375 -1157 0 feedthrough
rlabel pdiffusion 1382 -1157 1382 -1157 0 feedthrough
rlabel pdiffusion 1389 -1157 1389 -1157 0 feedthrough
rlabel pdiffusion 1396 -1157 1396 -1157 0 feedthrough
rlabel pdiffusion 1403 -1157 1403 -1157 0 feedthrough
rlabel pdiffusion 1410 -1157 1410 -1157 0 feedthrough
rlabel pdiffusion 1417 -1157 1417 -1157 0 feedthrough
rlabel pdiffusion 1424 -1157 1424 -1157 0 feedthrough
rlabel pdiffusion 1431 -1157 1431 -1157 0 feedthrough
rlabel pdiffusion 1438 -1157 1438 -1157 0 feedthrough
rlabel pdiffusion 1445 -1157 1445 -1157 0 feedthrough
rlabel pdiffusion 1452 -1157 1452 -1157 0 feedthrough
rlabel pdiffusion 1459 -1157 1459 -1157 0 feedthrough
rlabel pdiffusion 1466 -1157 1466 -1157 0 feedthrough
rlabel pdiffusion 1473 -1157 1473 -1157 0 feedthrough
rlabel pdiffusion 1480 -1157 1480 -1157 0 feedthrough
rlabel pdiffusion 1487 -1157 1487 -1157 0 feedthrough
rlabel pdiffusion 1494 -1157 1494 -1157 0 feedthrough
rlabel pdiffusion 1501 -1157 1501 -1157 0 feedthrough
rlabel pdiffusion 1508 -1157 1508 -1157 0 feedthrough
rlabel pdiffusion 1515 -1157 1515 -1157 0 feedthrough
rlabel pdiffusion 1522 -1157 1522 -1157 0 feedthrough
rlabel pdiffusion 1529 -1157 1529 -1157 0 feedthrough
rlabel pdiffusion 1536 -1157 1536 -1157 0 feedthrough
rlabel pdiffusion 1543 -1157 1543 -1157 0 feedthrough
rlabel pdiffusion 1550 -1157 1550 -1157 0 feedthrough
rlabel pdiffusion 1557 -1157 1557 -1157 0 feedthrough
rlabel pdiffusion 1564 -1157 1564 -1157 0 feedthrough
rlabel pdiffusion 1571 -1157 1571 -1157 0 feedthrough
rlabel pdiffusion 1578 -1157 1578 -1157 0 feedthrough
rlabel pdiffusion 1585 -1157 1585 -1157 0 feedthrough
rlabel pdiffusion 1592 -1157 1592 -1157 0 feedthrough
rlabel pdiffusion 1599 -1157 1599 -1157 0 feedthrough
rlabel pdiffusion 3 -1282 3 -1282 0 feedthrough
rlabel pdiffusion 10 -1282 10 -1282 0 feedthrough
rlabel pdiffusion 17 -1282 17 -1282 0 feedthrough
rlabel pdiffusion 24 -1282 24 -1282 0 feedthrough
rlabel pdiffusion 31 -1282 31 -1282 0 feedthrough
rlabel pdiffusion 38 -1282 38 -1282 0 feedthrough
rlabel pdiffusion 45 -1282 45 -1282 0 feedthrough
rlabel pdiffusion 52 -1282 52 -1282 0 feedthrough
rlabel pdiffusion 59 -1282 59 -1282 0 cellNo=71
rlabel pdiffusion 66 -1282 66 -1282 0 feedthrough
rlabel pdiffusion 73 -1282 73 -1282 0 feedthrough
rlabel pdiffusion 80 -1282 80 -1282 0 feedthrough
rlabel pdiffusion 87 -1282 87 -1282 0 feedthrough
rlabel pdiffusion 94 -1282 94 -1282 0 feedthrough
rlabel pdiffusion 101 -1282 101 -1282 0 cellNo=23
rlabel pdiffusion 108 -1282 108 -1282 0 feedthrough
rlabel pdiffusion 115 -1282 115 -1282 0 feedthrough
rlabel pdiffusion 122 -1282 122 -1282 0 feedthrough
rlabel pdiffusion 129 -1282 129 -1282 0 cellNo=171
rlabel pdiffusion 136 -1282 136 -1282 0 feedthrough
rlabel pdiffusion 143 -1282 143 -1282 0 feedthrough
rlabel pdiffusion 150 -1282 150 -1282 0 feedthrough
rlabel pdiffusion 157 -1282 157 -1282 0 feedthrough
rlabel pdiffusion 164 -1282 164 -1282 0 feedthrough
rlabel pdiffusion 171 -1282 171 -1282 0 cellNo=460
rlabel pdiffusion 178 -1282 178 -1282 0 feedthrough
rlabel pdiffusion 185 -1282 185 -1282 0 feedthrough
rlabel pdiffusion 192 -1282 192 -1282 0 feedthrough
rlabel pdiffusion 199 -1282 199 -1282 0 feedthrough
rlabel pdiffusion 206 -1282 206 -1282 0 feedthrough
rlabel pdiffusion 213 -1282 213 -1282 0 feedthrough
rlabel pdiffusion 220 -1282 220 -1282 0 feedthrough
rlabel pdiffusion 227 -1282 227 -1282 0 feedthrough
rlabel pdiffusion 234 -1282 234 -1282 0 feedthrough
rlabel pdiffusion 241 -1282 241 -1282 0 feedthrough
rlabel pdiffusion 248 -1282 248 -1282 0 feedthrough
rlabel pdiffusion 255 -1282 255 -1282 0 feedthrough
rlabel pdiffusion 262 -1282 262 -1282 0 feedthrough
rlabel pdiffusion 269 -1282 269 -1282 0 feedthrough
rlabel pdiffusion 276 -1282 276 -1282 0 feedthrough
rlabel pdiffusion 283 -1282 283 -1282 0 feedthrough
rlabel pdiffusion 290 -1282 290 -1282 0 feedthrough
rlabel pdiffusion 297 -1282 297 -1282 0 feedthrough
rlabel pdiffusion 304 -1282 304 -1282 0 feedthrough
rlabel pdiffusion 311 -1282 311 -1282 0 feedthrough
rlabel pdiffusion 318 -1282 318 -1282 0 cellNo=273
rlabel pdiffusion 325 -1282 325 -1282 0 feedthrough
rlabel pdiffusion 332 -1282 332 -1282 0 feedthrough
rlabel pdiffusion 339 -1282 339 -1282 0 cellNo=62
rlabel pdiffusion 346 -1282 346 -1282 0 feedthrough
rlabel pdiffusion 353 -1282 353 -1282 0 feedthrough
rlabel pdiffusion 360 -1282 360 -1282 0 cellNo=152
rlabel pdiffusion 367 -1282 367 -1282 0 feedthrough
rlabel pdiffusion 374 -1282 374 -1282 0 feedthrough
rlabel pdiffusion 381 -1282 381 -1282 0 feedthrough
rlabel pdiffusion 388 -1282 388 -1282 0 feedthrough
rlabel pdiffusion 395 -1282 395 -1282 0 feedthrough
rlabel pdiffusion 402 -1282 402 -1282 0 feedthrough
rlabel pdiffusion 409 -1282 409 -1282 0 feedthrough
rlabel pdiffusion 416 -1282 416 -1282 0 feedthrough
rlabel pdiffusion 423 -1282 423 -1282 0 feedthrough
rlabel pdiffusion 430 -1282 430 -1282 0 feedthrough
rlabel pdiffusion 437 -1282 437 -1282 0 feedthrough
rlabel pdiffusion 444 -1282 444 -1282 0 feedthrough
rlabel pdiffusion 451 -1282 451 -1282 0 feedthrough
rlabel pdiffusion 458 -1282 458 -1282 0 feedthrough
rlabel pdiffusion 465 -1282 465 -1282 0 feedthrough
rlabel pdiffusion 472 -1282 472 -1282 0 feedthrough
rlabel pdiffusion 479 -1282 479 -1282 0 cellNo=389
rlabel pdiffusion 486 -1282 486 -1282 0 feedthrough
rlabel pdiffusion 493 -1282 493 -1282 0 feedthrough
rlabel pdiffusion 500 -1282 500 -1282 0 feedthrough
rlabel pdiffusion 507 -1282 507 -1282 0 cellNo=162
rlabel pdiffusion 514 -1282 514 -1282 0 feedthrough
rlabel pdiffusion 521 -1282 521 -1282 0 cellNo=332
rlabel pdiffusion 528 -1282 528 -1282 0 cellNo=187
rlabel pdiffusion 535 -1282 535 -1282 0 feedthrough
rlabel pdiffusion 542 -1282 542 -1282 0 feedthrough
rlabel pdiffusion 549 -1282 549 -1282 0 cellNo=111
rlabel pdiffusion 556 -1282 556 -1282 0 cellNo=231
rlabel pdiffusion 563 -1282 563 -1282 0 feedthrough
rlabel pdiffusion 570 -1282 570 -1282 0 feedthrough
rlabel pdiffusion 577 -1282 577 -1282 0 feedthrough
rlabel pdiffusion 584 -1282 584 -1282 0 feedthrough
rlabel pdiffusion 591 -1282 591 -1282 0 feedthrough
rlabel pdiffusion 598 -1282 598 -1282 0 feedthrough
rlabel pdiffusion 605 -1282 605 -1282 0 cellNo=223
rlabel pdiffusion 612 -1282 612 -1282 0 feedthrough
rlabel pdiffusion 619 -1282 619 -1282 0 feedthrough
rlabel pdiffusion 626 -1282 626 -1282 0 feedthrough
rlabel pdiffusion 633 -1282 633 -1282 0 feedthrough
rlabel pdiffusion 640 -1282 640 -1282 0 feedthrough
rlabel pdiffusion 647 -1282 647 -1282 0 feedthrough
rlabel pdiffusion 654 -1282 654 -1282 0 feedthrough
rlabel pdiffusion 661 -1282 661 -1282 0 feedthrough
rlabel pdiffusion 668 -1282 668 -1282 0 feedthrough
rlabel pdiffusion 675 -1282 675 -1282 0 feedthrough
rlabel pdiffusion 682 -1282 682 -1282 0 feedthrough
rlabel pdiffusion 689 -1282 689 -1282 0 feedthrough
rlabel pdiffusion 696 -1282 696 -1282 0 feedthrough
rlabel pdiffusion 703 -1282 703 -1282 0 feedthrough
rlabel pdiffusion 710 -1282 710 -1282 0 feedthrough
rlabel pdiffusion 717 -1282 717 -1282 0 cellNo=380
rlabel pdiffusion 724 -1282 724 -1282 0 cellNo=323
rlabel pdiffusion 731 -1282 731 -1282 0 feedthrough
rlabel pdiffusion 738 -1282 738 -1282 0 feedthrough
rlabel pdiffusion 745 -1282 745 -1282 0 feedthrough
rlabel pdiffusion 752 -1282 752 -1282 0 cellNo=183
rlabel pdiffusion 759 -1282 759 -1282 0 feedthrough
rlabel pdiffusion 766 -1282 766 -1282 0 cellNo=365
rlabel pdiffusion 773 -1282 773 -1282 0 feedthrough
rlabel pdiffusion 780 -1282 780 -1282 0 cellNo=395
rlabel pdiffusion 787 -1282 787 -1282 0 feedthrough
rlabel pdiffusion 794 -1282 794 -1282 0 feedthrough
rlabel pdiffusion 801 -1282 801 -1282 0 feedthrough
rlabel pdiffusion 808 -1282 808 -1282 0 feedthrough
rlabel pdiffusion 815 -1282 815 -1282 0 feedthrough
rlabel pdiffusion 822 -1282 822 -1282 0 feedthrough
rlabel pdiffusion 829 -1282 829 -1282 0 feedthrough
rlabel pdiffusion 836 -1282 836 -1282 0 cellNo=21
rlabel pdiffusion 843 -1282 843 -1282 0 feedthrough
rlabel pdiffusion 850 -1282 850 -1282 0 feedthrough
rlabel pdiffusion 857 -1282 857 -1282 0 cellNo=473
rlabel pdiffusion 864 -1282 864 -1282 0 feedthrough
rlabel pdiffusion 871 -1282 871 -1282 0 feedthrough
rlabel pdiffusion 878 -1282 878 -1282 0 feedthrough
rlabel pdiffusion 885 -1282 885 -1282 0 feedthrough
rlabel pdiffusion 892 -1282 892 -1282 0 feedthrough
rlabel pdiffusion 899 -1282 899 -1282 0 feedthrough
rlabel pdiffusion 906 -1282 906 -1282 0 feedthrough
rlabel pdiffusion 913 -1282 913 -1282 0 feedthrough
rlabel pdiffusion 920 -1282 920 -1282 0 cellNo=73
rlabel pdiffusion 927 -1282 927 -1282 0 feedthrough
rlabel pdiffusion 934 -1282 934 -1282 0 cellNo=530
rlabel pdiffusion 941 -1282 941 -1282 0 feedthrough
rlabel pdiffusion 948 -1282 948 -1282 0 feedthrough
rlabel pdiffusion 955 -1282 955 -1282 0 feedthrough
rlabel pdiffusion 962 -1282 962 -1282 0 feedthrough
rlabel pdiffusion 969 -1282 969 -1282 0 feedthrough
rlabel pdiffusion 976 -1282 976 -1282 0 feedthrough
rlabel pdiffusion 983 -1282 983 -1282 0 feedthrough
rlabel pdiffusion 990 -1282 990 -1282 0 feedthrough
rlabel pdiffusion 997 -1282 997 -1282 0 feedthrough
rlabel pdiffusion 1004 -1282 1004 -1282 0 feedthrough
rlabel pdiffusion 1011 -1282 1011 -1282 0 feedthrough
rlabel pdiffusion 1018 -1282 1018 -1282 0 feedthrough
rlabel pdiffusion 1025 -1282 1025 -1282 0 feedthrough
rlabel pdiffusion 1032 -1282 1032 -1282 0 feedthrough
rlabel pdiffusion 1039 -1282 1039 -1282 0 feedthrough
rlabel pdiffusion 1046 -1282 1046 -1282 0 feedthrough
rlabel pdiffusion 1053 -1282 1053 -1282 0 cellNo=205
rlabel pdiffusion 1060 -1282 1060 -1282 0 feedthrough
rlabel pdiffusion 1067 -1282 1067 -1282 0 feedthrough
rlabel pdiffusion 1074 -1282 1074 -1282 0 feedthrough
rlabel pdiffusion 1081 -1282 1081 -1282 0 feedthrough
rlabel pdiffusion 1088 -1282 1088 -1282 0 feedthrough
rlabel pdiffusion 1095 -1282 1095 -1282 0 feedthrough
rlabel pdiffusion 1102 -1282 1102 -1282 0 feedthrough
rlabel pdiffusion 1109 -1282 1109 -1282 0 feedthrough
rlabel pdiffusion 1116 -1282 1116 -1282 0 feedthrough
rlabel pdiffusion 1123 -1282 1123 -1282 0 feedthrough
rlabel pdiffusion 1130 -1282 1130 -1282 0 feedthrough
rlabel pdiffusion 1137 -1282 1137 -1282 0 feedthrough
rlabel pdiffusion 1144 -1282 1144 -1282 0 feedthrough
rlabel pdiffusion 1151 -1282 1151 -1282 0 feedthrough
rlabel pdiffusion 1158 -1282 1158 -1282 0 feedthrough
rlabel pdiffusion 1165 -1282 1165 -1282 0 feedthrough
rlabel pdiffusion 1172 -1282 1172 -1282 0 cellNo=538
rlabel pdiffusion 1179 -1282 1179 -1282 0 feedthrough
rlabel pdiffusion 1186 -1282 1186 -1282 0 feedthrough
rlabel pdiffusion 1193 -1282 1193 -1282 0 feedthrough
rlabel pdiffusion 1200 -1282 1200 -1282 0 feedthrough
rlabel pdiffusion 1207 -1282 1207 -1282 0 feedthrough
rlabel pdiffusion 1214 -1282 1214 -1282 0 feedthrough
rlabel pdiffusion 1221 -1282 1221 -1282 0 feedthrough
rlabel pdiffusion 1228 -1282 1228 -1282 0 feedthrough
rlabel pdiffusion 1235 -1282 1235 -1282 0 feedthrough
rlabel pdiffusion 1242 -1282 1242 -1282 0 feedthrough
rlabel pdiffusion 1249 -1282 1249 -1282 0 feedthrough
rlabel pdiffusion 1256 -1282 1256 -1282 0 feedthrough
rlabel pdiffusion 1263 -1282 1263 -1282 0 feedthrough
rlabel pdiffusion 1270 -1282 1270 -1282 0 feedthrough
rlabel pdiffusion 1277 -1282 1277 -1282 0 feedthrough
rlabel pdiffusion 1284 -1282 1284 -1282 0 feedthrough
rlabel pdiffusion 1291 -1282 1291 -1282 0 feedthrough
rlabel pdiffusion 1298 -1282 1298 -1282 0 feedthrough
rlabel pdiffusion 1305 -1282 1305 -1282 0 feedthrough
rlabel pdiffusion 1312 -1282 1312 -1282 0 feedthrough
rlabel pdiffusion 1319 -1282 1319 -1282 0 feedthrough
rlabel pdiffusion 1326 -1282 1326 -1282 0 feedthrough
rlabel pdiffusion 1333 -1282 1333 -1282 0 feedthrough
rlabel pdiffusion 1340 -1282 1340 -1282 0 feedthrough
rlabel pdiffusion 1347 -1282 1347 -1282 0 feedthrough
rlabel pdiffusion 1354 -1282 1354 -1282 0 feedthrough
rlabel pdiffusion 1361 -1282 1361 -1282 0 feedthrough
rlabel pdiffusion 1368 -1282 1368 -1282 0 feedthrough
rlabel pdiffusion 1375 -1282 1375 -1282 0 feedthrough
rlabel pdiffusion 1382 -1282 1382 -1282 0 feedthrough
rlabel pdiffusion 1389 -1282 1389 -1282 0 feedthrough
rlabel pdiffusion 1396 -1282 1396 -1282 0 feedthrough
rlabel pdiffusion 1403 -1282 1403 -1282 0 feedthrough
rlabel pdiffusion 1410 -1282 1410 -1282 0 feedthrough
rlabel pdiffusion 1417 -1282 1417 -1282 0 feedthrough
rlabel pdiffusion 1424 -1282 1424 -1282 0 feedthrough
rlabel pdiffusion 1431 -1282 1431 -1282 0 feedthrough
rlabel pdiffusion 1438 -1282 1438 -1282 0 feedthrough
rlabel pdiffusion 1445 -1282 1445 -1282 0 feedthrough
rlabel pdiffusion 1452 -1282 1452 -1282 0 feedthrough
rlabel pdiffusion 1459 -1282 1459 -1282 0 feedthrough
rlabel pdiffusion 1466 -1282 1466 -1282 0 feedthrough
rlabel pdiffusion 1473 -1282 1473 -1282 0 feedthrough
rlabel pdiffusion 1480 -1282 1480 -1282 0 feedthrough
rlabel pdiffusion 1487 -1282 1487 -1282 0 feedthrough
rlabel pdiffusion 1494 -1282 1494 -1282 0 feedthrough
rlabel pdiffusion 1501 -1282 1501 -1282 0 feedthrough
rlabel pdiffusion 1508 -1282 1508 -1282 0 feedthrough
rlabel pdiffusion 1515 -1282 1515 -1282 0 feedthrough
rlabel pdiffusion 1522 -1282 1522 -1282 0 feedthrough
rlabel pdiffusion 1529 -1282 1529 -1282 0 feedthrough
rlabel pdiffusion 1536 -1282 1536 -1282 0 feedthrough
rlabel pdiffusion 1543 -1282 1543 -1282 0 feedthrough
rlabel pdiffusion 1550 -1282 1550 -1282 0 feedthrough
rlabel pdiffusion 1557 -1282 1557 -1282 0 feedthrough
rlabel pdiffusion 1564 -1282 1564 -1282 0 feedthrough
rlabel pdiffusion 3 -1401 3 -1401 0 feedthrough
rlabel pdiffusion 10 -1401 10 -1401 0 feedthrough
rlabel pdiffusion 17 -1401 17 -1401 0 feedthrough
rlabel pdiffusion 24 -1401 24 -1401 0 feedthrough
rlabel pdiffusion 31 -1401 31 -1401 0 feedthrough
rlabel pdiffusion 38 -1401 38 -1401 0 feedthrough
rlabel pdiffusion 45 -1401 45 -1401 0 feedthrough
rlabel pdiffusion 52 -1401 52 -1401 0 feedthrough
rlabel pdiffusion 59 -1401 59 -1401 0 feedthrough
rlabel pdiffusion 66 -1401 66 -1401 0 cellNo=387
rlabel pdiffusion 73 -1401 73 -1401 0 feedthrough
rlabel pdiffusion 80 -1401 80 -1401 0 cellNo=484
rlabel pdiffusion 87 -1401 87 -1401 0 feedthrough
rlabel pdiffusion 94 -1401 94 -1401 0 feedthrough
rlabel pdiffusion 101 -1401 101 -1401 0 feedthrough
rlabel pdiffusion 108 -1401 108 -1401 0 cellNo=173
rlabel pdiffusion 115 -1401 115 -1401 0 feedthrough
rlabel pdiffusion 122 -1401 122 -1401 0 feedthrough
rlabel pdiffusion 129 -1401 129 -1401 0 feedthrough
rlabel pdiffusion 136 -1401 136 -1401 0 feedthrough
rlabel pdiffusion 143 -1401 143 -1401 0 feedthrough
rlabel pdiffusion 150 -1401 150 -1401 0 feedthrough
rlabel pdiffusion 157 -1401 157 -1401 0 feedthrough
rlabel pdiffusion 164 -1401 164 -1401 0 feedthrough
rlabel pdiffusion 171 -1401 171 -1401 0 feedthrough
rlabel pdiffusion 178 -1401 178 -1401 0 feedthrough
rlabel pdiffusion 185 -1401 185 -1401 0 feedthrough
rlabel pdiffusion 192 -1401 192 -1401 0 feedthrough
rlabel pdiffusion 199 -1401 199 -1401 0 feedthrough
rlabel pdiffusion 206 -1401 206 -1401 0 feedthrough
rlabel pdiffusion 213 -1401 213 -1401 0 cellNo=514
rlabel pdiffusion 220 -1401 220 -1401 0 feedthrough
rlabel pdiffusion 227 -1401 227 -1401 0 feedthrough
rlabel pdiffusion 234 -1401 234 -1401 0 feedthrough
rlabel pdiffusion 241 -1401 241 -1401 0 feedthrough
rlabel pdiffusion 248 -1401 248 -1401 0 feedthrough
rlabel pdiffusion 255 -1401 255 -1401 0 feedthrough
rlabel pdiffusion 262 -1401 262 -1401 0 feedthrough
rlabel pdiffusion 269 -1401 269 -1401 0 feedthrough
rlabel pdiffusion 276 -1401 276 -1401 0 feedthrough
rlabel pdiffusion 283 -1401 283 -1401 0 feedthrough
rlabel pdiffusion 290 -1401 290 -1401 0 feedthrough
rlabel pdiffusion 297 -1401 297 -1401 0 feedthrough
rlabel pdiffusion 304 -1401 304 -1401 0 feedthrough
rlabel pdiffusion 311 -1401 311 -1401 0 feedthrough
rlabel pdiffusion 318 -1401 318 -1401 0 cellNo=188
rlabel pdiffusion 325 -1401 325 -1401 0 feedthrough
rlabel pdiffusion 332 -1401 332 -1401 0 feedthrough
rlabel pdiffusion 339 -1401 339 -1401 0 feedthrough
rlabel pdiffusion 346 -1401 346 -1401 0 feedthrough
rlabel pdiffusion 353 -1401 353 -1401 0 feedthrough
rlabel pdiffusion 360 -1401 360 -1401 0 feedthrough
rlabel pdiffusion 367 -1401 367 -1401 0 feedthrough
rlabel pdiffusion 374 -1401 374 -1401 0 feedthrough
rlabel pdiffusion 381 -1401 381 -1401 0 feedthrough
rlabel pdiffusion 388 -1401 388 -1401 0 cellNo=467
rlabel pdiffusion 395 -1401 395 -1401 0 feedthrough
rlabel pdiffusion 402 -1401 402 -1401 0 cellNo=167
rlabel pdiffusion 409 -1401 409 -1401 0 feedthrough
rlabel pdiffusion 416 -1401 416 -1401 0 cellNo=209
rlabel pdiffusion 423 -1401 423 -1401 0 feedthrough
rlabel pdiffusion 430 -1401 430 -1401 0 feedthrough
rlabel pdiffusion 437 -1401 437 -1401 0 feedthrough
rlabel pdiffusion 444 -1401 444 -1401 0 feedthrough
rlabel pdiffusion 451 -1401 451 -1401 0 feedthrough
rlabel pdiffusion 458 -1401 458 -1401 0 feedthrough
rlabel pdiffusion 465 -1401 465 -1401 0 cellNo=3
rlabel pdiffusion 472 -1401 472 -1401 0 feedthrough
rlabel pdiffusion 479 -1401 479 -1401 0 cellNo=204
rlabel pdiffusion 486 -1401 486 -1401 0 cellNo=193
rlabel pdiffusion 493 -1401 493 -1401 0 cellNo=203
rlabel pdiffusion 500 -1401 500 -1401 0 feedthrough
rlabel pdiffusion 507 -1401 507 -1401 0 feedthrough
rlabel pdiffusion 514 -1401 514 -1401 0 cellNo=37
rlabel pdiffusion 521 -1401 521 -1401 0 cellNo=454
rlabel pdiffusion 528 -1401 528 -1401 0 feedthrough
rlabel pdiffusion 535 -1401 535 -1401 0 feedthrough
rlabel pdiffusion 542 -1401 542 -1401 0 feedthrough
rlabel pdiffusion 549 -1401 549 -1401 0 feedthrough
rlabel pdiffusion 556 -1401 556 -1401 0 feedthrough
rlabel pdiffusion 563 -1401 563 -1401 0 feedthrough
rlabel pdiffusion 570 -1401 570 -1401 0 feedthrough
rlabel pdiffusion 577 -1401 577 -1401 0 feedthrough
rlabel pdiffusion 584 -1401 584 -1401 0 feedthrough
rlabel pdiffusion 591 -1401 591 -1401 0 feedthrough
rlabel pdiffusion 598 -1401 598 -1401 0 feedthrough
rlabel pdiffusion 605 -1401 605 -1401 0 feedthrough
rlabel pdiffusion 612 -1401 612 -1401 0 feedthrough
rlabel pdiffusion 619 -1401 619 -1401 0 feedthrough
rlabel pdiffusion 626 -1401 626 -1401 0 feedthrough
rlabel pdiffusion 633 -1401 633 -1401 0 feedthrough
rlabel pdiffusion 640 -1401 640 -1401 0 feedthrough
rlabel pdiffusion 647 -1401 647 -1401 0 cellNo=106
rlabel pdiffusion 654 -1401 654 -1401 0 feedthrough
rlabel pdiffusion 661 -1401 661 -1401 0 feedthrough
rlabel pdiffusion 668 -1401 668 -1401 0 feedthrough
rlabel pdiffusion 675 -1401 675 -1401 0 feedthrough
rlabel pdiffusion 682 -1401 682 -1401 0 feedthrough
rlabel pdiffusion 689 -1401 689 -1401 0 feedthrough
rlabel pdiffusion 696 -1401 696 -1401 0 feedthrough
rlabel pdiffusion 703 -1401 703 -1401 0 feedthrough
rlabel pdiffusion 710 -1401 710 -1401 0 cellNo=43
rlabel pdiffusion 717 -1401 717 -1401 0 feedthrough
rlabel pdiffusion 724 -1401 724 -1401 0 feedthrough
rlabel pdiffusion 731 -1401 731 -1401 0 feedthrough
rlabel pdiffusion 738 -1401 738 -1401 0 feedthrough
rlabel pdiffusion 745 -1401 745 -1401 0 feedthrough
rlabel pdiffusion 752 -1401 752 -1401 0 feedthrough
rlabel pdiffusion 759 -1401 759 -1401 0 feedthrough
rlabel pdiffusion 766 -1401 766 -1401 0 feedthrough
rlabel pdiffusion 773 -1401 773 -1401 0 feedthrough
rlabel pdiffusion 780 -1401 780 -1401 0 feedthrough
rlabel pdiffusion 787 -1401 787 -1401 0 feedthrough
rlabel pdiffusion 794 -1401 794 -1401 0 feedthrough
rlabel pdiffusion 801 -1401 801 -1401 0 feedthrough
rlabel pdiffusion 808 -1401 808 -1401 0 feedthrough
rlabel pdiffusion 815 -1401 815 -1401 0 feedthrough
rlabel pdiffusion 822 -1401 822 -1401 0 feedthrough
rlabel pdiffusion 829 -1401 829 -1401 0 feedthrough
rlabel pdiffusion 836 -1401 836 -1401 0 feedthrough
rlabel pdiffusion 843 -1401 843 -1401 0 cellNo=76
rlabel pdiffusion 850 -1401 850 -1401 0 feedthrough
rlabel pdiffusion 857 -1401 857 -1401 0 feedthrough
rlabel pdiffusion 864 -1401 864 -1401 0 feedthrough
rlabel pdiffusion 871 -1401 871 -1401 0 cellNo=197
rlabel pdiffusion 878 -1401 878 -1401 0 cellNo=33
rlabel pdiffusion 885 -1401 885 -1401 0 feedthrough
rlabel pdiffusion 892 -1401 892 -1401 0 feedthrough
rlabel pdiffusion 899 -1401 899 -1401 0 feedthrough
rlabel pdiffusion 906 -1401 906 -1401 0 feedthrough
rlabel pdiffusion 913 -1401 913 -1401 0 feedthrough
rlabel pdiffusion 920 -1401 920 -1401 0 cellNo=301
rlabel pdiffusion 927 -1401 927 -1401 0 feedthrough
rlabel pdiffusion 934 -1401 934 -1401 0 feedthrough
rlabel pdiffusion 941 -1401 941 -1401 0 feedthrough
rlabel pdiffusion 948 -1401 948 -1401 0 cellNo=381
rlabel pdiffusion 955 -1401 955 -1401 0 feedthrough
rlabel pdiffusion 962 -1401 962 -1401 0 feedthrough
rlabel pdiffusion 969 -1401 969 -1401 0 feedthrough
rlabel pdiffusion 976 -1401 976 -1401 0 cellNo=275
rlabel pdiffusion 983 -1401 983 -1401 0 feedthrough
rlabel pdiffusion 990 -1401 990 -1401 0 feedthrough
rlabel pdiffusion 997 -1401 997 -1401 0 feedthrough
rlabel pdiffusion 1004 -1401 1004 -1401 0 cellNo=221
rlabel pdiffusion 1011 -1401 1011 -1401 0 feedthrough
rlabel pdiffusion 1018 -1401 1018 -1401 0 cellNo=235
rlabel pdiffusion 1025 -1401 1025 -1401 0 feedthrough
rlabel pdiffusion 1032 -1401 1032 -1401 0 feedthrough
rlabel pdiffusion 1039 -1401 1039 -1401 0 feedthrough
rlabel pdiffusion 1046 -1401 1046 -1401 0 feedthrough
rlabel pdiffusion 1053 -1401 1053 -1401 0 feedthrough
rlabel pdiffusion 1060 -1401 1060 -1401 0 feedthrough
rlabel pdiffusion 1067 -1401 1067 -1401 0 feedthrough
rlabel pdiffusion 1074 -1401 1074 -1401 0 feedthrough
rlabel pdiffusion 1081 -1401 1081 -1401 0 feedthrough
rlabel pdiffusion 1088 -1401 1088 -1401 0 feedthrough
rlabel pdiffusion 1095 -1401 1095 -1401 0 feedthrough
rlabel pdiffusion 1102 -1401 1102 -1401 0 feedthrough
rlabel pdiffusion 1109 -1401 1109 -1401 0 feedthrough
rlabel pdiffusion 1116 -1401 1116 -1401 0 feedthrough
rlabel pdiffusion 1123 -1401 1123 -1401 0 feedthrough
rlabel pdiffusion 1130 -1401 1130 -1401 0 feedthrough
rlabel pdiffusion 1137 -1401 1137 -1401 0 feedthrough
rlabel pdiffusion 1144 -1401 1144 -1401 0 feedthrough
rlabel pdiffusion 1151 -1401 1151 -1401 0 feedthrough
rlabel pdiffusion 1158 -1401 1158 -1401 0 feedthrough
rlabel pdiffusion 1165 -1401 1165 -1401 0 feedthrough
rlabel pdiffusion 1172 -1401 1172 -1401 0 feedthrough
rlabel pdiffusion 1179 -1401 1179 -1401 0 feedthrough
rlabel pdiffusion 1186 -1401 1186 -1401 0 feedthrough
rlabel pdiffusion 1193 -1401 1193 -1401 0 feedthrough
rlabel pdiffusion 1200 -1401 1200 -1401 0 feedthrough
rlabel pdiffusion 1207 -1401 1207 -1401 0 feedthrough
rlabel pdiffusion 1214 -1401 1214 -1401 0 feedthrough
rlabel pdiffusion 1221 -1401 1221 -1401 0 feedthrough
rlabel pdiffusion 1228 -1401 1228 -1401 0 feedthrough
rlabel pdiffusion 1235 -1401 1235 -1401 0 feedthrough
rlabel pdiffusion 1242 -1401 1242 -1401 0 feedthrough
rlabel pdiffusion 1249 -1401 1249 -1401 0 feedthrough
rlabel pdiffusion 1256 -1401 1256 -1401 0 feedthrough
rlabel pdiffusion 1263 -1401 1263 -1401 0 feedthrough
rlabel pdiffusion 1270 -1401 1270 -1401 0 feedthrough
rlabel pdiffusion 1277 -1401 1277 -1401 0 feedthrough
rlabel pdiffusion 1284 -1401 1284 -1401 0 feedthrough
rlabel pdiffusion 1291 -1401 1291 -1401 0 feedthrough
rlabel pdiffusion 1298 -1401 1298 -1401 0 feedthrough
rlabel pdiffusion 1305 -1401 1305 -1401 0 feedthrough
rlabel pdiffusion 1312 -1401 1312 -1401 0 feedthrough
rlabel pdiffusion 1319 -1401 1319 -1401 0 feedthrough
rlabel pdiffusion 1326 -1401 1326 -1401 0 feedthrough
rlabel pdiffusion 1333 -1401 1333 -1401 0 feedthrough
rlabel pdiffusion 1340 -1401 1340 -1401 0 feedthrough
rlabel pdiffusion 1347 -1401 1347 -1401 0 feedthrough
rlabel pdiffusion 1354 -1401 1354 -1401 0 feedthrough
rlabel pdiffusion 1361 -1401 1361 -1401 0 feedthrough
rlabel pdiffusion 1368 -1401 1368 -1401 0 feedthrough
rlabel pdiffusion 1375 -1401 1375 -1401 0 feedthrough
rlabel pdiffusion 1382 -1401 1382 -1401 0 feedthrough
rlabel pdiffusion 1389 -1401 1389 -1401 0 feedthrough
rlabel pdiffusion 1396 -1401 1396 -1401 0 feedthrough
rlabel pdiffusion 1403 -1401 1403 -1401 0 feedthrough
rlabel pdiffusion 1410 -1401 1410 -1401 0 feedthrough
rlabel pdiffusion 1417 -1401 1417 -1401 0 feedthrough
rlabel pdiffusion 1424 -1401 1424 -1401 0 feedthrough
rlabel pdiffusion 1431 -1401 1431 -1401 0 feedthrough
rlabel pdiffusion 1438 -1401 1438 -1401 0 feedthrough
rlabel pdiffusion 1445 -1401 1445 -1401 0 feedthrough
rlabel pdiffusion 1452 -1401 1452 -1401 0 feedthrough
rlabel pdiffusion 1459 -1401 1459 -1401 0 feedthrough
rlabel pdiffusion 1466 -1401 1466 -1401 0 feedthrough
rlabel pdiffusion 1473 -1401 1473 -1401 0 feedthrough
rlabel pdiffusion 1480 -1401 1480 -1401 0 feedthrough
rlabel pdiffusion 1487 -1401 1487 -1401 0 feedthrough
rlabel pdiffusion 1494 -1401 1494 -1401 0 feedthrough
rlabel pdiffusion 1501 -1401 1501 -1401 0 feedthrough
rlabel pdiffusion 1508 -1401 1508 -1401 0 feedthrough
rlabel pdiffusion 1515 -1401 1515 -1401 0 feedthrough
rlabel pdiffusion 1522 -1401 1522 -1401 0 cellNo=32
rlabel pdiffusion 1529 -1401 1529 -1401 0 feedthrough
rlabel pdiffusion 1536 -1401 1536 -1401 0 feedthrough
rlabel pdiffusion 3 -1534 3 -1534 0 feedthrough
rlabel pdiffusion 10 -1534 10 -1534 0 feedthrough
rlabel pdiffusion 17 -1534 17 -1534 0 feedthrough
rlabel pdiffusion 24 -1534 24 -1534 0 feedthrough
rlabel pdiffusion 31 -1534 31 -1534 0 feedthrough
rlabel pdiffusion 38 -1534 38 -1534 0 feedthrough
rlabel pdiffusion 45 -1534 45 -1534 0 feedthrough
rlabel pdiffusion 52 -1534 52 -1534 0 cellNo=236
rlabel pdiffusion 59 -1534 59 -1534 0 feedthrough
rlabel pdiffusion 66 -1534 66 -1534 0 feedthrough
rlabel pdiffusion 73 -1534 73 -1534 0 feedthrough
rlabel pdiffusion 80 -1534 80 -1534 0 cellNo=490
rlabel pdiffusion 87 -1534 87 -1534 0 feedthrough
rlabel pdiffusion 94 -1534 94 -1534 0 feedthrough
rlabel pdiffusion 101 -1534 101 -1534 0 cellNo=284
rlabel pdiffusion 108 -1534 108 -1534 0 feedthrough
rlabel pdiffusion 115 -1534 115 -1534 0 feedthrough
rlabel pdiffusion 122 -1534 122 -1534 0 feedthrough
rlabel pdiffusion 129 -1534 129 -1534 0 feedthrough
rlabel pdiffusion 136 -1534 136 -1534 0 feedthrough
rlabel pdiffusion 143 -1534 143 -1534 0 feedthrough
rlabel pdiffusion 150 -1534 150 -1534 0 feedthrough
rlabel pdiffusion 157 -1534 157 -1534 0 feedthrough
rlabel pdiffusion 164 -1534 164 -1534 0 feedthrough
rlabel pdiffusion 171 -1534 171 -1534 0 cellNo=38
rlabel pdiffusion 178 -1534 178 -1534 0 feedthrough
rlabel pdiffusion 185 -1534 185 -1534 0 feedthrough
rlabel pdiffusion 192 -1534 192 -1534 0 feedthrough
rlabel pdiffusion 199 -1534 199 -1534 0 feedthrough
rlabel pdiffusion 206 -1534 206 -1534 0 feedthrough
rlabel pdiffusion 213 -1534 213 -1534 0 feedthrough
rlabel pdiffusion 220 -1534 220 -1534 0 feedthrough
rlabel pdiffusion 227 -1534 227 -1534 0 feedthrough
rlabel pdiffusion 234 -1534 234 -1534 0 feedthrough
rlabel pdiffusion 241 -1534 241 -1534 0 feedthrough
rlabel pdiffusion 248 -1534 248 -1534 0 feedthrough
rlabel pdiffusion 255 -1534 255 -1534 0 feedthrough
rlabel pdiffusion 262 -1534 262 -1534 0 feedthrough
rlabel pdiffusion 269 -1534 269 -1534 0 feedthrough
rlabel pdiffusion 276 -1534 276 -1534 0 feedthrough
rlabel pdiffusion 283 -1534 283 -1534 0 feedthrough
rlabel pdiffusion 290 -1534 290 -1534 0 feedthrough
rlabel pdiffusion 297 -1534 297 -1534 0 feedthrough
rlabel pdiffusion 304 -1534 304 -1534 0 feedthrough
rlabel pdiffusion 311 -1534 311 -1534 0 feedthrough
rlabel pdiffusion 318 -1534 318 -1534 0 feedthrough
rlabel pdiffusion 325 -1534 325 -1534 0 feedthrough
rlabel pdiffusion 332 -1534 332 -1534 0 feedthrough
rlabel pdiffusion 339 -1534 339 -1534 0 feedthrough
rlabel pdiffusion 346 -1534 346 -1534 0 feedthrough
rlabel pdiffusion 353 -1534 353 -1534 0 feedthrough
rlabel pdiffusion 360 -1534 360 -1534 0 feedthrough
rlabel pdiffusion 367 -1534 367 -1534 0 feedthrough
rlabel pdiffusion 374 -1534 374 -1534 0 feedthrough
rlabel pdiffusion 381 -1534 381 -1534 0 feedthrough
rlabel pdiffusion 388 -1534 388 -1534 0 feedthrough
rlabel pdiffusion 395 -1534 395 -1534 0 cellNo=86
rlabel pdiffusion 402 -1534 402 -1534 0 feedthrough
rlabel pdiffusion 409 -1534 409 -1534 0 feedthrough
rlabel pdiffusion 416 -1534 416 -1534 0 feedthrough
rlabel pdiffusion 423 -1534 423 -1534 0 feedthrough
rlabel pdiffusion 430 -1534 430 -1534 0 cellNo=85
rlabel pdiffusion 437 -1534 437 -1534 0 feedthrough
rlabel pdiffusion 444 -1534 444 -1534 0 feedthrough
rlabel pdiffusion 451 -1534 451 -1534 0 feedthrough
rlabel pdiffusion 458 -1534 458 -1534 0 feedthrough
rlabel pdiffusion 465 -1534 465 -1534 0 feedthrough
rlabel pdiffusion 472 -1534 472 -1534 0 cellNo=190
rlabel pdiffusion 479 -1534 479 -1534 0 feedthrough
rlabel pdiffusion 486 -1534 486 -1534 0 feedthrough
rlabel pdiffusion 493 -1534 493 -1534 0 feedthrough
rlabel pdiffusion 500 -1534 500 -1534 0 cellNo=434
rlabel pdiffusion 507 -1534 507 -1534 0 feedthrough
rlabel pdiffusion 514 -1534 514 -1534 0 feedthrough
rlabel pdiffusion 521 -1534 521 -1534 0 feedthrough
rlabel pdiffusion 528 -1534 528 -1534 0 feedthrough
rlabel pdiffusion 535 -1534 535 -1534 0 feedthrough
rlabel pdiffusion 542 -1534 542 -1534 0 feedthrough
rlabel pdiffusion 549 -1534 549 -1534 0 feedthrough
rlabel pdiffusion 556 -1534 556 -1534 0 feedthrough
rlabel pdiffusion 563 -1534 563 -1534 0 feedthrough
rlabel pdiffusion 570 -1534 570 -1534 0 feedthrough
rlabel pdiffusion 577 -1534 577 -1534 0 cellNo=316
rlabel pdiffusion 584 -1534 584 -1534 0 feedthrough
rlabel pdiffusion 591 -1534 591 -1534 0 feedthrough
rlabel pdiffusion 598 -1534 598 -1534 0 cellNo=44
rlabel pdiffusion 605 -1534 605 -1534 0 feedthrough
rlabel pdiffusion 612 -1534 612 -1534 0 feedthrough
rlabel pdiffusion 619 -1534 619 -1534 0 feedthrough
rlabel pdiffusion 626 -1534 626 -1534 0 feedthrough
rlabel pdiffusion 633 -1534 633 -1534 0 feedthrough
rlabel pdiffusion 640 -1534 640 -1534 0 feedthrough
rlabel pdiffusion 647 -1534 647 -1534 0 feedthrough
rlabel pdiffusion 654 -1534 654 -1534 0 feedthrough
rlabel pdiffusion 661 -1534 661 -1534 0 feedthrough
rlabel pdiffusion 668 -1534 668 -1534 0 feedthrough
rlabel pdiffusion 675 -1534 675 -1534 0 cellNo=325
rlabel pdiffusion 682 -1534 682 -1534 0 cellNo=158
rlabel pdiffusion 689 -1534 689 -1534 0 feedthrough
rlabel pdiffusion 696 -1534 696 -1534 0 feedthrough
rlabel pdiffusion 703 -1534 703 -1534 0 feedthrough
rlabel pdiffusion 710 -1534 710 -1534 0 feedthrough
rlabel pdiffusion 717 -1534 717 -1534 0 feedthrough
rlabel pdiffusion 724 -1534 724 -1534 0 cellNo=74
rlabel pdiffusion 731 -1534 731 -1534 0 feedthrough
rlabel pdiffusion 738 -1534 738 -1534 0 feedthrough
rlabel pdiffusion 745 -1534 745 -1534 0 feedthrough
rlabel pdiffusion 752 -1534 752 -1534 0 feedthrough
rlabel pdiffusion 759 -1534 759 -1534 0 feedthrough
rlabel pdiffusion 766 -1534 766 -1534 0 cellNo=525
rlabel pdiffusion 773 -1534 773 -1534 0 feedthrough
rlabel pdiffusion 780 -1534 780 -1534 0 feedthrough
rlabel pdiffusion 787 -1534 787 -1534 0 feedthrough
rlabel pdiffusion 794 -1534 794 -1534 0 feedthrough
rlabel pdiffusion 801 -1534 801 -1534 0 cellNo=41
rlabel pdiffusion 808 -1534 808 -1534 0 feedthrough
rlabel pdiffusion 815 -1534 815 -1534 0 cellNo=544
rlabel pdiffusion 822 -1534 822 -1534 0 feedthrough
rlabel pdiffusion 829 -1534 829 -1534 0 cellNo=526
rlabel pdiffusion 836 -1534 836 -1534 0 cellNo=177
rlabel pdiffusion 843 -1534 843 -1534 0 feedthrough
rlabel pdiffusion 850 -1534 850 -1534 0 feedthrough
rlabel pdiffusion 857 -1534 857 -1534 0 cellNo=499
rlabel pdiffusion 864 -1534 864 -1534 0 feedthrough
rlabel pdiffusion 871 -1534 871 -1534 0 feedthrough
rlabel pdiffusion 878 -1534 878 -1534 0 cellNo=186
rlabel pdiffusion 885 -1534 885 -1534 0 feedthrough
rlabel pdiffusion 892 -1534 892 -1534 0 feedthrough
rlabel pdiffusion 899 -1534 899 -1534 0 feedthrough
rlabel pdiffusion 906 -1534 906 -1534 0 feedthrough
rlabel pdiffusion 913 -1534 913 -1534 0 feedthrough
rlabel pdiffusion 920 -1534 920 -1534 0 feedthrough
rlabel pdiffusion 927 -1534 927 -1534 0 feedthrough
rlabel pdiffusion 934 -1534 934 -1534 0 feedthrough
rlabel pdiffusion 941 -1534 941 -1534 0 feedthrough
rlabel pdiffusion 948 -1534 948 -1534 0 feedthrough
rlabel pdiffusion 955 -1534 955 -1534 0 feedthrough
rlabel pdiffusion 962 -1534 962 -1534 0 feedthrough
rlabel pdiffusion 969 -1534 969 -1534 0 feedthrough
rlabel pdiffusion 976 -1534 976 -1534 0 feedthrough
rlabel pdiffusion 983 -1534 983 -1534 0 feedthrough
rlabel pdiffusion 990 -1534 990 -1534 0 cellNo=540
rlabel pdiffusion 997 -1534 997 -1534 0 cellNo=215
rlabel pdiffusion 1004 -1534 1004 -1534 0 feedthrough
rlabel pdiffusion 1011 -1534 1011 -1534 0 feedthrough
rlabel pdiffusion 1018 -1534 1018 -1534 0 feedthrough
rlabel pdiffusion 1025 -1534 1025 -1534 0 feedthrough
rlabel pdiffusion 1032 -1534 1032 -1534 0 feedthrough
rlabel pdiffusion 1039 -1534 1039 -1534 0 feedthrough
rlabel pdiffusion 1046 -1534 1046 -1534 0 feedthrough
rlabel pdiffusion 1053 -1534 1053 -1534 0 feedthrough
rlabel pdiffusion 1060 -1534 1060 -1534 0 feedthrough
rlabel pdiffusion 1067 -1534 1067 -1534 0 feedthrough
rlabel pdiffusion 1074 -1534 1074 -1534 0 cellNo=130
rlabel pdiffusion 1081 -1534 1081 -1534 0 feedthrough
rlabel pdiffusion 1088 -1534 1088 -1534 0 feedthrough
rlabel pdiffusion 1095 -1534 1095 -1534 0 feedthrough
rlabel pdiffusion 1102 -1534 1102 -1534 0 feedthrough
rlabel pdiffusion 1109 -1534 1109 -1534 0 feedthrough
rlabel pdiffusion 1116 -1534 1116 -1534 0 feedthrough
rlabel pdiffusion 1123 -1534 1123 -1534 0 cellNo=185
rlabel pdiffusion 1130 -1534 1130 -1534 0 feedthrough
rlabel pdiffusion 1137 -1534 1137 -1534 0 feedthrough
rlabel pdiffusion 1144 -1534 1144 -1534 0 feedthrough
rlabel pdiffusion 1151 -1534 1151 -1534 0 feedthrough
rlabel pdiffusion 1158 -1534 1158 -1534 0 feedthrough
rlabel pdiffusion 1165 -1534 1165 -1534 0 feedthrough
rlabel pdiffusion 1172 -1534 1172 -1534 0 feedthrough
rlabel pdiffusion 1179 -1534 1179 -1534 0 feedthrough
rlabel pdiffusion 1186 -1534 1186 -1534 0 feedthrough
rlabel pdiffusion 1193 -1534 1193 -1534 0 feedthrough
rlabel pdiffusion 1200 -1534 1200 -1534 0 feedthrough
rlabel pdiffusion 1207 -1534 1207 -1534 0 feedthrough
rlabel pdiffusion 1214 -1534 1214 -1534 0 feedthrough
rlabel pdiffusion 1221 -1534 1221 -1534 0 feedthrough
rlabel pdiffusion 1228 -1534 1228 -1534 0 feedthrough
rlabel pdiffusion 1235 -1534 1235 -1534 0 feedthrough
rlabel pdiffusion 1242 -1534 1242 -1534 0 feedthrough
rlabel pdiffusion 1249 -1534 1249 -1534 0 feedthrough
rlabel pdiffusion 1256 -1534 1256 -1534 0 feedthrough
rlabel pdiffusion 1263 -1534 1263 -1534 0 feedthrough
rlabel pdiffusion 1270 -1534 1270 -1534 0 feedthrough
rlabel pdiffusion 1277 -1534 1277 -1534 0 feedthrough
rlabel pdiffusion 1284 -1534 1284 -1534 0 feedthrough
rlabel pdiffusion 1291 -1534 1291 -1534 0 feedthrough
rlabel pdiffusion 1298 -1534 1298 -1534 0 feedthrough
rlabel pdiffusion 1305 -1534 1305 -1534 0 feedthrough
rlabel pdiffusion 1312 -1534 1312 -1534 0 feedthrough
rlabel pdiffusion 1319 -1534 1319 -1534 0 feedthrough
rlabel pdiffusion 1326 -1534 1326 -1534 0 feedthrough
rlabel pdiffusion 1333 -1534 1333 -1534 0 feedthrough
rlabel pdiffusion 1340 -1534 1340 -1534 0 feedthrough
rlabel pdiffusion 1347 -1534 1347 -1534 0 feedthrough
rlabel pdiffusion 1354 -1534 1354 -1534 0 feedthrough
rlabel pdiffusion 1361 -1534 1361 -1534 0 feedthrough
rlabel pdiffusion 1368 -1534 1368 -1534 0 feedthrough
rlabel pdiffusion 1375 -1534 1375 -1534 0 feedthrough
rlabel pdiffusion 1382 -1534 1382 -1534 0 feedthrough
rlabel pdiffusion 1389 -1534 1389 -1534 0 feedthrough
rlabel pdiffusion 1396 -1534 1396 -1534 0 feedthrough
rlabel pdiffusion 1403 -1534 1403 -1534 0 feedthrough
rlabel pdiffusion 1410 -1534 1410 -1534 0 feedthrough
rlabel pdiffusion 1417 -1534 1417 -1534 0 feedthrough
rlabel pdiffusion 1424 -1534 1424 -1534 0 feedthrough
rlabel pdiffusion 1431 -1534 1431 -1534 0 feedthrough
rlabel pdiffusion 1438 -1534 1438 -1534 0 feedthrough
rlabel pdiffusion 1445 -1534 1445 -1534 0 feedthrough
rlabel pdiffusion 1452 -1534 1452 -1534 0 feedthrough
rlabel pdiffusion 1459 -1534 1459 -1534 0 feedthrough
rlabel pdiffusion 1466 -1534 1466 -1534 0 feedthrough
rlabel pdiffusion 1473 -1534 1473 -1534 0 feedthrough
rlabel pdiffusion 1480 -1534 1480 -1534 0 feedthrough
rlabel pdiffusion 1487 -1534 1487 -1534 0 feedthrough
rlabel pdiffusion 1494 -1534 1494 -1534 0 feedthrough
rlabel pdiffusion 1501 -1534 1501 -1534 0 feedthrough
rlabel pdiffusion 1508 -1534 1508 -1534 0 feedthrough
rlabel pdiffusion 1515 -1534 1515 -1534 0 feedthrough
rlabel pdiffusion 1522 -1534 1522 -1534 0 cellNo=178
rlabel pdiffusion 1529 -1534 1529 -1534 0 feedthrough
rlabel pdiffusion 1536 -1534 1536 -1534 0 feedthrough
rlabel pdiffusion 3 -1641 3 -1641 0 feedthrough
rlabel pdiffusion 10 -1641 10 -1641 0 feedthrough
rlabel pdiffusion 17 -1641 17 -1641 0 feedthrough
rlabel pdiffusion 24 -1641 24 -1641 0 feedthrough
rlabel pdiffusion 31 -1641 31 -1641 0 feedthrough
rlabel pdiffusion 38 -1641 38 -1641 0 feedthrough
rlabel pdiffusion 45 -1641 45 -1641 0 feedthrough
rlabel pdiffusion 52 -1641 52 -1641 0 feedthrough
rlabel pdiffusion 59 -1641 59 -1641 0 feedthrough
rlabel pdiffusion 66 -1641 66 -1641 0 feedthrough
rlabel pdiffusion 73 -1641 73 -1641 0 cellNo=46
rlabel pdiffusion 80 -1641 80 -1641 0 feedthrough
rlabel pdiffusion 87 -1641 87 -1641 0 feedthrough
rlabel pdiffusion 94 -1641 94 -1641 0 feedthrough
rlabel pdiffusion 101 -1641 101 -1641 0 feedthrough
rlabel pdiffusion 108 -1641 108 -1641 0 cellNo=146
rlabel pdiffusion 115 -1641 115 -1641 0 feedthrough
rlabel pdiffusion 122 -1641 122 -1641 0 feedthrough
rlabel pdiffusion 129 -1641 129 -1641 0 cellNo=452
rlabel pdiffusion 136 -1641 136 -1641 0 feedthrough
rlabel pdiffusion 143 -1641 143 -1641 0 cellNo=445
rlabel pdiffusion 150 -1641 150 -1641 0 feedthrough
rlabel pdiffusion 157 -1641 157 -1641 0 feedthrough
rlabel pdiffusion 164 -1641 164 -1641 0 feedthrough
rlabel pdiffusion 171 -1641 171 -1641 0 feedthrough
rlabel pdiffusion 178 -1641 178 -1641 0 feedthrough
rlabel pdiffusion 185 -1641 185 -1641 0 feedthrough
rlabel pdiffusion 192 -1641 192 -1641 0 feedthrough
rlabel pdiffusion 199 -1641 199 -1641 0 feedthrough
rlabel pdiffusion 206 -1641 206 -1641 0 feedthrough
rlabel pdiffusion 213 -1641 213 -1641 0 feedthrough
rlabel pdiffusion 220 -1641 220 -1641 0 feedthrough
rlabel pdiffusion 227 -1641 227 -1641 0 feedthrough
rlabel pdiffusion 234 -1641 234 -1641 0 feedthrough
rlabel pdiffusion 241 -1641 241 -1641 0 feedthrough
rlabel pdiffusion 248 -1641 248 -1641 0 feedthrough
rlabel pdiffusion 255 -1641 255 -1641 0 feedthrough
rlabel pdiffusion 262 -1641 262 -1641 0 feedthrough
rlabel pdiffusion 269 -1641 269 -1641 0 cellNo=482
rlabel pdiffusion 276 -1641 276 -1641 0 feedthrough
rlabel pdiffusion 283 -1641 283 -1641 0 feedthrough
rlabel pdiffusion 290 -1641 290 -1641 0 feedthrough
rlabel pdiffusion 297 -1641 297 -1641 0 feedthrough
rlabel pdiffusion 304 -1641 304 -1641 0 feedthrough
rlabel pdiffusion 311 -1641 311 -1641 0 feedthrough
rlabel pdiffusion 318 -1641 318 -1641 0 feedthrough
rlabel pdiffusion 325 -1641 325 -1641 0 feedthrough
rlabel pdiffusion 332 -1641 332 -1641 0 feedthrough
rlabel pdiffusion 339 -1641 339 -1641 0 feedthrough
rlabel pdiffusion 346 -1641 346 -1641 0 cellNo=196
rlabel pdiffusion 353 -1641 353 -1641 0 feedthrough
rlabel pdiffusion 360 -1641 360 -1641 0 feedthrough
rlabel pdiffusion 367 -1641 367 -1641 0 cellNo=161
rlabel pdiffusion 374 -1641 374 -1641 0 feedthrough
rlabel pdiffusion 381 -1641 381 -1641 0 feedthrough
rlabel pdiffusion 388 -1641 388 -1641 0 feedthrough
rlabel pdiffusion 395 -1641 395 -1641 0 feedthrough
rlabel pdiffusion 402 -1641 402 -1641 0 feedthrough
rlabel pdiffusion 409 -1641 409 -1641 0 feedthrough
rlabel pdiffusion 416 -1641 416 -1641 0 feedthrough
rlabel pdiffusion 423 -1641 423 -1641 0 feedthrough
rlabel pdiffusion 430 -1641 430 -1641 0 feedthrough
rlabel pdiffusion 437 -1641 437 -1641 0 cellNo=308
rlabel pdiffusion 444 -1641 444 -1641 0 cellNo=542
rlabel pdiffusion 451 -1641 451 -1641 0 feedthrough
rlabel pdiffusion 458 -1641 458 -1641 0 feedthrough
rlabel pdiffusion 465 -1641 465 -1641 0 feedthrough
rlabel pdiffusion 472 -1641 472 -1641 0 cellNo=532
rlabel pdiffusion 479 -1641 479 -1641 0 feedthrough
rlabel pdiffusion 486 -1641 486 -1641 0 feedthrough
rlabel pdiffusion 493 -1641 493 -1641 0 feedthrough
rlabel pdiffusion 500 -1641 500 -1641 0 cellNo=142
rlabel pdiffusion 507 -1641 507 -1641 0 feedthrough
rlabel pdiffusion 514 -1641 514 -1641 0 feedthrough
rlabel pdiffusion 521 -1641 521 -1641 0 feedthrough
rlabel pdiffusion 528 -1641 528 -1641 0 feedthrough
rlabel pdiffusion 535 -1641 535 -1641 0 feedthrough
rlabel pdiffusion 542 -1641 542 -1641 0 feedthrough
rlabel pdiffusion 549 -1641 549 -1641 0 feedthrough
rlabel pdiffusion 556 -1641 556 -1641 0 cellNo=31
rlabel pdiffusion 563 -1641 563 -1641 0 cellNo=83
rlabel pdiffusion 570 -1641 570 -1641 0 feedthrough
rlabel pdiffusion 577 -1641 577 -1641 0 feedthrough
rlabel pdiffusion 584 -1641 584 -1641 0 feedthrough
rlabel pdiffusion 591 -1641 591 -1641 0 feedthrough
rlabel pdiffusion 598 -1641 598 -1641 0 feedthrough
rlabel pdiffusion 605 -1641 605 -1641 0 feedthrough
rlabel pdiffusion 612 -1641 612 -1641 0 feedthrough
rlabel pdiffusion 619 -1641 619 -1641 0 cellNo=260
rlabel pdiffusion 626 -1641 626 -1641 0 feedthrough
rlabel pdiffusion 633 -1641 633 -1641 0 feedthrough
rlabel pdiffusion 640 -1641 640 -1641 0 feedthrough
rlabel pdiffusion 647 -1641 647 -1641 0 cellNo=448
rlabel pdiffusion 654 -1641 654 -1641 0 feedthrough
rlabel pdiffusion 661 -1641 661 -1641 0 feedthrough
rlabel pdiffusion 668 -1641 668 -1641 0 feedthrough
rlabel pdiffusion 675 -1641 675 -1641 0 feedthrough
rlabel pdiffusion 682 -1641 682 -1641 0 feedthrough
rlabel pdiffusion 689 -1641 689 -1641 0 feedthrough
rlabel pdiffusion 696 -1641 696 -1641 0 feedthrough
rlabel pdiffusion 703 -1641 703 -1641 0 feedthrough
rlabel pdiffusion 710 -1641 710 -1641 0 feedthrough
rlabel pdiffusion 717 -1641 717 -1641 0 feedthrough
rlabel pdiffusion 724 -1641 724 -1641 0 feedthrough
rlabel pdiffusion 731 -1641 731 -1641 0 feedthrough
rlabel pdiffusion 738 -1641 738 -1641 0 cellNo=94
rlabel pdiffusion 745 -1641 745 -1641 0 feedthrough
rlabel pdiffusion 752 -1641 752 -1641 0 cellNo=408
rlabel pdiffusion 759 -1641 759 -1641 0 feedthrough
rlabel pdiffusion 766 -1641 766 -1641 0 feedthrough
rlabel pdiffusion 773 -1641 773 -1641 0 feedthrough
rlabel pdiffusion 780 -1641 780 -1641 0 cellNo=406
rlabel pdiffusion 787 -1641 787 -1641 0 feedthrough
rlabel pdiffusion 794 -1641 794 -1641 0 feedthrough
rlabel pdiffusion 801 -1641 801 -1641 0 feedthrough
rlabel pdiffusion 808 -1641 808 -1641 0 feedthrough
rlabel pdiffusion 815 -1641 815 -1641 0 cellNo=382
rlabel pdiffusion 822 -1641 822 -1641 0 feedthrough
rlabel pdiffusion 829 -1641 829 -1641 0 cellNo=93
rlabel pdiffusion 836 -1641 836 -1641 0 feedthrough
rlabel pdiffusion 843 -1641 843 -1641 0 feedthrough
rlabel pdiffusion 850 -1641 850 -1641 0 feedthrough
rlabel pdiffusion 857 -1641 857 -1641 0 feedthrough
rlabel pdiffusion 864 -1641 864 -1641 0 feedthrough
rlabel pdiffusion 871 -1641 871 -1641 0 feedthrough
rlabel pdiffusion 878 -1641 878 -1641 0 cellNo=336
rlabel pdiffusion 885 -1641 885 -1641 0 feedthrough
rlabel pdiffusion 892 -1641 892 -1641 0 feedthrough
rlabel pdiffusion 899 -1641 899 -1641 0 feedthrough
rlabel pdiffusion 906 -1641 906 -1641 0 feedthrough
rlabel pdiffusion 913 -1641 913 -1641 0 feedthrough
rlabel pdiffusion 920 -1641 920 -1641 0 feedthrough
rlabel pdiffusion 927 -1641 927 -1641 0 feedthrough
rlabel pdiffusion 934 -1641 934 -1641 0 feedthrough
rlabel pdiffusion 941 -1641 941 -1641 0 feedthrough
rlabel pdiffusion 948 -1641 948 -1641 0 feedthrough
rlabel pdiffusion 955 -1641 955 -1641 0 cellNo=270
rlabel pdiffusion 962 -1641 962 -1641 0 feedthrough
rlabel pdiffusion 969 -1641 969 -1641 0 feedthrough
rlabel pdiffusion 976 -1641 976 -1641 0 feedthrough
rlabel pdiffusion 983 -1641 983 -1641 0 feedthrough
rlabel pdiffusion 990 -1641 990 -1641 0 cellNo=155
rlabel pdiffusion 997 -1641 997 -1641 0 feedthrough
rlabel pdiffusion 1004 -1641 1004 -1641 0 feedthrough
rlabel pdiffusion 1011 -1641 1011 -1641 0 feedthrough
rlabel pdiffusion 1018 -1641 1018 -1641 0 feedthrough
rlabel pdiffusion 1025 -1641 1025 -1641 0 feedthrough
rlabel pdiffusion 1032 -1641 1032 -1641 0 feedthrough
rlabel pdiffusion 1039 -1641 1039 -1641 0 feedthrough
rlabel pdiffusion 1046 -1641 1046 -1641 0 feedthrough
rlabel pdiffusion 1053 -1641 1053 -1641 0 feedthrough
rlabel pdiffusion 1060 -1641 1060 -1641 0 feedthrough
rlabel pdiffusion 1067 -1641 1067 -1641 0 feedthrough
rlabel pdiffusion 1074 -1641 1074 -1641 0 feedthrough
rlabel pdiffusion 1081 -1641 1081 -1641 0 feedthrough
rlabel pdiffusion 1088 -1641 1088 -1641 0 feedthrough
rlabel pdiffusion 1095 -1641 1095 -1641 0 feedthrough
rlabel pdiffusion 1102 -1641 1102 -1641 0 feedthrough
rlabel pdiffusion 1109 -1641 1109 -1641 0 feedthrough
rlabel pdiffusion 1116 -1641 1116 -1641 0 feedthrough
rlabel pdiffusion 1123 -1641 1123 -1641 0 feedthrough
rlabel pdiffusion 1130 -1641 1130 -1641 0 feedthrough
rlabel pdiffusion 1137 -1641 1137 -1641 0 feedthrough
rlabel pdiffusion 1144 -1641 1144 -1641 0 feedthrough
rlabel pdiffusion 1151 -1641 1151 -1641 0 feedthrough
rlabel pdiffusion 1158 -1641 1158 -1641 0 feedthrough
rlabel pdiffusion 1165 -1641 1165 -1641 0 feedthrough
rlabel pdiffusion 1172 -1641 1172 -1641 0 feedthrough
rlabel pdiffusion 1179 -1641 1179 -1641 0 feedthrough
rlabel pdiffusion 1186 -1641 1186 -1641 0 feedthrough
rlabel pdiffusion 1193 -1641 1193 -1641 0 feedthrough
rlabel pdiffusion 1200 -1641 1200 -1641 0 feedthrough
rlabel pdiffusion 1207 -1641 1207 -1641 0 feedthrough
rlabel pdiffusion 1214 -1641 1214 -1641 0 feedthrough
rlabel pdiffusion 1221 -1641 1221 -1641 0 feedthrough
rlabel pdiffusion 1228 -1641 1228 -1641 0 feedthrough
rlabel pdiffusion 1235 -1641 1235 -1641 0 feedthrough
rlabel pdiffusion 1242 -1641 1242 -1641 0 feedthrough
rlabel pdiffusion 1249 -1641 1249 -1641 0 feedthrough
rlabel pdiffusion 1256 -1641 1256 -1641 0 feedthrough
rlabel pdiffusion 1263 -1641 1263 -1641 0 feedthrough
rlabel pdiffusion 1270 -1641 1270 -1641 0 feedthrough
rlabel pdiffusion 1277 -1641 1277 -1641 0 feedthrough
rlabel pdiffusion 1284 -1641 1284 -1641 0 feedthrough
rlabel pdiffusion 1291 -1641 1291 -1641 0 feedthrough
rlabel pdiffusion 1298 -1641 1298 -1641 0 feedthrough
rlabel pdiffusion 1305 -1641 1305 -1641 0 feedthrough
rlabel pdiffusion 1312 -1641 1312 -1641 0 feedthrough
rlabel pdiffusion 1319 -1641 1319 -1641 0 feedthrough
rlabel pdiffusion 1326 -1641 1326 -1641 0 feedthrough
rlabel pdiffusion 1333 -1641 1333 -1641 0 feedthrough
rlabel pdiffusion 1340 -1641 1340 -1641 0 feedthrough
rlabel pdiffusion 1347 -1641 1347 -1641 0 cellNo=100
rlabel pdiffusion 1354 -1641 1354 -1641 0 feedthrough
rlabel pdiffusion 1361 -1641 1361 -1641 0 feedthrough
rlabel pdiffusion 1368 -1641 1368 -1641 0 feedthrough
rlabel pdiffusion 1375 -1641 1375 -1641 0 feedthrough
rlabel pdiffusion 1382 -1641 1382 -1641 0 feedthrough
rlabel pdiffusion 1389 -1641 1389 -1641 0 feedthrough
rlabel pdiffusion 1396 -1641 1396 -1641 0 cellNo=431
rlabel pdiffusion 1403 -1641 1403 -1641 0 feedthrough
rlabel pdiffusion 1410 -1641 1410 -1641 0 feedthrough
rlabel pdiffusion 1417 -1641 1417 -1641 0 feedthrough
rlabel pdiffusion 1424 -1641 1424 -1641 0 feedthrough
rlabel pdiffusion 1431 -1641 1431 -1641 0 feedthrough
rlabel pdiffusion 1438 -1641 1438 -1641 0 feedthrough
rlabel pdiffusion 1452 -1641 1452 -1641 0 feedthrough
rlabel pdiffusion 10 -1766 10 -1766 0 feedthrough
rlabel pdiffusion 17 -1766 17 -1766 0 feedthrough
rlabel pdiffusion 24 -1766 24 -1766 0 feedthrough
rlabel pdiffusion 31 -1766 31 -1766 0 feedthrough
rlabel pdiffusion 38 -1766 38 -1766 0 feedthrough
rlabel pdiffusion 45 -1766 45 -1766 0 feedthrough
rlabel pdiffusion 52 -1766 52 -1766 0 feedthrough
rlabel pdiffusion 59 -1766 59 -1766 0 feedthrough
rlabel pdiffusion 66 -1766 66 -1766 0 feedthrough
rlabel pdiffusion 73 -1766 73 -1766 0 cellNo=135
rlabel pdiffusion 80 -1766 80 -1766 0 cellNo=246
rlabel pdiffusion 87 -1766 87 -1766 0 feedthrough
rlabel pdiffusion 94 -1766 94 -1766 0 feedthrough
rlabel pdiffusion 101 -1766 101 -1766 0 feedthrough
rlabel pdiffusion 108 -1766 108 -1766 0 cellNo=79
rlabel pdiffusion 115 -1766 115 -1766 0 feedthrough
rlabel pdiffusion 122 -1766 122 -1766 0 feedthrough
rlabel pdiffusion 129 -1766 129 -1766 0 feedthrough
rlabel pdiffusion 136 -1766 136 -1766 0 feedthrough
rlabel pdiffusion 143 -1766 143 -1766 0 feedthrough
rlabel pdiffusion 150 -1766 150 -1766 0 feedthrough
rlabel pdiffusion 157 -1766 157 -1766 0 feedthrough
rlabel pdiffusion 164 -1766 164 -1766 0 feedthrough
rlabel pdiffusion 171 -1766 171 -1766 0 feedthrough
rlabel pdiffusion 178 -1766 178 -1766 0 feedthrough
rlabel pdiffusion 185 -1766 185 -1766 0 feedthrough
rlabel pdiffusion 192 -1766 192 -1766 0 feedthrough
rlabel pdiffusion 199 -1766 199 -1766 0 feedthrough
rlabel pdiffusion 206 -1766 206 -1766 0 feedthrough
rlabel pdiffusion 213 -1766 213 -1766 0 feedthrough
rlabel pdiffusion 220 -1766 220 -1766 0 feedthrough
rlabel pdiffusion 227 -1766 227 -1766 0 feedthrough
rlabel pdiffusion 234 -1766 234 -1766 0 feedthrough
rlabel pdiffusion 241 -1766 241 -1766 0 feedthrough
rlabel pdiffusion 248 -1766 248 -1766 0 feedthrough
rlabel pdiffusion 255 -1766 255 -1766 0 feedthrough
rlabel pdiffusion 262 -1766 262 -1766 0 feedthrough
rlabel pdiffusion 269 -1766 269 -1766 0 feedthrough
rlabel pdiffusion 276 -1766 276 -1766 0 feedthrough
rlabel pdiffusion 283 -1766 283 -1766 0 feedthrough
rlabel pdiffusion 290 -1766 290 -1766 0 feedthrough
rlabel pdiffusion 297 -1766 297 -1766 0 feedthrough
rlabel pdiffusion 304 -1766 304 -1766 0 feedthrough
rlabel pdiffusion 311 -1766 311 -1766 0 feedthrough
rlabel pdiffusion 318 -1766 318 -1766 0 feedthrough
rlabel pdiffusion 325 -1766 325 -1766 0 feedthrough
rlabel pdiffusion 332 -1766 332 -1766 0 feedthrough
rlabel pdiffusion 339 -1766 339 -1766 0 cellNo=180
rlabel pdiffusion 346 -1766 346 -1766 0 feedthrough
rlabel pdiffusion 353 -1766 353 -1766 0 feedthrough
rlabel pdiffusion 360 -1766 360 -1766 0 feedthrough
rlabel pdiffusion 367 -1766 367 -1766 0 cellNo=375
rlabel pdiffusion 374 -1766 374 -1766 0 feedthrough
rlabel pdiffusion 381 -1766 381 -1766 0 feedthrough
rlabel pdiffusion 388 -1766 388 -1766 0 feedthrough
rlabel pdiffusion 395 -1766 395 -1766 0 feedthrough
rlabel pdiffusion 402 -1766 402 -1766 0 feedthrough
rlabel pdiffusion 409 -1766 409 -1766 0 feedthrough
rlabel pdiffusion 416 -1766 416 -1766 0 cellNo=299
rlabel pdiffusion 423 -1766 423 -1766 0 cellNo=462
rlabel pdiffusion 430 -1766 430 -1766 0 feedthrough
rlabel pdiffusion 437 -1766 437 -1766 0 feedthrough
rlabel pdiffusion 444 -1766 444 -1766 0 feedthrough
rlabel pdiffusion 451 -1766 451 -1766 0 feedthrough
rlabel pdiffusion 458 -1766 458 -1766 0 feedthrough
rlabel pdiffusion 465 -1766 465 -1766 0 feedthrough
rlabel pdiffusion 472 -1766 472 -1766 0 feedthrough
rlabel pdiffusion 479 -1766 479 -1766 0 feedthrough
rlabel pdiffusion 486 -1766 486 -1766 0 cellNo=472
rlabel pdiffusion 493 -1766 493 -1766 0 feedthrough
rlabel pdiffusion 500 -1766 500 -1766 0 feedthrough
rlabel pdiffusion 507 -1766 507 -1766 0 cellNo=168
rlabel pdiffusion 514 -1766 514 -1766 0 feedthrough
rlabel pdiffusion 521 -1766 521 -1766 0 cellNo=48
rlabel pdiffusion 528 -1766 528 -1766 0 cellNo=388
rlabel pdiffusion 535 -1766 535 -1766 0 feedthrough
rlabel pdiffusion 542 -1766 542 -1766 0 feedthrough
rlabel pdiffusion 549 -1766 549 -1766 0 feedthrough
rlabel pdiffusion 556 -1766 556 -1766 0 feedthrough
rlabel pdiffusion 563 -1766 563 -1766 0 feedthrough
rlabel pdiffusion 570 -1766 570 -1766 0 feedthrough
rlabel pdiffusion 577 -1766 577 -1766 0 feedthrough
rlabel pdiffusion 584 -1766 584 -1766 0 cellNo=582
rlabel pdiffusion 591 -1766 591 -1766 0 feedthrough
rlabel pdiffusion 598 -1766 598 -1766 0 feedthrough
rlabel pdiffusion 605 -1766 605 -1766 0 feedthrough
rlabel pdiffusion 612 -1766 612 -1766 0 feedthrough
rlabel pdiffusion 619 -1766 619 -1766 0 feedthrough
rlabel pdiffusion 626 -1766 626 -1766 0 feedthrough
rlabel pdiffusion 633 -1766 633 -1766 0 cellNo=370
rlabel pdiffusion 640 -1766 640 -1766 0 feedthrough
rlabel pdiffusion 647 -1766 647 -1766 0 feedthrough
rlabel pdiffusion 654 -1766 654 -1766 0 feedthrough
rlabel pdiffusion 661 -1766 661 -1766 0 feedthrough
rlabel pdiffusion 668 -1766 668 -1766 0 feedthrough
rlabel pdiffusion 675 -1766 675 -1766 0 feedthrough
rlabel pdiffusion 682 -1766 682 -1766 0 feedthrough
rlabel pdiffusion 689 -1766 689 -1766 0 feedthrough
rlabel pdiffusion 696 -1766 696 -1766 0 feedthrough
rlabel pdiffusion 703 -1766 703 -1766 0 feedthrough
rlabel pdiffusion 710 -1766 710 -1766 0 feedthrough
rlabel pdiffusion 717 -1766 717 -1766 0 cellNo=541
rlabel pdiffusion 724 -1766 724 -1766 0 feedthrough
rlabel pdiffusion 731 -1766 731 -1766 0 feedthrough
rlabel pdiffusion 738 -1766 738 -1766 0 feedthrough
rlabel pdiffusion 745 -1766 745 -1766 0 feedthrough
rlabel pdiffusion 752 -1766 752 -1766 0 feedthrough
rlabel pdiffusion 759 -1766 759 -1766 0 feedthrough
rlabel pdiffusion 766 -1766 766 -1766 0 feedthrough
rlabel pdiffusion 773 -1766 773 -1766 0 cellNo=57
rlabel pdiffusion 780 -1766 780 -1766 0 feedthrough
rlabel pdiffusion 787 -1766 787 -1766 0 feedthrough
rlabel pdiffusion 794 -1766 794 -1766 0 cellNo=488
rlabel pdiffusion 801 -1766 801 -1766 0 feedthrough
rlabel pdiffusion 808 -1766 808 -1766 0 cellNo=118
rlabel pdiffusion 815 -1766 815 -1766 0 feedthrough
rlabel pdiffusion 822 -1766 822 -1766 0 feedthrough
rlabel pdiffusion 829 -1766 829 -1766 0 feedthrough
rlabel pdiffusion 836 -1766 836 -1766 0 feedthrough
rlabel pdiffusion 843 -1766 843 -1766 0 cellNo=58
rlabel pdiffusion 850 -1766 850 -1766 0 feedthrough
rlabel pdiffusion 857 -1766 857 -1766 0 feedthrough
rlabel pdiffusion 864 -1766 864 -1766 0 feedthrough
rlabel pdiffusion 871 -1766 871 -1766 0 cellNo=403
rlabel pdiffusion 878 -1766 878 -1766 0 cellNo=217
rlabel pdiffusion 885 -1766 885 -1766 0 feedthrough
rlabel pdiffusion 892 -1766 892 -1766 0 feedthrough
rlabel pdiffusion 899 -1766 899 -1766 0 cellNo=138
rlabel pdiffusion 906 -1766 906 -1766 0 feedthrough
rlabel pdiffusion 913 -1766 913 -1766 0 feedthrough
rlabel pdiffusion 920 -1766 920 -1766 0 feedthrough
rlabel pdiffusion 927 -1766 927 -1766 0 feedthrough
rlabel pdiffusion 934 -1766 934 -1766 0 feedthrough
rlabel pdiffusion 941 -1766 941 -1766 0 feedthrough
rlabel pdiffusion 948 -1766 948 -1766 0 feedthrough
rlabel pdiffusion 955 -1766 955 -1766 0 feedthrough
rlabel pdiffusion 962 -1766 962 -1766 0 feedthrough
rlabel pdiffusion 969 -1766 969 -1766 0 feedthrough
rlabel pdiffusion 976 -1766 976 -1766 0 feedthrough
rlabel pdiffusion 983 -1766 983 -1766 0 feedthrough
rlabel pdiffusion 990 -1766 990 -1766 0 cellNo=524
rlabel pdiffusion 997 -1766 997 -1766 0 feedthrough
rlabel pdiffusion 1004 -1766 1004 -1766 0 cellNo=131
rlabel pdiffusion 1011 -1766 1011 -1766 0 feedthrough
rlabel pdiffusion 1018 -1766 1018 -1766 0 feedthrough
rlabel pdiffusion 1025 -1766 1025 -1766 0 feedthrough
rlabel pdiffusion 1032 -1766 1032 -1766 0 feedthrough
rlabel pdiffusion 1039 -1766 1039 -1766 0 feedthrough
rlabel pdiffusion 1046 -1766 1046 -1766 0 feedthrough
rlabel pdiffusion 1053 -1766 1053 -1766 0 feedthrough
rlabel pdiffusion 1060 -1766 1060 -1766 0 feedthrough
rlabel pdiffusion 1067 -1766 1067 -1766 0 feedthrough
rlabel pdiffusion 1074 -1766 1074 -1766 0 feedthrough
rlabel pdiffusion 1081 -1766 1081 -1766 0 feedthrough
rlabel pdiffusion 1088 -1766 1088 -1766 0 feedthrough
rlabel pdiffusion 1095 -1766 1095 -1766 0 feedthrough
rlabel pdiffusion 1102 -1766 1102 -1766 0 feedthrough
rlabel pdiffusion 1109 -1766 1109 -1766 0 feedthrough
rlabel pdiffusion 1116 -1766 1116 -1766 0 feedthrough
rlabel pdiffusion 1123 -1766 1123 -1766 0 feedthrough
rlabel pdiffusion 1130 -1766 1130 -1766 0 feedthrough
rlabel pdiffusion 1137 -1766 1137 -1766 0 feedthrough
rlabel pdiffusion 1144 -1766 1144 -1766 0 feedthrough
rlabel pdiffusion 1151 -1766 1151 -1766 0 feedthrough
rlabel pdiffusion 1158 -1766 1158 -1766 0 feedthrough
rlabel pdiffusion 1165 -1766 1165 -1766 0 feedthrough
rlabel pdiffusion 1172 -1766 1172 -1766 0 feedthrough
rlabel pdiffusion 1179 -1766 1179 -1766 0 feedthrough
rlabel pdiffusion 1186 -1766 1186 -1766 0 feedthrough
rlabel pdiffusion 1193 -1766 1193 -1766 0 feedthrough
rlabel pdiffusion 1200 -1766 1200 -1766 0 feedthrough
rlabel pdiffusion 1207 -1766 1207 -1766 0 feedthrough
rlabel pdiffusion 1214 -1766 1214 -1766 0 feedthrough
rlabel pdiffusion 1221 -1766 1221 -1766 0 feedthrough
rlabel pdiffusion 1228 -1766 1228 -1766 0 feedthrough
rlabel pdiffusion 1235 -1766 1235 -1766 0 feedthrough
rlabel pdiffusion 1242 -1766 1242 -1766 0 feedthrough
rlabel pdiffusion 1249 -1766 1249 -1766 0 feedthrough
rlabel pdiffusion 1256 -1766 1256 -1766 0 feedthrough
rlabel pdiffusion 1263 -1766 1263 -1766 0 feedthrough
rlabel pdiffusion 1270 -1766 1270 -1766 0 feedthrough
rlabel pdiffusion 1277 -1766 1277 -1766 0 feedthrough
rlabel pdiffusion 1284 -1766 1284 -1766 0 feedthrough
rlabel pdiffusion 1291 -1766 1291 -1766 0 feedthrough
rlabel pdiffusion 1298 -1766 1298 -1766 0 feedthrough
rlabel pdiffusion 1305 -1766 1305 -1766 0 feedthrough
rlabel pdiffusion 1312 -1766 1312 -1766 0 feedthrough
rlabel pdiffusion 1319 -1766 1319 -1766 0 feedthrough
rlabel pdiffusion 1326 -1766 1326 -1766 0 feedthrough
rlabel pdiffusion 1333 -1766 1333 -1766 0 feedthrough
rlabel pdiffusion 1340 -1766 1340 -1766 0 feedthrough
rlabel pdiffusion 1347 -1766 1347 -1766 0 feedthrough
rlabel pdiffusion 1354 -1766 1354 -1766 0 feedthrough
rlabel pdiffusion 1361 -1766 1361 -1766 0 feedthrough
rlabel pdiffusion 1368 -1766 1368 -1766 0 cellNo=305
rlabel pdiffusion 1375 -1766 1375 -1766 0 cellNo=228
rlabel pdiffusion 1382 -1766 1382 -1766 0 feedthrough
rlabel pdiffusion 1389 -1766 1389 -1766 0 feedthrough
rlabel pdiffusion 1396 -1766 1396 -1766 0 feedthrough
rlabel pdiffusion 1403 -1766 1403 -1766 0 feedthrough
rlabel pdiffusion 1410 -1766 1410 -1766 0 feedthrough
rlabel pdiffusion 1417 -1766 1417 -1766 0 feedthrough
rlabel pdiffusion 1424 -1766 1424 -1766 0 feedthrough
rlabel pdiffusion 3 -1863 3 -1863 0 feedthrough
rlabel pdiffusion 10 -1863 10 -1863 0 feedthrough
rlabel pdiffusion 17 -1863 17 -1863 0 cellNo=379
rlabel pdiffusion 24 -1863 24 -1863 0 feedthrough
rlabel pdiffusion 31 -1863 31 -1863 0 feedthrough
rlabel pdiffusion 38 -1863 38 -1863 0 feedthrough
rlabel pdiffusion 45 -1863 45 -1863 0 feedthrough
rlabel pdiffusion 52 -1863 52 -1863 0 feedthrough
rlabel pdiffusion 59 -1863 59 -1863 0 cellNo=150
rlabel pdiffusion 66 -1863 66 -1863 0 feedthrough
rlabel pdiffusion 73 -1863 73 -1863 0 feedthrough
rlabel pdiffusion 80 -1863 80 -1863 0 feedthrough
rlabel pdiffusion 87 -1863 87 -1863 0 cellNo=136
rlabel pdiffusion 94 -1863 94 -1863 0 feedthrough
rlabel pdiffusion 101 -1863 101 -1863 0 feedthrough
rlabel pdiffusion 108 -1863 108 -1863 0 feedthrough
rlabel pdiffusion 115 -1863 115 -1863 0 feedthrough
rlabel pdiffusion 122 -1863 122 -1863 0 feedthrough
rlabel pdiffusion 129 -1863 129 -1863 0 feedthrough
rlabel pdiffusion 136 -1863 136 -1863 0 cellNo=105
rlabel pdiffusion 143 -1863 143 -1863 0 feedthrough
rlabel pdiffusion 150 -1863 150 -1863 0 feedthrough
rlabel pdiffusion 157 -1863 157 -1863 0 feedthrough
rlabel pdiffusion 164 -1863 164 -1863 0 feedthrough
rlabel pdiffusion 171 -1863 171 -1863 0 feedthrough
rlabel pdiffusion 178 -1863 178 -1863 0 feedthrough
rlabel pdiffusion 185 -1863 185 -1863 0 feedthrough
rlabel pdiffusion 192 -1863 192 -1863 0 feedthrough
rlabel pdiffusion 199 -1863 199 -1863 0 feedthrough
rlabel pdiffusion 206 -1863 206 -1863 0 feedthrough
rlabel pdiffusion 213 -1863 213 -1863 0 feedthrough
rlabel pdiffusion 220 -1863 220 -1863 0 feedthrough
rlabel pdiffusion 227 -1863 227 -1863 0 feedthrough
rlabel pdiffusion 234 -1863 234 -1863 0 feedthrough
rlabel pdiffusion 241 -1863 241 -1863 0 feedthrough
rlabel pdiffusion 248 -1863 248 -1863 0 feedthrough
rlabel pdiffusion 255 -1863 255 -1863 0 feedthrough
rlabel pdiffusion 262 -1863 262 -1863 0 feedthrough
rlabel pdiffusion 269 -1863 269 -1863 0 feedthrough
rlabel pdiffusion 276 -1863 276 -1863 0 feedthrough
rlabel pdiffusion 283 -1863 283 -1863 0 feedthrough
rlabel pdiffusion 290 -1863 290 -1863 0 feedthrough
rlabel pdiffusion 297 -1863 297 -1863 0 cellNo=13
rlabel pdiffusion 304 -1863 304 -1863 0 feedthrough
rlabel pdiffusion 311 -1863 311 -1863 0 feedthrough
rlabel pdiffusion 318 -1863 318 -1863 0 feedthrough
rlabel pdiffusion 325 -1863 325 -1863 0 feedthrough
rlabel pdiffusion 332 -1863 332 -1863 0 feedthrough
rlabel pdiffusion 339 -1863 339 -1863 0 feedthrough
rlabel pdiffusion 346 -1863 346 -1863 0 cellNo=211
rlabel pdiffusion 353 -1863 353 -1863 0 feedthrough
rlabel pdiffusion 360 -1863 360 -1863 0 feedthrough
rlabel pdiffusion 367 -1863 367 -1863 0 feedthrough
rlabel pdiffusion 374 -1863 374 -1863 0 feedthrough
rlabel pdiffusion 381 -1863 381 -1863 0 feedthrough
rlabel pdiffusion 388 -1863 388 -1863 0 feedthrough
rlabel pdiffusion 395 -1863 395 -1863 0 cellNo=523
rlabel pdiffusion 402 -1863 402 -1863 0 feedthrough
rlabel pdiffusion 409 -1863 409 -1863 0 feedthrough
rlabel pdiffusion 416 -1863 416 -1863 0 feedthrough
rlabel pdiffusion 423 -1863 423 -1863 0 feedthrough
rlabel pdiffusion 430 -1863 430 -1863 0 cellNo=507
rlabel pdiffusion 437 -1863 437 -1863 0 feedthrough
rlabel pdiffusion 444 -1863 444 -1863 0 feedthrough
rlabel pdiffusion 451 -1863 451 -1863 0 feedthrough
rlabel pdiffusion 458 -1863 458 -1863 0 feedthrough
rlabel pdiffusion 465 -1863 465 -1863 0 feedthrough
rlabel pdiffusion 472 -1863 472 -1863 0 feedthrough
rlabel pdiffusion 479 -1863 479 -1863 0 feedthrough
rlabel pdiffusion 486 -1863 486 -1863 0 feedthrough
rlabel pdiffusion 493 -1863 493 -1863 0 feedthrough
rlabel pdiffusion 500 -1863 500 -1863 0 cellNo=226
rlabel pdiffusion 507 -1863 507 -1863 0 feedthrough
rlabel pdiffusion 514 -1863 514 -1863 0 feedthrough
rlabel pdiffusion 521 -1863 521 -1863 0 feedthrough
rlabel pdiffusion 528 -1863 528 -1863 0 feedthrough
rlabel pdiffusion 535 -1863 535 -1863 0 feedthrough
rlabel pdiffusion 542 -1863 542 -1863 0 feedthrough
rlabel pdiffusion 549 -1863 549 -1863 0 feedthrough
rlabel pdiffusion 556 -1863 556 -1863 0 cellNo=306
rlabel pdiffusion 563 -1863 563 -1863 0 feedthrough
rlabel pdiffusion 570 -1863 570 -1863 0 cellNo=459
rlabel pdiffusion 577 -1863 577 -1863 0 feedthrough
rlabel pdiffusion 584 -1863 584 -1863 0 feedthrough
rlabel pdiffusion 591 -1863 591 -1863 0 cellNo=27
rlabel pdiffusion 598 -1863 598 -1863 0 feedthrough
rlabel pdiffusion 605 -1863 605 -1863 0 feedthrough
rlabel pdiffusion 612 -1863 612 -1863 0 feedthrough
rlabel pdiffusion 619 -1863 619 -1863 0 feedthrough
rlabel pdiffusion 626 -1863 626 -1863 0 feedthrough
rlabel pdiffusion 633 -1863 633 -1863 0 feedthrough
rlabel pdiffusion 640 -1863 640 -1863 0 feedthrough
rlabel pdiffusion 647 -1863 647 -1863 0 feedthrough
rlabel pdiffusion 654 -1863 654 -1863 0 feedthrough
rlabel pdiffusion 661 -1863 661 -1863 0 cellNo=289
rlabel pdiffusion 668 -1863 668 -1863 0 feedthrough
rlabel pdiffusion 675 -1863 675 -1863 0 feedthrough
rlabel pdiffusion 682 -1863 682 -1863 0 cellNo=438
rlabel pdiffusion 689 -1863 689 -1863 0 cellNo=495
rlabel pdiffusion 696 -1863 696 -1863 0 feedthrough
rlabel pdiffusion 703 -1863 703 -1863 0 feedthrough
rlabel pdiffusion 710 -1863 710 -1863 0 feedthrough
rlabel pdiffusion 717 -1863 717 -1863 0 cellNo=279
rlabel pdiffusion 724 -1863 724 -1863 0 feedthrough
rlabel pdiffusion 731 -1863 731 -1863 0 feedthrough
rlabel pdiffusion 738 -1863 738 -1863 0 feedthrough
rlabel pdiffusion 745 -1863 745 -1863 0 feedthrough
rlabel pdiffusion 752 -1863 752 -1863 0 cellNo=558
rlabel pdiffusion 759 -1863 759 -1863 0 feedthrough
rlabel pdiffusion 766 -1863 766 -1863 0 feedthrough
rlabel pdiffusion 773 -1863 773 -1863 0 cellNo=521
rlabel pdiffusion 780 -1863 780 -1863 0 feedthrough
rlabel pdiffusion 787 -1863 787 -1863 0 feedthrough
rlabel pdiffusion 794 -1863 794 -1863 0 feedthrough
rlabel pdiffusion 801 -1863 801 -1863 0 cellNo=119
rlabel pdiffusion 808 -1863 808 -1863 0 feedthrough
rlabel pdiffusion 815 -1863 815 -1863 0 feedthrough
rlabel pdiffusion 822 -1863 822 -1863 0 feedthrough
rlabel pdiffusion 829 -1863 829 -1863 0 feedthrough
rlabel pdiffusion 836 -1863 836 -1863 0 feedthrough
rlabel pdiffusion 843 -1863 843 -1863 0 feedthrough
rlabel pdiffusion 850 -1863 850 -1863 0 feedthrough
rlabel pdiffusion 857 -1863 857 -1863 0 feedthrough
rlabel pdiffusion 864 -1863 864 -1863 0 feedthrough
rlabel pdiffusion 871 -1863 871 -1863 0 feedthrough
rlabel pdiffusion 878 -1863 878 -1863 0 feedthrough
rlabel pdiffusion 885 -1863 885 -1863 0 cellNo=520
rlabel pdiffusion 892 -1863 892 -1863 0 feedthrough
rlabel pdiffusion 899 -1863 899 -1863 0 feedthrough
rlabel pdiffusion 906 -1863 906 -1863 0 cellNo=250
rlabel pdiffusion 913 -1863 913 -1863 0 feedthrough
rlabel pdiffusion 920 -1863 920 -1863 0 feedthrough
rlabel pdiffusion 927 -1863 927 -1863 0 feedthrough
rlabel pdiffusion 934 -1863 934 -1863 0 cellNo=560
rlabel pdiffusion 941 -1863 941 -1863 0 feedthrough
rlabel pdiffusion 948 -1863 948 -1863 0 feedthrough
rlabel pdiffusion 955 -1863 955 -1863 0 feedthrough
rlabel pdiffusion 962 -1863 962 -1863 0 feedthrough
rlabel pdiffusion 969 -1863 969 -1863 0 feedthrough
rlabel pdiffusion 976 -1863 976 -1863 0 feedthrough
rlabel pdiffusion 983 -1863 983 -1863 0 feedthrough
rlabel pdiffusion 990 -1863 990 -1863 0 feedthrough
rlabel pdiffusion 997 -1863 997 -1863 0 feedthrough
rlabel pdiffusion 1004 -1863 1004 -1863 0 feedthrough
rlabel pdiffusion 1011 -1863 1011 -1863 0 feedthrough
rlabel pdiffusion 1018 -1863 1018 -1863 0 feedthrough
rlabel pdiffusion 1025 -1863 1025 -1863 0 feedthrough
rlabel pdiffusion 1032 -1863 1032 -1863 0 feedthrough
rlabel pdiffusion 1039 -1863 1039 -1863 0 feedthrough
rlabel pdiffusion 1046 -1863 1046 -1863 0 feedthrough
rlabel pdiffusion 1053 -1863 1053 -1863 0 feedthrough
rlabel pdiffusion 1060 -1863 1060 -1863 0 cellNo=84
rlabel pdiffusion 1067 -1863 1067 -1863 0 cellNo=242
rlabel pdiffusion 1074 -1863 1074 -1863 0 feedthrough
rlabel pdiffusion 1081 -1863 1081 -1863 0 feedthrough
rlabel pdiffusion 1088 -1863 1088 -1863 0 feedthrough
rlabel pdiffusion 1095 -1863 1095 -1863 0 feedthrough
rlabel pdiffusion 1102 -1863 1102 -1863 0 feedthrough
rlabel pdiffusion 1109 -1863 1109 -1863 0 feedthrough
rlabel pdiffusion 1116 -1863 1116 -1863 0 feedthrough
rlabel pdiffusion 1123 -1863 1123 -1863 0 feedthrough
rlabel pdiffusion 1130 -1863 1130 -1863 0 feedthrough
rlabel pdiffusion 1137 -1863 1137 -1863 0 feedthrough
rlabel pdiffusion 1144 -1863 1144 -1863 0 feedthrough
rlabel pdiffusion 1151 -1863 1151 -1863 0 feedthrough
rlabel pdiffusion 1158 -1863 1158 -1863 0 feedthrough
rlabel pdiffusion 1165 -1863 1165 -1863 0 feedthrough
rlabel pdiffusion 1172 -1863 1172 -1863 0 feedthrough
rlabel pdiffusion 1179 -1863 1179 -1863 0 feedthrough
rlabel pdiffusion 1186 -1863 1186 -1863 0 feedthrough
rlabel pdiffusion 1193 -1863 1193 -1863 0 feedthrough
rlabel pdiffusion 1200 -1863 1200 -1863 0 feedthrough
rlabel pdiffusion 1207 -1863 1207 -1863 0 feedthrough
rlabel pdiffusion 1214 -1863 1214 -1863 0 feedthrough
rlabel pdiffusion 1221 -1863 1221 -1863 0 feedthrough
rlabel pdiffusion 1228 -1863 1228 -1863 0 feedthrough
rlabel pdiffusion 1235 -1863 1235 -1863 0 feedthrough
rlabel pdiffusion 1242 -1863 1242 -1863 0 feedthrough
rlabel pdiffusion 1249 -1863 1249 -1863 0 feedthrough
rlabel pdiffusion 1256 -1863 1256 -1863 0 feedthrough
rlabel pdiffusion 1263 -1863 1263 -1863 0 feedthrough
rlabel pdiffusion 1270 -1863 1270 -1863 0 feedthrough
rlabel pdiffusion 1277 -1863 1277 -1863 0 feedthrough
rlabel pdiffusion 1284 -1863 1284 -1863 0 feedthrough
rlabel pdiffusion 1291 -1863 1291 -1863 0 feedthrough
rlabel pdiffusion 1298 -1863 1298 -1863 0 feedthrough
rlabel pdiffusion 1305 -1863 1305 -1863 0 feedthrough
rlabel pdiffusion 1312 -1863 1312 -1863 0 feedthrough
rlabel pdiffusion 1319 -1863 1319 -1863 0 feedthrough
rlabel pdiffusion 1326 -1863 1326 -1863 0 feedthrough
rlabel pdiffusion 1333 -1863 1333 -1863 0 feedthrough
rlabel pdiffusion 1340 -1863 1340 -1863 0 feedthrough
rlabel pdiffusion 1347 -1863 1347 -1863 0 feedthrough
rlabel pdiffusion 1354 -1863 1354 -1863 0 feedthrough
rlabel pdiffusion 1361 -1863 1361 -1863 0 feedthrough
rlabel pdiffusion 1368 -1863 1368 -1863 0 feedthrough
rlabel pdiffusion 1375 -1863 1375 -1863 0 feedthrough
rlabel pdiffusion 1382 -1863 1382 -1863 0 feedthrough
rlabel pdiffusion 1389 -1863 1389 -1863 0 feedthrough
rlabel pdiffusion 1396 -1863 1396 -1863 0 cellNo=163
rlabel pdiffusion 1403 -1863 1403 -1863 0 feedthrough
rlabel pdiffusion 1410 -1863 1410 -1863 0 feedthrough
rlabel pdiffusion 1417 -1863 1417 -1863 0 feedthrough
rlabel pdiffusion 1424 -1863 1424 -1863 0 feedthrough
rlabel pdiffusion 1431 -1863 1431 -1863 0 feedthrough
rlabel pdiffusion 3 -1990 3 -1990 0 feedthrough
rlabel pdiffusion 10 -1990 10 -1990 0 feedthrough
rlabel pdiffusion 17 -1990 17 -1990 0 feedthrough
rlabel pdiffusion 24 -1990 24 -1990 0 cellNo=255
rlabel pdiffusion 31 -1990 31 -1990 0 feedthrough
rlabel pdiffusion 38 -1990 38 -1990 0 cellNo=493
rlabel pdiffusion 45 -1990 45 -1990 0 feedthrough
rlabel pdiffusion 52 -1990 52 -1990 0 feedthrough
rlabel pdiffusion 59 -1990 59 -1990 0 feedthrough
rlabel pdiffusion 66 -1990 66 -1990 0 cellNo=537
rlabel pdiffusion 73 -1990 73 -1990 0 cellNo=436
rlabel pdiffusion 80 -1990 80 -1990 0 feedthrough
rlabel pdiffusion 87 -1990 87 -1990 0 feedthrough
rlabel pdiffusion 94 -1990 94 -1990 0 feedthrough
rlabel pdiffusion 101 -1990 101 -1990 0 feedthrough
rlabel pdiffusion 108 -1990 108 -1990 0 feedthrough
rlabel pdiffusion 115 -1990 115 -1990 0 feedthrough
rlabel pdiffusion 122 -1990 122 -1990 0 feedthrough
rlabel pdiffusion 129 -1990 129 -1990 0 feedthrough
rlabel pdiffusion 136 -1990 136 -1990 0 feedthrough
rlabel pdiffusion 143 -1990 143 -1990 0 feedthrough
rlabel pdiffusion 150 -1990 150 -1990 0 feedthrough
rlabel pdiffusion 157 -1990 157 -1990 0 feedthrough
rlabel pdiffusion 164 -1990 164 -1990 0 feedthrough
rlabel pdiffusion 171 -1990 171 -1990 0 cellNo=30
rlabel pdiffusion 178 -1990 178 -1990 0 feedthrough
rlabel pdiffusion 185 -1990 185 -1990 0 feedthrough
rlabel pdiffusion 192 -1990 192 -1990 0 feedthrough
rlabel pdiffusion 199 -1990 199 -1990 0 feedthrough
rlabel pdiffusion 206 -1990 206 -1990 0 feedthrough
rlabel pdiffusion 213 -1990 213 -1990 0 feedthrough
rlabel pdiffusion 220 -1990 220 -1990 0 feedthrough
rlabel pdiffusion 227 -1990 227 -1990 0 cellNo=433
rlabel pdiffusion 234 -1990 234 -1990 0 feedthrough
rlabel pdiffusion 241 -1990 241 -1990 0 feedthrough
rlabel pdiffusion 248 -1990 248 -1990 0 feedthrough
rlabel pdiffusion 255 -1990 255 -1990 0 feedthrough
rlabel pdiffusion 262 -1990 262 -1990 0 feedthrough
rlabel pdiffusion 269 -1990 269 -1990 0 feedthrough
rlabel pdiffusion 276 -1990 276 -1990 0 feedthrough
rlabel pdiffusion 283 -1990 283 -1990 0 feedthrough
rlabel pdiffusion 290 -1990 290 -1990 0 feedthrough
rlabel pdiffusion 297 -1990 297 -1990 0 feedthrough
rlabel pdiffusion 304 -1990 304 -1990 0 feedthrough
rlabel pdiffusion 311 -1990 311 -1990 0 feedthrough
rlabel pdiffusion 318 -1990 318 -1990 0 feedthrough
rlabel pdiffusion 325 -1990 325 -1990 0 feedthrough
rlabel pdiffusion 332 -1990 332 -1990 0 feedthrough
rlabel pdiffusion 339 -1990 339 -1990 0 feedthrough
rlabel pdiffusion 346 -1990 346 -1990 0 feedthrough
rlabel pdiffusion 353 -1990 353 -1990 0 cellNo=61
rlabel pdiffusion 360 -1990 360 -1990 0 feedthrough
rlabel pdiffusion 367 -1990 367 -1990 0 feedthrough
rlabel pdiffusion 374 -1990 374 -1990 0 cellNo=345
rlabel pdiffusion 381 -1990 381 -1990 0 feedthrough
rlabel pdiffusion 388 -1990 388 -1990 0 feedthrough
rlabel pdiffusion 395 -1990 395 -1990 0 feedthrough
rlabel pdiffusion 402 -1990 402 -1990 0 feedthrough
rlabel pdiffusion 409 -1990 409 -1990 0 cellNo=476
rlabel pdiffusion 416 -1990 416 -1990 0 feedthrough
rlabel pdiffusion 423 -1990 423 -1990 0 feedthrough
rlabel pdiffusion 430 -1990 430 -1990 0 feedthrough
rlabel pdiffusion 437 -1990 437 -1990 0 feedthrough
rlabel pdiffusion 444 -1990 444 -1990 0 feedthrough
rlabel pdiffusion 451 -1990 451 -1990 0 feedthrough
rlabel pdiffusion 458 -1990 458 -1990 0 feedthrough
rlabel pdiffusion 465 -1990 465 -1990 0 feedthrough
rlabel pdiffusion 472 -1990 472 -1990 0 feedthrough
rlabel pdiffusion 479 -1990 479 -1990 0 feedthrough
rlabel pdiffusion 486 -1990 486 -1990 0 feedthrough
rlabel pdiffusion 493 -1990 493 -1990 0 feedthrough
rlabel pdiffusion 500 -1990 500 -1990 0 feedthrough
rlabel pdiffusion 507 -1990 507 -1990 0 cellNo=300
rlabel pdiffusion 514 -1990 514 -1990 0 cellNo=587
rlabel pdiffusion 521 -1990 521 -1990 0 cellNo=556
rlabel pdiffusion 528 -1990 528 -1990 0 feedthrough
rlabel pdiffusion 535 -1990 535 -1990 0 feedthrough
rlabel pdiffusion 542 -1990 542 -1990 0 feedthrough
rlabel pdiffusion 549 -1990 549 -1990 0 feedthrough
rlabel pdiffusion 556 -1990 556 -1990 0 feedthrough
rlabel pdiffusion 563 -1990 563 -1990 0 cellNo=478
rlabel pdiffusion 570 -1990 570 -1990 0 feedthrough
rlabel pdiffusion 577 -1990 577 -1990 0 cellNo=586
rlabel pdiffusion 584 -1990 584 -1990 0 cellNo=573
rlabel pdiffusion 591 -1990 591 -1990 0 feedthrough
rlabel pdiffusion 598 -1990 598 -1990 0 feedthrough
rlabel pdiffusion 605 -1990 605 -1990 0 feedthrough
rlabel pdiffusion 612 -1990 612 -1990 0 cellNo=36
rlabel pdiffusion 619 -1990 619 -1990 0 feedthrough
rlabel pdiffusion 626 -1990 626 -1990 0 feedthrough
rlabel pdiffusion 633 -1990 633 -1990 0 feedthrough
rlabel pdiffusion 640 -1990 640 -1990 0 cellNo=398
rlabel pdiffusion 647 -1990 647 -1990 0 feedthrough
rlabel pdiffusion 654 -1990 654 -1990 0 feedthrough
rlabel pdiffusion 661 -1990 661 -1990 0 cellNo=464
rlabel pdiffusion 668 -1990 668 -1990 0 feedthrough
rlabel pdiffusion 675 -1990 675 -1990 0 feedthrough
rlabel pdiffusion 682 -1990 682 -1990 0 feedthrough
rlabel pdiffusion 689 -1990 689 -1990 0 feedthrough
rlabel pdiffusion 696 -1990 696 -1990 0 feedthrough
rlabel pdiffusion 703 -1990 703 -1990 0 cellNo=2
rlabel pdiffusion 710 -1990 710 -1990 0 feedthrough
rlabel pdiffusion 717 -1990 717 -1990 0 feedthrough
rlabel pdiffusion 724 -1990 724 -1990 0 cellNo=194
rlabel pdiffusion 731 -1990 731 -1990 0 feedthrough
rlabel pdiffusion 738 -1990 738 -1990 0 feedthrough
rlabel pdiffusion 745 -1990 745 -1990 0 feedthrough
rlabel pdiffusion 752 -1990 752 -1990 0 cellNo=232
rlabel pdiffusion 759 -1990 759 -1990 0 feedthrough
rlabel pdiffusion 766 -1990 766 -1990 0 feedthrough
rlabel pdiffusion 773 -1990 773 -1990 0 feedthrough
rlabel pdiffusion 780 -1990 780 -1990 0 cellNo=358
rlabel pdiffusion 787 -1990 787 -1990 0 feedthrough
rlabel pdiffusion 794 -1990 794 -1990 0 feedthrough
rlabel pdiffusion 801 -1990 801 -1990 0 feedthrough
rlabel pdiffusion 808 -1990 808 -1990 0 cellNo=517
rlabel pdiffusion 815 -1990 815 -1990 0 feedthrough
rlabel pdiffusion 822 -1990 822 -1990 0 feedthrough
rlabel pdiffusion 829 -1990 829 -1990 0 feedthrough
rlabel pdiffusion 836 -1990 836 -1990 0 feedthrough
rlabel pdiffusion 843 -1990 843 -1990 0 feedthrough
rlabel pdiffusion 850 -1990 850 -1990 0 cellNo=372
rlabel pdiffusion 857 -1990 857 -1990 0 feedthrough
rlabel pdiffusion 864 -1990 864 -1990 0 feedthrough
rlabel pdiffusion 871 -1990 871 -1990 0 feedthrough
rlabel pdiffusion 878 -1990 878 -1990 0 feedthrough
rlabel pdiffusion 885 -1990 885 -1990 0 feedthrough
rlabel pdiffusion 892 -1990 892 -1990 0 feedthrough
rlabel pdiffusion 899 -1990 899 -1990 0 feedthrough
rlabel pdiffusion 906 -1990 906 -1990 0 feedthrough
rlabel pdiffusion 913 -1990 913 -1990 0 feedthrough
rlabel pdiffusion 920 -1990 920 -1990 0 feedthrough
rlabel pdiffusion 927 -1990 927 -1990 0 feedthrough
rlabel pdiffusion 934 -1990 934 -1990 0 feedthrough
rlabel pdiffusion 941 -1990 941 -1990 0 feedthrough
rlabel pdiffusion 948 -1990 948 -1990 0 cellNo=475
rlabel pdiffusion 955 -1990 955 -1990 0 feedthrough
rlabel pdiffusion 962 -1990 962 -1990 0 feedthrough
rlabel pdiffusion 969 -1990 969 -1990 0 feedthrough
rlabel pdiffusion 976 -1990 976 -1990 0 feedthrough
rlabel pdiffusion 983 -1990 983 -1990 0 feedthrough
rlabel pdiffusion 990 -1990 990 -1990 0 feedthrough
rlabel pdiffusion 997 -1990 997 -1990 0 feedthrough
rlabel pdiffusion 1004 -1990 1004 -1990 0 feedthrough
rlabel pdiffusion 1011 -1990 1011 -1990 0 feedthrough
rlabel pdiffusion 1018 -1990 1018 -1990 0 feedthrough
rlabel pdiffusion 1025 -1990 1025 -1990 0 feedthrough
rlabel pdiffusion 1032 -1990 1032 -1990 0 feedthrough
rlabel pdiffusion 1039 -1990 1039 -1990 0 feedthrough
rlabel pdiffusion 1046 -1990 1046 -1990 0 feedthrough
rlabel pdiffusion 1053 -1990 1053 -1990 0 feedthrough
rlabel pdiffusion 1060 -1990 1060 -1990 0 feedthrough
rlabel pdiffusion 1067 -1990 1067 -1990 0 feedthrough
rlabel pdiffusion 1074 -1990 1074 -1990 0 feedthrough
rlabel pdiffusion 1081 -1990 1081 -1990 0 feedthrough
rlabel pdiffusion 1088 -1990 1088 -1990 0 feedthrough
rlabel pdiffusion 1095 -1990 1095 -1990 0 feedthrough
rlabel pdiffusion 1102 -1990 1102 -1990 0 feedthrough
rlabel pdiffusion 1109 -1990 1109 -1990 0 feedthrough
rlabel pdiffusion 1116 -1990 1116 -1990 0 feedthrough
rlabel pdiffusion 1123 -1990 1123 -1990 0 feedthrough
rlabel pdiffusion 1130 -1990 1130 -1990 0 feedthrough
rlabel pdiffusion 1137 -1990 1137 -1990 0 feedthrough
rlabel pdiffusion 1144 -1990 1144 -1990 0 feedthrough
rlabel pdiffusion 1151 -1990 1151 -1990 0 feedthrough
rlabel pdiffusion 1158 -1990 1158 -1990 0 feedthrough
rlabel pdiffusion 1165 -1990 1165 -1990 0 feedthrough
rlabel pdiffusion 1172 -1990 1172 -1990 0 feedthrough
rlabel pdiffusion 1179 -1990 1179 -1990 0 feedthrough
rlabel pdiffusion 1186 -1990 1186 -1990 0 feedthrough
rlabel pdiffusion 1193 -1990 1193 -1990 0 feedthrough
rlabel pdiffusion 1200 -1990 1200 -1990 0 feedthrough
rlabel pdiffusion 1207 -1990 1207 -1990 0 feedthrough
rlabel pdiffusion 1214 -1990 1214 -1990 0 feedthrough
rlabel pdiffusion 1221 -1990 1221 -1990 0 feedthrough
rlabel pdiffusion 1228 -1990 1228 -1990 0 feedthrough
rlabel pdiffusion 1235 -1990 1235 -1990 0 feedthrough
rlabel pdiffusion 1242 -1990 1242 -1990 0 feedthrough
rlabel pdiffusion 1249 -1990 1249 -1990 0 feedthrough
rlabel pdiffusion 1256 -1990 1256 -1990 0 feedthrough
rlabel pdiffusion 1263 -1990 1263 -1990 0 feedthrough
rlabel pdiffusion 1270 -1990 1270 -1990 0 feedthrough
rlabel pdiffusion 1277 -1990 1277 -1990 0 feedthrough
rlabel pdiffusion 1284 -1990 1284 -1990 0 feedthrough
rlabel pdiffusion 1291 -1990 1291 -1990 0 feedthrough
rlabel pdiffusion 1298 -1990 1298 -1990 0 feedthrough
rlabel pdiffusion 1305 -1990 1305 -1990 0 feedthrough
rlabel pdiffusion 1312 -1990 1312 -1990 0 feedthrough
rlabel pdiffusion 1319 -1990 1319 -1990 0 feedthrough
rlabel pdiffusion 1326 -1990 1326 -1990 0 feedthrough
rlabel pdiffusion 1333 -1990 1333 -1990 0 feedthrough
rlabel pdiffusion 1340 -1990 1340 -1990 0 feedthrough
rlabel pdiffusion 1347 -1990 1347 -1990 0 feedthrough
rlabel pdiffusion 1354 -1990 1354 -1990 0 feedthrough
rlabel pdiffusion 1361 -1990 1361 -1990 0 feedthrough
rlabel pdiffusion 1368 -1990 1368 -1990 0 feedthrough
rlabel pdiffusion 1375 -1990 1375 -1990 0 feedthrough
rlabel pdiffusion 1382 -1990 1382 -1990 0 feedthrough
rlabel pdiffusion 1389 -1990 1389 -1990 0 feedthrough
rlabel pdiffusion 1396 -1990 1396 -1990 0 feedthrough
rlabel pdiffusion 1403 -1990 1403 -1990 0 feedthrough
rlabel pdiffusion 3 -2109 3 -2109 0 cellNo=361
rlabel pdiffusion 10 -2109 10 -2109 0 cellNo=129
rlabel pdiffusion 17 -2109 17 -2109 0 feedthrough
rlabel pdiffusion 24 -2109 24 -2109 0 feedthrough
rlabel pdiffusion 31 -2109 31 -2109 0 feedthrough
rlabel pdiffusion 38 -2109 38 -2109 0 feedthrough
rlabel pdiffusion 45 -2109 45 -2109 0 feedthrough
rlabel pdiffusion 52 -2109 52 -2109 0 feedthrough
rlabel pdiffusion 59 -2109 59 -2109 0 feedthrough
rlabel pdiffusion 66 -2109 66 -2109 0 feedthrough
rlabel pdiffusion 73 -2109 73 -2109 0 feedthrough
rlabel pdiffusion 80 -2109 80 -2109 0 feedthrough
rlabel pdiffusion 87 -2109 87 -2109 0 feedthrough
rlabel pdiffusion 94 -2109 94 -2109 0 cellNo=147
rlabel pdiffusion 101 -2109 101 -2109 0 feedthrough
rlabel pdiffusion 108 -2109 108 -2109 0 cellNo=127
rlabel pdiffusion 115 -2109 115 -2109 0 feedthrough
rlabel pdiffusion 122 -2109 122 -2109 0 feedthrough
rlabel pdiffusion 129 -2109 129 -2109 0 cellNo=509
rlabel pdiffusion 136 -2109 136 -2109 0 feedthrough
rlabel pdiffusion 143 -2109 143 -2109 0 feedthrough
rlabel pdiffusion 150 -2109 150 -2109 0 feedthrough
rlabel pdiffusion 157 -2109 157 -2109 0 feedthrough
rlabel pdiffusion 164 -2109 164 -2109 0 cellNo=364
rlabel pdiffusion 171 -2109 171 -2109 0 cellNo=529
rlabel pdiffusion 178 -2109 178 -2109 0 feedthrough
rlabel pdiffusion 185 -2109 185 -2109 0 feedthrough
rlabel pdiffusion 192 -2109 192 -2109 0 feedthrough
rlabel pdiffusion 199 -2109 199 -2109 0 feedthrough
rlabel pdiffusion 206 -2109 206 -2109 0 feedthrough
rlabel pdiffusion 213 -2109 213 -2109 0 feedthrough
rlabel pdiffusion 220 -2109 220 -2109 0 feedthrough
rlabel pdiffusion 227 -2109 227 -2109 0 feedthrough
rlabel pdiffusion 234 -2109 234 -2109 0 feedthrough
rlabel pdiffusion 241 -2109 241 -2109 0 feedthrough
rlabel pdiffusion 248 -2109 248 -2109 0 feedthrough
rlabel pdiffusion 255 -2109 255 -2109 0 feedthrough
rlabel pdiffusion 262 -2109 262 -2109 0 feedthrough
rlabel pdiffusion 269 -2109 269 -2109 0 feedthrough
rlabel pdiffusion 276 -2109 276 -2109 0 feedthrough
rlabel pdiffusion 283 -2109 283 -2109 0 feedthrough
rlabel pdiffusion 290 -2109 290 -2109 0 feedthrough
rlabel pdiffusion 297 -2109 297 -2109 0 feedthrough
rlabel pdiffusion 304 -2109 304 -2109 0 feedthrough
rlabel pdiffusion 311 -2109 311 -2109 0 feedthrough
rlabel pdiffusion 318 -2109 318 -2109 0 cellNo=555
rlabel pdiffusion 325 -2109 325 -2109 0 feedthrough
rlabel pdiffusion 332 -2109 332 -2109 0 cellNo=594
rlabel pdiffusion 339 -2109 339 -2109 0 feedthrough
rlabel pdiffusion 346 -2109 346 -2109 0 cellNo=294
rlabel pdiffusion 353 -2109 353 -2109 0 feedthrough
rlabel pdiffusion 360 -2109 360 -2109 0 feedthrough
rlabel pdiffusion 367 -2109 367 -2109 0 feedthrough
rlabel pdiffusion 374 -2109 374 -2109 0 feedthrough
rlabel pdiffusion 381 -2109 381 -2109 0 feedthrough
rlabel pdiffusion 388 -2109 388 -2109 0 feedthrough
rlabel pdiffusion 395 -2109 395 -2109 0 feedthrough
rlabel pdiffusion 402 -2109 402 -2109 0 feedthrough
rlabel pdiffusion 409 -2109 409 -2109 0 feedthrough
rlabel pdiffusion 416 -2109 416 -2109 0 feedthrough
rlabel pdiffusion 423 -2109 423 -2109 0 feedthrough
rlabel pdiffusion 430 -2109 430 -2109 0 feedthrough
rlabel pdiffusion 437 -2109 437 -2109 0 feedthrough
rlabel pdiffusion 444 -2109 444 -2109 0 feedthrough
rlabel pdiffusion 451 -2109 451 -2109 0 cellNo=324
rlabel pdiffusion 458 -2109 458 -2109 0 feedthrough
rlabel pdiffusion 465 -2109 465 -2109 0 feedthrough
rlabel pdiffusion 472 -2109 472 -2109 0 feedthrough
rlabel pdiffusion 479 -2109 479 -2109 0 feedthrough
rlabel pdiffusion 486 -2109 486 -2109 0 cellNo=352
rlabel pdiffusion 493 -2109 493 -2109 0 feedthrough
rlabel pdiffusion 500 -2109 500 -2109 0 cellNo=572
rlabel pdiffusion 507 -2109 507 -2109 0 feedthrough
rlabel pdiffusion 514 -2109 514 -2109 0 feedthrough
rlabel pdiffusion 521 -2109 521 -2109 0 feedthrough
rlabel pdiffusion 528 -2109 528 -2109 0 feedthrough
rlabel pdiffusion 535 -2109 535 -2109 0 feedthrough
rlabel pdiffusion 542 -2109 542 -2109 0 feedthrough
rlabel pdiffusion 549 -2109 549 -2109 0 feedthrough
rlabel pdiffusion 556 -2109 556 -2109 0 feedthrough
rlabel pdiffusion 563 -2109 563 -2109 0 feedthrough
rlabel pdiffusion 570 -2109 570 -2109 0 feedthrough
rlabel pdiffusion 577 -2109 577 -2109 0 cellNo=543
rlabel pdiffusion 584 -2109 584 -2109 0 feedthrough
rlabel pdiffusion 591 -2109 591 -2109 0 feedthrough
rlabel pdiffusion 598 -2109 598 -2109 0 feedthrough
rlabel pdiffusion 605 -2109 605 -2109 0 feedthrough
rlabel pdiffusion 612 -2109 612 -2109 0 feedthrough
rlabel pdiffusion 619 -2109 619 -2109 0 cellNo=290
rlabel pdiffusion 626 -2109 626 -2109 0 feedthrough
rlabel pdiffusion 633 -2109 633 -2109 0 feedthrough
rlabel pdiffusion 640 -2109 640 -2109 0 feedthrough
rlabel pdiffusion 647 -2109 647 -2109 0 feedthrough
rlabel pdiffusion 654 -2109 654 -2109 0 feedthrough
rlabel pdiffusion 661 -2109 661 -2109 0 feedthrough
rlabel pdiffusion 668 -2109 668 -2109 0 cellNo=115
rlabel pdiffusion 675 -2109 675 -2109 0 feedthrough
rlabel pdiffusion 682 -2109 682 -2109 0 feedthrough
rlabel pdiffusion 689 -2109 689 -2109 0 cellNo=213
rlabel pdiffusion 696 -2109 696 -2109 0 feedthrough
rlabel pdiffusion 703 -2109 703 -2109 0 feedthrough
rlabel pdiffusion 710 -2109 710 -2109 0 feedthrough
rlabel pdiffusion 717 -2109 717 -2109 0 feedthrough
rlabel pdiffusion 724 -2109 724 -2109 0 feedthrough
rlabel pdiffusion 731 -2109 731 -2109 0 feedthrough
rlabel pdiffusion 738 -2109 738 -2109 0 feedthrough
rlabel pdiffusion 745 -2109 745 -2109 0 feedthrough
rlabel pdiffusion 752 -2109 752 -2109 0 feedthrough
rlabel pdiffusion 759 -2109 759 -2109 0 feedthrough
rlabel pdiffusion 766 -2109 766 -2109 0 feedthrough
rlabel pdiffusion 773 -2109 773 -2109 0 feedthrough
rlabel pdiffusion 780 -2109 780 -2109 0 cellNo=133
rlabel pdiffusion 787 -2109 787 -2109 0 feedthrough
rlabel pdiffusion 794 -2109 794 -2109 0 feedthrough
rlabel pdiffusion 801 -2109 801 -2109 0 feedthrough
rlabel pdiffusion 808 -2109 808 -2109 0 feedthrough
rlabel pdiffusion 815 -2109 815 -2109 0 cellNo=441
rlabel pdiffusion 822 -2109 822 -2109 0 cellNo=81
rlabel pdiffusion 829 -2109 829 -2109 0 feedthrough
rlabel pdiffusion 836 -2109 836 -2109 0 feedthrough
rlabel pdiffusion 843 -2109 843 -2109 0 feedthrough
rlabel pdiffusion 850 -2109 850 -2109 0 feedthrough
rlabel pdiffusion 857 -2109 857 -2109 0 feedthrough
rlabel pdiffusion 864 -2109 864 -2109 0 feedthrough
rlabel pdiffusion 871 -2109 871 -2109 0 feedthrough
rlabel pdiffusion 878 -2109 878 -2109 0 feedthrough
rlabel pdiffusion 885 -2109 885 -2109 0 feedthrough
rlabel pdiffusion 892 -2109 892 -2109 0 cellNo=293
rlabel pdiffusion 899 -2109 899 -2109 0 feedthrough
rlabel pdiffusion 906 -2109 906 -2109 0 feedthrough
rlabel pdiffusion 913 -2109 913 -2109 0 feedthrough
rlabel pdiffusion 920 -2109 920 -2109 0 feedthrough
rlabel pdiffusion 927 -2109 927 -2109 0 feedthrough
rlabel pdiffusion 934 -2109 934 -2109 0 feedthrough
rlabel pdiffusion 941 -2109 941 -2109 0 feedthrough
rlabel pdiffusion 948 -2109 948 -2109 0 feedthrough
rlabel pdiffusion 955 -2109 955 -2109 0 feedthrough
rlabel pdiffusion 962 -2109 962 -2109 0 feedthrough
rlabel pdiffusion 969 -2109 969 -2109 0 cellNo=593
rlabel pdiffusion 976 -2109 976 -2109 0 feedthrough
rlabel pdiffusion 983 -2109 983 -2109 0 feedthrough
rlabel pdiffusion 990 -2109 990 -2109 0 cellNo=208
rlabel pdiffusion 997 -2109 997 -2109 0 feedthrough
rlabel pdiffusion 1004 -2109 1004 -2109 0 feedthrough
rlabel pdiffusion 1011 -2109 1011 -2109 0 feedthrough
rlabel pdiffusion 1018 -2109 1018 -2109 0 feedthrough
rlabel pdiffusion 1025 -2109 1025 -2109 0 feedthrough
rlabel pdiffusion 1032 -2109 1032 -2109 0 feedthrough
rlabel pdiffusion 1039 -2109 1039 -2109 0 feedthrough
rlabel pdiffusion 1046 -2109 1046 -2109 0 feedthrough
rlabel pdiffusion 1053 -2109 1053 -2109 0 feedthrough
rlabel pdiffusion 1060 -2109 1060 -2109 0 feedthrough
rlabel pdiffusion 1067 -2109 1067 -2109 0 feedthrough
rlabel pdiffusion 1074 -2109 1074 -2109 0 feedthrough
rlabel pdiffusion 1081 -2109 1081 -2109 0 feedthrough
rlabel pdiffusion 1088 -2109 1088 -2109 0 feedthrough
rlabel pdiffusion 1095 -2109 1095 -2109 0 feedthrough
rlabel pdiffusion 1102 -2109 1102 -2109 0 feedthrough
rlabel pdiffusion 1109 -2109 1109 -2109 0 feedthrough
rlabel pdiffusion 1116 -2109 1116 -2109 0 cellNo=351
rlabel pdiffusion 1123 -2109 1123 -2109 0 feedthrough
rlabel pdiffusion 1130 -2109 1130 -2109 0 feedthrough
rlabel pdiffusion 1137 -2109 1137 -2109 0 cellNo=80
rlabel pdiffusion 1144 -2109 1144 -2109 0 feedthrough
rlabel pdiffusion 1151 -2109 1151 -2109 0 feedthrough
rlabel pdiffusion 1158 -2109 1158 -2109 0 feedthrough
rlabel pdiffusion 1165 -2109 1165 -2109 0 feedthrough
rlabel pdiffusion 1172 -2109 1172 -2109 0 feedthrough
rlabel pdiffusion 1179 -2109 1179 -2109 0 feedthrough
rlabel pdiffusion 1186 -2109 1186 -2109 0 feedthrough
rlabel pdiffusion 1193 -2109 1193 -2109 0 feedthrough
rlabel pdiffusion 1200 -2109 1200 -2109 0 feedthrough
rlabel pdiffusion 1207 -2109 1207 -2109 0 feedthrough
rlabel pdiffusion 1214 -2109 1214 -2109 0 feedthrough
rlabel pdiffusion 1221 -2109 1221 -2109 0 feedthrough
rlabel pdiffusion 1228 -2109 1228 -2109 0 feedthrough
rlabel pdiffusion 1235 -2109 1235 -2109 0 feedthrough
rlabel pdiffusion 1242 -2109 1242 -2109 0 feedthrough
rlabel pdiffusion 1249 -2109 1249 -2109 0 feedthrough
rlabel pdiffusion 1256 -2109 1256 -2109 0 feedthrough
rlabel pdiffusion 1263 -2109 1263 -2109 0 feedthrough
rlabel pdiffusion 1270 -2109 1270 -2109 0 feedthrough
rlabel pdiffusion 1277 -2109 1277 -2109 0 feedthrough
rlabel pdiffusion 1284 -2109 1284 -2109 0 feedthrough
rlabel pdiffusion 1291 -2109 1291 -2109 0 feedthrough
rlabel pdiffusion 1298 -2109 1298 -2109 0 feedthrough
rlabel pdiffusion 1305 -2109 1305 -2109 0 feedthrough
rlabel pdiffusion 1312 -2109 1312 -2109 0 feedthrough
rlabel pdiffusion 1319 -2109 1319 -2109 0 feedthrough
rlabel pdiffusion 1326 -2109 1326 -2109 0 feedthrough
rlabel pdiffusion 3 -2242 3 -2242 0 feedthrough
rlabel pdiffusion 10 -2242 10 -2242 0 feedthrough
rlabel pdiffusion 17 -2242 17 -2242 0 feedthrough
rlabel pdiffusion 24 -2242 24 -2242 0 cellNo=353
rlabel pdiffusion 31 -2242 31 -2242 0 cellNo=580
rlabel pdiffusion 38 -2242 38 -2242 0 cellNo=257
rlabel pdiffusion 45 -2242 45 -2242 0 feedthrough
rlabel pdiffusion 52 -2242 52 -2242 0 feedthrough
rlabel pdiffusion 59 -2242 59 -2242 0 feedthrough
rlabel pdiffusion 66 -2242 66 -2242 0 feedthrough
rlabel pdiffusion 73 -2242 73 -2242 0 cellNo=501
rlabel pdiffusion 80 -2242 80 -2242 0 feedthrough
rlabel pdiffusion 87 -2242 87 -2242 0 feedthrough
rlabel pdiffusion 94 -2242 94 -2242 0 feedthrough
rlabel pdiffusion 101 -2242 101 -2242 0 feedthrough
rlabel pdiffusion 108 -2242 108 -2242 0 feedthrough
rlabel pdiffusion 115 -2242 115 -2242 0 cellNo=321
rlabel pdiffusion 122 -2242 122 -2242 0 feedthrough
rlabel pdiffusion 129 -2242 129 -2242 0 feedthrough
rlabel pdiffusion 136 -2242 136 -2242 0 cellNo=569
rlabel pdiffusion 143 -2242 143 -2242 0 feedthrough
rlabel pdiffusion 150 -2242 150 -2242 0 cellNo=378
rlabel pdiffusion 157 -2242 157 -2242 0 feedthrough
rlabel pdiffusion 164 -2242 164 -2242 0 feedthrough
rlabel pdiffusion 171 -2242 171 -2242 0 feedthrough
rlabel pdiffusion 178 -2242 178 -2242 0 feedthrough
rlabel pdiffusion 185 -2242 185 -2242 0 feedthrough
rlabel pdiffusion 192 -2242 192 -2242 0 feedthrough
rlabel pdiffusion 199 -2242 199 -2242 0 feedthrough
rlabel pdiffusion 206 -2242 206 -2242 0 feedthrough
rlabel pdiffusion 213 -2242 213 -2242 0 feedthrough
rlabel pdiffusion 220 -2242 220 -2242 0 feedthrough
rlabel pdiffusion 227 -2242 227 -2242 0 feedthrough
rlabel pdiffusion 234 -2242 234 -2242 0 feedthrough
rlabel pdiffusion 241 -2242 241 -2242 0 feedthrough
rlabel pdiffusion 248 -2242 248 -2242 0 feedthrough
rlabel pdiffusion 255 -2242 255 -2242 0 feedthrough
rlabel pdiffusion 262 -2242 262 -2242 0 feedthrough
rlabel pdiffusion 269 -2242 269 -2242 0 feedthrough
rlabel pdiffusion 276 -2242 276 -2242 0 feedthrough
rlabel pdiffusion 283 -2242 283 -2242 0 feedthrough
rlabel pdiffusion 290 -2242 290 -2242 0 feedthrough
rlabel pdiffusion 297 -2242 297 -2242 0 cellNo=549
rlabel pdiffusion 304 -2242 304 -2242 0 feedthrough
rlabel pdiffusion 311 -2242 311 -2242 0 feedthrough
rlabel pdiffusion 318 -2242 318 -2242 0 feedthrough
rlabel pdiffusion 325 -2242 325 -2242 0 feedthrough
rlabel pdiffusion 332 -2242 332 -2242 0 feedthrough
rlabel pdiffusion 339 -2242 339 -2242 0 cellNo=384
rlabel pdiffusion 346 -2242 346 -2242 0 feedthrough
rlabel pdiffusion 353 -2242 353 -2242 0 feedthrough
rlabel pdiffusion 360 -2242 360 -2242 0 feedthrough
rlabel pdiffusion 367 -2242 367 -2242 0 feedthrough
rlabel pdiffusion 374 -2242 374 -2242 0 feedthrough
rlabel pdiffusion 381 -2242 381 -2242 0 feedthrough
rlabel pdiffusion 388 -2242 388 -2242 0 feedthrough
rlabel pdiffusion 395 -2242 395 -2242 0 cellNo=420
rlabel pdiffusion 402 -2242 402 -2242 0 cellNo=313
rlabel pdiffusion 409 -2242 409 -2242 0 cellNo=17
rlabel pdiffusion 416 -2242 416 -2242 0 feedthrough
rlabel pdiffusion 423 -2242 423 -2242 0 cellNo=512
rlabel pdiffusion 430 -2242 430 -2242 0 feedthrough
rlabel pdiffusion 437 -2242 437 -2242 0 feedthrough
rlabel pdiffusion 444 -2242 444 -2242 0 feedthrough
rlabel pdiffusion 451 -2242 451 -2242 0 cellNo=570
rlabel pdiffusion 458 -2242 458 -2242 0 feedthrough
rlabel pdiffusion 465 -2242 465 -2242 0 feedthrough
rlabel pdiffusion 472 -2242 472 -2242 0 feedthrough
rlabel pdiffusion 479 -2242 479 -2242 0 feedthrough
rlabel pdiffusion 486 -2242 486 -2242 0 feedthrough
rlabel pdiffusion 493 -2242 493 -2242 0 feedthrough
rlabel pdiffusion 500 -2242 500 -2242 0 feedthrough
rlabel pdiffusion 507 -2242 507 -2242 0 feedthrough
rlabel pdiffusion 514 -2242 514 -2242 0 feedthrough
rlabel pdiffusion 521 -2242 521 -2242 0 cellNo=317
rlabel pdiffusion 528 -2242 528 -2242 0 cellNo=266
rlabel pdiffusion 535 -2242 535 -2242 0 feedthrough
rlabel pdiffusion 542 -2242 542 -2242 0 feedthrough
rlabel pdiffusion 549 -2242 549 -2242 0 feedthrough
rlabel pdiffusion 556 -2242 556 -2242 0 cellNo=287
rlabel pdiffusion 563 -2242 563 -2242 0 feedthrough
rlabel pdiffusion 570 -2242 570 -2242 0 feedthrough
rlabel pdiffusion 577 -2242 577 -2242 0 feedthrough
rlabel pdiffusion 584 -2242 584 -2242 0 feedthrough
rlabel pdiffusion 591 -2242 591 -2242 0 feedthrough
rlabel pdiffusion 598 -2242 598 -2242 0 feedthrough
rlabel pdiffusion 605 -2242 605 -2242 0 feedthrough
rlabel pdiffusion 612 -2242 612 -2242 0 feedthrough
rlabel pdiffusion 619 -2242 619 -2242 0 cellNo=350
rlabel pdiffusion 626 -2242 626 -2242 0 cellNo=430
rlabel pdiffusion 633 -2242 633 -2242 0 feedthrough
rlabel pdiffusion 640 -2242 640 -2242 0 feedthrough
rlabel pdiffusion 647 -2242 647 -2242 0 cellNo=34
rlabel pdiffusion 654 -2242 654 -2242 0 feedthrough
rlabel pdiffusion 661 -2242 661 -2242 0 feedthrough
rlabel pdiffusion 668 -2242 668 -2242 0 feedthrough
rlabel pdiffusion 675 -2242 675 -2242 0 cellNo=442
rlabel pdiffusion 682 -2242 682 -2242 0 feedthrough
rlabel pdiffusion 689 -2242 689 -2242 0 feedthrough
rlabel pdiffusion 696 -2242 696 -2242 0 feedthrough
rlabel pdiffusion 703 -2242 703 -2242 0 feedthrough
rlabel pdiffusion 710 -2242 710 -2242 0 feedthrough
rlabel pdiffusion 717 -2242 717 -2242 0 feedthrough
rlabel pdiffusion 724 -2242 724 -2242 0 feedthrough
rlabel pdiffusion 731 -2242 731 -2242 0 feedthrough
rlabel pdiffusion 738 -2242 738 -2242 0 feedthrough
rlabel pdiffusion 745 -2242 745 -2242 0 feedthrough
rlabel pdiffusion 752 -2242 752 -2242 0 feedthrough
rlabel pdiffusion 759 -2242 759 -2242 0 feedthrough
rlabel pdiffusion 766 -2242 766 -2242 0 feedthrough
rlabel pdiffusion 773 -2242 773 -2242 0 feedthrough
rlabel pdiffusion 780 -2242 780 -2242 0 feedthrough
rlabel pdiffusion 787 -2242 787 -2242 0 feedthrough
rlabel pdiffusion 794 -2242 794 -2242 0 feedthrough
rlabel pdiffusion 801 -2242 801 -2242 0 feedthrough
rlabel pdiffusion 808 -2242 808 -2242 0 cellNo=391
rlabel pdiffusion 815 -2242 815 -2242 0 feedthrough
rlabel pdiffusion 822 -2242 822 -2242 0 feedthrough
rlabel pdiffusion 829 -2242 829 -2242 0 feedthrough
rlabel pdiffusion 836 -2242 836 -2242 0 feedthrough
rlabel pdiffusion 843 -2242 843 -2242 0 feedthrough
rlabel pdiffusion 850 -2242 850 -2242 0 feedthrough
rlabel pdiffusion 857 -2242 857 -2242 0 feedthrough
rlabel pdiffusion 864 -2242 864 -2242 0 feedthrough
rlabel pdiffusion 871 -2242 871 -2242 0 cellNo=212
rlabel pdiffusion 878 -2242 878 -2242 0 feedthrough
rlabel pdiffusion 885 -2242 885 -2242 0 feedthrough
rlabel pdiffusion 892 -2242 892 -2242 0 feedthrough
rlabel pdiffusion 899 -2242 899 -2242 0 feedthrough
rlabel pdiffusion 906 -2242 906 -2242 0 feedthrough
rlabel pdiffusion 913 -2242 913 -2242 0 feedthrough
rlabel pdiffusion 920 -2242 920 -2242 0 feedthrough
rlabel pdiffusion 927 -2242 927 -2242 0 feedthrough
rlabel pdiffusion 934 -2242 934 -2242 0 cellNo=456
rlabel pdiffusion 941 -2242 941 -2242 0 feedthrough
rlabel pdiffusion 948 -2242 948 -2242 0 feedthrough
rlabel pdiffusion 955 -2242 955 -2242 0 feedthrough
rlabel pdiffusion 962 -2242 962 -2242 0 feedthrough
rlabel pdiffusion 969 -2242 969 -2242 0 feedthrough
rlabel pdiffusion 976 -2242 976 -2242 0 feedthrough
rlabel pdiffusion 983 -2242 983 -2242 0 cellNo=396
rlabel pdiffusion 990 -2242 990 -2242 0 feedthrough
rlabel pdiffusion 997 -2242 997 -2242 0 feedthrough
rlabel pdiffusion 1004 -2242 1004 -2242 0 feedthrough
rlabel pdiffusion 1011 -2242 1011 -2242 0 feedthrough
rlabel pdiffusion 1018 -2242 1018 -2242 0 feedthrough
rlabel pdiffusion 1025 -2242 1025 -2242 0 feedthrough
rlabel pdiffusion 1032 -2242 1032 -2242 0 feedthrough
rlabel pdiffusion 1039 -2242 1039 -2242 0 feedthrough
rlabel pdiffusion 1046 -2242 1046 -2242 0 feedthrough
rlabel pdiffusion 1053 -2242 1053 -2242 0 feedthrough
rlabel pdiffusion 1060 -2242 1060 -2242 0 feedthrough
rlabel pdiffusion 1067 -2242 1067 -2242 0 feedthrough
rlabel pdiffusion 1074 -2242 1074 -2242 0 feedthrough
rlabel pdiffusion 1081 -2242 1081 -2242 0 feedthrough
rlabel pdiffusion 1088 -2242 1088 -2242 0 feedthrough
rlabel pdiffusion 1095 -2242 1095 -2242 0 feedthrough
rlabel pdiffusion 1102 -2242 1102 -2242 0 feedthrough
rlabel pdiffusion 1109 -2242 1109 -2242 0 feedthrough
rlabel pdiffusion 1116 -2242 1116 -2242 0 feedthrough
rlabel pdiffusion 1123 -2242 1123 -2242 0 feedthrough
rlabel pdiffusion 1130 -2242 1130 -2242 0 feedthrough
rlabel pdiffusion 1137 -2242 1137 -2242 0 feedthrough
rlabel pdiffusion 1144 -2242 1144 -2242 0 feedthrough
rlabel pdiffusion 1151 -2242 1151 -2242 0 feedthrough
rlabel pdiffusion 1158 -2242 1158 -2242 0 feedthrough
rlabel pdiffusion 1165 -2242 1165 -2242 0 feedthrough
rlabel pdiffusion 1172 -2242 1172 -2242 0 feedthrough
rlabel pdiffusion 1179 -2242 1179 -2242 0 feedthrough
rlabel pdiffusion 1186 -2242 1186 -2242 0 feedthrough
rlabel pdiffusion 1193 -2242 1193 -2242 0 feedthrough
rlabel pdiffusion 1200 -2242 1200 -2242 0 feedthrough
rlabel pdiffusion 1207 -2242 1207 -2242 0 feedthrough
rlabel pdiffusion 1214 -2242 1214 -2242 0 feedthrough
rlabel pdiffusion 1221 -2242 1221 -2242 0 feedthrough
rlabel pdiffusion 1228 -2242 1228 -2242 0 feedthrough
rlabel pdiffusion 1235 -2242 1235 -2242 0 feedthrough
rlabel pdiffusion 1242 -2242 1242 -2242 0 feedthrough
rlabel pdiffusion 1249 -2242 1249 -2242 0 feedthrough
rlabel pdiffusion 1256 -2242 1256 -2242 0 feedthrough
rlabel pdiffusion 1263 -2242 1263 -2242 0 feedthrough
rlabel pdiffusion 1270 -2242 1270 -2242 0 feedthrough
rlabel pdiffusion 1277 -2242 1277 -2242 0 feedthrough
rlabel pdiffusion 1284 -2242 1284 -2242 0 feedthrough
rlabel pdiffusion 1291 -2242 1291 -2242 0 feedthrough
rlabel pdiffusion 1298 -2242 1298 -2242 0 feedthrough
rlabel pdiffusion 1305 -2242 1305 -2242 0 feedthrough
rlabel pdiffusion 1312 -2242 1312 -2242 0 feedthrough
rlabel pdiffusion 3 -2367 3 -2367 0 cellNo=534
rlabel pdiffusion 10 -2367 10 -2367 0 feedthrough
rlabel pdiffusion 17 -2367 17 -2367 0 feedthrough
rlabel pdiffusion 24 -2367 24 -2367 0 feedthrough
rlabel pdiffusion 31 -2367 31 -2367 0 feedthrough
rlabel pdiffusion 38 -2367 38 -2367 0 cellNo=471
rlabel pdiffusion 45 -2367 45 -2367 0 feedthrough
rlabel pdiffusion 52 -2367 52 -2367 0 cellNo=121
rlabel pdiffusion 59 -2367 59 -2367 0 cellNo=443
rlabel pdiffusion 66 -2367 66 -2367 0 feedthrough
rlabel pdiffusion 73 -2367 73 -2367 0 feedthrough
rlabel pdiffusion 80 -2367 80 -2367 0 feedthrough
rlabel pdiffusion 87 -2367 87 -2367 0 feedthrough
rlabel pdiffusion 94 -2367 94 -2367 0 cellNo=272
rlabel pdiffusion 101 -2367 101 -2367 0 feedthrough
rlabel pdiffusion 108 -2367 108 -2367 0 feedthrough
rlabel pdiffusion 115 -2367 115 -2367 0 feedthrough
rlabel pdiffusion 122 -2367 122 -2367 0 feedthrough
rlabel pdiffusion 129 -2367 129 -2367 0 feedthrough
rlabel pdiffusion 136 -2367 136 -2367 0 cellNo=424
rlabel pdiffusion 143 -2367 143 -2367 0 feedthrough
rlabel pdiffusion 150 -2367 150 -2367 0 cellNo=42
rlabel pdiffusion 157 -2367 157 -2367 0 feedthrough
rlabel pdiffusion 164 -2367 164 -2367 0 feedthrough
rlabel pdiffusion 171 -2367 171 -2367 0 feedthrough
rlabel pdiffusion 178 -2367 178 -2367 0 feedthrough
rlabel pdiffusion 185 -2367 185 -2367 0 feedthrough
rlabel pdiffusion 192 -2367 192 -2367 0 feedthrough
rlabel pdiffusion 199 -2367 199 -2367 0 feedthrough
rlabel pdiffusion 206 -2367 206 -2367 0 feedthrough
rlabel pdiffusion 213 -2367 213 -2367 0 feedthrough
rlabel pdiffusion 220 -2367 220 -2367 0 feedthrough
rlabel pdiffusion 227 -2367 227 -2367 0 feedthrough
rlabel pdiffusion 234 -2367 234 -2367 0 feedthrough
rlabel pdiffusion 241 -2367 241 -2367 0 feedthrough
rlabel pdiffusion 248 -2367 248 -2367 0 feedthrough
rlabel pdiffusion 255 -2367 255 -2367 0 feedthrough
rlabel pdiffusion 262 -2367 262 -2367 0 feedthrough
rlabel pdiffusion 269 -2367 269 -2367 0 feedthrough
rlabel pdiffusion 276 -2367 276 -2367 0 feedthrough
rlabel pdiffusion 283 -2367 283 -2367 0 feedthrough
rlabel pdiffusion 290 -2367 290 -2367 0 feedthrough
rlabel pdiffusion 297 -2367 297 -2367 0 feedthrough
rlabel pdiffusion 304 -2367 304 -2367 0 cellNo=578
rlabel pdiffusion 311 -2367 311 -2367 0 feedthrough
rlabel pdiffusion 318 -2367 318 -2367 0 cellNo=16
rlabel pdiffusion 325 -2367 325 -2367 0 feedthrough
rlabel pdiffusion 332 -2367 332 -2367 0 feedthrough
rlabel pdiffusion 339 -2367 339 -2367 0 cellNo=545
rlabel pdiffusion 346 -2367 346 -2367 0 feedthrough
rlabel pdiffusion 353 -2367 353 -2367 0 feedthrough
rlabel pdiffusion 360 -2367 360 -2367 0 feedthrough
rlabel pdiffusion 367 -2367 367 -2367 0 feedthrough
rlabel pdiffusion 374 -2367 374 -2367 0 feedthrough
rlabel pdiffusion 381 -2367 381 -2367 0 feedthrough
rlabel pdiffusion 388 -2367 388 -2367 0 feedthrough
rlabel pdiffusion 395 -2367 395 -2367 0 cellNo=590
rlabel pdiffusion 402 -2367 402 -2367 0 feedthrough
rlabel pdiffusion 409 -2367 409 -2367 0 feedthrough
rlabel pdiffusion 416 -2367 416 -2367 0 feedthrough
rlabel pdiffusion 423 -2367 423 -2367 0 cellNo=120
rlabel pdiffusion 430 -2367 430 -2367 0 feedthrough
rlabel pdiffusion 437 -2367 437 -2367 0 cellNo=12
rlabel pdiffusion 444 -2367 444 -2367 0 feedthrough
rlabel pdiffusion 451 -2367 451 -2367 0 feedthrough
rlabel pdiffusion 458 -2367 458 -2367 0 feedthrough
rlabel pdiffusion 465 -2367 465 -2367 0 feedthrough
rlabel pdiffusion 472 -2367 472 -2367 0 feedthrough
rlabel pdiffusion 479 -2367 479 -2367 0 feedthrough
rlabel pdiffusion 486 -2367 486 -2367 0 feedthrough
rlabel pdiffusion 493 -2367 493 -2367 0 feedthrough
rlabel pdiffusion 500 -2367 500 -2367 0 feedthrough
rlabel pdiffusion 507 -2367 507 -2367 0 feedthrough
rlabel pdiffusion 514 -2367 514 -2367 0 cellNo=413
rlabel pdiffusion 521 -2367 521 -2367 0 feedthrough
rlabel pdiffusion 528 -2367 528 -2367 0 feedthrough
rlabel pdiffusion 535 -2367 535 -2367 0 feedthrough
rlabel pdiffusion 542 -2367 542 -2367 0 feedthrough
rlabel pdiffusion 549 -2367 549 -2367 0 feedthrough
rlabel pdiffusion 556 -2367 556 -2367 0 cellNo=339
rlabel pdiffusion 563 -2367 563 -2367 0 feedthrough
rlabel pdiffusion 570 -2367 570 -2367 0 feedthrough
rlabel pdiffusion 577 -2367 577 -2367 0 cellNo=439
rlabel pdiffusion 584 -2367 584 -2367 0 feedthrough
rlabel pdiffusion 591 -2367 591 -2367 0 cellNo=550
rlabel pdiffusion 598 -2367 598 -2367 0 feedthrough
rlabel pdiffusion 605 -2367 605 -2367 0 feedthrough
rlabel pdiffusion 612 -2367 612 -2367 0 feedthrough
rlabel pdiffusion 619 -2367 619 -2367 0 feedthrough
rlabel pdiffusion 626 -2367 626 -2367 0 feedthrough
rlabel pdiffusion 633 -2367 633 -2367 0 cellNo=470
rlabel pdiffusion 640 -2367 640 -2367 0 feedthrough
rlabel pdiffusion 647 -2367 647 -2367 0 feedthrough
rlabel pdiffusion 654 -2367 654 -2367 0 feedthrough
rlabel pdiffusion 661 -2367 661 -2367 0 cellNo=278
rlabel pdiffusion 668 -2367 668 -2367 0 feedthrough
rlabel pdiffusion 675 -2367 675 -2367 0 feedthrough
rlabel pdiffusion 682 -2367 682 -2367 0 feedthrough
rlabel pdiffusion 689 -2367 689 -2367 0 feedthrough
rlabel pdiffusion 696 -2367 696 -2367 0 feedthrough
rlabel pdiffusion 703 -2367 703 -2367 0 feedthrough
rlabel pdiffusion 710 -2367 710 -2367 0 feedthrough
rlabel pdiffusion 717 -2367 717 -2367 0 feedthrough
rlabel pdiffusion 724 -2367 724 -2367 0 cellNo=291
rlabel pdiffusion 731 -2367 731 -2367 0 feedthrough
rlabel pdiffusion 738 -2367 738 -2367 0 feedthrough
rlabel pdiffusion 745 -2367 745 -2367 0 cellNo=311
rlabel pdiffusion 752 -2367 752 -2367 0 feedthrough
rlabel pdiffusion 759 -2367 759 -2367 0 cellNo=598
rlabel pdiffusion 766 -2367 766 -2367 0 feedthrough
rlabel pdiffusion 773 -2367 773 -2367 0 feedthrough
rlabel pdiffusion 780 -2367 780 -2367 0 feedthrough
rlabel pdiffusion 787 -2367 787 -2367 0 feedthrough
rlabel pdiffusion 794 -2367 794 -2367 0 feedthrough
rlabel pdiffusion 801 -2367 801 -2367 0 feedthrough
rlabel pdiffusion 808 -2367 808 -2367 0 cellNo=577
rlabel pdiffusion 815 -2367 815 -2367 0 feedthrough
rlabel pdiffusion 822 -2367 822 -2367 0 feedthrough
rlabel pdiffusion 829 -2367 829 -2367 0 feedthrough
rlabel pdiffusion 836 -2367 836 -2367 0 feedthrough
rlabel pdiffusion 843 -2367 843 -2367 0 feedthrough
rlabel pdiffusion 850 -2367 850 -2367 0 cellNo=575
rlabel pdiffusion 857 -2367 857 -2367 0 feedthrough
rlabel pdiffusion 864 -2367 864 -2367 0 feedthrough
rlabel pdiffusion 871 -2367 871 -2367 0 feedthrough
rlabel pdiffusion 878 -2367 878 -2367 0 feedthrough
rlabel pdiffusion 885 -2367 885 -2367 0 feedthrough
rlabel pdiffusion 892 -2367 892 -2367 0 feedthrough
rlabel pdiffusion 899 -2367 899 -2367 0 feedthrough
rlabel pdiffusion 906 -2367 906 -2367 0 feedthrough
rlabel pdiffusion 913 -2367 913 -2367 0 feedthrough
rlabel pdiffusion 920 -2367 920 -2367 0 feedthrough
rlabel pdiffusion 927 -2367 927 -2367 0 feedthrough
rlabel pdiffusion 934 -2367 934 -2367 0 feedthrough
rlabel pdiffusion 941 -2367 941 -2367 0 feedthrough
rlabel pdiffusion 948 -2367 948 -2367 0 feedthrough
rlabel pdiffusion 955 -2367 955 -2367 0 feedthrough
rlabel pdiffusion 962 -2367 962 -2367 0 feedthrough
rlabel pdiffusion 969 -2367 969 -2367 0 feedthrough
rlabel pdiffusion 976 -2367 976 -2367 0 feedthrough
rlabel pdiffusion 983 -2367 983 -2367 0 feedthrough
rlabel pdiffusion 990 -2367 990 -2367 0 feedthrough
rlabel pdiffusion 997 -2367 997 -2367 0 feedthrough
rlabel pdiffusion 1004 -2367 1004 -2367 0 feedthrough
rlabel pdiffusion 1011 -2367 1011 -2367 0 feedthrough
rlabel pdiffusion 1018 -2367 1018 -2367 0 feedthrough
rlabel pdiffusion 1025 -2367 1025 -2367 0 feedthrough
rlabel pdiffusion 1032 -2367 1032 -2367 0 cellNo=567
rlabel pdiffusion 1039 -2367 1039 -2367 0 feedthrough
rlabel pdiffusion 1046 -2367 1046 -2367 0 feedthrough
rlabel pdiffusion 1053 -2367 1053 -2367 0 feedthrough
rlabel pdiffusion 1060 -2367 1060 -2367 0 feedthrough
rlabel pdiffusion 1067 -2367 1067 -2367 0 feedthrough
rlabel pdiffusion 1074 -2367 1074 -2367 0 feedthrough
rlabel pdiffusion 1081 -2367 1081 -2367 0 feedthrough
rlabel pdiffusion 1088 -2367 1088 -2367 0 feedthrough
rlabel pdiffusion 1095 -2367 1095 -2367 0 feedthrough
rlabel pdiffusion 1102 -2367 1102 -2367 0 feedthrough
rlabel pdiffusion 1109 -2367 1109 -2367 0 feedthrough
rlabel pdiffusion 1116 -2367 1116 -2367 0 feedthrough
rlabel pdiffusion 1123 -2367 1123 -2367 0 feedthrough
rlabel pdiffusion 1130 -2367 1130 -2367 0 feedthrough
rlabel pdiffusion 1137 -2367 1137 -2367 0 feedthrough
rlabel pdiffusion 1144 -2367 1144 -2367 0 feedthrough
rlabel pdiffusion 1151 -2367 1151 -2367 0 feedthrough
rlabel pdiffusion 1158 -2367 1158 -2367 0 feedthrough
rlabel pdiffusion 1165 -2367 1165 -2367 0 feedthrough
rlabel pdiffusion 1172 -2367 1172 -2367 0 feedthrough
rlabel pdiffusion 1179 -2367 1179 -2367 0 feedthrough
rlabel pdiffusion 1186 -2367 1186 -2367 0 feedthrough
rlabel pdiffusion 1193 -2367 1193 -2367 0 feedthrough
rlabel pdiffusion 1200 -2367 1200 -2367 0 feedthrough
rlabel pdiffusion 1207 -2367 1207 -2367 0 feedthrough
rlabel pdiffusion 1214 -2367 1214 -2367 0 feedthrough
rlabel pdiffusion 1221 -2367 1221 -2367 0 feedthrough
rlabel pdiffusion 1228 -2367 1228 -2367 0 feedthrough
rlabel pdiffusion 1235 -2367 1235 -2367 0 feedthrough
rlabel pdiffusion 1242 -2367 1242 -2367 0 feedthrough
rlabel pdiffusion 1249 -2367 1249 -2367 0 feedthrough
rlabel pdiffusion 59 -2464 59 -2464 0 feedthrough
rlabel pdiffusion 66 -2464 66 -2464 0 feedthrough
rlabel pdiffusion 73 -2464 73 -2464 0 feedthrough
rlabel pdiffusion 80 -2464 80 -2464 0 feedthrough
rlabel pdiffusion 87 -2464 87 -2464 0 feedthrough
rlabel pdiffusion 94 -2464 94 -2464 0 feedthrough
rlabel pdiffusion 101 -2464 101 -2464 0 feedthrough
rlabel pdiffusion 108 -2464 108 -2464 0 feedthrough
rlabel pdiffusion 115 -2464 115 -2464 0 feedthrough
rlabel pdiffusion 122 -2464 122 -2464 0 cellNo=371
rlabel pdiffusion 129 -2464 129 -2464 0 cellNo=574
rlabel pdiffusion 136 -2464 136 -2464 0 feedthrough
rlabel pdiffusion 143 -2464 143 -2464 0 feedthrough
rlabel pdiffusion 150 -2464 150 -2464 0 feedthrough
rlabel pdiffusion 157 -2464 157 -2464 0 feedthrough
rlabel pdiffusion 164 -2464 164 -2464 0 cellNo=264
rlabel pdiffusion 171 -2464 171 -2464 0 cellNo=8
rlabel pdiffusion 178 -2464 178 -2464 0 feedthrough
rlabel pdiffusion 185 -2464 185 -2464 0 feedthrough
rlabel pdiffusion 192 -2464 192 -2464 0 feedthrough
rlabel pdiffusion 199 -2464 199 -2464 0 cellNo=248
rlabel pdiffusion 206 -2464 206 -2464 0 feedthrough
rlabel pdiffusion 213 -2464 213 -2464 0 feedthrough
rlabel pdiffusion 220 -2464 220 -2464 0 feedthrough
rlabel pdiffusion 227 -2464 227 -2464 0 feedthrough
rlabel pdiffusion 234 -2464 234 -2464 0 feedthrough
rlabel pdiffusion 241 -2464 241 -2464 0 feedthrough
rlabel pdiffusion 248 -2464 248 -2464 0 feedthrough
rlabel pdiffusion 255 -2464 255 -2464 0 feedthrough
rlabel pdiffusion 262 -2464 262 -2464 0 feedthrough
rlabel pdiffusion 269 -2464 269 -2464 0 feedthrough
rlabel pdiffusion 276 -2464 276 -2464 0 feedthrough
rlabel pdiffusion 283 -2464 283 -2464 0 feedthrough
rlabel pdiffusion 290 -2464 290 -2464 0 feedthrough
rlabel pdiffusion 297 -2464 297 -2464 0 feedthrough
rlabel pdiffusion 304 -2464 304 -2464 0 feedthrough
rlabel pdiffusion 311 -2464 311 -2464 0 feedthrough
rlabel pdiffusion 318 -2464 318 -2464 0 feedthrough
rlabel pdiffusion 325 -2464 325 -2464 0 feedthrough
rlabel pdiffusion 332 -2464 332 -2464 0 feedthrough
rlabel pdiffusion 339 -2464 339 -2464 0 feedthrough
rlabel pdiffusion 346 -2464 346 -2464 0 feedthrough
rlabel pdiffusion 353 -2464 353 -2464 0 cellNo=455
rlabel pdiffusion 360 -2464 360 -2464 0 feedthrough
rlabel pdiffusion 367 -2464 367 -2464 0 feedthrough
rlabel pdiffusion 374 -2464 374 -2464 0 cellNo=123
rlabel pdiffusion 381 -2464 381 -2464 0 feedthrough
rlabel pdiffusion 388 -2464 388 -2464 0 feedthrough
rlabel pdiffusion 395 -2464 395 -2464 0 feedthrough
rlabel pdiffusion 402 -2464 402 -2464 0 feedthrough
rlabel pdiffusion 409 -2464 409 -2464 0 feedthrough
rlabel pdiffusion 416 -2464 416 -2464 0 feedthrough
rlabel pdiffusion 423 -2464 423 -2464 0 feedthrough
rlabel pdiffusion 430 -2464 430 -2464 0 feedthrough
rlabel pdiffusion 437 -2464 437 -2464 0 cellNo=67
rlabel pdiffusion 444 -2464 444 -2464 0 cellNo=547
rlabel pdiffusion 451 -2464 451 -2464 0 feedthrough
rlabel pdiffusion 458 -2464 458 -2464 0 feedthrough
rlabel pdiffusion 465 -2464 465 -2464 0 cellNo=498
rlabel pdiffusion 472 -2464 472 -2464 0 feedthrough
rlabel pdiffusion 479 -2464 479 -2464 0 feedthrough
rlabel pdiffusion 486 -2464 486 -2464 0 feedthrough
rlabel pdiffusion 493 -2464 493 -2464 0 feedthrough
rlabel pdiffusion 500 -2464 500 -2464 0 feedthrough
rlabel pdiffusion 507 -2464 507 -2464 0 feedthrough
rlabel pdiffusion 514 -2464 514 -2464 0 cellNo=216
rlabel pdiffusion 521 -2464 521 -2464 0 feedthrough
rlabel pdiffusion 528 -2464 528 -2464 0 feedthrough
rlabel pdiffusion 535 -2464 535 -2464 0 feedthrough
rlabel pdiffusion 542 -2464 542 -2464 0 feedthrough
rlabel pdiffusion 549 -2464 549 -2464 0 feedthrough
rlabel pdiffusion 556 -2464 556 -2464 0 feedthrough
rlabel pdiffusion 563 -2464 563 -2464 0 cellNo=330
rlabel pdiffusion 570 -2464 570 -2464 0 cellNo=360
rlabel pdiffusion 577 -2464 577 -2464 0 feedthrough
rlabel pdiffusion 584 -2464 584 -2464 0 feedthrough
rlabel pdiffusion 591 -2464 591 -2464 0 feedthrough
rlabel pdiffusion 598 -2464 598 -2464 0 feedthrough
rlabel pdiffusion 605 -2464 605 -2464 0 feedthrough
rlabel pdiffusion 612 -2464 612 -2464 0 cellNo=407
rlabel pdiffusion 619 -2464 619 -2464 0 feedthrough
rlabel pdiffusion 626 -2464 626 -2464 0 feedthrough
rlabel pdiffusion 633 -2464 633 -2464 0 feedthrough
rlabel pdiffusion 640 -2464 640 -2464 0 feedthrough
rlabel pdiffusion 647 -2464 647 -2464 0 feedthrough
rlabel pdiffusion 654 -2464 654 -2464 0 feedthrough
rlabel pdiffusion 661 -2464 661 -2464 0 cellNo=328
rlabel pdiffusion 668 -2464 668 -2464 0 feedthrough
rlabel pdiffusion 675 -2464 675 -2464 0 cellNo=45
rlabel pdiffusion 682 -2464 682 -2464 0 feedthrough
rlabel pdiffusion 689 -2464 689 -2464 0 feedthrough
rlabel pdiffusion 696 -2464 696 -2464 0 cellNo=296
rlabel pdiffusion 703 -2464 703 -2464 0 feedthrough
rlabel pdiffusion 710 -2464 710 -2464 0 feedthrough
rlabel pdiffusion 717 -2464 717 -2464 0 feedthrough
rlabel pdiffusion 724 -2464 724 -2464 0 cellNo=417
rlabel pdiffusion 731 -2464 731 -2464 0 feedthrough
rlabel pdiffusion 738 -2464 738 -2464 0 feedthrough
rlabel pdiffusion 745 -2464 745 -2464 0 feedthrough
rlabel pdiffusion 752 -2464 752 -2464 0 feedthrough
rlabel pdiffusion 759 -2464 759 -2464 0 feedthrough
rlabel pdiffusion 766 -2464 766 -2464 0 feedthrough
rlabel pdiffusion 773 -2464 773 -2464 0 feedthrough
rlabel pdiffusion 780 -2464 780 -2464 0 feedthrough
rlabel pdiffusion 787 -2464 787 -2464 0 feedthrough
rlabel pdiffusion 794 -2464 794 -2464 0 cellNo=531
rlabel pdiffusion 801 -2464 801 -2464 0 feedthrough
rlabel pdiffusion 808 -2464 808 -2464 0 feedthrough
rlabel pdiffusion 815 -2464 815 -2464 0 feedthrough
rlabel pdiffusion 822 -2464 822 -2464 0 feedthrough
rlabel pdiffusion 829 -2464 829 -2464 0 cellNo=318
rlabel pdiffusion 836 -2464 836 -2464 0 feedthrough
rlabel pdiffusion 843 -2464 843 -2464 0 feedthrough
rlabel pdiffusion 850 -2464 850 -2464 0 feedthrough
rlabel pdiffusion 857 -2464 857 -2464 0 feedthrough
rlabel pdiffusion 864 -2464 864 -2464 0 feedthrough
rlabel pdiffusion 871 -2464 871 -2464 0 feedthrough
rlabel pdiffusion 878 -2464 878 -2464 0 feedthrough
rlabel pdiffusion 885 -2464 885 -2464 0 feedthrough
rlabel pdiffusion 892 -2464 892 -2464 0 feedthrough
rlabel pdiffusion 899 -2464 899 -2464 0 feedthrough
rlabel pdiffusion 906 -2464 906 -2464 0 cellNo=528
rlabel pdiffusion 913 -2464 913 -2464 0 feedthrough
rlabel pdiffusion 920 -2464 920 -2464 0 feedthrough
rlabel pdiffusion 927 -2464 927 -2464 0 feedthrough
rlabel pdiffusion 934 -2464 934 -2464 0 feedthrough
rlabel pdiffusion 941 -2464 941 -2464 0 cellNo=409
rlabel pdiffusion 948 -2464 948 -2464 0 feedthrough
rlabel pdiffusion 955 -2464 955 -2464 0 feedthrough
rlabel pdiffusion 962 -2464 962 -2464 0 feedthrough
rlabel pdiffusion 969 -2464 969 -2464 0 feedthrough
rlabel pdiffusion 976 -2464 976 -2464 0 feedthrough
rlabel pdiffusion 983 -2464 983 -2464 0 feedthrough
rlabel pdiffusion 990 -2464 990 -2464 0 feedthrough
rlabel pdiffusion 997 -2464 997 -2464 0 feedthrough
rlabel pdiffusion 1004 -2464 1004 -2464 0 feedthrough
rlabel pdiffusion 1011 -2464 1011 -2464 0 cellNo=502
rlabel pdiffusion 1018 -2464 1018 -2464 0 feedthrough
rlabel pdiffusion 1025 -2464 1025 -2464 0 feedthrough
rlabel pdiffusion 1032 -2464 1032 -2464 0 feedthrough
rlabel pdiffusion 1060 -2464 1060 -2464 0 feedthrough
rlabel pdiffusion 1067 -2464 1067 -2464 0 feedthrough
rlabel pdiffusion 1074 -2464 1074 -2464 0 feedthrough
rlabel pdiffusion 1081 -2464 1081 -2464 0 feedthrough
rlabel pdiffusion 1088 -2464 1088 -2464 0 feedthrough
rlabel pdiffusion 1095 -2464 1095 -2464 0 feedthrough
rlabel pdiffusion 1102 -2464 1102 -2464 0 cellNo=487
rlabel pdiffusion 1109 -2464 1109 -2464 0 feedthrough
rlabel pdiffusion 1130 -2464 1130 -2464 0 feedthrough
rlabel pdiffusion 1193 -2464 1193 -2464 0 feedthrough
rlabel pdiffusion 129 -2547 129 -2547 0 feedthrough
rlabel pdiffusion 136 -2547 136 -2547 0 feedthrough
rlabel pdiffusion 227 -2547 227 -2547 0 feedthrough
rlabel pdiffusion 234 -2547 234 -2547 0 feedthrough
rlabel pdiffusion 248 -2547 248 -2547 0 feedthrough
rlabel pdiffusion 255 -2547 255 -2547 0 feedthrough
rlabel pdiffusion 262 -2547 262 -2547 0 feedthrough
rlabel pdiffusion 269 -2547 269 -2547 0 feedthrough
rlabel pdiffusion 276 -2547 276 -2547 0 cellNo=335
rlabel pdiffusion 283 -2547 283 -2547 0 feedthrough
rlabel pdiffusion 290 -2547 290 -2547 0 feedthrough
rlabel pdiffusion 297 -2547 297 -2547 0 feedthrough
rlabel pdiffusion 304 -2547 304 -2547 0 feedthrough
rlabel pdiffusion 311 -2547 311 -2547 0 feedthrough
rlabel pdiffusion 318 -2547 318 -2547 0 feedthrough
rlabel pdiffusion 325 -2547 325 -2547 0 cellNo=500
rlabel pdiffusion 332 -2547 332 -2547 0 feedthrough
rlabel pdiffusion 339 -2547 339 -2547 0 feedthrough
rlabel pdiffusion 346 -2547 346 -2547 0 feedthrough
rlabel pdiffusion 353 -2547 353 -2547 0 feedthrough
rlabel pdiffusion 360 -2547 360 -2547 0 feedthrough
rlabel pdiffusion 367 -2547 367 -2547 0 cellNo=97
rlabel pdiffusion 374 -2547 374 -2547 0 feedthrough
rlabel pdiffusion 381 -2547 381 -2547 0 feedthrough
rlabel pdiffusion 388 -2547 388 -2547 0 cellNo=505
rlabel pdiffusion 395 -2547 395 -2547 0 feedthrough
rlabel pdiffusion 402 -2547 402 -2547 0 feedthrough
rlabel pdiffusion 409 -2547 409 -2547 0 feedthrough
rlabel pdiffusion 416 -2547 416 -2547 0 feedthrough
rlabel pdiffusion 423 -2547 423 -2547 0 feedthrough
rlabel pdiffusion 430 -2547 430 -2547 0 feedthrough
rlabel pdiffusion 437 -2547 437 -2547 0 feedthrough
rlabel pdiffusion 444 -2547 444 -2547 0 feedthrough
rlabel pdiffusion 451 -2547 451 -2547 0 feedthrough
rlabel pdiffusion 458 -2547 458 -2547 0 cellNo=564
rlabel pdiffusion 465 -2547 465 -2547 0 feedthrough
rlabel pdiffusion 472 -2547 472 -2547 0 cellNo=568
rlabel pdiffusion 479 -2547 479 -2547 0 feedthrough
rlabel pdiffusion 486 -2547 486 -2547 0 cellNo=349
rlabel pdiffusion 493 -2547 493 -2547 0 feedthrough
rlabel pdiffusion 500 -2547 500 -2547 0 feedthrough
rlabel pdiffusion 507 -2547 507 -2547 0 cellNo=440
rlabel pdiffusion 514 -2547 514 -2547 0 feedthrough
rlabel pdiffusion 521 -2547 521 -2547 0 cellNo=463
rlabel pdiffusion 528 -2547 528 -2547 0 cellNo=366
rlabel pdiffusion 535 -2547 535 -2547 0 feedthrough
rlabel pdiffusion 542 -2547 542 -2547 0 cellNo=280
rlabel pdiffusion 549 -2547 549 -2547 0 cellNo=474
rlabel pdiffusion 556 -2547 556 -2547 0 feedthrough
rlabel pdiffusion 563 -2547 563 -2547 0 feedthrough
rlabel pdiffusion 570 -2547 570 -2547 0 cellNo=268
rlabel pdiffusion 577 -2547 577 -2547 0 feedthrough
rlabel pdiffusion 584 -2547 584 -2547 0 cellNo=581
rlabel pdiffusion 591 -2547 591 -2547 0 cellNo=546
rlabel pdiffusion 598 -2547 598 -2547 0 feedthrough
rlabel pdiffusion 605 -2547 605 -2547 0 feedthrough
rlabel pdiffusion 612 -2547 612 -2547 0 feedthrough
rlabel pdiffusion 619 -2547 619 -2547 0 cellNo=527
rlabel pdiffusion 626 -2547 626 -2547 0 feedthrough
rlabel pdiffusion 633 -2547 633 -2547 0 feedthrough
rlabel pdiffusion 640 -2547 640 -2547 0 feedthrough
rlabel pdiffusion 647 -2547 647 -2547 0 feedthrough
rlabel pdiffusion 654 -2547 654 -2547 0 feedthrough
rlabel pdiffusion 661 -2547 661 -2547 0 feedthrough
rlabel pdiffusion 668 -2547 668 -2547 0 feedthrough
rlabel pdiffusion 675 -2547 675 -2547 0 feedthrough
rlabel pdiffusion 682 -2547 682 -2547 0 cellNo=559
rlabel pdiffusion 689 -2547 689 -2547 0 cellNo=489
rlabel pdiffusion 696 -2547 696 -2547 0 feedthrough
rlabel pdiffusion 703 -2547 703 -2547 0 feedthrough
rlabel pdiffusion 710 -2547 710 -2547 0 feedthrough
rlabel pdiffusion 717 -2547 717 -2547 0 feedthrough
rlabel pdiffusion 724 -2547 724 -2547 0 feedthrough
rlabel pdiffusion 731 -2547 731 -2547 0 feedthrough
rlabel pdiffusion 738 -2547 738 -2547 0 cellNo=519
rlabel pdiffusion 745 -2547 745 -2547 0 cellNo=427
rlabel pdiffusion 752 -2547 752 -2547 0 feedthrough
rlabel pdiffusion 759 -2547 759 -2547 0 feedthrough
rlabel pdiffusion 766 -2547 766 -2547 0 feedthrough
rlabel pdiffusion 773 -2547 773 -2547 0 feedthrough
rlabel pdiffusion 780 -2547 780 -2547 0 feedthrough
rlabel pdiffusion 787 -2547 787 -2547 0 feedthrough
rlabel pdiffusion 794 -2547 794 -2547 0 feedthrough
rlabel pdiffusion 801 -2547 801 -2547 0 feedthrough
rlabel pdiffusion 808 -2547 808 -2547 0 cellNo=584
rlabel pdiffusion 829 -2547 829 -2547 0 feedthrough
rlabel pdiffusion 864 -2547 864 -2547 0 cellNo=561
rlabel pdiffusion 871 -2547 871 -2547 0 feedthrough
rlabel pdiffusion 913 -2547 913 -2547 0 feedthrough
rlabel pdiffusion 927 -2547 927 -2547 0 feedthrough
rlabel pdiffusion 934 -2547 934 -2547 0 feedthrough
rlabel pdiffusion 948 -2547 948 -2547 0 feedthrough
rlabel pdiffusion 955 -2547 955 -2547 0 feedthrough
rlabel pdiffusion 976 -2547 976 -2547 0 feedthrough
rlabel pdiffusion 1018 -2547 1018 -2547 0 feedthrough
rlabel pdiffusion 1032 -2547 1032 -2547 0 feedthrough
rlabel pdiffusion 1039 -2547 1039 -2547 0 feedthrough
rlabel pdiffusion 1053 -2547 1053 -2547 0 feedthrough
rlabel pdiffusion 1067 -2547 1067 -2547 0 feedthrough
rlabel pdiffusion 1095 -2547 1095 -2547 0 cellNo=425
rlabel pdiffusion 1144 -2547 1144 -2547 0 feedthrough
rlabel pdiffusion 1179 -2547 1179 -2547 0 cellNo=288
rlabel pdiffusion 1186 -2547 1186 -2547 0 feedthrough
rlabel pdiffusion 129 -2592 129 -2592 0 cellNo=68
rlabel pdiffusion 136 -2592 136 -2592 0 feedthrough
rlabel pdiffusion 255 -2592 255 -2592 0 cellNo=256
rlabel pdiffusion 325 -2592 325 -2592 0 feedthrough
rlabel pdiffusion 332 -2592 332 -2592 0 feedthrough
rlabel pdiffusion 339 -2592 339 -2592 0 feedthrough
rlabel pdiffusion 346 -2592 346 -2592 0 cellNo=343
rlabel pdiffusion 367 -2592 367 -2592 0 feedthrough
rlabel pdiffusion 374 -2592 374 -2592 0 cellNo=347
rlabel pdiffusion 381 -2592 381 -2592 0 cellNo=600
rlabel pdiffusion 444 -2592 444 -2592 0 feedthrough
rlabel pdiffusion 451 -2592 451 -2592 0 feedthrough
rlabel pdiffusion 472 -2592 472 -2592 0 feedthrough
rlabel pdiffusion 493 -2592 493 -2592 0 feedthrough
rlabel pdiffusion 500 -2592 500 -2592 0 feedthrough
rlabel pdiffusion 507 -2592 507 -2592 0 feedthrough
rlabel pdiffusion 514 -2592 514 -2592 0 cellNo=251
rlabel pdiffusion 528 -2592 528 -2592 0 cellNo=585
rlabel pdiffusion 535 -2592 535 -2592 0 feedthrough
rlabel pdiffusion 542 -2592 542 -2592 0 cellNo=303
rlabel pdiffusion 549 -2592 549 -2592 0 cellNo=269
rlabel pdiffusion 556 -2592 556 -2592 0 feedthrough
rlabel pdiffusion 563 -2592 563 -2592 0 cellNo=494
rlabel pdiffusion 570 -2592 570 -2592 0 feedthrough
rlabel pdiffusion 577 -2592 577 -2592 0 feedthrough
rlabel pdiffusion 598 -2592 598 -2592 0 cellNo=418
rlabel pdiffusion 647 -2592 647 -2592 0 cellNo=199
rlabel pdiffusion 661 -2592 661 -2592 0 cellNo=392
rlabel pdiffusion 668 -2592 668 -2592 0 feedthrough
rlabel pdiffusion 675 -2592 675 -2592 0 cellNo=143
rlabel pdiffusion 682 -2592 682 -2592 0 cellNo=557
rlabel pdiffusion 689 -2592 689 -2592 0 cellNo=447
rlabel pdiffusion 710 -2592 710 -2592 0 cellNo=229
rlabel pdiffusion 717 -2592 717 -2592 0 feedthrough
rlabel pdiffusion 724 -2592 724 -2592 0 feedthrough
rlabel pdiffusion 731 -2592 731 -2592 0 feedthrough
rlabel pdiffusion 752 -2592 752 -2592 0 feedthrough
rlabel pdiffusion 808 -2592 808 -2592 0 cellNo=479
rlabel pdiffusion 815 -2592 815 -2592 0 feedthrough
rlabel pdiffusion 885 -2592 885 -2592 0 cellNo=588
rlabel pdiffusion 899 -2592 899 -2592 0 feedthrough
rlabel pdiffusion 955 -2592 955 -2592 0 feedthrough
rlabel pdiffusion 962 -2592 962 -2592 0 cellNo=571
rlabel pdiffusion 969 -2592 969 -2592 0 feedthrough
rlabel pdiffusion 1011 -2592 1011 -2592 0 cellNo=492
rlabel pdiffusion 1018 -2592 1018 -2592 0 feedthrough
rlabel pdiffusion 1025 -2592 1025 -2592 0 feedthrough
rlabel pdiffusion 1046 -2592 1046 -2592 0 feedthrough
rlabel pdiffusion 1053 -2592 1053 -2592 0 cellNo=47
rlabel pdiffusion 1060 -2592 1060 -2592 0 feedthrough
rlabel polysilicon 156 -22 156 -22 0 3
rlabel polysilicon 215 -16 215 -16 0 2
rlabel polysilicon 215 -22 215 -22 0 4
rlabel polysilicon 240 -16 240 -16 0 1
rlabel polysilicon 240 -22 240 -22 0 3
rlabel polysilicon 247 -16 247 -16 0 1
rlabel polysilicon 247 -22 247 -22 0 3
rlabel polysilicon 261 -16 261 -16 0 1
rlabel polysilicon 261 -22 261 -22 0 3
rlabel polysilicon 268 -16 268 -16 0 1
rlabel polysilicon 275 -16 275 -16 0 1
rlabel polysilicon 275 -22 275 -22 0 3
rlabel polysilicon 282 -22 282 -22 0 3
rlabel polysilicon 285 -22 285 -22 0 4
rlabel polysilicon 338 -16 338 -16 0 1
rlabel polysilicon 338 -22 338 -22 0 3
rlabel polysilicon 373 -16 373 -16 0 1
rlabel polysilicon 373 -22 373 -22 0 3
rlabel polysilicon 380 -16 380 -16 0 1
rlabel polysilicon 380 -22 380 -22 0 3
rlabel polysilicon 383 -22 383 -22 0 4
rlabel polysilicon 387 -16 387 -16 0 1
rlabel polysilicon 387 -22 387 -22 0 3
rlabel polysilicon 397 -16 397 -16 0 2
rlabel polysilicon 397 -22 397 -22 0 4
rlabel polysilicon 401 -16 401 -16 0 1
rlabel polysilicon 401 -22 401 -22 0 3
rlabel polysilicon 404 -22 404 -22 0 4
rlabel polysilicon 408 -16 408 -16 0 1
rlabel polysilicon 411 -16 411 -16 0 2
rlabel polysilicon 408 -22 408 -22 0 3
rlabel polysilicon 415 -16 415 -16 0 1
rlabel polysilicon 415 -22 415 -22 0 3
rlabel polysilicon 425 -16 425 -16 0 2
rlabel polysilicon 425 -22 425 -22 0 4
rlabel polysilicon 429 -16 429 -16 0 1
rlabel polysilicon 429 -22 429 -22 0 3
rlabel polysilicon 457 -16 457 -16 0 1
rlabel polysilicon 457 -22 457 -22 0 3
rlabel polysilicon 460 -22 460 -22 0 4
rlabel polysilicon 464 -16 464 -16 0 1
rlabel polysilicon 467 -16 467 -16 0 2
rlabel polysilicon 467 -22 467 -22 0 4
rlabel polysilicon 478 -16 478 -16 0 1
rlabel polysilicon 478 -22 478 -22 0 3
rlabel polysilicon 481 -22 481 -22 0 4
rlabel polysilicon 485 -16 485 -16 0 1
rlabel polysilicon 485 -22 485 -22 0 3
rlabel polysilicon 499 -16 499 -16 0 1
rlabel polysilicon 499 -22 499 -22 0 3
rlabel polysilicon 506 -16 506 -16 0 1
rlabel polysilicon 506 -22 506 -22 0 3
rlabel polysilicon 516 -16 516 -16 0 2
rlabel polysilicon 513 -22 513 -22 0 3
rlabel polysilicon 516 -22 516 -22 0 4
rlabel polysilicon 527 -16 527 -16 0 1
rlabel polysilicon 527 -22 527 -22 0 3
rlabel polysilicon 548 -22 548 -22 0 3
rlabel polysilicon 551 -22 551 -22 0 4
rlabel polysilicon 562 -16 562 -16 0 1
rlabel polysilicon 562 -22 562 -22 0 3
rlabel polysilicon 569 -16 569 -16 0 1
rlabel polysilicon 569 -22 569 -22 0 3
rlabel polysilicon 576 -16 576 -16 0 1
rlabel polysilicon 576 -22 576 -22 0 3
rlabel polysilicon 583 -16 583 -16 0 1
rlabel polysilicon 586 -16 586 -16 0 2
rlabel polysilicon 583 -22 583 -22 0 3
rlabel polysilicon 604 -16 604 -16 0 1
rlabel polysilicon 607 -16 607 -16 0 2
rlabel polysilicon 607 -22 607 -22 0 4
rlabel polysilicon 639 -16 639 -16 0 1
rlabel polysilicon 639 -22 639 -22 0 3
rlabel polysilicon 667 -16 667 -16 0 1
rlabel polysilicon 667 -22 667 -22 0 3
rlabel polysilicon 681 -16 681 -16 0 1
rlabel polysilicon 681 -22 681 -22 0 3
rlabel polysilicon 702 -16 702 -16 0 1
rlabel polysilicon 702 -22 702 -22 0 3
rlabel polysilicon 709 -16 709 -16 0 1
rlabel polysilicon 709 -22 709 -22 0 3
rlabel polysilicon 765 -16 765 -16 0 1
rlabel polysilicon 765 -22 765 -22 0 3
rlabel polysilicon 800 -16 800 -16 0 1
rlabel polysilicon 803 -16 803 -16 0 2
rlabel polysilicon 800 -22 800 -22 0 3
rlabel polysilicon 828 -16 828 -16 0 1
rlabel polysilicon 828 -22 828 -22 0 3
rlabel polysilicon 149 -65 149 -65 0 3
rlabel polysilicon 152 -65 152 -65 0 4
rlabel polysilicon 156 -59 156 -59 0 1
rlabel polysilicon 159 -65 159 -65 0 4
rlabel polysilicon 163 -59 163 -59 0 1
rlabel polysilicon 163 -65 163 -65 0 3
rlabel polysilicon 191 -59 191 -59 0 1
rlabel polysilicon 191 -65 191 -65 0 3
rlabel polysilicon 219 -59 219 -59 0 1
rlabel polysilicon 219 -65 219 -65 0 3
rlabel polysilicon 226 -59 226 -59 0 1
rlabel polysilicon 226 -65 226 -65 0 3
rlabel polysilicon 233 -59 233 -59 0 1
rlabel polysilicon 233 -65 233 -65 0 3
rlabel polysilicon 247 -59 247 -59 0 1
rlabel polysilicon 247 -65 247 -65 0 3
rlabel polysilicon 254 -59 254 -59 0 1
rlabel polysilicon 254 -65 254 -65 0 3
rlabel polysilicon 261 -59 261 -59 0 1
rlabel polysilicon 261 -65 261 -65 0 3
rlabel polysilicon 268 -59 268 -59 0 1
rlabel polysilicon 268 -65 268 -65 0 3
rlabel polysilicon 275 -59 275 -59 0 1
rlabel polysilicon 275 -65 275 -65 0 3
rlabel polysilicon 282 -59 282 -59 0 1
rlabel polysilicon 282 -65 282 -65 0 3
rlabel polysilicon 292 -59 292 -59 0 2
rlabel polysilicon 289 -65 289 -65 0 3
rlabel polysilicon 292 -65 292 -65 0 4
rlabel polysilicon 296 -59 296 -59 0 1
rlabel polysilicon 296 -65 296 -65 0 3
rlabel polysilicon 303 -59 303 -59 0 1
rlabel polysilicon 303 -65 303 -65 0 3
rlabel polysilicon 310 -59 310 -59 0 1
rlabel polysilicon 310 -65 310 -65 0 3
rlabel polysilicon 317 -59 317 -59 0 1
rlabel polysilicon 317 -65 317 -65 0 3
rlabel polysilicon 324 -59 324 -59 0 1
rlabel polysilicon 324 -65 324 -65 0 3
rlabel polysilicon 331 -59 331 -59 0 1
rlabel polysilicon 331 -65 331 -65 0 3
rlabel polysilicon 338 -65 338 -65 0 3
rlabel polysilicon 341 -65 341 -65 0 4
rlabel polysilicon 345 -59 345 -59 0 1
rlabel polysilicon 345 -65 345 -65 0 3
rlabel polysilicon 348 -65 348 -65 0 4
rlabel polysilicon 355 -59 355 -59 0 2
rlabel polysilicon 352 -65 352 -65 0 3
rlabel polysilicon 355 -65 355 -65 0 4
rlabel polysilicon 359 -59 359 -59 0 1
rlabel polysilicon 359 -65 359 -65 0 3
rlabel polysilicon 366 -59 366 -59 0 1
rlabel polysilicon 366 -65 366 -65 0 3
rlabel polysilicon 373 -59 373 -59 0 1
rlabel polysilicon 373 -65 373 -65 0 3
rlabel polysilicon 380 -59 380 -59 0 1
rlabel polysilicon 383 -65 383 -65 0 4
rlabel polysilicon 387 -59 387 -59 0 1
rlabel polysilicon 387 -65 387 -65 0 3
rlabel polysilicon 394 -59 394 -59 0 1
rlabel polysilicon 394 -65 394 -65 0 3
rlabel polysilicon 401 -59 401 -59 0 1
rlabel polysilicon 401 -65 401 -65 0 3
rlabel polysilicon 411 -59 411 -59 0 2
rlabel polysilicon 411 -65 411 -65 0 4
rlabel polysilicon 418 -59 418 -59 0 2
rlabel polysilicon 415 -65 415 -65 0 3
rlabel polysilicon 418 -65 418 -65 0 4
rlabel polysilicon 422 -59 422 -59 0 1
rlabel polysilicon 422 -65 422 -65 0 3
rlabel polysilicon 429 -59 429 -59 0 1
rlabel polysilicon 429 -65 429 -65 0 3
rlabel polysilicon 436 -59 436 -59 0 1
rlabel polysilicon 436 -65 436 -65 0 3
rlabel polysilicon 443 -59 443 -59 0 1
rlabel polysilicon 443 -65 443 -65 0 3
rlabel polysilicon 450 -65 450 -65 0 3
rlabel polysilicon 453 -65 453 -65 0 4
rlabel polysilicon 457 -59 457 -59 0 1
rlabel polysilicon 457 -65 457 -65 0 3
rlabel polysilicon 464 -59 464 -59 0 1
rlabel polysilicon 464 -65 464 -65 0 3
rlabel polysilicon 471 -59 471 -59 0 1
rlabel polysilicon 471 -65 471 -65 0 3
rlabel polysilicon 478 -59 478 -59 0 1
rlabel polysilicon 478 -65 478 -65 0 3
rlabel polysilicon 481 -65 481 -65 0 4
rlabel polysilicon 485 -59 485 -59 0 1
rlabel polysilicon 485 -65 485 -65 0 3
rlabel polysilicon 492 -59 492 -59 0 1
rlabel polysilicon 492 -65 492 -65 0 3
rlabel polysilicon 499 -59 499 -59 0 1
rlabel polysilicon 502 -59 502 -59 0 2
rlabel polysilicon 499 -65 499 -65 0 3
rlabel polysilicon 506 -59 506 -59 0 1
rlabel polysilicon 506 -65 506 -65 0 3
rlabel polysilicon 513 -59 513 -59 0 1
rlabel polysilicon 513 -65 513 -65 0 3
rlabel polysilicon 520 -59 520 -59 0 1
rlabel polysilicon 520 -65 520 -65 0 3
rlabel polysilicon 527 -59 527 -59 0 1
rlabel polysilicon 527 -65 527 -65 0 3
rlabel polysilicon 534 -59 534 -59 0 1
rlabel polysilicon 537 -59 537 -59 0 2
rlabel polysilicon 537 -65 537 -65 0 4
rlabel polysilicon 541 -59 541 -59 0 1
rlabel polysilicon 541 -65 541 -65 0 3
rlabel polysilicon 548 -59 548 -59 0 1
rlabel polysilicon 548 -65 548 -65 0 3
rlabel polysilicon 555 -59 555 -59 0 1
rlabel polysilicon 555 -65 555 -65 0 3
rlabel polysilicon 558 -65 558 -65 0 4
rlabel polysilicon 562 -59 562 -59 0 1
rlabel polysilicon 562 -65 562 -65 0 3
rlabel polysilicon 569 -59 569 -59 0 1
rlabel polysilicon 569 -65 569 -65 0 3
rlabel polysilicon 579 -59 579 -59 0 2
rlabel polysilicon 576 -65 576 -65 0 3
rlabel polysilicon 579 -65 579 -65 0 4
rlabel polysilicon 583 -59 583 -59 0 1
rlabel polysilicon 583 -65 583 -65 0 3
rlabel polysilicon 593 -59 593 -59 0 2
rlabel polysilicon 590 -65 590 -65 0 3
rlabel polysilicon 593 -65 593 -65 0 4
rlabel polysilicon 597 -59 597 -59 0 1
rlabel polysilicon 597 -65 597 -65 0 3
rlabel polysilicon 604 -59 604 -59 0 1
rlabel polysilicon 604 -65 604 -65 0 3
rlabel polysilicon 611 -59 611 -59 0 1
rlabel polysilicon 611 -65 611 -65 0 3
rlabel polysilicon 618 -59 618 -59 0 1
rlabel polysilicon 621 -59 621 -59 0 2
rlabel polysilicon 618 -65 618 -65 0 3
rlabel polysilicon 625 -59 625 -59 0 1
rlabel polysilicon 625 -65 625 -65 0 3
rlabel polysilicon 632 -59 632 -59 0 1
rlabel polysilicon 632 -65 632 -65 0 3
rlabel polysilicon 639 -59 639 -59 0 1
rlabel polysilicon 639 -65 639 -65 0 3
rlabel polysilicon 646 -59 646 -59 0 1
rlabel polysilicon 646 -65 646 -65 0 3
rlabel polysilicon 653 -59 653 -59 0 1
rlabel polysilicon 653 -65 653 -65 0 3
rlabel polysilicon 660 -59 660 -59 0 1
rlabel polysilicon 660 -65 660 -65 0 3
rlabel polysilicon 667 -59 667 -59 0 1
rlabel polysilicon 670 -65 670 -65 0 4
rlabel polysilicon 674 -59 674 -59 0 1
rlabel polysilicon 674 -65 674 -65 0 3
rlabel polysilicon 681 -59 681 -59 0 1
rlabel polysilicon 681 -65 681 -65 0 3
rlabel polysilicon 688 -59 688 -59 0 1
rlabel polysilicon 688 -65 688 -65 0 3
rlabel polysilicon 702 -59 702 -59 0 1
rlabel polysilicon 702 -65 702 -65 0 3
rlabel polysilicon 716 -59 716 -59 0 1
rlabel polysilicon 719 -59 719 -59 0 2
rlabel polysilicon 719 -65 719 -65 0 4
rlabel polysilicon 723 -59 723 -59 0 1
rlabel polysilicon 723 -65 723 -65 0 3
rlabel polysilicon 751 -59 751 -59 0 1
rlabel polysilicon 751 -65 751 -65 0 3
rlabel polysilicon 758 -59 758 -59 0 1
rlabel polysilicon 758 -65 758 -65 0 3
rlabel polysilicon 772 -59 772 -59 0 1
rlabel polysilicon 772 -65 772 -65 0 3
rlabel polysilicon 828 -59 828 -59 0 1
rlabel polysilicon 828 -65 828 -65 0 3
rlabel polysilicon 849 -59 849 -59 0 1
rlabel polysilicon 849 -65 849 -65 0 3
rlabel polysilicon 877 -59 877 -59 0 1
rlabel polysilicon 877 -65 877 -65 0 3
rlabel polysilicon 905 -59 905 -59 0 1
rlabel polysilicon 905 -65 905 -65 0 3
rlabel polysilicon 23 -120 23 -120 0 1
rlabel polysilicon 23 -126 23 -126 0 3
rlabel polysilicon 30 -120 30 -120 0 1
rlabel polysilicon 30 -126 30 -126 0 3
rlabel polysilicon 37 -120 37 -120 0 1
rlabel polysilicon 37 -126 37 -126 0 3
rlabel polysilicon 44 -120 44 -120 0 1
rlabel polysilicon 44 -126 44 -126 0 3
rlabel polysilicon 51 -120 51 -120 0 1
rlabel polysilicon 51 -126 51 -126 0 3
rlabel polysilicon 58 -126 58 -126 0 3
rlabel polysilicon 61 -126 61 -126 0 4
rlabel polysilicon 65 -120 65 -120 0 1
rlabel polysilicon 68 -126 68 -126 0 4
rlabel polysilicon 75 -120 75 -120 0 2
rlabel polysilicon 75 -126 75 -126 0 4
rlabel polysilicon 79 -120 79 -120 0 1
rlabel polysilicon 79 -126 79 -126 0 3
rlabel polysilicon 86 -120 86 -120 0 1
rlabel polysilicon 89 -120 89 -120 0 2
rlabel polysilicon 89 -126 89 -126 0 4
rlabel polysilicon 93 -120 93 -120 0 1
rlabel polysilicon 93 -126 93 -126 0 3
rlabel polysilicon 100 -120 100 -120 0 1
rlabel polysilicon 100 -126 100 -126 0 3
rlabel polysilicon 107 -120 107 -120 0 1
rlabel polysilicon 107 -126 107 -126 0 3
rlabel polysilicon 114 -120 114 -120 0 1
rlabel polysilicon 117 -120 117 -120 0 2
rlabel polysilicon 117 -126 117 -126 0 4
rlabel polysilicon 121 -120 121 -120 0 1
rlabel polysilicon 121 -126 121 -126 0 3
rlabel polysilicon 128 -120 128 -120 0 1
rlabel polysilicon 131 -126 131 -126 0 4
rlabel polysilicon 135 -120 135 -120 0 1
rlabel polysilicon 135 -126 135 -126 0 3
rlabel polysilicon 142 -120 142 -120 0 1
rlabel polysilicon 142 -126 142 -126 0 3
rlabel polysilicon 149 -120 149 -120 0 1
rlabel polysilicon 149 -126 149 -126 0 3
rlabel polysilicon 156 -120 156 -120 0 1
rlabel polysilicon 156 -126 156 -126 0 3
rlabel polysilicon 163 -120 163 -120 0 1
rlabel polysilicon 163 -126 163 -126 0 3
rlabel polysilicon 170 -120 170 -120 0 1
rlabel polysilicon 170 -126 170 -126 0 3
rlabel polysilicon 177 -120 177 -120 0 1
rlabel polysilicon 177 -126 177 -126 0 3
rlabel polysilicon 184 -120 184 -120 0 1
rlabel polysilicon 187 -120 187 -120 0 2
rlabel polysilicon 187 -126 187 -126 0 4
rlabel polysilicon 194 -120 194 -120 0 2
rlabel polysilicon 191 -126 191 -126 0 3
rlabel polysilicon 194 -126 194 -126 0 4
rlabel polysilicon 198 -120 198 -120 0 1
rlabel polysilicon 198 -126 198 -126 0 3
rlabel polysilicon 205 -120 205 -120 0 1
rlabel polysilicon 205 -126 205 -126 0 3
rlabel polysilicon 212 -120 212 -120 0 1
rlabel polysilicon 212 -126 212 -126 0 3
rlabel polysilicon 219 -120 219 -120 0 1
rlabel polysilicon 219 -126 219 -126 0 3
rlabel polysilicon 226 -120 226 -120 0 1
rlabel polysilicon 226 -126 226 -126 0 3
rlabel polysilicon 233 -120 233 -120 0 1
rlabel polysilicon 233 -126 233 -126 0 3
rlabel polysilicon 240 -120 240 -120 0 1
rlabel polysilicon 240 -126 240 -126 0 3
rlabel polysilicon 247 -120 247 -120 0 1
rlabel polysilicon 247 -126 247 -126 0 3
rlabel polysilicon 254 -120 254 -120 0 1
rlabel polysilicon 254 -126 254 -126 0 3
rlabel polysilicon 261 -120 261 -120 0 1
rlabel polysilicon 261 -126 261 -126 0 3
rlabel polysilicon 268 -120 268 -120 0 1
rlabel polysilicon 271 -120 271 -120 0 2
rlabel polysilicon 268 -126 268 -126 0 3
rlabel polysilicon 271 -126 271 -126 0 4
rlabel polysilicon 275 -120 275 -120 0 1
rlabel polysilicon 275 -126 275 -126 0 3
rlabel polysilicon 282 -120 282 -120 0 1
rlabel polysilicon 282 -126 282 -126 0 3
rlabel polysilicon 289 -120 289 -120 0 1
rlabel polysilicon 289 -126 289 -126 0 3
rlabel polysilicon 299 -120 299 -120 0 2
rlabel polysilicon 296 -126 296 -126 0 3
rlabel polysilicon 299 -126 299 -126 0 4
rlabel polysilicon 303 -120 303 -120 0 1
rlabel polysilicon 303 -126 303 -126 0 3
rlabel polysilicon 310 -120 310 -120 0 1
rlabel polysilicon 313 -120 313 -120 0 2
rlabel polysilicon 310 -126 310 -126 0 3
rlabel polysilicon 317 -120 317 -120 0 1
rlabel polysilicon 317 -126 317 -126 0 3
rlabel polysilicon 327 -120 327 -120 0 2
rlabel polysilicon 324 -126 324 -126 0 3
rlabel polysilicon 327 -126 327 -126 0 4
rlabel polysilicon 331 -120 331 -120 0 1
rlabel polysilicon 331 -126 331 -126 0 3
rlabel polysilicon 338 -120 338 -120 0 1
rlabel polysilicon 338 -126 338 -126 0 3
rlabel polysilicon 345 -120 345 -120 0 1
rlabel polysilicon 345 -126 345 -126 0 3
rlabel polysilicon 352 -120 352 -120 0 1
rlabel polysilicon 352 -126 352 -126 0 3
rlabel polysilicon 359 -120 359 -120 0 1
rlabel polysilicon 362 -126 362 -126 0 4
rlabel polysilicon 366 -120 366 -120 0 1
rlabel polysilicon 366 -126 366 -126 0 3
rlabel polysilicon 373 -120 373 -120 0 1
rlabel polysilicon 373 -126 373 -126 0 3
rlabel polysilicon 380 -120 380 -120 0 1
rlabel polysilicon 380 -126 380 -126 0 3
rlabel polysilicon 387 -120 387 -120 0 1
rlabel polysilicon 387 -126 387 -126 0 3
rlabel polysilicon 394 -120 394 -120 0 1
rlabel polysilicon 397 -120 397 -120 0 2
rlabel polysilicon 397 -126 397 -126 0 4
rlabel polysilicon 401 -120 401 -120 0 1
rlabel polysilicon 404 -120 404 -120 0 2
rlabel polysilicon 401 -126 401 -126 0 3
rlabel polysilicon 408 -120 408 -120 0 1
rlabel polysilicon 408 -126 408 -126 0 3
rlabel polysilicon 415 -120 415 -120 0 1
rlabel polysilicon 415 -126 415 -126 0 3
rlabel polysilicon 422 -120 422 -120 0 1
rlabel polysilicon 422 -126 422 -126 0 3
rlabel polysilicon 429 -120 429 -120 0 1
rlabel polysilicon 429 -126 429 -126 0 3
rlabel polysilicon 436 -120 436 -120 0 1
rlabel polysilicon 439 -120 439 -120 0 2
rlabel polysilicon 436 -126 436 -126 0 3
rlabel polysilicon 439 -126 439 -126 0 4
rlabel polysilicon 443 -120 443 -120 0 1
rlabel polysilicon 443 -126 443 -126 0 3
rlabel polysilicon 450 -120 450 -120 0 1
rlabel polysilicon 450 -126 450 -126 0 3
rlabel polysilicon 457 -120 457 -120 0 1
rlabel polysilicon 457 -126 457 -126 0 3
rlabel polysilicon 464 -120 464 -120 0 1
rlabel polysilicon 464 -126 464 -126 0 3
rlabel polysilicon 471 -120 471 -120 0 1
rlabel polysilicon 471 -126 471 -126 0 3
rlabel polysilicon 478 -120 478 -120 0 1
rlabel polysilicon 478 -126 478 -126 0 3
rlabel polysilicon 485 -120 485 -120 0 1
rlabel polysilicon 485 -126 485 -126 0 3
rlabel polysilicon 492 -120 492 -120 0 1
rlabel polysilicon 492 -126 492 -126 0 3
rlabel polysilicon 499 -120 499 -120 0 1
rlabel polysilicon 499 -126 499 -126 0 3
rlabel polysilicon 506 -120 506 -120 0 1
rlabel polysilicon 506 -126 506 -126 0 3
rlabel polysilicon 513 -120 513 -120 0 1
rlabel polysilicon 513 -126 513 -126 0 3
rlabel polysilicon 520 -120 520 -120 0 1
rlabel polysilicon 520 -126 520 -126 0 3
rlabel polysilicon 530 -120 530 -120 0 2
rlabel polysilicon 527 -126 527 -126 0 3
rlabel polysilicon 530 -126 530 -126 0 4
rlabel polysilicon 534 -120 534 -120 0 1
rlabel polysilicon 534 -126 534 -126 0 3
rlabel polysilicon 541 -120 541 -120 0 1
rlabel polysilicon 541 -126 541 -126 0 3
rlabel polysilicon 548 -120 548 -120 0 1
rlabel polysilicon 548 -126 548 -126 0 3
rlabel polysilicon 555 -120 555 -120 0 1
rlabel polysilicon 555 -126 555 -126 0 3
rlabel polysilicon 562 -120 562 -120 0 1
rlabel polysilicon 562 -126 562 -126 0 3
rlabel polysilicon 569 -120 569 -120 0 1
rlabel polysilicon 569 -126 569 -126 0 3
rlabel polysilicon 576 -120 576 -120 0 1
rlabel polysilicon 576 -126 576 -126 0 3
rlabel polysilicon 583 -120 583 -120 0 1
rlabel polysilicon 583 -126 583 -126 0 3
rlabel polysilicon 590 -120 590 -120 0 1
rlabel polysilicon 590 -126 590 -126 0 3
rlabel polysilicon 597 -120 597 -120 0 1
rlabel polysilicon 597 -126 597 -126 0 3
rlabel polysilicon 604 -120 604 -120 0 1
rlabel polysilicon 607 -120 607 -120 0 2
rlabel polysilicon 607 -126 607 -126 0 4
rlabel polysilicon 611 -120 611 -120 0 1
rlabel polysilicon 611 -126 611 -126 0 3
rlabel polysilicon 618 -120 618 -120 0 1
rlabel polysilicon 618 -126 618 -126 0 3
rlabel polysilicon 625 -120 625 -120 0 1
rlabel polysilicon 625 -126 625 -126 0 3
rlabel polysilicon 632 -120 632 -120 0 1
rlabel polysilicon 632 -126 632 -126 0 3
rlabel polysilicon 639 -120 639 -120 0 1
rlabel polysilicon 639 -126 639 -126 0 3
rlabel polysilicon 646 -120 646 -120 0 1
rlabel polysilicon 646 -126 646 -126 0 3
rlabel polysilicon 653 -120 653 -120 0 1
rlabel polysilicon 653 -126 653 -126 0 3
rlabel polysilicon 660 -120 660 -120 0 1
rlabel polysilicon 663 -120 663 -120 0 2
rlabel polysilicon 663 -126 663 -126 0 4
rlabel polysilicon 667 -120 667 -120 0 1
rlabel polysilicon 667 -126 667 -126 0 3
rlabel polysilicon 674 -120 674 -120 0 1
rlabel polysilicon 674 -126 674 -126 0 3
rlabel polysilicon 681 -120 681 -120 0 1
rlabel polysilicon 681 -126 681 -126 0 3
rlabel polysilicon 688 -120 688 -120 0 1
rlabel polysilicon 688 -126 688 -126 0 3
rlabel polysilicon 695 -120 695 -120 0 1
rlabel polysilicon 695 -126 695 -126 0 3
rlabel polysilicon 702 -120 702 -120 0 1
rlabel polysilicon 702 -126 702 -126 0 3
rlabel polysilicon 709 -120 709 -120 0 1
rlabel polysilicon 709 -126 709 -126 0 3
rlabel polysilicon 716 -120 716 -120 0 1
rlabel polysilicon 716 -126 716 -126 0 3
rlabel polysilicon 723 -120 723 -120 0 1
rlabel polysilicon 723 -126 723 -126 0 3
rlabel polysilicon 730 -120 730 -120 0 1
rlabel polysilicon 730 -126 730 -126 0 3
rlabel polysilicon 737 -120 737 -120 0 1
rlabel polysilicon 737 -126 737 -126 0 3
rlabel polysilicon 744 -120 744 -120 0 1
rlabel polysilicon 744 -126 744 -126 0 3
rlabel polysilicon 751 -120 751 -120 0 1
rlabel polysilicon 751 -126 751 -126 0 3
rlabel polysilicon 761 -120 761 -120 0 2
rlabel polysilicon 765 -120 765 -120 0 1
rlabel polysilicon 765 -126 765 -126 0 3
rlabel polysilicon 772 -120 772 -120 0 1
rlabel polysilicon 772 -126 772 -126 0 3
rlabel polysilicon 779 -120 779 -120 0 1
rlabel polysilicon 779 -126 779 -126 0 3
rlabel polysilicon 786 -120 786 -120 0 1
rlabel polysilicon 786 -126 786 -126 0 3
rlabel polysilicon 793 -120 793 -120 0 1
rlabel polysilicon 793 -126 793 -126 0 3
rlabel polysilicon 800 -120 800 -120 0 1
rlabel polysilicon 800 -126 800 -126 0 3
rlabel polysilicon 807 -120 807 -120 0 1
rlabel polysilicon 807 -126 807 -126 0 3
rlabel polysilicon 814 -120 814 -120 0 1
rlabel polysilicon 814 -126 814 -126 0 3
rlabel polysilicon 821 -120 821 -120 0 1
rlabel polysilicon 821 -126 821 -126 0 3
rlabel polysilicon 849 -120 849 -120 0 1
rlabel polysilicon 849 -126 849 -126 0 3
rlabel polysilicon 856 -120 856 -120 0 1
rlabel polysilicon 856 -126 856 -126 0 3
rlabel polysilicon 870 -120 870 -120 0 1
rlabel polysilicon 870 -126 870 -126 0 3
rlabel polysilicon 877 -120 877 -120 0 1
rlabel polysilicon 877 -126 877 -126 0 3
rlabel polysilicon 940 -120 940 -120 0 1
rlabel polysilicon 940 -126 940 -126 0 3
rlabel polysilicon 947 -120 947 -120 0 1
rlabel polysilicon 947 -126 947 -126 0 3
rlabel polysilicon 1500 -120 1500 -120 0 1
rlabel polysilicon 1500 -126 1500 -126 0 3
rlabel polysilicon 1507 -120 1507 -120 0 1
rlabel polysilicon 9 -199 9 -199 0 1
rlabel polysilicon 9 -205 9 -205 0 3
rlabel polysilicon 16 -199 16 -199 0 1
rlabel polysilicon 16 -205 16 -205 0 3
rlabel polysilicon 23 -199 23 -199 0 1
rlabel polysilicon 23 -205 23 -205 0 3
rlabel polysilicon 30 -199 30 -199 0 1
rlabel polysilicon 30 -205 30 -205 0 3
rlabel polysilicon 37 -199 37 -199 0 1
rlabel polysilicon 37 -205 37 -205 0 3
rlabel polysilicon 44 -199 44 -199 0 1
rlabel polysilicon 44 -205 44 -205 0 3
rlabel polysilicon 51 -199 51 -199 0 1
rlabel polysilicon 54 -199 54 -199 0 2
rlabel polysilicon 51 -205 51 -205 0 3
rlabel polysilicon 54 -205 54 -205 0 4
rlabel polysilicon 58 -199 58 -199 0 1
rlabel polysilicon 58 -205 58 -205 0 3
rlabel polysilicon 65 -199 65 -199 0 1
rlabel polysilicon 65 -205 65 -205 0 3
rlabel polysilicon 72 -199 72 -199 0 1
rlabel polysilicon 72 -205 72 -205 0 3
rlabel polysilicon 79 -199 79 -199 0 1
rlabel polysilicon 79 -205 79 -205 0 3
rlabel polysilicon 86 -199 86 -199 0 1
rlabel polysilicon 86 -205 86 -205 0 3
rlabel polysilicon 93 -199 93 -199 0 1
rlabel polysilicon 93 -205 93 -205 0 3
rlabel polysilicon 100 -199 100 -199 0 1
rlabel polysilicon 103 -199 103 -199 0 2
rlabel polysilicon 103 -205 103 -205 0 4
rlabel polysilicon 107 -199 107 -199 0 1
rlabel polysilicon 107 -205 107 -205 0 3
rlabel polysilicon 114 -199 114 -199 0 1
rlabel polysilicon 114 -205 114 -205 0 3
rlabel polysilicon 121 -199 121 -199 0 1
rlabel polysilicon 121 -205 121 -205 0 3
rlabel polysilicon 128 -199 128 -199 0 1
rlabel polysilicon 128 -205 128 -205 0 3
rlabel polysilicon 135 -199 135 -199 0 1
rlabel polysilicon 135 -205 135 -205 0 3
rlabel polysilicon 142 -199 142 -199 0 1
rlabel polysilicon 145 -199 145 -199 0 2
rlabel polysilicon 142 -205 142 -205 0 3
rlabel polysilicon 149 -199 149 -199 0 1
rlabel polysilicon 152 -199 152 -199 0 2
rlabel polysilicon 149 -205 149 -205 0 3
rlabel polysilicon 156 -199 156 -199 0 1
rlabel polysilicon 156 -205 156 -205 0 3
rlabel polysilicon 159 -205 159 -205 0 4
rlabel polysilicon 163 -199 163 -199 0 1
rlabel polysilicon 163 -205 163 -205 0 3
rlabel polysilicon 170 -199 170 -199 0 1
rlabel polysilicon 170 -205 170 -205 0 3
rlabel polysilicon 177 -199 177 -199 0 1
rlabel polysilicon 177 -205 177 -205 0 3
rlabel polysilicon 184 -199 184 -199 0 1
rlabel polysilicon 184 -205 184 -205 0 3
rlabel polysilicon 191 -199 191 -199 0 1
rlabel polysilicon 191 -205 191 -205 0 3
rlabel polysilicon 198 -199 198 -199 0 1
rlabel polysilicon 198 -205 198 -205 0 3
rlabel polysilicon 205 -199 205 -199 0 1
rlabel polysilicon 205 -205 205 -205 0 3
rlabel polysilicon 212 -199 212 -199 0 1
rlabel polysilicon 212 -205 212 -205 0 3
rlabel polysilicon 219 -199 219 -199 0 1
rlabel polysilicon 219 -205 219 -205 0 3
rlabel polysilicon 226 -199 226 -199 0 1
rlabel polysilicon 226 -205 226 -205 0 3
rlabel polysilicon 233 -199 233 -199 0 1
rlabel polysilicon 233 -205 233 -205 0 3
rlabel polysilicon 240 -199 240 -199 0 1
rlabel polysilicon 240 -205 240 -205 0 3
rlabel polysilicon 243 -205 243 -205 0 4
rlabel polysilicon 247 -199 247 -199 0 1
rlabel polysilicon 247 -205 247 -205 0 3
rlabel polysilicon 254 -199 254 -199 0 1
rlabel polysilicon 254 -205 254 -205 0 3
rlabel polysilicon 261 -199 261 -199 0 1
rlabel polysilicon 261 -205 261 -205 0 3
rlabel polysilicon 268 -199 268 -199 0 1
rlabel polysilicon 271 -199 271 -199 0 2
rlabel polysilicon 268 -205 268 -205 0 3
rlabel polysilicon 271 -205 271 -205 0 4
rlabel polysilicon 275 -199 275 -199 0 1
rlabel polysilicon 275 -205 275 -205 0 3
rlabel polysilicon 282 -199 282 -199 0 1
rlabel polysilicon 282 -205 282 -205 0 3
rlabel polysilicon 289 -199 289 -199 0 1
rlabel polysilicon 289 -205 289 -205 0 3
rlabel polysilicon 296 -199 296 -199 0 1
rlabel polysilicon 296 -205 296 -205 0 3
rlabel polysilicon 303 -199 303 -199 0 1
rlabel polysilicon 306 -199 306 -199 0 2
rlabel polysilicon 303 -205 303 -205 0 3
rlabel polysilicon 310 -199 310 -199 0 1
rlabel polysilicon 310 -205 310 -205 0 3
rlabel polysilicon 317 -199 317 -199 0 1
rlabel polysilicon 320 -199 320 -199 0 2
rlabel polysilicon 317 -205 317 -205 0 3
rlabel polysilicon 320 -205 320 -205 0 4
rlabel polysilicon 324 -199 324 -199 0 1
rlabel polysilicon 324 -205 324 -205 0 3
rlabel polysilicon 331 -199 331 -199 0 1
rlabel polysilicon 334 -199 334 -199 0 2
rlabel polysilicon 334 -205 334 -205 0 4
rlabel polysilicon 338 -199 338 -199 0 1
rlabel polysilicon 338 -205 338 -205 0 3
rlabel polysilicon 345 -199 345 -199 0 1
rlabel polysilicon 345 -205 345 -205 0 3
rlabel polysilicon 352 -199 352 -199 0 1
rlabel polysilicon 352 -205 352 -205 0 3
rlabel polysilicon 359 -199 359 -199 0 1
rlabel polysilicon 359 -205 359 -205 0 3
rlabel polysilicon 366 -199 366 -199 0 1
rlabel polysilicon 366 -205 366 -205 0 3
rlabel polysilicon 373 -199 373 -199 0 1
rlabel polysilicon 373 -205 373 -205 0 3
rlabel polysilicon 380 -199 380 -199 0 1
rlabel polysilicon 380 -205 380 -205 0 3
rlabel polysilicon 387 -199 387 -199 0 1
rlabel polysilicon 390 -199 390 -199 0 2
rlabel polysilicon 387 -205 387 -205 0 3
rlabel polysilicon 390 -205 390 -205 0 4
rlabel polysilicon 394 -199 394 -199 0 1
rlabel polysilicon 394 -205 394 -205 0 3
rlabel polysilicon 401 -199 401 -199 0 1
rlabel polysilicon 401 -205 401 -205 0 3
rlabel polysilicon 408 -199 408 -199 0 1
rlabel polysilicon 408 -205 408 -205 0 3
rlabel polysilicon 415 -199 415 -199 0 1
rlabel polysilicon 415 -205 415 -205 0 3
rlabel polysilicon 422 -199 422 -199 0 1
rlabel polysilicon 422 -205 422 -205 0 3
rlabel polysilicon 429 -199 429 -199 0 1
rlabel polysilicon 429 -205 429 -205 0 3
rlabel polysilicon 436 -199 436 -199 0 1
rlabel polysilicon 439 -199 439 -199 0 2
rlabel polysilicon 436 -205 436 -205 0 3
rlabel polysilicon 439 -205 439 -205 0 4
rlabel polysilicon 443 -199 443 -199 0 1
rlabel polysilicon 443 -205 443 -205 0 3
rlabel polysilicon 446 -205 446 -205 0 4
rlabel polysilicon 450 -199 450 -199 0 1
rlabel polysilicon 450 -205 450 -205 0 3
rlabel polysilicon 457 -199 457 -199 0 1
rlabel polysilicon 460 -199 460 -199 0 2
rlabel polysilicon 457 -205 457 -205 0 3
rlabel polysilicon 464 -199 464 -199 0 1
rlabel polysilicon 464 -205 464 -205 0 3
rlabel polysilicon 471 -199 471 -199 0 1
rlabel polysilicon 471 -205 471 -205 0 3
rlabel polysilicon 478 -199 478 -199 0 1
rlabel polysilicon 478 -205 478 -205 0 3
rlabel polysilicon 485 -199 485 -199 0 1
rlabel polysilicon 488 -199 488 -199 0 2
rlabel polysilicon 485 -205 485 -205 0 3
rlabel polysilicon 492 -199 492 -199 0 1
rlabel polysilicon 492 -205 492 -205 0 3
rlabel polysilicon 499 -199 499 -199 0 1
rlabel polysilicon 499 -205 499 -205 0 3
rlabel polysilicon 506 -199 506 -199 0 1
rlabel polysilicon 506 -205 506 -205 0 3
rlabel polysilicon 516 -199 516 -199 0 2
rlabel polysilicon 513 -205 513 -205 0 3
rlabel polysilicon 516 -205 516 -205 0 4
rlabel polysilicon 520 -199 520 -199 0 1
rlabel polysilicon 520 -205 520 -205 0 3
rlabel polysilicon 527 -199 527 -199 0 1
rlabel polysilicon 527 -205 527 -205 0 3
rlabel polysilicon 534 -199 534 -199 0 1
rlabel polysilicon 537 -199 537 -199 0 2
rlabel polysilicon 534 -205 534 -205 0 3
rlabel polysilicon 537 -205 537 -205 0 4
rlabel polysilicon 541 -199 541 -199 0 1
rlabel polysilicon 541 -205 541 -205 0 3
rlabel polysilicon 548 -199 548 -199 0 1
rlabel polysilicon 548 -205 548 -205 0 3
rlabel polysilicon 555 -199 555 -199 0 1
rlabel polysilicon 555 -205 555 -205 0 3
rlabel polysilicon 562 -199 562 -199 0 1
rlabel polysilicon 562 -205 562 -205 0 3
rlabel polysilicon 569 -199 569 -199 0 1
rlabel polysilicon 569 -205 569 -205 0 3
rlabel polysilicon 576 -199 576 -199 0 1
rlabel polysilicon 576 -205 576 -205 0 3
rlabel polysilicon 583 -199 583 -199 0 1
rlabel polysilicon 583 -205 583 -205 0 3
rlabel polysilicon 590 -199 590 -199 0 1
rlabel polysilicon 590 -205 590 -205 0 3
rlabel polysilicon 597 -199 597 -199 0 1
rlabel polysilicon 597 -205 597 -205 0 3
rlabel polysilicon 604 -199 604 -199 0 1
rlabel polysilicon 607 -199 607 -199 0 2
rlabel polysilicon 604 -205 604 -205 0 3
rlabel polysilicon 607 -205 607 -205 0 4
rlabel polysilicon 611 -199 611 -199 0 1
rlabel polysilicon 611 -205 611 -205 0 3
rlabel polysilicon 618 -199 618 -199 0 1
rlabel polysilicon 618 -205 618 -205 0 3
rlabel polysilicon 625 -199 625 -199 0 1
rlabel polysilicon 625 -205 625 -205 0 3
rlabel polysilicon 632 -199 632 -199 0 1
rlabel polysilicon 632 -205 632 -205 0 3
rlabel polysilicon 639 -199 639 -199 0 1
rlabel polysilicon 639 -205 639 -205 0 3
rlabel polysilicon 646 -199 646 -199 0 1
rlabel polysilicon 646 -205 646 -205 0 3
rlabel polysilicon 653 -199 653 -199 0 1
rlabel polysilicon 653 -205 653 -205 0 3
rlabel polysilicon 660 -199 660 -199 0 1
rlabel polysilicon 660 -205 660 -205 0 3
rlabel polysilicon 667 -199 667 -199 0 1
rlabel polysilicon 667 -205 667 -205 0 3
rlabel polysilicon 674 -199 674 -199 0 1
rlabel polysilicon 674 -205 674 -205 0 3
rlabel polysilicon 681 -199 681 -199 0 1
rlabel polysilicon 681 -205 681 -205 0 3
rlabel polysilicon 688 -199 688 -199 0 1
rlabel polysilicon 688 -205 688 -205 0 3
rlabel polysilicon 695 -199 695 -199 0 1
rlabel polysilicon 695 -205 695 -205 0 3
rlabel polysilicon 702 -199 702 -199 0 1
rlabel polysilicon 702 -205 702 -205 0 3
rlabel polysilicon 709 -199 709 -199 0 1
rlabel polysilicon 709 -205 709 -205 0 3
rlabel polysilicon 719 -199 719 -199 0 2
rlabel polysilicon 716 -205 716 -205 0 3
rlabel polysilicon 719 -205 719 -205 0 4
rlabel polysilicon 723 -199 723 -199 0 1
rlabel polysilicon 723 -205 723 -205 0 3
rlabel polysilicon 730 -199 730 -199 0 1
rlabel polysilicon 730 -205 730 -205 0 3
rlabel polysilicon 737 -199 737 -199 0 1
rlabel polysilicon 737 -205 737 -205 0 3
rlabel polysilicon 744 -199 744 -199 0 1
rlabel polysilicon 744 -205 744 -205 0 3
rlabel polysilicon 751 -199 751 -199 0 1
rlabel polysilicon 751 -205 751 -205 0 3
rlabel polysilicon 758 -199 758 -199 0 1
rlabel polysilicon 758 -205 758 -205 0 3
rlabel polysilicon 765 -199 765 -199 0 1
rlabel polysilicon 765 -205 765 -205 0 3
rlabel polysilicon 772 -199 772 -199 0 1
rlabel polysilicon 772 -205 772 -205 0 3
rlabel polysilicon 779 -199 779 -199 0 1
rlabel polysilicon 779 -205 779 -205 0 3
rlabel polysilicon 786 -199 786 -199 0 1
rlabel polysilicon 786 -205 786 -205 0 3
rlabel polysilicon 793 -199 793 -199 0 1
rlabel polysilicon 793 -205 793 -205 0 3
rlabel polysilicon 800 -199 800 -199 0 1
rlabel polysilicon 800 -205 800 -205 0 3
rlabel polysilicon 807 -199 807 -199 0 1
rlabel polysilicon 807 -205 807 -205 0 3
rlabel polysilicon 814 -199 814 -199 0 1
rlabel polysilicon 814 -205 814 -205 0 3
rlabel polysilicon 821 -199 821 -199 0 1
rlabel polysilicon 821 -205 821 -205 0 3
rlabel polysilicon 828 -199 828 -199 0 1
rlabel polysilicon 828 -205 828 -205 0 3
rlabel polysilicon 835 -199 835 -199 0 1
rlabel polysilicon 835 -205 835 -205 0 3
rlabel polysilicon 842 -199 842 -199 0 1
rlabel polysilicon 842 -205 842 -205 0 3
rlabel polysilicon 849 -199 849 -199 0 1
rlabel polysilicon 849 -205 849 -205 0 3
rlabel polysilicon 856 -199 856 -199 0 1
rlabel polysilicon 856 -205 856 -205 0 3
rlabel polysilicon 863 -199 863 -199 0 1
rlabel polysilicon 863 -205 863 -205 0 3
rlabel polysilicon 870 -199 870 -199 0 1
rlabel polysilicon 870 -205 870 -205 0 3
rlabel polysilicon 877 -199 877 -199 0 1
rlabel polysilicon 877 -205 877 -205 0 3
rlabel polysilicon 884 -199 884 -199 0 1
rlabel polysilicon 884 -205 884 -205 0 3
rlabel polysilicon 891 -199 891 -199 0 1
rlabel polysilicon 891 -205 891 -205 0 3
rlabel polysilicon 898 -199 898 -199 0 1
rlabel polysilicon 898 -205 898 -205 0 3
rlabel polysilicon 905 -199 905 -199 0 1
rlabel polysilicon 905 -205 905 -205 0 3
rlabel polysilicon 912 -199 912 -199 0 1
rlabel polysilicon 912 -205 912 -205 0 3
rlabel polysilicon 919 -199 919 -199 0 1
rlabel polysilicon 919 -205 919 -205 0 3
rlabel polysilicon 926 -199 926 -199 0 1
rlabel polysilicon 926 -205 926 -205 0 3
rlabel polysilicon 933 -199 933 -199 0 1
rlabel polysilicon 933 -205 933 -205 0 3
rlabel polysilicon 940 -199 940 -199 0 1
rlabel polysilicon 940 -205 940 -205 0 3
rlabel polysilicon 947 -199 947 -199 0 1
rlabel polysilicon 947 -205 947 -205 0 3
rlabel polysilicon 954 -199 954 -199 0 1
rlabel polysilicon 954 -205 954 -205 0 3
rlabel polysilicon 961 -199 961 -199 0 1
rlabel polysilicon 961 -205 961 -205 0 3
rlabel polysilicon 968 -199 968 -199 0 1
rlabel polysilicon 968 -205 968 -205 0 3
rlabel polysilicon 975 -199 975 -199 0 1
rlabel polysilicon 978 -199 978 -199 0 2
rlabel polysilicon 975 -205 975 -205 0 3
rlabel polysilicon 978 -205 978 -205 0 4
rlabel polysilicon 982 -199 982 -199 0 1
rlabel polysilicon 985 -199 985 -199 0 2
rlabel polysilicon 982 -205 982 -205 0 3
rlabel polysilicon 989 -199 989 -199 0 1
rlabel polysilicon 992 -205 992 -205 0 4
rlabel polysilicon 996 -199 996 -199 0 1
rlabel polysilicon 996 -205 996 -205 0 3
rlabel polysilicon 1024 -199 1024 -199 0 1
rlabel polysilicon 1024 -205 1024 -205 0 3
rlabel polysilicon 1500 -199 1500 -199 0 1
rlabel polysilicon 1500 -205 1500 -205 0 3
rlabel polysilicon 2 -310 2 -310 0 1
rlabel polysilicon 2 -316 2 -316 0 3
rlabel polysilicon 9 -310 9 -310 0 1
rlabel polysilicon 9 -316 9 -316 0 3
rlabel polysilicon 16 -310 16 -310 0 1
rlabel polysilicon 16 -316 16 -316 0 3
rlabel polysilicon 26 -310 26 -310 0 2
rlabel polysilicon 23 -316 23 -316 0 3
rlabel polysilicon 26 -316 26 -316 0 4
rlabel polysilicon 30 -310 30 -310 0 1
rlabel polysilicon 33 -310 33 -310 0 2
rlabel polysilicon 33 -316 33 -316 0 4
rlabel polysilicon 37 -310 37 -310 0 1
rlabel polysilicon 40 -310 40 -310 0 2
rlabel polysilicon 37 -316 37 -316 0 3
rlabel polysilicon 44 -310 44 -310 0 1
rlabel polysilicon 44 -316 44 -316 0 3
rlabel polysilicon 51 -310 51 -310 0 1
rlabel polysilicon 54 -310 54 -310 0 2
rlabel polysilicon 51 -316 51 -316 0 3
rlabel polysilicon 58 -310 58 -310 0 1
rlabel polysilicon 58 -316 58 -316 0 3
rlabel polysilicon 65 -310 65 -310 0 1
rlabel polysilicon 68 -310 68 -310 0 2
rlabel polysilicon 68 -316 68 -316 0 4
rlabel polysilicon 72 -310 72 -310 0 1
rlabel polysilicon 72 -316 72 -316 0 3
rlabel polysilicon 82 -310 82 -310 0 2
rlabel polysilicon 79 -316 79 -316 0 3
rlabel polysilicon 82 -316 82 -316 0 4
rlabel polysilicon 86 -310 86 -310 0 1
rlabel polysilicon 86 -316 86 -316 0 3
rlabel polysilicon 93 -310 93 -310 0 1
rlabel polysilicon 96 -310 96 -310 0 2
rlabel polysilicon 93 -316 93 -316 0 3
rlabel polysilicon 96 -316 96 -316 0 4
rlabel polysilicon 100 -310 100 -310 0 1
rlabel polysilicon 100 -316 100 -316 0 3
rlabel polysilicon 107 -310 107 -310 0 1
rlabel polysilicon 107 -316 107 -316 0 3
rlabel polysilicon 114 -310 114 -310 0 1
rlabel polysilicon 114 -316 114 -316 0 3
rlabel polysilicon 121 -310 121 -310 0 1
rlabel polysilicon 124 -310 124 -310 0 2
rlabel polysilicon 121 -316 121 -316 0 3
rlabel polysilicon 124 -316 124 -316 0 4
rlabel polysilicon 128 -310 128 -310 0 1
rlabel polysilicon 128 -316 128 -316 0 3
rlabel polysilicon 135 -310 135 -310 0 1
rlabel polysilicon 135 -316 135 -316 0 3
rlabel polysilicon 142 -310 142 -310 0 1
rlabel polysilicon 142 -316 142 -316 0 3
rlabel polysilicon 149 -310 149 -310 0 1
rlabel polysilicon 149 -316 149 -316 0 3
rlabel polysilicon 156 -310 156 -310 0 1
rlabel polysilicon 156 -316 156 -316 0 3
rlabel polysilicon 163 -310 163 -310 0 1
rlabel polysilicon 163 -316 163 -316 0 3
rlabel polysilicon 170 -310 170 -310 0 1
rlabel polysilicon 170 -316 170 -316 0 3
rlabel polysilicon 177 -310 177 -310 0 1
rlabel polysilicon 177 -316 177 -316 0 3
rlabel polysilicon 184 -310 184 -310 0 1
rlabel polysilicon 184 -316 184 -316 0 3
rlabel polysilicon 191 -310 191 -310 0 1
rlabel polysilicon 191 -316 191 -316 0 3
rlabel polysilicon 198 -310 198 -310 0 1
rlabel polysilicon 198 -316 198 -316 0 3
rlabel polysilicon 205 -310 205 -310 0 1
rlabel polysilicon 205 -316 205 -316 0 3
rlabel polysilicon 212 -310 212 -310 0 1
rlabel polysilicon 212 -316 212 -316 0 3
rlabel polysilicon 219 -310 219 -310 0 1
rlabel polysilicon 219 -316 219 -316 0 3
rlabel polysilicon 226 -310 226 -310 0 1
rlabel polysilicon 226 -316 226 -316 0 3
rlabel polysilicon 233 -310 233 -310 0 1
rlabel polysilicon 233 -316 233 -316 0 3
rlabel polysilicon 240 -310 240 -310 0 1
rlabel polysilicon 240 -316 240 -316 0 3
rlabel polysilicon 247 -310 247 -310 0 1
rlabel polysilicon 247 -316 247 -316 0 3
rlabel polysilicon 254 -310 254 -310 0 1
rlabel polysilicon 254 -316 254 -316 0 3
rlabel polysilicon 261 -310 261 -310 0 1
rlabel polysilicon 261 -316 261 -316 0 3
rlabel polysilicon 268 -310 268 -310 0 1
rlabel polysilicon 268 -316 268 -316 0 3
rlabel polysilicon 275 -310 275 -310 0 1
rlabel polysilicon 275 -316 275 -316 0 3
rlabel polysilicon 282 -310 282 -310 0 1
rlabel polysilicon 285 -310 285 -310 0 2
rlabel polysilicon 282 -316 282 -316 0 3
rlabel polysilicon 285 -316 285 -316 0 4
rlabel polysilicon 289 -310 289 -310 0 1
rlabel polysilicon 289 -316 289 -316 0 3
rlabel polysilicon 296 -310 296 -310 0 1
rlabel polysilicon 296 -316 296 -316 0 3
rlabel polysilicon 303 -310 303 -310 0 1
rlabel polysilicon 303 -316 303 -316 0 3
rlabel polysilicon 310 -310 310 -310 0 1
rlabel polysilicon 313 -310 313 -310 0 2
rlabel polysilicon 313 -316 313 -316 0 4
rlabel polysilicon 317 -310 317 -310 0 1
rlabel polysilicon 320 -310 320 -310 0 2
rlabel polysilicon 317 -316 317 -316 0 3
rlabel polysilicon 320 -316 320 -316 0 4
rlabel polysilicon 324 -310 324 -310 0 1
rlabel polysilicon 327 -310 327 -310 0 2
rlabel polysilicon 324 -316 324 -316 0 3
rlabel polysilicon 327 -316 327 -316 0 4
rlabel polysilicon 331 -310 331 -310 0 1
rlabel polysilicon 331 -316 331 -316 0 3
rlabel polysilicon 338 -310 338 -310 0 1
rlabel polysilicon 338 -316 338 -316 0 3
rlabel polysilicon 345 -310 345 -310 0 1
rlabel polysilicon 345 -316 345 -316 0 3
rlabel polysilicon 352 -310 352 -310 0 1
rlabel polysilicon 352 -316 352 -316 0 3
rlabel polysilicon 359 -310 359 -310 0 1
rlabel polysilicon 362 -310 362 -310 0 2
rlabel polysilicon 359 -316 359 -316 0 3
rlabel polysilicon 366 -310 366 -310 0 1
rlabel polysilicon 366 -316 366 -316 0 3
rlabel polysilicon 373 -310 373 -310 0 1
rlabel polysilicon 373 -316 373 -316 0 3
rlabel polysilicon 380 -310 380 -310 0 1
rlabel polysilicon 380 -316 380 -316 0 3
rlabel polysilicon 387 -310 387 -310 0 1
rlabel polysilicon 387 -316 387 -316 0 3
rlabel polysilicon 394 -310 394 -310 0 1
rlabel polysilicon 394 -316 394 -316 0 3
rlabel polysilicon 401 -310 401 -310 0 1
rlabel polysilicon 401 -316 401 -316 0 3
rlabel polysilicon 408 -310 408 -310 0 1
rlabel polysilicon 408 -316 408 -316 0 3
rlabel polysilicon 411 -316 411 -316 0 4
rlabel polysilicon 415 -310 415 -310 0 1
rlabel polysilicon 415 -316 415 -316 0 3
rlabel polysilicon 422 -310 422 -310 0 1
rlabel polysilicon 425 -310 425 -310 0 2
rlabel polysilicon 422 -316 422 -316 0 3
rlabel polysilicon 429 -310 429 -310 0 1
rlabel polysilicon 429 -316 429 -316 0 3
rlabel polysilicon 436 -310 436 -310 0 1
rlabel polysilicon 436 -316 436 -316 0 3
rlabel polysilicon 443 -310 443 -310 0 1
rlabel polysilicon 443 -316 443 -316 0 3
rlabel polysilicon 450 -310 450 -310 0 1
rlabel polysilicon 453 -310 453 -310 0 2
rlabel polysilicon 450 -316 450 -316 0 3
rlabel polysilicon 453 -316 453 -316 0 4
rlabel polysilicon 457 -310 457 -310 0 1
rlabel polysilicon 457 -316 457 -316 0 3
rlabel polysilicon 464 -310 464 -310 0 1
rlabel polysilicon 464 -316 464 -316 0 3
rlabel polysilicon 471 -310 471 -310 0 1
rlabel polysilicon 471 -316 471 -316 0 3
rlabel polysilicon 478 -310 478 -310 0 1
rlabel polysilicon 478 -316 478 -316 0 3
rlabel polysilicon 485 -310 485 -310 0 1
rlabel polysilicon 485 -316 485 -316 0 3
rlabel polysilicon 492 -310 492 -310 0 1
rlabel polysilicon 492 -316 492 -316 0 3
rlabel polysilicon 499 -310 499 -310 0 1
rlabel polysilicon 499 -316 499 -316 0 3
rlabel polysilicon 506 -310 506 -310 0 1
rlabel polysilicon 506 -316 506 -316 0 3
rlabel polysilicon 513 -310 513 -310 0 1
rlabel polysilicon 513 -316 513 -316 0 3
rlabel polysilicon 520 -310 520 -310 0 1
rlabel polysilicon 520 -316 520 -316 0 3
rlabel polysilicon 527 -310 527 -310 0 1
rlabel polysilicon 527 -316 527 -316 0 3
rlabel polysilicon 534 -310 534 -310 0 1
rlabel polysilicon 534 -316 534 -316 0 3
rlabel polysilicon 541 -310 541 -310 0 1
rlabel polysilicon 544 -310 544 -310 0 2
rlabel polysilicon 544 -316 544 -316 0 4
rlabel polysilicon 548 -310 548 -310 0 1
rlabel polysilicon 548 -316 548 -316 0 3
rlabel polysilicon 555 -310 555 -310 0 1
rlabel polysilicon 555 -316 555 -316 0 3
rlabel polysilicon 562 -310 562 -310 0 1
rlabel polysilicon 562 -316 562 -316 0 3
rlabel polysilicon 569 -310 569 -310 0 1
rlabel polysilicon 569 -316 569 -316 0 3
rlabel polysilicon 576 -310 576 -310 0 1
rlabel polysilicon 579 -310 579 -310 0 2
rlabel polysilicon 576 -316 576 -316 0 3
rlabel polysilicon 579 -316 579 -316 0 4
rlabel polysilicon 583 -310 583 -310 0 1
rlabel polysilicon 583 -316 583 -316 0 3
rlabel polysilicon 586 -316 586 -316 0 4
rlabel polysilicon 590 -310 590 -310 0 1
rlabel polysilicon 590 -316 590 -316 0 3
rlabel polysilicon 597 -310 597 -310 0 1
rlabel polysilicon 597 -316 597 -316 0 3
rlabel polysilicon 604 -310 604 -310 0 1
rlabel polysilicon 607 -310 607 -310 0 2
rlabel polysilicon 611 -310 611 -310 0 1
rlabel polysilicon 611 -316 611 -316 0 3
rlabel polysilicon 618 -310 618 -310 0 1
rlabel polysilicon 618 -316 618 -316 0 3
rlabel polysilicon 625 -310 625 -310 0 1
rlabel polysilicon 625 -316 625 -316 0 3
rlabel polysilicon 632 -310 632 -310 0 1
rlabel polysilicon 632 -316 632 -316 0 3
rlabel polysilicon 639 -310 639 -310 0 1
rlabel polysilicon 639 -316 639 -316 0 3
rlabel polysilicon 646 -310 646 -310 0 1
rlabel polysilicon 646 -316 646 -316 0 3
rlabel polysilicon 653 -310 653 -310 0 1
rlabel polysilicon 653 -316 653 -316 0 3
rlabel polysilicon 660 -310 660 -310 0 1
rlabel polysilicon 660 -316 660 -316 0 3
rlabel polysilicon 667 -310 667 -310 0 1
rlabel polysilicon 667 -316 667 -316 0 3
rlabel polysilicon 674 -310 674 -310 0 1
rlabel polysilicon 674 -316 674 -316 0 3
rlabel polysilicon 681 -310 681 -310 0 1
rlabel polysilicon 681 -316 681 -316 0 3
rlabel polysilicon 688 -310 688 -310 0 1
rlabel polysilicon 688 -316 688 -316 0 3
rlabel polysilicon 695 -310 695 -310 0 1
rlabel polysilicon 698 -310 698 -310 0 2
rlabel polysilicon 695 -316 695 -316 0 3
rlabel polysilicon 698 -316 698 -316 0 4
rlabel polysilicon 705 -310 705 -310 0 2
rlabel polysilicon 702 -316 702 -316 0 3
rlabel polysilicon 709 -310 709 -310 0 1
rlabel polysilicon 709 -316 709 -316 0 3
rlabel polysilicon 716 -310 716 -310 0 1
rlabel polysilicon 716 -316 716 -316 0 3
rlabel polysilicon 723 -310 723 -310 0 1
rlabel polysilicon 723 -316 723 -316 0 3
rlabel polysilicon 730 -310 730 -310 0 1
rlabel polysilicon 730 -316 730 -316 0 3
rlabel polysilicon 737 -310 737 -310 0 1
rlabel polysilicon 737 -316 737 -316 0 3
rlabel polysilicon 744 -310 744 -310 0 1
rlabel polysilicon 744 -316 744 -316 0 3
rlabel polysilicon 751 -310 751 -310 0 1
rlabel polysilicon 751 -316 751 -316 0 3
rlabel polysilicon 758 -310 758 -310 0 1
rlabel polysilicon 758 -316 758 -316 0 3
rlabel polysilicon 765 -310 765 -310 0 1
rlabel polysilicon 765 -316 765 -316 0 3
rlabel polysilicon 772 -310 772 -310 0 1
rlabel polysilicon 772 -316 772 -316 0 3
rlabel polysilicon 779 -310 779 -310 0 1
rlabel polysilicon 779 -316 779 -316 0 3
rlabel polysilicon 786 -310 786 -310 0 1
rlabel polysilicon 786 -316 786 -316 0 3
rlabel polysilicon 793 -310 793 -310 0 1
rlabel polysilicon 793 -316 793 -316 0 3
rlabel polysilicon 800 -310 800 -310 0 1
rlabel polysilicon 800 -316 800 -316 0 3
rlabel polysilicon 807 -310 807 -310 0 1
rlabel polysilicon 807 -316 807 -316 0 3
rlabel polysilicon 814 -310 814 -310 0 1
rlabel polysilicon 814 -316 814 -316 0 3
rlabel polysilicon 821 -310 821 -310 0 1
rlabel polysilicon 821 -316 821 -316 0 3
rlabel polysilicon 828 -310 828 -310 0 1
rlabel polysilicon 828 -316 828 -316 0 3
rlabel polysilicon 835 -310 835 -310 0 1
rlabel polysilicon 835 -316 835 -316 0 3
rlabel polysilicon 842 -310 842 -310 0 1
rlabel polysilicon 842 -316 842 -316 0 3
rlabel polysilicon 849 -310 849 -310 0 1
rlabel polysilicon 849 -316 849 -316 0 3
rlabel polysilicon 856 -310 856 -310 0 1
rlabel polysilicon 856 -316 856 -316 0 3
rlabel polysilicon 863 -310 863 -310 0 1
rlabel polysilicon 863 -316 863 -316 0 3
rlabel polysilicon 870 -310 870 -310 0 1
rlabel polysilicon 870 -316 870 -316 0 3
rlabel polysilicon 877 -310 877 -310 0 1
rlabel polysilicon 877 -316 877 -316 0 3
rlabel polysilicon 884 -310 884 -310 0 1
rlabel polysilicon 884 -316 884 -316 0 3
rlabel polysilicon 891 -310 891 -310 0 1
rlabel polysilicon 891 -316 891 -316 0 3
rlabel polysilicon 898 -310 898 -310 0 1
rlabel polysilicon 898 -316 898 -316 0 3
rlabel polysilicon 905 -310 905 -310 0 1
rlabel polysilicon 905 -316 905 -316 0 3
rlabel polysilicon 912 -310 912 -310 0 1
rlabel polysilicon 912 -316 912 -316 0 3
rlabel polysilicon 919 -310 919 -310 0 1
rlabel polysilicon 919 -316 919 -316 0 3
rlabel polysilicon 926 -310 926 -310 0 1
rlabel polysilicon 926 -316 926 -316 0 3
rlabel polysilicon 933 -310 933 -310 0 1
rlabel polysilicon 933 -316 933 -316 0 3
rlabel polysilicon 940 -310 940 -310 0 1
rlabel polysilicon 940 -316 940 -316 0 3
rlabel polysilicon 947 -310 947 -310 0 1
rlabel polysilicon 947 -316 947 -316 0 3
rlabel polysilicon 954 -310 954 -310 0 1
rlabel polysilicon 954 -316 954 -316 0 3
rlabel polysilicon 961 -310 961 -310 0 1
rlabel polysilicon 961 -316 961 -316 0 3
rlabel polysilicon 968 -310 968 -310 0 1
rlabel polysilicon 968 -316 968 -316 0 3
rlabel polysilicon 975 -310 975 -310 0 1
rlabel polysilicon 975 -316 975 -316 0 3
rlabel polysilicon 982 -310 982 -310 0 1
rlabel polysilicon 982 -316 982 -316 0 3
rlabel polysilicon 989 -310 989 -310 0 1
rlabel polysilicon 989 -316 989 -316 0 3
rlabel polysilicon 996 -310 996 -310 0 1
rlabel polysilicon 996 -316 996 -316 0 3
rlabel polysilicon 1003 -310 1003 -310 0 1
rlabel polysilicon 1003 -316 1003 -316 0 3
rlabel polysilicon 1010 -310 1010 -310 0 1
rlabel polysilicon 1010 -316 1010 -316 0 3
rlabel polysilicon 1017 -310 1017 -310 0 1
rlabel polysilicon 1017 -316 1017 -316 0 3
rlabel polysilicon 1024 -310 1024 -310 0 1
rlabel polysilicon 1024 -316 1024 -316 0 3
rlabel polysilicon 1031 -310 1031 -310 0 1
rlabel polysilicon 1031 -316 1031 -316 0 3
rlabel polysilicon 1038 -310 1038 -310 0 1
rlabel polysilicon 1038 -316 1038 -316 0 3
rlabel polysilicon 1045 -310 1045 -310 0 1
rlabel polysilicon 1045 -316 1045 -316 0 3
rlabel polysilicon 1052 -310 1052 -310 0 1
rlabel polysilicon 1052 -316 1052 -316 0 3
rlabel polysilicon 1059 -310 1059 -310 0 1
rlabel polysilicon 1059 -316 1059 -316 0 3
rlabel polysilicon 1066 -310 1066 -310 0 1
rlabel polysilicon 1066 -316 1066 -316 0 3
rlabel polysilicon 1073 -310 1073 -310 0 1
rlabel polysilicon 1073 -316 1073 -316 0 3
rlabel polysilicon 1080 -310 1080 -310 0 1
rlabel polysilicon 1080 -316 1080 -316 0 3
rlabel polysilicon 1087 -310 1087 -310 0 1
rlabel polysilicon 1087 -316 1087 -316 0 3
rlabel polysilicon 1094 -310 1094 -310 0 1
rlabel polysilicon 1094 -316 1094 -316 0 3
rlabel polysilicon 1101 -310 1101 -310 0 1
rlabel polysilicon 1101 -316 1101 -316 0 3
rlabel polysilicon 1108 -310 1108 -310 0 1
rlabel polysilicon 1108 -316 1108 -316 0 3
rlabel polysilicon 1115 -310 1115 -310 0 1
rlabel polysilicon 1115 -316 1115 -316 0 3
rlabel polysilicon 1122 -310 1122 -310 0 1
rlabel polysilicon 1122 -316 1122 -316 0 3
rlabel polysilicon 1129 -310 1129 -310 0 1
rlabel polysilicon 1129 -316 1129 -316 0 3
rlabel polysilicon 1136 -310 1136 -310 0 1
rlabel polysilicon 1136 -316 1136 -316 0 3
rlabel polysilicon 1143 -310 1143 -310 0 1
rlabel polysilicon 1143 -316 1143 -316 0 3
rlabel polysilicon 1150 -310 1150 -310 0 1
rlabel polysilicon 1153 -310 1153 -310 0 2
rlabel polysilicon 1178 -310 1178 -310 0 1
rlabel polysilicon 1178 -316 1178 -316 0 3
rlabel polysilicon 1500 -310 1500 -310 0 1
rlabel polysilicon 1500 -316 1500 -316 0 3
rlabel polysilicon 2 -399 2 -399 0 1
rlabel polysilicon 2 -405 2 -405 0 3
rlabel polysilicon 9 -399 9 -399 0 1
rlabel polysilicon 9 -405 9 -405 0 3
rlabel polysilicon 16 -399 16 -399 0 1
rlabel polysilicon 16 -405 16 -405 0 3
rlabel polysilicon 23 -399 23 -399 0 1
rlabel polysilicon 26 -399 26 -399 0 2
rlabel polysilicon 23 -405 23 -405 0 3
rlabel polysilicon 26 -405 26 -405 0 4
rlabel polysilicon 30 -399 30 -399 0 1
rlabel polysilicon 30 -405 30 -405 0 3
rlabel polysilicon 37 -399 37 -399 0 1
rlabel polysilicon 40 -399 40 -399 0 2
rlabel polysilicon 37 -405 37 -405 0 3
rlabel polysilicon 44 -399 44 -399 0 1
rlabel polysilicon 47 -399 47 -399 0 2
rlabel polysilicon 44 -405 44 -405 0 3
rlabel polysilicon 47 -405 47 -405 0 4
rlabel polysilicon 51 -399 51 -399 0 1
rlabel polysilicon 51 -405 51 -405 0 3
rlabel polysilicon 58 -399 58 -399 0 1
rlabel polysilicon 61 -399 61 -399 0 2
rlabel polysilicon 58 -405 58 -405 0 3
rlabel polysilicon 61 -405 61 -405 0 4
rlabel polysilicon 65 -399 65 -399 0 1
rlabel polysilicon 65 -405 65 -405 0 3
rlabel polysilicon 72 -399 72 -399 0 1
rlabel polysilicon 75 -399 75 -399 0 2
rlabel polysilicon 75 -405 75 -405 0 4
rlabel polysilicon 79 -399 79 -399 0 1
rlabel polysilicon 82 -399 82 -399 0 2
rlabel polysilicon 79 -405 79 -405 0 3
rlabel polysilicon 82 -405 82 -405 0 4
rlabel polysilicon 86 -399 86 -399 0 1
rlabel polysilicon 89 -399 89 -399 0 2
rlabel polysilicon 86 -405 86 -405 0 3
rlabel polysilicon 89 -405 89 -405 0 4
rlabel polysilicon 93 -399 93 -399 0 1
rlabel polysilicon 93 -405 93 -405 0 3
rlabel polysilicon 100 -399 100 -399 0 1
rlabel polysilicon 100 -405 100 -405 0 3
rlabel polysilicon 107 -399 107 -399 0 1
rlabel polysilicon 107 -405 107 -405 0 3
rlabel polysilicon 114 -399 114 -399 0 1
rlabel polysilicon 114 -405 114 -405 0 3
rlabel polysilicon 121 -399 121 -399 0 1
rlabel polysilicon 124 -399 124 -399 0 2
rlabel polysilicon 124 -405 124 -405 0 4
rlabel polysilicon 128 -399 128 -399 0 1
rlabel polysilicon 128 -405 128 -405 0 3
rlabel polysilicon 135 -399 135 -399 0 1
rlabel polysilicon 135 -405 135 -405 0 3
rlabel polysilicon 142 -399 142 -399 0 1
rlabel polysilicon 142 -405 142 -405 0 3
rlabel polysilicon 149 -399 149 -399 0 1
rlabel polysilicon 149 -405 149 -405 0 3
rlabel polysilicon 156 -399 156 -399 0 1
rlabel polysilicon 156 -405 156 -405 0 3
rlabel polysilicon 163 -399 163 -399 0 1
rlabel polysilicon 163 -405 163 -405 0 3
rlabel polysilicon 170 -399 170 -399 0 1
rlabel polysilicon 170 -405 170 -405 0 3
rlabel polysilicon 177 -399 177 -399 0 1
rlabel polysilicon 177 -405 177 -405 0 3
rlabel polysilicon 184 -399 184 -399 0 1
rlabel polysilicon 184 -405 184 -405 0 3
rlabel polysilicon 191 -399 191 -399 0 1
rlabel polysilicon 191 -405 191 -405 0 3
rlabel polysilicon 198 -399 198 -399 0 1
rlabel polysilicon 198 -405 198 -405 0 3
rlabel polysilicon 205 -399 205 -399 0 1
rlabel polysilicon 205 -405 205 -405 0 3
rlabel polysilicon 212 -399 212 -399 0 1
rlabel polysilicon 212 -405 212 -405 0 3
rlabel polysilicon 219 -399 219 -399 0 1
rlabel polysilicon 219 -405 219 -405 0 3
rlabel polysilicon 226 -399 226 -399 0 1
rlabel polysilicon 226 -405 226 -405 0 3
rlabel polysilicon 233 -399 233 -399 0 1
rlabel polysilicon 233 -405 233 -405 0 3
rlabel polysilicon 240 -399 240 -399 0 1
rlabel polysilicon 240 -405 240 -405 0 3
rlabel polysilicon 247 -399 247 -399 0 1
rlabel polysilicon 247 -405 247 -405 0 3
rlabel polysilicon 254 -399 254 -399 0 1
rlabel polysilicon 254 -405 254 -405 0 3
rlabel polysilicon 261 -399 261 -399 0 1
rlabel polysilicon 264 -399 264 -399 0 2
rlabel polysilicon 261 -405 261 -405 0 3
rlabel polysilicon 264 -405 264 -405 0 4
rlabel polysilicon 268 -399 268 -399 0 1
rlabel polysilicon 268 -405 268 -405 0 3
rlabel polysilicon 275 -399 275 -399 0 1
rlabel polysilicon 275 -405 275 -405 0 3
rlabel polysilicon 282 -399 282 -399 0 1
rlabel polysilicon 282 -405 282 -405 0 3
rlabel polysilicon 289 -399 289 -399 0 1
rlabel polysilicon 289 -405 289 -405 0 3
rlabel polysilicon 296 -399 296 -399 0 1
rlabel polysilicon 296 -405 296 -405 0 3
rlabel polysilicon 303 -399 303 -399 0 1
rlabel polysilicon 303 -405 303 -405 0 3
rlabel polysilicon 310 -399 310 -399 0 1
rlabel polysilicon 310 -405 310 -405 0 3
rlabel polysilicon 317 -399 317 -399 0 1
rlabel polysilicon 317 -405 317 -405 0 3
rlabel polysilicon 324 -399 324 -399 0 1
rlabel polysilicon 324 -405 324 -405 0 3
rlabel polysilicon 331 -399 331 -399 0 1
rlabel polysilicon 331 -405 331 -405 0 3
rlabel polysilicon 338 -399 338 -399 0 1
rlabel polysilicon 338 -405 338 -405 0 3
rlabel polysilicon 345 -399 345 -399 0 1
rlabel polysilicon 345 -405 345 -405 0 3
rlabel polysilicon 352 -399 352 -399 0 1
rlabel polysilicon 352 -405 352 -405 0 3
rlabel polysilicon 359 -399 359 -399 0 1
rlabel polysilicon 359 -405 359 -405 0 3
rlabel polysilicon 366 -399 366 -399 0 1
rlabel polysilicon 366 -405 366 -405 0 3
rlabel polysilicon 373 -399 373 -399 0 1
rlabel polysilicon 373 -405 373 -405 0 3
rlabel polysilicon 380 -399 380 -399 0 1
rlabel polysilicon 380 -405 380 -405 0 3
rlabel polysilicon 387 -399 387 -399 0 1
rlabel polysilicon 387 -405 387 -405 0 3
rlabel polysilicon 397 -399 397 -399 0 2
rlabel polysilicon 394 -405 394 -405 0 3
rlabel polysilicon 397 -405 397 -405 0 4
rlabel polysilicon 401 -399 401 -399 0 1
rlabel polysilicon 401 -405 401 -405 0 3
rlabel polysilicon 408 -399 408 -399 0 1
rlabel polysilicon 411 -399 411 -399 0 2
rlabel polysilicon 408 -405 408 -405 0 3
rlabel polysilicon 411 -405 411 -405 0 4
rlabel polysilicon 415 -399 415 -399 0 1
rlabel polysilicon 415 -405 415 -405 0 3
rlabel polysilicon 422 -399 422 -399 0 1
rlabel polysilicon 422 -405 422 -405 0 3
rlabel polysilicon 429 -399 429 -399 0 1
rlabel polysilicon 429 -405 429 -405 0 3
rlabel polysilicon 436 -399 436 -399 0 1
rlabel polysilicon 436 -405 436 -405 0 3
rlabel polysilicon 443 -399 443 -399 0 1
rlabel polysilicon 443 -405 443 -405 0 3
rlabel polysilicon 450 -399 450 -399 0 1
rlabel polysilicon 450 -405 450 -405 0 3
rlabel polysilicon 457 -399 457 -399 0 1
rlabel polysilicon 457 -405 457 -405 0 3
rlabel polysilicon 464 -399 464 -399 0 1
rlabel polysilicon 464 -405 464 -405 0 3
rlabel polysilicon 471 -399 471 -399 0 1
rlabel polysilicon 471 -405 471 -405 0 3
rlabel polysilicon 478 -399 478 -399 0 1
rlabel polysilicon 478 -405 478 -405 0 3
rlabel polysilicon 485 -399 485 -399 0 1
rlabel polysilicon 485 -405 485 -405 0 3
rlabel polysilicon 492 -399 492 -399 0 1
rlabel polysilicon 492 -405 492 -405 0 3
rlabel polysilicon 499 -399 499 -399 0 1
rlabel polysilicon 502 -399 502 -399 0 2
rlabel polysilicon 499 -405 499 -405 0 3
rlabel polysilicon 502 -405 502 -405 0 4
rlabel polysilicon 506 -399 506 -399 0 1
rlabel polysilicon 509 -399 509 -399 0 2
rlabel polysilicon 513 -399 513 -399 0 1
rlabel polysilicon 516 -399 516 -399 0 2
rlabel polysilicon 516 -405 516 -405 0 4
rlabel polysilicon 520 -399 520 -399 0 1
rlabel polysilicon 520 -405 520 -405 0 3
rlabel polysilicon 527 -399 527 -399 0 1
rlabel polysilicon 527 -405 527 -405 0 3
rlabel polysilicon 534 -399 534 -399 0 1
rlabel polysilicon 534 -405 534 -405 0 3
rlabel polysilicon 541 -399 541 -399 0 1
rlabel polysilicon 541 -405 541 -405 0 3
rlabel polysilicon 548 -399 548 -399 0 1
rlabel polysilicon 551 -399 551 -399 0 2
rlabel polysilicon 548 -405 548 -405 0 3
rlabel polysilicon 551 -405 551 -405 0 4
rlabel polysilicon 555 -399 555 -399 0 1
rlabel polysilicon 555 -405 555 -405 0 3
rlabel polysilicon 565 -399 565 -399 0 2
rlabel polysilicon 562 -405 562 -405 0 3
rlabel polysilicon 565 -405 565 -405 0 4
rlabel polysilicon 569 -399 569 -399 0 1
rlabel polysilicon 572 -399 572 -399 0 2
rlabel polysilicon 569 -405 569 -405 0 3
rlabel polysilicon 572 -405 572 -405 0 4
rlabel polysilicon 576 -399 576 -399 0 1
rlabel polysilicon 576 -405 576 -405 0 3
rlabel polysilicon 583 -399 583 -399 0 1
rlabel polysilicon 583 -405 583 -405 0 3
rlabel polysilicon 590 -399 590 -399 0 1
rlabel polysilicon 590 -405 590 -405 0 3
rlabel polysilicon 593 -405 593 -405 0 4
rlabel polysilicon 597 -399 597 -399 0 1
rlabel polysilicon 597 -405 597 -405 0 3
rlabel polysilicon 604 -399 604 -399 0 1
rlabel polysilicon 604 -405 604 -405 0 3
rlabel polysilicon 611 -399 611 -399 0 1
rlabel polysilicon 611 -405 611 -405 0 3
rlabel polysilicon 618 -399 618 -399 0 1
rlabel polysilicon 618 -405 618 -405 0 3
rlabel polysilicon 625 -399 625 -399 0 1
rlabel polysilicon 625 -405 625 -405 0 3
rlabel polysilicon 632 -399 632 -399 0 1
rlabel polysilicon 632 -405 632 -405 0 3
rlabel polysilicon 639 -399 639 -399 0 1
rlabel polysilicon 642 -399 642 -399 0 2
rlabel polysilicon 642 -405 642 -405 0 4
rlabel polysilicon 646 -399 646 -399 0 1
rlabel polysilicon 646 -405 646 -405 0 3
rlabel polysilicon 653 -399 653 -399 0 1
rlabel polysilicon 653 -405 653 -405 0 3
rlabel polysilicon 660 -399 660 -399 0 1
rlabel polysilicon 660 -405 660 -405 0 3
rlabel polysilicon 663 -405 663 -405 0 4
rlabel polysilicon 667 -399 667 -399 0 1
rlabel polysilicon 670 -399 670 -399 0 2
rlabel polysilicon 667 -405 667 -405 0 3
rlabel polysilicon 670 -405 670 -405 0 4
rlabel polysilicon 674 -399 674 -399 0 1
rlabel polysilicon 674 -405 674 -405 0 3
rlabel polysilicon 681 -399 681 -399 0 1
rlabel polysilicon 681 -405 681 -405 0 3
rlabel polysilicon 688 -399 688 -399 0 1
rlabel polysilicon 688 -405 688 -405 0 3
rlabel polysilicon 695 -399 695 -399 0 1
rlabel polysilicon 695 -405 695 -405 0 3
rlabel polysilicon 702 -399 702 -399 0 1
rlabel polysilicon 702 -405 702 -405 0 3
rlabel polysilicon 709 -399 709 -399 0 1
rlabel polysilicon 709 -405 709 -405 0 3
rlabel polysilicon 716 -399 716 -399 0 1
rlabel polysilicon 716 -405 716 -405 0 3
rlabel polysilicon 723 -399 723 -399 0 1
rlabel polysilicon 723 -405 723 -405 0 3
rlabel polysilicon 730 -399 730 -399 0 1
rlabel polysilicon 730 -405 730 -405 0 3
rlabel polysilicon 737 -399 737 -399 0 1
rlabel polysilicon 737 -405 737 -405 0 3
rlabel polysilicon 744 -399 744 -399 0 1
rlabel polysilicon 744 -405 744 -405 0 3
rlabel polysilicon 751 -399 751 -399 0 1
rlabel polysilicon 751 -405 751 -405 0 3
rlabel polysilicon 758 -399 758 -399 0 1
rlabel polysilicon 758 -405 758 -405 0 3
rlabel polysilicon 765 -399 765 -399 0 1
rlabel polysilicon 765 -405 765 -405 0 3
rlabel polysilicon 772 -399 772 -399 0 1
rlabel polysilicon 772 -405 772 -405 0 3
rlabel polysilicon 779 -399 779 -399 0 1
rlabel polysilicon 779 -405 779 -405 0 3
rlabel polysilicon 786 -399 786 -399 0 1
rlabel polysilicon 786 -405 786 -405 0 3
rlabel polysilicon 793 -399 793 -399 0 1
rlabel polysilicon 793 -405 793 -405 0 3
rlabel polysilicon 800 -399 800 -399 0 1
rlabel polysilicon 800 -405 800 -405 0 3
rlabel polysilicon 807 -399 807 -399 0 1
rlabel polysilicon 807 -405 807 -405 0 3
rlabel polysilicon 814 -399 814 -399 0 1
rlabel polysilicon 814 -405 814 -405 0 3
rlabel polysilicon 821 -399 821 -399 0 1
rlabel polysilicon 821 -405 821 -405 0 3
rlabel polysilicon 828 -399 828 -399 0 1
rlabel polysilicon 828 -405 828 -405 0 3
rlabel polysilicon 835 -399 835 -399 0 1
rlabel polysilicon 835 -405 835 -405 0 3
rlabel polysilicon 842 -399 842 -399 0 1
rlabel polysilicon 842 -405 842 -405 0 3
rlabel polysilicon 849 -399 849 -399 0 1
rlabel polysilicon 849 -405 849 -405 0 3
rlabel polysilicon 856 -399 856 -399 0 1
rlabel polysilicon 856 -405 856 -405 0 3
rlabel polysilicon 863 -399 863 -399 0 1
rlabel polysilicon 863 -405 863 -405 0 3
rlabel polysilicon 870 -399 870 -399 0 1
rlabel polysilicon 870 -405 870 -405 0 3
rlabel polysilicon 877 -399 877 -399 0 1
rlabel polysilicon 877 -405 877 -405 0 3
rlabel polysilicon 884 -399 884 -399 0 1
rlabel polysilicon 884 -405 884 -405 0 3
rlabel polysilicon 891 -399 891 -399 0 1
rlabel polysilicon 891 -405 891 -405 0 3
rlabel polysilicon 898 -399 898 -399 0 1
rlabel polysilicon 898 -405 898 -405 0 3
rlabel polysilicon 905 -399 905 -399 0 1
rlabel polysilicon 905 -405 905 -405 0 3
rlabel polysilicon 912 -399 912 -399 0 1
rlabel polysilicon 912 -405 912 -405 0 3
rlabel polysilicon 919 -399 919 -399 0 1
rlabel polysilicon 919 -405 919 -405 0 3
rlabel polysilicon 926 -399 926 -399 0 1
rlabel polysilicon 926 -405 926 -405 0 3
rlabel polysilicon 933 -399 933 -399 0 1
rlabel polysilicon 933 -405 933 -405 0 3
rlabel polysilicon 940 -399 940 -399 0 1
rlabel polysilicon 940 -405 940 -405 0 3
rlabel polysilicon 947 -399 947 -399 0 1
rlabel polysilicon 947 -405 947 -405 0 3
rlabel polysilicon 954 -399 954 -399 0 1
rlabel polysilicon 954 -405 954 -405 0 3
rlabel polysilicon 961 -399 961 -399 0 1
rlabel polysilicon 961 -405 961 -405 0 3
rlabel polysilicon 968 -399 968 -399 0 1
rlabel polysilicon 968 -405 968 -405 0 3
rlabel polysilicon 975 -399 975 -399 0 1
rlabel polysilicon 975 -405 975 -405 0 3
rlabel polysilicon 982 -399 982 -399 0 1
rlabel polysilicon 982 -405 982 -405 0 3
rlabel polysilicon 989 -399 989 -399 0 1
rlabel polysilicon 989 -405 989 -405 0 3
rlabel polysilicon 996 -399 996 -399 0 1
rlabel polysilicon 996 -405 996 -405 0 3
rlabel polysilicon 1003 -399 1003 -399 0 1
rlabel polysilicon 1003 -405 1003 -405 0 3
rlabel polysilicon 1010 -399 1010 -399 0 1
rlabel polysilicon 1010 -405 1010 -405 0 3
rlabel polysilicon 1017 -399 1017 -399 0 1
rlabel polysilicon 1017 -405 1017 -405 0 3
rlabel polysilicon 1024 -399 1024 -399 0 1
rlabel polysilicon 1024 -405 1024 -405 0 3
rlabel polysilicon 1031 -399 1031 -399 0 1
rlabel polysilicon 1031 -405 1031 -405 0 3
rlabel polysilicon 1038 -399 1038 -399 0 1
rlabel polysilicon 1038 -405 1038 -405 0 3
rlabel polysilicon 1045 -399 1045 -399 0 1
rlabel polysilicon 1045 -405 1045 -405 0 3
rlabel polysilicon 1052 -399 1052 -399 0 1
rlabel polysilicon 1052 -405 1052 -405 0 3
rlabel polysilicon 1059 -399 1059 -399 0 1
rlabel polysilicon 1059 -405 1059 -405 0 3
rlabel polysilicon 1066 -399 1066 -399 0 1
rlabel polysilicon 1066 -405 1066 -405 0 3
rlabel polysilicon 1073 -399 1073 -399 0 1
rlabel polysilicon 1073 -405 1073 -405 0 3
rlabel polysilicon 1080 -399 1080 -399 0 1
rlabel polysilicon 1080 -405 1080 -405 0 3
rlabel polysilicon 1087 -399 1087 -399 0 1
rlabel polysilicon 1087 -405 1087 -405 0 3
rlabel polysilicon 1094 -399 1094 -399 0 1
rlabel polysilicon 1094 -405 1094 -405 0 3
rlabel polysilicon 1101 -399 1101 -399 0 1
rlabel polysilicon 1101 -405 1101 -405 0 3
rlabel polysilicon 1108 -399 1108 -399 0 1
rlabel polysilicon 1108 -405 1108 -405 0 3
rlabel polysilicon 1115 -399 1115 -399 0 1
rlabel polysilicon 1115 -405 1115 -405 0 3
rlabel polysilicon 1122 -399 1122 -399 0 1
rlabel polysilicon 1122 -405 1122 -405 0 3
rlabel polysilicon 1129 -399 1129 -399 0 1
rlabel polysilicon 1129 -405 1129 -405 0 3
rlabel polysilicon 1136 -399 1136 -399 0 1
rlabel polysilicon 1136 -405 1136 -405 0 3
rlabel polysilicon 1143 -399 1143 -399 0 1
rlabel polysilicon 1143 -405 1143 -405 0 3
rlabel polysilicon 1150 -399 1150 -399 0 1
rlabel polysilicon 1150 -405 1150 -405 0 3
rlabel polysilicon 1157 -399 1157 -399 0 1
rlabel polysilicon 1157 -405 1157 -405 0 3
rlabel polysilicon 1164 -399 1164 -399 0 1
rlabel polysilicon 1164 -405 1164 -405 0 3
rlabel polysilicon 1171 -399 1171 -399 0 1
rlabel polysilicon 1171 -405 1171 -405 0 3
rlabel polysilicon 1178 -399 1178 -399 0 1
rlabel polysilicon 1178 -405 1178 -405 0 3
rlabel polysilicon 1185 -399 1185 -399 0 1
rlabel polysilicon 1185 -405 1185 -405 0 3
rlabel polysilicon 1192 -399 1192 -399 0 1
rlabel polysilicon 1192 -405 1192 -405 0 3
rlabel polysilicon 1202 -399 1202 -399 0 2
rlabel polysilicon 1199 -405 1199 -405 0 3
rlabel polysilicon 1202 -405 1202 -405 0 4
rlabel polysilicon 1209 -399 1209 -399 0 2
rlabel polysilicon 1209 -405 1209 -405 0 4
rlabel polysilicon 1500 -399 1500 -399 0 1
rlabel polysilicon 1500 -405 1500 -405 0 3
rlabel polysilicon 2 -520 2 -520 0 3
rlabel polysilicon 5 -520 5 -520 0 4
rlabel polysilicon 9 -514 9 -514 0 1
rlabel polysilicon 9 -520 9 -520 0 3
rlabel polysilicon 16 -514 16 -514 0 1
rlabel polysilicon 16 -520 16 -520 0 3
rlabel polysilicon 23 -514 23 -514 0 1
rlabel polysilicon 23 -520 23 -520 0 3
rlabel polysilicon 30 -514 30 -514 0 1
rlabel polysilicon 33 -514 33 -514 0 2
rlabel polysilicon 33 -520 33 -520 0 4
rlabel polysilicon 37 -514 37 -514 0 1
rlabel polysilicon 40 -514 40 -514 0 2
rlabel polysilicon 37 -520 37 -520 0 3
rlabel polysilicon 40 -520 40 -520 0 4
rlabel polysilicon 44 -514 44 -514 0 1
rlabel polysilicon 44 -520 44 -520 0 3
rlabel polysilicon 51 -514 51 -514 0 1
rlabel polysilicon 51 -520 51 -520 0 3
rlabel polysilicon 58 -514 58 -514 0 1
rlabel polysilicon 58 -520 58 -520 0 3
rlabel polysilicon 65 -514 65 -514 0 1
rlabel polysilicon 65 -520 65 -520 0 3
rlabel polysilicon 72 -514 72 -514 0 1
rlabel polysilicon 75 -514 75 -514 0 2
rlabel polysilicon 72 -520 72 -520 0 3
rlabel polysilicon 79 -514 79 -514 0 1
rlabel polysilicon 79 -520 79 -520 0 3
rlabel polysilicon 86 -514 86 -514 0 1
rlabel polysilicon 89 -514 89 -514 0 2
rlabel polysilicon 86 -520 86 -520 0 3
rlabel polysilicon 89 -520 89 -520 0 4
rlabel polysilicon 93 -514 93 -514 0 1
rlabel polysilicon 93 -520 93 -520 0 3
rlabel polysilicon 100 -514 100 -514 0 1
rlabel polysilicon 100 -520 100 -520 0 3
rlabel polysilicon 107 -514 107 -514 0 1
rlabel polysilicon 110 -514 110 -514 0 2
rlabel polysilicon 107 -520 107 -520 0 3
rlabel polysilicon 110 -520 110 -520 0 4
rlabel polysilicon 114 -514 114 -514 0 1
rlabel polysilicon 114 -520 114 -520 0 3
rlabel polysilicon 121 -514 121 -514 0 1
rlabel polysilicon 121 -520 121 -520 0 3
rlabel polysilicon 128 -514 128 -514 0 1
rlabel polysilicon 128 -520 128 -520 0 3
rlabel polysilicon 135 -514 135 -514 0 1
rlabel polysilicon 138 -514 138 -514 0 2
rlabel polysilicon 135 -520 135 -520 0 3
rlabel polysilicon 138 -520 138 -520 0 4
rlabel polysilicon 142 -514 142 -514 0 1
rlabel polysilicon 145 -514 145 -514 0 2
rlabel polysilicon 142 -520 142 -520 0 3
rlabel polysilicon 145 -520 145 -520 0 4
rlabel polysilicon 149 -514 149 -514 0 1
rlabel polysilicon 149 -520 149 -520 0 3
rlabel polysilicon 159 -514 159 -514 0 2
rlabel polysilicon 156 -520 156 -520 0 3
rlabel polysilicon 159 -520 159 -520 0 4
rlabel polysilicon 163 -514 163 -514 0 1
rlabel polysilicon 163 -520 163 -520 0 3
rlabel polysilicon 170 -514 170 -514 0 1
rlabel polysilicon 170 -520 170 -520 0 3
rlabel polysilicon 177 -514 177 -514 0 1
rlabel polysilicon 177 -520 177 -520 0 3
rlabel polysilicon 184 -514 184 -514 0 1
rlabel polysilicon 184 -520 184 -520 0 3
rlabel polysilicon 191 -514 191 -514 0 1
rlabel polysilicon 191 -520 191 -520 0 3
rlabel polysilicon 198 -514 198 -514 0 1
rlabel polysilicon 201 -514 201 -514 0 2
rlabel polysilicon 198 -520 198 -520 0 3
rlabel polysilicon 201 -520 201 -520 0 4
rlabel polysilicon 205 -514 205 -514 0 1
rlabel polysilicon 205 -520 205 -520 0 3
rlabel polysilicon 212 -514 212 -514 0 1
rlabel polysilicon 212 -520 212 -520 0 3
rlabel polysilicon 219 -514 219 -514 0 1
rlabel polysilicon 219 -520 219 -520 0 3
rlabel polysilicon 226 -514 226 -514 0 1
rlabel polysilicon 226 -520 226 -520 0 3
rlabel polysilicon 233 -514 233 -514 0 1
rlabel polysilicon 233 -520 233 -520 0 3
rlabel polysilicon 240 -514 240 -514 0 1
rlabel polysilicon 240 -520 240 -520 0 3
rlabel polysilicon 247 -520 247 -520 0 3
rlabel polysilicon 250 -520 250 -520 0 4
rlabel polysilicon 254 -520 254 -520 0 3
rlabel polysilicon 257 -520 257 -520 0 4
rlabel polysilicon 261 -514 261 -514 0 1
rlabel polysilicon 261 -520 261 -520 0 3
rlabel polysilicon 268 -514 268 -514 0 1
rlabel polysilicon 268 -520 268 -520 0 3
rlabel polysilicon 275 -514 275 -514 0 1
rlabel polysilicon 275 -520 275 -520 0 3
rlabel polysilicon 282 -514 282 -514 0 1
rlabel polysilicon 282 -520 282 -520 0 3
rlabel polysilicon 289 -514 289 -514 0 1
rlabel polysilicon 289 -520 289 -520 0 3
rlabel polysilicon 296 -514 296 -514 0 1
rlabel polysilicon 296 -520 296 -520 0 3
rlabel polysilicon 303 -514 303 -514 0 1
rlabel polysilicon 303 -520 303 -520 0 3
rlabel polysilicon 310 -514 310 -514 0 1
rlabel polysilicon 310 -520 310 -520 0 3
rlabel polysilicon 317 -514 317 -514 0 1
rlabel polysilicon 317 -520 317 -520 0 3
rlabel polysilicon 324 -514 324 -514 0 1
rlabel polysilicon 324 -520 324 -520 0 3
rlabel polysilicon 331 -514 331 -514 0 1
rlabel polysilicon 331 -520 331 -520 0 3
rlabel polysilicon 338 -514 338 -514 0 1
rlabel polysilicon 338 -520 338 -520 0 3
rlabel polysilicon 345 -514 345 -514 0 1
rlabel polysilicon 345 -520 345 -520 0 3
rlabel polysilicon 352 -514 352 -514 0 1
rlabel polysilicon 352 -520 352 -520 0 3
rlabel polysilicon 359 -514 359 -514 0 1
rlabel polysilicon 359 -520 359 -520 0 3
rlabel polysilicon 366 -514 366 -514 0 1
rlabel polysilicon 366 -520 366 -520 0 3
rlabel polysilicon 373 -514 373 -514 0 1
rlabel polysilicon 373 -520 373 -520 0 3
rlabel polysilicon 380 -514 380 -514 0 1
rlabel polysilicon 383 -514 383 -514 0 2
rlabel polysilicon 380 -520 380 -520 0 3
rlabel polysilicon 383 -520 383 -520 0 4
rlabel polysilicon 387 -514 387 -514 0 1
rlabel polysilicon 387 -520 387 -520 0 3
rlabel polysilicon 394 -514 394 -514 0 1
rlabel polysilicon 394 -520 394 -520 0 3
rlabel polysilicon 401 -514 401 -514 0 1
rlabel polysilicon 401 -520 401 -520 0 3
rlabel polysilicon 408 -514 408 -514 0 1
rlabel polysilicon 408 -520 408 -520 0 3
rlabel polysilicon 415 -514 415 -514 0 1
rlabel polysilicon 415 -520 415 -520 0 3
rlabel polysilicon 418 -520 418 -520 0 4
rlabel polysilicon 422 -514 422 -514 0 1
rlabel polysilicon 425 -514 425 -514 0 2
rlabel polysilicon 422 -520 422 -520 0 3
rlabel polysilicon 425 -520 425 -520 0 4
rlabel polysilicon 429 -514 429 -514 0 1
rlabel polysilicon 429 -520 429 -520 0 3
rlabel polysilicon 436 -514 436 -514 0 1
rlabel polysilicon 436 -520 436 -520 0 3
rlabel polysilicon 443 -514 443 -514 0 1
rlabel polysilicon 443 -520 443 -520 0 3
rlabel polysilicon 450 -514 450 -514 0 1
rlabel polysilicon 450 -520 450 -520 0 3
rlabel polysilicon 457 -514 457 -514 0 1
rlabel polysilicon 460 -514 460 -514 0 2
rlabel polysilicon 457 -520 457 -520 0 3
rlabel polysilicon 460 -520 460 -520 0 4
rlabel polysilicon 464 -514 464 -514 0 1
rlabel polysilicon 464 -520 464 -520 0 3
rlabel polysilicon 471 -514 471 -514 0 1
rlabel polysilicon 471 -520 471 -520 0 3
rlabel polysilicon 478 -514 478 -514 0 1
rlabel polysilicon 478 -520 478 -520 0 3
rlabel polysilicon 485 -514 485 -514 0 1
rlabel polysilicon 485 -520 485 -520 0 3
rlabel polysilicon 492 -514 492 -514 0 1
rlabel polysilicon 492 -520 492 -520 0 3
rlabel polysilicon 499 -514 499 -514 0 1
rlabel polysilicon 502 -514 502 -514 0 2
rlabel polysilicon 499 -520 499 -520 0 3
rlabel polysilicon 502 -520 502 -520 0 4
rlabel polysilicon 506 -514 506 -514 0 1
rlabel polysilicon 509 -514 509 -514 0 2
rlabel polysilicon 506 -520 506 -520 0 3
rlabel polysilicon 509 -520 509 -520 0 4
rlabel polysilicon 513 -514 513 -514 0 1
rlabel polysilicon 513 -520 513 -520 0 3
rlabel polysilicon 520 -514 520 -514 0 1
rlabel polysilicon 520 -520 520 -520 0 3
rlabel polysilicon 527 -514 527 -514 0 1
rlabel polysilicon 530 -514 530 -514 0 2
rlabel polysilicon 530 -520 530 -520 0 4
rlabel polysilicon 534 -514 534 -514 0 1
rlabel polysilicon 537 -514 537 -514 0 2
rlabel polysilicon 534 -520 534 -520 0 3
rlabel polysilicon 541 -514 541 -514 0 1
rlabel polysilicon 541 -520 541 -520 0 3
rlabel polysilicon 548 -514 548 -514 0 1
rlabel polysilicon 548 -520 548 -520 0 3
rlabel polysilicon 555 -514 555 -514 0 1
rlabel polysilicon 555 -520 555 -520 0 3
rlabel polysilicon 562 -514 562 -514 0 1
rlabel polysilicon 562 -520 562 -520 0 3
rlabel polysilicon 569 -514 569 -514 0 1
rlabel polysilicon 569 -520 569 -520 0 3
rlabel polysilicon 576 -514 576 -514 0 1
rlabel polysilicon 576 -520 576 -520 0 3
rlabel polysilicon 583 -514 583 -514 0 1
rlabel polysilicon 583 -520 583 -520 0 3
rlabel polysilicon 590 -514 590 -514 0 1
rlabel polysilicon 590 -520 590 -520 0 3
rlabel polysilicon 597 -514 597 -514 0 1
rlabel polysilicon 600 -514 600 -514 0 2
rlabel polysilicon 597 -520 597 -520 0 3
rlabel polysilicon 600 -520 600 -520 0 4
rlabel polysilicon 604 -514 604 -514 0 1
rlabel polysilicon 604 -520 604 -520 0 3
rlabel polysilicon 611 -514 611 -514 0 1
rlabel polysilicon 614 -514 614 -514 0 2
rlabel polysilicon 611 -520 611 -520 0 3
rlabel polysilicon 614 -520 614 -520 0 4
rlabel polysilicon 618 -514 618 -514 0 1
rlabel polysilicon 618 -520 618 -520 0 3
rlabel polysilicon 625 -514 625 -514 0 1
rlabel polysilicon 625 -520 625 -520 0 3
rlabel polysilicon 632 -514 632 -514 0 1
rlabel polysilicon 632 -520 632 -520 0 3
rlabel polysilicon 639 -514 639 -514 0 1
rlabel polysilicon 639 -520 639 -520 0 3
rlabel polysilicon 646 -514 646 -514 0 1
rlabel polysilicon 646 -520 646 -520 0 3
rlabel polysilicon 653 -514 653 -514 0 1
rlabel polysilicon 653 -520 653 -520 0 3
rlabel polysilicon 660 -514 660 -514 0 1
rlabel polysilicon 663 -514 663 -514 0 2
rlabel polysilicon 660 -520 660 -520 0 3
rlabel polysilicon 663 -520 663 -520 0 4
rlabel polysilicon 667 -514 667 -514 0 1
rlabel polysilicon 667 -520 667 -520 0 3
rlabel polysilicon 674 -514 674 -514 0 1
rlabel polysilicon 674 -520 674 -520 0 3
rlabel polysilicon 681 -514 681 -514 0 1
rlabel polysilicon 681 -520 681 -520 0 3
rlabel polysilicon 688 -514 688 -514 0 1
rlabel polysilicon 688 -520 688 -520 0 3
rlabel polysilicon 698 -514 698 -514 0 2
rlabel polysilicon 695 -520 695 -520 0 3
rlabel polysilicon 698 -520 698 -520 0 4
rlabel polysilicon 702 -514 702 -514 0 1
rlabel polysilicon 705 -514 705 -514 0 2
rlabel polysilicon 702 -520 702 -520 0 3
rlabel polysilicon 705 -520 705 -520 0 4
rlabel polysilicon 709 -514 709 -514 0 1
rlabel polysilicon 709 -520 709 -520 0 3
rlabel polysilicon 716 -514 716 -514 0 1
rlabel polysilicon 716 -520 716 -520 0 3
rlabel polysilicon 723 -514 723 -514 0 1
rlabel polysilicon 723 -520 723 -520 0 3
rlabel polysilicon 730 -514 730 -514 0 1
rlabel polysilicon 730 -520 730 -520 0 3
rlabel polysilicon 737 -514 737 -514 0 1
rlabel polysilicon 737 -520 737 -520 0 3
rlabel polysilicon 744 -514 744 -514 0 1
rlabel polysilicon 744 -520 744 -520 0 3
rlabel polysilicon 751 -514 751 -514 0 1
rlabel polysilicon 751 -520 751 -520 0 3
rlabel polysilicon 758 -514 758 -514 0 1
rlabel polysilicon 758 -520 758 -520 0 3
rlabel polysilicon 765 -514 765 -514 0 1
rlabel polysilicon 765 -520 765 -520 0 3
rlabel polysilicon 772 -514 772 -514 0 1
rlabel polysilicon 772 -520 772 -520 0 3
rlabel polysilicon 779 -514 779 -514 0 1
rlabel polysilicon 779 -520 779 -520 0 3
rlabel polysilicon 786 -514 786 -514 0 1
rlabel polysilicon 786 -520 786 -520 0 3
rlabel polysilicon 793 -514 793 -514 0 1
rlabel polysilicon 793 -520 793 -520 0 3
rlabel polysilicon 800 -514 800 -514 0 1
rlabel polysilicon 800 -520 800 -520 0 3
rlabel polysilicon 807 -514 807 -514 0 1
rlabel polysilicon 807 -520 807 -520 0 3
rlabel polysilicon 814 -514 814 -514 0 1
rlabel polysilicon 814 -520 814 -520 0 3
rlabel polysilicon 821 -514 821 -514 0 1
rlabel polysilicon 821 -520 821 -520 0 3
rlabel polysilicon 828 -514 828 -514 0 1
rlabel polysilicon 828 -520 828 -520 0 3
rlabel polysilicon 835 -514 835 -514 0 1
rlabel polysilicon 835 -520 835 -520 0 3
rlabel polysilicon 842 -514 842 -514 0 1
rlabel polysilicon 842 -520 842 -520 0 3
rlabel polysilicon 849 -514 849 -514 0 1
rlabel polysilicon 849 -520 849 -520 0 3
rlabel polysilicon 856 -514 856 -514 0 1
rlabel polysilicon 856 -520 856 -520 0 3
rlabel polysilicon 863 -514 863 -514 0 1
rlabel polysilicon 863 -520 863 -520 0 3
rlabel polysilicon 870 -514 870 -514 0 1
rlabel polysilicon 870 -520 870 -520 0 3
rlabel polysilicon 877 -514 877 -514 0 1
rlabel polysilicon 877 -520 877 -520 0 3
rlabel polysilicon 884 -514 884 -514 0 1
rlabel polysilicon 884 -520 884 -520 0 3
rlabel polysilicon 891 -514 891 -514 0 1
rlabel polysilicon 891 -520 891 -520 0 3
rlabel polysilicon 898 -514 898 -514 0 1
rlabel polysilicon 898 -520 898 -520 0 3
rlabel polysilicon 905 -514 905 -514 0 1
rlabel polysilicon 905 -520 905 -520 0 3
rlabel polysilicon 912 -514 912 -514 0 1
rlabel polysilicon 912 -520 912 -520 0 3
rlabel polysilicon 919 -514 919 -514 0 1
rlabel polysilicon 919 -520 919 -520 0 3
rlabel polysilicon 926 -514 926 -514 0 1
rlabel polysilicon 926 -520 926 -520 0 3
rlabel polysilicon 933 -514 933 -514 0 1
rlabel polysilicon 933 -520 933 -520 0 3
rlabel polysilicon 940 -514 940 -514 0 1
rlabel polysilicon 940 -520 940 -520 0 3
rlabel polysilicon 947 -514 947 -514 0 1
rlabel polysilicon 947 -520 947 -520 0 3
rlabel polysilicon 954 -514 954 -514 0 1
rlabel polysilicon 954 -520 954 -520 0 3
rlabel polysilicon 961 -514 961 -514 0 1
rlabel polysilicon 961 -520 961 -520 0 3
rlabel polysilicon 968 -514 968 -514 0 1
rlabel polysilicon 968 -520 968 -520 0 3
rlabel polysilicon 975 -514 975 -514 0 1
rlabel polysilicon 975 -520 975 -520 0 3
rlabel polysilicon 982 -514 982 -514 0 1
rlabel polysilicon 982 -520 982 -520 0 3
rlabel polysilicon 989 -514 989 -514 0 1
rlabel polysilicon 989 -520 989 -520 0 3
rlabel polysilicon 996 -514 996 -514 0 1
rlabel polysilicon 996 -520 996 -520 0 3
rlabel polysilicon 1003 -514 1003 -514 0 1
rlabel polysilicon 1003 -520 1003 -520 0 3
rlabel polysilicon 1010 -514 1010 -514 0 1
rlabel polysilicon 1010 -520 1010 -520 0 3
rlabel polysilicon 1017 -514 1017 -514 0 1
rlabel polysilicon 1017 -520 1017 -520 0 3
rlabel polysilicon 1024 -514 1024 -514 0 1
rlabel polysilicon 1024 -520 1024 -520 0 3
rlabel polysilicon 1031 -514 1031 -514 0 1
rlabel polysilicon 1031 -520 1031 -520 0 3
rlabel polysilicon 1038 -514 1038 -514 0 1
rlabel polysilicon 1038 -520 1038 -520 0 3
rlabel polysilicon 1045 -514 1045 -514 0 1
rlabel polysilicon 1045 -520 1045 -520 0 3
rlabel polysilicon 1052 -514 1052 -514 0 1
rlabel polysilicon 1052 -520 1052 -520 0 3
rlabel polysilicon 1059 -514 1059 -514 0 1
rlabel polysilicon 1059 -520 1059 -520 0 3
rlabel polysilicon 1066 -514 1066 -514 0 1
rlabel polysilicon 1066 -520 1066 -520 0 3
rlabel polysilicon 1073 -514 1073 -514 0 1
rlabel polysilicon 1073 -520 1073 -520 0 3
rlabel polysilicon 1080 -514 1080 -514 0 1
rlabel polysilicon 1080 -520 1080 -520 0 3
rlabel polysilicon 1087 -514 1087 -514 0 1
rlabel polysilicon 1087 -520 1087 -520 0 3
rlabel polysilicon 1094 -514 1094 -514 0 1
rlabel polysilicon 1094 -520 1094 -520 0 3
rlabel polysilicon 1101 -514 1101 -514 0 1
rlabel polysilicon 1101 -520 1101 -520 0 3
rlabel polysilicon 1108 -514 1108 -514 0 1
rlabel polysilicon 1108 -520 1108 -520 0 3
rlabel polysilicon 1115 -514 1115 -514 0 1
rlabel polysilicon 1115 -520 1115 -520 0 3
rlabel polysilicon 1122 -514 1122 -514 0 1
rlabel polysilicon 1122 -520 1122 -520 0 3
rlabel polysilicon 1129 -514 1129 -514 0 1
rlabel polysilicon 1129 -520 1129 -520 0 3
rlabel polysilicon 1136 -514 1136 -514 0 1
rlabel polysilicon 1136 -520 1136 -520 0 3
rlabel polysilicon 1143 -514 1143 -514 0 1
rlabel polysilicon 1143 -520 1143 -520 0 3
rlabel polysilicon 1150 -514 1150 -514 0 1
rlabel polysilicon 1150 -520 1150 -520 0 3
rlabel polysilicon 1157 -514 1157 -514 0 1
rlabel polysilicon 1157 -520 1157 -520 0 3
rlabel polysilicon 1164 -514 1164 -514 0 1
rlabel polysilicon 1164 -520 1164 -520 0 3
rlabel polysilicon 1171 -514 1171 -514 0 1
rlabel polysilicon 1171 -520 1171 -520 0 3
rlabel polysilicon 1178 -514 1178 -514 0 1
rlabel polysilicon 1178 -520 1178 -520 0 3
rlabel polysilicon 1185 -514 1185 -514 0 1
rlabel polysilicon 1185 -520 1185 -520 0 3
rlabel polysilicon 1192 -514 1192 -514 0 1
rlabel polysilicon 1192 -520 1192 -520 0 3
rlabel polysilicon 1199 -514 1199 -514 0 1
rlabel polysilicon 1199 -520 1199 -520 0 3
rlabel polysilicon 1206 -514 1206 -514 0 1
rlabel polysilicon 1206 -520 1206 -520 0 3
rlabel polysilicon 1213 -514 1213 -514 0 1
rlabel polysilicon 1213 -520 1213 -520 0 3
rlabel polysilicon 1220 -514 1220 -514 0 1
rlabel polysilicon 1220 -520 1220 -520 0 3
rlabel polysilicon 1227 -514 1227 -514 0 1
rlabel polysilicon 1227 -520 1227 -520 0 3
rlabel polysilicon 1234 -514 1234 -514 0 1
rlabel polysilicon 1234 -520 1234 -520 0 3
rlabel polysilicon 1241 -514 1241 -514 0 1
rlabel polysilicon 1241 -520 1241 -520 0 3
rlabel polysilicon 1248 -514 1248 -514 0 1
rlabel polysilicon 1248 -520 1248 -520 0 3
rlabel polysilicon 1255 -514 1255 -514 0 1
rlabel polysilicon 1255 -520 1255 -520 0 3
rlabel polysilicon 1262 -514 1262 -514 0 1
rlabel polysilicon 1262 -520 1262 -520 0 3
rlabel polysilicon 1395 -514 1395 -514 0 1
rlabel polysilicon 1395 -520 1395 -520 0 3
rlabel polysilicon 1500 -514 1500 -514 0 1
rlabel polysilicon 1500 -520 1500 -520 0 3
rlabel polysilicon 2 -629 2 -629 0 1
rlabel polysilicon 2 -635 2 -635 0 3
rlabel polysilicon 9 -629 9 -629 0 1
rlabel polysilicon 9 -635 9 -635 0 3
rlabel polysilicon 19 -629 19 -629 0 2
rlabel polysilicon 16 -635 16 -635 0 3
rlabel polysilicon 19 -635 19 -635 0 4
rlabel polysilicon 23 -629 23 -629 0 1
rlabel polysilicon 23 -635 23 -635 0 3
rlabel polysilicon 30 -629 30 -629 0 1
rlabel polysilicon 30 -635 30 -635 0 3
rlabel polysilicon 37 -629 37 -629 0 1
rlabel polysilicon 40 -629 40 -629 0 2
rlabel polysilicon 44 -629 44 -629 0 1
rlabel polysilicon 47 -629 47 -629 0 2
rlabel polysilicon 44 -635 44 -635 0 3
rlabel polysilicon 47 -635 47 -635 0 4
rlabel polysilicon 51 -629 51 -629 0 1
rlabel polysilicon 51 -635 51 -635 0 3
rlabel polysilicon 58 -629 58 -629 0 1
rlabel polysilicon 58 -635 58 -635 0 3
rlabel polysilicon 65 -629 65 -629 0 1
rlabel polysilicon 65 -635 65 -635 0 3
rlabel polysilicon 72 -629 72 -629 0 1
rlabel polysilicon 75 -629 75 -629 0 2
rlabel polysilicon 72 -635 72 -635 0 3
rlabel polysilicon 75 -635 75 -635 0 4
rlabel polysilicon 79 -629 79 -629 0 1
rlabel polysilicon 79 -635 79 -635 0 3
rlabel polysilicon 86 -629 86 -629 0 1
rlabel polysilicon 86 -635 86 -635 0 3
rlabel polysilicon 93 -629 93 -629 0 1
rlabel polysilicon 96 -629 96 -629 0 2
rlabel polysilicon 93 -635 93 -635 0 3
rlabel polysilicon 96 -635 96 -635 0 4
rlabel polysilicon 100 -629 100 -629 0 1
rlabel polysilicon 100 -635 100 -635 0 3
rlabel polysilicon 107 -629 107 -629 0 1
rlabel polysilicon 107 -635 107 -635 0 3
rlabel polysilicon 114 -629 114 -629 0 1
rlabel polysilicon 117 -629 117 -629 0 2
rlabel polysilicon 114 -635 114 -635 0 3
rlabel polysilicon 117 -635 117 -635 0 4
rlabel polysilicon 121 -629 121 -629 0 1
rlabel polysilicon 121 -635 121 -635 0 3
rlabel polysilicon 128 -629 128 -629 0 1
rlabel polysilicon 128 -635 128 -635 0 3
rlabel polysilicon 135 -629 135 -629 0 1
rlabel polysilicon 135 -635 135 -635 0 3
rlabel polysilicon 142 -629 142 -629 0 1
rlabel polysilicon 142 -635 142 -635 0 3
rlabel polysilicon 149 -629 149 -629 0 1
rlabel polysilicon 149 -635 149 -635 0 3
rlabel polysilicon 156 -629 156 -629 0 1
rlabel polysilicon 156 -635 156 -635 0 3
rlabel polysilicon 163 -629 163 -629 0 1
rlabel polysilicon 163 -635 163 -635 0 3
rlabel polysilicon 170 -629 170 -629 0 1
rlabel polysilicon 170 -635 170 -635 0 3
rlabel polysilicon 173 -635 173 -635 0 4
rlabel polysilicon 177 -629 177 -629 0 1
rlabel polysilicon 177 -635 177 -635 0 3
rlabel polysilicon 184 -629 184 -629 0 1
rlabel polysilicon 184 -635 184 -635 0 3
rlabel polysilicon 191 -629 191 -629 0 1
rlabel polysilicon 191 -635 191 -635 0 3
rlabel polysilicon 198 -629 198 -629 0 1
rlabel polysilicon 198 -635 198 -635 0 3
rlabel polysilicon 205 -629 205 -629 0 1
rlabel polysilicon 205 -635 205 -635 0 3
rlabel polysilicon 212 -629 212 -629 0 1
rlabel polysilicon 212 -635 212 -635 0 3
rlabel polysilicon 219 -629 219 -629 0 1
rlabel polysilicon 219 -635 219 -635 0 3
rlabel polysilicon 226 -629 226 -629 0 1
rlabel polysilicon 226 -635 226 -635 0 3
rlabel polysilicon 233 -629 233 -629 0 1
rlabel polysilicon 233 -635 233 -635 0 3
rlabel polysilicon 240 -629 240 -629 0 1
rlabel polysilicon 240 -635 240 -635 0 3
rlabel polysilicon 247 -629 247 -629 0 1
rlabel polysilicon 247 -635 247 -635 0 3
rlabel polysilicon 254 -629 254 -629 0 1
rlabel polysilicon 254 -635 254 -635 0 3
rlabel polysilicon 261 -629 261 -629 0 1
rlabel polysilicon 261 -635 261 -635 0 3
rlabel polysilicon 268 -629 268 -629 0 1
rlabel polysilicon 271 -629 271 -629 0 2
rlabel polysilicon 271 -635 271 -635 0 4
rlabel polysilicon 275 -629 275 -629 0 1
rlabel polysilicon 275 -635 275 -635 0 3
rlabel polysilicon 282 -629 282 -629 0 1
rlabel polysilicon 282 -635 282 -635 0 3
rlabel polysilicon 289 -629 289 -629 0 1
rlabel polysilicon 289 -635 289 -635 0 3
rlabel polysilicon 296 -629 296 -629 0 1
rlabel polysilicon 296 -635 296 -635 0 3
rlabel polysilicon 303 -629 303 -629 0 1
rlabel polysilicon 303 -635 303 -635 0 3
rlabel polysilicon 310 -635 310 -635 0 3
rlabel polysilicon 313 -635 313 -635 0 4
rlabel polysilicon 317 -629 317 -629 0 1
rlabel polysilicon 317 -635 317 -635 0 3
rlabel polysilicon 324 -629 324 -629 0 1
rlabel polysilicon 324 -635 324 -635 0 3
rlabel polysilicon 331 -629 331 -629 0 1
rlabel polysilicon 331 -635 331 -635 0 3
rlabel polysilicon 338 -629 338 -629 0 1
rlabel polysilicon 338 -635 338 -635 0 3
rlabel polysilicon 348 -629 348 -629 0 2
rlabel polysilicon 345 -635 345 -635 0 3
rlabel polysilicon 348 -635 348 -635 0 4
rlabel polysilicon 352 -629 352 -629 0 1
rlabel polysilicon 355 -635 355 -635 0 4
rlabel polysilicon 359 -629 359 -629 0 1
rlabel polysilicon 359 -635 359 -635 0 3
rlabel polysilicon 366 -629 366 -629 0 1
rlabel polysilicon 366 -635 366 -635 0 3
rlabel polysilicon 373 -629 373 -629 0 1
rlabel polysilicon 373 -635 373 -635 0 3
rlabel polysilicon 380 -629 380 -629 0 1
rlabel polysilicon 380 -635 380 -635 0 3
rlabel polysilicon 383 -635 383 -635 0 4
rlabel polysilicon 387 -629 387 -629 0 1
rlabel polysilicon 390 -629 390 -629 0 2
rlabel polysilicon 387 -635 387 -635 0 3
rlabel polysilicon 390 -635 390 -635 0 4
rlabel polysilicon 394 -629 394 -629 0 1
rlabel polysilicon 394 -635 394 -635 0 3
rlabel polysilicon 401 -629 401 -629 0 1
rlabel polysilicon 401 -635 401 -635 0 3
rlabel polysilicon 408 -629 408 -629 0 1
rlabel polysilicon 408 -635 408 -635 0 3
rlabel polysilicon 415 -629 415 -629 0 1
rlabel polysilicon 418 -629 418 -629 0 2
rlabel polysilicon 415 -635 415 -635 0 3
rlabel polysilicon 418 -635 418 -635 0 4
rlabel polysilicon 422 -629 422 -629 0 1
rlabel polysilicon 422 -635 422 -635 0 3
rlabel polysilicon 429 -629 429 -629 0 1
rlabel polysilicon 429 -635 429 -635 0 3
rlabel polysilicon 436 -629 436 -629 0 1
rlabel polysilicon 436 -635 436 -635 0 3
rlabel polysilicon 443 -629 443 -629 0 1
rlabel polysilicon 446 -629 446 -629 0 2
rlabel polysilicon 443 -635 443 -635 0 3
rlabel polysilicon 446 -635 446 -635 0 4
rlabel polysilicon 450 -629 450 -629 0 1
rlabel polysilicon 450 -635 450 -635 0 3
rlabel polysilicon 457 -629 457 -629 0 1
rlabel polysilicon 457 -635 457 -635 0 3
rlabel polysilicon 464 -629 464 -629 0 1
rlabel polysilicon 464 -635 464 -635 0 3
rlabel polysilicon 471 -629 471 -629 0 1
rlabel polysilicon 471 -635 471 -635 0 3
rlabel polysilicon 481 -629 481 -629 0 2
rlabel polysilicon 478 -635 478 -635 0 3
rlabel polysilicon 481 -635 481 -635 0 4
rlabel polysilicon 485 -629 485 -629 0 1
rlabel polysilicon 485 -635 485 -635 0 3
rlabel polysilicon 492 -629 492 -629 0 1
rlabel polysilicon 492 -635 492 -635 0 3
rlabel polysilicon 499 -629 499 -629 0 1
rlabel polysilicon 499 -635 499 -635 0 3
rlabel polysilicon 506 -629 506 -629 0 1
rlabel polysilicon 509 -629 509 -629 0 2
rlabel polysilicon 506 -635 506 -635 0 3
rlabel polysilicon 509 -635 509 -635 0 4
rlabel polysilicon 513 -629 513 -629 0 1
rlabel polysilicon 513 -635 513 -635 0 3
rlabel polysilicon 520 -629 520 -629 0 1
rlabel polysilicon 520 -635 520 -635 0 3
rlabel polysilicon 527 -629 527 -629 0 1
rlabel polysilicon 527 -635 527 -635 0 3
rlabel polysilicon 534 -629 534 -629 0 1
rlabel polysilicon 534 -635 534 -635 0 3
rlabel polysilicon 541 -629 541 -629 0 1
rlabel polysilicon 541 -635 541 -635 0 3
rlabel polysilicon 548 -629 548 -629 0 1
rlabel polysilicon 548 -635 548 -635 0 3
rlabel polysilicon 555 -629 555 -629 0 1
rlabel polysilicon 555 -635 555 -635 0 3
rlabel polysilicon 562 -629 562 -629 0 1
rlabel polysilicon 565 -629 565 -629 0 2
rlabel polysilicon 562 -635 562 -635 0 3
rlabel polysilicon 569 -629 569 -629 0 1
rlabel polysilicon 569 -635 569 -635 0 3
rlabel polysilicon 576 -629 576 -629 0 1
rlabel polysilicon 576 -635 576 -635 0 3
rlabel polysilicon 583 -629 583 -629 0 1
rlabel polysilicon 583 -635 583 -635 0 3
rlabel polysilicon 590 -629 590 -629 0 1
rlabel polysilicon 590 -635 590 -635 0 3
rlabel polysilicon 597 -629 597 -629 0 1
rlabel polysilicon 597 -635 597 -635 0 3
rlabel polysilicon 604 -629 604 -629 0 1
rlabel polysilicon 604 -635 604 -635 0 3
rlabel polysilicon 611 -629 611 -629 0 1
rlabel polysilicon 614 -629 614 -629 0 2
rlabel polysilicon 611 -635 611 -635 0 3
rlabel polysilicon 614 -635 614 -635 0 4
rlabel polysilicon 618 -629 618 -629 0 1
rlabel polysilicon 618 -635 618 -635 0 3
rlabel polysilicon 625 -629 625 -629 0 1
rlabel polysilicon 628 -629 628 -629 0 2
rlabel polysilicon 625 -635 625 -635 0 3
rlabel polysilicon 628 -635 628 -635 0 4
rlabel polysilicon 632 -629 632 -629 0 1
rlabel polysilicon 635 -629 635 -629 0 2
rlabel polysilicon 632 -635 632 -635 0 3
rlabel polysilicon 635 -635 635 -635 0 4
rlabel polysilicon 639 -629 639 -629 0 1
rlabel polysilicon 639 -635 639 -635 0 3
rlabel polysilicon 646 -629 646 -629 0 1
rlabel polysilicon 646 -635 646 -635 0 3
rlabel polysilicon 653 -629 653 -629 0 1
rlabel polysilicon 653 -635 653 -635 0 3
rlabel polysilicon 660 -629 660 -629 0 1
rlabel polysilicon 660 -635 660 -635 0 3
rlabel polysilicon 667 -629 667 -629 0 1
rlabel polysilicon 670 -629 670 -629 0 2
rlabel polysilicon 667 -635 667 -635 0 3
rlabel polysilicon 674 -629 674 -629 0 1
rlabel polysilicon 674 -635 674 -635 0 3
rlabel polysilicon 681 -629 681 -629 0 1
rlabel polysilicon 681 -635 681 -635 0 3
rlabel polysilicon 688 -629 688 -629 0 1
rlabel polysilicon 688 -635 688 -635 0 3
rlabel polysilicon 695 -629 695 -629 0 1
rlabel polysilicon 695 -635 695 -635 0 3
rlabel polysilicon 702 -629 702 -629 0 1
rlabel polysilicon 702 -635 702 -635 0 3
rlabel polysilicon 709 -629 709 -629 0 1
rlabel polysilicon 709 -635 709 -635 0 3
rlabel polysilicon 716 -629 716 -629 0 1
rlabel polysilicon 716 -635 716 -635 0 3
rlabel polysilicon 723 -629 723 -629 0 1
rlabel polysilicon 723 -635 723 -635 0 3
rlabel polysilicon 730 -629 730 -629 0 1
rlabel polysilicon 730 -635 730 -635 0 3
rlabel polysilicon 737 -629 737 -629 0 1
rlabel polysilicon 737 -635 737 -635 0 3
rlabel polysilicon 747 -629 747 -629 0 2
rlabel polysilicon 744 -635 744 -635 0 3
rlabel polysilicon 747 -635 747 -635 0 4
rlabel polysilicon 751 -629 751 -629 0 1
rlabel polysilicon 751 -635 751 -635 0 3
rlabel polysilicon 758 -629 758 -629 0 1
rlabel polysilicon 758 -635 758 -635 0 3
rlabel polysilicon 765 -629 765 -629 0 1
rlabel polysilicon 765 -635 765 -635 0 3
rlabel polysilicon 772 -629 772 -629 0 1
rlabel polysilicon 772 -635 772 -635 0 3
rlabel polysilicon 779 -629 779 -629 0 1
rlabel polysilicon 779 -635 779 -635 0 3
rlabel polysilicon 786 -629 786 -629 0 1
rlabel polysilicon 786 -635 786 -635 0 3
rlabel polysilicon 793 -629 793 -629 0 1
rlabel polysilicon 793 -635 793 -635 0 3
rlabel polysilicon 800 -629 800 -629 0 1
rlabel polysilicon 800 -635 800 -635 0 3
rlabel polysilicon 807 -629 807 -629 0 1
rlabel polysilicon 807 -635 807 -635 0 3
rlabel polysilicon 814 -629 814 -629 0 1
rlabel polysilicon 814 -635 814 -635 0 3
rlabel polysilicon 821 -629 821 -629 0 1
rlabel polysilicon 821 -635 821 -635 0 3
rlabel polysilicon 828 -629 828 -629 0 1
rlabel polysilicon 828 -635 828 -635 0 3
rlabel polysilicon 835 -629 835 -629 0 1
rlabel polysilicon 835 -635 835 -635 0 3
rlabel polysilicon 842 -629 842 -629 0 1
rlabel polysilicon 842 -635 842 -635 0 3
rlabel polysilicon 849 -629 849 -629 0 1
rlabel polysilicon 849 -635 849 -635 0 3
rlabel polysilicon 856 -629 856 -629 0 1
rlabel polysilicon 856 -635 856 -635 0 3
rlabel polysilicon 863 -629 863 -629 0 1
rlabel polysilicon 863 -635 863 -635 0 3
rlabel polysilicon 870 -629 870 -629 0 1
rlabel polysilicon 870 -635 870 -635 0 3
rlabel polysilicon 877 -629 877 -629 0 1
rlabel polysilicon 877 -635 877 -635 0 3
rlabel polysilicon 884 -629 884 -629 0 1
rlabel polysilicon 884 -635 884 -635 0 3
rlabel polysilicon 891 -629 891 -629 0 1
rlabel polysilicon 891 -635 891 -635 0 3
rlabel polysilicon 898 -629 898 -629 0 1
rlabel polysilicon 898 -635 898 -635 0 3
rlabel polysilicon 905 -629 905 -629 0 1
rlabel polysilicon 905 -635 905 -635 0 3
rlabel polysilicon 912 -629 912 -629 0 1
rlabel polysilicon 912 -635 912 -635 0 3
rlabel polysilicon 919 -629 919 -629 0 1
rlabel polysilicon 919 -635 919 -635 0 3
rlabel polysilicon 926 -629 926 -629 0 1
rlabel polysilicon 926 -635 926 -635 0 3
rlabel polysilicon 933 -629 933 -629 0 1
rlabel polysilicon 933 -635 933 -635 0 3
rlabel polysilicon 940 -629 940 -629 0 1
rlabel polysilicon 940 -635 940 -635 0 3
rlabel polysilicon 947 -629 947 -629 0 1
rlabel polysilicon 947 -635 947 -635 0 3
rlabel polysilicon 954 -629 954 -629 0 1
rlabel polysilicon 954 -635 954 -635 0 3
rlabel polysilicon 961 -629 961 -629 0 1
rlabel polysilicon 961 -635 961 -635 0 3
rlabel polysilicon 964 -635 964 -635 0 4
rlabel polysilicon 968 -629 968 -629 0 1
rlabel polysilicon 968 -635 968 -635 0 3
rlabel polysilicon 975 -629 975 -629 0 1
rlabel polysilicon 975 -635 975 -635 0 3
rlabel polysilicon 982 -629 982 -629 0 1
rlabel polysilicon 982 -635 982 -635 0 3
rlabel polysilicon 989 -629 989 -629 0 1
rlabel polysilicon 989 -635 989 -635 0 3
rlabel polysilicon 996 -629 996 -629 0 1
rlabel polysilicon 996 -635 996 -635 0 3
rlabel polysilicon 1003 -629 1003 -629 0 1
rlabel polysilicon 1003 -635 1003 -635 0 3
rlabel polysilicon 1010 -629 1010 -629 0 1
rlabel polysilicon 1010 -635 1010 -635 0 3
rlabel polysilicon 1017 -629 1017 -629 0 1
rlabel polysilicon 1017 -635 1017 -635 0 3
rlabel polysilicon 1024 -629 1024 -629 0 1
rlabel polysilicon 1024 -635 1024 -635 0 3
rlabel polysilicon 1031 -629 1031 -629 0 1
rlabel polysilicon 1034 -629 1034 -629 0 2
rlabel polysilicon 1034 -635 1034 -635 0 4
rlabel polysilicon 1038 -629 1038 -629 0 1
rlabel polysilicon 1038 -635 1038 -635 0 3
rlabel polysilicon 1045 -629 1045 -629 0 1
rlabel polysilicon 1045 -635 1045 -635 0 3
rlabel polysilicon 1052 -629 1052 -629 0 1
rlabel polysilicon 1052 -635 1052 -635 0 3
rlabel polysilicon 1059 -629 1059 -629 0 1
rlabel polysilicon 1059 -635 1059 -635 0 3
rlabel polysilicon 1066 -629 1066 -629 0 1
rlabel polysilicon 1066 -635 1066 -635 0 3
rlabel polysilicon 1073 -629 1073 -629 0 1
rlabel polysilicon 1073 -635 1073 -635 0 3
rlabel polysilicon 1080 -629 1080 -629 0 1
rlabel polysilicon 1080 -635 1080 -635 0 3
rlabel polysilicon 1087 -629 1087 -629 0 1
rlabel polysilicon 1087 -635 1087 -635 0 3
rlabel polysilicon 1094 -629 1094 -629 0 1
rlabel polysilicon 1094 -635 1094 -635 0 3
rlabel polysilicon 1101 -629 1101 -629 0 1
rlabel polysilicon 1101 -635 1101 -635 0 3
rlabel polysilicon 1108 -629 1108 -629 0 1
rlabel polysilicon 1108 -635 1108 -635 0 3
rlabel polysilicon 1115 -629 1115 -629 0 1
rlabel polysilicon 1115 -635 1115 -635 0 3
rlabel polysilicon 1122 -629 1122 -629 0 1
rlabel polysilicon 1122 -635 1122 -635 0 3
rlabel polysilicon 1129 -629 1129 -629 0 1
rlabel polysilicon 1129 -635 1129 -635 0 3
rlabel polysilicon 1136 -629 1136 -629 0 1
rlabel polysilicon 1136 -635 1136 -635 0 3
rlabel polysilicon 1143 -629 1143 -629 0 1
rlabel polysilicon 1143 -635 1143 -635 0 3
rlabel polysilicon 1150 -629 1150 -629 0 1
rlabel polysilicon 1150 -635 1150 -635 0 3
rlabel polysilicon 1157 -629 1157 -629 0 1
rlabel polysilicon 1157 -635 1157 -635 0 3
rlabel polysilicon 1164 -629 1164 -629 0 1
rlabel polysilicon 1164 -635 1164 -635 0 3
rlabel polysilicon 1171 -629 1171 -629 0 1
rlabel polysilicon 1171 -635 1171 -635 0 3
rlabel polysilicon 1178 -629 1178 -629 0 1
rlabel polysilicon 1178 -635 1178 -635 0 3
rlabel polysilicon 1185 -629 1185 -629 0 1
rlabel polysilicon 1185 -635 1185 -635 0 3
rlabel polysilicon 1192 -629 1192 -629 0 1
rlabel polysilicon 1192 -635 1192 -635 0 3
rlabel polysilicon 1199 -629 1199 -629 0 1
rlabel polysilicon 1199 -635 1199 -635 0 3
rlabel polysilicon 1206 -629 1206 -629 0 1
rlabel polysilicon 1206 -635 1206 -635 0 3
rlabel polysilicon 1213 -629 1213 -629 0 1
rlabel polysilicon 1213 -635 1213 -635 0 3
rlabel polysilicon 1220 -629 1220 -629 0 1
rlabel polysilicon 1220 -635 1220 -635 0 3
rlabel polysilicon 1227 -629 1227 -629 0 1
rlabel polysilicon 1227 -635 1227 -635 0 3
rlabel polysilicon 1234 -629 1234 -629 0 1
rlabel polysilicon 1234 -635 1234 -635 0 3
rlabel polysilicon 1241 -629 1241 -629 0 1
rlabel polysilicon 1241 -635 1241 -635 0 3
rlabel polysilicon 1248 -629 1248 -629 0 1
rlabel polysilicon 1248 -635 1248 -635 0 3
rlabel polysilicon 1255 -629 1255 -629 0 1
rlabel polysilicon 1255 -635 1255 -635 0 3
rlabel polysilicon 1262 -629 1262 -629 0 1
rlabel polysilicon 1262 -635 1262 -635 0 3
rlabel polysilicon 1269 -629 1269 -629 0 1
rlabel polysilicon 1269 -635 1269 -635 0 3
rlabel polysilicon 1276 -629 1276 -629 0 1
rlabel polysilicon 1276 -635 1276 -635 0 3
rlabel polysilicon 1283 -629 1283 -629 0 1
rlabel polysilicon 1283 -635 1283 -635 0 3
rlabel polysilicon 1290 -629 1290 -629 0 1
rlabel polysilicon 1290 -635 1290 -635 0 3
rlabel polysilicon 1297 -629 1297 -629 0 1
rlabel polysilicon 1297 -635 1297 -635 0 3
rlabel polysilicon 1304 -629 1304 -629 0 1
rlabel polysilicon 1304 -635 1304 -635 0 3
rlabel polysilicon 1311 -629 1311 -629 0 1
rlabel polysilicon 1311 -635 1311 -635 0 3
rlabel polysilicon 1318 -629 1318 -629 0 1
rlabel polysilicon 1318 -635 1318 -635 0 3
rlabel polysilicon 1325 -629 1325 -629 0 1
rlabel polysilicon 1325 -635 1325 -635 0 3
rlabel polysilicon 1332 -629 1332 -629 0 1
rlabel polysilicon 1332 -635 1332 -635 0 3
rlabel polysilicon 1339 -629 1339 -629 0 1
rlabel polysilicon 1339 -635 1339 -635 0 3
rlabel polysilicon 1346 -629 1346 -629 0 1
rlabel polysilicon 1346 -635 1346 -635 0 3
rlabel polysilicon 1353 -629 1353 -629 0 1
rlabel polysilicon 1353 -635 1353 -635 0 3
rlabel polysilicon 1360 -629 1360 -629 0 1
rlabel polysilicon 1360 -635 1360 -635 0 3
rlabel polysilicon 1367 -629 1367 -629 0 1
rlabel polysilicon 1367 -635 1367 -635 0 3
rlabel polysilicon 1374 -629 1374 -629 0 1
rlabel polysilicon 1374 -635 1374 -635 0 3
rlabel polysilicon 1472 -629 1472 -629 0 1
rlabel polysilicon 1472 -635 1472 -635 0 3
rlabel polysilicon 1507 -629 1507 -629 0 1
rlabel polysilicon 1507 -635 1507 -635 0 3
rlabel polysilicon 5 -748 5 -748 0 2
rlabel polysilicon 2 -754 2 -754 0 3
rlabel polysilicon 12 -748 12 -748 0 2
rlabel polysilicon 9 -754 9 -754 0 3
rlabel polysilicon 12 -754 12 -754 0 4
rlabel polysilicon 16 -748 16 -748 0 1
rlabel polysilicon 16 -754 16 -754 0 3
rlabel polysilicon 23 -748 23 -748 0 1
rlabel polysilicon 23 -754 23 -754 0 3
rlabel polysilicon 30 -748 30 -748 0 1
rlabel polysilicon 30 -754 30 -754 0 3
rlabel polysilicon 37 -748 37 -748 0 1
rlabel polysilicon 37 -754 37 -754 0 3
rlabel polysilicon 44 -748 44 -748 0 1
rlabel polysilicon 44 -754 44 -754 0 3
rlabel polysilicon 51 -748 51 -748 0 1
rlabel polysilicon 51 -754 51 -754 0 3
rlabel polysilicon 58 -748 58 -748 0 1
rlabel polysilicon 61 -748 61 -748 0 2
rlabel polysilicon 58 -754 58 -754 0 3
rlabel polysilicon 61 -754 61 -754 0 4
rlabel polysilicon 65 -748 65 -748 0 1
rlabel polysilicon 65 -754 65 -754 0 3
rlabel polysilicon 72 -748 72 -748 0 1
rlabel polysilicon 75 -748 75 -748 0 2
rlabel polysilicon 72 -754 72 -754 0 3
rlabel polysilicon 75 -754 75 -754 0 4
rlabel polysilicon 79 -748 79 -748 0 1
rlabel polysilicon 79 -754 79 -754 0 3
rlabel polysilicon 86 -748 86 -748 0 1
rlabel polysilicon 86 -754 86 -754 0 3
rlabel polysilicon 93 -748 93 -748 0 1
rlabel polysilicon 93 -754 93 -754 0 3
rlabel polysilicon 100 -748 100 -748 0 1
rlabel polysilicon 103 -748 103 -748 0 2
rlabel polysilicon 100 -754 100 -754 0 3
rlabel polysilicon 103 -754 103 -754 0 4
rlabel polysilicon 107 -748 107 -748 0 1
rlabel polysilicon 107 -754 107 -754 0 3
rlabel polysilicon 114 -748 114 -748 0 1
rlabel polysilicon 117 -748 117 -748 0 2
rlabel polysilicon 114 -754 114 -754 0 3
rlabel polysilicon 117 -754 117 -754 0 4
rlabel polysilicon 121 -748 121 -748 0 1
rlabel polysilicon 121 -754 121 -754 0 3
rlabel polysilicon 128 -748 128 -748 0 1
rlabel polysilicon 128 -754 128 -754 0 3
rlabel polysilicon 135 -754 135 -754 0 3
rlabel polysilicon 138 -754 138 -754 0 4
rlabel polysilicon 142 -748 142 -748 0 1
rlabel polysilicon 142 -754 142 -754 0 3
rlabel polysilicon 149 -748 149 -748 0 1
rlabel polysilicon 149 -754 149 -754 0 3
rlabel polysilicon 156 -748 156 -748 0 1
rlabel polysilicon 156 -754 156 -754 0 3
rlabel polysilicon 163 -748 163 -748 0 1
rlabel polysilicon 163 -754 163 -754 0 3
rlabel polysilicon 170 -748 170 -748 0 1
rlabel polysilicon 170 -754 170 -754 0 3
rlabel polysilicon 177 -748 177 -748 0 1
rlabel polysilicon 177 -754 177 -754 0 3
rlabel polysilicon 184 -748 184 -748 0 1
rlabel polysilicon 184 -754 184 -754 0 3
rlabel polysilicon 191 -748 191 -748 0 1
rlabel polysilicon 191 -754 191 -754 0 3
rlabel polysilicon 198 -748 198 -748 0 1
rlabel polysilicon 198 -754 198 -754 0 3
rlabel polysilicon 205 -748 205 -748 0 1
rlabel polysilicon 205 -754 205 -754 0 3
rlabel polysilicon 212 -748 212 -748 0 1
rlabel polysilicon 212 -754 212 -754 0 3
rlabel polysilicon 219 -748 219 -748 0 1
rlabel polysilicon 219 -754 219 -754 0 3
rlabel polysilicon 226 -748 226 -748 0 1
rlabel polysilicon 226 -754 226 -754 0 3
rlabel polysilicon 233 -748 233 -748 0 1
rlabel polysilicon 233 -754 233 -754 0 3
rlabel polysilicon 240 -748 240 -748 0 1
rlabel polysilicon 240 -754 240 -754 0 3
rlabel polysilicon 247 -748 247 -748 0 1
rlabel polysilicon 247 -754 247 -754 0 3
rlabel polysilicon 254 -748 254 -748 0 1
rlabel polysilicon 254 -754 254 -754 0 3
rlabel polysilicon 261 -748 261 -748 0 1
rlabel polysilicon 261 -754 261 -754 0 3
rlabel polysilicon 268 -748 268 -748 0 1
rlabel polysilicon 271 -748 271 -748 0 2
rlabel polysilicon 268 -754 268 -754 0 3
rlabel polysilicon 271 -754 271 -754 0 4
rlabel polysilicon 275 -748 275 -748 0 1
rlabel polysilicon 275 -754 275 -754 0 3
rlabel polysilicon 282 -748 282 -748 0 1
rlabel polysilicon 282 -754 282 -754 0 3
rlabel polysilicon 289 -748 289 -748 0 1
rlabel polysilicon 289 -754 289 -754 0 3
rlabel polysilicon 296 -748 296 -748 0 1
rlabel polysilicon 296 -754 296 -754 0 3
rlabel polysilicon 303 -748 303 -748 0 1
rlabel polysilicon 303 -754 303 -754 0 3
rlabel polysilicon 310 -748 310 -748 0 1
rlabel polysilicon 310 -754 310 -754 0 3
rlabel polysilicon 317 -748 317 -748 0 1
rlabel polysilicon 317 -754 317 -754 0 3
rlabel polysilicon 324 -748 324 -748 0 1
rlabel polysilicon 324 -754 324 -754 0 3
rlabel polysilicon 331 -748 331 -748 0 1
rlabel polysilicon 331 -754 331 -754 0 3
rlabel polysilicon 338 -748 338 -748 0 1
rlabel polysilicon 338 -754 338 -754 0 3
rlabel polysilicon 345 -748 345 -748 0 1
rlabel polysilicon 345 -754 345 -754 0 3
rlabel polysilicon 352 -748 352 -748 0 1
rlabel polysilicon 355 -748 355 -748 0 2
rlabel polysilicon 352 -754 352 -754 0 3
rlabel polysilicon 355 -754 355 -754 0 4
rlabel polysilicon 359 -748 359 -748 0 1
rlabel polysilicon 359 -754 359 -754 0 3
rlabel polysilicon 366 -748 366 -748 0 1
rlabel polysilicon 366 -754 366 -754 0 3
rlabel polysilicon 369 -754 369 -754 0 4
rlabel polysilicon 373 -748 373 -748 0 1
rlabel polysilicon 373 -754 373 -754 0 3
rlabel polysilicon 380 -748 380 -748 0 1
rlabel polysilicon 380 -754 380 -754 0 3
rlabel polysilicon 387 -748 387 -748 0 1
rlabel polysilicon 387 -754 387 -754 0 3
rlabel polysilicon 394 -748 394 -748 0 1
rlabel polysilicon 394 -754 394 -754 0 3
rlabel polysilicon 401 -748 401 -748 0 1
rlabel polysilicon 401 -754 401 -754 0 3
rlabel polysilicon 408 -748 408 -748 0 1
rlabel polysilicon 408 -754 408 -754 0 3
rlabel polysilicon 415 -748 415 -748 0 1
rlabel polysilicon 422 -748 422 -748 0 1
rlabel polysilicon 425 -748 425 -748 0 2
rlabel polysilicon 422 -754 422 -754 0 3
rlabel polysilicon 425 -754 425 -754 0 4
rlabel polysilicon 429 -748 429 -748 0 1
rlabel polysilicon 429 -754 429 -754 0 3
rlabel polysilicon 436 -748 436 -748 0 1
rlabel polysilicon 436 -754 436 -754 0 3
rlabel polysilicon 443 -748 443 -748 0 1
rlabel polysilicon 443 -754 443 -754 0 3
rlabel polysilicon 450 -748 450 -748 0 1
rlabel polysilicon 450 -754 450 -754 0 3
rlabel polysilicon 457 -748 457 -748 0 1
rlabel polysilicon 457 -754 457 -754 0 3
rlabel polysilicon 464 -748 464 -748 0 1
rlabel polysilicon 464 -754 464 -754 0 3
rlabel polysilicon 471 -748 471 -748 0 1
rlabel polysilicon 471 -754 471 -754 0 3
rlabel polysilicon 478 -748 478 -748 0 1
rlabel polysilicon 478 -754 478 -754 0 3
rlabel polysilicon 485 -748 485 -748 0 1
rlabel polysilicon 485 -754 485 -754 0 3
rlabel polysilicon 492 -748 492 -748 0 1
rlabel polysilicon 492 -754 492 -754 0 3
rlabel polysilicon 499 -748 499 -748 0 1
rlabel polysilicon 499 -754 499 -754 0 3
rlabel polysilicon 506 -748 506 -748 0 1
rlabel polysilicon 506 -754 506 -754 0 3
rlabel polysilicon 513 -748 513 -748 0 1
rlabel polysilicon 513 -754 513 -754 0 3
rlabel polysilicon 523 -748 523 -748 0 2
rlabel polysilicon 520 -754 520 -754 0 3
rlabel polysilicon 523 -754 523 -754 0 4
rlabel polysilicon 527 -748 527 -748 0 1
rlabel polysilicon 527 -754 527 -754 0 3
rlabel polysilicon 530 -754 530 -754 0 4
rlabel polysilicon 534 -748 534 -748 0 1
rlabel polysilicon 537 -748 537 -748 0 2
rlabel polysilicon 534 -754 534 -754 0 3
rlabel polysilicon 537 -754 537 -754 0 4
rlabel polysilicon 541 -748 541 -748 0 1
rlabel polysilicon 544 -748 544 -748 0 2
rlabel polysilicon 541 -754 541 -754 0 3
rlabel polysilicon 544 -754 544 -754 0 4
rlabel polysilicon 548 -748 548 -748 0 1
rlabel polysilicon 548 -754 548 -754 0 3
rlabel polysilicon 555 -748 555 -748 0 1
rlabel polysilicon 555 -754 555 -754 0 3
rlabel polysilicon 562 -748 562 -748 0 1
rlabel polysilicon 565 -748 565 -748 0 2
rlabel polysilicon 562 -754 562 -754 0 3
rlabel polysilicon 569 -748 569 -748 0 1
rlabel polysilicon 569 -754 569 -754 0 3
rlabel polysilicon 576 -748 576 -748 0 1
rlabel polysilicon 576 -754 576 -754 0 3
rlabel polysilicon 583 -748 583 -748 0 1
rlabel polysilicon 583 -754 583 -754 0 3
rlabel polysilicon 590 -748 590 -748 0 1
rlabel polysilicon 590 -754 590 -754 0 3
rlabel polysilicon 600 -748 600 -748 0 2
rlabel polysilicon 597 -754 597 -754 0 3
rlabel polysilicon 600 -754 600 -754 0 4
rlabel polysilicon 604 -748 604 -748 0 1
rlabel polysilicon 604 -754 604 -754 0 3
rlabel polysilicon 611 -748 611 -748 0 1
rlabel polysilicon 614 -748 614 -748 0 2
rlabel polysilicon 611 -754 611 -754 0 3
rlabel polysilicon 614 -754 614 -754 0 4
rlabel polysilicon 618 -748 618 -748 0 1
rlabel polysilicon 621 -748 621 -748 0 2
rlabel polysilicon 618 -754 618 -754 0 3
rlabel polysilicon 628 -748 628 -748 0 2
rlabel polysilicon 625 -754 625 -754 0 3
rlabel polysilicon 632 -748 632 -748 0 1
rlabel polysilicon 632 -754 632 -754 0 3
rlabel polysilicon 639 -748 639 -748 0 1
rlabel polysilicon 639 -754 639 -754 0 3
rlabel polysilicon 646 -748 646 -748 0 1
rlabel polysilicon 646 -754 646 -754 0 3
rlabel polysilicon 653 -748 653 -748 0 1
rlabel polysilicon 653 -754 653 -754 0 3
rlabel polysilicon 660 -748 660 -748 0 1
rlabel polysilicon 663 -748 663 -748 0 2
rlabel polysilicon 660 -754 660 -754 0 3
rlabel polysilicon 663 -754 663 -754 0 4
rlabel polysilicon 667 -748 667 -748 0 1
rlabel polysilicon 667 -754 667 -754 0 3
rlabel polysilicon 674 -748 674 -748 0 1
rlabel polysilicon 674 -754 674 -754 0 3
rlabel polysilicon 681 -748 681 -748 0 1
rlabel polysilicon 681 -754 681 -754 0 3
rlabel polysilicon 688 -748 688 -748 0 1
rlabel polysilicon 688 -754 688 -754 0 3
rlabel polysilicon 695 -748 695 -748 0 1
rlabel polysilicon 695 -754 695 -754 0 3
rlabel polysilicon 702 -748 702 -748 0 1
rlabel polysilicon 702 -754 702 -754 0 3
rlabel polysilicon 709 -748 709 -748 0 1
rlabel polysilicon 709 -754 709 -754 0 3
rlabel polysilicon 716 -748 716 -748 0 1
rlabel polysilicon 716 -754 716 -754 0 3
rlabel polysilicon 723 -748 723 -748 0 1
rlabel polysilicon 723 -754 723 -754 0 3
rlabel polysilicon 730 -748 730 -748 0 1
rlabel polysilicon 730 -754 730 -754 0 3
rlabel polysilicon 737 -748 737 -748 0 1
rlabel polysilicon 737 -754 737 -754 0 3
rlabel polysilicon 744 -748 744 -748 0 1
rlabel polysilicon 747 -748 747 -748 0 2
rlabel polysilicon 744 -754 744 -754 0 3
rlabel polysilicon 747 -754 747 -754 0 4
rlabel polysilicon 751 -748 751 -748 0 1
rlabel polysilicon 751 -754 751 -754 0 3
rlabel polysilicon 758 -748 758 -748 0 1
rlabel polysilicon 761 -748 761 -748 0 2
rlabel polysilicon 758 -754 758 -754 0 3
rlabel polysilicon 761 -754 761 -754 0 4
rlabel polysilicon 765 -748 765 -748 0 1
rlabel polysilicon 765 -754 765 -754 0 3
rlabel polysilicon 772 -748 772 -748 0 1
rlabel polysilicon 772 -754 772 -754 0 3
rlabel polysilicon 775 -754 775 -754 0 4
rlabel polysilicon 779 -748 779 -748 0 1
rlabel polysilicon 779 -754 779 -754 0 3
rlabel polysilicon 786 -748 786 -748 0 1
rlabel polysilicon 786 -754 786 -754 0 3
rlabel polysilicon 793 -748 793 -748 0 1
rlabel polysilicon 793 -754 793 -754 0 3
rlabel polysilicon 800 -748 800 -748 0 1
rlabel polysilicon 800 -754 800 -754 0 3
rlabel polysilicon 807 -748 807 -748 0 1
rlabel polysilicon 807 -754 807 -754 0 3
rlabel polysilicon 814 -748 814 -748 0 1
rlabel polysilicon 814 -754 814 -754 0 3
rlabel polysilicon 821 -748 821 -748 0 1
rlabel polysilicon 821 -754 821 -754 0 3
rlabel polysilicon 828 -748 828 -748 0 1
rlabel polysilicon 828 -754 828 -754 0 3
rlabel polysilicon 835 -748 835 -748 0 1
rlabel polysilicon 835 -754 835 -754 0 3
rlabel polysilicon 842 -748 842 -748 0 1
rlabel polysilicon 842 -754 842 -754 0 3
rlabel polysilicon 849 -748 849 -748 0 1
rlabel polysilicon 849 -754 849 -754 0 3
rlabel polysilicon 856 -748 856 -748 0 1
rlabel polysilicon 856 -754 856 -754 0 3
rlabel polysilicon 863 -748 863 -748 0 1
rlabel polysilicon 863 -754 863 -754 0 3
rlabel polysilicon 870 -748 870 -748 0 1
rlabel polysilicon 870 -754 870 -754 0 3
rlabel polysilicon 877 -748 877 -748 0 1
rlabel polysilicon 877 -754 877 -754 0 3
rlabel polysilicon 884 -748 884 -748 0 1
rlabel polysilicon 887 -748 887 -748 0 2
rlabel polysilicon 884 -754 884 -754 0 3
rlabel polysilicon 887 -754 887 -754 0 4
rlabel polysilicon 891 -748 891 -748 0 1
rlabel polysilicon 891 -754 891 -754 0 3
rlabel polysilicon 898 -748 898 -748 0 1
rlabel polysilicon 898 -754 898 -754 0 3
rlabel polysilicon 905 -748 905 -748 0 1
rlabel polysilicon 905 -754 905 -754 0 3
rlabel polysilicon 912 -748 912 -748 0 1
rlabel polysilicon 912 -754 912 -754 0 3
rlabel polysilicon 919 -748 919 -748 0 1
rlabel polysilicon 919 -754 919 -754 0 3
rlabel polysilicon 926 -748 926 -748 0 1
rlabel polysilicon 926 -754 926 -754 0 3
rlabel polysilicon 933 -748 933 -748 0 1
rlabel polysilicon 933 -754 933 -754 0 3
rlabel polysilicon 940 -748 940 -748 0 1
rlabel polysilicon 943 -748 943 -748 0 2
rlabel polysilicon 940 -754 940 -754 0 3
rlabel polysilicon 943 -754 943 -754 0 4
rlabel polysilicon 947 -748 947 -748 0 1
rlabel polysilicon 947 -754 947 -754 0 3
rlabel polysilicon 954 -748 954 -748 0 1
rlabel polysilicon 954 -754 954 -754 0 3
rlabel polysilicon 961 -748 961 -748 0 1
rlabel polysilicon 961 -754 961 -754 0 3
rlabel polysilicon 968 -748 968 -748 0 1
rlabel polysilicon 968 -754 968 -754 0 3
rlabel polysilicon 975 -748 975 -748 0 1
rlabel polysilicon 975 -754 975 -754 0 3
rlabel polysilicon 982 -748 982 -748 0 1
rlabel polysilicon 982 -754 982 -754 0 3
rlabel polysilicon 989 -748 989 -748 0 1
rlabel polysilicon 989 -754 989 -754 0 3
rlabel polysilicon 996 -748 996 -748 0 1
rlabel polysilicon 996 -754 996 -754 0 3
rlabel polysilicon 1003 -748 1003 -748 0 1
rlabel polysilicon 1003 -754 1003 -754 0 3
rlabel polysilicon 1010 -748 1010 -748 0 1
rlabel polysilicon 1010 -754 1010 -754 0 3
rlabel polysilicon 1017 -748 1017 -748 0 1
rlabel polysilicon 1017 -754 1017 -754 0 3
rlabel polysilicon 1024 -748 1024 -748 0 1
rlabel polysilicon 1024 -754 1024 -754 0 3
rlabel polysilicon 1031 -748 1031 -748 0 1
rlabel polysilicon 1031 -754 1031 -754 0 3
rlabel polysilicon 1038 -748 1038 -748 0 1
rlabel polysilicon 1038 -754 1038 -754 0 3
rlabel polysilicon 1045 -748 1045 -748 0 1
rlabel polysilicon 1045 -754 1045 -754 0 3
rlabel polysilicon 1052 -748 1052 -748 0 1
rlabel polysilicon 1052 -754 1052 -754 0 3
rlabel polysilicon 1059 -748 1059 -748 0 1
rlabel polysilicon 1059 -754 1059 -754 0 3
rlabel polysilicon 1066 -748 1066 -748 0 1
rlabel polysilicon 1066 -754 1066 -754 0 3
rlabel polysilicon 1073 -748 1073 -748 0 1
rlabel polysilicon 1073 -754 1073 -754 0 3
rlabel polysilicon 1080 -748 1080 -748 0 1
rlabel polysilicon 1080 -754 1080 -754 0 3
rlabel polysilicon 1087 -748 1087 -748 0 1
rlabel polysilicon 1087 -754 1087 -754 0 3
rlabel polysilicon 1094 -748 1094 -748 0 1
rlabel polysilicon 1094 -754 1094 -754 0 3
rlabel polysilicon 1101 -748 1101 -748 0 1
rlabel polysilicon 1101 -754 1101 -754 0 3
rlabel polysilicon 1108 -748 1108 -748 0 1
rlabel polysilicon 1108 -754 1108 -754 0 3
rlabel polysilicon 1115 -748 1115 -748 0 1
rlabel polysilicon 1115 -754 1115 -754 0 3
rlabel polysilicon 1122 -748 1122 -748 0 1
rlabel polysilicon 1122 -754 1122 -754 0 3
rlabel polysilicon 1129 -748 1129 -748 0 1
rlabel polysilicon 1129 -754 1129 -754 0 3
rlabel polysilicon 1136 -748 1136 -748 0 1
rlabel polysilicon 1136 -754 1136 -754 0 3
rlabel polysilicon 1143 -748 1143 -748 0 1
rlabel polysilicon 1143 -754 1143 -754 0 3
rlabel polysilicon 1150 -748 1150 -748 0 1
rlabel polysilicon 1150 -754 1150 -754 0 3
rlabel polysilicon 1157 -748 1157 -748 0 1
rlabel polysilicon 1157 -754 1157 -754 0 3
rlabel polysilicon 1164 -748 1164 -748 0 1
rlabel polysilicon 1164 -754 1164 -754 0 3
rlabel polysilicon 1171 -748 1171 -748 0 1
rlabel polysilicon 1171 -754 1171 -754 0 3
rlabel polysilicon 1178 -748 1178 -748 0 1
rlabel polysilicon 1178 -754 1178 -754 0 3
rlabel polysilicon 1185 -748 1185 -748 0 1
rlabel polysilicon 1185 -754 1185 -754 0 3
rlabel polysilicon 1192 -748 1192 -748 0 1
rlabel polysilicon 1192 -754 1192 -754 0 3
rlabel polysilicon 1199 -748 1199 -748 0 1
rlabel polysilicon 1199 -754 1199 -754 0 3
rlabel polysilicon 1206 -748 1206 -748 0 1
rlabel polysilicon 1206 -754 1206 -754 0 3
rlabel polysilicon 1213 -748 1213 -748 0 1
rlabel polysilicon 1213 -754 1213 -754 0 3
rlabel polysilicon 1220 -748 1220 -748 0 1
rlabel polysilicon 1220 -754 1220 -754 0 3
rlabel polysilicon 1227 -748 1227 -748 0 1
rlabel polysilicon 1227 -754 1227 -754 0 3
rlabel polysilicon 1234 -748 1234 -748 0 1
rlabel polysilicon 1234 -754 1234 -754 0 3
rlabel polysilicon 1241 -748 1241 -748 0 1
rlabel polysilicon 1241 -754 1241 -754 0 3
rlabel polysilicon 1248 -748 1248 -748 0 1
rlabel polysilicon 1248 -754 1248 -754 0 3
rlabel polysilicon 1255 -748 1255 -748 0 1
rlabel polysilicon 1255 -754 1255 -754 0 3
rlabel polysilicon 1262 -748 1262 -748 0 1
rlabel polysilicon 1262 -754 1262 -754 0 3
rlabel polysilicon 1269 -748 1269 -748 0 1
rlabel polysilicon 1269 -754 1269 -754 0 3
rlabel polysilicon 1276 -748 1276 -748 0 1
rlabel polysilicon 1276 -754 1276 -754 0 3
rlabel polysilicon 1283 -748 1283 -748 0 1
rlabel polysilicon 1283 -754 1283 -754 0 3
rlabel polysilicon 1290 -748 1290 -748 0 1
rlabel polysilicon 1290 -754 1290 -754 0 3
rlabel polysilicon 1297 -748 1297 -748 0 1
rlabel polysilicon 1297 -754 1297 -754 0 3
rlabel polysilicon 1304 -748 1304 -748 0 1
rlabel polysilicon 1304 -754 1304 -754 0 3
rlabel polysilicon 1311 -748 1311 -748 0 1
rlabel polysilicon 1311 -754 1311 -754 0 3
rlabel polysilicon 1318 -748 1318 -748 0 1
rlabel polysilicon 1318 -754 1318 -754 0 3
rlabel polysilicon 1325 -748 1325 -748 0 1
rlabel polysilicon 1325 -754 1325 -754 0 3
rlabel polysilicon 1332 -748 1332 -748 0 1
rlabel polysilicon 1332 -754 1332 -754 0 3
rlabel polysilicon 1339 -748 1339 -748 0 1
rlabel polysilicon 1339 -754 1339 -754 0 3
rlabel polysilicon 1346 -748 1346 -748 0 1
rlabel polysilicon 1346 -754 1346 -754 0 3
rlabel polysilicon 1353 -748 1353 -748 0 1
rlabel polysilicon 1353 -754 1353 -754 0 3
rlabel polysilicon 1360 -748 1360 -748 0 1
rlabel polysilicon 1360 -754 1360 -754 0 3
rlabel polysilicon 1367 -748 1367 -748 0 1
rlabel polysilicon 1367 -754 1367 -754 0 3
rlabel polysilicon 1374 -748 1374 -748 0 1
rlabel polysilicon 1374 -754 1374 -754 0 3
rlabel polysilicon 1381 -748 1381 -748 0 1
rlabel polysilicon 1381 -754 1381 -754 0 3
rlabel polysilicon 1388 -748 1388 -748 0 1
rlabel polysilicon 1388 -754 1388 -754 0 3
rlabel polysilicon 1395 -748 1395 -748 0 1
rlabel polysilicon 1395 -754 1395 -754 0 3
rlabel polysilicon 1402 -748 1402 -748 0 1
rlabel polysilicon 1402 -754 1402 -754 0 3
rlabel polysilicon 1409 -748 1409 -748 0 1
rlabel polysilicon 1409 -754 1409 -754 0 3
rlabel polysilicon 1416 -748 1416 -748 0 1
rlabel polysilicon 1416 -754 1416 -754 0 3
rlabel polysilicon 1423 -748 1423 -748 0 1
rlabel polysilicon 1423 -754 1423 -754 0 3
rlabel polysilicon 1430 -748 1430 -748 0 1
rlabel polysilicon 1430 -754 1430 -754 0 3
rlabel polysilicon 1437 -748 1437 -748 0 1
rlabel polysilicon 1437 -754 1437 -754 0 3
rlabel polysilicon 1444 -748 1444 -748 0 1
rlabel polysilicon 1444 -754 1444 -754 0 3
rlabel polysilicon 1451 -748 1451 -748 0 1
rlabel polysilicon 1451 -754 1451 -754 0 3
rlabel polysilicon 1458 -748 1458 -748 0 1
rlabel polysilicon 1458 -754 1458 -754 0 3
rlabel polysilicon 1465 -748 1465 -748 0 1
rlabel polysilicon 1465 -754 1465 -754 0 3
rlabel polysilicon 1472 -748 1472 -748 0 1
rlabel polysilicon 1472 -754 1472 -754 0 3
rlabel polysilicon 1479 -748 1479 -748 0 1
rlabel polysilicon 1479 -754 1479 -754 0 3
rlabel polysilicon 1486 -748 1486 -748 0 1
rlabel polysilicon 1486 -754 1486 -754 0 3
rlabel polysilicon 1493 -748 1493 -748 0 1
rlabel polysilicon 1493 -754 1493 -754 0 3
rlabel polysilicon 1500 -748 1500 -748 0 1
rlabel polysilicon 1500 -754 1500 -754 0 3
rlabel polysilicon 1507 -748 1507 -748 0 1
rlabel polysilicon 1507 -754 1507 -754 0 3
rlabel polysilicon 1514 -748 1514 -748 0 1
rlabel polysilicon 1514 -754 1514 -754 0 3
rlabel polysilicon 1521 -748 1521 -748 0 1
rlabel polysilicon 1521 -754 1521 -754 0 3
rlabel polysilicon 1528 -748 1528 -748 0 1
rlabel polysilicon 1528 -754 1528 -754 0 3
rlabel polysilicon 2 -889 2 -889 0 1
rlabel polysilicon 2 -895 2 -895 0 3
rlabel polysilicon 9 -889 9 -889 0 1
rlabel polysilicon 9 -895 9 -895 0 3
rlabel polysilicon 16 -889 16 -889 0 1
rlabel polysilicon 16 -895 16 -895 0 3
rlabel polysilicon 23 -889 23 -889 0 1
rlabel polysilicon 23 -895 23 -895 0 3
rlabel polysilicon 30 -889 30 -889 0 1
rlabel polysilicon 30 -895 30 -895 0 3
rlabel polysilicon 40 -889 40 -889 0 2
rlabel polysilicon 37 -895 37 -895 0 3
rlabel polysilicon 40 -895 40 -895 0 4
rlabel polysilicon 44 -889 44 -889 0 1
rlabel polysilicon 47 -889 47 -889 0 2
rlabel polysilicon 44 -895 44 -895 0 3
rlabel polysilicon 51 -889 51 -889 0 1
rlabel polysilicon 51 -895 51 -895 0 3
rlabel polysilicon 58 -889 58 -889 0 1
rlabel polysilicon 58 -895 58 -895 0 3
rlabel polysilicon 65 -889 65 -889 0 1
rlabel polysilicon 65 -895 65 -895 0 3
rlabel polysilicon 72 -889 72 -889 0 1
rlabel polysilicon 72 -895 72 -895 0 3
rlabel polysilicon 79 -889 79 -889 0 1
rlabel polysilicon 79 -895 79 -895 0 3
rlabel polysilicon 86 -889 86 -889 0 1
rlabel polysilicon 86 -895 86 -895 0 3
rlabel polysilicon 93 -889 93 -889 0 1
rlabel polysilicon 93 -895 93 -895 0 3
rlabel polysilicon 100 -889 100 -889 0 1
rlabel polysilicon 100 -895 100 -895 0 3
rlabel polysilicon 107 -889 107 -889 0 1
rlabel polysilicon 107 -895 107 -895 0 3
rlabel polysilicon 114 -889 114 -889 0 1
rlabel polysilicon 114 -895 114 -895 0 3
rlabel polysilicon 121 -889 121 -889 0 1
rlabel polysilicon 121 -895 121 -895 0 3
rlabel polysilicon 128 -889 128 -889 0 1
rlabel polysilicon 131 -889 131 -889 0 2
rlabel polysilicon 128 -895 128 -895 0 3
rlabel polysilicon 131 -895 131 -895 0 4
rlabel polysilicon 135 -889 135 -889 0 1
rlabel polysilicon 135 -895 135 -895 0 3
rlabel polysilicon 142 -889 142 -889 0 1
rlabel polysilicon 142 -895 142 -895 0 3
rlabel polysilicon 149 -889 149 -889 0 1
rlabel polysilicon 149 -895 149 -895 0 3
rlabel polysilicon 156 -889 156 -889 0 1
rlabel polysilicon 156 -895 156 -895 0 3
rlabel polysilicon 163 -889 163 -889 0 1
rlabel polysilicon 166 -889 166 -889 0 2
rlabel polysilicon 163 -895 163 -895 0 3
rlabel polysilicon 170 -889 170 -889 0 1
rlabel polysilicon 170 -895 170 -895 0 3
rlabel polysilicon 177 -889 177 -889 0 1
rlabel polysilicon 177 -895 177 -895 0 3
rlabel polysilicon 184 -889 184 -889 0 1
rlabel polysilicon 184 -895 184 -895 0 3
rlabel polysilicon 191 -889 191 -889 0 1
rlabel polysilicon 191 -895 191 -895 0 3
rlabel polysilicon 198 -889 198 -889 0 1
rlabel polysilicon 198 -895 198 -895 0 3
rlabel polysilicon 205 -889 205 -889 0 1
rlabel polysilicon 205 -895 205 -895 0 3
rlabel polysilicon 212 -889 212 -889 0 1
rlabel polysilicon 212 -895 212 -895 0 3
rlabel polysilicon 219 -889 219 -889 0 1
rlabel polysilicon 219 -895 219 -895 0 3
rlabel polysilicon 226 -889 226 -889 0 1
rlabel polysilicon 226 -895 226 -895 0 3
rlabel polysilicon 233 -889 233 -889 0 1
rlabel polysilicon 236 -889 236 -889 0 2
rlabel polysilicon 233 -895 233 -895 0 3
rlabel polysilicon 236 -895 236 -895 0 4
rlabel polysilicon 240 -889 240 -889 0 1
rlabel polysilicon 240 -895 240 -895 0 3
rlabel polysilicon 247 -889 247 -889 0 1
rlabel polysilicon 247 -895 247 -895 0 3
rlabel polysilicon 254 -889 254 -889 0 1
rlabel polysilicon 254 -895 254 -895 0 3
rlabel polysilicon 261 -889 261 -889 0 1
rlabel polysilicon 261 -895 261 -895 0 3
rlabel polysilicon 268 -889 268 -889 0 1
rlabel polysilicon 268 -895 268 -895 0 3
rlabel polysilicon 275 -889 275 -889 0 1
rlabel polysilicon 275 -895 275 -895 0 3
rlabel polysilicon 282 -889 282 -889 0 1
rlabel polysilicon 282 -895 282 -895 0 3
rlabel polysilicon 289 -889 289 -889 0 1
rlabel polysilicon 289 -895 289 -895 0 3
rlabel polysilicon 296 -889 296 -889 0 1
rlabel polysilicon 296 -895 296 -895 0 3
rlabel polysilicon 303 -889 303 -889 0 1
rlabel polysilicon 303 -895 303 -895 0 3
rlabel polysilicon 310 -889 310 -889 0 1
rlabel polysilicon 310 -895 310 -895 0 3
rlabel polysilicon 317 -889 317 -889 0 1
rlabel polysilicon 317 -895 317 -895 0 3
rlabel polysilicon 324 -889 324 -889 0 1
rlabel polysilicon 324 -895 324 -895 0 3
rlabel polysilicon 331 -889 331 -889 0 1
rlabel polysilicon 331 -895 331 -895 0 3
rlabel polysilicon 338 -889 338 -889 0 1
rlabel polysilicon 338 -895 338 -895 0 3
rlabel polysilicon 345 -889 345 -889 0 1
rlabel polysilicon 345 -895 345 -895 0 3
rlabel polysilicon 352 -889 352 -889 0 1
rlabel polysilicon 352 -895 352 -895 0 3
rlabel polysilicon 359 -889 359 -889 0 1
rlabel polysilicon 359 -895 359 -895 0 3
rlabel polysilicon 366 -889 366 -889 0 1
rlabel polysilicon 369 -889 369 -889 0 2
rlabel polysilicon 366 -895 366 -895 0 3
rlabel polysilicon 369 -895 369 -895 0 4
rlabel polysilicon 373 -889 373 -889 0 1
rlabel polysilicon 373 -895 373 -895 0 3
rlabel polysilicon 380 -889 380 -889 0 1
rlabel polysilicon 380 -895 380 -895 0 3
rlabel polysilicon 387 -889 387 -889 0 1
rlabel polysilicon 387 -895 387 -895 0 3
rlabel polysilicon 394 -889 394 -889 0 1
rlabel polysilicon 394 -895 394 -895 0 3
rlabel polysilicon 401 -889 401 -889 0 1
rlabel polysilicon 401 -895 401 -895 0 3
rlabel polysilicon 408 -889 408 -889 0 1
rlabel polysilicon 408 -895 408 -895 0 3
rlabel polysilicon 415 -895 415 -895 0 3
rlabel polysilicon 422 -889 422 -889 0 1
rlabel polysilicon 422 -895 422 -895 0 3
rlabel polysilicon 429 -889 429 -889 0 1
rlabel polysilicon 429 -895 429 -895 0 3
rlabel polysilicon 436 -889 436 -889 0 1
rlabel polysilicon 439 -889 439 -889 0 2
rlabel polysilicon 436 -895 436 -895 0 3
rlabel polysilicon 443 -889 443 -889 0 1
rlabel polysilicon 443 -895 443 -895 0 3
rlabel polysilicon 450 -889 450 -889 0 1
rlabel polysilicon 450 -895 450 -895 0 3
rlabel polysilicon 457 -889 457 -889 0 1
rlabel polysilicon 460 -889 460 -889 0 2
rlabel polysilicon 457 -895 457 -895 0 3
rlabel polysilicon 460 -895 460 -895 0 4
rlabel polysilicon 464 -889 464 -889 0 1
rlabel polysilicon 467 -889 467 -889 0 2
rlabel polysilicon 464 -895 464 -895 0 3
rlabel polysilicon 467 -895 467 -895 0 4
rlabel polysilicon 471 -889 471 -889 0 1
rlabel polysilicon 471 -895 471 -895 0 3
rlabel polysilicon 478 -889 478 -889 0 1
rlabel polysilicon 478 -895 478 -895 0 3
rlabel polysilicon 485 -889 485 -889 0 1
rlabel polysilicon 485 -895 485 -895 0 3
rlabel polysilicon 492 -889 492 -889 0 1
rlabel polysilicon 492 -895 492 -895 0 3
rlabel polysilicon 499 -889 499 -889 0 1
rlabel polysilicon 499 -895 499 -895 0 3
rlabel polysilicon 506 -889 506 -889 0 1
rlabel polysilicon 509 -889 509 -889 0 2
rlabel polysilicon 506 -895 506 -895 0 3
rlabel polysilicon 509 -895 509 -895 0 4
rlabel polysilicon 513 -889 513 -889 0 1
rlabel polysilicon 513 -895 513 -895 0 3
rlabel polysilicon 520 -889 520 -889 0 1
rlabel polysilicon 520 -895 520 -895 0 3
rlabel polysilicon 527 -889 527 -889 0 1
rlabel polysilicon 530 -889 530 -889 0 2
rlabel polysilicon 527 -895 527 -895 0 3
rlabel polysilicon 534 -889 534 -889 0 1
rlabel polysilicon 537 -889 537 -889 0 2
rlabel polysilicon 534 -895 534 -895 0 3
rlabel polysilicon 537 -895 537 -895 0 4
rlabel polysilicon 541 -889 541 -889 0 1
rlabel polysilicon 541 -895 541 -895 0 3
rlabel polysilicon 544 -895 544 -895 0 4
rlabel polysilicon 548 -889 548 -889 0 1
rlabel polysilicon 551 -889 551 -889 0 2
rlabel polysilicon 548 -895 548 -895 0 3
rlabel polysilicon 551 -895 551 -895 0 4
rlabel polysilicon 555 -889 555 -889 0 1
rlabel polysilicon 555 -895 555 -895 0 3
rlabel polysilicon 562 -889 562 -889 0 1
rlabel polysilicon 562 -895 562 -895 0 3
rlabel polysilicon 569 -889 569 -889 0 1
rlabel polysilicon 569 -895 569 -895 0 3
rlabel polysilicon 576 -889 576 -889 0 1
rlabel polysilicon 576 -895 576 -895 0 3
rlabel polysilicon 583 -889 583 -889 0 1
rlabel polysilicon 583 -895 583 -895 0 3
rlabel polysilicon 590 -889 590 -889 0 1
rlabel polysilicon 590 -895 590 -895 0 3
rlabel polysilicon 597 -889 597 -889 0 1
rlabel polysilicon 597 -895 597 -895 0 3
rlabel polysilicon 604 -889 604 -889 0 1
rlabel polysilicon 604 -895 604 -895 0 3
rlabel polysilicon 611 -889 611 -889 0 1
rlabel polysilicon 611 -895 611 -895 0 3
rlabel polysilicon 618 -889 618 -889 0 1
rlabel polysilicon 618 -895 618 -895 0 3
rlabel polysilicon 625 -889 625 -889 0 1
rlabel polysilicon 625 -895 625 -895 0 3
rlabel polysilicon 632 -889 632 -889 0 1
rlabel polysilicon 632 -895 632 -895 0 3
rlabel polysilicon 639 -889 639 -889 0 1
rlabel polysilicon 642 -889 642 -889 0 2
rlabel polysilicon 639 -895 639 -895 0 3
rlabel polysilicon 642 -895 642 -895 0 4
rlabel polysilicon 646 -889 646 -889 0 1
rlabel polysilicon 649 -889 649 -889 0 2
rlabel polysilicon 646 -895 646 -895 0 3
rlabel polysilicon 649 -895 649 -895 0 4
rlabel polysilicon 653 -889 653 -889 0 1
rlabel polysilicon 656 -889 656 -889 0 2
rlabel polysilicon 653 -895 653 -895 0 3
rlabel polysilicon 656 -895 656 -895 0 4
rlabel polysilicon 660 -889 660 -889 0 1
rlabel polysilicon 663 -889 663 -889 0 2
rlabel polysilicon 660 -895 660 -895 0 3
rlabel polysilicon 667 -889 667 -889 0 1
rlabel polysilicon 667 -895 667 -895 0 3
rlabel polysilicon 674 -889 674 -889 0 1
rlabel polysilicon 674 -895 674 -895 0 3
rlabel polysilicon 681 -889 681 -889 0 1
rlabel polysilicon 681 -895 681 -895 0 3
rlabel polysilicon 691 -889 691 -889 0 2
rlabel polysilicon 688 -895 688 -895 0 3
rlabel polysilicon 691 -895 691 -895 0 4
rlabel polysilicon 695 -889 695 -889 0 1
rlabel polysilicon 695 -895 695 -895 0 3
rlabel polysilicon 702 -889 702 -889 0 1
rlabel polysilicon 702 -895 702 -895 0 3
rlabel polysilicon 709 -889 709 -889 0 1
rlabel polysilicon 712 -889 712 -889 0 2
rlabel polysilicon 709 -895 709 -895 0 3
rlabel polysilicon 712 -895 712 -895 0 4
rlabel polysilicon 716 -889 716 -889 0 1
rlabel polysilicon 716 -895 716 -895 0 3
rlabel polysilicon 723 -889 723 -889 0 1
rlabel polysilicon 723 -895 723 -895 0 3
rlabel polysilicon 730 -889 730 -889 0 1
rlabel polysilicon 730 -895 730 -895 0 3
rlabel polysilicon 737 -889 737 -889 0 1
rlabel polysilicon 737 -895 737 -895 0 3
rlabel polysilicon 744 -889 744 -889 0 1
rlabel polysilicon 744 -895 744 -895 0 3
rlabel polysilicon 751 -889 751 -889 0 1
rlabel polysilicon 751 -895 751 -895 0 3
rlabel polysilicon 758 -889 758 -889 0 1
rlabel polysilicon 758 -895 758 -895 0 3
rlabel polysilicon 765 -889 765 -889 0 1
rlabel polysilicon 768 -889 768 -889 0 2
rlabel polysilicon 765 -895 765 -895 0 3
rlabel polysilicon 768 -895 768 -895 0 4
rlabel polysilicon 772 -889 772 -889 0 1
rlabel polysilicon 772 -895 772 -895 0 3
rlabel polysilicon 779 -889 779 -889 0 1
rlabel polysilicon 779 -895 779 -895 0 3
rlabel polysilicon 786 -889 786 -889 0 1
rlabel polysilicon 786 -895 786 -895 0 3
rlabel polysilicon 793 -889 793 -889 0 1
rlabel polysilicon 793 -895 793 -895 0 3
rlabel polysilicon 800 -889 800 -889 0 1
rlabel polysilicon 800 -895 800 -895 0 3
rlabel polysilicon 807 -889 807 -889 0 1
rlabel polysilicon 807 -895 807 -895 0 3
rlabel polysilicon 810 -895 810 -895 0 4
rlabel polysilicon 814 -889 814 -889 0 1
rlabel polysilicon 814 -895 814 -895 0 3
rlabel polysilicon 821 -889 821 -889 0 1
rlabel polysilicon 821 -895 821 -895 0 3
rlabel polysilicon 828 -889 828 -889 0 1
rlabel polysilicon 828 -895 828 -895 0 3
rlabel polysilicon 835 -889 835 -889 0 1
rlabel polysilicon 838 -889 838 -889 0 2
rlabel polysilicon 835 -895 835 -895 0 3
rlabel polysilicon 838 -895 838 -895 0 4
rlabel polysilicon 842 -889 842 -889 0 1
rlabel polysilicon 842 -895 842 -895 0 3
rlabel polysilicon 849 -889 849 -889 0 1
rlabel polysilicon 849 -895 849 -895 0 3
rlabel polysilicon 856 -889 856 -889 0 1
rlabel polysilicon 856 -895 856 -895 0 3
rlabel polysilicon 863 -889 863 -889 0 1
rlabel polysilicon 863 -895 863 -895 0 3
rlabel polysilicon 870 -889 870 -889 0 1
rlabel polysilicon 870 -895 870 -895 0 3
rlabel polysilicon 877 -889 877 -889 0 1
rlabel polysilicon 877 -895 877 -895 0 3
rlabel polysilicon 884 -889 884 -889 0 1
rlabel polysilicon 884 -895 884 -895 0 3
rlabel polysilicon 891 -889 891 -889 0 1
rlabel polysilicon 891 -895 891 -895 0 3
rlabel polysilicon 898 -889 898 -889 0 1
rlabel polysilicon 898 -895 898 -895 0 3
rlabel polysilicon 905 -889 905 -889 0 1
rlabel polysilicon 905 -895 905 -895 0 3
rlabel polysilicon 912 -889 912 -889 0 1
rlabel polysilicon 912 -895 912 -895 0 3
rlabel polysilicon 919 -889 919 -889 0 1
rlabel polysilicon 919 -895 919 -895 0 3
rlabel polysilicon 926 -889 926 -889 0 1
rlabel polysilicon 926 -895 926 -895 0 3
rlabel polysilicon 933 -889 933 -889 0 1
rlabel polysilicon 933 -895 933 -895 0 3
rlabel polysilicon 943 -889 943 -889 0 2
rlabel polysilicon 943 -895 943 -895 0 4
rlabel polysilicon 947 -889 947 -889 0 1
rlabel polysilicon 947 -895 947 -895 0 3
rlabel polysilicon 954 -889 954 -889 0 1
rlabel polysilicon 954 -895 954 -895 0 3
rlabel polysilicon 961 -889 961 -889 0 1
rlabel polysilicon 961 -895 961 -895 0 3
rlabel polysilicon 968 -889 968 -889 0 1
rlabel polysilicon 968 -895 968 -895 0 3
rlabel polysilicon 975 -889 975 -889 0 1
rlabel polysilicon 975 -895 975 -895 0 3
rlabel polysilicon 982 -889 982 -889 0 1
rlabel polysilicon 989 -889 989 -889 0 1
rlabel polysilicon 989 -895 989 -895 0 3
rlabel polysilicon 996 -889 996 -889 0 1
rlabel polysilicon 999 -889 999 -889 0 2
rlabel polysilicon 996 -895 996 -895 0 3
rlabel polysilicon 1003 -889 1003 -889 0 1
rlabel polysilicon 1003 -895 1003 -895 0 3
rlabel polysilicon 1010 -889 1010 -889 0 1
rlabel polysilicon 1010 -895 1010 -895 0 3
rlabel polysilicon 1017 -889 1017 -889 0 1
rlabel polysilicon 1017 -895 1017 -895 0 3
rlabel polysilicon 1024 -889 1024 -889 0 1
rlabel polysilicon 1024 -895 1024 -895 0 3
rlabel polysilicon 1031 -889 1031 -889 0 1
rlabel polysilicon 1031 -895 1031 -895 0 3
rlabel polysilicon 1038 -889 1038 -889 0 1
rlabel polysilicon 1038 -895 1038 -895 0 3
rlabel polysilicon 1045 -889 1045 -889 0 1
rlabel polysilicon 1045 -895 1045 -895 0 3
rlabel polysilicon 1052 -889 1052 -889 0 1
rlabel polysilicon 1052 -895 1052 -895 0 3
rlabel polysilicon 1059 -889 1059 -889 0 1
rlabel polysilicon 1059 -895 1059 -895 0 3
rlabel polysilicon 1066 -889 1066 -889 0 1
rlabel polysilicon 1066 -895 1066 -895 0 3
rlabel polysilicon 1069 -895 1069 -895 0 4
rlabel polysilicon 1073 -889 1073 -889 0 1
rlabel polysilicon 1073 -895 1073 -895 0 3
rlabel polysilicon 1080 -889 1080 -889 0 1
rlabel polysilicon 1080 -895 1080 -895 0 3
rlabel polysilicon 1087 -889 1087 -889 0 1
rlabel polysilicon 1087 -895 1087 -895 0 3
rlabel polysilicon 1094 -889 1094 -889 0 1
rlabel polysilicon 1094 -895 1094 -895 0 3
rlabel polysilicon 1101 -889 1101 -889 0 1
rlabel polysilicon 1101 -895 1101 -895 0 3
rlabel polysilicon 1108 -889 1108 -889 0 1
rlabel polysilicon 1108 -895 1108 -895 0 3
rlabel polysilicon 1115 -889 1115 -889 0 1
rlabel polysilicon 1115 -895 1115 -895 0 3
rlabel polysilicon 1122 -889 1122 -889 0 1
rlabel polysilicon 1122 -895 1122 -895 0 3
rlabel polysilicon 1129 -889 1129 -889 0 1
rlabel polysilicon 1129 -895 1129 -895 0 3
rlabel polysilicon 1136 -889 1136 -889 0 1
rlabel polysilicon 1136 -895 1136 -895 0 3
rlabel polysilicon 1143 -889 1143 -889 0 1
rlabel polysilicon 1143 -895 1143 -895 0 3
rlabel polysilicon 1150 -889 1150 -889 0 1
rlabel polysilicon 1150 -895 1150 -895 0 3
rlabel polysilicon 1157 -889 1157 -889 0 1
rlabel polysilicon 1157 -895 1157 -895 0 3
rlabel polysilicon 1164 -889 1164 -889 0 1
rlabel polysilicon 1164 -895 1164 -895 0 3
rlabel polysilicon 1171 -889 1171 -889 0 1
rlabel polysilicon 1171 -895 1171 -895 0 3
rlabel polysilicon 1178 -889 1178 -889 0 1
rlabel polysilicon 1178 -895 1178 -895 0 3
rlabel polysilicon 1185 -889 1185 -889 0 1
rlabel polysilicon 1185 -895 1185 -895 0 3
rlabel polysilicon 1192 -889 1192 -889 0 1
rlabel polysilicon 1192 -895 1192 -895 0 3
rlabel polysilicon 1199 -889 1199 -889 0 1
rlabel polysilicon 1199 -895 1199 -895 0 3
rlabel polysilicon 1206 -889 1206 -889 0 1
rlabel polysilicon 1206 -895 1206 -895 0 3
rlabel polysilicon 1213 -889 1213 -889 0 1
rlabel polysilicon 1213 -895 1213 -895 0 3
rlabel polysilicon 1220 -889 1220 -889 0 1
rlabel polysilicon 1220 -895 1220 -895 0 3
rlabel polysilicon 1227 -889 1227 -889 0 1
rlabel polysilicon 1227 -895 1227 -895 0 3
rlabel polysilicon 1234 -889 1234 -889 0 1
rlabel polysilicon 1234 -895 1234 -895 0 3
rlabel polysilicon 1241 -889 1241 -889 0 1
rlabel polysilicon 1241 -895 1241 -895 0 3
rlabel polysilicon 1248 -889 1248 -889 0 1
rlabel polysilicon 1248 -895 1248 -895 0 3
rlabel polysilicon 1255 -889 1255 -889 0 1
rlabel polysilicon 1255 -895 1255 -895 0 3
rlabel polysilicon 1262 -889 1262 -889 0 1
rlabel polysilicon 1262 -895 1262 -895 0 3
rlabel polysilicon 1269 -889 1269 -889 0 1
rlabel polysilicon 1269 -895 1269 -895 0 3
rlabel polysilicon 1276 -889 1276 -889 0 1
rlabel polysilicon 1276 -895 1276 -895 0 3
rlabel polysilicon 1283 -889 1283 -889 0 1
rlabel polysilicon 1283 -895 1283 -895 0 3
rlabel polysilicon 1290 -889 1290 -889 0 1
rlabel polysilicon 1290 -895 1290 -895 0 3
rlabel polysilicon 1297 -889 1297 -889 0 1
rlabel polysilicon 1297 -895 1297 -895 0 3
rlabel polysilicon 1304 -889 1304 -889 0 1
rlabel polysilicon 1304 -895 1304 -895 0 3
rlabel polysilicon 1311 -889 1311 -889 0 1
rlabel polysilicon 1311 -895 1311 -895 0 3
rlabel polysilicon 1318 -889 1318 -889 0 1
rlabel polysilicon 1318 -895 1318 -895 0 3
rlabel polysilicon 1325 -889 1325 -889 0 1
rlabel polysilicon 1325 -895 1325 -895 0 3
rlabel polysilicon 1332 -889 1332 -889 0 1
rlabel polysilicon 1332 -895 1332 -895 0 3
rlabel polysilicon 1339 -889 1339 -889 0 1
rlabel polysilicon 1339 -895 1339 -895 0 3
rlabel polysilicon 1346 -889 1346 -889 0 1
rlabel polysilicon 1346 -895 1346 -895 0 3
rlabel polysilicon 1353 -889 1353 -889 0 1
rlabel polysilicon 1353 -895 1353 -895 0 3
rlabel polysilicon 1360 -889 1360 -889 0 1
rlabel polysilicon 1360 -895 1360 -895 0 3
rlabel polysilicon 1367 -889 1367 -889 0 1
rlabel polysilicon 1367 -895 1367 -895 0 3
rlabel polysilicon 1374 -889 1374 -889 0 1
rlabel polysilicon 1374 -895 1374 -895 0 3
rlabel polysilicon 1381 -889 1381 -889 0 1
rlabel polysilicon 1381 -895 1381 -895 0 3
rlabel polysilicon 1388 -889 1388 -889 0 1
rlabel polysilicon 1388 -895 1388 -895 0 3
rlabel polysilicon 1395 -889 1395 -889 0 1
rlabel polysilicon 1395 -895 1395 -895 0 3
rlabel polysilicon 1402 -889 1402 -889 0 1
rlabel polysilicon 1402 -895 1402 -895 0 3
rlabel polysilicon 1409 -889 1409 -889 0 1
rlabel polysilicon 1409 -895 1409 -895 0 3
rlabel polysilicon 1416 -889 1416 -889 0 1
rlabel polysilicon 1416 -895 1416 -895 0 3
rlabel polysilicon 1423 -889 1423 -889 0 1
rlabel polysilicon 1423 -895 1423 -895 0 3
rlabel polysilicon 1430 -889 1430 -889 0 1
rlabel polysilicon 1430 -895 1430 -895 0 3
rlabel polysilicon 1437 -889 1437 -889 0 1
rlabel polysilicon 1437 -895 1437 -895 0 3
rlabel polysilicon 1444 -889 1444 -889 0 1
rlabel polysilicon 1444 -895 1444 -895 0 3
rlabel polysilicon 1451 -889 1451 -889 0 1
rlabel polysilicon 1451 -895 1451 -895 0 3
rlabel polysilicon 1458 -889 1458 -889 0 1
rlabel polysilicon 1458 -895 1458 -895 0 3
rlabel polysilicon 1465 -889 1465 -889 0 1
rlabel polysilicon 1465 -895 1465 -895 0 3
rlabel polysilicon 1472 -889 1472 -889 0 1
rlabel polysilicon 1472 -895 1472 -895 0 3
rlabel polysilicon 1479 -889 1479 -889 0 1
rlabel polysilicon 1479 -895 1479 -895 0 3
rlabel polysilicon 1486 -889 1486 -889 0 1
rlabel polysilicon 1486 -895 1486 -895 0 3
rlabel polysilicon 1493 -889 1493 -889 0 1
rlabel polysilicon 1493 -895 1493 -895 0 3
rlabel polysilicon 1500 -889 1500 -889 0 1
rlabel polysilicon 1503 -889 1503 -889 0 2
rlabel polysilicon 1500 -895 1500 -895 0 3
rlabel polysilicon 1503 -895 1503 -895 0 4
rlabel polysilicon 1514 -889 1514 -889 0 1
rlabel polysilicon 1514 -895 1514 -895 0 3
rlabel polysilicon 2 -1006 2 -1006 0 1
rlabel polysilicon 2 -1012 2 -1012 0 3
rlabel polysilicon 9 -1006 9 -1006 0 1
rlabel polysilicon 9 -1012 9 -1012 0 3
rlabel polysilicon 16 -1006 16 -1006 0 1
rlabel polysilicon 16 -1012 16 -1012 0 3
rlabel polysilicon 23 -1006 23 -1006 0 1
rlabel polysilicon 23 -1012 23 -1012 0 3
rlabel polysilicon 30 -1006 30 -1006 0 1
rlabel polysilicon 30 -1012 30 -1012 0 3
rlabel polysilicon 37 -1006 37 -1006 0 1
rlabel polysilicon 37 -1012 37 -1012 0 3
rlabel polysilicon 44 -1006 44 -1006 0 1
rlabel polysilicon 44 -1012 44 -1012 0 3
rlabel polysilicon 51 -1006 51 -1006 0 1
rlabel polysilicon 51 -1012 51 -1012 0 3
rlabel polysilicon 58 -1006 58 -1006 0 1
rlabel polysilicon 58 -1012 58 -1012 0 3
rlabel polysilicon 65 -1006 65 -1006 0 1
rlabel polysilicon 65 -1012 65 -1012 0 3
rlabel polysilicon 72 -1006 72 -1006 0 1
rlabel polysilicon 72 -1012 72 -1012 0 3
rlabel polysilicon 79 -1006 79 -1006 0 1
rlabel polysilicon 79 -1012 79 -1012 0 3
rlabel polysilicon 86 -1006 86 -1006 0 1
rlabel polysilicon 86 -1012 86 -1012 0 3
rlabel polysilicon 93 -1006 93 -1006 0 1
rlabel polysilicon 96 -1006 96 -1006 0 2
rlabel polysilicon 93 -1012 93 -1012 0 3
rlabel polysilicon 96 -1012 96 -1012 0 4
rlabel polysilicon 100 -1006 100 -1006 0 1
rlabel polysilicon 100 -1012 100 -1012 0 3
rlabel polysilicon 107 -1006 107 -1006 0 1
rlabel polysilicon 107 -1012 107 -1012 0 3
rlabel polysilicon 114 -1006 114 -1006 0 1
rlabel polysilicon 114 -1012 114 -1012 0 3
rlabel polysilicon 121 -1006 121 -1006 0 1
rlabel polysilicon 121 -1012 121 -1012 0 3
rlabel polysilicon 128 -1006 128 -1006 0 1
rlabel polysilicon 128 -1012 128 -1012 0 3
rlabel polysilicon 135 -1006 135 -1006 0 1
rlabel polysilicon 135 -1012 135 -1012 0 3
rlabel polysilicon 142 -1006 142 -1006 0 1
rlabel polysilicon 145 -1006 145 -1006 0 2
rlabel polysilicon 142 -1012 142 -1012 0 3
rlabel polysilicon 145 -1012 145 -1012 0 4
rlabel polysilicon 149 -1006 149 -1006 0 1
rlabel polysilicon 149 -1012 149 -1012 0 3
rlabel polysilicon 156 -1006 156 -1006 0 1
rlabel polysilicon 156 -1012 156 -1012 0 3
rlabel polysilicon 163 -1006 163 -1006 0 1
rlabel polysilicon 163 -1012 163 -1012 0 3
rlabel polysilicon 170 -1006 170 -1006 0 1
rlabel polysilicon 170 -1012 170 -1012 0 3
rlabel polysilicon 177 -1006 177 -1006 0 1
rlabel polysilicon 177 -1012 177 -1012 0 3
rlabel polysilicon 184 -1006 184 -1006 0 1
rlabel polysilicon 184 -1012 184 -1012 0 3
rlabel polysilicon 191 -1006 191 -1006 0 1
rlabel polysilicon 191 -1012 191 -1012 0 3
rlabel polysilicon 198 -1006 198 -1006 0 1
rlabel polysilicon 198 -1012 198 -1012 0 3
rlabel polysilicon 205 -1006 205 -1006 0 1
rlabel polysilicon 205 -1012 205 -1012 0 3
rlabel polysilicon 212 -1006 212 -1006 0 1
rlabel polysilicon 212 -1012 212 -1012 0 3
rlabel polysilicon 219 -1006 219 -1006 0 1
rlabel polysilicon 219 -1012 219 -1012 0 3
rlabel polysilicon 226 -1006 226 -1006 0 1
rlabel polysilicon 226 -1012 226 -1012 0 3
rlabel polysilicon 233 -1006 233 -1006 0 1
rlabel polysilicon 233 -1012 233 -1012 0 3
rlabel polysilicon 243 -1006 243 -1006 0 2
rlabel polysilicon 240 -1012 240 -1012 0 3
rlabel polysilicon 243 -1012 243 -1012 0 4
rlabel polysilicon 247 -1006 247 -1006 0 1
rlabel polysilicon 247 -1012 247 -1012 0 3
rlabel polysilicon 254 -1006 254 -1006 0 1
rlabel polysilicon 254 -1012 254 -1012 0 3
rlabel polysilicon 261 -1006 261 -1006 0 1
rlabel polysilicon 261 -1012 261 -1012 0 3
rlabel polysilicon 268 -1006 268 -1006 0 1
rlabel polysilicon 268 -1012 268 -1012 0 3
rlabel polysilicon 275 -1006 275 -1006 0 1
rlabel polysilicon 275 -1012 275 -1012 0 3
rlabel polysilicon 282 -1006 282 -1006 0 1
rlabel polysilicon 282 -1012 282 -1012 0 3
rlabel polysilicon 289 -1006 289 -1006 0 1
rlabel polysilicon 289 -1012 289 -1012 0 3
rlabel polysilicon 296 -1006 296 -1006 0 1
rlabel polysilicon 299 -1006 299 -1006 0 2
rlabel polysilicon 296 -1012 296 -1012 0 3
rlabel polysilicon 299 -1012 299 -1012 0 4
rlabel polysilicon 303 -1006 303 -1006 0 1
rlabel polysilicon 303 -1012 303 -1012 0 3
rlabel polysilicon 310 -1006 310 -1006 0 1
rlabel polysilicon 310 -1012 310 -1012 0 3
rlabel polysilicon 317 -1006 317 -1006 0 1
rlabel polysilicon 317 -1012 317 -1012 0 3
rlabel polysilicon 324 -1006 324 -1006 0 1
rlabel polysilicon 324 -1012 324 -1012 0 3
rlabel polysilicon 334 -1006 334 -1006 0 2
rlabel polysilicon 331 -1012 331 -1012 0 3
rlabel polysilicon 334 -1012 334 -1012 0 4
rlabel polysilicon 338 -1006 338 -1006 0 1
rlabel polysilicon 338 -1012 338 -1012 0 3
rlabel polysilicon 345 -1006 345 -1006 0 1
rlabel polysilicon 345 -1012 345 -1012 0 3
rlabel polysilicon 352 -1006 352 -1006 0 1
rlabel polysilicon 352 -1012 352 -1012 0 3
rlabel polysilicon 359 -1006 359 -1006 0 1
rlabel polysilicon 359 -1012 359 -1012 0 3
rlabel polysilicon 366 -1006 366 -1006 0 1
rlabel polysilicon 366 -1012 366 -1012 0 3
rlabel polysilicon 373 -1006 373 -1006 0 1
rlabel polysilicon 376 -1006 376 -1006 0 2
rlabel polysilicon 373 -1012 373 -1012 0 3
rlabel polysilicon 376 -1012 376 -1012 0 4
rlabel polysilicon 380 -1006 380 -1006 0 1
rlabel polysilicon 380 -1012 380 -1012 0 3
rlabel polysilicon 387 -1006 387 -1006 0 1
rlabel polysilicon 387 -1012 387 -1012 0 3
rlabel polysilicon 394 -1006 394 -1006 0 1
rlabel polysilicon 394 -1012 394 -1012 0 3
rlabel polysilicon 401 -1006 401 -1006 0 1
rlabel polysilicon 401 -1012 401 -1012 0 3
rlabel polysilicon 408 -1006 408 -1006 0 1
rlabel polysilicon 408 -1012 408 -1012 0 3
rlabel polysilicon 415 -1006 415 -1006 0 1
rlabel polysilicon 415 -1012 415 -1012 0 3
rlabel polysilicon 422 -1006 422 -1006 0 1
rlabel polysilicon 422 -1012 422 -1012 0 3
rlabel polysilicon 429 -1006 429 -1006 0 1
rlabel polysilicon 429 -1012 429 -1012 0 3
rlabel polysilicon 436 -1006 436 -1006 0 1
rlabel polysilicon 436 -1012 436 -1012 0 3
rlabel polysilicon 443 -1006 443 -1006 0 1
rlabel polysilicon 443 -1012 443 -1012 0 3
rlabel polysilicon 450 -1006 450 -1006 0 1
rlabel polysilicon 450 -1012 450 -1012 0 3
rlabel polysilicon 457 -1006 457 -1006 0 1
rlabel polysilicon 457 -1012 457 -1012 0 3
rlabel polysilicon 464 -1006 464 -1006 0 1
rlabel polysilicon 464 -1012 464 -1012 0 3
rlabel polysilicon 471 -1006 471 -1006 0 1
rlabel polysilicon 471 -1012 471 -1012 0 3
rlabel polysilicon 478 -1006 478 -1006 0 1
rlabel polysilicon 478 -1012 478 -1012 0 3
rlabel polysilicon 481 -1012 481 -1012 0 4
rlabel polysilicon 485 -1006 485 -1006 0 1
rlabel polysilicon 485 -1012 485 -1012 0 3
rlabel polysilicon 492 -1006 492 -1006 0 1
rlabel polysilicon 495 -1006 495 -1006 0 2
rlabel polysilicon 492 -1012 492 -1012 0 3
rlabel polysilicon 495 -1012 495 -1012 0 4
rlabel polysilicon 499 -1006 499 -1006 0 1
rlabel polysilicon 499 -1012 499 -1012 0 3
rlabel polysilicon 506 -1006 506 -1006 0 1
rlabel polysilicon 506 -1012 506 -1012 0 3
rlabel polysilicon 513 -1006 513 -1006 0 1
rlabel polysilicon 513 -1012 513 -1012 0 3
rlabel polysilicon 520 -1006 520 -1006 0 1
rlabel polysilicon 520 -1012 520 -1012 0 3
rlabel polysilicon 527 -1006 527 -1006 0 1
rlabel polysilicon 527 -1012 527 -1012 0 3
rlabel polysilicon 534 -1006 534 -1006 0 1
rlabel polysilicon 537 -1006 537 -1006 0 2
rlabel polysilicon 534 -1012 534 -1012 0 3
rlabel polysilicon 537 -1012 537 -1012 0 4
rlabel polysilicon 541 -1006 541 -1006 0 1
rlabel polysilicon 544 -1006 544 -1006 0 2
rlabel polysilicon 541 -1012 541 -1012 0 3
rlabel polysilicon 544 -1012 544 -1012 0 4
rlabel polysilicon 548 -1006 548 -1006 0 1
rlabel polysilicon 551 -1006 551 -1006 0 2
rlabel polysilicon 548 -1012 548 -1012 0 3
rlabel polysilicon 551 -1012 551 -1012 0 4
rlabel polysilicon 555 -1006 555 -1006 0 1
rlabel polysilicon 555 -1012 555 -1012 0 3
rlabel polysilicon 562 -1006 562 -1006 0 1
rlabel polysilicon 562 -1012 562 -1012 0 3
rlabel polysilicon 569 -1006 569 -1006 0 1
rlabel polysilicon 569 -1012 569 -1012 0 3
rlabel polysilicon 576 -1006 576 -1006 0 1
rlabel polysilicon 576 -1012 576 -1012 0 3
rlabel polysilicon 583 -1006 583 -1006 0 1
rlabel polysilicon 583 -1012 583 -1012 0 3
rlabel polysilicon 590 -1006 590 -1006 0 1
rlabel polysilicon 590 -1012 590 -1012 0 3
rlabel polysilicon 597 -1006 597 -1006 0 1
rlabel polysilicon 600 -1006 600 -1006 0 2
rlabel polysilicon 597 -1012 597 -1012 0 3
rlabel polysilicon 600 -1012 600 -1012 0 4
rlabel polysilicon 604 -1006 604 -1006 0 1
rlabel polysilicon 604 -1012 604 -1012 0 3
rlabel polysilicon 611 -1006 611 -1006 0 1
rlabel polysilicon 611 -1012 611 -1012 0 3
rlabel polysilicon 618 -1006 618 -1006 0 1
rlabel polysilicon 618 -1012 618 -1012 0 3
rlabel polysilicon 625 -1006 625 -1006 0 1
rlabel polysilicon 625 -1012 625 -1012 0 3
rlabel polysilicon 632 -1006 632 -1006 0 1
rlabel polysilicon 632 -1012 632 -1012 0 3
rlabel polysilicon 639 -1006 639 -1006 0 1
rlabel polysilicon 639 -1012 639 -1012 0 3
rlabel polysilicon 646 -1006 646 -1006 0 1
rlabel polysilicon 646 -1012 646 -1012 0 3
rlabel polysilicon 653 -1006 653 -1006 0 1
rlabel polysilicon 653 -1012 653 -1012 0 3
rlabel polysilicon 660 -1006 660 -1006 0 1
rlabel polysilicon 660 -1012 660 -1012 0 3
rlabel polysilicon 667 -1006 667 -1006 0 1
rlabel polysilicon 667 -1012 667 -1012 0 3
rlabel polysilicon 674 -1006 674 -1006 0 1
rlabel polysilicon 677 -1006 677 -1006 0 2
rlabel polysilicon 674 -1012 674 -1012 0 3
rlabel polysilicon 677 -1012 677 -1012 0 4
rlabel polysilicon 681 -1006 681 -1006 0 1
rlabel polysilicon 681 -1012 681 -1012 0 3
rlabel polysilicon 688 -1006 688 -1006 0 1
rlabel polysilicon 691 -1006 691 -1006 0 2
rlabel polysilicon 691 -1012 691 -1012 0 4
rlabel polysilicon 695 -1006 695 -1006 0 1
rlabel polysilicon 695 -1012 695 -1012 0 3
rlabel polysilicon 702 -1006 702 -1006 0 1
rlabel polysilicon 705 -1006 705 -1006 0 2
rlabel polysilicon 702 -1012 702 -1012 0 3
rlabel polysilicon 705 -1012 705 -1012 0 4
rlabel polysilicon 709 -1006 709 -1006 0 1
rlabel polysilicon 709 -1012 709 -1012 0 3
rlabel polysilicon 716 -1006 716 -1006 0 1
rlabel polysilicon 716 -1012 716 -1012 0 3
rlabel polysilicon 723 -1006 723 -1006 0 1
rlabel polysilicon 723 -1012 723 -1012 0 3
rlabel polysilicon 730 -1006 730 -1006 0 1
rlabel polysilicon 730 -1012 730 -1012 0 3
rlabel polysilicon 737 -1006 737 -1006 0 1
rlabel polysilicon 737 -1012 737 -1012 0 3
rlabel polysilicon 744 -1006 744 -1006 0 1
rlabel polysilicon 747 -1006 747 -1006 0 2
rlabel polysilicon 744 -1012 744 -1012 0 3
rlabel polysilicon 747 -1012 747 -1012 0 4
rlabel polysilicon 751 -1006 751 -1006 0 1
rlabel polysilicon 754 -1006 754 -1006 0 2
rlabel polysilicon 751 -1012 751 -1012 0 3
rlabel polysilicon 754 -1012 754 -1012 0 4
rlabel polysilicon 758 -1006 758 -1006 0 1
rlabel polysilicon 761 -1006 761 -1006 0 2
rlabel polysilicon 758 -1012 758 -1012 0 3
rlabel polysilicon 761 -1012 761 -1012 0 4
rlabel polysilicon 765 -1006 765 -1006 0 1
rlabel polysilicon 765 -1012 765 -1012 0 3
rlabel polysilicon 772 -1006 772 -1006 0 1
rlabel polysilicon 772 -1012 772 -1012 0 3
rlabel polysilicon 779 -1006 779 -1006 0 1
rlabel polysilicon 779 -1012 779 -1012 0 3
rlabel polysilicon 786 -1006 786 -1006 0 1
rlabel polysilicon 786 -1012 786 -1012 0 3
rlabel polysilicon 793 -1006 793 -1006 0 1
rlabel polysilicon 793 -1012 793 -1012 0 3
rlabel polysilicon 800 -1006 800 -1006 0 1
rlabel polysilicon 800 -1012 800 -1012 0 3
rlabel polysilicon 807 -1006 807 -1006 0 1
rlabel polysilicon 807 -1012 807 -1012 0 3
rlabel polysilicon 814 -1006 814 -1006 0 1
rlabel polysilicon 814 -1012 814 -1012 0 3
rlabel polysilicon 821 -1006 821 -1006 0 1
rlabel polysilicon 824 -1006 824 -1006 0 2
rlabel polysilicon 821 -1012 821 -1012 0 3
rlabel polysilicon 824 -1012 824 -1012 0 4
rlabel polysilicon 828 -1006 828 -1006 0 1
rlabel polysilicon 831 -1006 831 -1006 0 2
rlabel polysilicon 828 -1012 828 -1012 0 3
rlabel polysilicon 831 -1012 831 -1012 0 4
rlabel polysilicon 835 -1006 835 -1006 0 1
rlabel polysilicon 835 -1012 835 -1012 0 3
rlabel polysilicon 842 -1006 842 -1006 0 1
rlabel polysilicon 842 -1012 842 -1012 0 3
rlabel polysilicon 849 -1006 849 -1006 0 1
rlabel polysilicon 849 -1012 849 -1012 0 3
rlabel polysilicon 856 -1006 856 -1006 0 1
rlabel polysilicon 859 -1006 859 -1006 0 2
rlabel polysilicon 856 -1012 856 -1012 0 3
rlabel polysilicon 859 -1012 859 -1012 0 4
rlabel polysilicon 863 -1006 863 -1006 0 1
rlabel polysilicon 863 -1012 863 -1012 0 3
rlabel polysilicon 870 -1006 870 -1006 0 1
rlabel polysilicon 870 -1012 870 -1012 0 3
rlabel polysilicon 873 -1012 873 -1012 0 4
rlabel polysilicon 877 -1006 877 -1006 0 1
rlabel polysilicon 877 -1012 877 -1012 0 3
rlabel polysilicon 884 -1006 884 -1006 0 1
rlabel polysilicon 884 -1012 884 -1012 0 3
rlabel polysilicon 891 -1006 891 -1006 0 1
rlabel polysilicon 891 -1012 891 -1012 0 3
rlabel polysilicon 898 -1006 898 -1006 0 1
rlabel polysilicon 898 -1012 898 -1012 0 3
rlabel polysilicon 905 -1006 905 -1006 0 1
rlabel polysilicon 908 -1006 908 -1006 0 2
rlabel polysilicon 908 -1012 908 -1012 0 4
rlabel polysilicon 912 -1006 912 -1006 0 1
rlabel polysilicon 912 -1012 912 -1012 0 3
rlabel polysilicon 919 -1006 919 -1006 0 1
rlabel polysilicon 919 -1012 919 -1012 0 3
rlabel polysilicon 926 -1006 926 -1006 0 1
rlabel polysilicon 926 -1012 926 -1012 0 3
rlabel polysilicon 933 -1006 933 -1006 0 1
rlabel polysilicon 933 -1012 933 -1012 0 3
rlabel polysilicon 940 -1006 940 -1006 0 1
rlabel polysilicon 940 -1012 940 -1012 0 3
rlabel polysilicon 947 -1006 947 -1006 0 1
rlabel polysilicon 947 -1012 947 -1012 0 3
rlabel polysilicon 954 -1006 954 -1006 0 1
rlabel polysilicon 954 -1012 954 -1012 0 3
rlabel polysilicon 961 -1006 961 -1006 0 1
rlabel polysilicon 961 -1012 961 -1012 0 3
rlabel polysilicon 968 -1006 968 -1006 0 1
rlabel polysilicon 968 -1012 968 -1012 0 3
rlabel polysilicon 975 -1006 975 -1006 0 1
rlabel polysilicon 975 -1012 975 -1012 0 3
rlabel polysilicon 982 -1012 982 -1012 0 3
rlabel polysilicon 992 -1006 992 -1006 0 2
rlabel polysilicon 989 -1012 989 -1012 0 3
rlabel polysilicon 992 -1012 992 -1012 0 4
rlabel polysilicon 996 -1006 996 -1006 0 1
rlabel polysilicon 996 -1012 996 -1012 0 3
rlabel polysilicon 1003 -1006 1003 -1006 0 1
rlabel polysilicon 1003 -1012 1003 -1012 0 3
rlabel polysilicon 1010 -1006 1010 -1006 0 1
rlabel polysilicon 1010 -1012 1010 -1012 0 3
rlabel polysilicon 1017 -1006 1017 -1006 0 1
rlabel polysilicon 1017 -1012 1017 -1012 0 3
rlabel polysilicon 1024 -1006 1024 -1006 0 1
rlabel polysilicon 1024 -1012 1024 -1012 0 3
rlabel polysilicon 1031 -1006 1031 -1006 0 1
rlabel polysilicon 1031 -1012 1031 -1012 0 3
rlabel polysilicon 1038 -1006 1038 -1006 0 1
rlabel polysilicon 1038 -1012 1038 -1012 0 3
rlabel polysilicon 1045 -1006 1045 -1006 0 1
rlabel polysilicon 1045 -1012 1045 -1012 0 3
rlabel polysilicon 1052 -1006 1052 -1006 0 1
rlabel polysilicon 1052 -1012 1052 -1012 0 3
rlabel polysilicon 1059 -1006 1059 -1006 0 1
rlabel polysilicon 1059 -1012 1059 -1012 0 3
rlabel polysilicon 1066 -1006 1066 -1006 0 1
rlabel polysilicon 1069 -1006 1069 -1006 0 2
rlabel polysilicon 1066 -1012 1066 -1012 0 3
rlabel polysilicon 1073 -1006 1073 -1006 0 1
rlabel polysilicon 1073 -1012 1073 -1012 0 3
rlabel polysilicon 1080 -1006 1080 -1006 0 1
rlabel polysilicon 1080 -1012 1080 -1012 0 3
rlabel polysilicon 1087 -1006 1087 -1006 0 1
rlabel polysilicon 1087 -1012 1087 -1012 0 3
rlabel polysilicon 1094 -1006 1094 -1006 0 1
rlabel polysilicon 1094 -1012 1094 -1012 0 3
rlabel polysilicon 1101 -1006 1101 -1006 0 1
rlabel polysilicon 1101 -1012 1101 -1012 0 3
rlabel polysilicon 1108 -1006 1108 -1006 0 1
rlabel polysilicon 1108 -1012 1108 -1012 0 3
rlabel polysilicon 1115 -1006 1115 -1006 0 1
rlabel polysilicon 1115 -1012 1115 -1012 0 3
rlabel polysilicon 1122 -1006 1122 -1006 0 1
rlabel polysilicon 1122 -1012 1122 -1012 0 3
rlabel polysilicon 1129 -1006 1129 -1006 0 1
rlabel polysilicon 1129 -1012 1129 -1012 0 3
rlabel polysilicon 1136 -1006 1136 -1006 0 1
rlabel polysilicon 1136 -1012 1136 -1012 0 3
rlabel polysilicon 1143 -1006 1143 -1006 0 1
rlabel polysilicon 1143 -1012 1143 -1012 0 3
rlabel polysilicon 1150 -1006 1150 -1006 0 1
rlabel polysilicon 1150 -1012 1150 -1012 0 3
rlabel polysilicon 1157 -1006 1157 -1006 0 1
rlabel polysilicon 1157 -1012 1157 -1012 0 3
rlabel polysilicon 1164 -1006 1164 -1006 0 1
rlabel polysilicon 1164 -1012 1164 -1012 0 3
rlabel polysilicon 1171 -1006 1171 -1006 0 1
rlabel polysilicon 1171 -1012 1171 -1012 0 3
rlabel polysilicon 1178 -1006 1178 -1006 0 1
rlabel polysilicon 1178 -1012 1178 -1012 0 3
rlabel polysilicon 1185 -1006 1185 -1006 0 1
rlabel polysilicon 1185 -1012 1185 -1012 0 3
rlabel polysilicon 1192 -1006 1192 -1006 0 1
rlabel polysilicon 1192 -1012 1192 -1012 0 3
rlabel polysilicon 1199 -1006 1199 -1006 0 1
rlabel polysilicon 1199 -1012 1199 -1012 0 3
rlabel polysilicon 1206 -1006 1206 -1006 0 1
rlabel polysilicon 1206 -1012 1206 -1012 0 3
rlabel polysilicon 1213 -1006 1213 -1006 0 1
rlabel polysilicon 1213 -1012 1213 -1012 0 3
rlabel polysilicon 1220 -1006 1220 -1006 0 1
rlabel polysilicon 1220 -1012 1220 -1012 0 3
rlabel polysilicon 1227 -1006 1227 -1006 0 1
rlabel polysilicon 1227 -1012 1227 -1012 0 3
rlabel polysilicon 1234 -1006 1234 -1006 0 1
rlabel polysilicon 1234 -1012 1234 -1012 0 3
rlabel polysilicon 1241 -1006 1241 -1006 0 1
rlabel polysilicon 1241 -1012 1241 -1012 0 3
rlabel polysilicon 1248 -1006 1248 -1006 0 1
rlabel polysilicon 1248 -1012 1248 -1012 0 3
rlabel polysilicon 1255 -1006 1255 -1006 0 1
rlabel polysilicon 1255 -1012 1255 -1012 0 3
rlabel polysilicon 1262 -1006 1262 -1006 0 1
rlabel polysilicon 1262 -1012 1262 -1012 0 3
rlabel polysilicon 1269 -1006 1269 -1006 0 1
rlabel polysilicon 1269 -1012 1269 -1012 0 3
rlabel polysilicon 1276 -1006 1276 -1006 0 1
rlabel polysilicon 1276 -1012 1276 -1012 0 3
rlabel polysilicon 1283 -1006 1283 -1006 0 1
rlabel polysilicon 1283 -1012 1283 -1012 0 3
rlabel polysilicon 1290 -1006 1290 -1006 0 1
rlabel polysilicon 1290 -1012 1290 -1012 0 3
rlabel polysilicon 1297 -1006 1297 -1006 0 1
rlabel polysilicon 1297 -1012 1297 -1012 0 3
rlabel polysilicon 1304 -1006 1304 -1006 0 1
rlabel polysilicon 1304 -1012 1304 -1012 0 3
rlabel polysilicon 1311 -1006 1311 -1006 0 1
rlabel polysilicon 1311 -1012 1311 -1012 0 3
rlabel polysilicon 1318 -1006 1318 -1006 0 1
rlabel polysilicon 1318 -1012 1318 -1012 0 3
rlabel polysilicon 1325 -1006 1325 -1006 0 1
rlabel polysilicon 1325 -1012 1325 -1012 0 3
rlabel polysilicon 1332 -1006 1332 -1006 0 1
rlabel polysilicon 1332 -1012 1332 -1012 0 3
rlabel polysilicon 1339 -1006 1339 -1006 0 1
rlabel polysilicon 1339 -1012 1339 -1012 0 3
rlabel polysilicon 1346 -1006 1346 -1006 0 1
rlabel polysilicon 1346 -1012 1346 -1012 0 3
rlabel polysilicon 1353 -1006 1353 -1006 0 1
rlabel polysilicon 1353 -1012 1353 -1012 0 3
rlabel polysilicon 1360 -1006 1360 -1006 0 1
rlabel polysilicon 1360 -1012 1360 -1012 0 3
rlabel polysilicon 1367 -1006 1367 -1006 0 1
rlabel polysilicon 1367 -1012 1367 -1012 0 3
rlabel polysilicon 1374 -1006 1374 -1006 0 1
rlabel polysilicon 1374 -1012 1374 -1012 0 3
rlabel polysilicon 1381 -1006 1381 -1006 0 1
rlabel polysilicon 1381 -1012 1381 -1012 0 3
rlabel polysilicon 1388 -1006 1388 -1006 0 1
rlabel polysilicon 1388 -1012 1388 -1012 0 3
rlabel polysilicon 1395 -1006 1395 -1006 0 1
rlabel polysilicon 1395 -1012 1395 -1012 0 3
rlabel polysilicon 1402 -1006 1402 -1006 0 1
rlabel polysilicon 1402 -1012 1402 -1012 0 3
rlabel polysilicon 1409 -1006 1409 -1006 0 1
rlabel polysilicon 1409 -1012 1409 -1012 0 3
rlabel polysilicon 1416 -1006 1416 -1006 0 1
rlabel polysilicon 1416 -1012 1416 -1012 0 3
rlabel polysilicon 1423 -1006 1423 -1006 0 1
rlabel polysilicon 1426 -1006 1426 -1006 0 2
rlabel polysilicon 1423 -1012 1423 -1012 0 3
rlabel polysilicon 1426 -1012 1426 -1012 0 4
rlabel polysilicon 1430 -1006 1430 -1006 0 1
rlabel polysilicon 1430 -1012 1430 -1012 0 3
rlabel polysilicon 1437 -1006 1437 -1006 0 1
rlabel polysilicon 1437 -1012 1437 -1012 0 3
rlabel polysilicon 1444 -1006 1444 -1006 0 1
rlabel polysilicon 1444 -1012 1444 -1012 0 3
rlabel polysilicon 1451 -1006 1451 -1006 0 1
rlabel polysilicon 1451 -1012 1451 -1012 0 3
rlabel polysilicon 1458 -1006 1458 -1006 0 1
rlabel polysilicon 1458 -1012 1458 -1012 0 3
rlabel polysilicon 2 -1153 2 -1153 0 1
rlabel polysilicon 2 -1159 2 -1159 0 3
rlabel polysilicon 9 -1153 9 -1153 0 1
rlabel polysilicon 9 -1159 9 -1159 0 3
rlabel polysilicon 12 -1159 12 -1159 0 4
rlabel polysilicon 16 -1153 16 -1153 0 1
rlabel polysilicon 16 -1159 16 -1159 0 3
rlabel polysilicon 23 -1153 23 -1153 0 1
rlabel polysilicon 23 -1159 23 -1159 0 3
rlabel polysilicon 30 -1153 30 -1153 0 1
rlabel polysilicon 33 -1153 33 -1153 0 2
rlabel polysilicon 33 -1159 33 -1159 0 4
rlabel polysilicon 37 -1153 37 -1153 0 1
rlabel polysilicon 40 -1153 40 -1153 0 2
rlabel polysilicon 37 -1159 37 -1159 0 3
rlabel polysilicon 40 -1159 40 -1159 0 4
rlabel polysilicon 44 -1153 44 -1153 0 1
rlabel polysilicon 44 -1159 44 -1159 0 3
rlabel polysilicon 51 -1153 51 -1153 0 1
rlabel polysilicon 51 -1159 51 -1159 0 3
rlabel polysilicon 58 -1153 58 -1153 0 1
rlabel polysilicon 58 -1159 58 -1159 0 3
rlabel polysilicon 65 -1153 65 -1153 0 1
rlabel polysilicon 65 -1159 65 -1159 0 3
rlabel polysilicon 72 -1153 72 -1153 0 1
rlabel polysilicon 72 -1159 72 -1159 0 3
rlabel polysilicon 79 -1153 79 -1153 0 1
rlabel polysilicon 82 -1153 82 -1153 0 2
rlabel polysilicon 79 -1159 79 -1159 0 3
rlabel polysilicon 82 -1159 82 -1159 0 4
rlabel polysilicon 86 -1153 86 -1153 0 1
rlabel polysilicon 86 -1159 86 -1159 0 3
rlabel polysilicon 93 -1153 93 -1153 0 1
rlabel polysilicon 93 -1159 93 -1159 0 3
rlabel polysilicon 100 -1153 100 -1153 0 1
rlabel polysilicon 100 -1159 100 -1159 0 3
rlabel polysilicon 107 -1153 107 -1153 0 1
rlabel polysilicon 107 -1159 107 -1159 0 3
rlabel polysilicon 114 -1153 114 -1153 0 1
rlabel polysilicon 114 -1159 114 -1159 0 3
rlabel polysilicon 121 -1153 121 -1153 0 1
rlabel polysilicon 121 -1159 121 -1159 0 3
rlabel polysilicon 128 -1153 128 -1153 0 1
rlabel polysilicon 128 -1159 128 -1159 0 3
rlabel polysilicon 135 -1153 135 -1153 0 1
rlabel polysilicon 135 -1159 135 -1159 0 3
rlabel polysilicon 142 -1153 142 -1153 0 1
rlabel polysilicon 142 -1159 142 -1159 0 3
rlabel polysilicon 149 -1153 149 -1153 0 1
rlabel polysilicon 149 -1159 149 -1159 0 3
rlabel polysilicon 156 -1153 156 -1153 0 1
rlabel polysilicon 156 -1159 156 -1159 0 3
rlabel polysilicon 166 -1153 166 -1153 0 2
rlabel polysilicon 163 -1159 163 -1159 0 3
rlabel polysilicon 166 -1159 166 -1159 0 4
rlabel polysilicon 170 -1153 170 -1153 0 1
rlabel polysilicon 170 -1159 170 -1159 0 3
rlabel polysilicon 177 -1153 177 -1153 0 1
rlabel polysilicon 177 -1159 177 -1159 0 3
rlabel polysilicon 184 -1153 184 -1153 0 1
rlabel polysilicon 184 -1159 184 -1159 0 3
rlabel polysilicon 191 -1153 191 -1153 0 1
rlabel polysilicon 191 -1159 191 -1159 0 3
rlabel polysilicon 198 -1153 198 -1153 0 1
rlabel polysilicon 201 -1153 201 -1153 0 2
rlabel polysilicon 198 -1159 198 -1159 0 3
rlabel polysilicon 205 -1153 205 -1153 0 1
rlabel polysilicon 205 -1159 205 -1159 0 3
rlabel polysilicon 212 -1153 212 -1153 0 1
rlabel polysilicon 212 -1159 212 -1159 0 3
rlabel polysilicon 219 -1153 219 -1153 0 1
rlabel polysilicon 219 -1159 219 -1159 0 3
rlabel polysilicon 226 -1153 226 -1153 0 1
rlabel polysilicon 226 -1159 226 -1159 0 3
rlabel polysilicon 233 -1153 233 -1153 0 1
rlabel polysilicon 233 -1159 233 -1159 0 3
rlabel polysilicon 240 -1153 240 -1153 0 1
rlabel polysilicon 240 -1159 240 -1159 0 3
rlabel polysilicon 247 -1153 247 -1153 0 1
rlabel polysilicon 247 -1159 247 -1159 0 3
rlabel polysilicon 254 -1153 254 -1153 0 1
rlabel polysilicon 254 -1159 254 -1159 0 3
rlabel polysilicon 261 -1153 261 -1153 0 1
rlabel polysilicon 261 -1159 261 -1159 0 3
rlabel polysilicon 268 -1153 268 -1153 0 1
rlabel polysilicon 268 -1159 268 -1159 0 3
rlabel polysilicon 275 -1153 275 -1153 0 1
rlabel polysilicon 275 -1159 275 -1159 0 3
rlabel polysilicon 282 -1153 282 -1153 0 1
rlabel polysilicon 282 -1159 282 -1159 0 3
rlabel polysilicon 289 -1153 289 -1153 0 1
rlabel polysilicon 289 -1159 289 -1159 0 3
rlabel polysilicon 296 -1153 296 -1153 0 1
rlabel polysilicon 296 -1159 296 -1159 0 3
rlabel polysilicon 303 -1153 303 -1153 0 1
rlabel polysilicon 303 -1159 303 -1159 0 3
rlabel polysilicon 310 -1153 310 -1153 0 1
rlabel polysilicon 310 -1159 310 -1159 0 3
rlabel polysilicon 317 -1153 317 -1153 0 1
rlabel polysilicon 317 -1159 317 -1159 0 3
rlabel polysilicon 324 -1153 324 -1153 0 1
rlabel polysilicon 324 -1159 324 -1159 0 3
rlabel polysilicon 331 -1153 331 -1153 0 1
rlabel polysilicon 331 -1159 331 -1159 0 3
rlabel polysilicon 338 -1153 338 -1153 0 1
rlabel polysilicon 338 -1159 338 -1159 0 3
rlabel polysilicon 345 -1153 345 -1153 0 1
rlabel polysilicon 345 -1159 345 -1159 0 3
rlabel polysilicon 352 -1153 352 -1153 0 1
rlabel polysilicon 355 -1153 355 -1153 0 2
rlabel polysilicon 352 -1159 352 -1159 0 3
rlabel polysilicon 355 -1159 355 -1159 0 4
rlabel polysilicon 359 -1153 359 -1153 0 1
rlabel polysilicon 359 -1159 359 -1159 0 3
rlabel polysilicon 366 -1153 366 -1153 0 1
rlabel polysilicon 366 -1159 366 -1159 0 3
rlabel polysilicon 373 -1153 373 -1153 0 1
rlabel polysilicon 373 -1159 373 -1159 0 3
rlabel polysilicon 380 -1153 380 -1153 0 1
rlabel polysilicon 380 -1159 380 -1159 0 3
rlabel polysilicon 387 -1153 387 -1153 0 1
rlabel polysilicon 390 -1153 390 -1153 0 2
rlabel polysilicon 387 -1159 387 -1159 0 3
rlabel polysilicon 390 -1159 390 -1159 0 4
rlabel polysilicon 394 -1153 394 -1153 0 1
rlabel polysilicon 394 -1159 394 -1159 0 3
rlabel polysilicon 401 -1153 401 -1153 0 1
rlabel polysilicon 401 -1159 401 -1159 0 3
rlabel polysilicon 408 -1153 408 -1153 0 1
rlabel polysilicon 408 -1159 408 -1159 0 3
rlabel polysilicon 415 -1153 415 -1153 0 1
rlabel polysilicon 415 -1159 415 -1159 0 3
rlabel polysilicon 422 -1153 422 -1153 0 1
rlabel polysilicon 422 -1159 422 -1159 0 3
rlabel polysilicon 432 -1153 432 -1153 0 2
rlabel polysilicon 429 -1159 429 -1159 0 3
rlabel polysilicon 436 -1153 436 -1153 0 1
rlabel polysilicon 436 -1159 436 -1159 0 3
rlabel polysilicon 443 -1153 443 -1153 0 1
rlabel polysilicon 446 -1153 446 -1153 0 2
rlabel polysilicon 443 -1159 443 -1159 0 3
rlabel polysilicon 446 -1159 446 -1159 0 4
rlabel polysilicon 450 -1153 450 -1153 0 1
rlabel polysilicon 450 -1159 450 -1159 0 3
rlabel polysilicon 457 -1153 457 -1153 0 1
rlabel polysilicon 460 -1153 460 -1153 0 2
rlabel polysilicon 457 -1159 457 -1159 0 3
rlabel polysilicon 460 -1159 460 -1159 0 4
rlabel polysilicon 464 -1153 464 -1153 0 1
rlabel polysilicon 464 -1159 464 -1159 0 3
rlabel polysilicon 471 -1153 471 -1153 0 1
rlabel polysilicon 471 -1159 471 -1159 0 3
rlabel polysilicon 478 -1153 478 -1153 0 1
rlabel polysilicon 478 -1159 478 -1159 0 3
rlabel polysilicon 485 -1153 485 -1153 0 1
rlabel polysilicon 485 -1159 485 -1159 0 3
rlabel polysilicon 492 -1153 492 -1153 0 1
rlabel polysilicon 492 -1159 492 -1159 0 3
rlabel polysilicon 499 -1153 499 -1153 0 1
rlabel polysilicon 499 -1159 499 -1159 0 3
rlabel polysilicon 506 -1153 506 -1153 0 1
rlabel polysilicon 506 -1159 506 -1159 0 3
rlabel polysilicon 513 -1153 513 -1153 0 1
rlabel polysilicon 513 -1159 513 -1159 0 3
rlabel polysilicon 520 -1153 520 -1153 0 1
rlabel polysilicon 520 -1159 520 -1159 0 3
rlabel polysilicon 527 -1153 527 -1153 0 1
rlabel polysilicon 527 -1159 527 -1159 0 3
rlabel polysilicon 534 -1153 534 -1153 0 1
rlabel polysilicon 534 -1159 534 -1159 0 3
rlabel polysilicon 541 -1153 541 -1153 0 1
rlabel polysilicon 541 -1159 541 -1159 0 3
rlabel polysilicon 548 -1153 548 -1153 0 1
rlabel polysilicon 548 -1159 548 -1159 0 3
rlabel polysilicon 555 -1153 555 -1153 0 1
rlabel polysilicon 555 -1159 555 -1159 0 3
rlabel polysilicon 562 -1153 562 -1153 0 1
rlabel polysilicon 562 -1159 562 -1159 0 3
rlabel polysilicon 569 -1153 569 -1153 0 1
rlabel polysilicon 569 -1159 569 -1159 0 3
rlabel polysilicon 576 -1153 576 -1153 0 1
rlabel polysilicon 576 -1159 576 -1159 0 3
rlabel polysilicon 583 -1153 583 -1153 0 1
rlabel polysilicon 583 -1159 583 -1159 0 3
rlabel polysilicon 590 -1153 590 -1153 0 1
rlabel polysilicon 593 -1153 593 -1153 0 2
rlabel polysilicon 590 -1159 590 -1159 0 3
rlabel polysilicon 593 -1159 593 -1159 0 4
rlabel polysilicon 597 -1153 597 -1153 0 1
rlabel polysilicon 597 -1159 597 -1159 0 3
rlabel polysilicon 604 -1153 604 -1153 0 1
rlabel polysilicon 607 -1153 607 -1153 0 2
rlabel polysilicon 604 -1159 604 -1159 0 3
rlabel polysilicon 611 -1153 611 -1153 0 1
rlabel polysilicon 611 -1159 611 -1159 0 3
rlabel polysilicon 618 -1153 618 -1153 0 1
rlabel polysilicon 618 -1159 618 -1159 0 3
rlabel polysilicon 625 -1153 625 -1153 0 1
rlabel polysilicon 628 -1153 628 -1153 0 2
rlabel polysilicon 625 -1159 625 -1159 0 3
rlabel polysilicon 628 -1159 628 -1159 0 4
rlabel polysilicon 632 -1153 632 -1153 0 1
rlabel polysilicon 632 -1159 632 -1159 0 3
rlabel polysilicon 639 -1153 639 -1153 0 1
rlabel polysilicon 639 -1159 639 -1159 0 3
rlabel polysilicon 646 -1153 646 -1153 0 1
rlabel polysilicon 646 -1159 646 -1159 0 3
rlabel polysilicon 653 -1153 653 -1153 0 1
rlabel polysilicon 653 -1159 653 -1159 0 3
rlabel polysilicon 660 -1153 660 -1153 0 1
rlabel polysilicon 663 -1153 663 -1153 0 2
rlabel polysilicon 660 -1159 660 -1159 0 3
rlabel polysilicon 663 -1159 663 -1159 0 4
rlabel polysilicon 667 -1153 667 -1153 0 1
rlabel polysilicon 670 -1153 670 -1153 0 2
rlabel polysilicon 667 -1159 667 -1159 0 3
rlabel polysilicon 670 -1159 670 -1159 0 4
rlabel polysilicon 674 -1153 674 -1153 0 1
rlabel polysilicon 674 -1159 674 -1159 0 3
rlabel polysilicon 681 -1153 681 -1153 0 1
rlabel polysilicon 681 -1159 681 -1159 0 3
rlabel polysilicon 688 -1153 688 -1153 0 1
rlabel polysilicon 688 -1159 688 -1159 0 3
rlabel polysilicon 695 -1153 695 -1153 0 1
rlabel polysilicon 695 -1159 695 -1159 0 3
rlabel polysilicon 702 -1153 702 -1153 0 1
rlabel polysilicon 702 -1159 702 -1159 0 3
rlabel polysilicon 709 -1153 709 -1153 0 1
rlabel polysilicon 709 -1159 709 -1159 0 3
rlabel polysilicon 716 -1153 716 -1153 0 1
rlabel polysilicon 719 -1153 719 -1153 0 2
rlabel polysilicon 716 -1159 716 -1159 0 3
rlabel polysilicon 719 -1159 719 -1159 0 4
rlabel polysilicon 723 -1153 723 -1153 0 1
rlabel polysilicon 723 -1159 723 -1159 0 3
rlabel polysilicon 730 -1153 730 -1153 0 1
rlabel polysilicon 733 -1153 733 -1153 0 2
rlabel polysilicon 730 -1159 730 -1159 0 3
rlabel polysilicon 733 -1159 733 -1159 0 4
rlabel polysilicon 737 -1153 737 -1153 0 1
rlabel polysilicon 737 -1159 737 -1159 0 3
rlabel polysilicon 744 -1153 744 -1153 0 1
rlabel polysilicon 744 -1159 744 -1159 0 3
rlabel polysilicon 751 -1153 751 -1153 0 1
rlabel polysilicon 754 -1153 754 -1153 0 2
rlabel polysilicon 751 -1159 751 -1159 0 3
rlabel polysilicon 754 -1159 754 -1159 0 4
rlabel polysilicon 758 -1153 758 -1153 0 1
rlabel polysilicon 758 -1159 758 -1159 0 3
rlabel polysilicon 765 -1153 765 -1153 0 1
rlabel polysilicon 765 -1159 765 -1159 0 3
rlabel polysilicon 772 -1153 772 -1153 0 1
rlabel polysilicon 772 -1159 772 -1159 0 3
rlabel polysilicon 779 -1153 779 -1153 0 1
rlabel polysilicon 779 -1159 779 -1159 0 3
rlabel polysilicon 786 -1153 786 -1153 0 1
rlabel polysilicon 786 -1159 786 -1159 0 3
rlabel polysilicon 793 -1153 793 -1153 0 1
rlabel polysilicon 796 -1153 796 -1153 0 2
rlabel polysilicon 793 -1159 793 -1159 0 3
rlabel polysilicon 796 -1159 796 -1159 0 4
rlabel polysilicon 800 -1153 800 -1153 0 1
rlabel polysilicon 800 -1159 800 -1159 0 3
rlabel polysilicon 807 -1153 807 -1153 0 1
rlabel polysilicon 807 -1159 807 -1159 0 3
rlabel polysilicon 814 -1153 814 -1153 0 1
rlabel polysilicon 814 -1159 814 -1159 0 3
rlabel polysilicon 821 -1153 821 -1153 0 1
rlabel polysilicon 821 -1159 821 -1159 0 3
rlabel polysilicon 828 -1153 828 -1153 0 1
rlabel polysilicon 831 -1153 831 -1153 0 2
rlabel polysilicon 828 -1159 828 -1159 0 3
rlabel polysilicon 831 -1159 831 -1159 0 4
rlabel polysilicon 835 -1153 835 -1153 0 1
rlabel polysilicon 835 -1159 835 -1159 0 3
rlabel polysilicon 842 -1153 842 -1153 0 1
rlabel polysilicon 842 -1159 842 -1159 0 3
rlabel polysilicon 849 -1153 849 -1153 0 1
rlabel polysilicon 849 -1159 849 -1159 0 3
rlabel polysilicon 856 -1153 856 -1153 0 1
rlabel polysilicon 859 -1153 859 -1153 0 2
rlabel polysilicon 856 -1159 856 -1159 0 3
rlabel polysilicon 859 -1159 859 -1159 0 4
rlabel polysilicon 863 -1153 863 -1153 0 1
rlabel polysilicon 863 -1159 863 -1159 0 3
rlabel polysilicon 870 -1153 870 -1153 0 1
rlabel polysilicon 870 -1159 870 -1159 0 3
rlabel polysilicon 877 -1153 877 -1153 0 1
rlabel polysilicon 877 -1159 877 -1159 0 3
rlabel polysilicon 884 -1153 884 -1153 0 1
rlabel polysilicon 884 -1159 884 -1159 0 3
rlabel polysilicon 894 -1153 894 -1153 0 2
rlabel polysilicon 891 -1159 891 -1159 0 3
rlabel polysilicon 894 -1159 894 -1159 0 4
rlabel polysilicon 898 -1153 898 -1153 0 1
rlabel polysilicon 898 -1159 898 -1159 0 3
rlabel polysilicon 905 -1153 905 -1153 0 1
rlabel polysilicon 905 -1159 905 -1159 0 3
rlabel polysilicon 912 -1153 912 -1153 0 1
rlabel polysilicon 912 -1159 912 -1159 0 3
rlabel polysilicon 919 -1153 919 -1153 0 1
rlabel polysilicon 919 -1159 919 -1159 0 3
rlabel polysilicon 926 -1153 926 -1153 0 1
rlabel polysilicon 926 -1159 926 -1159 0 3
rlabel polysilicon 933 -1153 933 -1153 0 1
rlabel polysilicon 936 -1153 936 -1153 0 2
rlabel polysilicon 933 -1159 933 -1159 0 3
rlabel polysilicon 936 -1159 936 -1159 0 4
rlabel polysilicon 940 -1153 940 -1153 0 1
rlabel polysilicon 940 -1159 940 -1159 0 3
rlabel polysilicon 947 -1153 947 -1153 0 1
rlabel polysilicon 947 -1159 947 -1159 0 3
rlabel polysilicon 954 -1153 954 -1153 0 1
rlabel polysilicon 957 -1153 957 -1153 0 2
rlabel polysilicon 954 -1159 954 -1159 0 3
rlabel polysilicon 957 -1159 957 -1159 0 4
rlabel polysilicon 961 -1153 961 -1153 0 1
rlabel polysilicon 961 -1159 961 -1159 0 3
rlabel polysilicon 968 -1153 968 -1153 0 1
rlabel polysilicon 968 -1159 968 -1159 0 3
rlabel polysilicon 975 -1153 975 -1153 0 1
rlabel polysilicon 975 -1159 975 -1159 0 3
rlabel polysilicon 982 -1153 982 -1153 0 1
rlabel polysilicon 982 -1159 982 -1159 0 3
rlabel polysilicon 989 -1153 989 -1153 0 1
rlabel polysilicon 989 -1159 989 -1159 0 3
rlabel polysilicon 996 -1153 996 -1153 0 1
rlabel polysilicon 996 -1159 996 -1159 0 3
rlabel polysilicon 1003 -1153 1003 -1153 0 1
rlabel polysilicon 1003 -1159 1003 -1159 0 3
rlabel polysilicon 1010 -1153 1010 -1153 0 1
rlabel polysilicon 1010 -1159 1010 -1159 0 3
rlabel polysilicon 1017 -1153 1017 -1153 0 1
rlabel polysilicon 1017 -1159 1017 -1159 0 3
rlabel polysilicon 1024 -1153 1024 -1153 0 1
rlabel polysilicon 1024 -1159 1024 -1159 0 3
rlabel polysilicon 1031 -1153 1031 -1153 0 1
rlabel polysilicon 1038 -1153 1038 -1153 0 1
rlabel polysilicon 1038 -1159 1038 -1159 0 3
rlabel polysilicon 1045 -1153 1045 -1153 0 1
rlabel polysilicon 1045 -1159 1045 -1159 0 3
rlabel polysilicon 1052 -1153 1052 -1153 0 1
rlabel polysilicon 1052 -1159 1052 -1159 0 3
rlabel polysilicon 1059 -1153 1059 -1153 0 1
rlabel polysilicon 1059 -1159 1059 -1159 0 3
rlabel polysilicon 1066 -1153 1066 -1153 0 1
rlabel polysilicon 1066 -1159 1066 -1159 0 3
rlabel polysilicon 1073 -1153 1073 -1153 0 1
rlabel polysilicon 1073 -1159 1073 -1159 0 3
rlabel polysilicon 1080 -1153 1080 -1153 0 1
rlabel polysilicon 1080 -1159 1080 -1159 0 3
rlabel polysilicon 1087 -1153 1087 -1153 0 1
rlabel polysilicon 1087 -1159 1087 -1159 0 3
rlabel polysilicon 1094 -1153 1094 -1153 0 1
rlabel polysilicon 1094 -1159 1094 -1159 0 3
rlabel polysilicon 1101 -1153 1101 -1153 0 1
rlabel polysilicon 1101 -1159 1101 -1159 0 3
rlabel polysilicon 1108 -1153 1108 -1153 0 1
rlabel polysilicon 1108 -1159 1108 -1159 0 3
rlabel polysilicon 1115 -1153 1115 -1153 0 1
rlabel polysilicon 1115 -1159 1115 -1159 0 3
rlabel polysilicon 1122 -1153 1122 -1153 0 1
rlabel polysilicon 1122 -1159 1122 -1159 0 3
rlabel polysilicon 1129 -1153 1129 -1153 0 1
rlabel polysilicon 1129 -1159 1129 -1159 0 3
rlabel polysilicon 1136 -1153 1136 -1153 0 1
rlabel polysilicon 1136 -1159 1136 -1159 0 3
rlabel polysilicon 1143 -1153 1143 -1153 0 1
rlabel polysilicon 1143 -1159 1143 -1159 0 3
rlabel polysilicon 1150 -1153 1150 -1153 0 1
rlabel polysilicon 1150 -1159 1150 -1159 0 3
rlabel polysilicon 1157 -1153 1157 -1153 0 1
rlabel polysilicon 1157 -1159 1157 -1159 0 3
rlabel polysilicon 1164 -1153 1164 -1153 0 1
rlabel polysilicon 1164 -1159 1164 -1159 0 3
rlabel polysilicon 1171 -1153 1171 -1153 0 1
rlabel polysilicon 1171 -1159 1171 -1159 0 3
rlabel polysilicon 1178 -1153 1178 -1153 0 1
rlabel polysilicon 1178 -1159 1178 -1159 0 3
rlabel polysilicon 1185 -1153 1185 -1153 0 1
rlabel polysilicon 1185 -1159 1185 -1159 0 3
rlabel polysilicon 1192 -1153 1192 -1153 0 1
rlabel polysilicon 1192 -1159 1192 -1159 0 3
rlabel polysilicon 1199 -1153 1199 -1153 0 1
rlabel polysilicon 1199 -1159 1199 -1159 0 3
rlabel polysilicon 1206 -1153 1206 -1153 0 1
rlabel polysilicon 1206 -1159 1206 -1159 0 3
rlabel polysilicon 1213 -1153 1213 -1153 0 1
rlabel polysilicon 1213 -1159 1213 -1159 0 3
rlabel polysilicon 1220 -1153 1220 -1153 0 1
rlabel polysilicon 1220 -1159 1220 -1159 0 3
rlabel polysilicon 1227 -1153 1227 -1153 0 1
rlabel polysilicon 1227 -1159 1227 -1159 0 3
rlabel polysilicon 1234 -1153 1234 -1153 0 1
rlabel polysilicon 1234 -1159 1234 -1159 0 3
rlabel polysilicon 1241 -1153 1241 -1153 0 1
rlabel polysilicon 1241 -1159 1241 -1159 0 3
rlabel polysilicon 1248 -1153 1248 -1153 0 1
rlabel polysilicon 1248 -1159 1248 -1159 0 3
rlabel polysilicon 1251 -1159 1251 -1159 0 4
rlabel polysilicon 1255 -1153 1255 -1153 0 1
rlabel polysilicon 1255 -1159 1255 -1159 0 3
rlabel polysilicon 1262 -1153 1262 -1153 0 1
rlabel polysilicon 1262 -1159 1262 -1159 0 3
rlabel polysilicon 1269 -1153 1269 -1153 0 1
rlabel polysilicon 1269 -1159 1269 -1159 0 3
rlabel polysilicon 1276 -1153 1276 -1153 0 1
rlabel polysilicon 1276 -1159 1276 -1159 0 3
rlabel polysilicon 1283 -1153 1283 -1153 0 1
rlabel polysilicon 1283 -1159 1283 -1159 0 3
rlabel polysilicon 1290 -1153 1290 -1153 0 1
rlabel polysilicon 1290 -1159 1290 -1159 0 3
rlabel polysilicon 1297 -1153 1297 -1153 0 1
rlabel polysilicon 1297 -1159 1297 -1159 0 3
rlabel polysilicon 1304 -1153 1304 -1153 0 1
rlabel polysilicon 1304 -1159 1304 -1159 0 3
rlabel polysilicon 1311 -1153 1311 -1153 0 1
rlabel polysilicon 1311 -1159 1311 -1159 0 3
rlabel polysilicon 1318 -1153 1318 -1153 0 1
rlabel polysilicon 1318 -1159 1318 -1159 0 3
rlabel polysilicon 1325 -1153 1325 -1153 0 1
rlabel polysilicon 1325 -1159 1325 -1159 0 3
rlabel polysilicon 1332 -1153 1332 -1153 0 1
rlabel polysilicon 1332 -1159 1332 -1159 0 3
rlabel polysilicon 1339 -1153 1339 -1153 0 1
rlabel polysilicon 1339 -1159 1339 -1159 0 3
rlabel polysilicon 1346 -1153 1346 -1153 0 1
rlabel polysilicon 1346 -1159 1346 -1159 0 3
rlabel polysilicon 1353 -1153 1353 -1153 0 1
rlabel polysilicon 1353 -1159 1353 -1159 0 3
rlabel polysilicon 1360 -1153 1360 -1153 0 1
rlabel polysilicon 1360 -1159 1360 -1159 0 3
rlabel polysilicon 1367 -1153 1367 -1153 0 1
rlabel polysilicon 1367 -1159 1367 -1159 0 3
rlabel polysilicon 1374 -1153 1374 -1153 0 1
rlabel polysilicon 1374 -1159 1374 -1159 0 3
rlabel polysilicon 1381 -1153 1381 -1153 0 1
rlabel polysilicon 1381 -1159 1381 -1159 0 3
rlabel polysilicon 1388 -1153 1388 -1153 0 1
rlabel polysilicon 1388 -1159 1388 -1159 0 3
rlabel polysilicon 1395 -1153 1395 -1153 0 1
rlabel polysilicon 1395 -1159 1395 -1159 0 3
rlabel polysilicon 1402 -1153 1402 -1153 0 1
rlabel polysilicon 1402 -1159 1402 -1159 0 3
rlabel polysilicon 1409 -1153 1409 -1153 0 1
rlabel polysilicon 1409 -1159 1409 -1159 0 3
rlabel polysilicon 1416 -1153 1416 -1153 0 1
rlabel polysilicon 1416 -1159 1416 -1159 0 3
rlabel polysilicon 1423 -1153 1423 -1153 0 1
rlabel polysilicon 1423 -1159 1423 -1159 0 3
rlabel polysilicon 1430 -1153 1430 -1153 0 1
rlabel polysilicon 1430 -1159 1430 -1159 0 3
rlabel polysilicon 1437 -1153 1437 -1153 0 1
rlabel polysilicon 1437 -1159 1437 -1159 0 3
rlabel polysilicon 1444 -1153 1444 -1153 0 1
rlabel polysilicon 1444 -1159 1444 -1159 0 3
rlabel polysilicon 1451 -1153 1451 -1153 0 1
rlabel polysilicon 1451 -1159 1451 -1159 0 3
rlabel polysilicon 1458 -1153 1458 -1153 0 1
rlabel polysilicon 1458 -1159 1458 -1159 0 3
rlabel polysilicon 1465 -1153 1465 -1153 0 1
rlabel polysilicon 1465 -1159 1465 -1159 0 3
rlabel polysilicon 1472 -1153 1472 -1153 0 1
rlabel polysilicon 1472 -1159 1472 -1159 0 3
rlabel polysilicon 1479 -1153 1479 -1153 0 1
rlabel polysilicon 1479 -1159 1479 -1159 0 3
rlabel polysilicon 1486 -1153 1486 -1153 0 1
rlabel polysilicon 1486 -1159 1486 -1159 0 3
rlabel polysilicon 1493 -1153 1493 -1153 0 1
rlabel polysilicon 1493 -1159 1493 -1159 0 3
rlabel polysilicon 1500 -1153 1500 -1153 0 1
rlabel polysilicon 1500 -1159 1500 -1159 0 3
rlabel polysilicon 1507 -1153 1507 -1153 0 1
rlabel polysilicon 1507 -1159 1507 -1159 0 3
rlabel polysilicon 1514 -1153 1514 -1153 0 1
rlabel polysilicon 1514 -1159 1514 -1159 0 3
rlabel polysilicon 1521 -1153 1521 -1153 0 1
rlabel polysilicon 1521 -1159 1521 -1159 0 3
rlabel polysilicon 1528 -1153 1528 -1153 0 1
rlabel polysilicon 1528 -1159 1528 -1159 0 3
rlabel polysilicon 1535 -1153 1535 -1153 0 1
rlabel polysilicon 1535 -1159 1535 -1159 0 3
rlabel polysilicon 1542 -1153 1542 -1153 0 1
rlabel polysilicon 1542 -1159 1542 -1159 0 3
rlabel polysilicon 1549 -1153 1549 -1153 0 1
rlabel polysilicon 1549 -1159 1549 -1159 0 3
rlabel polysilicon 1556 -1153 1556 -1153 0 1
rlabel polysilicon 1556 -1159 1556 -1159 0 3
rlabel polysilicon 1563 -1153 1563 -1153 0 1
rlabel polysilicon 1563 -1159 1563 -1159 0 3
rlabel polysilicon 1570 -1153 1570 -1153 0 1
rlabel polysilicon 1570 -1159 1570 -1159 0 3
rlabel polysilicon 1577 -1153 1577 -1153 0 1
rlabel polysilicon 1577 -1159 1577 -1159 0 3
rlabel polysilicon 1584 -1153 1584 -1153 0 1
rlabel polysilicon 1584 -1159 1584 -1159 0 3
rlabel polysilicon 1591 -1153 1591 -1153 0 1
rlabel polysilicon 1591 -1159 1591 -1159 0 3
rlabel polysilicon 1598 -1153 1598 -1153 0 1
rlabel polysilicon 1598 -1159 1598 -1159 0 3
rlabel polysilicon 2 -1278 2 -1278 0 1
rlabel polysilicon 2 -1284 2 -1284 0 3
rlabel polysilicon 9 -1278 9 -1278 0 1
rlabel polysilicon 9 -1284 9 -1284 0 3
rlabel polysilicon 16 -1278 16 -1278 0 1
rlabel polysilicon 16 -1284 16 -1284 0 3
rlabel polysilicon 23 -1278 23 -1278 0 1
rlabel polysilicon 23 -1284 23 -1284 0 3
rlabel polysilicon 30 -1278 30 -1278 0 1
rlabel polysilicon 30 -1284 30 -1284 0 3
rlabel polysilicon 37 -1278 37 -1278 0 1
rlabel polysilicon 37 -1284 37 -1284 0 3
rlabel polysilicon 44 -1278 44 -1278 0 1
rlabel polysilicon 44 -1284 44 -1284 0 3
rlabel polysilicon 51 -1278 51 -1278 0 1
rlabel polysilicon 51 -1284 51 -1284 0 3
rlabel polysilicon 58 -1278 58 -1278 0 1
rlabel polysilicon 61 -1278 61 -1278 0 2
rlabel polysilicon 58 -1284 58 -1284 0 3
rlabel polysilicon 61 -1284 61 -1284 0 4
rlabel polysilicon 65 -1278 65 -1278 0 1
rlabel polysilicon 65 -1284 65 -1284 0 3
rlabel polysilicon 72 -1278 72 -1278 0 1
rlabel polysilicon 72 -1284 72 -1284 0 3
rlabel polysilicon 79 -1278 79 -1278 0 1
rlabel polysilicon 79 -1284 79 -1284 0 3
rlabel polysilicon 86 -1278 86 -1278 0 1
rlabel polysilicon 86 -1284 86 -1284 0 3
rlabel polysilicon 93 -1278 93 -1278 0 1
rlabel polysilicon 93 -1284 93 -1284 0 3
rlabel polysilicon 100 -1278 100 -1278 0 1
rlabel polysilicon 103 -1278 103 -1278 0 2
rlabel polysilicon 100 -1284 100 -1284 0 3
rlabel polysilicon 103 -1284 103 -1284 0 4
rlabel polysilicon 107 -1278 107 -1278 0 1
rlabel polysilicon 107 -1284 107 -1284 0 3
rlabel polysilicon 114 -1278 114 -1278 0 1
rlabel polysilicon 114 -1284 114 -1284 0 3
rlabel polysilicon 121 -1278 121 -1278 0 1
rlabel polysilicon 121 -1284 121 -1284 0 3
rlabel polysilicon 128 -1278 128 -1278 0 1
rlabel polysilicon 131 -1278 131 -1278 0 2
rlabel polysilicon 128 -1284 128 -1284 0 3
rlabel polysilicon 131 -1284 131 -1284 0 4
rlabel polysilicon 135 -1278 135 -1278 0 1
rlabel polysilicon 135 -1284 135 -1284 0 3
rlabel polysilicon 142 -1278 142 -1278 0 1
rlabel polysilicon 142 -1284 142 -1284 0 3
rlabel polysilicon 149 -1278 149 -1278 0 1
rlabel polysilicon 149 -1284 149 -1284 0 3
rlabel polysilicon 156 -1278 156 -1278 0 1
rlabel polysilicon 156 -1284 156 -1284 0 3
rlabel polysilicon 163 -1278 163 -1278 0 1
rlabel polysilicon 163 -1284 163 -1284 0 3
rlabel polysilicon 170 -1278 170 -1278 0 1
rlabel polysilicon 173 -1278 173 -1278 0 2
rlabel polysilicon 170 -1284 170 -1284 0 3
rlabel polysilicon 177 -1278 177 -1278 0 1
rlabel polysilicon 177 -1284 177 -1284 0 3
rlabel polysilicon 184 -1278 184 -1278 0 1
rlabel polysilicon 184 -1284 184 -1284 0 3
rlabel polysilicon 191 -1278 191 -1278 0 1
rlabel polysilicon 191 -1284 191 -1284 0 3
rlabel polysilicon 198 -1278 198 -1278 0 1
rlabel polysilicon 198 -1284 198 -1284 0 3
rlabel polysilicon 205 -1278 205 -1278 0 1
rlabel polysilicon 205 -1284 205 -1284 0 3
rlabel polysilicon 212 -1278 212 -1278 0 1
rlabel polysilicon 212 -1284 212 -1284 0 3
rlabel polysilicon 219 -1278 219 -1278 0 1
rlabel polysilicon 219 -1284 219 -1284 0 3
rlabel polysilicon 226 -1278 226 -1278 0 1
rlabel polysilicon 226 -1284 226 -1284 0 3
rlabel polysilicon 233 -1278 233 -1278 0 1
rlabel polysilicon 233 -1284 233 -1284 0 3
rlabel polysilicon 240 -1278 240 -1278 0 1
rlabel polysilicon 240 -1284 240 -1284 0 3
rlabel polysilicon 247 -1278 247 -1278 0 1
rlabel polysilicon 247 -1284 247 -1284 0 3
rlabel polysilicon 254 -1278 254 -1278 0 1
rlabel polysilicon 254 -1284 254 -1284 0 3
rlabel polysilicon 261 -1278 261 -1278 0 1
rlabel polysilicon 261 -1284 261 -1284 0 3
rlabel polysilicon 268 -1278 268 -1278 0 1
rlabel polysilicon 268 -1284 268 -1284 0 3
rlabel polysilicon 275 -1278 275 -1278 0 1
rlabel polysilicon 275 -1284 275 -1284 0 3
rlabel polysilicon 282 -1278 282 -1278 0 1
rlabel polysilicon 282 -1284 282 -1284 0 3
rlabel polysilicon 289 -1278 289 -1278 0 1
rlabel polysilicon 289 -1284 289 -1284 0 3
rlabel polysilicon 296 -1278 296 -1278 0 1
rlabel polysilicon 296 -1284 296 -1284 0 3
rlabel polysilicon 303 -1278 303 -1278 0 1
rlabel polysilicon 303 -1284 303 -1284 0 3
rlabel polysilicon 310 -1278 310 -1278 0 1
rlabel polysilicon 310 -1284 310 -1284 0 3
rlabel polysilicon 317 -1278 317 -1278 0 1
rlabel polysilicon 320 -1278 320 -1278 0 2
rlabel polysilicon 317 -1284 317 -1284 0 3
rlabel polysilicon 320 -1284 320 -1284 0 4
rlabel polysilicon 324 -1278 324 -1278 0 1
rlabel polysilicon 324 -1284 324 -1284 0 3
rlabel polysilicon 331 -1278 331 -1278 0 1
rlabel polysilicon 331 -1284 331 -1284 0 3
rlabel polysilicon 338 -1278 338 -1278 0 1
rlabel polysilicon 341 -1278 341 -1278 0 2
rlabel polysilicon 345 -1278 345 -1278 0 1
rlabel polysilicon 345 -1284 345 -1284 0 3
rlabel polysilicon 352 -1278 352 -1278 0 1
rlabel polysilicon 352 -1284 352 -1284 0 3
rlabel polysilicon 359 -1278 359 -1278 0 1
rlabel polysilicon 362 -1278 362 -1278 0 2
rlabel polysilicon 359 -1284 359 -1284 0 3
rlabel polysilicon 362 -1284 362 -1284 0 4
rlabel polysilicon 366 -1278 366 -1278 0 1
rlabel polysilicon 366 -1284 366 -1284 0 3
rlabel polysilicon 373 -1278 373 -1278 0 1
rlabel polysilicon 373 -1284 373 -1284 0 3
rlabel polysilicon 380 -1278 380 -1278 0 1
rlabel polysilicon 380 -1284 380 -1284 0 3
rlabel polysilicon 387 -1278 387 -1278 0 1
rlabel polysilicon 387 -1284 387 -1284 0 3
rlabel polysilicon 394 -1278 394 -1278 0 1
rlabel polysilicon 394 -1284 394 -1284 0 3
rlabel polysilicon 401 -1278 401 -1278 0 1
rlabel polysilicon 401 -1284 401 -1284 0 3
rlabel polysilicon 408 -1278 408 -1278 0 1
rlabel polysilicon 408 -1284 408 -1284 0 3
rlabel polysilicon 415 -1278 415 -1278 0 1
rlabel polysilicon 415 -1284 415 -1284 0 3
rlabel polysilicon 422 -1278 422 -1278 0 1
rlabel polysilicon 422 -1284 422 -1284 0 3
rlabel polysilicon 429 -1278 429 -1278 0 1
rlabel polysilicon 429 -1284 429 -1284 0 3
rlabel polysilicon 436 -1278 436 -1278 0 1
rlabel polysilicon 436 -1284 436 -1284 0 3
rlabel polysilicon 443 -1278 443 -1278 0 1
rlabel polysilicon 443 -1284 443 -1284 0 3
rlabel polysilicon 450 -1278 450 -1278 0 1
rlabel polysilicon 450 -1284 450 -1284 0 3
rlabel polysilicon 457 -1278 457 -1278 0 1
rlabel polysilicon 457 -1284 457 -1284 0 3
rlabel polysilicon 464 -1278 464 -1278 0 1
rlabel polysilicon 464 -1284 464 -1284 0 3
rlabel polysilicon 471 -1278 471 -1278 0 1
rlabel polysilicon 471 -1284 471 -1284 0 3
rlabel polysilicon 478 -1278 478 -1278 0 1
rlabel polysilicon 481 -1278 481 -1278 0 2
rlabel polysilicon 478 -1284 478 -1284 0 3
rlabel polysilicon 481 -1284 481 -1284 0 4
rlabel polysilicon 485 -1278 485 -1278 0 1
rlabel polysilicon 485 -1284 485 -1284 0 3
rlabel polysilicon 492 -1278 492 -1278 0 1
rlabel polysilicon 492 -1284 492 -1284 0 3
rlabel polysilicon 499 -1278 499 -1278 0 1
rlabel polysilicon 499 -1284 499 -1284 0 3
rlabel polysilicon 506 -1278 506 -1278 0 1
rlabel polysilicon 509 -1278 509 -1278 0 2
rlabel polysilicon 506 -1284 506 -1284 0 3
rlabel polysilicon 509 -1284 509 -1284 0 4
rlabel polysilicon 513 -1278 513 -1278 0 1
rlabel polysilicon 513 -1284 513 -1284 0 3
rlabel polysilicon 520 -1278 520 -1278 0 1
rlabel polysilicon 520 -1284 520 -1284 0 3
rlabel polysilicon 523 -1284 523 -1284 0 4
rlabel polysilicon 527 -1278 527 -1278 0 1
rlabel polysilicon 530 -1278 530 -1278 0 2
rlabel polysilicon 527 -1284 527 -1284 0 3
rlabel polysilicon 530 -1284 530 -1284 0 4
rlabel polysilicon 534 -1278 534 -1278 0 1
rlabel polysilicon 534 -1284 534 -1284 0 3
rlabel polysilicon 541 -1278 541 -1278 0 1
rlabel polysilicon 541 -1284 541 -1284 0 3
rlabel polysilicon 548 -1278 548 -1278 0 1
rlabel polysilicon 548 -1284 548 -1284 0 3
rlabel polysilicon 551 -1284 551 -1284 0 4
rlabel polysilicon 555 -1278 555 -1278 0 1
rlabel polysilicon 558 -1278 558 -1278 0 2
rlabel polysilicon 555 -1284 555 -1284 0 3
rlabel polysilicon 558 -1284 558 -1284 0 4
rlabel polysilicon 562 -1278 562 -1278 0 1
rlabel polysilicon 562 -1284 562 -1284 0 3
rlabel polysilicon 569 -1278 569 -1278 0 1
rlabel polysilicon 569 -1284 569 -1284 0 3
rlabel polysilicon 576 -1278 576 -1278 0 1
rlabel polysilicon 576 -1284 576 -1284 0 3
rlabel polysilicon 583 -1278 583 -1278 0 1
rlabel polysilicon 583 -1284 583 -1284 0 3
rlabel polysilicon 590 -1278 590 -1278 0 1
rlabel polysilicon 590 -1284 590 -1284 0 3
rlabel polysilicon 597 -1278 597 -1278 0 1
rlabel polysilicon 597 -1284 597 -1284 0 3
rlabel polysilicon 604 -1278 604 -1278 0 1
rlabel polysilicon 607 -1278 607 -1278 0 2
rlabel polysilicon 604 -1284 604 -1284 0 3
rlabel polysilicon 607 -1284 607 -1284 0 4
rlabel polysilicon 611 -1278 611 -1278 0 1
rlabel polysilicon 611 -1284 611 -1284 0 3
rlabel polysilicon 618 -1278 618 -1278 0 1
rlabel polysilicon 618 -1284 618 -1284 0 3
rlabel polysilicon 625 -1278 625 -1278 0 1
rlabel polysilicon 625 -1284 625 -1284 0 3
rlabel polysilicon 632 -1278 632 -1278 0 1
rlabel polysilicon 632 -1284 632 -1284 0 3
rlabel polysilicon 639 -1278 639 -1278 0 1
rlabel polysilicon 639 -1284 639 -1284 0 3
rlabel polysilicon 646 -1278 646 -1278 0 1
rlabel polysilicon 646 -1284 646 -1284 0 3
rlabel polysilicon 653 -1278 653 -1278 0 1
rlabel polysilicon 653 -1284 653 -1284 0 3
rlabel polysilicon 660 -1278 660 -1278 0 1
rlabel polysilicon 660 -1284 660 -1284 0 3
rlabel polysilicon 667 -1278 667 -1278 0 1
rlabel polysilicon 667 -1284 667 -1284 0 3
rlabel polysilicon 674 -1278 674 -1278 0 1
rlabel polysilicon 674 -1284 674 -1284 0 3
rlabel polysilicon 681 -1278 681 -1278 0 1
rlabel polysilicon 681 -1284 681 -1284 0 3
rlabel polysilicon 688 -1278 688 -1278 0 1
rlabel polysilicon 688 -1284 688 -1284 0 3
rlabel polysilicon 695 -1278 695 -1278 0 1
rlabel polysilicon 695 -1284 695 -1284 0 3
rlabel polysilicon 702 -1278 702 -1278 0 1
rlabel polysilicon 702 -1284 702 -1284 0 3
rlabel polysilicon 709 -1278 709 -1278 0 1
rlabel polysilicon 709 -1284 709 -1284 0 3
rlabel polysilicon 716 -1278 716 -1278 0 1
rlabel polysilicon 719 -1278 719 -1278 0 2
rlabel polysilicon 716 -1284 716 -1284 0 3
rlabel polysilicon 719 -1284 719 -1284 0 4
rlabel polysilicon 723 -1278 723 -1278 0 1
rlabel polysilicon 726 -1278 726 -1278 0 2
rlabel polysilicon 723 -1284 723 -1284 0 3
rlabel polysilicon 726 -1284 726 -1284 0 4
rlabel polysilicon 730 -1278 730 -1278 0 1
rlabel polysilicon 730 -1284 730 -1284 0 3
rlabel polysilicon 737 -1278 737 -1278 0 1
rlabel polysilicon 737 -1284 737 -1284 0 3
rlabel polysilicon 744 -1278 744 -1278 0 1
rlabel polysilicon 744 -1284 744 -1284 0 3
rlabel polysilicon 751 -1278 751 -1278 0 1
rlabel polysilicon 754 -1278 754 -1278 0 2
rlabel polysilicon 751 -1284 751 -1284 0 3
rlabel polysilicon 754 -1284 754 -1284 0 4
rlabel polysilicon 758 -1278 758 -1278 0 1
rlabel polysilicon 758 -1284 758 -1284 0 3
rlabel polysilicon 765 -1278 765 -1278 0 1
rlabel polysilicon 768 -1278 768 -1278 0 2
rlabel polysilicon 765 -1284 765 -1284 0 3
rlabel polysilicon 768 -1284 768 -1284 0 4
rlabel polysilicon 772 -1278 772 -1278 0 1
rlabel polysilicon 772 -1284 772 -1284 0 3
rlabel polysilicon 779 -1278 779 -1278 0 1
rlabel polysilicon 782 -1278 782 -1278 0 2
rlabel polysilicon 779 -1284 779 -1284 0 3
rlabel polysilicon 782 -1284 782 -1284 0 4
rlabel polysilicon 786 -1278 786 -1278 0 1
rlabel polysilicon 786 -1284 786 -1284 0 3
rlabel polysilicon 793 -1278 793 -1278 0 1
rlabel polysilicon 793 -1284 793 -1284 0 3
rlabel polysilicon 800 -1278 800 -1278 0 1
rlabel polysilicon 800 -1284 800 -1284 0 3
rlabel polysilicon 807 -1278 807 -1278 0 1
rlabel polysilicon 807 -1284 807 -1284 0 3
rlabel polysilicon 814 -1278 814 -1278 0 1
rlabel polysilicon 814 -1284 814 -1284 0 3
rlabel polysilicon 821 -1278 821 -1278 0 1
rlabel polysilicon 821 -1284 821 -1284 0 3
rlabel polysilicon 828 -1278 828 -1278 0 1
rlabel polysilicon 828 -1284 828 -1284 0 3
rlabel polysilicon 835 -1278 835 -1278 0 1
rlabel polysilicon 838 -1278 838 -1278 0 2
rlabel polysilicon 835 -1284 835 -1284 0 3
rlabel polysilicon 838 -1284 838 -1284 0 4
rlabel polysilicon 842 -1278 842 -1278 0 1
rlabel polysilicon 842 -1284 842 -1284 0 3
rlabel polysilicon 849 -1278 849 -1278 0 1
rlabel polysilicon 849 -1284 849 -1284 0 3
rlabel polysilicon 856 -1278 856 -1278 0 1
rlabel polysilicon 859 -1278 859 -1278 0 2
rlabel polysilicon 856 -1284 856 -1284 0 3
rlabel polysilicon 859 -1284 859 -1284 0 4
rlabel polysilicon 863 -1278 863 -1278 0 1
rlabel polysilicon 863 -1284 863 -1284 0 3
rlabel polysilicon 870 -1278 870 -1278 0 1
rlabel polysilicon 870 -1284 870 -1284 0 3
rlabel polysilicon 877 -1278 877 -1278 0 1
rlabel polysilicon 877 -1284 877 -1284 0 3
rlabel polysilicon 884 -1278 884 -1278 0 1
rlabel polysilicon 884 -1284 884 -1284 0 3
rlabel polysilicon 891 -1278 891 -1278 0 1
rlabel polysilicon 891 -1284 891 -1284 0 3
rlabel polysilicon 898 -1278 898 -1278 0 1
rlabel polysilicon 898 -1284 898 -1284 0 3
rlabel polysilicon 905 -1278 905 -1278 0 1
rlabel polysilicon 905 -1284 905 -1284 0 3
rlabel polysilicon 912 -1278 912 -1278 0 1
rlabel polysilicon 912 -1284 912 -1284 0 3
rlabel polysilicon 919 -1278 919 -1278 0 1
rlabel polysilicon 922 -1278 922 -1278 0 2
rlabel polysilicon 922 -1284 922 -1284 0 4
rlabel polysilicon 926 -1278 926 -1278 0 1
rlabel polysilicon 926 -1284 926 -1284 0 3
rlabel polysilicon 933 -1278 933 -1278 0 1
rlabel polysilicon 936 -1278 936 -1278 0 2
rlabel polysilicon 933 -1284 933 -1284 0 3
rlabel polysilicon 940 -1278 940 -1278 0 1
rlabel polysilicon 940 -1284 940 -1284 0 3
rlabel polysilicon 947 -1278 947 -1278 0 1
rlabel polysilicon 947 -1284 947 -1284 0 3
rlabel polysilicon 954 -1278 954 -1278 0 1
rlabel polysilicon 954 -1284 954 -1284 0 3
rlabel polysilicon 961 -1278 961 -1278 0 1
rlabel polysilicon 961 -1284 961 -1284 0 3
rlabel polysilicon 968 -1278 968 -1278 0 1
rlabel polysilicon 968 -1284 968 -1284 0 3
rlabel polysilicon 975 -1278 975 -1278 0 1
rlabel polysilicon 975 -1284 975 -1284 0 3
rlabel polysilicon 982 -1278 982 -1278 0 1
rlabel polysilicon 982 -1284 982 -1284 0 3
rlabel polysilicon 989 -1278 989 -1278 0 1
rlabel polysilicon 989 -1284 989 -1284 0 3
rlabel polysilicon 996 -1278 996 -1278 0 1
rlabel polysilicon 996 -1284 996 -1284 0 3
rlabel polysilicon 1003 -1278 1003 -1278 0 1
rlabel polysilicon 1003 -1284 1003 -1284 0 3
rlabel polysilicon 1010 -1278 1010 -1278 0 1
rlabel polysilicon 1010 -1284 1010 -1284 0 3
rlabel polysilicon 1017 -1278 1017 -1278 0 1
rlabel polysilicon 1017 -1284 1017 -1284 0 3
rlabel polysilicon 1024 -1278 1024 -1278 0 1
rlabel polysilicon 1024 -1284 1024 -1284 0 3
rlabel polysilicon 1031 -1284 1031 -1284 0 3
rlabel polysilicon 1038 -1278 1038 -1278 0 1
rlabel polysilicon 1038 -1284 1038 -1284 0 3
rlabel polysilicon 1045 -1278 1045 -1278 0 1
rlabel polysilicon 1045 -1284 1045 -1284 0 3
rlabel polysilicon 1052 -1278 1052 -1278 0 1
rlabel polysilicon 1055 -1278 1055 -1278 0 2
rlabel polysilicon 1052 -1284 1052 -1284 0 3
rlabel polysilicon 1055 -1284 1055 -1284 0 4
rlabel polysilicon 1059 -1278 1059 -1278 0 1
rlabel polysilicon 1059 -1284 1059 -1284 0 3
rlabel polysilicon 1066 -1278 1066 -1278 0 1
rlabel polysilicon 1066 -1284 1066 -1284 0 3
rlabel polysilicon 1073 -1278 1073 -1278 0 1
rlabel polysilicon 1073 -1284 1073 -1284 0 3
rlabel polysilicon 1080 -1278 1080 -1278 0 1
rlabel polysilicon 1080 -1284 1080 -1284 0 3
rlabel polysilicon 1087 -1278 1087 -1278 0 1
rlabel polysilicon 1087 -1284 1087 -1284 0 3
rlabel polysilicon 1094 -1278 1094 -1278 0 1
rlabel polysilicon 1094 -1284 1094 -1284 0 3
rlabel polysilicon 1101 -1278 1101 -1278 0 1
rlabel polysilicon 1101 -1284 1101 -1284 0 3
rlabel polysilicon 1108 -1278 1108 -1278 0 1
rlabel polysilicon 1108 -1284 1108 -1284 0 3
rlabel polysilicon 1115 -1278 1115 -1278 0 1
rlabel polysilicon 1115 -1284 1115 -1284 0 3
rlabel polysilicon 1122 -1278 1122 -1278 0 1
rlabel polysilicon 1122 -1284 1122 -1284 0 3
rlabel polysilicon 1129 -1278 1129 -1278 0 1
rlabel polysilicon 1129 -1284 1129 -1284 0 3
rlabel polysilicon 1136 -1278 1136 -1278 0 1
rlabel polysilicon 1136 -1284 1136 -1284 0 3
rlabel polysilicon 1143 -1278 1143 -1278 0 1
rlabel polysilicon 1143 -1284 1143 -1284 0 3
rlabel polysilicon 1150 -1278 1150 -1278 0 1
rlabel polysilicon 1150 -1284 1150 -1284 0 3
rlabel polysilicon 1157 -1278 1157 -1278 0 1
rlabel polysilicon 1157 -1284 1157 -1284 0 3
rlabel polysilicon 1164 -1278 1164 -1278 0 1
rlabel polysilicon 1164 -1284 1164 -1284 0 3
rlabel polysilicon 1174 -1278 1174 -1278 0 2
rlabel polysilicon 1171 -1284 1171 -1284 0 3
rlabel polysilicon 1178 -1278 1178 -1278 0 1
rlabel polysilicon 1178 -1284 1178 -1284 0 3
rlabel polysilicon 1185 -1278 1185 -1278 0 1
rlabel polysilicon 1185 -1284 1185 -1284 0 3
rlabel polysilicon 1192 -1278 1192 -1278 0 1
rlabel polysilicon 1192 -1284 1192 -1284 0 3
rlabel polysilicon 1199 -1278 1199 -1278 0 1
rlabel polysilicon 1199 -1284 1199 -1284 0 3
rlabel polysilicon 1206 -1278 1206 -1278 0 1
rlabel polysilicon 1206 -1284 1206 -1284 0 3
rlabel polysilicon 1213 -1278 1213 -1278 0 1
rlabel polysilicon 1213 -1284 1213 -1284 0 3
rlabel polysilicon 1220 -1278 1220 -1278 0 1
rlabel polysilicon 1220 -1284 1220 -1284 0 3
rlabel polysilicon 1227 -1278 1227 -1278 0 1
rlabel polysilicon 1227 -1284 1227 -1284 0 3
rlabel polysilicon 1234 -1278 1234 -1278 0 1
rlabel polysilicon 1234 -1284 1234 -1284 0 3
rlabel polysilicon 1241 -1278 1241 -1278 0 1
rlabel polysilicon 1241 -1284 1241 -1284 0 3
rlabel polysilicon 1248 -1278 1248 -1278 0 1
rlabel polysilicon 1251 -1278 1251 -1278 0 2
rlabel polysilicon 1248 -1284 1248 -1284 0 3
rlabel polysilicon 1255 -1278 1255 -1278 0 1
rlabel polysilicon 1255 -1284 1255 -1284 0 3
rlabel polysilicon 1262 -1278 1262 -1278 0 1
rlabel polysilicon 1262 -1284 1262 -1284 0 3
rlabel polysilicon 1269 -1278 1269 -1278 0 1
rlabel polysilicon 1269 -1284 1269 -1284 0 3
rlabel polysilicon 1276 -1278 1276 -1278 0 1
rlabel polysilicon 1276 -1284 1276 -1284 0 3
rlabel polysilicon 1283 -1278 1283 -1278 0 1
rlabel polysilicon 1283 -1284 1283 -1284 0 3
rlabel polysilicon 1290 -1278 1290 -1278 0 1
rlabel polysilicon 1290 -1284 1290 -1284 0 3
rlabel polysilicon 1297 -1278 1297 -1278 0 1
rlabel polysilicon 1297 -1284 1297 -1284 0 3
rlabel polysilicon 1304 -1278 1304 -1278 0 1
rlabel polysilicon 1304 -1284 1304 -1284 0 3
rlabel polysilicon 1311 -1278 1311 -1278 0 1
rlabel polysilicon 1311 -1284 1311 -1284 0 3
rlabel polysilicon 1318 -1278 1318 -1278 0 1
rlabel polysilicon 1318 -1284 1318 -1284 0 3
rlabel polysilicon 1325 -1278 1325 -1278 0 1
rlabel polysilicon 1325 -1284 1325 -1284 0 3
rlabel polysilicon 1332 -1278 1332 -1278 0 1
rlabel polysilicon 1332 -1284 1332 -1284 0 3
rlabel polysilicon 1339 -1278 1339 -1278 0 1
rlabel polysilicon 1339 -1284 1339 -1284 0 3
rlabel polysilicon 1346 -1278 1346 -1278 0 1
rlabel polysilicon 1346 -1284 1346 -1284 0 3
rlabel polysilicon 1353 -1278 1353 -1278 0 1
rlabel polysilicon 1353 -1284 1353 -1284 0 3
rlabel polysilicon 1360 -1278 1360 -1278 0 1
rlabel polysilicon 1360 -1284 1360 -1284 0 3
rlabel polysilicon 1367 -1278 1367 -1278 0 1
rlabel polysilicon 1367 -1284 1367 -1284 0 3
rlabel polysilicon 1374 -1278 1374 -1278 0 1
rlabel polysilicon 1374 -1284 1374 -1284 0 3
rlabel polysilicon 1381 -1278 1381 -1278 0 1
rlabel polysilicon 1381 -1284 1381 -1284 0 3
rlabel polysilicon 1388 -1278 1388 -1278 0 1
rlabel polysilicon 1388 -1284 1388 -1284 0 3
rlabel polysilicon 1395 -1278 1395 -1278 0 1
rlabel polysilicon 1395 -1284 1395 -1284 0 3
rlabel polysilicon 1402 -1278 1402 -1278 0 1
rlabel polysilicon 1402 -1284 1402 -1284 0 3
rlabel polysilicon 1409 -1278 1409 -1278 0 1
rlabel polysilicon 1409 -1284 1409 -1284 0 3
rlabel polysilicon 1416 -1278 1416 -1278 0 1
rlabel polysilicon 1416 -1284 1416 -1284 0 3
rlabel polysilicon 1423 -1278 1423 -1278 0 1
rlabel polysilicon 1423 -1284 1423 -1284 0 3
rlabel polysilicon 1430 -1278 1430 -1278 0 1
rlabel polysilicon 1430 -1284 1430 -1284 0 3
rlabel polysilicon 1437 -1278 1437 -1278 0 1
rlabel polysilicon 1437 -1284 1437 -1284 0 3
rlabel polysilicon 1444 -1278 1444 -1278 0 1
rlabel polysilicon 1444 -1284 1444 -1284 0 3
rlabel polysilicon 1451 -1278 1451 -1278 0 1
rlabel polysilicon 1451 -1284 1451 -1284 0 3
rlabel polysilicon 1458 -1278 1458 -1278 0 1
rlabel polysilicon 1458 -1284 1458 -1284 0 3
rlabel polysilicon 1465 -1278 1465 -1278 0 1
rlabel polysilicon 1465 -1284 1465 -1284 0 3
rlabel polysilicon 1472 -1278 1472 -1278 0 1
rlabel polysilicon 1472 -1284 1472 -1284 0 3
rlabel polysilicon 1479 -1278 1479 -1278 0 1
rlabel polysilicon 1479 -1284 1479 -1284 0 3
rlabel polysilicon 1486 -1278 1486 -1278 0 1
rlabel polysilicon 1486 -1284 1486 -1284 0 3
rlabel polysilicon 1493 -1278 1493 -1278 0 1
rlabel polysilicon 1493 -1284 1493 -1284 0 3
rlabel polysilicon 1500 -1278 1500 -1278 0 1
rlabel polysilicon 1500 -1284 1500 -1284 0 3
rlabel polysilicon 1507 -1278 1507 -1278 0 1
rlabel polysilicon 1507 -1284 1507 -1284 0 3
rlabel polysilicon 1514 -1278 1514 -1278 0 1
rlabel polysilicon 1514 -1284 1514 -1284 0 3
rlabel polysilicon 1521 -1278 1521 -1278 0 1
rlabel polysilicon 1521 -1284 1521 -1284 0 3
rlabel polysilicon 1528 -1278 1528 -1278 0 1
rlabel polysilicon 1528 -1284 1528 -1284 0 3
rlabel polysilicon 1535 -1278 1535 -1278 0 1
rlabel polysilicon 1535 -1284 1535 -1284 0 3
rlabel polysilicon 1542 -1278 1542 -1278 0 1
rlabel polysilicon 1542 -1284 1542 -1284 0 3
rlabel polysilicon 1549 -1278 1549 -1278 0 1
rlabel polysilicon 1549 -1284 1549 -1284 0 3
rlabel polysilicon 1556 -1278 1556 -1278 0 1
rlabel polysilicon 1556 -1284 1556 -1284 0 3
rlabel polysilicon 1563 -1278 1563 -1278 0 1
rlabel polysilicon 1563 -1284 1563 -1284 0 3
rlabel polysilicon 2 -1397 2 -1397 0 1
rlabel polysilicon 2 -1403 2 -1403 0 3
rlabel polysilicon 9 -1397 9 -1397 0 1
rlabel polysilicon 9 -1403 9 -1403 0 3
rlabel polysilicon 16 -1397 16 -1397 0 1
rlabel polysilicon 16 -1403 16 -1403 0 3
rlabel polysilicon 23 -1397 23 -1397 0 1
rlabel polysilicon 23 -1403 23 -1403 0 3
rlabel polysilicon 30 -1397 30 -1397 0 1
rlabel polysilicon 30 -1403 30 -1403 0 3
rlabel polysilicon 37 -1397 37 -1397 0 1
rlabel polysilicon 37 -1403 37 -1403 0 3
rlabel polysilicon 44 -1397 44 -1397 0 1
rlabel polysilicon 44 -1403 44 -1403 0 3
rlabel polysilicon 51 -1397 51 -1397 0 1
rlabel polysilicon 51 -1403 51 -1403 0 3
rlabel polysilicon 58 -1397 58 -1397 0 1
rlabel polysilicon 58 -1403 58 -1403 0 3
rlabel polysilicon 65 -1397 65 -1397 0 1
rlabel polysilicon 68 -1397 68 -1397 0 2
rlabel polysilicon 65 -1403 65 -1403 0 3
rlabel polysilicon 68 -1403 68 -1403 0 4
rlabel polysilicon 72 -1397 72 -1397 0 1
rlabel polysilicon 72 -1403 72 -1403 0 3
rlabel polysilicon 79 -1397 79 -1397 0 1
rlabel polysilicon 82 -1397 82 -1397 0 2
rlabel polysilicon 79 -1403 79 -1403 0 3
rlabel polysilicon 82 -1403 82 -1403 0 4
rlabel polysilicon 86 -1397 86 -1397 0 1
rlabel polysilicon 86 -1403 86 -1403 0 3
rlabel polysilicon 93 -1397 93 -1397 0 1
rlabel polysilicon 93 -1403 93 -1403 0 3
rlabel polysilicon 100 -1397 100 -1397 0 1
rlabel polysilicon 100 -1403 100 -1403 0 3
rlabel polysilicon 107 -1397 107 -1397 0 1
rlabel polysilicon 110 -1397 110 -1397 0 2
rlabel polysilicon 107 -1403 107 -1403 0 3
rlabel polysilicon 110 -1403 110 -1403 0 4
rlabel polysilicon 114 -1397 114 -1397 0 1
rlabel polysilicon 114 -1403 114 -1403 0 3
rlabel polysilicon 121 -1397 121 -1397 0 1
rlabel polysilicon 121 -1403 121 -1403 0 3
rlabel polysilicon 128 -1397 128 -1397 0 1
rlabel polysilicon 128 -1403 128 -1403 0 3
rlabel polysilicon 135 -1397 135 -1397 0 1
rlabel polysilicon 135 -1403 135 -1403 0 3
rlabel polysilicon 142 -1397 142 -1397 0 1
rlabel polysilicon 142 -1403 142 -1403 0 3
rlabel polysilicon 149 -1397 149 -1397 0 1
rlabel polysilicon 149 -1403 149 -1403 0 3
rlabel polysilicon 156 -1397 156 -1397 0 1
rlabel polysilicon 156 -1403 156 -1403 0 3
rlabel polysilicon 163 -1397 163 -1397 0 1
rlabel polysilicon 163 -1403 163 -1403 0 3
rlabel polysilicon 170 -1397 170 -1397 0 1
rlabel polysilicon 170 -1403 170 -1403 0 3
rlabel polysilicon 177 -1397 177 -1397 0 1
rlabel polysilicon 177 -1403 177 -1403 0 3
rlabel polysilicon 184 -1397 184 -1397 0 1
rlabel polysilicon 184 -1403 184 -1403 0 3
rlabel polysilicon 191 -1397 191 -1397 0 1
rlabel polysilicon 191 -1403 191 -1403 0 3
rlabel polysilicon 198 -1397 198 -1397 0 1
rlabel polysilicon 198 -1403 198 -1403 0 3
rlabel polysilicon 205 -1397 205 -1397 0 1
rlabel polysilicon 205 -1403 205 -1403 0 3
rlabel polysilicon 212 -1397 212 -1397 0 1
rlabel polysilicon 215 -1397 215 -1397 0 2
rlabel polysilicon 212 -1403 212 -1403 0 3
rlabel polysilicon 219 -1397 219 -1397 0 1
rlabel polysilicon 219 -1403 219 -1403 0 3
rlabel polysilicon 226 -1397 226 -1397 0 1
rlabel polysilicon 226 -1403 226 -1403 0 3
rlabel polysilicon 233 -1397 233 -1397 0 1
rlabel polysilicon 233 -1403 233 -1403 0 3
rlabel polysilicon 240 -1397 240 -1397 0 1
rlabel polysilicon 240 -1403 240 -1403 0 3
rlabel polysilicon 247 -1397 247 -1397 0 1
rlabel polysilicon 247 -1403 247 -1403 0 3
rlabel polysilicon 254 -1397 254 -1397 0 1
rlabel polysilicon 254 -1403 254 -1403 0 3
rlabel polysilicon 261 -1397 261 -1397 0 1
rlabel polysilicon 261 -1403 261 -1403 0 3
rlabel polysilicon 268 -1397 268 -1397 0 1
rlabel polysilicon 268 -1403 268 -1403 0 3
rlabel polysilicon 275 -1397 275 -1397 0 1
rlabel polysilicon 275 -1403 275 -1403 0 3
rlabel polysilicon 282 -1397 282 -1397 0 1
rlabel polysilicon 282 -1403 282 -1403 0 3
rlabel polysilicon 289 -1397 289 -1397 0 1
rlabel polysilicon 289 -1403 289 -1403 0 3
rlabel polysilicon 296 -1397 296 -1397 0 1
rlabel polysilicon 296 -1403 296 -1403 0 3
rlabel polysilicon 303 -1397 303 -1397 0 1
rlabel polysilicon 303 -1403 303 -1403 0 3
rlabel polysilicon 310 -1397 310 -1397 0 1
rlabel polysilicon 310 -1403 310 -1403 0 3
rlabel polysilicon 317 -1397 317 -1397 0 1
rlabel polysilicon 320 -1397 320 -1397 0 2
rlabel polysilicon 317 -1403 317 -1403 0 3
rlabel polysilicon 320 -1403 320 -1403 0 4
rlabel polysilicon 324 -1397 324 -1397 0 1
rlabel polysilicon 324 -1403 324 -1403 0 3
rlabel polysilicon 331 -1397 331 -1397 0 1
rlabel polysilicon 331 -1403 331 -1403 0 3
rlabel polysilicon 338 -1397 338 -1397 0 1
rlabel polysilicon 338 -1403 338 -1403 0 3
rlabel polysilicon 345 -1397 345 -1397 0 1
rlabel polysilicon 345 -1403 345 -1403 0 3
rlabel polysilicon 352 -1397 352 -1397 0 1
rlabel polysilicon 352 -1403 352 -1403 0 3
rlabel polysilicon 359 -1397 359 -1397 0 1
rlabel polysilicon 359 -1403 359 -1403 0 3
rlabel polysilicon 366 -1397 366 -1397 0 1
rlabel polysilicon 366 -1403 366 -1403 0 3
rlabel polysilicon 373 -1397 373 -1397 0 1
rlabel polysilicon 373 -1403 373 -1403 0 3
rlabel polysilicon 380 -1397 380 -1397 0 1
rlabel polysilicon 380 -1403 380 -1403 0 3
rlabel polysilicon 387 -1397 387 -1397 0 1
rlabel polysilicon 390 -1397 390 -1397 0 2
rlabel polysilicon 387 -1403 387 -1403 0 3
rlabel polysilicon 390 -1403 390 -1403 0 4
rlabel polysilicon 394 -1397 394 -1397 0 1
rlabel polysilicon 394 -1403 394 -1403 0 3
rlabel polysilicon 404 -1397 404 -1397 0 2
rlabel polysilicon 401 -1403 401 -1403 0 3
rlabel polysilicon 404 -1403 404 -1403 0 4
rlabel polysilicon 408 -1397 408 -1397 0 1
rlabel polysilicon 408 -1403 408 -1403 0 3
rlabel polysilicon 418 -1397 418 -1397 0 2
rlabel polysilicon 415 -1403 415 -1403 0 3
rlabel polysilicon 418 -1403 418 -1403 0 4
rlabel polysilicon 422 -1397 422 -1397 0 1
rlabel polysilicon 422 -1403 422 -1403 0 3
rlabel polysilicon 429 -1397 429 -1397 0 1
rlabel polysilicon 429 -1403 429 -1403 0 3
rlabel polysilicon 436 -1397 436 -1397 0 1
rlabel polysilicon 436 -1403 436 -1403 0 3
rlabel polysilicon 443 -1397 443 -1397 0 1
rlabel polysilicon 443 -1403 443 -1403 0 3
rlabel polysilicon 450 -1397 450 -1397 0 1
rlabel polysilicon 450 -1403 450 -1403 0 3
rlabel polysilicon 457 -1397 457 -1397 0 1
rlabel polysilicon 457 -1403 457 -1403 0 3
rlabel polysilicon 464 -1397 464 -1397 0 1
rlabel polysilicon 467 -1397 467 -1397 0 2
rlabel polysilicon 464 -1403 464 -1403 0 3
rlabel polysilicon 467 -1403 467 -1403 0 4
rlabel polysilicon 471 -1397 471 -1397 0 1
rlabel polysilicon 471 -1403 471 -1403 0 3
rlabel polysilicon 478 -1397 478 -1397 0 1
rlabel polysilicon 481 -1397 481 -1397 0 2
rlabel polysilicon 478 -1403 478 -1403 0 3
rlabel polysilicon 481 -1403 481 -1403 0 4
rlabel polysilicon 485 -1397 485 -1397 0 1
rlabel polysilicon 488 -1397 488 -1397 0 2
rlabel polysilicon 485 -1403 485 -1403 0 3
rlabel polysilicon 488 -1403 488 -1403 0 4
rlabel polysilicon 492 -1397 492 -1397 0 1
rlabel polysilicon 495 -1397 495 -1397 0 2
rlabel polysilicon 492 -1403 492 -1403 0 3
rlabel polysilicon 495 -1403 495 -1403 0 4
rlabel polysilicon 499 -1397 499 -1397 0 1
rlabel polysilicon 499 -1403 499 -1403 0 3
rlabel polysilicon 506 -1397 506 -1397 0 1
rlabel polysilicon 506 -1403 506 -1403 0 3
rlabel polysilicon 513 -1397 513 -1397 0 1
rlabel polysilicon 516 -1397 516 -1397 0 2
rlabel polysilicon 513 -1403 513 -1403 0 3
rlabel polysilicon 516 -1403 516 -1403 0 4
rlabel polysilicon 520 -1397 520 -1397 0 1
rlabel polysilicon 523 -1397 523 -1397 0 2
rlabel polysilicon 520 -1403 520 -1403 0 3
rlabel polysilicon 523 -1403 523 -1403 0 4
rlabel polysilicon 527 -1397 527 -1397 0 1
rlabel polysilicon 527 -1403 527 -1403 0 3
rlabel polysilicon 534 -1397 534 -1397 0 1
rlabel polysilicon 534 -1403 534 -1403 0 3
rlabel polysilicon 541 -1397 541 -1397 0 1
rlabel polysilicon 541 -1403 541 -1403 0 3
rlabel polysilicon 548 -1397 548 -1397 0 1
rlabel polysilicon 548 -1403 548 -1403 0 3
rlabel polysilicon 555 -1397 555 -1397 0 1
rlabel polysilicon 555 -1403 555 -1403 0 3
rlabel polysilicon 562 -1397 562 -1397 0 1
rlabel polysilicon 562 -1403 562 -1403 0 3
rlabel polysilicon 569 -1397 569 -1397 0 1
rlabel polysilicon 569 -1403 569 -1403 0 3
rlabel polysilicon 576 -1397 576 -1397 0 1
rlabel polysilicon 576 -1403 576 -1403 0 3
rlabel polysilicon 583 -1397 583 -1397 0 1
rlabel polysilicon 583 -1403 583 -1403 0 3
rlabel polysilicon 590 -1397 590 -1397 0 1
rlabel polysilicon 590 -1403 590 -1403 0 3
rlabel polysilicon 597 -1397 597 -1397 0 1
rlabel polysilicon 597 -1403 597 -1403 0 3
rlabel polysilicon 604 -1397 604 -1397 0 1
rlabel polysilicon 604 -1403 604 -1403 0 3
rlabel polysilicon 611 -1397 611 -1397 0 1
rlabel polysilicon 611 -1403 611 -1403 0 3
rlabel polysilicon 618 -1397 618 -1397 0 1
rlabel polysilicon 618 -1403 618 -1403 0 3
rlabel polysilicon 625 -1397 625 -1397 0 1
rlabel polysilicon 625 -1403 625 -1403 0 3
rlabel polysilicon 632 -1397 632 -1397 0 1
rlabel polysilicon 632 -1403 632 -1403 0 3
rlabel polysilicon 639 -1397 639 -1397 0 1
rlabel polysilicon 639 -1403 639 -1403 0 3
rlabel polysilicon 646 -1397 646 -1397 0 1
rlabel polysilicon 649 -1397 649 -1397 0 2
rlabel polysilicon 646 -1403 646 -1403 0 3
rlabel polysilicon 649 -1403 649 -1403 0 4
rlabel polysilicon 653 -1397 653 -1397 0 1
rlabel polysilicon 653 -1403 653 -1403 0 3
rlabel polysilicon 660 -1397 660 -1397 0 1
rlabel polysilicon 660 -1403 660 -1403 0 3
rlabel polysilicon 667 -1397 667 -1397 0 1
rlabel polysilicon 667 -1403 667 -1403 0 3
rlabel polysilicon 674 -1397 674 -1397 0 1
rlabel polysilicon 674 -1403 674 -1403 0 3
rlabel polysilicon 681 -1397 681 -1397 0 1
rlabel polysilicon 681 -1403 681 -1403 0 3
rlabel polysilicon 688 -1397 688 -1397 0 1
rlabel polysilicon 688 -1403 688 -1403 0 3
rlabel polysilicon 695 -1397 695 -1397 0 1
rlabel polysilicon 695 -1403 695 -1403 0 3
rlabel polysilicon 702 -1397 702 -1397 0 1
rlabel polysilicon 702 -1403 702 -1403 0 3
rlabel polysilicon 709 -1397 709 -1397 0 1
rlabel polysilicon 712 -1397 712 -1397 0 2
rlabel polysilicon 709 -1403 709 -1403 0 3
rlabel polysilicon 712 -1403 712 -1403 0 4
rlabel polysilicon 716 -1397 716 -1397 0 1
rlabel polysilicon 716 -1403 716 -1403 0 3
rlabel polysilicon 723 -1397 723 -1397 0 1
rlabel polysilicon 723 -1403 723 -1403 0 3
rlabel polysilicon 730 -1397 730 -1397 0 1
rlabel polysilicon 730 -1403 730 -1403 0 3
rlabel polysilicon 737 -1397 737 -1397 0 1
rlabel polysilicon 737 -1403 737 -1403 0 3
rlabel polysilicon 744 -1397 744 -1397 0 1
rlabel polysilicon 744 -1403 744 -1403 0 3
rlabel polysilicon 751 -1397 751 -1397 0 1
rlabel polysilicon 751 -1403 751 -1403 0 3
rlabel polysilicon 758 -1397 758 -1397 0 1
rlabel polysilicon 758 -1403 758 -1403 0 3
rlabel polysilicon 765 -1397 765 -1397 0 1
rlabel polysilicon 765 -1403 765 -1403 0 3
rlabel polysilicon 772 -1397 772 -1397 0 1
rlabel polysilicon 772 -1403 772 -1403 0 3
rlabel polysilicon 779 -1397 779 -1397 0 1
rlabel polysilicon 779 -1403 779 -1403 0 3
rlabel polysilicon 786 -1397 786 -1397 0 1
rlabel polysilicon 786 -1403 786 -1403 0 3
rlabel polysilicon 793 -1397 793 -1397 0 1
rlabel polysilicon 793 -1403 793 -1403 0 3
rlabel polysilicon 800 -1397 800 -1397 0 1
rlabel polysilicon 800 -1403 800 -1403 0 3
rlabel polysilicon 807 -1397 807 -1397 0 1
rlabel polysilicon 807 -1403 807 -1403 0 3
rlabel polysilicon 814 -1397 814 -1397 0 1
rlabel polysilicon 814 -1403 814 -1403 0 3
rlabel polysilicon 821 -1397 821 -1397 0 1
rlabel polysilicon 821 -1403 821 -1403 0 3
rlabel polysilicon 828 -1397 828 -1397 0 1
rlabel polysilicon 828 -1403 828 -1403 0 3
rlabel polysilicon 835 -1397 835 -1397 0 1
rlabel polysilicon 835 -1403 835 -1403 0 3
rlabel polysilicon 842 -1397 842 -1397 0 1
rlabel polysilicon 845 -1397 845 -1397 0 2
rlabel polysilicon 842 -1403 842 -1403 0 3
rlabel polysilicon 845 -1403 845 -1403 0 4
rlabel polysilicon 849 -1397 849 -1397 0 1
rlabel polysilicon 849 -1403 849 -1403 0 3
rlabel polysilicon 856 -1397 856 -1397 0 1
rlabel polysilicon 856 -1403 856 -1403 0 3
rlabel polysilicon 863 -1397 863 -1397 0 1
rlabel polysilicon 863 -1403 863 -1403 0 3
rlabel polysilicon 870 -1397 870 -1397 0 1
rlabel polysilicon 873 -1397 873 -1397 0 2
rlabel polysilicon 870 -1403 870 -1403 0 3
rlabel polysilicon 873 -1403 873 -1403 0 4
rlabel polysilicon 877 -1397 877 -1397 0 1
rlabel polysilicon 880 -1397 880 -1397 0 2
rlabel polysilicon 877 -1403 877 -1403 0 3
rlabel polysilicon 880 -1403 880 -1403 0 4
rlabel polysilicon 884 -1397 884 -1397 0 1
rlabel polysilicon 884 -1403 884 -1403 0 3
rlabel polysilicon 891 -1397 891 -1397 0 1
rlabel polysilicon 891 -1403 891 -1403 0 3
rlabel polysilicon 898 -1397 898 -1397 0 1
rlabel polysilicon 898 -1403 898 -1403 0 3
rlabel polysilicon 905 -1397 905 -1397 0 1
rlabel polysilicon 905 -1403 905 -1403 0 3
rlabel polysilicon 912 -1397 912 -1397 0 1
rlabel polysilicon 912 -1403 912 -1403 0 3
rlabel polysilicon 919 -1397 919 -1397 0 1
rlabel polysilicon 922 -1397 922 -1397 0 2
rlabel polysilicon 919 -1403 919 -1403 0 3
rlabel polysilicon 922 -1403 922 -1403 0 4
rlabel polysilicon 926 -1397 926 -1397 0 1
rlabel polysilicon 926 -1403 926 -1403 0 3
rlabel polysilicon 933 -1397 933 -1397 0 1
rlabel polysilicon 933 -1403 933 -1403 0 3
rlabel polysilicon 940 -1397 940 -1397 0 1
rlabel polysilicon 940 -1403 940 -1403 0 3
rlabel polysilicon 947 -1397 947 -1397 0 1
rlabel polysilicon 950 -1397 950 -1397 0 2
rlabel polysilicon 947 -1403 947 -1403 0 3
rlabel polysilicon 950 -1403 950 -1403 0 4
rlabel polysilicon 954 -1397 954 -1397 0 1
rlabel polysilicon 954 -1403 954 -1403 0 3
rlabel polysilicon 961 -1397 961 -1397 0 1
rlabel polysilicon 961 -1403 961 -1403 0 3
rlabel polysilicon 968 -1397 968 -1397 0 1
rlabel polysilicon 968 -1403 968 -1403 0 3
rlabel polysilicon 975 -1397 975 -1397 0 1
rlabel polysilicon 978 -1397 978 -1397 0 2
rlabel polysilicon 975 -1403 975 -1403 0 3
rlabel polysilicon 978 -1403 978 -1403 0 4
rlabel polysilicon 982 -1397 982 -1397 0 1
rlabel polysilicon 982 -1403 982 -1403 0 3
rlabel polysilicon 989 -1397 989 -1397 0 1
rlabel polysilicon 989 -1403 989 -1403 0 3
rlabel polysilicon 996 -1397 996 -1397 0 1
rlabel polysilicon 996 -1403 996 -1403 0 3
rlabel polysilicon 1003 -1397 1003 -1397 0 1
rlabel polysilicon 1006 -1397 1006 -1397 0 2
rlabel polysilicon 1006 -1403 1006 -1403 0 4
rlabel polysilicon 1010 -1397 1010 -1397 0 1
rlabel polysilicon 1010 -1403 1010 -1403 0 3
rlabel polysilicon 1017 -1397 1017 -1397 0 1
rlabel polysilicon 1017 -1403 1017 -1403 0 3
rlabel polysilicon 1020 -1403 1020 -1403 0 4
rlabel polysilicon 1024 -1397 1024 -1397 0 1
rlabel polysilicon 1024 -1403 1024 -1403 0 3
rlabel polysilicon 1031 -1397 1031 -1397 0 1
rlabel polysilicon 1031 -1403 1031 -1403 0 3
rlabel polysilicon 1038 -1397 1038 -1397 0 1
rlabel polysilicon 1038 -1403 1038 -1403 0 3
rlabel polysilicon 1045 -1397 1045 -1397 0 1
rlabel polysilicon 1045 -1403 1045 -1403 0 3
rlabel polysilicon 1052 -1397 1052 -1397 0 1
rlabel polysilicon 1052 -1403 1052 -1403 0 3
rlabel polysilicon 1059 -1397 1059 -1397 0 1
rlabel polysilicon 1059 -1403 1059 -1403 0 3
rlabel polysilicon 1066 -1397 1066 -1397 0 1
rlabel polysilicon 1066 -1403 1066 -1403 0 3
rlabel polysilicon 1073 -1397 1073 -1397 0 1
rlabel polysilicon 1073 -1403 1073 -1403 0 3
rlabel polysilicon 1080 -1397 1080 -1397 0 1
rlabel polysilicon 1080 -1403 1080 -1403 0 3
rlabel polysilicon 1087 -1397 1087 -1397 0 1
rlabel polysilicon 1087 -1403 1087 -1403 0 3
rlabel polysilicon 1094 -1397 1094 -1397 0 1
rlabel polysilicon 1094 -1403 1094 -1403 0 3
rlabel polysilicon 1101 -1397 1101 -1397 0 1
rlabel polysilicon 1101 -1403 1101 -1403 0 3
rlabel polysilicon 1108 -1397 1108 -1397 0 1
rlabel polysilicon 1108 -1403 1108 -1403 0 3
rlabel polysilicon 1115 -1397 1115 -1397 0 1
rlabel polysilicon 1115 -1403 1115 -1403 0 3
rlabel polysilicon 1122 -1397 1122 -1397 0 1
rlabel polysilicon 1122 -1403 1122 -1403 0 3
rlabel polysilicon 1129 -1397 1129 -1397 0 1
rlabel polysilicon 1129 -1403 1129 -1403 0 3
rlabel polysilicon 1136 -1397 1136 -1397 0 1
rlabel polysilicon 1136 -1403 1136 -1403 0 3
rlabel polysilicon 1143 -1397 1143 -1397 0 1
rlabel polysilicon 1143 -1403 1143 -1403 0 3
rlabel polysilicon 1150 -1397 1150 -1397 0 1
rlabel polysilicon 1150 -1403 1150 -1403 0 3
rlabel polysilicon 1157 -1397 1157 -1397 0 1
rlabel polysilicon 1157 -1403 1157 -1403 0 3
rlabel polysilicon 1164 -1397 1164 -1397 0 1
rlabel polysilicon 1164 -1403 1164 -1403 0 3
rlabel polysilicon 1171 -1397 1171 -1397 0 1
rlabel polysilicon 1171 -1403 1171 -1403 0 3
rlabel polysilicon 1178 -1397 1178 -1397 0 1
rlabel polysilicon 1178 -1403 1178 -1403 0 3
rlabel polysilicon 1185 -1397 1185 -1397 0 1
rlabel polysilicon 1185 -1403 1185 -1403 0 3
rlabel polysilicon 1192 -1397 1192 -1397 0 1
rlabel polysilicon 1192 -1403 1192 -1403 0 3
rlabel polysilicon 1199 -1397 1199 -1397 0 1
rlabel polysilicon 1199 -1403 1199 -1403 0 3
rlabel polysilicon 1206 -1397 1206 -1397 0 1
rlabel polysilicon 1206 -1403 1206 -1403 0 3
rlabel polysilicon 1213 -1397 1213 -1397 0 1
rlabel polysilicon 1213 -1403 1213 -1403 0 3
rlabel polysilicon 1220 -1397 1220 -1397 0 1
rlabel polysilicon 1220 -1403 1220 -1403 0 3
rlabel polysilicon 1227 -1397 1227 -1397 0 1
rlabel polysilicon 1227 -1403 1227 -1403 0 3
rlabel polysilicon 1234 -1397 1234 -1397 0 1
rlabel polysilicon 1234 -1403 1234 -1403 0 3
rlabel polysilicon 1241 -1397 1241 -1397 0 1
rlabel polysilicon 1241 -1403 1241 -1403 0 3
rlabel polysilicon 1248 -1397 1248 -1397 0 1
rlabel polysilicon 1248 -1403 1248 -1403 0 3
rlabel polysilicon 1255 -1397 1255 -1397 0 1
rlabel polysilicon 1255 -1403 1255 -1403 0 3
rlabel polysilicon 1262 -1397 1262 -1397 0 1
rlabel polysilicon 1262 -1403 1262 -1403 0 3
rlabel polysilicon 1269 -1397 1269 -1397 0 1
rlabel polysilicon 1269 -1403 1269 -1403 0 3
rlabel polysilicon 1276 -1397 1276 -1397 0 1
rlabel polysilicon 1276 -1403 1276 -1403 0 3
rlabel polysilicon 1283 -1397 1283 -1397 0 1
rlabel polysilicon 1283 -1403 1283 -1403 0 3
rlabel polysilicon 1290 -1397 1290 -1397 0 1
rlabel polysilicon 1290 -1403 1290 -1403 0 3
rlabel polysilicon 1297 -1397 1297 -1397 0 1
rlabel polysilicon 1297 -1403 1297 -1403 0 3
rlabel polysilicon 1304 -1397 1304 -1397 0 1
rlabel polysilicon 1304 -1403 1304 -1403 0 3
rlabel polysilicon 1311 -1397 1311 -1397 0 1
rlabel polysilicon 1311 -1403 1311 -1403 0 3
rlabel polysilicon 1318 -1397 1318 -1397 0 1
rlabel polysilicon 1318 -1403 1318 -1403 0 3
rlabel polysilicon 1325 -1397 1325 -1397 0 1
rlabel polysilicon 1325 -1403 1325 -1403 0 3
rlabel polysilicon 1332 -1397 1332 -1397 0 1
rlabel polysilicon 1332 -1403 1332 -1403 0 3
rlabel polysilicon 1339 -1397 1339 -1397 0 1
rlabel polysilicon 1339 -1403 1339 -1403 0 3
rlabel polysilicon 1346 -1397 1346 -1397 0 1
rlabel polysilicon 1346 -1403 1346 -1403 0 3
rlabel polysilicon 1353 -1397 1353 -1397 0 1
rlabel polysilicon 1353 -1403 1353 -1403 0 3
rlabel polysilicon 1360 -1397 1360 -1397 0 1
rlabel polysilicon 1360 -1403 1360 -1403 0 3
rlabel polysilicon 1367 -1397 1367 -1397 0 1
rlabel polysilicon 1367 -1403 1367 -1403 0 3
rlabel polysilicon 1374 -1397 1374 -1397 0 1
rlabel polysilicon 1374 -1403 1374 -1403 0 3
rlabel polysilicon 1381 -1397 1381 -1397 0 1
rlabel polysilicon 1381 -1403 1381 -1403 0 3
rlabel polysilicon 1388 -1397 1388 -1397 0 1
rlabel polysilicon 1388 -1403 1388 -1403 0 3
rlabel polysilicon 1395 -1397 1395 -1397 0 1
rlabel polysilicon 1395 -1403 1395 -1403 0 3
rlabel polysilicon 1402 -1397 1402 -1397 0 1
rlabel polysilicon 1402 -1403 1402 -1403 0 3
rlabel polysilicon 1409 -1397 1409 -1397 0 1
rlabel polysilicon 1409 -1403 1409 -1403 0 3
rlabel polysilicon 1416 -1397 1416 -1397 0 1
rlabel polysilicon 1416 -1403 1416 -1403 0 3
rlabel polysilicon 1423 -1397 1423 -1397 0 1
rlabel polysilicon 1423 -1403 1423 -1403 0 3
rlabel polysilicon 1430 -1397 1430 -1397 0 1
rlabel polysilicon 1430 -1403 1430 -1403 0 3
rlabel polysilicon 1437 -1397 1437 -1397 0 1
rlabel polysilicon 1437 -1403 1437 -1403 0 3
rlabel polysilicon 1444 -1397 1444 -1397 0 1
rlabel polysilicon 1444 -1403 1444 -1403 0 3
rlabel polysilicon 1451 -1397 1451 -1397 0 1
rlabel polysilicon 1451 -1403 1451 -1403 0 3
rlabel polysilicon 1458 -1397 1458 -1397 0 1
rlabel polysilicon 1458 -1403 1458 -1403 0 3
rlabel polysilicon 1465 -1397 1465 -1397 0 1
rlabel polysilicon 1465 -1403 1465 -1403 0 3
rlabel polysilicon 1472 -1397 1472 -1397 0 1
rlabel polysilicon 1472 -1403 1472 -1403 0 3
rlabel polysilicon 1479 -1397 1479 -1397 0 1
rlabel polysilicon 1479 -1403 1479 -1403 0 3
rlabel polysilicon 1486 -1397 1486 -1397 0 1
rlabel polysilicon 1486 -1403 1486 -1403 0 3
rlabel polysilicon 1493 -1397 1493 -1397 0 1
rlabel polysilicon 1493 -1403 1493 -1403 0 3
rlabel polysilicon 1500 -1397 1500 -1397 0 1
rlabel polysilicon 1500 -1403 1500 -1403 0 3
rlabel polysilicon 1507 -1397 1507 -1397 0 1
rlabel polysilicon 1507 -1403 1507 -1403 0 3
rlabel polysilicon 1514 -1397 1514 -1397 0 1
rlabel polysilicon 1514 -1403 1514 -1403 0 3
rlabel polysilicon 1521 -1397 1521 -1397 0 1
rlabel polysilicon 1521 -1403 1521 -1403 0 3
rlabel polysilicon 1524 -1403 1524 -1403 0 4
rlabel polysilicon 1528 -1397 1528 -1397 0 1
rlabel polysilicon 1528 -1403 1528 -1403 0 3
rlabel polysilicon 1535 -1397 1535 -1397 0 1
rlabel polysilicon 1535 -1403 1535 -1403 0 3
rlabel polysilicon 2 -1530 2 -1530 0 1
rlabel polysilicon 2 -1536 2 -1536 0 3
rlabel polysilicon 9 -1530 9 -1530 0 1
rlabel polysilicon 9 -1536 9 -1536 0 3
rlabel polysilicon 16 -1530 16 -1530 0 1
rlabel polysilicon 16 -1536 16 -1536 0 3
rlabel polysilicon 23 -1530 23 -1530 0 1
rlabel polysilicon 23 -1536 23 -1536 0 3
rlabel polysilicon 30 -1530 30 -1530 0 1
rlabel polysilicon 30 -1536 30 -1536 0 3
rlabel polysilicon 37 -1530 37 -1530 0 1
rlabel polysilicon 37 -1536 37 -1536 0 3
rlabel polysilicon 44 -1530 44 -1530 0 1
rlabel polysilicon 44 -1536 44 -1536 0 3
rlabel polysilicon 51 -1530 51 -1530 0 1
rlabel polysilicon 54 -1530 54 -1530 0 2
rlabel polysilicon 51 -1536 51 -1536 0 3
rlabel polysilicon 54 -1536 54 -1536 0 4
rlabel polysilicon 58 -1530 58 -1530 0 1
rlabel polysilicon 58 -1536 58 -1536 0 3
rlabel polysilicon 65 -1530 65 -1530 0 1
rlabel polysilicon 65 -1536 65 -1536 0 3
rlabel polysilicon 72 -1530 72 -1530 0 1
rlabel polysilicon 72 -1536 72 -1536 0 3
rlabel polysilicon 79 -1530 79 -1530 0 1
rlabel polysilicon 82 -1530 82 -1530 0 2
rlabel polysilicon 82 -1536 82 -1536 0 4
rlabel polysilicon 86 -1530 86 -1530 0 1
rlabel polysilicon 86 -1536 86 -1536 0 3
rlabel polysilicon 93 -1530 93 -1530 0 1
rlabel polysilicon 93 -1536 93 -1536 0 3
rlabel polysilicon 100 -1530 100 -1530 0 1
rlabel polysilicon 103 -1530 103 -1530 0 2
rlabel polysilicon 100 -1536 100 -1536 0 3
rlabel polysilicon 103 -1536 103 -1536 0 4
rlabel polysilicon 107 -1530 107 -1530 0 1
rlabel polysilicon 107 -1536 107 -1536 0 3
rlabel polysilicon 114 -1530 114 -1530 0 1
rlabel polysilicon 114 -1536 114 -1536 0 3
rlabel polysilicon 121 -1530 121 -1530 0 1
rlabel polysilicon 121 -1536 121 -1536 0 3
rlabel polysilicon 128 -1530 128 -1530 0 1
rlabel polysilicon 128 -1536 128 -1536 0 3
rlabel polysilicon 135 -1530 135 -1530 0 1
rlabel polysilicon 135 -1536 135 -1536 0 3
rlabel polysilicon 142 -1530 142 -1530 0 1
rlabel polysilicon 142 -1536 142 -1536 0 3
rlabel polysilicon 149 -1530 149 -1530 0 1
rlabel polysilicon 149 -1536 149 -1536 0 3
rlabel polysilicon 156 -1530 156 -1530 0 1
rlabel polysilicon 156 -1536 156 -1536 0 3
rlabel polysilicon 163 -1530 163 -1530 0 1
rlabel polysilicon 163 -1536 163 -1536 0 3
rlabel polysilicon 173 -1530 173 -1530 0 2
rlabel polysilicon 170 -1536 170 -1536 0 3
rlabel polysilicon 173 -1536 173 -1536 0 4
rlabel polysilicon 177 -1530 177 -1530 0 1
rlabel polysilicon 177 -1536 177 -1536 0 3
rlabel polysilicon 184 -1530 184 -1530 0 1
rlabel polysilicon 184 -1536 184 -1536 0 3
rlabel polysilicon 191 -1530 191 -1530 0 1
rlabel polysilicon 191 -1536 191 -1536 0 3
rlabel polysilicon 198 -1530 198 -1530 0 1
rlabel polysilicon 198 -1536 198 -1536 0 3
rlabel polysilicon 205 -1530 205 -1530 0 1
rlabel polysilicon 205 -1536 205 -1536 0 3
rlabel polysilicon 212 -1530 212 -1530 0 1
rlabel polysilicon 212 -1536 212 -1536 0 3
rlabel polysilicon 219 -1530 219 -1530 0 1
rlabel polysilicon 219 -1536 219 -1536 0 3
rlabel polysilicon 226 -1530 226 -1530 0 1
rlabel polysilicon 226 -1536 226 -1536 0 3
rlabel polysilicon 233 -1530 233 -1530 0 1
rlabel polysilicon 233 -1536 233 -1536 0 3
rlabel polysilicon 240 -1530 240 -1530 0 1
rlabel polysilicon 240 -1536 240 -1536 0 3
rlabel polysilicon 247 -1530 247 -1530 0 1
rlabel polysilicon 247 -1536 247 -1536 0 3
rlabel polysilicon 254 -1530 254 -1530 0 1
rlabel polysilicon 254 -1536 254 -1536 0 3
rlabel polysilicon 261 -1530 261 -1530 0 1
rlabel polysilicon 261 -1536 261 -1536 0 3
rlabel polysilicon 268 -1530 268 -1530 0 1
rlabel polysilicon 268 -1536 268 -1536 0 3
rlabel polysilicon 275 -1530 275 -1530 0 1
rlabel polysilicon 275 -1536 275 -1536 0 3
rlabel polysilicon 282 -1530 282 -1530 0 1
rlabel polysilicon 282 -1536 282 -1536 0 3
rlabel polysilicon 289 -1530 289 -1530 0 1
rlabel polysilicon 289 -1536 289 -1536 0 3
rlabel polysilicon 296 -1530 296 -1530 0 1
rlabel polysilicon 296 -1536 296 -1536 0 3
rlabel polysilicon 303 -1530 303 -1530 0 1
rlabel polysilicon 303 -1536 303 -1536 0 3
rlabel polysilicon 310 -1530 310 -1530 0 1
rlabel polysilicon 310 -1536 310 -1536 0 3
rlabel polysilicon 317 -1530 317 -1530 0 1
rlabel polysilicon 317 -1536 317 -1536 0 3
rlabel polysilicon 324 -1530 324 -1530 0 1
rlabel polysilicon 324 -1536 324 -1536 0 3
rlabel polysilicon 331 -1530 331 -1530 0 1
rlabel polysilicon 331 -1536 331 -1536 0 3
rlabel polysilicon 338 -1530 338 -1530 0 1
rlabel polysilicon 338 -1536 338 -1536 0 3
rlabel polysilicon 345 -1530 345 -1530 0 1
rlabel polysilicon 345 -1536 345 -1536 0 3
rlabel polysilicon 352 -1530 352 -1530 0 1
rlabel polysilicon 352 -1536 352 -1536 0 3
rlabel polysilicon 359 -1530 359 -1530 0 1
rlabel polysilicon 359 -1536 359 -1536 0 3
rlabel polysilicon 366 -1530 366 -1530 0 1
rlabel polysilicon 366 -1536 366 -1536 0 3
rlabel polysilicon 373 -1530 373 -1530 0 1
rlabel polysilicon 373 -1536 373 -1536 0 3
rlabel polysilicon 380 -1530 380 -1530 0 1
rlabel polysilicon 380 -1536 380 -1536 0 3
rlabel polysilicon 387 -1530 387 -1530 0 1
rlabel polysilicon 387 -1536 387 -1536 0 3
rlabel polysilicon 394 -1530 394 -1530 0 1
rlabel polysilicon 397 -1530 397 -1530 0 2
rlabel polysilicon 394 -1536 394 -1536 0 3
rlabel polysilicon 397 -1536 397 -1536 0 4
rlabel polysilicon 401 -1530 401 -1530 0 1
rlabel polysilicon 401 -1536 401 -1536 0 3
rlabel polysilicon 408 -1530 408 -1530 0 1
rlabel polysilicon 408 -1536 408 -1536 0 3
rlabel polysilicon 415 -1530 415 -1530 0 1
rlabel polysilicon 415 -1536 415 -1536 0 3
rlabel polysilicon 422 -1530 422 -1530 0 1
rlabel polysilicon 422 -1536 422 -1536 0 3
rlabel polysilicon 429 -1530 429 -1530 0 1
rlabel polysilicon 432 -1530 432 -1530 0 2
rlabel polysilicon 432 -1536 432 -1536 0 4
rlabel polysilicon 436 -1530 436 -1530 0 1
rlabel polysilicon 436 -1536 436 -1536 0 3
rlabel polysilicon 443 -1530 443 -1530 0 1
rlabel polysilicon 443 -1536 443 -1536 0 3
rlabel polysilicon 450 -1530 450 -1530 0 1
rlabel polysilicon 450 -1536 450 -1536 0 3
rlabel polysilicon 457 -1530 457 -1530 0 1
rlabel polysilicon 457 -1536 457 -1536 0 3
rlabel polysilicon 464 -1530 464 -1530 0 1
rlabel polysilicon 464 -1536 464 -1536 0 3
rlabel polysilicon 471 -1530 471 -1530 0 1
rlabel polysilicon 474 -1530 474 -1530 0 2
rlabel polysilicon 471 -1536 471 -1536 0 3
rlabel polysilicon 474 -1536 474 -1536 0 4
rlabel polysilicon 478 -1530 478 -1530 0 1
rlabel polysilicon 478 -1536 478 -1536 0 3
rlabel polysilicon 485 -1530 485 -1530 0 1
rlabel polysilicon 485 -1536 485 -1536 0 3
rlabel polysilicon 492 -1530 492 -1530 0 1
rlabel polysilicon 492 -1536 492 -1536 0 3
rlabel polysilicon 499 -1530 499 -1530 0 1
rlabel polysilicon 502 -1530 502 -1530 0 2
rlabel polysilicon 499 -1536 499 -1536 0 3
rlabel polysilicon 502 -1536 502 -1536 0 4
rlabel polysilicon 506 -1530 506 -1530 0 1
rlabel polysilicon 506 -1536 506 -1536 0 3
rlabel polysilicon 513 -1530 513 -1530 0 1
rlabel polysilicon 513 -1536 513 -1536 0 3
rlabel polysilicon 520 -1530 520 -1530 0 1
rlabel polysilicon 520 -1536 520 -1536 0 3
rlabel polysilicon 527 -1530 527 -1530 0 1
rlabel polysilicon 527 -1536 527 -1536 0 3
rlabel polysilicon 534 -1530 534 -1530 0 1
rlabel polysilicon 534 -1536 534 -1536 0 3
rlabel polysilicon 541 -1530 541 -1530 0 1
rlabel polysilicon 541 -1536 541 -1536 0 3
rlabel polysilicon 548 -1530 548 -1530 0 1
rlabel polysilicon 548 -1536 548 -1536 0 3
rlabel polysilicon 555 -1530 555 -1530 0 1
rlabel polysilicon 555 -1536 555 -1536 0 3
rlabel polysilicon 562 -1530 562 -1530 0 1
rlabel polysilicon 562 -1536 562 -1536 0 3
rlabel polysilicon 569 -1530 569 -1530 0 1
rlabel polysilicon 569 -1536 569 -1536 0 3
rlabel polysilicon 576 -1530 576 -1530 0 1
rlabel polysilicon 579 -1530 579 -1530 0 2
rlabel polysilicon 576 -1536 576 -1536 0 3
rlabel polysilicon 579 -1536 579 -1536 0 4
rlabel polysilicon 583 -1530 583 -1530 0 1
rlabel polysilicon 583 -1536 583 -1536 0 3
rlabel polysilicon 590 -1530 590 -1530 0 1
rlabel polysilicon 590 -1536 590 -1536 0 3
rlabel polysilicon 597 -1530 597 -1530 0 1
rlabel polysilicon 600 -1530 600 -1530 0 2
rlabel polysilicon 600 -1536 600 -1536 0 4
rlabel polysilicon 604 -1530 604 -1530 0 1
rlabel polysilicon 604 -1536 604 -1536 0 3
rlabel polysilicon 611 -1530 611 -1530 0 1
rlabel polysilicon 611 -1536 611 -1536 0 3
rlabel polysilicon 618 -1530 618 -1530 0 1
rlabel polysilicon 618 -1536 618 -1536 0 3
rlabel polysilicon 625 -1530 625 -1530 0 1
rlabel polysilicon 625 -1536 625 -1536 0 3
rlabel polysilicon 632 -1530 632 -1530 0 1
rlabel polysilicon 632 -1536 632 -1536 0 3
rlabel polysilicon 639 -1530 639 -1530 0 1
rlabel polysilicon 639 -1536 639 -1536 0 3
rlabel polysilicon 646 -1530 646 -1530 0 1
rlabel polysilicon 646 -1536 646 -1536 0 3
rlabel polysilicon 653 -1530 653 -1530 0 1
rlabel polysilicon 653 -1536 653 -1536 0 3
rlabel polysilicon 660 -1530 660 -1530 0 1
rlabel polysilicon 660 -1536 660 -1536 0 3
rlabel polysilicon 667 -1530 667 -1530 0 1
rlabel polysilicon 667 -1536 667 -1536 0 3
rlabel polysilicon 674 -1530 674 -1530 0 1
rlabel polysilicon 677 -1530 677 -1530 0 2
rlabel polysilicon 674 -1536 674 -1536 0 3
rlabel polysilicon 677 -1536 677 -1536 0 4
rlabel polysilicon 681 -1530 681 -1530 0 1
rlabel polysilicon 684 -1530 684 -1530 0 2
rlabel polysilicon 681 -1536 681 -1536 0 3
rlabel polysilicon 684 -1536 684 -1536 0 4
rlabel polysilicon 688 -1530 688 -1530 0 1
rlabel polysilicon 688 -1536 688 -1536 0 3
rlabel polysilicon 695 -1530 695 -1530 0 1
rlabel polysilicon 695 -1536 695 -1536 0 3
rlabel polysilicon 702 -1530 702 -1530 0 1
rlabel polysilicon 702 -1536 702 -1536 0 3
rlabel polysilicon 709 -1530 709 -1530 0 1
rlabel polysilicon 709 -1536 709 -1536 0 3
rlabel polysilicon 716 -1530 716 -1530 0 1
rlabel polysilicon 716 -1536 716 -1536 0 3
rlabel polysilicon 723 -1530 723 -1530 0 1
rlabel polysilicon 726 -1530 726 -1530 0 2
rlabel polysilicon 723 -1536 723 -1536 0 3
rlabel polysilicon 726 -1536 726 -1536 0 4
rlabel polysilicon 730 -1530 730 -1530 0 1
rlabel polysilicon 730 -1536 730 -1536 0 3
rlabel polysilicon 737 -1530 737 -1530 0 1
rlabel polysilicon 737 -1536 737 -1536 0 3
rlabel polysilicon 744 -1530 744 -1530 0 1
rlabel polysilicon 744 -1536 744 -1536 0 3
rlabel polysilicon 751 -1530 751 -1530 0 1
rlabel polysilicon 751 -1536 751 -1536 0 3
rlabel polysilicon 758 -1530 758 -1530 0 1
rlabel polysilicon 758 -1536 758 -1536 0 3
rlabel polysilicon 765 -1530 765 -1530 0 1
rlabel polysilicon 768 -1530 768 -1530 0 2
rlabel polysilicon 765 -1536 765 -1536 0 3
rlabel polysilicon 768 -1536 768 -1536 0 4
rlabel polysilicon 772 -1530 772 -1530 0 1
rlabel polysilicon 772 -1536 772 -1536 0 3
rlabel polysilicon 779 -1530 779 -1530 0 1
rlabel polysilicon 779 -1536 779 -1536 0 3
rlabel polysilicon 786 -1530 786 -1530 0 1
rlabel polysilicon 786 -1536 786 -1536 0 3
rlabel polysilicon 793 -1530 793 -1530 0 1
rlabel polysilicon 793 -1536 793 -1536 0 3
rlabel polysilicon 800 -1530 800 -1530 0 1
rlabel polysilicon 803 -1530 803 -1530 0 2
rlabel polysilicon 800 -1536 800 -1536 0 3
rlabel polysilicon 803 -1536 803 -1536 0 4
rlabel polysilicon 807 -1530 807 -1530 0 1
rlabel polysilicon 807 -1536 807 -1536 0 3
rlabel polysilicon 814 -1530 814 -1530 0 1
rlabel polysilicon 817 -1530 817 -1530 0 2
rlabel polysilicon 814 -1536 814 -1536 0 3
rlabel polysilicon 817 -1536 817 -1536 0 4
rlabel polysilicon 821 -1530 821 -1530 0 1
rlabel polysilicon 821 -1536 821 -1536 0 3
rlabel polysilicon 828 -1530 828 -1530 0 1
rlabel polysilicon 831 -1530 831 -1530 0 2
rlabel polysilicon 828 -1536 828 -1536 0 3
rlabel polysilicon 831 -1536 831 -1536 0 4
rlabel polysilicon 835 -1530 835 -1530 0 1
rlabel polysilicon 838 -1530 838 -1530 0 2
rlabel polysilicon 835 -1536 835 -1536 0 3
rlabel polysilicon 838 -1536 838 -1536 0 4
rlabel polysilicon 842 -1530 842 -1530 0 1
rlabel polysilicon 842 -1536 842 -1536 0 3
rlabel polysilicon 849 -1530 849 -1530 0 1
rlabel polysilicon 849 -1536 849 -1536 0 3
rlabel polysilicon 856 -1530 856 -1530 0 1
rlabel polysilicon 859 -1530 859 -1530 0 2
rlabel polysilicon 859 -1536 859 -1536 0 4
rlabel polysilicon 863 -1530 863 -1530 0 1
rlabel polysilicon 863 -1536 863 -1536 0 3
rlabel polysilicon 870 -1530 870 -1530 0 1
rlabel polysilicon 870 -1536 870 -1536 0 3
rlabel polysilicon 877 -1530 877 -1530 0 1
rlabel polysilicon 880 -1530 880 -1530 0 2
rlabel polysilicon 877 -1536 877 -1536 0 3
rlabel polysilicon 884 -1530 884 -1530 0 1
rlabel polysilicon 884 -1536 884 -1536 0 3
rlabel polysilicon 891 -1530 891 -1530 0 1
rlabel polysilicon 891 -1536 891 -1536 0 3
rlabel polysilicon 898 -1530 898 -1530 0 1
rlabel polysilicon 898 -1536 898 -1536 0 3
rlabel polysilicon 905 -1530 905 -1530 0 1
rlabel polysilicon 905 -1536 905 -1536 0 3
rlabel polysilicon 912 -1530 912 -1530 0 1
rlabel polysilicon 912 -1536 912 -1536 0 3
rlabel polysilicon 919 -1530 919 -1530 0 1
rlabel polysilicon 919 -1536 919 -1536 0 3
rlabel polysilicon 926 -1530 926 -1530 0 1
rlabel polysilicon 926 -1536 926 -1536 0 3
rlabel polysilicon 933 -1530 933 -1530 0 1
rlabel polysilicon 933 -1536 933 -1536 0 3
rlabel polysilicon 940 -1530 940 -1530 0 1
rlabel polysilicon 940 -1536 940 -1536 0 3
rlabel polysilicon 947 -1530 947 -1530 0 1
rlabel polysilicon 947 -1536 947 -1536 0 3
rlabel polysilicon 954 -1530 954 -1530 0 1
rlabel polysilicon 954 -1536 954 -1536 0 3
rlabel polysilicon 961 -1530 961 -1530 0 1
rlabel polysilicon 961 -1536 961 -1536 0 3
rlabel polysilicon 968 -1530 968 -1530 0 1
rlabel polysilicon 968 -1536 968 -1536 0 3
rlabel polysilicon 975 -1530 975 -1530 0 1
rlabel polysilicon 975 -1536 975 -1536 0 3
rlabel polysilicon 982 -1530 982 -1530 0 1
rlabel polysilicon 982 -1536 982 -1536 0 3
rlabel polysilicon 989 -1530 989 -1530 0 1
rlabel polysilicon 992 -1530 992 -1530 0 2
rlabel polysilicon 989 -1536 989 -1536 0 3
rlabel polysilicon 992 -1536 992 -1536 0 4
rlabel polysilicon 999 -1530 999 -1530 0 2
rlabel polysilicon 996 -1536 996 -1536 0 3
rlabel polysilicon 999 -1536 999 -1536 0 4
rlabel polysilicon 1003 -1530 1003 -1530 0 1
rlabel polysilicon 1003 -1536 1003 -1536 0 3
rlabel polysilicon 1010 -1530 1010 -1530 0 1
rlabel polysilicon 1010 -1536 1010 -1536 0 3
rlabel polysilicon 1017 -1530 1017 -1530 0 1
rlabel polysilicon 1017 -1536 1017 -1536 0 3
rlabel polysilicon 1024 -1530 1024 -1530 0 1
rlabel polysilicon 1024 -1536 1024 -1536 0 3
rlabel polysilicon 1031 -1530 1031 -1530 0 1
rlabel polysilicon 1031 -1536 1031 -1536 0 3
rlabel polysilicon 1038 -1530 1038 -1530 0 1
rlabel polysilicon 1038 -1536 1038 -1536 0 3
rlabel polysilicon 1045 -1530 1045 -1530 0 1
rlabel polysilicon 1045 -1536 1045 -1536 0 3
rlabel polysilicon 1052 -1530 1052 -1530 0 1
rlabel polysilicon 1052 -1536 1052 -1536 0 3
rlabel polysilicon 1059 -1530 1059 -1530 0 1
rlabel polysilicon 1059 -1536 1059 -1536 0 3
rlabel polysilicon 1066 -1530 1066 -1530 0 1
rlabel polysilicon 1066 -1536 1066 -1536 0 3
rlabel polysilicon 1073 -1530 1073 -1530 0 1
rlabel polysilicon 1076 -1530 1076 -1530 0 2
rlabel polysilicon 1073 -1536 1073 -1536 0 3
rlabel polysilicon 1076 -1536 1076 -1536 0 4
rlabel polysilicon 1080 -1530 1080 -1530 0 1
rlabel polysilicon 1080 -1536 1080 -1536 0 3
rlabel polysilicon 1087 -1530 1087 -1530 0 1
rlabel polysilicon 1087 -1536 1087 -1536 0 3
rlabel polysilicon 1094 -1530 1094 -1530 0 1
rlabel polysilicon 1094 -1536 1094 -1536 0 3
rlabel polysilicon 1101 -1530 1101 -1530 0 1
rlabel polysilicon 1101 -1536 1101 -1536 0 3
rlabel polysilicon 1108 -1530 1108 -1530 0 1
rlabel polysilicon 1108 -1536 1108 -1536 0 3
rlabel polysilicon 1115 -1530 1115 -1530 0 1
rlabel polysilicon 1115 -1536 1115 -1536 0 3
rlabel polysilicon 1122 -1530 1122 -1530 0 1
rlabel polysilicon 1125 -1530 1125 -1530 0 2
rlabel polysilicon 1122 -1536 1122 -1536 0 3
rlabel polysilicon 1129 -1530 1129 -1530 0 1
rlabel polysilicon 1129 -1536 1129 -1536 0 3
rlabel polysilicon 1136 -1530 1136 -1530 0 1
rlabel polysilicon 1136 -1536 1136 -1536 0 3
rlabel polysilicon 1143 -1530 1143 -1530 0 1
rlabel polysilicon 1143 -1536 1143 -1536 0 3
rlabel polysilicon 1150 -1530 1150 -1530 0 1
rlabel polysilicon 1150 -1536 1150 -1536 0 3
rlabel polysilicon 1153 -1536 1153 -1536 0 4
rlabel polysilicon 1157 -1530 1157 -1530 0 1
rlabel polysilicon 1157 -1536 1157 -1536 0 3
rlabel polysilicon 1164 -1530 1164 -1530 0 1
rlabel polysilicon 1164 -1536 1164 -1536 0 3
rlabel polysilicon 1171 -1530 1171 -1530 0 1
rlabel polysilicon 1171 -1536 1171 -1536 0 3
rlabel polysilicon 1178 -1530 1178 -1530 0 1
rlabel polysilicon 1178 -1536 1178 -1536 0 3
rlabel polysilicon 1185 -1530 1185 -1530 0 1
rlabel polysilicon 1185 -1536 1185 -1536 0 3
rlabel polysilicon 1192 -1530 1192 -1530 0 1
rlabel polysilicon 1192 -1536 1192 -1536 0 3
rlabel polysilicon 1199 -1530 1199 -1530 0 1
rlabel polysilicon 1199 -1536 1199 -1536 0 3
rlabel polysilicon 1206 -1530 1206 -1530 0 1
rlabel polysilicon 1206 -1536 1206 -1536 0 3
rlabel polysilicon 1213 -1530 1213 -1530 0 1
rlabel polysilicon 1213 -1536 1213 -1536 0 3
rlabel polysilicon 1220 -1530 1220 -1530 0 1
rlabel polysilicon 1220 -1536 1220 -1536 0 3
rlabel polysilicon 1227 -1530 1227 -1530 0 1
rlabel polysilicon 1227 -1536 1227 -1536 0 3
rlabel polysilicon 1234 -1530 1234 -1530 0 1
rlabel polysilicon 1234 -1536 1234 -1536 0 3
rlabel polysilicon 1241 -1530 1241 -1530 0 1
rlabel polysilicon 1241 -1536 1241 -1536 0 3
rlabel polysilicon 1248 -1530 1248 -1530 0 1
rlabel polysilicon 1248 -1536 1248 -1536 0 3
rlabel polysilicon 1255 -1530 1255 -1530 0 1
rlabel polysilicon 1255 -1536 1255 -1536 0 3
rlabel polysilicon 1262 -1530 1262 -1530 0 1
rlabel polysilicon 1262 -1536 1262 -1536 0 3
rlabel polysilicon 1269 -1530 1269 -1530 0 1
rlabel polysilicon 1269 -1536 1269 -1536 0 3
rlabel polysilicon 1276 -1530 1276 -1530 0 1
rlabel polysilicon 1276 -1536 1276 -1536 0 3
rlabel polysilicon 1283 -1530 1283 -1530 0 1
rlabel polysilicon 1283 -1536 1283 -1536 0 3
rlabel polysilicon 1290 -1530 1290 -1530 0 1
rlabel polysilicon 1290 -1536 1290 -1536 0 3
rlabel polysilicon 1297 -1530 1297 -1530 0 1
rlabel polysilicon 1297 -1536 1297 -1536 0 3
rlabel polysilicon 1304 -1530 1304 -1530 0 1
rlabel polysilicon 1304 -1536 1304 -1536 0 3
rlabel polysilicon 1311 -1530 1311 -1530 0 1
rlabel polysilicon 1311 -1536 1311 -1536 0 3
rlabel polysilicon 1318 -1530 1318 -1530 0 1
rlabel polysilicon 1318 -1536 1318 -1536 0 3
rlabel polysilicon 1325 -1530 1325 -1530 0 1
rlabel polysilicon 1325 -1536 1325 -1536 0 3
rlabel polysilicon 1332 -1530 1332 -1530 0 1
rlabel polysilicon 1332 -1536 1332 -1536 0 3
rlabel polysilicon 1339 -1530 1339 -1530 0 1
rlabel polysilicon 1339 -1536 1339 -1536 0 3
rlabel polysilicon 1346 -1530 1346 -1530 0 1
rlabel polysilicon 1346 -1536 1346 -1536 0 3
rlabel polysilicon 1353 -1530 1353 -1530 0 1
rlabel polysilicon 1353 -1536 1353 -1536 0 3
rlabel polysilicon 1360 -1530 1360 -1530 0 1
rlabel polysilicon 1360 -1536 1360 -1536 0 3
rlabel polysilicon 1367 -1530 1367 -1530 0 1
rlabel polysilicon 1367 -1536 1367 -1536 0 3
rlabel polysilicon 1374 -1530 1374 -1530 0 1
rlabel polysilicon 1374 -1536 1374 -1536 0 3
rlabel polysilicon 1381 -1530 1381 -1530 0 1
rlabel polysilicon 1381 -1536 1381 -1536 0 3
rlabel polysilicon 1388 -1530 1388 -1530 0 1
rlabel polysilicon 1388 -1536 1388 -1536 0 3
rlabel polysilicon 1395 -1530 1395 -1530 0 1
rlabel polysilicon 1395 -1536 1395 -1536 0 3
rlabel polysilicon 1402 -1530 1402 -1530 0 1
rlabel polysilicon 1402 -1536 1402 -1536 0 3
rlabel polysilicon 1409 -1530 1409 -1530 0 1
rlabel polysilicon 1409 -1536 1409 -1536 0 3
rlabel polysilicon 1416 -1530 1416 -1530 0 1
rlabel polysilicon 1416 -1536 1416 -1536 0 3
rlabel polysilicon 1423 -1530 1423 -1530 0 1
rlabel polysilicon 1423 -1536 1423 -1536 0 3
rlabel polysilicon 1430 -1530 1430 -1530 0 1
rlabel polysilicon 1430 -1536 1430 -1536 0 3
rlabel polysilicon 1437 -1530 1437 -1530 0 1
rlabel polysilicon 1437 -1536 1437 -1536 0 3
rlabel polysilicon 1444 -1530 1444 -1530 0 1
rlabel polysilicon 1444 -1536 1444 -1536 0 3
rlabel polysilicon 1451 -1530 1451 -1530 0 1
rlabel polysilicon 1451 -1536 1451 -1536 0 3
rlabel polysilicon 1458 -1530 1458 -1530 0 1
rlabel polysilicon 1458 -1536 1458 -1536 0 3
rlabel polysilicon 1465 -1530 1465 -1530 0 1
rlabel polysilicon 1465 -1536 1465 -1536 0 3
rlabel polysilicon 1472 -1530 1472 -1530 0 1
rlabel polysilicon 1472 -1536 1472 -1536 0 3
rlabel polysilicon 1479 -1530 1479 -1530 0 1
rlabel polysilicon 1479 -1536 1479 -1536 0 3
rlabel polysilicon 1486 -1530 1486 -1530 0 1
rlabel polysilicon 1486 -1536 1486 -1536 0 3
rlabel polysilicon 1493 -1530 1493 -1530 0 1
rlabel polysilicon 1493 -1536 1493 -1536 0 3
rlabel polysilicon 1500 -1530 1500 -1530 0 1
rlabel polysilicon 1500 -1536 1500 -1536 0 3
rlabel polysilicon 1507 -1530 1507 -1530 0 1
rlabel polysilicon 1507 -1536 1507 -1536 0 3
rlabel polysilicon 1514 -1530 1514 -1530 0 1
rlabel polysilicon 1514 -1536 1514 -1536 0 3
rlabel polysilicon 1521 -1530 1521 -1530 0 1
rlabel polysilicon 1524 -1530 1524 -1530 0 2
rlabel polysilicon 1521 -1536 1521 -1536 0 3
rlabel polysilicon 1524 -1536 1524 -1536 0 4
rlabel polysilicon 1528 -1530 1528 -1530 0 1
rlabel polysilicon 1528 -1536 1528 -1536 0 3
rlabel polysilicon 1535 -1530 1535 -1530 0 1
rlabel polysilicon 1535 -1536 1535 -1536 0 3
rlabel polysilicon 2 -1637 2 -1637 0 1
rlabel polysilicon 2 -1643 2 -1643 0 3
rlabel polysilicon 9 -1637 9 -1637 0 1
rlabel polysilicon 9 -1643 9 -1643 0 3
rlabel polysilicon 16 -1637 16 -1637 0 1
rlabel polysilicon 16 -1643 16 -1643 0 3
rlabel polysilicon 23 -1637 23 -1637 0 1
rlabel polysilicon 23 -1643 23 -1643 0 3
rlabel polysilicon 30 -1637 30 -1637 0 1
rlabel polysilicon 30 -1643 30 -1643 0 3
rlabel polysilicon 37 -1637 37 -1637 0 1
rlabel polysilicon 37 -1643 37 -1643 0 3
rlabel polysilicon 44 -1637 44 -1637 0 1
rlabel polysilicon 44 -1643 44 -1643 0 3
rlabel polysilicon 51 -1637 51 -1637 0 1
rlabel polysilicon 51 -1643 51 -1643 0 3
rlabel polysilicon 58 -1637 58 -1637 0 1
rlabel polysilicon 58 -1643 58 -1643 0 3
rlabel polysilicon 65 -1637 65 -1637 0 1
rlabel polysilicon 65 -1643 65 -1643 0 3
rlabel polysilicon 72 -1637 72 -1637 0 1
rlabel polysilicon 75 -1637 75 -1637 0 2
rlabel polysilicon 72 -1643 72 -1643 0 3
rlabel polysilicon 75 -1643 75 -1643 0 4
rlabel polysilicon 79 -1637 79 -1637 0 1
rlabel polysilicon 79 -1643 79 -1643 0 3
rlabel polysilicon 86 -1637 86 -1637 0 1
rlabel polysilicon 86 -1643 86 -1643 0 3
rlabel polysilicon 93 -1637 93 -1637 0 1
rlabel polysilicon 93 -1643 93 -1643 0 3
rlabel polysilicon 100 -1637 100 -1637 0 1
rlabel polysilicon 100 -1643 100 -1643 0 3
rlabel polysilicon 107 -1637 107 -1637 0 1
rlabel polysilicon 107 -1643 107 -1643 0 3
rlabel polysilicon 110 -1643 110 -1643 0 4
rlabel polysilicon 114 -1637 114 -1637 0 1
rlabel polysilicon 114 -1643 114 -1643 0 3
rlabel polysilicon 121 -1637 121 -1637 0 1
rlabel polysilicon 121 -1643 121 -1643 0 3
rlabel polysilicon 128 -1637 128 -1637 0 1
rlabel polysilicon 131 -1637 131 -1637 0 2
rlabel polysilicon 128 -1643 128 -1643 0 3
rlabel polysilicon 131 -1643 131 -1643 0 4
rlabel polysilicon 135 -1637 135 -1637 0 1
rlabel polysilicon 135 -1643 135 -1643 0 3
rlabel polysilicon 142 -1637 142 -1637 0 1
rlabel polysilicon 145 -1637 145 -1637 0 2
rlabel polysilicon 142 -1643 142 -1643 0 3
rlabel polysilicon 145 -1643 145 -1643 0 4
rlabel polysilicon 149 -1637 149 -1637 0 1
rlabel polysilicon 149 -1643 149 -1643 0 3
rlabel polysilicon 156 -1637 156 -1637 0 1
rlabel polysilicon 156 -1643 156 -1643 0 3
rlabel polysilicon 163 -1637 163 -1637 0 1
rlabel polysilicon 163 -1643 163 -1643 0 3
rlabel polysilicon 170 -1637 170 -1637 0 1
rlabel polysilicon 170 -1643 170 -1643 0 3
rlabel polysilicon 177 -1637 177 -1637 0 1
rlabel polysilicon 177 -1643 177 -1643 0 3
rlabel polysilicon 184 -1637 184 -1637 0 1
rlabel polysilicon 184 -1643 184 -1643 0 3
rlabel polysilicon 191 -1637 191 -1637 0 1
rlabel polysilicon 191 -1643 191 -1643 0 3
rlabel polysilicon 198 -1637 198 -1637 0 1
rlabel polysilicon 198 -1643 198 -1643 0 3
rlabel polysilicon 205 -1637 205 -1637 0 1
rlabel polysilicon 205 -1643 205 -1643 0 3
rlabel polysilicon 212 -1637 212 -1637 0 1
rlabel polysilicon 212 -1643 212 -1643 0 3
rlabel polysilicon 219 -1637 219 -1637 0 1
rlabel polysilicon 219 -1643 219 -1643 0 3
rlabel polysilicon 226 -1637 226 -1637 0 1
rlabel polysilicon 226 -1643 226 -1643 0 3
rlabel polysilicon 233 -1637 233 -1637 0 1
rlabel polysilicon 233 -1643 233 -1643 0 3
rlabel polysilicon 240 -1637 240 -1637 0 1
rlabel polysilicon 240 -1643 240 -1643 0 3
rlabel polysilicon 247 -1637 247 -1637 0 1
rlabel polysilicon 247 -1643 247 -1643 0 3
rlabel polysilicon 254 -1637 254 -1637 0 1
rlabel polysilicon 254 -1643 254 -1643 0 3
rlabel polysilicon 261 -1637 261 -1637 0 1
rlabel polysilicon 261 -1643 261 -1643 0 3
rlabel polysilicon 268 -1637 268 -1637 0 1
rlabel polysilicon 271 -1637 271 -1637 0 2
rlabel polysilicon 268 -1643 268 -1643 0 3
rlabel polysilicon 271 -1643 271 -1643 0 4
rlabel polysilicon 275 -1637 275 -1637 0 1
rlabel polysilicon 275 -1643 275 -1643 0 3
rlabel polysilicon 282 -1637 282 -1637 0 1
rlabel polysilicon 282 -1643 282 -1643 0 3
rlabel polysilicon 289 -1637 289 -1637 0 1
rlabel polysilicon 289 -1643 289 -1643 0 3
rlabel polysilicon 296 -1637 296 -1637 0 1
rlabel polysilicon 296 -1643 296 -1643 0 3
rlabel polysilicon 303 -1637 303 -1637 0 1
rlabel polysilicon 303 -1643 303 -1643 0 3
rlabel polysilicon 310 -1637 310 -1637 0 1
rlabel polysilicon 310 -1643 310 -1643 0 3
rlabel polysilicon 317 -1637 317 -1637 0 1
rlabel polysilicon 317 -1643 317 -1643 0 3
rlabel polysilicon 324 -1637 324 -1637 0 1
rlabel polysilicon 324 -1643 324 -1643 0 3
rlabel polysilicon 331 -1637 331 -1637 0 1
rlabel polysilicon 331 -1643 331 -1643 0 3
rlabel polysilicon 338 -1637 338 -1637 0 1
rlabel polysilicon 338 -1643 338 -1643 0 3
rlabel polysilicon 348 -1637 348 -1637 0 2
rlabel polysilicon 345 -1643 345 -1643 0 3
rlabel polysilicon 352 -1637 352 -1637 0 1
rlabel polysilicon 352 -1643 352 -1643 0 3
rlabel polysilicon 359 -1637 359 -1637 0 1
rlabel polysilicon 359 -1643 359 -1643 0 3
rlabel polysilicon 366 -1637 366 -1637 0 1
rlabel polysilicon 369 -1637 369 -1637 0 2
rlabel polysilicon 366 -1643 366 -1643 0 3
rlabel polysilicon 369 -1643 369 -1643 0 4
rlabel polysilicon 373 -1637 373 -1637 0 1
rlabel polysilicon 373 -1643 373 -1643 0 3
rlabel polysilicon 380 -1637 380 -1637 0 1
rlabel polysilicon 380 -1643 380 -1643 0 3
rlabel polysilicon 387 -1637 387 -1637 0 1
rlabel polysilicon 387 -1643 387 -1643 0 3
rlabel polysilicon 394 -1637 394 -1637 0 1
rlabel polysilicon 394 -1643 394 -1643 0 3
rlabel polysilicon 401 -1637 401 -1637 0 1
rlabel polysilicon 401 -1643 401 -1643 0 3
rlabel polysilicon 408 -1637 408 -1637 0 1
rlabel polysilicon 408 -1643 408 -1643 0 3
rlabel polysilicon 415 -1637 415 -1637 0 1
rlabel polysilicon 415 -1643 415 -1643 0 3
rlabel polysilicon 422 -1637 422 -1637 0 1
rlabel polysilicon 422 -1643 422 -1643 0 3
rlabel polysilicon 429 -1637 429 -1637 0 1
rlabel polysilicon 429 -1643 429 -1643 0 3
rlabel polysilicon 439 -1637 439 -1637 0 2
rlabel polysilicon 436 -1643 436 -1643 0 3
rlabel polysilicon 443 -1637 443 -1637 0 1
rlabel polysilicon 446 -1637 446 -1637 0 2
rlabel polysilicon 446 -1643 446 -1643 0 4
rlabel polysilicon 450 -1637 450 -1637 0 1
rlabel polysilicon 450 -1643 450 -1643 0 3
rlabel polysilicon 457 -1637 457 -1637 0 1
rlabel polysilicon 457 -1643 457 -1643 0 3
rlabel polysilicon 464 -1637 464 -1637 0 1
rlabel polysilicon 464 -1643 464 -1643 0 3
rlabel polysilicon 471 -1637 471 -1637 0 1
rlabel polysilicon 474 -1637 474 -1637 0 2
rlabel polysilicon 471 -1643 471 -1643 0 3
rlabel polysilicon 474 -1643 474 -1643 0 4
rlabel polysilicon 478 -1637 478 -1637 0 1
rlabel polysilicon 478 -1643 478 -1643 0 3
rlabel polysilicon 485 -1637 485 -1637 0 1
rlabel polysilicon 485 -1643 485 -1643 0 3
rlabel polysilicon 492 -1637 492 -1637 0 1
rlabel polysilicon 492 -1643 492 -1643 0 3
rlabel polysilicon 499 -1637 499 -1637 0 1
rlabel polysilicon 502 -1637 502 -1637 0 2
rlabel polysilicon 499 -1643 499 -1643 0 3
rlabel polysilicon 502 -1643 502 -1643 0 4
rlabel polysilicon 506 -1637 506 -1637 0 1
rlabel polysilicon 506 -1643 506 -1643 0 3
rlabel polysilicon 513 -1637 513 -1637 0 1
rlabel polysilicon 513 -1643 513 -1643 0 3
rlabel polysilicon 520 -1637 520 -1637 0 1
rlabel polysilicon 520 -1643 520 -1643 0 3
rlabel polysilicon 527 -1637 527 -1637 0 1
rlabel polysilicon 527 -1643 527 -1643 0 3
rlabel polysilicon 534 -1637 534 -1637 0 1
rlabel polysilicon 534 -1643 534 -1643 0 3
rlabel polysilicon 541 -1637 541 -1637 0 1
rlabel polysilicon 541 -1643 541 -1643 0 3
rlabel polysilicon 548 -1637 548 -1637 0 1
rlabel polysilicon 548 -1643 548 -1643 0 3
rlabel polysilicon 555 -1637 555 -1637 0 1
rlabel polysilicon 558 -1637 558 -1637 0 2
rlabel polysilicon 555 -1643 555 -1643 0 3
rlabel polysilicon 562 -1637 562 -1637 0 1
rlabel polysilicon 565 -1637 565 -1637 0 2
rlabel polysilicon 562 -1643 562 -1643 0 3
rlabel polysilicon 565 -1643 565 -1643 0 4
rlabel polysilicon 569 -1637 569 -1637 0 1
rlabel polysilicon 569 -1643 569 -1643 0 3
rlabel polysilicon 576 -1637 576 -1637 0 1
rlabel polysilicon 576 -1643 576 -1643 0 3
rlabel polysilicon 583 -1637 583 -1637 0 1
rlabel polysilicon 583 -1643 583 -1643 0 3
rlabel polysilicon 590 -1637 590 -1637 0 1
rlabel polysilicon 590 -1643 590 -1643 0 3
rlabel polysilicon 597 -1643 597 -1643 0 3
rlabel polysilicon 604 -1637 604 -1637 0 1
rlabel polysilicon 604 -1643 604 -1643 0 3
rlabel polysilicon 611 -1637 611 -1637 0 1
rlabel polysilicon 611 -1643 611 -1643 0 3
rlabel polysilicon 618 -1637 618 -1637 0 1
rlabel polysilicon 621 -1637 621 -1637 0 2
rlabel polysilicon 618 -1643 618 -1643 0 3
rlabel polysilicon 621 -1643 621 -1643 0 4
rlabel polysilicon 625 -1637 625 -1637 0 1
rlabel polysilicon 625 -1643 625 -1643 0 3
rlabel polysilicon 632 -1637 632 -1637 0 1
rlabel polysilicon 632 -1643 632 -1643 0 3
rlabel polysilicon 639 -1637 639 -1637 0 1
rlabel polysilicon 639 -1643 639 -1643 0 3
rlabel polysilicon 646 -1637 646 -1637 0 1
rlabel polysilicon 649 -1637 649 -1637 0 2
rlabel polysilicon 646 -1643 646 -1643 0 3
rlabel polysilicon 649 -1643 649 -1643 0 4
rlabel polysilicon 653 -1637 653 -1637 0 1
rlabel polysilicon 653 -1643 653 -1643 0 3
rlabel polysilicon 660 -1637 660 -1637 0 1
rlabel polysilicon 660 -1643 660 -1643 0 3
rlabel polysilicon 667 -1637 667 -1637 0 1
rlabel polysilicon 667 -1643 667 -1643 0 3
rlabel polysilicon 674 -1637 674 -1637 0 1
rlabel polysilicon 674 -1643 674 -1643 0 3
rlabel polysilicon 681 -1637 681 -1637 0 1
rlabel polysilicon 681 -1643 681 -1643 0 3
rlabel polysilicon 688 -1637 688 -1637 0 1
rlabel polysilicon 688 -1643 688 -1643 0 3
rlabel polysilicon 695 -1637 695 -1637 0 1
rlabel polysilicon 695 -1643 695 -1643 0 3
rlabel polysilicon 702 -1637 702 -1637 0 1
rlabel polysilicon 702 -1643 702 -1643 0 3
rlabel polysilicon 709 -1637 709 -1637 0 1
rlabel polysilicon 709 -1643 709 -1643 0 3
rlabel polysilicon 716 -1637 716 -1637 0 1
rlabel polysilicon 716 -1643 716 -1643 0 3
rlabel polysilicon 723 -1637 723 -1637 0 1
rlabel polysilicon 723 -1643 723 -1643 0 3
rlabel polysilicon 730 -1637 730 -1637 0 1
rlabel polysilicon 730 -1643 730 -1643 0 3
rlabel polysilicon 737 -1637 737 -1637 0 1
rlabel polysilicon 740 -1637 740 -1637 0 2
rlabel polysilicon 737 -1643 737 -1643 0 3
rlabel polysilicon 740 -1643 740 -1643 0 4
rlabel polysilicon 744 -1637 744 -1637 0 1
rlabel polysilicon 744 -1643 744 -1643 0 3
rlabel polysilicon 751 -1637 751 -1637 0 1
rlabel polysilicon 754 -1637 754 -1637 0 2
rlabel polysilicon 751 -1643 751 -1643 0 3
rlabel polysilicon 754 -1643 754 -1643 0 4
rlabel polysilicon 758 -1637 758 -1637 0 1
rlabel polysilicon 758 -1643 758 -1643 0 3
rlabel polysilicon 765 -1637 765 -1637 0 1
rlabel polysilicon 765 -1643 765 -1643 0 3
rlabel polysilicon 772 -1637 772 -1637 0 1
rlabel polysilicon 772 -1643 772 -1643 0 3
rlabel polysilicon 779 -1637 779 -1637 0 1
rlabel polysilicon 782 -1637 782 -1637 0 2
rlabel polysilicon 779 -1643 779 -1643 0 3
rlabel polysilicon 782 -1643 782 -1643 0 4
rlabel polysilicon 786 -1637 786 -1637 0 1
rlabel polysilicon 786 -1643 786 -1643 0 3
rlabel polysilicon 793 -1637 793 -1637 0 1
rlabel polysilicon 793 -1643 793 -1643 0 3
rlabel polysilicon 800 -1637 800 -1637 0 1
rlabel polysilicon 800 -1643 800 -1643 0 3
rlabel polysilicon 807 -1637 807 -1637 0 1
rlabel polysilicon 807 -1643 807 -1643 0 3
rlabel polysilicon 814 -1637 814 -1637 0 1
rlabel polysilicon 817 -1637 817 -1637 0 2
rlabel polysilicon 817 -1643 817 -1643 0 4
rlabel polysilicon 821 -1637 821 -1637 0 1
rlabel polysilicon 821 -1643 821 -1643 0 3
rlabel polysilicon 828 -1637 828 -1637 0 1
rlabel polysilicon 831 -1637 831 -1637 0 2
rlabel polysilicon 828 -1643 828 -1643 0 3
rlabel polysilicon 831 -1643 831 -1643 0 4
rlabel polysilicon 835 -1637 835 -1637 0 1
rlabel polysilicon 835 -1643 835 -1643 0 3
rlabel polysilicon 842 -1637 842 -1637 0 1
rlabel polysilicon 842 -1643 842 -1643 0 3
rlabel polysilicon 849 -1637 849 -1637 0 1
rlabel polysilicon 849 -1643 849 -1643 0 3
rlabel polysilicon 856 -1637 856 -1637 0 1
rlabel polysilicon 856 -1643 856 -1643 0 3
rlabel polysilicon 863 -1637 863 -1637 0 1
rlabel polysilicon 863 -1643 863 -1643 0 3
rlabel polysilicon 870 -1637 870 -1637 0 1
rlabel polysilicon 870 -1643 870 -1643 0 3
rlabel polysilicon 877 -1637 877 -1637 0 1
rlabel polysilicon 880 -1637 880 -1637 0 2
rlabel polysilicon 877 -1643 877 -1643 0 3
rlabel polysilicon 880 -1643 880 -1643 0 4
rlabel polysilicon 884 -1637 884 -1637 0 1
rlabel polysilicon 884 -1643 884 -1643 0 3
rlabel polysilicon 891 -1637 891 -1637 0 1
rlabel polysilicon 891 -1643 891 -1643 0 3
rlabel polysilicon 898 -1637 898 -1637 0 1
rlabel polysilicon 898 -1643 898 -1643 0 3
rlabel polysilicon 905 -1637 905 -1637 0 1
rlabel polysilicon 905 -1643 905 -1643 0 3
rlabel polysilicon 912 -1637 912 -1637 0 1
rlabel polysilicon 912 -1643 912 -1643 0 3
rlabel polysilicon 919 -1637 919 -1637 0 1
rlabel polysilicon 919 -1643 919 -1643 0 3
rlabel polysilicon 926 -1637 926 -1637 0 1
rlabel polysilicon 926 -1643 926 -1643 0 3
rlabel polysilicon 933 -1637 933 -1637 0 1
rlabel polysilicon 933 -1643 933 -1643 0 3
rlabel polysilicon 940 -1637 940 -1637 0 1
rlabel polysilicon 940 -1643 940 -1643 0 3
rlabel polysilicon 947 -1637 947 -1637 0 1
rlabel polysilicon 947 -1643 947 -1643 0 3
rlabel polysilicon 954 -1637 954 -1637 0 1
rlabel polysilicon 957 -1637 957 -1637 0 2
rlabel polysilicon 954 -1643 954 -1643 0 3
rlabel polysilicon 961 -1637 961 -1637 0 1
rlabel polysilicon 961 -1643 961 -1643 0 3
rlabel polysilicon 968 -1637 968 -1637 0 1
rlabel polysilicon 968 -1643 968 -1643 0 3
rlabel polysilicon 975 -1637 975 -1637 0 1
rlabel polysilicon 975 -1643 975 -1643 0 3
rlabel polysilicon 982 -1637 982 -1637 0 1
rlabel polysilicon 982 -1643 982 -1643 0 3
rlabel polysilicon 989 -1637 989 -1637 0 1
rlabel polysilicon 992 -1637 992 -1637 0 2
rlabel polysilicon 992 -1643 992 -1643 0 4
rlabel polysilicon 996 -1637 996 -1637 0 1
rlabel polysilicon 996 -1643 996 -1643 0 3
rlabel polysilicon 1003 -1637 1003 -1637 0 1
rlabel polysilicon 1003 -1643 1003 -1643 0 3
rlabel polysilicon 1010 -1637 1010 -1637 0 1
rlabel polysilicon 1010 -1643 1010 -1643 0 3
rlabel polysilicon 1017 -1637 1017 -1637 0 1
rlabel polysilicon 1017 -1643 1017 -1643 0 3
rlabel polysilicon 1024 -1637 1024 -1637 0 1
rlabel polysilicon 1024 -1643 1024 -1643 0 3
rlabel polysilicon 1031 -1637 1031 -1637 0 1
rlabel polysilicon 1031 -1643 1031 -1643 0 3
rlabel polysilicon 1038 -1637 1038 -1637 0 1
rlabel polysilicon 1038 -1643 1038 -1643 0 3
rlabel polysilicon 1045 -1637 1045 -1637 0 1
rlabel polysilicon 1045 -1643 1045 -1643 0 3
rlabel polysilicon 1052 -1637 1052 -1637 0 1
rlabel polysilicon 1052 -1643 1052 -1643 0 3
rlabel polysilicon 1059 -1637 1059 -1637 0 1
rlabel polysilicon 1059 -1643 1059 -1643 0 3
rlabel polysilicon 1066 -1637 1066 -1637 0 1
rlabel polysilicon 1066 -1643 1066 -1643 0 3
rlabel polysilicon 1073 -1637 1073 -1637 0 1
rlabel polysilicon 1073 -1643 1073 -1643 0 3
rlabel polysilicon 1080 -1637 1080 -1637 0 1
rlabel polysilicon 1080 -1643 1080 -1643 0 3
rlabel polysilicon 1087 -1637 1087 -1637 0 1
rlabel polysilicon 1087 -1643 1087 -1643 0 3
rlabel polysilicon 1094 -1637 1094 -1637 0 1
rlabel polysilicon 1094 -1643 1094 -1643 0 3
rlabel polysilicon 1101 -1637 1101 -1637 0 1
rlabel polysilicon 1101 -1643 1101 -1643 0 3
rlabel polysilicon 1108 -1637 1108 -1637 0 1
rlabel polysilicon 1108 -1643 1108 -1643 0 3
rlabel polysilicon 1115 -1637 1115 -1637 0 1
rlabel polysilicon 1115 -1643 1115 -1643 0 3
rlabel polysilicon 1122 -1637 1122 -1637 0 1
rlabel polysilicon 1122 -1643 1122 -1643 0 3
rlabel polysilicon 1129 -1637 1129 -1637 0 1
rlabel polysilicon 1129 -1643 1129 -1643 0 3
rlabel polysilicon 1136 -1637 1136 -1637 0 1
rlabel polysilicon 1136 -1643 1136 -1643 0 3
rlabel polysilicon 1143 -1637 1143 -1637 0 1
rlabel polysilicon 1143 -1643 1143 -1643 0 3
rlabel polysilicon 1150 -1637 1150 -1637 0 1
rlabel polysilicon 1153 -1637 1153 -1637 0 2
rlabel polysilicon 1150 -1643 1150 -1643 0 3
rlabel polysilicon 1157 -1637 1157 -1637 0 1
rlabel polysilicon 1157 -1643 1157 -1643 0 3
rlabel polysilicon 1164 -1637 1164 -1637 0 1
rlabel polysilicon 1164 -1643 1164 -1643 0 3
rlabel polysilicon 1171 -1637 1171 -1637 0 1
rlabel polysilicon 1171 -1643 1171 -1643 0 3
rlabel polysilicon 1178 -1637 1178 -1637 0 1
rlabel polysilicon 1178 -1643 1178 -1643 0 3
rlabel polysilicon 1185 -1637 1185 -1637 0 1
rlabel polysilicon 1185 -1643 1185 -1643 0 3
rlabel polysilicon 1192 -1637 1192 -1637 0 1
rlabel polysilicon 1192 -1643 1192 -1643 0 3
rlabel polysilicon 1199 -1637 1199 -1637 0 1
rlabel polysilicon 1199 -1643 1199 -1643 0 3
rlabel polysilicon 1206 -1637 1206 -1637 0 1
rlabel polysilicon 1206 -1643 1206 -1643 0 3
rlabel polysilicon 1213 -1637 1213 -1637 0 1
rlabel polysilicon 1213 -1643 1213 -1643 0 3
rlabel polysilicon 1220 -1637 1220 -1637 0 1
rlabel polysilicon 1220 -1643 1220 -1643 0 3
rlabel polysilicon 1227 -1637 1227 -1637 0 1
rlabel polysilicon 1227 -1643 1227 -1643 0 3
rlabel polysilicon 1234 -1637 1234 -1637 0 1
rlabel polysilicon 1234 -1643 1234 -1643 0 3
rlabel polysilicon 1241 -1637 1241 -1637 0 1
rlabel polysilicon 1241 -1643 1241 -1643 0 3
rlabel polysilicon 1248 -1637 1248 -1637 0 1
rlabel polysilicon 1248 -1643 1248 -1643 0 3
rlabel polysilicon 1255 -1637 1255 -1637 0 1
rlabel polysilicon 1255 -1643 1255 -1643 0 3
rlabel polysilicon 1262 -1637 1262 -1637 0 1
rlabel polysilicon 1262 -1643 1262 -1643 0 3
rlabel polysilicon 1269 -1637 1269 -1637 0 1
rlabel polysilicon 1269 -1643 1269 -1643 0 3
rlabel polysilicon 1276 -1637 1276 -1637 0 1
rlabel polysilicon 1276 -1643 1276 -1643 0 3
rlabel polysilicon 1283 -1637 1283 -1637 0 1
rlabel polysilicon 1283 -1643 1283 -1643 0 3
rlabel polysilicon 1290 -1637 1290 -1637 0 1
rlabel polysilicon 1290 -1643 1290 -1643 0 3
rlabel polysilicon 1297 -1637 1297 -1637 0 1
rlabel polysilicon 1297 -1643 1297 -1643 0 3
rlabel polysilicon 1304 -1637 1304 -1637 0 1
rlabel polysilicon 1304 -1643 1304 -1643 0 3
rlabel polysilicon 1311 -1637 1311 -1637 0 1
rlabel polysilicon 1311 -1643 1311 -1643 0 3
rlabel polysilicon 1318 -1637 1318 -1637 0 1
rlabel polysilicon 1318 -1643 1318 -1643 0 3
rlabel polysilicon 1325 -1637 1325 -1637 0 1
rlabel polysilicon 1325 -1643 1325 -1643 0 3
rlabel polysilicon 1332 -1637 1332 -1637 0 1
rlabel polysilicon 1332 -1643 1332 -1643 0 3
rlabel polysilicon 1339 -1637 1339 -1637 0 1
rlabel polysilicon 1339 -1643 1339 -1643 0 3
rlabel polysilicon 1346 -1637 1346 -1637 0 1
rlabel polysilicon 1349 -1637 1349 -1637 0 2
rlabel polysilicon 1346 -1643 1346 -1643 0 3
rlabel polysilicon 1349 -1643 1349 -1643 0 4
rlabel polysilicon 1353 -1637 1353 -1637 0 1
rlabel polysilicon 1353 -1643 1353 -1643 0 3
rlabel polysilicon 1360 -1637 1360 -1637 0 1
rlabel polysilicon 1360 -1643 1360 -1643 0 3
rlabel polysilicon 1367 -1637 1367 -1637 0 1
rlabel polysilicon 1367 -1643 1367 -1643 0 3
rlabel polysilicon 1374 -1637 1374 -1637 0 1
rlabel polysilicon 1374 -1643 1374 -1643 0 3
rlabel polysilicon 1381 -1637 1381 -1637 0 1
rlabel polysilicon 1381 -1643 1381 -1643 0 3
rlabel polysilicon 1388 -1637 1388 -1637 0 1
rlabel polysilicon 1388 -1643 1388 -1643 0 3
rlabel polysilicon 1395 -1637 1395 -1637 0 1
rlabel polysilicon 1395 -1643 1395 -1643 0 3
rlabel polysilicon 1402 -1637 1402 -1637 0 1
rlabel polysilicon 1402 -1643 1402 -1643 0 3
rlabel polysilicon 1409 -1637 1409 -1637 0 1
rlabel polysilicon 1409 -1643 1409 -1643 0 3
rlabel polysilicon 1416 -1637 1416 -1637 0 1
rlabel polysilicon 1416 -1643 1416 -1643 0 3
rlabel polysilicon 1423 -1637 1423 -1637 0 1
rlabel polysilicon 1423 -1643 1423 -1643 0 3
rlabel polysilicon 1430 -1637 1430 -1637 0 1
rlabel polysilicon 1430 -1643 1430 -1643 0 3
rlabel polysilicon 1437 -1637 1437 -1637 0 1
rlabel polysilicon 1437 -1643 1437 -1643 0 3
rlabel polysilicon 1451 -1637 1451 -1637 0 1
rlabel polysilicon 1451 -1643 1451 -1643 0 3
rlabel polysilicon 9 -1762 9 -1762 0 1
rlabel polysilicon 9 -1768 9 -1768 0 3
rlabel polysilicon 16 -1762 16 -1762 0 1
rlabel polysilicon 16 -1768 16 -1768 0 3
rlabel polysilicon 23 -1762 23 -1762 0 1
rlabel polysilicon 23 -1768 23 -1768 0 3
rlabel polysilicon 30 -1762 30 -1762 0 1
rlabel polysilicon 30 -1768 30 -1768 0 3
rlabel polysilicon 37 -1762 37 -1762 0 1
rlabel polysilicon 37 -1768 37 -1768 0 3
rlabel polysilicon 44 -1762 44 -1762 0 1
rlabel polysilicon 44 -1768 44 -1768 0 3
rlabel polysilicon 51 -1762 51 -1762 0 1
rlabel polysilicon 51 -1768 51 -1768 0 3
rlabel polysilicon 58 -1762 58 -1762 0 1
rlabel polysilicon 58 -1768 58 -1768 0 3
rlabel polysilicon 65 -1762 65 -1762 0 1
rlabel polysilicon 65 -1768 65 -1768 0 3
rlabel polysilicon 72 -1762 72 -1762 0 1
rlabel polysilicon 75 -1762 75 -1762 0 2
rlabel polysilicon 72 -1768 72 -1768 0 3
rlabel polysilicon 75 -1768 75 -1768 0 4
rlabel polysilicon 79 -1762 79 -1762 0 1
rlabel polysilicon 82 -1762 82 -1762 0 2
rlabel polysilicon 79 -1768 79 -1768 0 3
rlabel polysilicon 82 -1768 82 -1768 0 4
rlabel polysilicon 86 -1762 86 -1762 0 1
rlabel polysilicon 86 -1768 86 -1768 0 3
rlabel polysilicon 93 -1762 93 -1762 0 1
rlabel polysilicon 93 -1768 93 -1768 0 3
rlabel polysilicon 100 -1762 100 -1762 0 1
rlabel polysilicon 100 -1768 100 -1768 0 3
rlabel polysilicon 107 -1762 107 -1762 0 1
rlabel polysilicon 110 -1762 110 -1762 0 2
rlabel polysilicon 107 -1768 107 -1768 0 3
rlabel polysilicon 114 -1762 114 -1762 0 1
rlabel polysilicon 114 -1768 114 -1768 0 3
rlabel polysilicon 121 -1762 121 -1762 0 1
rlabel polysilicon 121 -1768 121 -1768 0 3
rlabel polysilicon 128 -1762 128 -1762 0 1
rlabel polysilicon 128 -1768 128 -1768 0 3
rlabel polysilicon 135 -1762 135 -1762 0 1
rlabel polysilicon 135 -1768 135 -1768 0 3
rlabel polysilicon 142 -1762 142 -1762 0 1
rlabel polysilicon 142 -1768 142 -1768 0 3
rlabel polysilicon 149 -1762 149 -1762 0 1
rlabel polysilicon 149 -1768 149 -1768 0 3
rlabel polysilicon 156 -1762 156 -1762 0 1
rlabel polysilicon 156 -1768 156 -1768 0 3
rlabel polysilicon 163 -1762 163 -1762 0 1
rlabel polysilicon 163 -1768 163 -1768 0 3
rlabel polysilicon 170 -1762 170 -1762 0 1
rlabel polysilicon 170 -1768 170 -1768 0 3
rlabel polysilicon 177 -1762 177 -1762 0 1
rlabel polysilicon 177 -1768 177 -1768 0 3
rlabel polysilicon 184 -1762 184 -1762 0 1
rlabel polysilicon 184 -1768 184 -1768 0 3
rlabel polysilicon 191 -1762 191 -1762 0 1
rlabel polysilicon 191 -1768 191 -1768 0 3
rlabel polysilicon 198 -1762 198 -1762 0 1
rlabel polysilicon 198 -1768 198 -1768 0 3
rlabel polysilicon 205 -1762 205 -1762 0 1
rlabel polysilicon 205 -1768 205 -1768 0 3
rlabel polysilicon 212 -1762 212 -1762 0 1
rlabel polysilicon 212 -1768 212 -1768 0 3
rlabel polysilicon 219 -1762 219 -1762 0 1
rlabel polysilicon 219 -1768 219 -1768 0 3
rlabel polysilicon 226 -1762 226 -1762 0 1
rlabel polysilicon 226 -1768 226 -1768 0 3
rlabel polysilicon 233 -1762 233 -1762 0 1
rlabel polysilicon 233 -1768 233 -1768 0 3
rlabel polysilicon 240 -1762 240 -1762 0 1
rlabel polysilicon 240 -1768 240 -1768 0 3
rlabel polysilicon 247 -1762 247 -1762 0 1
rlabel polysilicon 247 -1768 247 -1768 0 3
rlabel polysilicon 254 -1762 254 -1762 0 1
rlabel polysilicon 254 -1768 254 -1768 0 3
rlabel polysilicon 261 -1762 261 -1762 0 1
rlabel polysilicon 261 -1768 261 -1768 0 3
rlabel polysilicon 268 -1762 268 -1762 0 1
rlabel polysilicon 268 -1768 268 -1768 0 3
rlabel polysilicon 275 -1762 275 -1762 0 1
rlabel polysilicon 275 -1768 275 -1768 0 3
rlabel polysilicon 282 -1762 282 -1762 0 1
rlabel polysilicon 282 -1768 282 -1768 0 3
rlabel polysilicon 289 -1762 289 -1762 0 1
rlabel polysilicon 289 -1768 289 -1768 0 3
rlabel polysilicon 296 -1762 296 -1762 0 1
rlabel polysilicon 296 -1768 296 -1768 0 3
rlabel polysilicon 303 -1762 303 -1762 0 1
rlabel polysilicon 303 -1768 303 -1768 0 3
rlabel polysilicon 310 -1762 310 -1762 0 1
rlabel polysilicon 310 -1768 310 -1768 0 3
rlabel polysilicon 317 -1762 317 -1762 0 1
rlabel polysilicon 317 -1768 317 -1768 0 3
rlabel polysilicon 324 -1762 324 -1762 0 1
rlabel polysilicon 324 -1768 324 -1768 0 3
rlabel polysilicon 331 -1762 331 -1762 0 1
rlabel polysilicon 331 -1768 331 -1768 0 3
rlabel polysilicon 338 -1762 338 -1762 0 1
rlabel polysilicon 341 -1762 341 -1762 0 2
rlabel polysilicon 338 -1768 338 -1768 0 3
rlabel polysilicon 341 -1768 341 -1768 0 4
rlabel polysilicon 345 -1762 345 -1762 0 1
rlabel polysilicon 345 -1768 345 -1768 0 3
rlabel polysilicon 352 -1762 352 -1762 0 1
rlabel polysilicon 352 -1768 352 -1768 0 3
rlabel polysilicon 359 -1762 359 -1762 0 1
rlabel polysilicon 359 -1768 359 -1768 0 3
rlabel polysilicon 366 -1762 366 -1762 0 1
rlabel polysilicon 369 -1762 369 -1762 0 2
rlabel polysilicon 366 -1768 366 -1768 0 3
rlabel polysilicon 369 -1768 369 -1768 0 4
rlabel polysilicon 373 -1762 373 -1762 0 1
rlabel polysilicon 373 -1768 373 -1768 0 3
rlabel polysilicon 380 -1762 380 -1762 0 1
rlabel polysilicon 380 -1768 380 -1768 0 3
rlabel polysilicon 387 -1762 387 -1762 0 1
rlabel polysilicon 387 -1768 387 -1768 0 3
rlabel polysilicon 394 -1762 394 -1762 0 1
rlabel polysilicon 394 -1768 394 -1768 0 3
rlabel polysilicon 401 -1762 401 -1762 0 1
rlabel polysilicon 401 -1768 401 -1768 0 3
rlabel polysilicon 408 -1762 408 -1762 0 1
rlabel polysilicon 408 -1768 408 -1768 0 3
rlabel polysilicon 415 -1762 415 -1762 0 1
rlabel polysilicon 418 -1762 418 -1762 0 2
rlabel polysilicon 415 -1768 415 -1768 0 3
rlabel polysilicon 418 -1768 418 -1768 0 4
rlabel polysilicon 422 -1762 422 -1762 0 1
rlabel polysilicon 425 -1762 425 -1762 0 2
rlabel polysilicon 422 -1768 422 -1768 0 3
rlabel polysilicon 429 -1762 429 -1762 0 1
rlabel polysilicon 429 -1768 429 -1768 0 3
rlabel polysilicon 436 -1762 436 -1762 0 1
rlabel polysilicon 436 -1768 436 -1768 0 3
rlabel polysilicon 443 -1762 443 -1762 0 1
rlabel polysilicon 443 -1768 443 -1768 0 3
rlabel polysilicon 450 -1762 450 -1762 0 1
rlabel polysilicon 450 -1768 450 -1768 0 3
rlabel polysilicon 457 -1762 457 -1762 0 1
rlabel polysilicon 464 -1762 464 -1762 0 1
rlabel polysilicon 464 -1768 464 -1768 0 3
rlabel polysilicon 471 -1762 471 -1762 0 1
rlabel polysilicon 471 -1768 471 -1768 0 3
rlabel polysilicon 478 -1762 478 -1762 0 1
rlabel polysilicon 478 -1768 478 -1768 0 3
rlabel polysilicon 488 -1762 488 -1762 0 2
rlabel polysilicon 485 -1768 485 -1768 0 3
rlabel polysilicon 488 -1768 488 -1768 0 4
rlabel polysilicon 492 -1762 492 -1762 0 1
rlabel polysilicon 492 -1768 492 -1768 0 3
rlabel polysilicon 499 -1762 499 -1762 0 1
rlabel polysilicon 499 -1768 499 -1768 0 3
rlabel polysilicon 506 -1762 506 -1762 0 1
rlabel polysilicon 509 -1762 509 -1762 0 2
rlabel polysilicon 506 -1768 506 -1768 0 3
rlabel polysilicon 509 -1768 509 -1768 0 4
rlabel polysilicon 513 -1762 513 -1762 0 1
rlabel polysilicon 513 -1768 513 -1768 0 3
rlabel polysilicon 520 -1762 520 -1762 0 1
rlabel polysilicon 523 -1762 523 -1762 0 2
rlabel polysilicon 527 -1762 527 -1762 0 1
rlabel polysilicon 530 -1762 530 -1762 0 2
rlabel polysilicon 527 -1768 527 -1768 0 3
rlabel polysilicon 530 -1768 530 -1768 0 4
rlabel polysilicon 534 -1762 534 -1762 0 1
rlabel polysilicon 534 -1768 534 -1768 0 3
rlabel polysilicon 541 -1762 541 -1762 0 1
rlabel polysilicon 541 -1768 541 -1768 0 3
rlabel polysilicon 548 -1762 548 -1762 0 1
rlabel polysilicon 548 -1768 548 -1768 0 3
rlabel polysilicon 555 -1762 555 -1762 0 1
rlabel polysilicon 555 -1768 555 -1768 0 3
rlabel polysilicon 562 -1762 562 -1762 0 1
rlabel polysilicon 562 -1768 562 -1768 0 3
rlabel polysilicon 569 -1762 569 -1762 0 1
rlabel polysilicon 569 -1768 569 -1768 0 3
rlabel polysilicon 576 -1762 576 -1762 0 1
rlabel polysilicon 576 -1768 576 -1768 0 3
rlabel polysilicon 583 -1762 583 -1762 0 1
rlabel polysilicon 586 -1762 586 -1762 0 2
rlabel polysilicon 583 -1768 583 -1768 0 3
rlabel polysilicon 586 -1768 586 -1768 0 4
rlabel polysilicon 590 -1762 590 -1762 0 1
rlabel polysilicon 590 -1768 590 -1768 0 3
rlabel polysilicon 597 -1762 597 -1762 0 1
rlabel polysilicon 597 -1768 597 -1768 0 3
rlabel polysilicon 604 -1762 604 -1762 0 1
rlabel polysilicon 604 -1768 604 -1768 0 3
rlabel polysilicon 611 -1762 611 -1762 0 1
rlabel polysilicon 611 -1768 611 -1768 0 3
rlabel polysilicon 618 -1762 618 -1762 0 1
rlabel polysilicon 618 -1768 618 -1768 0 3
rlabel polysilicon 625 -1762 625 -1762 0 1
rlabel polysilicon 625 -1768 625 -1768 0 3
rlabel polysilicon 632 -1762 632 -1762 0 1
rlabel polysilicon 635 -1762 635 -1762 0 2
rlabel polysilicon 632 -1768 632 -1768 0 3
rlabel polysilicon 635 -1768 635 -1768 0 4
rlabel polysilicon 639 -1762 639 -1762 0 1
rlabel polysilicon 639 -1768 639 -1768 0 3
rlabel polysilicon 646 -1762 646 -1762 0 1
rlabel polysilicon 646 -1768 646 -1768 0 3
rlabel polysilicon 653 -1762 653 -1762 0 1
rlabel polysilicon 653 -1768 653 -1768 0 3
rlabel polysilicon 660 -1762 660 -1762 0 1
rlabel polysilicon 660 -1768 660 -1768 0 3
rlabel polysilicon 667 -1762 667 -1762 0 1
rlabel polysilicon 667 -1768 667 -1768 0 3
rlabel polysilicon 674 -1762 674 -1762 0 1
rlabel polysilicon 674 -1768 674 -1768 0 3
rlabel polysilicon 681 -1762 681 -1762 0 1
rlabel polysilicon 681 -1768 681 -1768 0 3
rlabel polysilicon 688 -1762 688 -1762 0 1
rlabel polysilicon 688 -1768 688 -1768 0 3
rlabel polysilicon 695 -1762 695 -1762 0 1
rlabel polysilicon 695 -1768 695 -1768 0 3
rlabel polysilicon 702 -1762 702 -1762 0 1
rlabel polysilicon 702 -1768 702 -1768 0 3
rlabel polysilicon 709 -1762 709 -1762 0 1
rlabel polysilicon 709 -1768 709 -1768 0 3
rlabel polysilicon 716 -1762 716 -1762 0 1
rlabel polysilicon 719 -1762 719 -1762 0 2
rlabel polysilicon 716 -1768 716 -1768 0 3
rlabel polysilicon 719 -1768 719 -1768 0 4
rlabel polysilicon 723 -1762 723 -1762 0 1
rlabel polysilicon 723 -1768 723 -1768 0 3
rlabel polysilicon 730 -1762 730 -1762 0 1
rlabel polysilicon 730 -1768 730 -1768 0 3
rlabel polysilicon 737 -1762 737 -1762 0 1
rlabel polysilicon 737 -1768 737 -1768 0 3
rlabel polysilicon 744 -1762 744 -1762 0 1
rlabel polysilicon 744 -1768 744 -1768 0 3
rlabel polysilicon 751 -1762 751 -1762 0 1
rlabel polysilicon 751 -1768 751 -1768 0 3
rlabel polysilicon 758 -1762 758 -1762 0 1
rlabel polysilicon 758 -1768 758 -1768 0 3
rlabel polysilicon 765 -1762 765 -1762 0 1
rlabel polysilicon 765 -1768 765 -1768 0 3
rlabel polysilicon 772 -1762 772 -1762 0 1
rlabel polysilicon 775 -1762 775 -1762 0 2
rlabel polysilicon 772 -1768 772 -1768 0 3
rlabel polysilicon 775 -1768 775 -1768 0 4
rlabel polysilicon 779 -1762 779 -1762 0 1
rlabel polysilicon 779 -1768 779 -1768 0 3
rlabel polysilicon 786 -1762 786 -1762 0 1
rlabel polysilicon 786 -1768 786 -1768 0 3
rlabel polysilicon 793 -1762 793 -1762 0 1
rlabel polysilicon 796 -1762 796 -1762 0 2
rlabel polysilicon 793 -1768 793 -1768 0 3
rlabel polysilicon 796 -1768 796 -1768 0 4
rlabel polysilicon 800 -1762 800 -1762 0 1
rlabel polysilicon 800 -1768 800 -1768 0 3
rlabel polysilicon 810 -1762 810 -1762 0 2
rlabel polysilicon 807 -1768 807 -1768 0 3
rlabel polysilicon 810 -1768 810 -1768 0 4
rlabel polysilicon 814 -1762 814 -1762 0 1
rlabel polysilicon 814 -1768 814 -1768 0 3
rlabel polysilicon 821 -1762 821 -1762 0 1
rlabel polysilicon 821 -1768 821 -1768 0 3
rlabel polysilicon 828 -1762 828 -1762 0 1
rlabel polysilicon 828 -1768 828 -1768 0 3
rlabel polysilicon 835 -1762 835 -1762 0 1
rlabel polysilicon 835 -1768 835 -1768 0 3
rlabel polysilicon 842 -1762 842 -1762 0 1
rlabel polysilicon 845 -1762 845 -1762 0 2
rlabel polysilicon 842 -1768 842 -1768 0 3
rlabel polysilicon 845 -1768 845 -1768 0 4
rlabel polysilicon 849 -1762 849 -1762 0 1
rlabel polysilicon 849 -1768 849 -1768 0 3
rlabel polysilicon 856 -1762 856 -1762 0 1
rlabel polysilicon 856 -1768 856 -1768 0 3
rlabel polysilicon 863 -1762 863 -1762 0 1
rlabel polysilicon 863 -1768 863 -1768 0 3
rlabel polysilicon 870 -1762 870 -1762 0 1
rlabel polysilicon 873 -1762 873 -1762 0 2
rlabel polysilicon 870 -1768 870 -1768 0 3
rlabel polysilicon 873 -1768 873 -1768 0 4
rlabel polysilicon 877 -1762 877 -1762 0 1
rlabel polysilicon 880 -1762 880 -1762 0 2
rlabel polysilicon 877 -1768 877 -1768 0 3
rlabel polysilicon 880 -1768 880 -1768 0 4
rlabel polysilicon 884 -1762 884 -1762 0 1
rlabel polysilicon 884 -1768 884 -1768 0 3
rlabel polysilicon 891 -1762 891 -1762 0 1
rlabel polysilicon 891 -1768 891 -1768 0 3
rlabel polysilicon 898 -1762 898 -1762 0 1
rlabel polysilicon 901 -1762 901 -1762 0 2
rlabel polysilicon 898 -1768 898 -1768 0 3
rlabel polysilicon 901 -1768 901 -1768 0 4
rlabel polysilicon 905 -1762 905 -1762 0 1
rlabel polysilicon 905 -1768 905 -1768 0 3
rlabel polysilicon 912 -1762 912 -1762 0 1
rlabel polysilicon 912 -1768 912 -1768 0 3
rlabel polysilicon 919 -1762 919 -1762 0 1
rlabel polysilicon 919 -1768 919 -1768 0 3
rlabel polysilicon 926 -1762 926 -1762 0 1
rlabel polysilicon 926 -1768 926 -1768 0 3
rlabel polysilicon 933 -1762 933 -1762 0 1
rlabel polysilicon 933 -1768 933 -1768 0 3
rlabel polysilicon 940 -1762 940 -1762 0 1
rlabel polysilicon 940 -1768 940 -1768 0 3
rlabel polysilicon 947 -1762 947 -1762 0 1
rlabel polysilicon 947 -1768 947 -1768 0 3
rlabel polysilicon 954 -1762 954 -1762 0 1
rlabel polysilicon 954 -1768 954 -1768 0 3
rlabel polysilicon 961 -1762 961 -1762 0 1
rlabel polysilicon 961 -1768 961 -1768 0 3
rlabel polysilicon 968 -1762 968 -1762 0 1
rlabel polysilicon 968 -1768 968 -1768 0 3
rlabel polysilicon 975 -1762 975 -1762 0 1
rlabel polysilicon 975 -1768 975 -1768 0 3
rlabel polysilicon 982 -1762 982 -1762 0 1
rlabel polysilicon 982 -1768 982 -1768 0 3
rlabel polysilicon 989 -1762 989 -1762 0 1
rlabel polysilicon 992 -1762 992 -1762 0 2
rlabel polysilicon 989 -1768 989 -1768 0 3
rlabel polysilicon 996 -1762 996 -1762 0 1
rlabel polysilicon 996 -1768 996 -1768 0 3
rlabel polysilicon 1003 -1762 1003 -1762 0 1
rlabel polysilicon 1006 -1762 1006 -1762 0 2
rlabel polysilicon 1003 -1768 1003 -1768 0 3
rlabel polysilicon 1006 -1768 1006 -1768 0 4
rlabel polysilicon 1010 -1762 1010 -1762 0 1
rlabel polysilicon 1010 -1768 1010 -1768 0 3
rlabel polysilicon 1017 -1762 1017 -1762 0 1
rlabel polysilicon 1017 -1768 1017 -1768 0 3
rlabel polysilicon 1024 -1762 1024 -1762 0 1
rlabel polysilicon 1024 -1768 1024 -1768 0 3
rlabel polysilicon 1031 -1762 1031 -1762 0 1
rlabel polysilicon 1031 -1768 1031 -1768 0 3
rlabel polysilicon 1038 -1762 1038 -1762 0 1
rlabel polysilicon 1038 -1768 1038 -1768 0 3
rlabel polysilicon 1045 -1762 1045 -1762 0 1
rlabel polysilicon 1045 -1768 1045 -1768 0 3
rlabel polysilicon 1052 -1762 1052 -1762 0 1
rlabel polysilicon 1052 -1768 1052 -1768 0 3
rlabel polysilicon 1059 -1762 1059 -1762 0 1
rlabel polysilicon 1059 -1768 1059 -1768 0 3
rlabel polysilicon 1066 -1762 1066 -1762 0 1
rlabel polysilicon 1066 -1768 1066 -1768 0 3
rlabel polysilicon 1073 -1762 1073 -1762 0 1
rlabel polysilicon 1073 -1768 1073 -1768 0 3
rlabel polysilicon 1080 -1762 1080 -1762 0 1
rlabel polysilicon 1080 -1768 1080 -1768 0 3
rlabel polysilicon 1087 -1762 1087 -1762 0 1
rlabel polysilicon 1087 -1768 1087 -1768 0 3
rlabel polysilicon 1094 -1762 1094 -1762 0 1
rlabel polysilicon 1094 -1768 1094 -1768 0 3
rlabel polysilicon 1101 -1762 1101 -1762 0 1
rlabel polysilicon 1101 -1768 1101 -1768 0 3
rlabel polysilicon 1108 -1762 1108 -1762 0 1
rlabel polysilicon 1108 -1768 1108 -1768 0 3
rlabel polysilicon 1115 -1762 1115 -1762 0 1
rlabel polysilicon 1115 -1768 1115 -1768 0 3
rlabel polysilicon 1122 -1762 1122 -1762 0 1
rlabel polysilicon 1122 -1768 1122 -1768 0 3
rlabel polysilicon 1129 -1762 1129 -1762 0 1
rlabel polysilicon 1129 -1768 1129 -1768 0 3
rlabel polysilicon 1136 -1762 1136 -1762 0 1
rlabel polysilicon 1136 -1768 1136 -1768 0 3
rlabel polysilicon 1143 -1762 1143 -1762 0 1
rlabel polysilicon 1143 -1768 1143 -1768 0 3
rlabel polysilicon 1150 -1762 1150 -1762 0 1
rlabel polysilicon 1150 -1768 1150 -1768 0 3
rlabel polysilicon 1157 -1762 1157 -1762 0 1
rlabel polysilicon 1157 -1768 1157 -1768 0 3
rlabel polysilicon 1164 -1762 1164 -1762 0 1
rlabel polysilicon 1164 -1768 1164 -1768 0 3
rlabel polysilicon 1171 -1762 1171 -1762 0 1
rlabel polysilicon 1171 -1768 1171 -1768 0 3
rlabel polysilicon 1178 -1762 1178 -1762 0 1
rlabel polysilicon 1178 -1768 1178 -1768 0 3
rlabel polysilicon 1185 -1762 1185 -1762 0 1
rlabel polysilicon 1185 -1768 1185 -1768 0 3
rlabel polysilicon 1192 -1762 1192 -1762 0 1
rlabel polysilicon 1192 -1768 1192 -1768 0 3
rlabel polysilicon 1199 -1762 1199 -1762 0 1
rlabel polysilicon 1199 -1768 1199 -1768 0 3
rlabel polysilicon 1206 -1762 1206 -1762 0 1
rlabel polysilicon 1206 -1768 1206 -1768 0 3
rlabel polysilicon 1213 -1762 1213 -1762 0 1
rlabel polysilicon 1213 -1768 1213 -1768 0 3
rlabel polysilicon 1220 -1762 1220 -1762 0 1
rlabel polysilicon 1220 -1768 1220 -1768 0 3
rlabel polysilicon 1227 -1762 1227 -1762 0 1
rlabel polysilicon 1227 -1768 1227 -1768 0 3
rlabel polysilicon 1234 -1762 1234 -1762 0 1
rlabel polysilicon 1234 -1768 1234 -1768 0 3
rlabel polysilicon 1241 -1762 1241 -1762 0 1
rlabel polysilicon 1241 -1768 1241 -1768 0 3
rlabel polysilicon 1248 -1762 1248 -1762 0 1
rlabel polysilicon 1248 -1768 1248 -1768 0 3
rlabel polysilicon 1255 -1762 1255 -1762 0 1
rlabel polysilicon 1255 -1768 1255 -1768 0 3
rlabel polysilicon 1258 -1768 1258 -1768 0 4
rlabel polysilicon 1262 -1762 1262 -1762 0 1
rlabel polysilicon 1262 -1768 1262 -1768 0 3
rlabel polysilicon 1269 -1762 1269 -1762 0 1
rlabel polysilicon 1269 -1768 1269 -1768 0 3
rlabel polysilicon 1276 -1762 1276 -1762 0 1
rlabel polysilicon 1276 -1768 1276 -1768 0 3
rlabel polysilicon 1283 -1762 1283 -1762 0 1
rlabel polysilicon 1283 -1768 1283 -1768 0 3
rlabel polysilicon 1290 -1762 1290 -1762 0 1
rlabel polysilicon 1290 -1768 1290 -1768 0 3
rlabel polysilicon 1297 -1762 1297 -1762 0 1
rlabel polysilicon 1297 -1768 1297 -1768 0 3
rlabel polysilicon 1304 -1762 1304 -1762 0 1
rlabel polysilicon 1304 -1768 1304 -1768 0 3
rlabel polysilicon 1311 -1762 1311 -1762 0 1
rlabel polysilicon 1311 -1768 1311 -1768 0 3
rlabel polysilicon 1318 -1762 1318 -1762 0 1
rlabel polysilicon 1318 -1768 1318 -1768 0 3
rlabel polysilicon 1325 -1762 1325 -1762 0 1
rlabel polysilicon 1325 -1768 1325 -1768 0 3
rlabel polysilicon 1332 -1762 1332 -1762 0 1
rlabel polysilicon 1332 -1768 1332 -1768 0 3
rlabel polysilicon 1339 -1762 1339 -1762 0 1
rlabel polysilicon 1339 -1768 1339 -1768 0 3
rlabel polysilicon 1346 -1762 1346 -1762 0 1
rlabel polysilicon 1346 -1768 1346 -1768 0 3
rlabel polysilicon 1353 -1762 1353 -1762 0 1
rlabel polysilicon 1353 -1768 1353 -1768 0 3
rlabel polysilicon 1360 -1762 1360 -1762 0 1
rlabel polysilicon 1360 -1768 1360 -1768 0 3
rlabel polysilicon 1367 -1762 1367 -1762 0 1
rlabel polysilicon 1370 -1762 1370 -1762 0 2
rlabel polysilicon 1367 -1768 1367 -1768 0 3
rlabel polysilicon 1370 -1768 1370 -1768 0 4
rlabel polysilicon 1374 -1762 1374 -1762 0 1
rlabel polysilicon 1377 -1762 1377 -1762 0 2
rlabel polysilicon 1374 -1768 1374 -1768 0 3
rlabel polysilicon 1377 -1768 1377 -1768 0 4
rlabel polysilicon 1381 -1762 1381 -1762 0 1
rlabel polysilicon 1381 -1768 1381 -1768 0 3
rlabel polysilicon 1388 -1762 1388 -1762 0 1
rlabel polysilicon 1388 -1768 1388 -1768 0 3
rlabel polysilicon 1395 -1762 1395 -1762 0 1
rlabel polysilicon 1395 -1768 1395 -1768 0 3
rlabel polysilicon 1402 -1762 1402 -1762 0 1
rlabel polysilicon 1402 -1768 1402 -1768 0 3
rlabel polysilicon 1409 -1762 1409 -1762 0 1
rlabel polysilicon 1409 -1768 1409 -1768 0 3
rlabel polysilicon 1416 -1762 1416 -1762 0 1
rlabel polysilicon 1416 -1768 1416 -1768 0 3
rlabel polysilicon 1423 -1762 1423 -1762 0 1
rlabel polysilicon 1423 -1768 1423 -1768 0 3
rlabel polysilicon 2 -1859 2 -1859 0 1
rlabel polysilicon 2 -1865 2 -1865 0 3
rlabel polysilicon 9 -1859 9 -1859 0 1
rlabel polysilicon 9 -1865 9 -1865 0 3
rlabel polysilicon 19 -1859 19 -1859 0 2
rlabel polysilicon 16 -1865 16 -1865 0 3
rlabel polysilicon 19 -1865 19 -1865 0 4
rlabel polysilicon 23 -1859 23 -1859 0 1
rlabel polysilicon 23 -1865 23 -1865 0 3
rlabel polysilicon 30 -1859 30 -1859 0 1
rlabel polysilicon 30 -1865 30 -1865 0 3
rlabel polysilicon 37 -1859 37 -1859 0 1
rlabel polysilicon 37 -1865 37 -1865 0 3
rlabel polysilicon 44 -1859 44 -1859 0 1
rlabel polysilicon 44 -1865 44 -1865 0 3
rlabel polysilicon 51 -1859 51 -1859 0 1
rlabel polysilicon 51 -1865 51 -1865 0 3
rlabel polysilicon 58 -1859 58 -1859 0 1
rlabel polysilicon 61 -1859 61 -1859 0 2
rlabel polysilicon 58 -1865 58 -1865 0 3
rlabel polysilicon 61 -1865 61 -1865 0 4
rlabel polysilicon 65 -1859 65 -1859 0 1
rlabel polysilicon 65 -1865 65 -1865 0 3
rlabel polysilicon 72 -1859 72 -1859 0 1
rlabel polysilicon 72 -1865 72 -1865 0 3
rlabel polysilicon 79 -1859 79 -1859 0 1
rlabel polysilicon 79 -1865 79 -1865 0 3
rlabel polysilicon 86 -1859 86 -1859 0 1
rlabel polysilicon 89 -1859 89 -1859 0 2
rlabel polysilicon 86 -1865 86 -1865 0 3
rlabel polysilicon 89 -1865 89 -1865 0 4
rlabel polysilicon 93 -1859 93 -1859 0 1
rlabel polysilicon 93 -1865 93 -1865 0 3
rlabel polysilicon 100 -1859 100 -1859 0 1
rlabel polysilicon 100 -1865 100 -1865 0 3
rlabel polysilicon 107 -1859 107 -1859 0 1
rlabel polysilicon 107 -1865 107 -1865 0 3
rlabel polysilicon 114 -1859 114 -1859 0 1
rlabel polysilicon 114 -1865 114 -1865 0 3
rlabel polysilicon 121 -1859 121 -1859 0 1
rlabel polysilicon 121 -1865 121 -1865 0 3
rlabel polysilicon 128 -1859 128 -1859 0 1
rlabel polysilicon 128 -1865 128 -1865 0 3
rlabel polysilicon 135 -1859 135 -1859 0 1
rlabel polysilicon 138 -1859 138 -1859 0 2
rlabel polysilicon 135 -1865 135 -1865 0 3
rlabel polysilicon 138 -1865 138 -1865 0 4
rlabel polysilicon 142 -1859 142 -1859 0 1
rlabel polysilicon 142 -1865 142 -1865 0 3
rlabel polysilicon 149 -1859 149 -1859 0 1
rlabel polysilicon 149 -1865 149 -1865 0 3
rlabel polysilicon 156 -1859 156 -1859 0 1
rlabel polysilicon 156 -1865 156 -1865 0 3
rlabel polysilicon 163 -1859 163 -1859 0 1
rlabel polysilicon 163 -1865 163 -1865 0 3
rlabel polysilicon 170 -1859 170 -1859 0 1
rlabel polysilicon 170 -1865 170 -1865 0 3
rlabel polysilicon 177 -1859 177 -1859 0 1
rlabel polysilicon 177 -1865 177 -1865 0 3
rlabel polysilicon 184 -1859 184 -1859 0 1
rlabel polysilicon 184 -1865 184 -1865 0 3
rlabel polysilicon 191 -1859 191 -1859 0 1
rlabel polysilicon 191 -1865 191 -1865 0 3
rlabel polysilicon 198 -1859 198 -1859 0 1
rlabel polysilicon 198 -1865 198 -1865 0 3
rlabel polysilicon 205 -1859 205 -1859 0 1
rlabel polysilicon 205 -1865 205 -1865 0 3
rlabel polysilicon 212 -1859 212 -1859 0 1
rlabel polysilicon 212 -1865 212 -1865 0 3
rlabel polysilicon 219 -1859 219 -1859 0 1
rlabel polysilicon 219 -1865 219 -1865 0 3
rlabel polysilicon 226 -1859 226 -1859 0 1
rlabel polysilicon 226 -1865 226 -1865 0 3
rlabel polysilicon 233 -1859 233 -1859 0 1
rlabel polysilicon 233 -1865 233 -1865 0 3
rlabel polysilicon 240 -1859 240 -1859 0 1
rlabel polysilicon 240 -1865 240 -1865 0 3
rlabel polysilicon 247 -1859 247 -1859 0 1
rlabel polysilicon 247 -1865 247 -1865 0 3
rlabel polysilicon 254 -1859 254 -1859 0 1
rlabel polysilicon 254 -1865 254 -1865 0 3
rlabel polysilicon 261 -1859 261 -1859 0 1
rlabel polysilicon 261 -1865 261 -1865 0 3
rlabel polysilicon 268 -1859 268 -1859 0 1
rlabel polysilicon 268 -1865 268 -1865 0 3
rlabel polysilicon 275 -1859 275 -1859 0 1
rlabel polysilicon 275 -1865 275 -1865 0 3
rlabel polysilicon 282 -1859 282 -1859 0 1
rlabel polysilicon 282 -1865 282 -1865 0 3
rlabel polysilicon 289 -1859 289 -1859 0 1
rlabel polysilicon 289 -1865 289 -1865 0 3
rlabel polysilicon 296 -1859 296 -1859 0 1
rlabel polysilicon 299 -1859 299 -1859 0 2
rlabel polysilicon 296 -1865 296 -1865 0 3
rlabel polysilicon 299 -1865 299 -1865 0 4
rlabel polysilicon 303 -1859 303 -1859 0 1
rlabel polysilicon 303 -1865 303 -1865 0 3
rlabel polysilicon 310 -1859 310 -1859 0 1
rlabel polysilicon 310 -1865 310 -1865 0 3
rlabel polysilicon 317 -1859 317 -1859 0 1
rlabel polysilicon 317 -1865 317 -1865 0 3
rlabel polysilicon 324 -1859 324 -1859 0 1
rlabel polysilicon 324 -1865 324 -1865 0 3
rlabel polysilicon 331 -1859 331 -1859 0 1
rlabel polysilicon 331 -1865 331 -1865 0 3
rlabel polysilicon 338 -1859 338 -1859 0 1
rlabel polysilicon 338 -1865 338 -1865 0 3
rlabel polysilicon 345 -1859 345 -1859 0 1
rlabel polysilicon 345 -1865 345 -1865 0 3
rlabel polysilicon 348 -1865 348 -1865 0 4
rlabel polysilicon 352 -1859 352 -1859 0 1
rlabel polysilicon 352 -1865 352 -1865 0 3
rlabel polysilicon 359 -1859 359 -1859 0 1
rlabel polysilicon 359 -1865 359 -1865 0 3
rlabel polysilicon 366 -1859 366 -1859 0 1
rlabel polysilicon 366 -1865 366 -1865 0 3
rlabel polysilicon 373 -1859 373 -1859 0 1
rlabel polysilicon 373 -1865 373 -1865 0 3
rlabel polysilicon 380 -1859 380 -1859 0 1
rlabel polysilicon 380 -1865 380 -1865 0 3
rlabel polysilicon 387 -1859 387 -1859 0 1
rlabel polysilicon 387 -1865 387 -1865 0 3
rlabel polysilicon 394 -1859 394 -1859 0 1
rlabel polysilicon 397 -1859 397 -1859 0 2
rlabel polysilicon 394 -1865 394 -1865 0 3
rlabel polysilicon 397 -1865 397 -1865 0 4
rlabel polysilicon 401 -1859 401 -1859 0 1
rlabel polysilicon 401 -1865 401 -1865 0 3
rlabel polysilicon 408 -1859 408 -1859 0 1
rlabel polysilicon 408 -1865 408 -1865 0 3
rlabel polysilicon 415 -1859 415 -1859 0 1
rlabel polysilicon 415 -1865 415 -1865 0 3
rlabel polysilicon 422 -1859 422 -1859 0 1
rlabel polysilicon 422 -1865 422 -1865 0 3
rlabel polysilicon 432 -1859 432 -1859 0 2
rlabel polysilicon 429 -1865 429 -1865 0 3
rlabel polysilicon 432 -1865 432 -1865 0 4
rlabel polysilicon 436 -1859 436 -1859 0 1
rlabel polysilicon 436 -1865 436 -1865 0 3
rlabel polysilicon 443 -1859 443 -1859 0 1
rlabel polysilicon 443 -1865 443 -1865 0 3
rlabel polysilicon 450 -1859 450 -1859 0 1
rlabel polysilicon 450 -1865 450 -1865 0 3
rlabel polysilicon 457 -1865 457 -1865 0 3
rlabel polysilicon 464 -1859 464 -1859 0 1
rlabel polysilicon 464 -1865 464 -1865 0 3
rlabel polysilicon 471 -1859 471 -1859 0 1
rlabel polysilicon 471 -1865 471 -1865 0 3
rlabel polysilicon 478 -1859 478 -1859 0 1
rlabel polysilicon 478 -1865 478 -1865 0 3
rlabel polysilicon 485 -1859 485 -1859 0 1
rlabel polysilicon 485 -1865 485 -1865 0 3
rlabel polysilicon 492 -1859 492 -1859 0 1
rlabel polysilicon 492 -1865 492 -1865 0 3
rlabel polysilicon 499 -1859 499 -1859 0 1
rlabel polysilicon 502 -1859 502 -1859 0 2
rlabel polysilicon 499 -1865 499 -1865 0 3
rlabel polysilicon 502 -1865 502 -1865 0 4
rlabel polysilicon 506 -1859 506 -1859 0 1
rlabel polysilicon 506 -1865 506 -1865 0 3
rlabel polysilicon 513 -1859 513 -1859 0 1
rlabel polysilicon 513 -1865 513 -1865 0 3
rlabel polysilicon 520 -1859 520 -1859 0 1
rlabel polysilicon 520 -1865 520 -1865 0 3
rlabel polysilicon 527 -1859 527 -1859 0 1
rlabel polysilicon 527 -1865 527 -1865 0 3
rlabel polysilicon 534 -1859 534 -1859 0 1
rlabel polysilicon 534 -1865 534 -1865 0 3
rlabel polysilicon 541 -1859 541 -1859 0 1
rlabel polysilicon 541 -1865 541 -1865 0 3
rlabel polysilicon 548 -1859 548 -1859 0 1
rlabel polysilicon 548 -1865 548 -1865 0 3
rlabel polysilicon 555 -1859 555 -1859 0 1
rlabel polysilicon 558 -1859 558 -1859 0 2
rlabel polysilicon 558 -1865 558 -1865 0 4
rlabel polysilicon 562 -1859 562 -1859 0 1
rlabel polysilicon 562 -1865 562 -1865 0 3
rlabel polysilicon 569 -1859 569 -1859 0 1
rlabel polysilicon 572 -1859 572 -1859 0 2
rlabel polysilicon 569 -1865 569 -1865 0 3
rlabel polysilicon 572 -1865 572 -1865 0 4
rlabel polysilicon 576 -1859 576 -1859 0 1
rlabel polysilicon 576 -1865 576 -1865 0 3
rlabel polysilicon 583 -1859 583 -1859 0 1
rlabel polysilicon 583 -1865 583 -1865 0 3
rlabel polysilicon 590 -1859 590 -1859 0 1
rlabel polysilicon 593 -1859 593 -1859 0 2
rlabel polysilicon 590 -1865 590 -1865 0 3
rlabel polysilicon 593 -1865 593 -1865 0 4
rlabel polysilicon 597 -1859 597 -1859 0 1
rlabel polysilicon 597 -1865 597 -1865 0 3
rlabel polysilicon 604 -1859 604 -1859 0 1
rlabel polysilicon 604 -1865 604 -1865 0 3
rlabel polysilicon 611 -1859 611 -1859 0 1
rlabel polysilicon 611 -1865 611 -1865 0 3
rlabel polysilicon 618 -1859 618 -1859 0 1
rlabel polysilicon 618 -1865 618 -1865 0 3
rlabel polysilicon 625 -1859 625 -1859 0 1
rlabel polysilicon 625 -1865 625 -1865 0 3
rlabel polysilicon 632 -1859 632 -1859 0 1
rlabel polysilicon 632 -1865 632 -1865 0 3
rlabel polysilicon 639 -1859 639 -1859 0 1
rlabel polysilicon 639 -1865 639 -1865 0 3
rlabel polysilicon 646 -1859 646 -1859 0 1
rlabel polysilicon 646 -1865 646 -1865 0 3
rlabel polysilicon 653 -1859 653 -1859 0 1
rlabel polysilicon 653 -1865 653 -1865 0 3
rlabel polysilicon 660 -1859 660 -1859 0 1
rlabel polysilicon 663 -1859 663 -1859 0 2
rlabel polysilicon 660 -1865 660 -1865 0 3
rlabel polysilicon 663 -1865 663 -1865 0 4
rlabel polysilicon 667 -1859 667 -1859 0 1
rlabel polysilicon 667 -1865 667 -1865 0 3
rlabel polysilicon 674 -1859 674 -1859 0 1
rlabel polysilicon 674 -1865 674 -1865 0 3
rlabel polysilicon 681 -1859 681 -1859 0 1
rlabel polysilicon 684 -1859 684 -1859 0 2
rlabel polysilicon 681 -1865 681 -1865 0 3
rlabel polysilicon 684 -1865 684 -1865 0 4
rlabel polysilicon 688 -1859 688 -1859 0 1
rlabel polysilicon 691 -1859 691 -1859 0 2
rlabel polysilicon 688 -1865 688 -1865 0 3
rlabel polysilicon 691 -1865 691 -1865 0 4
rlabel polysilicon 695 -1859 695 -1859 0 1
rlabel polysilicon 695 -1865 695 -1865 0 3
rlabel polysilicon 702 -1859 702 -1859 0 1
rlabel polysilicon 702 -1865 702 -1865 0 3
rlabel polysilicon 709 -1859 709 -1859 0 1
rlabel polysilicon 709 -1865 709 -1865 0 3
rlabel polysilicon 716 -1859 716 -1859 0 1
rlabel polysilicon 719 -1859 719 -1859 0 2
rlabel polysilicon 716 -1865 716 -1865 0 3
rlabel polysilicon 719 -1865 719 -1865 0 4
rlabel polysilicon 723 -1859 723 -1859 0 1
rlabel polysilicon 723 -1865 723 -1865 0 3
rlabel polysilicon 730 -1859 730 -1859 0 1
rlabel polysilicon 730 -1865 730 -1865 0 3
rlabel polysilicon 737 -1859 737 -1859 0 1
rlabel polysilicon 737 -1865 737 -1865 0 3
rlabel polysilicon 744 -1859 744 -1859 0 1
rlabel polysilicon 744 -1865 744 -1865 0 3
rlabel polysilicon 751 -1859 751 -1859 0 1
rlabel polysilicon 754 -1859 754 -1859 0 2
rlabel polysilicon 751 -1865 751 -1865 0 3
rlabel polysilicon 754 -1865 754 -1865 0 4
rlabel polysilicon 758 -1859 758 -1859 0 1
rlabel polysilicon 758 -1865 758 -1865 0 3
rlabel polysilicon 765 -1859 765 -1859 0 1
rlabel polysilicon 765 -1865 765 -1865 0 3
rlabel polysilicon 772 -1859 772 -1859 0 1
rlabel polysilicon 772 -1865 772 -1865 0 3
rlabel polysilicon 775 -1865 775 -1865 0 4
rlabel polysilicon 779 -1859 779 -1859 0 1
rlabel polysilicon 779 -1865 779 -1865 0 3
rlabel polysilicon 786 -1859 786 -1859 0 1
rlabel polysilicon 786 -1865 786 -1865 0 3
rlabel polysilicon 793 -1859 793 -1859 0 1
rlabel polysilicon 793 -1865 793 -1865 0 3
rlabel polysilicon 800 -1859 800 -1859 0 1
rlabel polysilicon 803 -1859 803 -1859 0 2
rlabel polysilicon 800 -1865 800 -1865 0 3
rlabel polysilicon 803 -1865 803 -1865 0 4
rlabel polysilicon 807 -1859 807 -1859 0 1
rlabel polysilicon 807 -1865 807 -1865 0 3
rlabel polysilicon 814 -1859 814 -1859 0 1
rlabel polysilicon 814 -1865 814 -1865 0 3
rlabel polysilicon 821 -1859 821 -1859 0 1
rlabel polysilicon 821 -1865 821 -1865 0 3
rlabel polysilicon 828 -1859 828 -1859 0 1
rlabel polysilicon 828 -1865 828 -1865 0 3
rlabel polysilicon 835 -1859 835 -1859 0 1
rlabel polysilicon 835 -1865 835 -1865 0 3
rlabel polysilicon 842 -1859 842 -1859 0 1
rlabel polysilicon 842 -1865 842 -1865 0 3
rlabel polysilicon 849 -1859 849 -1859 0 1
rlabel polysilicon 849 -1865 849 -1865 0 3
rlabel polysilicon 856 -1859 856 -1859 0 1
rlabel polysilicon 856 -1865 856 -1865 0 3
rlabel polysilicon 863 -1859 863 -1859 0 1
rlabel polysilicon 863 -1865 863 -1865 0 3
rlabel polysilicon 870 -1859 870 -1859 0 1
rlabel polysilicon 870 -1865 870 -1865 0 3
rlabel polysilicon 877 -1859 877 -1859 0 1
rlabel polysilicon 877 -1865 877 -1865 0 3
rlabel polysilicon 884 -1859 884 -1859 0 1
rlabel polysilicon 887 -1859 887 -1859 0 2
rlabel polysilicon 884 -1865 884 -1865 0 3
rlabel polysilicon 887 -1865 887 -1865 0 4
rlabel polysilicon 891 -1859 891 -1859 0 1
rlabel polysilicon 891 -1865 891 -1865 0 3
rlabel polysilicon 898 -1859 898 -1859 0 1
rlabel polysilicon 898 -1865 898 -1865 0 3
rlabel polysilicon 905 -1859 905 -1859 0 1
rlabel polysilicon 908 -1859 908 -1859 0 2
rlabel polysilicon 908 -1865 908 -1865 0 4
rlabel polysilicon 912 -1859 912 -1859 0 1
rlabel polysilicon 912 -1865 912 -1865 0 3
rlabel polysilicon 919 -1859 919 -1859 0 1
rlabel polysilicon 919 -1865 919 -1865 0 3
rlabel polysilicon 926 -1859 926 -1859 0 1
rlabel polysilicon 926 -1865 926 -1865 0 3
rlabel polysilicon 933 -1859 933 -1859 0 1
rlabel polysilicon 936 -1859 936 -1859 0 2
rlabel polysilicon 933 -1865 933 -1865 0 3
rlabel polysilicon 936 -1865 936 -1865 0 4
rlabel polysilicon 940 -1859 940 -1859 0 1
rlabel polysilicon 940 -1865 940 -1865 0 3
rlabel polysilicon 947 -1859 947 -1859 0 1
rlabel polysilicon 947 -1865 947 -1865 0 3
rlabel polysilicon 954 -1859 954 -1859 0 1
rlabel polysilicon 954 -1865 954 -1865 0 3
rlabel polysilicon 961 -1859 961 -1859 0 1
rlabel polysilicon 961 -1865 961 -1865 0 3
rlabel polysilicon 968 -1859 968 -1859 0 1
rlabel polysilicon 968 -1865 968 -1865 0 3
rlabel polysilicon 975 -1859 975 -1859 0 1
rlabel polysilicon 975 -1865 975 -1865 0 3
rlabel polysilicon 982 -1859 982 -1859 0 1
rlabel polysilicon 982 -1865 982 -1865 0 3
rlabel polysilicon 989 -1859 989 -1859 0 1
rlabel polysilicon 989 -1865 989 -1865 0 3
rlabel polysilicon 996 -1859 996 -1859 0 1
rlabel polysilicon 996 -1865 996 -1865 0 3
rlabel polysilicon 1003 -1859 1003 -1859 0 1
rlabel polysilicon 1003 -1865 1003 -1865 0 3
rlabel polysilicon 1010 -1859 1010 -1859 0 1
rlabel polysilicon 1010 -1865 1010 -1865 0 3
rlabel polysilicon 1017 -1859 1017 -1859 0 1
rlabel polysilicon 1017 -1865 1017 -1865 0 3
rlabel polysilicon 1024 -1859 1024 -1859 0 1
rlabel polysilicon 1024 -1865 1024 -1865 0 3
rlabel polysilicon 1031 -1859 1031 -1859 0 1
rlabel polysilicon 1031 -1865 1031 -1865 0 3
rlabel polysilicon 1038 -1859 1038 -1859 0 1
rlabel polysilicon 1038 -1865 1038 -1865 0 3
rlabel polysilicon 1045 -1859 1045 -1859 0 1
rlabel polysilicon 1045 -1865 1045 -1865 0 3
rlabel polysilicon 1052 -1859 1052 -1859 0 1
rlabel polysilicon 1052 -1865 1052 -1865 0 3
rlabel polysilicon 1062 -1859 1062 -1859 0 2
rlabel polysilicon 1059 -1865 1059 -1865 0 3
rlabel polysilicon 1062 -1865 1062 -1865 0 4
rlabel polysilicon 1066 -1859 1066 -1859 0 1
rlabel polysilicon 1066 -1865 1066 -1865 0 3
rlabel polysilicon 1073 -1859 1073 -1859 0 1
rlabel polysilicon 1073 -1865 1073 -1865 0 3
rlabel polysilicon 1080 -1859 1080 -1859 0 1
rlabel polysilicon 1080 -1865 1080 -1865 0 3
rlabel polysilicon 1087 -1859 1087 -1859 0 1
rlabel polysilicon 1087 -1865 1087 -1865 0 3
rlabel polysilicon 1094 -1859 1094 -1859 0 1
rlabel polysilicon 1094 -1865 1094 -1865 0 3
rlabel polysilicon 1101 -1859 1101 -1859 0 1
rlabel polysilicon 1101 -1865 1101 -1865 0 3
rlabel polysilicon 1108 -1859 1108 -1859 0 1
rlabel polysilicon 1108 -1865 1108 -1865 0 3
rlabel polysilicon 1115 -1859 1115 -1859 0 1
rlabel polysilicon 1115 -1865 1115 -1865 0 3
rlabel polysilicon 1122 -1859 1122 -1859 0 1
rlabel polysilicon 1122 -1865 1122 -1865 0 3
rlabel polysilicon 1129 -1859 1129 -1859 0 1
rlabel polysilicon 1129 -1865 1129 -1865 0 3
rlabel polysilicon 1136 -1859 1136 -1859 0 1
rlabel polysilicon 1136 -1865 1136 -1865 0 3
rlabel polysilicon 1143 -1859 1143 -1859 0 1
rlabel polysilicon 1143 -1865 1143 -1865 0 3
rlabel polysilicon 1150 -1859 1150 -1859 0 1
rlabel polysilicon 1150 -1865 1150 -1865 0 3
rlabel polysilicon 1157 -1859 1157 -1859 0 1
rlabel polysilicon 1157 -1865 1157 -1865 0 3
rlabel polysilicon 1164 -1859 1164 -1859 0 1
rlabel polysilicon 1164 -1865 1164 -1865 0 3
rlabel polysilicon 1171 -1859 1171 -1859 0 1
rlabel polysilicon 1171 -1865 1171 -1865 0 3
rlabel polysilicon 1178 -1859 1178 -1859 0 1
rlabel polysilicon 1178 -1865 1178 -1865 0 3
rlabel polysilicon 1185 -1859 1185 -1859 0 1
rlabel polysilicon 1185 -1865 1185 -1865 0 3
rlabel polysilicon 1192 -1859 1192 -1859 0 1
rlabel polysilicon 1192 -1865 1192 -1865 0 3
rlabel polysilicon 1199 -1859 1199 -1859 0 1
rlabel polysilicon 1199 -1865 1199 -1865 0 3
rlabel polysilicon 1206 -1859 1206 -1859 0 1
rlabel polysilicon 1206 -1865 1206 -1865 0 3
rlabel polysilicon 1213 -1859 1213 -1859 0 1
rlabel polysilicon 1213 -1865 1213 -1865 0 3
rlabel polysilicon 1220 -1859 1220 -1859 0 1
rlabel polysilicon 1220 -1865 1220 -1865 0 3
rlabel polysilicon 1227 -1859 1227 -1859 0 1
rlabel polysilicon 1227 -1865 1227 -1865 0 3
rlabel polysilicon 1234 -1859 1234 -1859 0 1
rlabel polysilicon 1234 -1865 1234 -1865 0 3
rlabel polysilicon 1241 -1859 1241 -1859 0 1
rlabel polysilicon 1241 -1865 1241 -1865 0 3
rlabel polysilicon 1248 -1859 1248 -1859 0 1
rlabel polysilicon 1248 -1865 1248 -1865 0 3
rlabel polysilicon 1255 -1859 1255 -1859 0 1
rlabel polysilicon 1258 -1859 1258 -1859 0 2
rlabel polysilicon 1255 -1865 1255 -1865 0 3
rlabel polysilicon 1262 -1859 1262 -1859 0 1
rlabel polysilicon 1262 -1865 1262 -1865 0 3
rlabel polysilicon 1269 -1859 1269 -1859 0 1
rlabel polysilicon 1269 -1865 1269 -1865 0 3
rlabel polysilicon 1276 -1859 1276 -1859 0 1
rlabel polysilicon 1276 -1865 1276 -1865 0 3
rlabel polysilicon 1283 -1859 1283 -1859 0 1
rlabel polysilicon 1283 -1865 1283 -1865 0 3
rlabel polysilicon 1290 -1859 1290 -1859 0 1
rlabel polysilicon 1290 -1865 1290 -1865 0 3
rlabel polysilicon 1297 -1859 1297 -1859 0 1
rlabel polysilicon 1297 -1865 1297 -1865 0 3
rlabel polysilicon 1304 -1859 1304 -1859 0 1
rlabel polysilicon 1304 -1865 1304 -1865 0 3
rlabel polysilicon 1311 -1859 1311 -1859 0 1
rlabel polysilicon 1311 -1865 1311 -1865 0 3
rlabel polysilicon 1318 -1859 1318 -1859 0 1
rlabel polysilicon 1318 -1865 1318 -1865 0 3
rlabel polysilicon 1325 -1859 1325 -1859 0 1
rlabel polysilicon 1325 -1865 1325 -1865 0 3
rlabel polysilicon 1332 -1859 1332 -1859 0 1
rlabel polysilicon 1332 -1865 1332 -1865 0 3
rlabel polysilicon 1339 -1859 1339 -1859 0 1
rlabel polysilicon 1339 -1865 1339 -1865 0 3
rlabel polysilicon 1346 -1859 1346 -1859 0 1
rlabel polysilicon 1346 -1865 1346 -1865 0 3
rlabel polysilicon 1353 -1859 1353 -1859 0 1
rlabel polysilicon 1353 -1865 1353 -1865 0 3
rlabel polysilicon 1360 -1859 1360 -1859 0 1
rlabel polysilicon 1360 -1865 1360 -1865 0 3
rlabel polysilicon 1367 -1859 1367 -1859 0 1
rlabel polysilicon 1367 -1865 1367 -1865 0 3
rlabel polysilicon 1374 -1859 1374 -1859 0 1
rlabel polysilicon 1374 -1865 1374 -1865 0 3
rlabel polysilicon 1381 -1859 1381 -1859 0 1
rlabel polysilicon 1381 -1865 1381 -1865 0 3
rlabel polysilicon 1388 -1859 1388 -1859 0 1
rlabel polysilicon 1388 -1865 1388 -1865 0 3
rlabel polysilicon 1395 -1859 1395 -1859 0 1
rlabel polysilicon 1395 -1865 1395 -1865 0 3
rlabel polysilicon 1398 -1865 1398 -1865 0 4
rlabel polysilicon 1402 -1859 1402 -1859 0 1
rlabel polysilicon 1402 -1865 1402 -1865 0 3
rlabel polysilicon 1409 -1859 1409 -1859 0 1
rlabel polysilicon 1409 -1865 1409 -1865 0 3
rlabel polysilicon 1416 -1859 1416 -1859 0 1
rlabel polysilicon 1416 -1865 1416 -1865 0 3
rlabel polysilicon 1423 -1859 1423 -1859 0 1
rlabel polysilicon 1423 -1865 1423 -1865 0 3
rlabel polysilicon 1430 -1859 1430 -1859 0 1
rlabel polysilicon 1430 -1865 1430 -1865 0 3
rlabel polysilicon 2 -1986 2 -1986 0 1
rlabel polysilicon 2 -1992 2 -1992 0 3
rlabel polysilicon 9 -1986 9 -1986 0 1
rlabel polysilicon 9 -1992 9 -1992 0 3
rlabel polysilicon 16 -1986 16 -1986 0 1
rlabel polysilicon 16 -1992 16 -1992 0 3
rlabel polysilicon 23 -1986 23 -1986 0 1
rlabel polysilicon 26 -1986 26 -1986 0 2
rlabel polysilicon 23 -1992 23 -1992 0 3
rlabel polysilicon 30 -1986 30 -1986 0 1
rlabel polysilicon 30 -1992 30 -1992 0 3
rlabel polysilicon 37 -1986 37 -1986 0 1
rlabel polysilicon 40 -1986 40 -1986 0 2
rlabel polysilicon 37 -1992 37 -1992 0 3
rlabel polysilicon 40 -1992 40 -1992 0 4
rlabel polysilicon 44 -1986 44 -1986 0 1
rlabel polysilicon 44 -1992 44 -1992 0 3
rlabel polysilicon 51 -1986 51 -1986 0 1
rlabel polysilicon 51 -1992 51 -1992 0 3
rlabel polysilicon 58 -1986 58 -1986 0 1
rlabel polysilicon 58 -1992 58 -1992 0 3
rlabel polysilicon 65 -1986 65 -1986 0 1
rlabel polysilicon 68 -1986 68 -1986 0 2
rlabel polysilicon 65 -1992 65 -1992 0 3
rlabel polysilicon 68 -1992 68 -1992 0 4
rlabel polysilicon 72 -1986 72 -1986 0 1
rlabel polysilicon 75 -1986 75 -1986 0 2
rlabel polysilicon 72 -1992 72 -1992 0 3
rlabel polysilicon 75 -1992 75 -1992 0 4
rlabel polysilicon 79 -1986 79 -1986 0 1
rlabel polysilicon 79 -1992 79 -1992 0 3
rlabel polysilicon 86 -1986 86 -1986 0 1
rlabel polysilicon 86 -1992 86 -1992 0 3
rlabel polysilicon 93 -1986 93 -1986 0 1
rlabel polysilicon 93 -1992 93 -1992 0 3
rlabel polysilicon 100 -1986 100 -1986 0 1
rlabel polysilicon 100 -1992 100 -1992 0 3
rlabel polysilicon 107 -1986 107 -1986 0 1
rlabel polysilicon 107 -1992 107 -1992 0 3
rlabel polysilicon 114 -1986 114 -1986 0 1
rlabel polysilicon 114 -1992 114 -1992 0 3
rlabel polysilicon 121 -1986 121 -1986 0 1
rlabel polysilicon 121 -1992 121 -1992 0 3
rlabel polysilicon 128 -1986 128 -1986 0 1
rlabel polysilicon 128 -1992 128 -1992 0 3
rlabel polysilicon 135 -1986 135 -1986 0 1
rlabel polysilicon 135 -1992 135 -1992 0 3
rlabel polysilicon 142 -1986 142 -1986 0 1
rlabel polysilicon 142 -1992 142 -1992 0 3
rlabel polysilicon 149 -1986 149 -1986 0 1
rlabel polysilicon 149 -1992 149 -1992 0 3
rlabel polysilicon 156 -1986 156 -1986 0 1
rlabel polysilicon 156 -1992 156 -1992 0 3
rlabel polysilicon 163 -1986 163 -1986 0 1
rlabel polysilicon 163 -1992 163 -1992 0 3
rlabel polysilicon 170 -1986 170 -1986 0 1
rlabel polysilicon 173 -1986 173 -1986 0 2
rlabel polysilicon 170 -1992 170 -1992 0 3
rlabel polysilicon 173 -1992 173 -1992 0 4
rlabel polysilicon 177 -1986 177 -1986 0 1
rlabel polysilicon 177 -1992 177 -1992 0 3
rlabel polysilicon 184 -1986 184 -1986 0 1
rlabel polysilicon 184 -1992 184 -1992 0 3
rlabel polysilicon 191 -1986 191 -1986 0 1
rlabel polysilicon 191 -1992 191 -1992 0 3
rlabel polysilicon 198 -1986 198 -1986 0 1
rlabel polysilicon 198 -1992 198 -1992 0 3
rlabel polysilicon 205 -1986 205 -1986 0 1
rlabel polysilicon 205 -1992 205 -1992 0 3
rlabel polysilicon 212 -1986 212 -1986 0 1
rlabel polysilicon 212 -1992 212 -1992 0 3
rlabel polysilicon 219 -1986 219 -1986 0 1
rlabel polysilicon 219 -1992 219 -1992 0 3
rlabel polysilicon 226 -1986 226 -1986 0 1
rlabel polysilicon 229 -1986 229 -1986 0 2
rlabel polysilicon 226 -1992 226 -1992 0 3
rlabel polysilicon 229 -1992 229 -1992 0 4
rlabel polysilicon 233 -1986 233 -1986 0 1
rlabel polysilicon 233 -1992 233 -1992 0 3
rlabel polysilicon 240 -1986 240 -1986 0 1
rlabel polysilicon 240 -1992 240 -1992 0 3
rlabel polysilicon 247 -1986 247 -1986 0 1
rlabel polysilicon 247 -1992 247 -1992 0 3
rlabel polysilicon 254 -1986 254 -1986 0 1
rlabel polysilicon 254 -1992 254 -1992 0 3
rlabel polysilicon 261 -1986 261 -1986 0 1
rlabel polysilicon 261 -1992 261 -1992 0 3
rlabel polysilicon 268 -1986 268 -1986 0 1
rlabel polysilicon 268 -1992 268 -1992 0 3
rlabel polysilicon 275 -1986 275 -1986 0 1
rlabel polysilicon 275 -1992 275 -1992 0 3
rlabel polysilicon 282 -1986 282 -1986 0 1
rlabel polysilicon 282 -1992 282 -1992 0 3
rlabel polysilicon 289 -1986 289 -1986 0 1
rlabel polysilicon 289 -1992 289 -1992 0 3
rlabel polysilicon 296 -1986 296 -1986 0 1
rlabel polysilicon 296 -1992 296 -1992 0 3
rlabel polysilicon 303 -1986 303 -1986 0 1
rlabel polysilicon 303 -1992 303 -1992 0 3
rlabel polysilicon 310 -1986 310 -1986 0 1
rlabel polysilicon 310 -1992 310 -1992 0 3
rlabel polysilicon 317 -1986 317 -1986 0 1
rlabel polysilicon 317 -1992 317 -1992 0 3
rlabel polysilicon 324 -1986 324 -1986 0 1
rlabel polysilicon 324 -1992 324 -1992 0 3
rlabel polysilicon 331 -1986 331 -1986 0 1
rlabel polysilicon 331 -1992 331 -1992 0 3
rlabel polysilicon 338 -1986 338 -1986 0 1
rlabel polysilicon 338 -1992 338 -1992 0 3
rlabel polysilicon 345 -1986 345 -1986 0 1
rlabel polysilicon 345 -1992 345 -1992 0 3
rlabel polysilicon 352 -1986 352 -1986 0 1
rlabel polysilicon 355 -1986 355 -1986 0 2
rlabel polysilicon 352 -1992 352 -1992 0 3
rlabel polysilicon 355 -1992 355 -1992 0 4
rlabel polysilicon 359 -1986 359 -1986 0 1
rlabel polysilicon 359 -1992 359 -1992 0 3
rlabel polysilicon 366 -1986 366 -1986 0 1
rlabel polysilicon 366 -1992 366 -1992 0 3
rlabel polysilicon 373 -1986 373 -1986 0 1
rlabel polysilicon 373 -1992 373 -1992 0 3
rlabel polysilicon 376 -1992 376 -1992 0 4
rlabel polysilicon 380 -1986 380 -1986 0 1
rlabel polysilicon 380 -1992 380 -1992 0 3
rlabel polysilicon 387 -1986 387 -1986 0 1
rlabel polysilicon 387 -1992 387 -1992 0 3
rlabel polysilicon 394 -1986 394 -1986 0 1
rlabel polysilicon 394 -1992 394 -1992 0 3
rlabel polysilicon 401 -1986 401 -1986 0 1
rlabel polysilicon 401 -1992 401 -1992 0 3
rlabel polysilicon 408 -1986 408 -1986 0 1
rlabel polysilicon 411 -1986 411 -1986 0 2
rlabel polysilicon 408 -1992 408 -1992 0 3
rlabel polysilicon 411 -1992 411 -1992 0 4
rlabel polysilicon 415 -1986 415 -1986 0 1
rlabel polysilicon 415 -1992 415 -1992 0 3
rlabel polysilicon 422 -1986 422 -1986 0 1
rlabel polysilicon 422 -1992 422 -1992 0 3
rlabel polysilicon 429 -1986 429 -1986 0 1
rlabel polysilicon 429 -1992 429 -1992 0 3
rlabel polysilicon 436 -1986 436 -1986 0 1
rlabel polysilicon 436 -1992 436 -1992 0 3
rlabel polysilicon 443 -1986 443 -1986 0 1
rlabel polysilicon 443 -1992 443 -1992 0 3
rlabel polysilicon 450 -1986 450 -1986 0 1
rlabel polysilicon 450 -1992 450 -1992 0 3
rlabel polysilicon 457 -1986 457 -1986 0 1
rlabel polysilicon 457 -1992 457 -1992 0 3
rlabel polysilicon 464 -1986 464 -1986 0 1
rlabel polysilicon 464 -1992 464 -1992 0 3
rlabel polysilicon 471 -1986 471 -1986 0 1
rlabel polysilicon 471 -1992 471 -1992 0 3
rlabel polysilicon 478 -1986 478 -1986 0 1
rlabel polysilicon 478 -1992 478 -1992 0 3
rlabel polysilicon 485 -1986 485 -1986 0 1
rlabel polysilicon 485 -1992 485 -1992 0 3
rlabel polysilicon 492 -1986 492 -1986 0 1
rlabel polysilicon 492 -1992 492 -1992 0 3
rlabel polysilicon 499 -1986 499 -1986 0 1
rlabel polysilicon 499 -1992 499 -1992 0 3
rlabel polysilicon 506 -1986 506 -1986 0 1
rlabel polysilicon 509 -1986 509 -1986 0 2
rlabel polysilicon 506 -1992 506 -1992 0 3
rlabel polysilicon 509 -1992 509 -1992 0 4
rlabel polysilicon 513 -1986 513 -1986 0 1
rlabel polysilicon 516 -1986 516 -1986 0 2
rlabel polysilicon 513 -1992 513 -1992 0 3
rlabel polysilicon 516 -1992 516 -1992 0 4
rlabel polysilicon 520 -1986 520 -1986 0 1
rlabel polysilicon 523 -1986 523 -1986 0 2
rlabel polysilicon 520 -1992 520 -1992 0 3
rlabel polysilicon 523 -1992 523 -1992 0 4
rlabel polysilicon 527 -1986 527 -1986 0 1
rlabel polysilicon 527 -1992 527 -1992 0 3
rlabel polysilicon 534 -1986 534 -1986 0 1
rlabel polysilicon 534 -1992 534 -1992 0 3
rlabel polysilicon 541 -1986 541 -1986 0 1
rlabel polysilicon 541 -1992 541 -1992 0 3
rlabel polysilicon 548 -1986 548 -1986 0 1
rlabel polysilicon 548 -1992 548 -1992 0 3
rlabel polysilicon 555 -1986 555 -1986 0 1
rlabel polysilicon 555 -1992 555 -1992 0 3
rlabel polysilicon 562 -1986 562 -1986 0 1
rlabel polysilicon 565 -1986 565 -1986 0 2
rlabel polysilicon 562 -1992 562 -1992 0 3
rlabel polysilicon 569 -1986 569 -1986 0 1
rlabel polysilicon 569 -1992 569 -1992 0 3
rlabel polysilicon 576 -1986 576 -1986 0 1
rlabel polysilicon 579 -1986 579 -1986 0 2
rlabel polysilicon 576 -1992 576 -1992 0 3
rlabel polysilicon 579 -1992 579 -1992 0 4
rlabel polysilicon 583 -1986 583 -1986 0 1
rlabel polysilicon 583 -1992 583 -1992 0 3
rlabel polysilicon 586 -1992 586 -1992 0 4
rlabel polysilicon 590 -1986 590 -1986 0 1
rlabel polysilicon 590 -1992 590 -1992 0 3
rlabel polysilicon 597 -1986 597 -1986 0 1
rlabel polysilicon 597 -1992 597 -1992 0 3
rlabel polysilicon 604 -1986 604 -1986 0 1
rlabel polysilicon 604 -1992 604 -1992 0 3
rlabel polysilicon 611 -1986 611 -1986 0 1
rlabel polysilicon 614 -1986 614 -1986 0 2
rlabel polysilicon 611 -1992 611 -1992 0 3
rlabel polysilicon 614 -1992 614 -1992 0 4
rlabel polysilicon 618 -1986 618 -1986 0 1
rlabel polysilicon 618 -1992 618 -1992 0 3
rlabel polysilicon 625 -1986 625 -1986 0 1
rlabel polysilicon 625 -1992 625 -1992 0 3
rlabel polysilicon 632 -1986 632 -1986 0 1
rlabel polysilicon 632 -1992 632 -1992 0 3
rlabel polysilicon 639 -1986 639 -1986 0 1
rlabel polysilicon 642 -1986 642 -1986 0 2
rlabel polysilicon 639 -1992 639 -1992 0 3
rlabel polysilicon 642 -1992 642 -1992 0 4
rlabel polysilicon 646 -1986 646 -1986 0 1
rlabel polysilicon 646 -1992 646 -1992 0 3
rlabel polysilicon 653 -1986 653 -1986 0 1
rlabel polysilicon 653 -1992 653 -1992 0 3
rlabel polysilicon 660 -1986 660 -1986 0 1
rlabel polysilicon 663 -1986 663 -1986 0 2
rlabel polysilicon 660 -1992 660 -1992 0 3
rlabel polysilicon 663 -1992 663 -1992 0 4
rlabel polysilicon 667 -1986 667 -1986 0 1
rlabel polysilicon 667 -1992 667 -1992 0 3
rlabel polysilicon 674 -1986 674 -1986 0 1
rlabel polysilicon 674 -1992 674 -1992 0 3
rlabel polysilicon 681 -1986 681 -1986 0 1
rlabel polysilicon 681 -1992 681 -1992 0 3
rlabel polysilicon 688 -1986 688 -1986 0 1
rlabel polysilicon 688 -1992 688 -1992 0 3
rlabel polysilicon 695 -1986 695 -1986 0 1
rlabel polysilicon 695 -1992 695 -1992 0 3
rlabel polysilicon 702 -1986 702 -1986 0 1
rlabel polysilicon 705 -1986 705 -1986 0 2
rlabel polysilicon 702 -1992 702 -1992 0 3
rlabel polysilicon 705 -1992 705 -1992 0 4
rlabel polysilicon 709 -1986 709 -1986 0 1
rlabel polysilicon 709 -1992 709 -1992 0 3
rlabel polysilicon 716 -1986 716 -1986 0 1
rlabel polysilicon 716 -1992 716 -1992 0 3
rlabel polysilicon 723 -1986 723 -1986 0 1
rlabel polysilicon 726 -1986 726 -1986 0 2
rlabel polysilicon 723 -1992 723 -1992 0 3
rlabel polysilicon 726 -1992 726 -1992 0 4
rlabel polysilicon 730 -1986 730 -1986 0 1
rlabel polysilicon 730 -1992 730 -1992 0 3
rlabel polysilicon 737 -1986 737 -1986 0 1
rlabel polysilicon 737 -1992 737 -1992 0 3
rlabel polysilicon 744 -1986 744 -1986 0 1
rlabel polysilicon 744 -1992 744 -1992 0 3
rlabel polysilicon 751 -1986 751 -1986 0 1
rlabel polysilicon 754 -1986 754 -1986 0 2
rlabel polysilicon 751 -1992 751 -1992 0 3
rlabel polysilicon 754 -1992 754 -1992 0 4
rlabel polysilicon 758 -1986 758 -1986 0 1
rlabel polysilicon 758 -1992 758 -1992 0 3
rlabel polysilicon 765 -1986 765 -1986 0 1
rlabel polysilicon 765 -1992 765 -1992 0 3
rlabel polysilicon 772 -1986 772 -1986 0 1
rlabel polysilicon 772 -1992 772 -1992 0 3
rlabel polysilicon 779 -1986 779 -1986 0 1
rlabel polysilicon 782 -1986 782 -1986 0 2
rlabel polysilicon 779 -1992 779 -1992 0 3
rlabel polysilicon 782 -1992 782 -1992 0 4
rlabel polysilicon 786 -1986 786 -1986 0 1
rlabel polysilicon 786 -1992 786 -1992 0 3
rlabel polysilicon 793 -1986 793 -1986 0 1
rlabel polysilicon 793 -1992 793 -1992 0 3
rlabel polysilicon 800 -1986 800 -1986 0 1
rlabel polysilicon 800 -1992 800 -1992 0 3
rlabel polysilicon 807 -1986 807 -1986 0 1
rlabel polysilicon 807 -1992 807 -1992 0 3
rlabel polysilicon 810 -1992 810 -1992 0 4
rlabel polysilicon 814 -1986 814 -1986 0 1
rlabel polysilicon 814 -1992 814 -1992 0 3
rlabel polysilicon 821 -1986 821 -1986 0 1
rlabel polysilicon 821 -1992 821 -1992 0 3
rlabel polysilicon 828 -1986 828 -1986 0 1
rlabel polysilicon 828 -1992 828 -1992 0 3
rlabel polysilicon 835 -1986 835 -1986 0 1
rlabel polysilicon 835 -1992 835 -1992 0 3
rlabel polysilicon 842 -1986 842 -1986 0 1
rlabel polysilicon 842 -1992 842 -1992 0 3
rlabel polysilicon 852 -1986 852 -1986 0 2
rlabel polysilicon 849 -1992 849 -1992 0 3
rlabel polysilicon 852 -1992 852 -1992 0 4
rlabel polysilicon 856 -1986 856 -1986 0 1
rlabel polysilicon 856 -1992 856 -1992 0 3
rlabel polysilicon 863 -1986 863 -1986 0 1
rlabel polysilicon 863 -1992 863 -1992 0 3
rlabel polysilicon 870 -1986 870 -1986 0 1
rlabel polysilicon 870 -1992 870 -1992 0 3
rlabel polysilicon 877 -1986 877 -1986 0 1
rlabel polysilicon 877 -1992 877 -1992 0 3
rlabel polysilicon 884 -1986 884 -1986 0 1
rlabel polysilicon 884 -1992 884 -1992 0 3
rlabel polysilicon 891 -1986 891 -1986 0 1
rlabel polysilicon 891 -1992 891 -1992 0 3
rlabel polysilicon 898 -1986 898 -1986 0 1
rlabel polysilicon 898 -1992 898 -1992 0 3
rlabel polysilicon 905 -1986 905 -1986 0 1
rlabel polysilicon 905 -1992 905 -1992 0 3
rlabel polysilicon 912 -1986 912 -1986 0 1
rlabel polysilicon 912 -1992 912 -1992 0 3
rlabel polysilicon 919 -1986 919 -1986 0 1
rlabel polysilicon 919 -1992 919 -1992 0 3
rlabel polysilicon 926 -1986 926 -1986 0 1
rlabel polysilicon 926 -1992 926 -1992 0 3
rlabel polysilicon 933 -1986 933 -1986 0 1
rlabel polysilicon 933 -1992 933 -1992 0 3
rlabel polysilicon 940 -1986 940 -1986 0 1
rlabel polysilicon 940 -1992 940 -1992 0 3
rlabel polysilicon 947 -1986 947 -1986 0 1
rlabel polysilicon 947 -1992 947 -1992 0 3
rlabel polysilicon 954 -1986 954 -1986 0 1
rlabel polysilicon 954 -1992 954 -1992 0 3
rlabel polysilicon 961 -1986 961 -1986 0 1
rlabel polysilicon 961 -1992 961 -1992 0 3
rlabel polysilicon 968 -1986 968 -1986 0 1
rlabel polysilicon 968 -1992 968 -1992 0 3
rlabel polysilicon 975 -1986 975 -1986 0 1
rlabel polysilicon 975 -1992 975 -1992 0 3
rlabel polysilicon 982 -1986 982 -1986 0 1
rlabel polysilicon 982 -1992 982 -1992 0 3
rlabel polysilicon 989 -1986 989 -1986 0 1
rlabel polysilicon 989 -1992 989 -1992 0 3
rlabel polysilicon 996 -1986 996 -1986 0 1
rlabel polysilicon 996 -1992 996 -1992 0 3
rlabel polysilicon 1003 -1986 1003 -1986 0 1
rlabel polysilicon 1003 -1992 1003 -1992 0 3
rlabel polysilicon 1010 -1986 1010 -1986 0 1
rlabel polysilicon 1010 -1992 1010 -1992 0 3
rlabel polysilicon 1017 -1986 1017 -1986 0 1
rlabel polysilicon 1017 -1992 1017 -1992 0 3
rlabel polysilicon 1024 -1986 1024 -1986 0 1
rlabel polysilicon 1024 -1992 1024 -1992 0 3
rlabel polysilicon 1031 -1986 1031 -1986 0 1
rlabel polysilicon 1031 -1992 1031 -1992 0 3
rlabel polysilicon 1038 -1986 1038 -1986 0 1
rlabel polysilicon 1038 -1992 1038 -1992 0 3
rlabel polysilicon 1045 -1986 1045 -1986 0 1
rlabel polysilicon 1045 -1992 1045 -1992 0 3
rlabel polysilicon 1052 -1986 1052 -1986 0 1
rlabel polysilicon 1052 -1992 1052 -1992 0 3
rlabel polysilicon 1059 -1986 1059 -1986 0 1
rlabel polysilicon 1059 -1992 1059 -1992 0 3
rlabel polysilicon 1066 -1986 1066 -1986 0 1
rlabel polysilicon 1066 -1992 1066 -1992 0 3
rlabel polysilicon 1073 -1986 1073 -1986 0 1
rlabel polysilicon 1073 -1992 1073 -1992 0 3
rlabel polysilicon 1080 -1986 1080 -1986 0 1
rlabel polysilicon 1080 -1992 1080 -1992 0 3
rlabel polysilicon 1087 -1986 1087 -1986 0 1
rlabel polysilicon 1087 -1992 1087 -1992 0 3
rlabel polysilicon 1094 -1986 1094 -1986 0 1
rlabel polysilicon 1094 -1992 1094 -1992 0 3
rlabel polysilicon 1101 -1986 1101 -1986 0 1
rlabel polysilicon 1101 -1992 1101 -1992 0 3
rlabel polysilicon 1108 -1986 1108 -1986 0 1
rlabel polysilicon 1108 -1992 1108 -1992 0 3
rlabel polysilicon 1115 -1986 1115 -1986 0 1
rlabel polysilicon 1115 -1992 1115 -1992 0 3
rlabel polysilicon 1122 -1986 1122 -1986 0 1
rlabel polysilicon 1122 -1992 1122 -1992 0 3
rlabel polysilicon 1129 -1986 1129 -1986 0 1
rlabel polysilicon 1129 -1992 1129 -1992 0 3
rlabel polysilicon 1136 -1986 1136 -1986 0 1
rlabel polysilicon 1136 -1992 1136 -1992 0 3
rlabel polysilicon 1143 -1986 1143 -1986 0 1
rlabel polysilicon 1143 -1992 1143 -1992 0 3
rlabel polysilicon 1150 -1986 1150 -1986 0 1
rlabel polysilicon 1150 -1992 1150 -1992 0 3
rlabel polysilicon 1157 -1986 1157 -1986 0 1
rlabel polysilicon 1157 -1992 1157 -1992 0 3
rlabel polysilicon 1164 -1986 1164 -1986 0 1
rlabel polysilicon 1164 -1992 1164 -1992 0 3
rlabel polysilicon 1171 -1986 1171 -1986 0 1
rlabel polysilicon 1171 -1992 1171 -1992 0 3
rlabel polysilicon 1178 -1986 1178 -1986 0 1
rlabel polysilicon 1178 -1992 1178 -1992 0 3
rlabel polysilicon 1185 -1986 1185 -1986 0 1
rlabel polysilicon 1185 -1992 1185 -1992 0 3
rlabel polysilicon 1192 -1986 1192 -1986 0 1
rlabel polysilicon 1192 -1992 1192 -1992 0 3
rlabel polysilicon 1199 -1986 1199 -1986 0 1
rlabel polysilicon 1199 -1992 1199 -1992 0 3
rlabel polysilicon 1206 -1986 1206 -1986 0 1
rlabel polysilicon 1206 -1992 1206 -1992 0 3
rlabel polysilicon 1213 -1986 1213 -1986 0 1
rlabel polysilicon 1213 -1992 1213 -1992 0 3
rlabel polysilicon 1220 -1986 1220 -1986 0 1
rlabel polysilicon 1220 -1992 1220 -1992 0 3
rlabel polysilicon 1227 -1986 1227 -1986 0 1
rlabel polysilicon 1227 -1992 1227 -1992 0 3
rlabel polysilicon 1234 -1986 1234 -1986 0 1
rlabel polysilicon 1234 -1992 1234 -1992 0 3
rlabel polysilicon 1241 -1986 1241 -1986 0 1
rlabel polysilicon 1241 -1992 1241 -1992 0 3
rlabel polysilicon 1248 -1986 1248 -1986 0 1
rlabel polysilicon 1248 -1992 1248 -1992 0 3
rlabel polysilicon 1255 -1986 1255 -1986 0 1
rlabel polysilicon 1255 -1992 1255 -1992 0 3
rlabel polysilicon 1262 -1986 1262 -1986 0 1
rlabel polysilicon 1262 -1992 1262 -1992 0 3
rlabel polysilicon 1269 -1986 1269 -1986 0 1
rlabel polysilicon 1269 -1992 1269 -1992 0 3
rlabel polysilicon 1276 -1986 1276 -1986 0 1
rlabel polysilicon 1276 -1992 1276 -1992 0 3
rlabel polysilicon 1283 -1986 1283 -1986 0 1
rlabel polysilicon 1283 -1992 1283 -1992 0 3
rlabel polysilicon 1290 -1986 1290 -1986 0 1
rlabel polysilicon 1290 -1992 1290 -1992 0 3
rlabel polysilicon 1297 -1986 1297 -1986 0 1
rlabel polysilicon 1297 -1992 1297 -1992 0 3
rlabel polysilicon 1304 -1986 1304 -1986 0 1
rlabel polysilicon 1304 -1992 1304 -1992 0 3
rlabel polysilicon 1311 -1986 1311 -1986 0 1
rlabel polysilicon 1311 -1992 1311 -1992 0 3
rlabel polysilicon 1318 -1986 1318 -1986 0 1
rlabel polysilicon 1318 -1992 1318 -1992 0 3
rlabel polysilicon 1325 -1986 1325 -1986 0 1
rlabel polysilicon 1325 -1992 1325 -1992 0 3
rlabel polysilicon 1332 -1986 1332 -1986 0 1
rlabel polysilicon 1332 -1992 1332 -1992 0 3
rlabel polysilicon 1339 -1986 1339 -1986 0 1
rlabel polysilicon 1339 -1992 1339 -1992 0 3
rlabel polysilicon 1346 -1986 1346 -1986 0 1
rlabel polysilicon 1346 -1992 1346 -1992 0 3
rlabel polysilicon 1353 -1986 1353 -1986 0 1
rlabel polysilicon 1353 -1992 1353 -1992 0 3
rlabel polysilicon 1360 -1986 1360 -1986 0 1
rlabel polysilicon 1360 -1992 1360 -1992 0 3
rlabel polysilicon 1367 -1986 1367 -1986 0 1
rlabel polysilicon 1367 -1992 1367 -1992 0 3
rlabel polysilicon 1374 -1986 1374 -1986 0 1
rlabel polysilicon 1374 -1992 1374 -1992 0 3
rlabel polysilicon 1381 -1986 1381 -1986 0 1
rlabel polysilicon 1381 -1992 1381 -1992 0 3
rlabel polysilicon 1388 -1986 1388 -1986 0 1
rlabel polysilicon 1388 -1992 1388 -1992 0 3
rlabel polysilicon 1395 -1986 1395 -1986 0 1
rlabel polysilicon 1395 -1992 1395 -1992 0 3
rlabel polysilicon 1402 -1986 1402 -1986 0 1
rlabel polysilicon 1402 -1992 1402 -1992 0 3
rlabel polysilicon 2 -2105 2 -2105 0 1
rlabel polysilicon 5 -2105 5 -2105 0 2
rlabel polysilicon 5 -2111 5 -2111 0 4
rlabel polysilicon 9 -2105 9 -2105 0 1
rlabel polysilicon 9 -2111 9 -2111 0 3
rlabel polysilicon 16 -2105 16 -2105 0 1
rlabel polysilicon 16 -2111 16 -2111 0 3
rlabel polysilicon 23 -2105 23 -2105 0 1
rlabel polysilicon 23 -2111 23 -2111 0 3
rlabel polysilicon 30 -2105 30 -2105 0 1
rlabel polysilicon 30 -2111 30 -2111 0 3
rlabel polysilicon 37 -2105 37 -2105 0 1
rlabel polysilicon 37 -2111 37 -2111 0 3
rlabel polysilicon 44 -2105 44 -2105 0 1
rlabel polysilicon 44 -2111 44 -2111 0 3
rlabel polysilicon 51 -2105 51 -2105 0 1
rlabel polysilicon 51 -2111 51 -2111 0 3
rlabel polysilicon 58 -2105 58 -2105 0 1
rlabel polysilicon 58 -2111 58 -2111 0 3
rlabel polysilicon 65 -2105 65 -2105 0 1
rlabel polysilicon 65 -2111 65 -2111 0 3
rlabel polysilicon 72 -2105 72 -2105 0 1
rlabel polysilicon 72 -2111 72 -2111 0 3
rlabel polysilicon 79 -2105 79 -2105 0 1
rlabel polysilicon 79 -2111 79 -2111 0 3
rlabel polysilicon 86 -2105 86 -2105 0 1
rlabel polysilicon 86 -2111 86 -2111 0 3
rlabel polysilicon 93 -2105 93 -2105 0 1
rlabel polysilicon 96 -2105 96 -2105 0 2
rlabel polysilicon 93 -2111 93 -2111 0 3
rlabel polysilicon 100 -2105 100 -2105 0 1
rlabel polysilicon 100 -2111 100 -2111 0 3
rlabel polysilicon 107 -2105 107 -2105 0 1
rlabel polysilicon 110 -2105 110 -2105 0 2
rlabel polysilicon 107 -2111 107 -2111 0 3
rlabel polysilicon 110 -2111 110 -2111 0 4
rlabel polysilicon 114 -2105 114 -2105 0 1
rlabel polysilicon 114 -2111 114 -2111 0 3
rlabel polysilicon 121 -2105 121 -2105 0 1
rlabel polysilicon 121 -2111 121 -2111 0 3
rlabel polysilicon 128 -2105 128 -2105 0 1
rlabel polysilicon 131 -2105 131 -2105 0 2
rlabel polysilicon 128 -2111 128 -2111 0 3
rlabel polysilicon 131 -2111 131 -2111 0 4
rlabel polysilicon 135 -2105 135 -2105 0 1
rlabel polysilicon 135 -2111 135 -2111 0 3
rlabel polysilicon 142 -2105 142 -2105 0 1
rlabel polysilicon 142 -2111 142 -2111 0 3
rlabel polysilicon 149 -2105 149 -2105 0 1
rlabel polysilicon 149 -2111 149 -2111 0 3
rlabel polysilicon 156 -2105 156 -2105 0 1
rlabel polysilicon 156 -2111 156 -2111 0 3
rlabel polysilicon 163 -2105 163 -2105 0 1
rlabel polysilicon 166 -2105 166 -2105 0 2
rlabel polysilicon 170 -2105 170 -2105 0 1
rlabel polysilicon 173 -2105 173 -2105 0 2
rlabel polysilicon 170 -2111 170 -2111 0 3
rlabel polysilicon 177 -2105 177 -2105 0 1
rlabel polysilicon 177 -2111 177 -2111 0 3
rlabel polysilicon 184 -2105 184 -2105 0 1
rlabel polysilicon 184 -2111 184 -2111 0 3
rlabel polysilicon 191 -2105 191 -2105 0 1
rlabel polysilicon 191 -2111 191 -2111 0 3
rlabel polysilicon 198 -2105 198 -2105 0 1
rlabel polysilicon 198 -2111 198 -2111 0 3
rlabel polysilicon 205 -2105 205 -2105 0 1
rlabel polysilicon 205 -2111 205 -2111 0 3
rlabel polysilicon 212 -2105 212 -2105 0 1
rlabel polysilicon 212 -2111 212 -2111 0 3
rlabel polysilicon 219 -2105 219 -2105 0 1
rlabel polysilicon 219 -2111 219 -2111 0 3
rlabel polysilicon 226 -2105 226 -2105 0 1
rlabel polysilicon 226 -2111 226 -2111 0 3
rlabel polysilicon 233 -2105 233 -2105 0 1
rlabel polysilicon 240 -2105 240 -2105 0 1
rlabel polysilicon 240 -2111 240 -2111 0 3
rlabel polysilicon 247 -2105 247 -2105 0 1
rlabel polysilicon 247 -2111 247 -2111 0 3
rlabel polysilicon 254 -2105 254 -2105 0 1
rlabel polysilicon 254 -2111 254 -2111 0 3
rlabel polysilicon 261 -2105 261 -2105 0 1
rlabel polysilicon 261 -2111 261 -2111 0 3
rlabel polysilicon 268 -2105 268 -2105 0 1
rlabel polysilicon 268 -2111 268 -2111 0 3
rlabel polysilicon 275 -2105 275 -2105 0 1
rlabel polysilicon 275 -2111 275 -2111 0 3
rlabel polysilicon 282 -2105 282 -2105 0 1
rlabel polysilicon 282 -2111 282 -2111 0 3
rlabel polysilicon 289 -2105 289 -2105 0 1
rlabel polysilicon 289 -2111 289 -2111 0 3
rlabel polysilicon 296 -2105 296 -2105 0 1
rlabel polysilicon 296 -2111 296 -2111 0 3
rlabel polysilicon 303 -2105 303 -2105 0 1
rlabel polysilicon 303 -2111 303 -2111 0 3
rlabel polysilicon 310 -2105 310 -2105 0 1
rlabel polysilicon 310 -2111 310 -2111 0 3
rlabel polysilicon 317 -2105 317 -2105 0 1
rlabel polysilicon 320 -2105 320 -2105 0 2
rlabel polysilicon 317 -2111 317 -2111 0 3
rlabel polysilicon 320 -2111 320 -2111 0 4
rlabel polysilicon 324 -2105 324 -2105 0 1
rlabel polysilicon 324 -2111 324 -2111 0 3
rlabel polysilicon 331 -2105 331 -2105 0 1
rlabel polysilicon 334 -2105 334 -2105 0 2
rlabel polysilicon 331 -2111 331 -2111 0 3
rlabel polysilicon 334 -2111 334 -2111 0 4
rlabel polysilicon 338 -2105 338 -2105 0 1
rlabel polysilicon 338 -2111 338 -2111 0 3
rlabel polysilicon 345 -2105 345 -2105 0 1
rlabel polysilicon 348 -2111 348 -2111 0 4
rlabel polysilicon 352 -2105 352 -2105 0 1
rlabel polysilicon 352 -2111 352 -2111 0 3
rlabel polysilicon 359 -2105 359 -2105 0 1
rlabel polysilicon 359 -2111 359 -2111 0 3
rlabel polysilicon 366 -2105 366 -2105 0 1
rlabel polysilicon 366 -2111 366 -2111 0 3
rlabel polysilicon 373 -2105 373 -2105 0 1
rlabel polysilicon 373 -2111 373 -2111 0 3
rlabel polysilicon 380 -2105 380 -2105 0 1
rlabel polysilicon 380 -2111 380 -2111 0 3
rlabel polysilicon 387 -2105 387 -2105 0 1
rlabel polysilicon 387 -2111 387 -2111 0 3
rlabel polysilicon 394 -2105 394 -2105 0 1
rlabel polysilicon 394 -2111 394 -2111 0 3
rlabel polysilicon 401 -2105 401 -2105 0 1
rlabel polysilicon 401 -2111 401 -2111 0 3
rlabel polysilicon 408 -2105 408 -2105 0 1
rlabel polysilicon 408 -2111 408 -2111 0 3
rlabel polysilicon 415 -2105 415 -2105 0 1
rlabel polysilicon 415 -2111 415 -2111 0 3
rlabel polysilicon 422 -2105 422 -2105 0 1
rlabel polysilicon 422 -2111 422 -2111 0 3
rlabel polysilicon 429 -2105 429 -2105 0 1
rlabel polysilicon 429 -2111 429 -2111 0 3
rlabel polysilicon 436 -2105 436 -2105 0 1
rlabel polysilicon 436 -2111 436 -2111 0 3
rlabel polysilicon 443 -2105 443 -2105 0 1
rlabel polysilicon 443 -2111 443 -2111 0 3
rlabel polysilicon 450 -2105 450 -2105 0 1
rlabel polysilicon 453 -2105 453 -2105 0 2
rlabel polysilicon 450 -2111 450 -2111 0 3
rlabel polysilicon 453 -2111 453 -2111 0 4
rlabel polysilicon 457 -2105 457 -2105 0 1
rlabel polysilicon 457 -2111 457 -2111 0 3
rlabel polysilicon 464 -2105 464 -2105 0 1
rlabel polysilicon 464 -2111 464 -2111 0 3
rlabel polysilicon 471 -2105 471 -2105 0 1
rlabel polysilicon 471 -2111 471 -2111 0 3
rlabel polysilicon 478 -2105 478 -2105 0 1
rlabel polysilicon 478 -2111 478 -2111 0 3
rlabel polysilicon 485 -2105 485 -2105 0 1
rlabel polysilicon 488 -2105 488 -2105 0 2
rlabel polysilicon 485 -2111 485 -2111 0 3
rlabel polysilicon 488 -2111 488 -2111 0 4
rlabel polysilicon 492 -2105 492 -2105 0 1
rlabel polysilicon 492 -2111 492 -2111 0 3
rlabel polysilicon 499 -2105 499 -2105 0 1
rlabel polysilicon 502 -2105 502 -2105 0 2
rlabel polysilicon 499 -2111 499 -2111 0 3
rlabel polysilicon 502 -2111 502 -2111 0 4
rlabel polysilicon 506 -2105 506 -2105 0 1
rlabel polysilicon 506 -2111 506 -2111 0 3
rlabel polysilicon 513 -2105 513 -2105 0 1
rlabel polysilicon 513 -2111 513 -2111 0 3
rlabel polysilicon 520 -2105 520 -2105 0 1
rlabel polysilicon 520 -2111 520 -2111 0 3
rlabel polysilicon 527 -2105 527 -2105 0 1
rlabel polysilicon 527 -2111 527 -2111 0 3
rlabel polysilicon 534 -2105 534 -2105 0 1
rlabel polysilicon 534 -2111 534 -2111 0 3
rlabel polysilicon 541 -2105 541 -2105 0 1
rlabel polysilicon 541 -2111 541 -2111 0 3
rlabel polysilicon 548 -2105 548 -2105 0 1
rlabel polysilicon 548 -2111 548 -2111 0 3
rlabel polysilicon 555 -2105 555 -2105 0 1
rlabel polysilicon 555 -2111 555 -2111 0 3
rlabel polysilicon 562 -2105 562 -2105 0 1
rlabel polysilicon 562 -2111 562 -2111 0 3
rlabel polysilicon 569 -2105 569 -2105 0 1
rlabel polysilicon 569 -2111 569 -2111 0 3
rlabel polysilicon 576 -2105 576 -2105 0 1
rlabel polysilicon 579 -2105 579 -2105 0 2
rlabel polysilicon 576 -2111 576 -2111 0 3
rlabel polysilicon 579 -2111 579 -2111 0 4
rlabel polysilicon 583 -2105 583 -2105 0 1
rlabel polysilicon 583 -2111 583 -2111 0 3
rlabel polysilicon 590 -2105 590 -2105 0 1
rlabel polysilicon 590 -2111 590 -2111 0 3
rlabel polysilicon 597 -2105 597 -2105 0 1
rlabel polysilicon 597 -2111 597 -2111 0 3
rlabel polysilicon 604 -2105 604 -2105 0 1
rlabel polysilicon 604 -2111 604 -2111 0 3
rlabel polysilicon 611 -2105 611 -2105 0 1
rlabel polysilicon 611 -2111 611 -2111 0 3
rlabel polysilicon 618 -2105 618 -2105 0 1
rlabel polysilicon 621 -2105 621 -2105 0 2
rlabel polysilicon 618 -2111 618 -2111 0 3
rlabel polysilicon 621 -2111 621 -2111 0 4
rlabel polysilicon 625 -2105 625 -2105 0 1
rlabel polysilicon 625 -2111 625 -2111 0 3
rlabel polysilicon 632 -2105 632 -2105 0 1
rlabel polysilicon 632 -2111 632 -2111 0 3
rlabel polysilicon 639 -2105 639 -2105 0 1
rlabel polysilicon 639 -2111 639 -2111 0 3
rlabel polysilicon 646 -2105 646 -2105 0 1
rlabel polysilicon 646 -2111 646 -2111 0 3
rlabel polysilicon 653 -2105 653 -2105 0 1
rlabel polysilicon 653 -2111 653 -2111 0 3
rlabel polysilicon 660 -2105 660 -2105 0 1
rlabel polysilicon 660 -2111 660 -2111 0 3
rlabel polysilicon 667 -2105 667 -2105 0 1
rlabel polysilicon 670 -2105 670 -2105 0 2
rlabel polysilicon 667 -2111 667 -2111 0 3
rlabel polysilicon 674 -2105 674 -2105 0 1
rlabel polysilicon 674 -2111 674 -2111 0 3
rlabel polysilicon 681 -2105 681 -2105 0 1
rlabel polysilicon 681 -2111 681 -2111 0 3
rlabel polysilicon 688 -2105 688 -2105 0 1
rlabel polysilicon 691 -2105 691 -2105 0 2
rlabel polysilicon 688 -2111 688 -2111 0 3
rlabel polysilicon 691 -2111 691 -2111 0 4
rlabel polysilicon 695 -2105 695 -2105 0 1
rlabel polysilicon 695 -2111 695 -2111 0 3
rlabel polysilicon 702 -2105 702 -2105 0 1
rlabel polysilicon 702 -2111 702 -2111 0 3
rlabel polysilicon 709 -2105 709 -2105 0 1
rlabel polysilicon 709 -2111 709 -2111 0 3
rlabel polysilicon 716 -2105 716 -2105 0 1
rlabel polysilicon 716 -2111 716 -2111 0 3
rlabel polysilicon 723 -2105 723 -2105 0 1
rlabel polysilicon 723 -2111 723 -2111 0 3
rlabel polysilicon 730 -2105 730 -2105 0 1
rlabel polysilicon 730 -2111 730 -2111 0 3
rlabel polysilicon 737 -2105 737 -2105 0 1
rlabel polysilicon 737 -2111 737 -2111 0 3
rlabel polysilicon 744 -2105 744 -2105 0 1
rlabel polysilicon 744 -2111 744 -2111 0 3
rlabel polysilicon 751 -2105 751 -2105 0 1
rlabel polysilicon 751 -2111 751 -2111 0 3
rlabel polysilicon 758 -2105 758 -2105 0 1
rlabel polysilicon 758 -2111 758 -2111 0 3
rlabel polysilicon 765 -2105 765 -2105 0 1
rlabel polysilicon 765 -2111 765 -2111 0 3
rlabel polysilicon 768 -2111 768 -2111 0 4
rlabel polysilicon 772 -2105 772 -2105 0 1
rlabel polysilicon 772 -2111 772 -2111 0 3
rlabel polysilicon 779 -2105 779 -2105 0 1
rlabel polysilicon 782 -2105 782 -2105 0 2
rlabel polysilicon 782 -2111 782 -2111 0 4
rlabel polysilicon 786 -2105 786 -2105 0 1
rlabel polysilicon 786 -2111 786 -2111 0 3
rlabel polysilicon 793 -2105 793 -2105 0 1
rlabel polysilicon 793 -2111 793 -2111 0 3
rlabel polysilicon 800 -2105 800 -2105 0 1
rlabel polysilicon 800 -2111 800 -2111 0 3
rlabel polysilicon 807 -2105 807 -2105 0 1
rlabel polysilicon 807 -2111 807 -2111 0 3
rlabel polysilicon 814 -2105 814 -2105 0 1
rlabel polysilicon 817 -2105 817 -2105 0 2
rlabel polysilicon 814 -2111 814 -2111 0 3
rlabel polysilicon 817 -2111 817 -2111 0 4
rlabel polysilicon 821 -2105 821 -2105 0 1
rlabel polysilicon 824 -2105 824 -2105 0 2
rlabel polysilicon 824 -2111 824 -2111 0 4
rlabel polysilicon 828 -2105 828 -2105 0 1
rlabel polysilicon 828 -2111 828 -2111 0 3
rlabel polysilicon 835 -2105 835 -2105 0 1
rlabel polysilicon 835 -2111 835 -2111 0 3
rlabel polysilicon 842 -2105 842 -2105 0 1
rlabel polysilicon 842 -2111 842 -2111 0 3
rlabel polysilicon 849 -2105 849 -2105 0 1
rlabel polysilicon 849 -2111 849 -2111 0 3
rlabel polysilicon 856 -2105 856 -2105 0 1
rlabel polysilicon 856 -2111 856 -2111 0 3
rlabel polysilicon 863 -2105 863 -2105 0 1
rlabel polysilicon 863 -2111 863 -2111 0 3
rlabel polysilicon 870 -2105 870 -2105 0 1
rlabel polysilicon 870 -2111 870 -2111 0 3
rlabel polysilicon 877 -2105 877 -2105 0 1
rlabel polysilicon 877 -2111 877 -2111 0 3
rlabel polysilicon 884 -2105 884 -2105 0 1
rlabel polysilicon 884 -2111 884 -2111 0 3
rlabel polysilicon 894 -2105 894 -2105 0 2
rlabel polysilicon 891 -2111 891 -2111 0 3
rlabel polysilicon 894 -2111 894 -2111 0 4
rlabel polysilicon 898 -2105 898 -2105 0 1
rlabel polysilicon 898 -2111 898 -2111 0 3
rlabel polysilicon 905 -2105 905 -2105 0 1
rlabel polysilicon 905 -2111 905 -2111 0 3
rlabel polysilicon 912 -2105 912 -2105 0 1
rlabel polysilicon 912 -2111 912 -2111 0 3
rlabel polysilicon 919 -2105 919 -2105 0 1
rlabel polysilicon 919 -2111 919 -2111 0 3
rlabel polysilicon 926 -2105 926 -2105 0 1
rlabel polysilicon 926 -2111 926 -2111 0 3
rlabel polysilicon 933 -2105 933 -2105 0 1
rlabel polysilicon 933 -2111 933 -2111 0 3
rlabel polysilicon 940 -2105 940 -2105 0 1
rlabel polysilicon 940 -2111 940 -2111 0 3
rlabel polysilicon 947 -2105 947 -2105 0 1
rlabel polysilicon 947 -2111 947 -2111 0 3
rlabel polysilicon 954 -2105 954 -2105 0 1
rlabel polysilicon 954 -2111 954 -2111 0 3
rlabel polysilicon 961 -2105 961 -2105 0 1
rlabel polysilicon 961 -2111 961 -2111 0 3
rlabel polysilicon 968 -2105 968 -2105 0 1
rlabel polysilicon 971 -2105 971 -2105 0 2
rlabel polysilicon 968 -2111 968 -2111 0 3
rlabel polysilicon 971 -2111 971 -2111 0 4
rlabel polysilicon 975 -2105 975 -2105 0 1
rlabel polysilicon 975 -2111 975 -2111 0 3
rlabel polysilicon 982 -2105 982 -2105 0 1
rlabel polysilicon 982 -2111 982 -2111 0 3
rlabel polysilicon 992 -2105 992 -2105 0 2
rlabel polysilicon 989 -2111 989 -2111 0 3
rlabel polysilicon 992 -2111 992 -2111 0 4
rlabel polysilicon 996 -2105 996 -2105 0 1
rlabel polysilicon 996 -2111 996 -2111 0 3
rlabel polysilicon 1003 -2105 1003 -2105 0 1
rlabel polysilicon 1003 -2111 1003 -2111 0 3
rlabel polysilicon 1010 -2105 1010 -2105 0 1
rlabel polysilicon 1010 -2111 1010 -2111 0 3
rlabel polysilicon 1017 -2105 1017 -2105 0 1
rlabel polysilicon 1017 -2111 1017 -2111 0 3
rlabel polysilicon 1024 -2105 1024 -2105 0 1
rlabel polysilicon 1024 -2111 1024 -2111 0 3
rlabel polysilicon 1031 -2105 1031 -2105 0 1
rlabel polysilicon 1031 -2111 1031 -2111 0 3
rlabel polysilicon 1038 -2105 1038 -2105 0 1
rlabel polysilicon 1038 -2111 1038 -2111 0 3
rlabel polysilicon 1045 -2105 1045 -2105 0 1
rlabel polysilicon 1045 -2111 1045 -2111 0 3
rlabel polysilicon 1052 -2105 1052 -2105 0 1
rlabel polysilicon 1052 -2111 1052 -2111 0 3
rlabel polysilicon 1059 -2105 1059 -2105 0 1
rlabel polysilicon 1059 -2111 1059 -2111 0 3
rlabel polysilicon 1066 -2105 1066 -2105 0 1
rlabel polysilicon 1066 -2111 1066 -2111 0 3
rlabel polysilicon 1073 -2105 1073 -2105 0 1
rlabel polysilicon 1073 -2111 1073 -2111 0 3
rlabel polysilicon 1080 -2105 1080 -2105 0 1
rlabel polysilicon 1080 -2111 1080 -2111 0 3
rlabel polysilicon 1087 -2105 1087 -2105 0 1
rlabel polysilicon 1087 -2111 1087 -2111 0 3
rlabel polysilicon 1094 -2105 1094 -2105 0 1
rlabel polysilicon 1094 -2111 1094 -2111 0 3
rlabel polysilicon 1101 -2105 1101 -2105 0 1
rlabel polysilicon 1101 -2111 1101 -2111 0 3
rlabel polysilicon 1108 -2105 1108 -2105 0 1
rlabel polysilicon 1108 -2111 1108 -2111 0 3
rlabel polysilicon 1115 -2105 1115 -2105 0 1
rlabel polysilicon 1115 -2111 1115 -2111 0 3
rlabel polysilicon 1118 -2111 1118 -2111 0 4
rlabel polysilicon 1122 -2105 1122 -2105 0 1
rlabel polysilicon 1122 -2111 1122 -2111 0 3
rlabel polysilicon 1129 -2105 1129 -2105 0 1
rlabel polysilicon 1129 -2111 1129 -2111 0 3
rlabel polysilicon 1139 -2105 1139 -2105 0 2
rlabel polysilicon 1136 -2111 1136 -2111 0 3
rlabel polysilicon 1139 -2111 1139 -2111 0 4
rlabel polysilicon 1143 -2105 1143 -2105 0 1
rlabel polysilicon 1143 -2111 1143 -2111 0 3
rlabel polysilicon 1150 -2105 1150 -2105 0 1
rlabel polysilicon 1150 -2111 1150 -2111 0 3
rlabel polysilicon 1157 -2105 1157 -2105 0 1
rlabel polysilicon 1157 -2111 1157 -2111 0 3
rlabel polysilicon 1164 -2105 1164 -2105 0 1
rlabel polysilicon 1164 -2111 1164 -2111 0 3
rlabel polysilicon 1171 -2105 1171 -2105 0 1
rlabel polysilicon 1171 -2111 1171 -2111 0 3
rlabel polysilicon 1178 -2105 1178 -2105 0 1
rlabel polysilicon 1178 -2111 1178 -2111 0 3
rlabel polysilicon 1185 -2105 1185 -2105 0 1
rlabel polysilicon 1185 -2111 1185 -2111 0 3
rlabel polysilicon 1192 -2105 1192 -2105 0 1
rlabel polysilicon 1192 -2111 1192 -2111 0 3
rlabel polysilicon 1199 -2105 1199 -2105 0 1
rlabel polysilicon 1199 -2111 1199 -2111 0 3
rlabel polysilicon 1206 -2105 1206 -2105 0 1
rlabel polysilicon 1206 -2111 1206 -2111 0 3
rlabel polysilicon 1213 -2105 1213 -2105 0 1
rlabel polysilicon 1213 -2111 1213 -2111 0 3
rlabel polysilicon 1220 -2105 1220 -2105 0 1
rlabel polysilicon 1220 -2111 1220 -2111 0 3
rlabel polysilicon 1227 -2105 1227 -2105 0 1
rlabel polysilicon 1227 -2111 1227 -2111 0 3
rlabel polysilicon 1234 -2105 1234 -2105 0 1
rlabel polysilicon 1234 -2111 1234 -2111 0 3
rlabel polysilicon 1241 -2105 1241 -2105 0 1
rlabel polysilicon 1241 -2111 1241 -2111 0 3
rlabel polysilicon 1248 -2105 1248 -2105 0 1
rlabel polysilicon 1248 -2111 1248 -2111 0 3
rlabel polysilicon 1255 -2105 1255 -2105 0 1
rlabel polysilicon 1255 -2111 1255 -2111 0 3
rlabel polysilicon 1262 -2105 1262 -2105 0 1
rlabel polysilicon 1262 -2111 1262 -2111 0 3
rlabel polysilicon 1269 -2105 1269 -2105 0 1
rlabel polysilicon 1269 -2111 1269 -2111 0 3
rlabel polysilicon 1276 -2105 1276 -2105 0 1
rlabel polysilicon 1276 -2111 1276 -2111 0 3
rlabel polysilicon 1283 -2105 1283 -2105 0 1
rlabel polysilicon 1283 -2111 1283 -2111 0 3
rlabel polysilicon 1290 -2105 1290 -2105 0 1
rlabel polysilicon 1290 -2111 1290 -2111 0 3
rlabel polysilicon 1297 -2105 1297 -2105 0 1
rlabel polysilicon 1297 -2111 1297 -2111 0 3
rlabel polysilicon 1304 -2105 1304 -2105 0 1
rlabel polysilicon 1304 -2111 1304 -2111 0 3
rlabel polysilicon 1311 -2105 1311 -2105 0 1
rlabel polysilicon 1311 -2111 1311 -2111 0 3
rlabel polysilicon 1318 -2105 1318 -2105 0 1
rlabel polysilicon 1318 -2111 1318 -2111 0 3
rlabel polysilicon 1325 -2105 1325 -2105 0 1
rlabel polysilicon 1325 -2111 1325 -2111 0 3
rlabel polysilicon 2 -2238 2 -2238 0 1
rlabel polysilicon 2 -2244 2 -2244 0 3
rlabel polysilicon 9 -2238 9 -2238 0 1
rlabel polysilicon 9 -2244 9 -2244 0 3
rlabel polysilicon 16 -2238 16 -2238 0 1
rlabel polysilicon 16 -2244 16 -2244 0 3
rlabel polysilicon 23 -2238 23 -2238 0 1
rlabel polysilicon 26 -2238 26 -2238 0 2
rlabel polysilicon 23 -2244 23 -2244 0 3
rlabel polysilicon 30 -2244 30 -2244 0 3
rlabel polysilicon 33 -2244 33 -2244 0 4
rlabel polysilicon 37 -2238 37 -2238 0 1
rlabel polysilicon 40 -2238 40 -2238 0 2
rlabel polysilicon 37 -2244 37 -2244 0 3
rlabel polysilicon 40 -2244 40 -2244 0 4
rlabel polysilicon 44 -2238 44 -2238 0 1
rlabel polysilicon 44 -2244 44 -2244 0 3
rlabel polysilicon 51 -2238 51 -2238 0 1
rlabel polysilicon 51 -2244 51 -2244 0 3
rlabel polysilicon 58 -2238 58 -2238 0 1
rlabel polysilicon 58 -2244 58 -2244 0 3
rlabel polysilicon 65 -2238 65 -2238 0 1
rlabel polysilicon 65 -2244 65 -2244 0 3
rlabel polysilicon 72 -2238 72 -2238 0 1
rlabel polysilicon 75 -2238 75 -2238 0 2
rlabel polysilicon 72 -2244 72 -2244 0 3
rlabel polysilicon 75 -2244 75 -2244 0 4
rlabel polysilicon 79 -2238 79 -2238 0 1
rlabel polysilicon 79 -2244 79 -2244 0 3
rlabel polysilicon 86 -2238 86 -2238 0 1
rlabel polysilicon 86 -2244 86 -2244 0 3
rlabel polysilicon 93 -2238 93 -2238 0 1
rlabel polysilicon 93 -2244 93 -2244 0 3
rlabel polysilicon 100 -2238 100 -2238 0 1
rlabel polysilicon 100 -2244 100 -2244 0 3
rlabel polysilicon 107 -2238 107 -2238 0 1
rlabel polysilicon 107 -2244 107 -2244 0 3
rlabel polysilicon 117 -2238 117 -2238 0 2
rlabel polysilicon 114 -2244 114 -2244 0 3
rlabel polysilicon 117 -2244 117 -2244 0 4
rlabel polysilicon 121 -2238 121 -2238 0 1
rlabel polysilicon 121 -2244 121 -2244 0 3
rlabel polysilicon 128 -2238 128 -2238 0 1
rlabel polysilicon 128 -2244 128 -2244 0 3
rlabel polysilicon 135 -2238 135 -2238 0 1
rlabel polysilicon 138 -2238 138 -2238 0 2
rlabel polysilicon 135 -2244 135 -2244 0 3
rlabel polysilicon 138 -2244 138 -2244 0 4
rlabel polysilicon 142 -2238 142 -2238 0 1
rlabel polysilicon 142 -2244 142 -2244 0 3
rlabel polysilicon 149 -2238 149 -2238 0 1
rlabel polysilicon 152 -2238 152 -2238 0 2
rlabel polysilicon 149 -2244 149 -2244 0 3
rlabel polysilicon 156 -2238 156 -2238 0 1
rlabel polysilicon 156 -2244 156 -2244 0 3
rlabel polysilicon 163 -2238 163 -2238 0 1
rlabel polysilicon 163 -2244 163 -2244 0 3
rlabel polysilicon 170 -2238 170 -2238 0 1
rlabel polysilicon 170 -2244 170 -2244 0 3
rlabel polysilicon 177 -2238 177 -2238 0 1
rlabel polysilicon 177 -2244 177 -2244 0 3
rlabel polysilicon 184 -2238 184 -2238 0 1
rlabel polysilicon 184 -2244 184 -2244 0 3
rlabel polysilicon 191 -2238 191 -2238 0 1
rlabel polysilicon 191 -2244 191 -2244 0 3
rlabel polysilicon 198 -2238 198 -2238 0 1
rlabel polysilicon 198 -2244 198 -2244 0 3
rlabel polysilicon 205 -2238 205 -2238 0 1
rlabel polysilicon 205 -2244 205 -2244 0 3
rlabel polysilicon 212 -2238 212 -2238 0 1
rlabel polysilicon 212 -2244 212 -2244 0 3
rlabel polysilicon 219 -2238 219 -2238 0 1
rlabel polysilicon 219 -2244 219 -2244 0 3
rlabel polysilicon 226 -2238 226 -2238 0 1
rlabel polysilicon 226 -2244 226 -2244 0 3
rlabel polysilicon 233 -2244 233 -2244 0 3
rlabel polysilicon 240 -2238 240 -2238 0 1
rlabel polysilicon 240 -2244 240 -2244 0 3
rlabel polysilicon 247 -2238 247 -2238 0 1
rlabel polysilicon 247 -2244 247 -2244 0 3
rlabel polysilicon 254 -2238 254 -2238 0 1
rlabel polysilicon 254 -2244 254 -2244 0 3
rlabel polysilicon 261 -2238 261 -2238 0 1
rlabel polysilicon 261 -2244 261 -2244 0 3
rlabel polysilicon 268 -2238 268 -2238 0 1
rlabel polysilicon 268 -2244 268 -2244 0 3
rlabel polysilicon 275 -2238 275 -2238 0 1
rlabel polysilicon 275 -2244 275 -2244 0 3
rlabel polysilicon 282 -2238 282 -2238 0 1
rlabel polysilicon 282 -2244 282 -2244 0 3
rlabel polysilicon 289 -2238 289 -2238 0 1
rlabel polysilicon 289 -2244 289 -2244 0 3
rlabel polysilicon 296 -2238 296 -2238 0 1
rlabel polysilicon 299 -2238 299 -2238 0 2
rlabel polysilicon 296 -2244 296 -2244 0 3
rlabel polysilicon 299 -2244 299 -2244 0 4
rlabel polysilicon 303 -2238 303 -2238 0 1
rlabel polysilicon 303 -2244 303 -2244 0 3
rlabel polysilicon 310 -2238 310 -2238 0 1
rlabel polysilicon 310 -2244 310 -2244 0 3
rlabel polysilicon 317 -2238 317 -2238 0 1
rlabel polysilicon 317 -2244 317 -2244 0 3
rlabel polysilicon 324 -2238 324 -2238 0 1
rlabel polysilicon 324 -2244 324 -2244 0 3
rlabel polysilicon 331 -2238 331 -2238 0 1
rlabel polysilicon 331 -2244 331 -2244 0 3
rlabel polysilicon 338 -2238 338 -2238 0 1
rlabel polysilicon 338 -2244 338 -2244 0 3
rlabel polysilicon 341 -2244 341 -2244 0 4
rlabel polysilicon 345 -2238 345 -2238 0 1
rlabel polysilicon 345 -2244 345 -2244 0 3
rlabel polysilicon 352 -2238 352 -2238 0 1
rlabel polysilicon 352 -2244 352 -2244 0 3
rlabel polysilicon 359 -2238 359 -2238 0 1
rlabel polysilicon 359 -2244 359 -2244 0 3
rlabel polysilicon 366 -2238 366 -2238 0 1
rlabel polysilicon 366 -2244 366 -2244 0 3
rlabel polysilicon 373 -2238 373 -2238 0 1
rlabel polysilicon 373 -2244 373 -2244 0 3
rlabel polysilicon 380 -2238 380 -2238 0 1
rlabel polysilicon 380 -2244 380 -2244 0 3
rlabel polysilicon 387 -2238 387 -2238 0 1
rlabel polysilicon 387 -2244 387 -2244 0 3
rlabel polysilicon 394 -2238 394 -2238 0 1
rlabel polysilicon 397 -2238 397 -2238 0 2
rlabel polysilicon 394 -2244 394 -2244 0 3
rlabel polysilicon 397 -2244 397 -2244 0 4
rlabel polysilicon 401 -2238 401 -2238 0 1
rlabel polysilicon 404 -2238 404 -2238 0 2
rlabel polysilicon 401 -2244 401 -2244 0 3
rlabel polysilicon 404 -2244 404 -2244 0 4
rlabel polysilicon 408 -2238 408 -2238 0 1
rlabel polysilicon 411 -2238 411 -2238 0 2
rlabel polysilicon 408 -2244 408 -2244 0 3
rlabel polysilicon 411 -2244 411 -2244 0 4
rlabel polysilicon 415 -2238 415 -2238 0 1
rlabel polysilicon 415 -2244 415 -2244 0 3
rlabel polysilicon 425 -2238 425 -2238 0 2
rlabel polysilicon 422 -2244 422 -2244 0 3
rlabel polysilicon 425 -2244 425 -2244 0 4
rlabel polysilicon 429 -2238 429 -2238 0 1
rlabel polysilicon 429 -2244 429 -2244 0 3
rlabel polysilicon 436 -2238 436 -2238 0 1
rlabel polysilicon 436 -2244 436 -2244 0 3
rlabel polysilicon 443 -2238 443 -2238 0 1
rlabel polysilicon 443 -2244 443 -2244 0 3
rlabel polysilicon 450 -2238 450 -2238 0 1
rlabel polysilicon 453 -2238 453 -2238 0 2
rlabel polysilicon 450 -2244 450 -2244 0 3
rlabel polysilicon 453 -2244 453 -2244 0 4
rlabel polysilicon 457 -2238 457 -2238 0 1
rlabel polysilicon 457 -2244 457 -2244 0 3
rlabel polysilicon 464 -2238 464 -2238 0 1
rlabel polysilicon 464 -2244 464 -2244 0 3
rlabel polysilicon 471 -2238 471 -2238 0 1
rlabel polysilicon 471 -2244 471 -2244 0 3
rlabel polysilicon 478 -2238 478 -2238 0 1
rlabel polysilicon 478 -2244 478 -2244 0 3
rlabel polysilicon 485 -2238 485 -2238 0 1
rlabel polysilicon 485 -2244 485 -2244 0 3
rlabel polysilicon 492 -2238 492 -2238 0 1
rlabel polysilicon 492 -2244 492 -2244 0 3
rlabel polysilicon 499 -2238 499 -2238 0 1
rlabel polysilicon 499 -2244 499 -2244 0 3
rlabel polysilicon 506 -2238 506 -2238 0 1
rlabel polysilicon 506 -2244 506 -2244 0 3
rlabel polysilicon 513 -2238 513 -2238 0 1
rlabel polysilicon 513 -2244 513 -2244 0 3
rlabel polysilicon 520 -2238 520 -2238 0 1
rlabel polysilicon 523 -2238 523 -2238 0 2
rlabel polysilicon 520 -2244 520 -2244 0 3
rlabel polysilicon 523 -2244 523 -2244 0 4
rlabel polysilicon 527 -2238 527 -2238 0 1
rlabel polysilicon 530 -2238 530 -2238 0 2
rlabel polysilicon 527 -2244 527 -2244 0 3
rlabel polysilicon 530 -2244 530 -2244 0 4
rlabel polysilicon 534 -2238 534 -2238 0 1
rlabel polysilicon 534 -2244 534 -2244 0 3
rlabel polysilicon 541 -2238 541 -2238 0 1
rlabel polysilicon 541 -2244 541 -2244 0 3
rlabel polysilicon 548 -2238 548 -2238 0 1
rlabel polysilicon 548 -2244 548 -2244 0 3
rlabel polysilicon 555 -2238 555 -2238 0 1
rlabel polysilicon 555 -2244 555 -2244 0 3
rlabel polysilicon 558 -2244 558 -2244 0 4
rlabel polysilicon 562 -2238 562 -2238 0 1
rlabel polysilicon 562 -2244 562 -2244 0 3
rlabel polysilicon 569 -2238 569 -2238 0 1
rlabel polysilicon 569 -2244 569 -2244 0 3
rlabel polysilicon 576 -2238 576 -2238 0 1
rlabel polysilicon 576 -2244 576 -2244 0 3
rlabel polysilicon 583 -2238 583 -2238 0 1
rlabel polysilicon 583 -2244 583 -2244 0 3
rlabel polysilicon 590 -2238 590 -2238 0 1
rlabel polysilicon 590 -2244 590 -2244 0 3
rlabel polysilicon 597 -2238 597 -2238 0 1
rlabel polysilicon 597 -2244 597 -2244 0 3
rlabel polysilicon 604 -2238 604 -2238 0 1
rlabel polysilicon 604 -2244 604 -2244 0 3
rlabel polysilicon 611 -2238 611 -2238 0 1
rlabel polysilicon 611 -2244 611 -2244 0 3
rlabel polysilicon 618 -2238 618 -2238 0 1
rlabel polysilicon 621 -2238 621 -2238 0 2
rlabel polysilicon 618 -2244 618 -2244 0 3
rlabel polysilicon 621 -2244 621 -2244 0 4
rlabel polysilicon 625 -2238 625 -2238 0 1
rlabel polysilicon 628 -2238 628 -2238 0 2
rlabel polysilicon 628 -2244 628 -2244 0 4
rlabel polysilicon 632 -2238 632 -2238 0 1
rlabel polysilicon 632 -2244 632 -2244 0 3
rlabel polysilicon 639 -2238 639 -2238 0 1
rlabel polysilicon 639 -2244 639 -2244 0 3
rlabel polysilicon 646 -2238 646 -2238 0 1
rlabel polysilicon 649 -2238 649 -2238 0 2
rlabel polysilicon 646 -2244 646 -2244 0 3
rlabel polysilicon 653 -2238 653 -2238 0 1
rlabel polysilicon 653 -2244 653 -2244 0 3
rlabel polysilicon 660 -2238 660 -2238 0 1
rlabel polysilicon 660 -2244 660 -2244 0 3
rlabel polysilicon 667 -2238 667 -2238 0 1
rlabel polysilicon 667 -2244 667 -2244 0 3
rlabel polysilicon 677 -2238 677 -2238 0 2
rlabel polysilicon 677 -2244 677 -2244 0 4
rlabel polysilicon 681 -2238 681 -2238 0 1
rlabel polysilicon 681 -2244 681 -2244 0 3
rlabel polysilicon 688 -2238 688 -2238 0 1
rlabel polysilicon 688 -2244 688 -2244 0 3
rlabel polysilicon 695 -2238 695 -2238 0 1
rlabel polysilicon 695 -2244 695 -2244 0 3
rlabel polysilicon 702 -2238 702 -2238 0 1
rlabel polysilicon 702 -2244 702 -2244 0 3
rlabel polysilicon 709 -2238 709 -2238 0 1
rlabel polysilicon 709 -2244 709 -2244 0 3
rlabel polysilicon 716 -2238 716 -2238 0 1
rlabel polysilicon 716 -2244 716 -2244 0 3
rlabel polysilicon 723 -2238 723 -2238 0 1
rlabel polysilicon 723 -2244 723 -2244 0 3
rlabel polysilicon 730 -2238 730 -2238 0 1
rlabel polysilicon 730 -2244 730 -2244 0 3
rlabel polysilicon 737 -2238 737 -2238 0 1
rlabel polysilicon 737 -2244 737 -2244 0 3
rlabel polysilicon 744 -2238 744 -2238 0 1
rlabel polysilicon 744 -2244 744 -2244 0 3
rlabel polysilicon 751 -2238 751 -2238 0 1
rlabel polysilicon 751 -2244 751 -2244 0 3
rlabel polysilicon 758 -2238 758 -2238 0 1
rlabel polysilicon 758 -2244 758 -2244 0 3
rlabel polysilicon 765 -2238 765 -2238 0 1
rlabel polysilicon 768 -2238 768 -2238 0 2
rlabel polysilicon 765 -2244 765 -2244 0 3
rlabel polysilicon 772 -2238 772 -2238 0 1
rlabel polysilicon 772 -2244 772 -2244 0 3
rlabel polysilicon 779 -2238 779 -2238 0 1
rlabel polysilicon 779 -2244 779 -2244 0 3
rlabel polysilicon 786 -2238 786 -2238 0 1
rlabel polysilicon 786 -2244 786 -2244 0 3
rlabel polysilicon 793 -2238 793 -2238 0 1
rlabel polysilicon 793 -2244 793 -2244 0 3
rlabel polysilicon 800 -2238 800 -2238 0 1
rlabel polysilicon 800 -2244 800 -2244 0 3
rlabel polysilicon 807 -2238 807 -2238 0 1
rlabel polysilicon 810 -2238 810 -2238 0 2
rlabel polysilicon 807 -2244 807 -2244 0 3
rlabel polysilicon 810 -2244 810 -2244 0 4
rlabel polysilicon 814 -2238 814 -2238 0 1
rlabel polysilicon 814 -2244 814 -2244 0 3
rlabel polysilicon 821 -2238 821 -2238 0 1
rlabel polysilicon 821 -2244 821 -2244 0 3
rlabel polysilicon 828 -2238 828 -2238 0 1
rlabel polysilicon 828 -2244 828 -2244 0 3
rlabel polysilicon 835 -2238 835 -2238 0 1
rlabel polysilicon 835 -2244 835 -2244 0 3
rlabel polysilicon 842 -2238 842 -2238 0 1
rlabel polysilicon 842 -2244 842 -2244 0 3
rlabel polysilicon 849 -2238 849 -2238 0 1
rlabel polysilicon 849 -2244 849 -2244 0 3
rlabel polysilicon 856 -2238 856 -2238 0 1
rlabel polysilicon 856 -2244 856 -2244 0 3
rlabel polysilicon 863 -2238 863 -2238 0 1
rlabel polysilicon 863 -2244 863 -2244 0 3
rlabel polysilicon 870 -2238 870 -2238 0 1
rlabel polysilicon 870 -2244 870 -2244 0 3
rlabel polysilicon 873 -2244 873 -2244 0 4
rlabel polysilicon 877 -2238 877 -2238 0 1
rlabel polysilicon 877 -2244 877 -2244 0 3
rlabel polysilicon 884 -2238 884 -2238 0 1
rlabel polysilicon 884 -2244 884 -2244 0 3
rlabel polysilicon 891 -2238 891 -2238 0 1
rlabel polysilicon 891 -2244 891 -2244 0 3
rlabel polysilicon 898 -2238 898 -2238 0 1
rlabel polysilicon 898 -2244 898 -2244 0 3
rlabel polysilicon 905 -2238 905 -2238 0 1
rlabel polysilicon 905 -2244 905 -2244 0 3
rlabel polysilicon 912 -2238 912 -2238 0 1
rlabel polysilicon 912 -2244 912 -2244 0 3
rlabel polysilicon 919 -2238 919 -2238 0 1
rlabel polysilicon 919 -2244 919 -2244 0 3
rlabel polysilicon 926 -2238 926 -2238 0 1
rlabel polysilicon 926 -2244 926 -2244 0 3
rlabel polysilicon 933 -2238 933 -2238 0 1
rlabel polysilicon 936 -2238 936 -2238 0 2
rlabel polysilicon 933 -2244 933 -2244 0 3
rlabel polysilicon 940 -2238 940 -2238 0 1
rlabel polysilicon 940 -2244 940 -2244 0 3
rlabel polysilicon 947 -2238 947 -2238 0 1
rlabel polysilicon 947 -2244 947 -2244 0 3
rlabel polysilicon 954 -2238 954 -2238 0 1
rlabel polysilicon 954 -2244 954 -2244 0 3
rlabel polysilicon 961 -2238 961 -2238 0 1
rlabel polysilicon 961 -2244 961 -2244 0 3
rlabel polysilicon 968 -2238 968 -2238 0 1
rlabel polysilicon 968 -2244 968 -2244 0 3
rlabel polysilicon 975 -2238 975 -2238 0 1
rlabel polysilicon 975 -2244 975 -2244 0 3
rlabel polysilicon 982 -2238 982 -2238 0 1
rlabel polysilicon 985 -2238 985 -2238 0 2
rlabel polysilicon 982 -2244 982 -2244 0 3
rlabel polysilicon 985 -2244 985 -2244 0 4
rlabel polysilicon 989 -2238 989 -2238 0 1
rlabel polysilicon 989 -2244 989 -2244 0 3
rlabel polysilicon 996 -2238 996 -2238 0 1
rlabel polysilicon 996 -2244 996 -2244 0 3
rlabel polysilicon 1003 -2238 1003 -2238 0 1
rlabel polysilicon 1003 -2244 1003 -2244 0 3
rlabel polysilicon 1010 -2238 1010 -2238 0 1
rlabel polysilicon 1010 -2244 1010 -2244 0 3
rlabel polysilicon 1017 -2238 1017 -2238 0 1
rlabel polysilicon 1017 -2244 1017 -2244 0 3
rlabel polysilicon 1024 -2238 1024 -2238 0 1
rlabel polysilicon 1024 -2244 1024 -2244 0 3
rlabel polysilicon 1031 -2238 1031 -2238 0 1
rlabel polysilicon 1031 -2244 1031 -2244 0 3
rlabel polysilicon 1038 -2238 1038 -2238 0 1
rlabel polysilicon 1038 -2244 1038 -2244 0 3
rlabel polysilicon 1045 -2238 1045 -2238 0 1
rlabel polysilicon 1045 -2244 1045 -2244 0 3
rlabel polysilicon 1052 -2238 1052 -2238 0 1
rlabel polysilicon 1052 -2244 1052 -2244 0 3
rlabel polysilicon 1059 -2238 1059 -2238 0 1
rlabel polysilicon 1059 -2244 1059 -2244 0 3
rlabel polysilicon 1066 -2238 1066 -2238 0 1
rlabel polysilicon 1066 -2244 1066 -2244 0 3
rlabel polysilicon 1073 -2238 1073 -2238 0 1
rlabel polysilicon 1073 -2244 1073 -2244 0 3
rlabel polysilicon 1080 -2238 1080 -2238 0 1
rlabel polysilicon 1080 -2244 1080 -2244 0 3
rlabel polysilicon 1087 -2238 1087 -2238 0 1
rlabel polysilicon 1087 -2244 1087 -2244 0 3
rlabel polysilicon 1094 -2238 1094 -2238 0 1
rlabel polysilicon 1094 -2244 1094 -2244 0 3
rlabel polysilicon 1101 -2238 1101 -2238 0 1
rlabel polysilicon 1101 -2244 1101 -2244 0 3
rlabel polysilicon 1108 -2238 1108 -2238 0 1
rlabel polysilicon 1108 -2244 1108 -2244 0 3
rlabel polysilicon 1115 -2238 1115 -2238 0 1
rlabel polysilicon 1115 -2244 1115 -2244 0 3
rlabel polysilicon 1122 -2238 1122 -2238 0 1
rlabel polysilicon 1122 -2244 1122 -2244 0 3
rlabel polysilicon 1129 -2238 1129 -2238 0 1
rlabel polysilicon 1129 -2244 1129 -2244 0 3
rlabel polysilicon 1136 -2238 1136 -2238 0 1
rlabel polysilicon 1136 -2244 1136 -2244 0 3
rlabel polysilicon 1143 -2238 1143 -2238 0 1
rlabel polysilicon 1143 -2244 1143 -2244 0 3
rlabel polysilicon 1150 -2238 1150 -2238 0 1
rlabel polysilicon 1150 -2244 1150 -2244 0 3
rlabel polysilicon 1157 -2238 1157 -2238 0 1
rlabel polysilicon 1157 -2244 1157 -2244 0 3
rlabel polysilicon 1164 -2238 1164 -2238 0 1
rlabel polysilicon 1164 -2244 1164 -2244 0 3
rlabel polysilicon 1171 -2238 1171 -2238 0 1
rlabel polysilicon 1171 -2244 1171 -2244 0 3
rlabel polysilicon 1178 -2238 1178 -2238 0 1
rlabel polysilicon 1178 -2244 1178 -2244 0 3
rlabel polysilicon 1185 -2238 1185 -2238 0 1
rlabel polysilicon 1185 -2244 1185 -2244 0 3
rlabel polysilicon 1192 -2238 1192 -2238 0 1
rlabel polysilicon 1192 -2244 1192 -2244 0 3
rlabel polysilicon 1199 -2238 1199 -2238 0 1
rlabel polysilicon 1199 -2244 1199 -2244 0 3
rlabel polysilicon 1206 -2238 1206 -2238 0 1
rlabel polysilicon 1206 -2244 1206 -2244 0 3
rlabel polysilicon 1213 -2238 1213 -2238 0 1
rlabel polysilicon 1213 -2244 1213 -2244 0 3
rlabel polysilicon 1220 -2238 1220 -2238 0 1
rlabel polysilicon 1220 -2244 1220 -2244 0 3
rlabel polysilicon 1227 -2238 1227 -2238 0 1
rlabel polysilicon 1227 -2244 1227 -2244 0 3
rlabel polysilicon 1234 -2238 1234 -2238 0 1
rlabel polysilicon 1234 -2244 1234 -2244 0 3
rlabel polysilicon 1241 -2238 1241 -2238 0 1
rlabel polysilicon 1241 -2244 1241 -2244 0 3
rlabel polysilicon 1248 -2238 1248 -2238 0 1
rlabel polysilicon 1248 -2244 1248 -2244 0 3
rlabel polysilicon 1255 -2238 1255 -2238 0 1
rlabel polysilicon 1255 -2244 1255 -2244 0 3
rlabel polysilicon 1262 -2238 1262 -2238 0 1
rlabel polysilicon 1262 -2244 1262 -2244 0 3
rlabel polysilicon 1269 -2238 1269 -2238 0 1
rlabel polysilicon 1269 -2244 1269 -2244 0 3
rlabel polysilicon 1276 -2238 1276 -2238 0 1
rlabel polysilicon 1276 -2244 1276 -2244 0 3
rlabel polysilicon 1283 -2238 1283 -2238 0 1
rlabel polysilicon 1283 -2244 1283 -2244 0 3
rlabel polysilicon 1290 -2238 1290 -2238 0 1
rlabel polysilicon 1290 -2244 1290 -2244 0 3
rlabel polysilicon 1297 -2238 1297 -2238 0 1
rlabel polysilicon 1297 -2244 1297 -2244 0 3
rlabel polysilicon 1304 -2238 1304 -2238 0 1
rlabel polysilicon 1304 -2244 1304 -2244 0 3
rlabel polysilicon 1311 -2238 1311 -2238 0 1
rlabel polysilicon 1311 -2244 1311 -2244 0 3
rlabel polysilicon 2 -2363 2 -2363 0 1
rlabel polysilicon 5 -2363 5 -2363 0 2
rlabel polysilicon 9 -2363 9 -2363 0 1
rlabel polysilicon 9 -2369 9 -2369 0 3
rlabel polysilicon 16 -2363 16 -2363 0 1
rlabel polysilicon 16 -2369 16 -2369 0 3
rlabel polysilicon 23 -2363 23 -2363 0 1
rlabel polysilicon 23 -2369 23 -2369 0 3
rlabel polysilicon 30 -2363 30 -2363 0 1
rlabel polysilicon 30 -2369 30 -2369 0 3
rlabel polysilicon 37 -2363 37 -2363 0 1
rlabel polysilicon 40 -2363 40 -2363 0 2
rlabel polysilicon 37 -2369 37 -2369 0 3
rlabel polysilicon 40 -2369 40 -2369 0 4
rlabel polysilicon 44 -2363 44 -2363 0 1
rlabel polysilicon 44 -2369 44 -2369 0 3
rlabel polysilicon 51 -2363 51 -2363 0 1
rlabel polysilicon 51 -2369 51 -2369 0 3
rlabel polysilicon 54 -2369 54 -2369 0 4
rlabel polysilicon 58 -2363 58 -2363 0 1
rlabel polysilicon 61 -2363 61 -2363 0 2
rlabel polysilicon 58 -2369 58 -2369 0 3
rlabel polysilicon 61 -2369 61 -2369 0 4
rlabel polysilicon 65 -2363 65 -2363 0 1
rlabel polysilicon 65 -2369 65 -2369 0 3
rlabel polysilicon 72 -2363 72 -2363 0 1
rlabel polysilicon 72 -2369 72 -2369 0 3
rlabel polysilicon 79 -2363 79 -2363 0 1
rlabel polysilicon 79 -2369 79 -2369 0 3
rlabel polysilicon 86 -2363 86 -2363 0 1
rlabel polysilicon 86 -2369 86 -2369 0 3
rlabel polysilicon 93 -2363 93 -2363 0 1
rlabel polysilicon 96 -2363 96 -2363 0 2
rlabel polysilicon 93 -2369 93 -2369 0 3
rlabel polysilicon 100 -2363 100 -2363 0 1
rlabel polysilicon 100 -2369 100 -2369 0 3
rlabel polysilicon 107 -2363 107 -2363 0 1
rlabel polysilicon 107 -2369 107 -2369 0 3
rlabel polysilicon 114 -2363 114 -2363 0 1
rlabel polysilicon 114 -2369 114 -2369 0 3
rlabel polysilicon 121 -2363 121 -2363 0 1
rlabel polysilicon 121 -2369 121 -2369 0 3
rlabel polysilicon 128 -2363 128 -2363 0 1
rlabel polysilicon 128 -2369 128 -2369 0 3
rlabel polysilicon 135 -2363 135 -2363 0 1
rlabel polysilicon 138 -2363 138 -2363 0 2
rlabel polysilicon 135 -2369 135 -2369 0 3
rlabel polysilicon 138 -2369 138 -2369 0 4
rlabel polysilicon 142 -2363 142 -2363 0 1
rlabel polysilicon 142 -2369 142 -2369 0 3
rlabel polysilicon 149 -2363 149 -2363 0 1
rlabel polysilicon 152 -2363 152 -2363 0 2
rlabel polysilicon 156 -2363 156 -2363 0 1
rlabel polysilicon 156 -2369 156 -2369 0 3
rlabel polysilicon 163 -2363 163 -2363 0 1
rlabel polysilicon 163 -2369 163 -2369 0 3
rlabel polysilicon 170 -2363 170 -2363 0 1
rlabel polysilicon 170 -2369 170 -2369 0 3
rlabel polysilicon 177 -2363 177 -2363 0 1
rlabel polysilicon 177 -2369 177 -2369 0 3
rlabel polysilicon 184 -2363 184 -2363 0 1
rlabel polysilicon 184 -2369 184 -2369 0 3
rlabel polysilicon 191 -2363 191 -2363 0 1
rlabel polysilicon 191 -2369 191 -2369 0 3
rlabel polysilicon 198 -2363 198 -2363 0 1
rlabel polysilicon 198 -2369 198 -2369 0 3
rlabel polysilicon 205 -2363 205 -2363 0 1
rlabel polysilicon 205 -2369 205 -2369 0 3
rlabel polysilicon 212 -2363 212 -2363 0 1
rlabel polysilicon 212 -2369 212 -2369 0 3
rlabel polysilicon 219 -2363 219 -2363 0 1
rlabel polysilicon 219 -2369 219 -2369 0 3
rlabel polysilicon 226 -2363 226 -2363 0 1
rlabel polysilicon 226 -2369 226 -2369 0 3
rlabel polysilicon 233 -2363 233 -2363 0 1
rlabel polysilicon 233 -2369 233 -2369 0 3
rlabel polysilicon 240 -2363 240 -2363 0 1
rlabel polysilicon 240 -2369 240 -2369 0 3
rlabel polysilicon 247 -2363 247 -2363 0 1
rlabel polysilicon 247 -2369 247 -2369 0 3
rlabel polysilicon 254 -2363 254 -2363 0 1
rlabel polysilicon 254 -2369 254 -2369 0 3
rlabel polysilicon 261 -2363 261 -2363 0 1
rlabel polysilicon 261 -2369 261 -2369 0 3
rlabel polysilicon 268 -2363 268 -2363 0 1
rlabel polysilicon 268 -2369 268 -2369 0 3
rlabel polysilicon 275 -2363 275 -2363 0 1
rlabel polysilicon 275 -2369 275 -2369 0 3
rlabel polysilicon 282 -2363 282 -2363 0 1
rlabel polysilicon 282 -2369 282 -2369 0 3
rlabel polysilicon 289 -2363 289 -2363 0 1
rlabel polysilicon 289 -2369 289 -2369 0 3
rlabel polysilicon 296 -2363 296 -2363 0 1
rlabel polysilicon 296 -2369 296 -2369 0 3
rlabel polysilicon 306 -2363 306 -2363 0 2
rlabel polysilicon 303 -2369 303 -2369 0 3
rlabel polysilicon 306 -2369 306 -2369 0 4
rlabel polysilicon 310 -2363 310 -2363 0 1
rlabel polysilicon 310 -2369 310 -2369 0 3
rlabel polysilicon 317 -2363 317 -2363 0 1
rlabel polysilicon 320 -2363 320 -2363 0 2
rlabel polysilicon 317 -2369 317 -2369 0 3
rlabel polysilicon 320 -2369 320 -2369 0 4
rlabel polysilicon 324 -2363 324 -2363 0 1
rlabel polysilicon 324 -2369 324 -2369 0 3
rlabel polysilicon 331 -2363 331 -2363 0 1
rlabel polysilicon 331 -2369 331 -2369 0 3
rlabel polysilicon 338 -2363 338 -2363 0 1
rlabel polysilicon 341 -2363 341 -2363 0 2
rlabel polysilicon 341 -2369 341 -2369 0 4
rlabel polysilicon 345 -2363 345 -2363 0 1
rlabel polysilicon 345 -2369 345 -2369 0 3
rlabel polysilicon 352 -2363 352 -2363 0 1
rlabel polysilicon 352 -2369 352 -2369 0 3
rlabel polysilicon 359 -2363 359 -2363 0 1
rlabel polysilicon 359 -2369 359 -2369 0 3
rlabel polysilicon 366 -2363 366 -2363 0 1
rlabel polysilicon 366 -2369 366 -2369 0 3
rlabel polysilicon 373 -2363 373 -2363 0 1
rlabel polysilicon 373 -2369 373 -2369 0 3
rlabel polysilicon 380 -2363 380 -2363 0 1
rlabel polysilicon 380 -2369 380 -2369 0 3
rlabel polysilicon 387 -2363 387 -2363 0 1
rlabel polysilicon 387 -2369 387 -2369 0 3
rlabel polysilicon 394 -2363 394 -2363 0 1
rlabel polysilicon 397 -2363 397 -2363 0 2
rlabel polysilicon 394 -2369 394 -2369 0 3
rlabel polysilicon 397 -2369 397 -2369 0 4
rlabel polysilicon 401 -2363 401 -2363 0 1
rlabel polysilicon 401 -2369 401 -2369 0 3
rlabel polysilicon 408 -2363 408 -2363 0 1
rlabel polysilicon 408 -2369 408 -2369 0 3
rlabel polysilicon 415 -2363 415 -2363 0 1
rlabel polysilicon 415 -2369 415 -2369 0 3
rlabel polysilicon 425 -2363 425 -2363 0 2
rlabel polysilicon 422 -2369 422 -2369 0 3
rlabel polysilicon 425 -2369 425 -2369 0 4
rlabel polysilicon 429 -2363 429 -2363 0 1
rlabel polysilicon 429 -2369 429 -2369 0 3
rlabel polysilicon 436 -2363 436 -2363 0 1
rlabel polysilicon 436 -2369 436 -2369 0 3
rlabel polysilicon 439 -2369 439 -2369 0 4
rlabel polysilicon 443 -2363 443 -2363 0 1
rlabel polysilicon 443 -2369 443 -2369 0 3
rlabel polysilicon 450 -2363 450 -2363 0 1
rlabel polysilicon 450 -2369 450 -2369 0 3
rlabel polysilicon 457 -2363 457 -2363 0 1
rlabel polysilicon 457 -2369 457 -2369 0 3
rlabel polysilicon 464 -2363 464 -2363 0 1
rlabel polysilicon 464 -2369 464 -2369 0 3
rlabel polysilicon 471 -2363 471 -2363 0 1
rlabel polysilicon 471 -2369 471 -2369 0 3
rlabel polysilicon 478 -2363 478 -2363 0 1
rlabel polysilicon 478 -2369 478 -2369 0 3
rlabel polysilicon 485 -2363 485 -2363 0 1
rlabel polysilicon 485 -2369 485 -2369 0 3
rlabel polysilicon 492 -2363 492 -2363 0 1
rlabel polysilicon 492 -2369 492 -2369 0 3
rlabel polysilicon 499 -2363 499 -2363 0 1
rlabel polysilicon 499 -2369 499 -2369 0 3
rlabel polysilicon 506 -2363 506 -2363 0 1
rlabel polysilicon 506 -2369 506 -2369 0 3
rlabel polysilicon 513 -2363 513 -2363 0 1
rlabel polysilicon 516 -2363 516 -2363 0 2
rlabel polysilicon 513 -2369 513 -2369 0 3
rlabel polysilicon 516 -2369 516 -2369 0 4
rlabel polysilicon 520 -2363 520 -2363 0 1
rlabel polysilicon 520 -2369 520 -2369 0 3
rlabel polysilicon 527 -2363 527 -2363 0 1
rlabel polysilicon 527 -2369 527 -2369 0 3
rlabel polysilicon 534 -2363 534 -2363 0 1
rlabel polysilicon 534 -2369 534 -2369 0 3
rlabel polysilicon 541 -2363 541 -2363 0 1
rlabel polysilicon 541 -2369 541 -2369 0 3
rlabel polysilicon 548 -2363 548 -2363 0 1
rlabel polysilicon 548 -2369 548 -2369 0 3
rlabel polysilicon 555 -2363 555 -2363 0 1
rlabel polysilicon 558 -2369 558 -2369 0 4
rlabel polysilicon 562 -2363 562 -2363 0 1
rlabel polysilicon 562 -2369 562 -2369 0 3
rlabel polysilicon 569 -2363 569 -2363 0 1
rlabel polysilicon 569 -2369 569 -2369 0 3
rlabel polysilicon 576 -2363 576 -2363 0 1
rlabel polysilicon 579 -2363 579 -2363 0 2
rlabel polysilicon 576 -2369 576 -2369 0 3
rlabel polysilicon 579 -2369 579 -2369 0 4
rlabel polysilicon 583 -2363 583 -2363 0 1
rlabel polysilicon 583 -2369 583 -2369 0 3
rlabel polysilicon 590 -2363 590 -2363 0 1
rlabel polysilicon 593 -2363 593 -2363 0 2
rlabel polysilicon 590 -2369 590 -2369 0 3
rlabel polysilicon 593 -2369 593 -2369 0 4
rlabel polysilicon 597 -2363 597 -2363 0 1
rlabel polysilicon 597 -2369 597 -2369 0 3
rlabel polysilicon 604 -2363 604 -2363 0 1
rlabel polysilicon 604 -2369 604 -2369 0 3
rlabel polysilicon 611 -2363 611 -2363 0 1
rlabel polysilicon 611 -2369 611 -2369 0 3
rlabel polysilicon 618 -2363 618 -2363 0 1
rlabel polysilicon 618 -2369 618 -2369 0 3
rlabel polysilicon 625 -2363 625 -2363 0 1
rlabel polysilicon 625 -2369 625 -2369 0 3
rlabel polysilicon 632 -2363 632 -2363 0 1
rlabel polysilicon 635 -2363 635 -2363 0 2
rlabel polysilicon 632 -2369 632 -2369 0 3
rlabel polysilicon 635 -2369 635 -2369 0 4
rlabel polysilicon 639 -2363 639 -2363 0 1
rlabel polysilicon 639 -2369 639 -2369 0 3
rlabel polysilicon 646 -2363 646 -2363 0 1
rlabel polysilicon 646 -2369 646 -2369 0 3
rlabel polysilicon 653 -2363 653 -2363 0 1
rlabel polysilicon 653 -2369 653 -2369 0 3
rlabel polysilicon 660 -2363 660 -2363 0 1
rlabel polysilicon 663 -2363 663 -2363 0 2
rlabel polysilicon 660 -2369 660 -2369 0 3
rlabel polysilicon 667 -2363 667 -2363 0 1
rlabel polysilicon 667 -2369 667 -2369 0 3
rlabel polysilicon 674 -2363 674 -2363 0 1
rlabel polysilicon 674 -2369 674 -2369 0 3
rlabel polysilicon 681 -2363 681 -2363 0 1
rlabel polysilicon 681 -2369 681 -2369 0 3
rlabel polysilicon 688 -2363 688 -2363 0 1
rlabel polysilicon 688 -2369 688 -2369 0 3
rlabel polysilicon 695 -2363 695 -2363 0 1
rlabel polysilicon 695 -2369 695 -2369 0 3
rlabel polysilicon 702 -2363 702 -2363 0 1
rlabel polysilicon 702 -2369 702 -2369 0 3
rlabel polysilicon 709 -2363 709 -2363 0 1
rlabel polysilicon 709 -2369 709 -2369 0 3
rlabel polysilicon 716 -2363 716 -2363 0 1
rlabel polysilicon 716 -2369 716 -2369 0 3
rlabel polysilicon 726 -2363 726 -2363 0 2
rlabel polysilicon 723 -2369 723 -2369 0 3
rlabel polysilicon 726 -2369 726 -2369 0 4
rlabel polysilicon 730 -2363 730 -2363 0 1
rlabel polysilicon 730 -2369 730 -2369 0 3
rlabel polysilicon 737 -2363 737 -2363 0 1
rlabel polysilicon 737 -2369 737 -2369 0 3
rlabel polysilicon 744 -2363 744 -2363 0 1
rlabel polysilicon 747 -2363 747 -2363 0 2
rlabel polysilicon 744 -2369 744 -2369 0 3
rlabel polysilicon 751 -2363 751 -2363 0 1
rlabel polysilicon 751 -2369 751 -2369 0 3
rlabel polysilicon 758 -2363 758 -2363 0 1
rlabel polysilicon 761 -2363 761 -2363 0 2
rlabel polysilicon 758 -2369 758 -2369 0 3
rlabel polysilicon 761 -2369 761 -2369 0 4
rlabel polysilicon 765 -2363 765 -2363 0 1
rlabel polysilicon 765 -2369 765 -2369 0 3
rlabel polysilicon 772 -2363 772 -2363 0 1
rlabel polysilicon 772 -2369 772 -2369 0 3
rlabel polysilicon 779 -2363 779 -2363 0 1
rlabel polysilicon 779 -2369 779 -2369 0 3
rlabel polysilicon 786 -2363 786 -2363 0 1
rlabel polysilicon 786 -2369 786 -2369 0 3
rlabel polysilicon 793 -2363 793 -2363 0 1
rlabel polysilicon 793 -2369 793 -2369 0 3
rlabel polysilicon 800 -2363 800 -2363 0 1
rlabel polysilicon 800 -2369 800 -2369 0 3
rlabel polysilicon 807 -2363 807 -2363 0 1
rlabel polysilicon 810 -2363 810 -2363 0 2
rlabel polysilicon 807 -2369 807 -2369 0 3
rlabel polysilicon 810 -2369 810 -2369 0 4
rlabel polysilicon 814 -2363 814 -2363 0 1
rlabel polysilicon 814 -2369 814 -2369 0 3
rlabel polysilicon 821 -2363 821 -2363 0 1
rlabel polysilicon 821 -2369 821 -2369 0 3
rlabel polysilicon 828 -2363 828 -2363 0 1
rlabel polysilicon 828 -2369 828 -2369 0 3
rlabel polysilicon 835 -2363 835 -2363 0 1
rlabel polysilicon 835 -2369 835 -2369 0 3
rlabel polysilicon 842 -2363 842 -2363 0 1
rlabel polysilicon 842 -2369 842 -2369 0 3
rlabel polysilicon 849 -2363 849 -2363 0 1
rlabel polysilicon 849 -2369 849 -2369 0 3
rlabel polysilicon 852 -2369 852 -2369 0 4
rlabel polysilicon 856 -2363 856 -2363 0 1
rlabel polysilicon 856 -2369 856 -2369 0 3
rlabel polysilicon 863 -2363 863 -2363 0 1
rlabel polysilicon 863 -2369 863 -2369 0 3
rlabel polysilicon 870 -2363 870 -2363 0 1
rlabel polysilicon 870 -2369 870 -2369 0 3
rlabel polysilicon 877 -2363 877 -2363 0 1
rlabel polysilicon 877 -2369 877 -2369 0 3
rlabel polysilicon 884 -2363 884 -2363 0 1
rlabel polysilicon 884 -2369 884 -2369 0 3
rlabel polysilicon 891 -2363 891 -2363 0 1
rlabel polysilicon 891 -2369 891 -2369 0 3
rlabel polysilicon 898 -2363 898 -2363 0 1
rlabel polysilicon 898 -2369 898 -2369 0 3
rlabel polysilicon 905 -2363 905 -2363 0 1
rlabel polysilicon 905 -2369 905 -2369 0 3
rlabel polysilicon 912 -2363 912 -2363 0 1
rlabel polysilicon 912 -2369 912 -2369 0 3
rlabel polysilicon 919 -2363 919 -2363 0 1
rlabel polysilicon 919 -2369 919 -2369 0 3
rlabel polysilicon 926 -2363 926 -2363 0 1
rlabel polysilicon 926 -2369 926 -2369 0 3
rlabel polysilicon 933 -2363 933 -2363 0 1
rlabel polysilicon 933 -2369 933 -2369 0 3
rlabel polysilicon 940 -2363 940 -2363 0 1
rlabel polysilicon 940 -2369 940 -2369 0 3
rlabel polysilicon 947 -2363 947 -2363 0 1
rlabel polysilicon 947 -2369 947 -2369 0 3
rlabel polysilicon 954 -2363 954 -2363 0 1
rlabel polysilicon 954 -2369 954 -2369 0 3
rlabel polysilicon 961 -2363 961 -2363 0 1
rlabel polysilicon 961 -2369 961 -2369 0 3
rlabel polysilicon 968 -2363 968 -2363 0 1
rlabel polysilicon 968 -2369 968 -2369 0 3
rlabel polysilicon 975 -2363 975 -2363 0 1
rlabel polysilicon 975 -2369 975 -2369 0 3
rlabel polysilicon 982 -2363 982 -2363 0 1
rlabel polysilicon 982 -2369 982 -2369 0 3
rlabel polysilicon 989 -2363 989 -2363 0 1
rlabel polysilicon 989 -2369 989 -2369 0 3
rlabel polysilicon 996 -2363 996 -2363 0 1
rlabel polysilicon 996 -2369 996 -2369 0 3
rlabel polysilicon 1003 -2363 1003 -2363 0 1
rlabel polysilicon 1003 -2369 1003 -2369 0 3
rlabel polysilicon 1010 -2363 1010 -2363 0 1
rlabel polysilicon 1010 -2369 1010 -2369 0 3
rlabel polysilicon 1017 -2363 1017 -2363 0 1
rlabel polysilicon 1017 -2369 1017 -2369 0 3
rlabel polysilicon 1024 -2363 1024 -2363 0 1
rlabel polysilicon 1024 -2369 1024 -2369 0 3
rlabel polysilicon 1031 -2363 1031 -2363 0 1
rlabel polysilicon 1034 -2363 1034 -2363 0 2
rlabel polysilicon 1034 -2369 1034 -2369 0 4
rlabel polysilicon 1038 -2363 1038 -2363 0 1
rlabel polysilicon 1038 -2369 1038 -2369 0 3
rlabel polysilicon 1045 -2363 1045 -2363 0 1
rlabel polysilicon 1045 -2369 1045 -2369 0 3
rlabel polysilicon 1052 -2363 1052 -2363 0 1
rlabel polysilicon 1052 -2369 1052 -2369 0 3
rlabel polysilicon 1059 -2363 1059 -2363 0 1
rlabel polysilicon 1059 -2369 1059 -2369 0 3
rlabel polysilicon 1066 -2363 1066 -2363 0 1
rlabel polysilicon 1066 -2369 1066 -2369 0 3
rlabel polysilicon 1073 -2363 1073 -2363 0 1
rlabel polysilicon 1073 -2369 1073 -2369 0 3
rlabel polysilicon 1080 -2363 1080 -2363 0 1
rlabel polysilicon 1080 -2369 1080 -2369 0 3
rlabel polysilicon 1087 -2363 1087 -2363 0 1
rlabel polysilicon 1087 -2369 1087 -2369 0 3
rlabel polysilicon 1094 -2363 1094 -2363 0 1
rlabel polysilicon 1094 -2369 1094 -2369 0 3
rlabel polysilicon 1101 -2363 1101 -2363 0 1
rlabel polysilicon 1101 -2369 1101 -2369 0 3
rlabel polysilicon 1108 -2363 1108 -2363 0 1
rlabel polysilicon 1108 -2369 1108 -2369 0 3
rlabel polysilicon 1115 -2363 1115 -2363 0 1
rlabel polysilicon 1115 -2369 1115 -2369 0 3
rlabel polysilicon 1122 -2363 1122 -2363 0 1
rlabel polysilicon 1122 -2369 1122 -2369 0 3
rlabel polysilicon 1129 -2363 1129 -2363 0 1
rlabel polysilicon 1129 -2369 1129 -2369 0 3
rlabel polysilicon 1136 -2363 1136 -2363 0 1
rlabel polysilicon 1136 -2369 1136 -2369 0 3
rlabel polysilicon 1143 -2363 1143 -2363 0 1
rlabel polysilicon 1143 -2369 1143 -2369 0 3
rlabel polysilicon 1150 -2363 1150 -2363 0 1
rlabel polysilicon 1150 -2369 1150 -2369 0 3
rlabel polysilicon 1157 -2363 1157 -2363 0 1
rlabel polysilicon 1157 -2369 1157 -2369 0 3
rlabel polysilicon 1164 -2363 1164 -2363 0 1
rlabel polysilicon 1164 -2369 1164 -2369 0 3
rlabel polysilicon 1171 -2363 1171 -2363 0 1
rlabel polysilicon 1171 -2369 1171 -2369 0 3
rlabel polysilicon 1178 -2363 1178 -2363 0 1
rlabel polysilicon 1178 -2369 1178 -2369 0 3
rlabel polysilicon 1185 -2363 1185 -2363 0 1
rlabel polysilicon 1185 -2369 1185 -2369 0 3
rlabel polysilicon 1192 -2363 1192 -2363 0 1
rlabel polysilicon 1192 -2369 1192 -2369 0 3
rlabel polysilicon 1199 -2363 1199 -2363 0 1
rlabel polysilicon 1199 -2369 1199 -2369 0 3
rlabel polysilicon 1206 -2363 1206 -2363 0 1
rlabel polysilicon 1206 -2369 1206 -2369 0 3
rlabel polysilicon 1213 -2363 1213 -2363 0 1
rlabel polysilicon 1213 -2369 1213 -2369 0 3
rlabel polysilicon 1220 -2363 1220 -2363 0 1
rlabel polysilicon 1220 -2369 1220 -2369 0 3
rlabel polysilicon 1227 -2363 1227 -2363 0 1
rlabel polysilicon 1227 -2369 1227 -2369 0 3
rlabel polysilicon 1234 -2363 1234 -2363 0 1
rlabel polysilicon 1234 -2369 1234 -2369 0 3
rlabel polysilicon 1241 -2363 1241 -2363 0 1
rlabel polysilicon 1241 -2369 1241 -2369 0 3
rlabel polysilicon 1248 -2363 1248 -2363 0 1
rlabel polysilicon 1248 -2369 1248 -2369 0 3
rlabel polysilicon 58 -2460 58 -2460 0 1
rlabel polysilicon 58 -2466 58 -2466 0 3
rlabel polysilicon 65 -2460 65 -2460 0 1
rlabel polysilicon 65 -2466 65 -2466 0 3
rlabel polysilicon 72 -2460 72 -2460 0 1
rlabel polysilicon 72 -2466 72 -2466 0 3
rlabel polysilicon 79 -2460 79 -2460 0 1
rlabel polysilicon 79 -2466 79 -2466 0 3
rlabel polysilicon 86 -2460 86 -2460 0 1
rlabel polysilicon 86 -2466 86 -2466 0 3
rlabel polysilicon 93 -2460 93 -2460 0 1
rlabel polysilicon 93 -2466 93 -2466 0 3
rlabel polysilicon 100 -2460 100 -2460 0 1
rlabel polysilicon 100 -2466 100 -2466 0 3
rlabel polysilicon 107 -2460 107 -2460 0 1
rlabel polysilicon 107 -2466 107 -2466 0 3
rlabel polysilicon 114 -2460 114 -2460 0 1
rlabel polysilicon 114 -2466 114 -2466 0 3
rlabel polysilicon 124 -2460 124 -2460 0 2
rlabel polysilicon 121 -2466 121 -2466 0 3
rlabel polysilicon 124 -2466 124 -2466 0 4
rlabel polysilicon 128 -2460 128 -2460 0 1
rlabel polysilicon 131 -2460 131 -2460 0 2
rlabel polysilicon 128 -2466 128 -2466 0 3
rlabel polysilicon 131 -2466 131 -2466 0 4
rlabel polysilicon 135 -2460 135 -2460 0 1
rlabel polysilicon 135 -2466 135 -2466 0 3
rlabel polysilicon 142 -2460 142 -2460 0 1
rlabel polysilicon 142 -2466 142 -2466 0 3
rlabel polysilicon 149 -2460 149 -2460 0 1
rlabel polysilicon 149 -2466 149 -2466 0 3
rlabel polysilicon 156 -2460 156 -2460 0 1
rlabel polysilicon 156 -2466 156 -2466 0 3
rlabel polysilicon 163 -2460 163 -2460 0 1
rlabel polysilicon 166 -2466 166 -2466 0 4
rlabel polysilicon 170 -2460 170 -2460 0 1
rlabel polysilicon 170 -2466 170 -2466 0 3
rlabel polysilicon 173 -2466 173 -2466 0 4
rlabel polysilicon 177 -2460 177 -2460 0 1
rlabel polysilicon 177 -2466 177 -2466 0 3
rlabel polysilicon 184 -2460 184 -2460 0 1
rlabel polysilicon 184 -2466 184 -2466 0 3
rlabel polysilicon 191 -2460 191 -2460 0 1
rlabel polysilicon 191 -2466 191 -2466 0 3
rlabel polysilicon 198 -2460 198 -2460 0 1
rlabel polysilicon 201 -2460 201 -2460 0 2
rlabel polysilicon 201 -2466 201 -2466 0 4
rlabel polysilicon 205 -2460 205 -2460 0 1
rlabel polysilicon 205 -2466 205 -2466 0 3
rlabel polysilicon 212 -2460 212 -2460 0 1
rlabel polysilicon 212 -2466 212 -2466 0 3
rlabel polysilicon 219 -2460 219 -2460 0 1
rlabel polysilicon 219 -2466 219 -2466 0 3
rlabel polysilicon 226 -2460 226 -2460 0 1
rlabel polysilicon 226 -2466 226 -2466 0 3
rlabel polysilicon 233 -2460 233 -2460 0 1
rlabel polysilicon 233 -2466 233 -2466 0 3
rlabel polysilicon 240 -2460 240 -2460 0 1
rlabel polysilicon 240 -2466 240 -2466 0 3
rlabel polysilicon 247 -2460 247 -2460 0 1
rlabel polysilicon 247 -2466 247 -2466 0 3
rlabel polysilicon 254 -2460 254 -2460 0 1
rlabel polysilicon 254 -2466 254 -2466 0 3
rlabel polysilicon 261 -2460 261 -2460 0 1
rlabel polysilicon 261 -2466 261 -2466 0 3
rlabel polysilicon 268 -2460 268 -2460 0 1
rlabel polysilicon 268 -2466 268 -2466 0 3
rlabel polysilicon 275 -2460 275 -2460 0 1
rlabel polysilicon 275 -2466 275 -2466 0 3
rlabel polysilicon 282 -2460 282 -2460 0 1
rlabel polysilicon 282 -2466 282 -2466 0 3
rlabel polysilicon 289 -2460 289 -2460 0 1
rlabel polysilicon 289 -2466 289 -2466 0 3
rlabel polysilicon 296 -2460 296 -2460 0 1
rlabel polysilicon 296 -2466 296 -2466 0 3
rlabel polysilicon 303 -2460 303 -2460 0 1
rlabel polysilicon 303 -2466 303 -2466 0 3
rlabel polysilicon 310 -2460 310 -2460 0 1
rlabel polysilicon 310 -2466 310 -2466 0 3
rlabel polysilicon 317 -2460 317 -2460 0 1
rlabel polysilicon 317 -2466 317 -2466 0 3
rlabel polysilicon 324 -2460 324 -2460 0 1
rlabel polysilicon 324 -2466 324 -2466 0 3
rlabel polysilicon 331 -2460 331 -2460 0 1
rlabel polysilicon 331 -2466 331 -2466 0 3
rlabel polysilicon 338 -2460 338 -2460 0 1
rlabel polysilicon 338 -2466 338 -2466 0 3
rlabel polysilicon 345 -2460 345 -2460 0 1
rlabel polysilicon 345 -2466 345 -2466 0 3
rlabel polysilicon 352 -2460 352 -2460 0 1
rlabel polysilicon 352 -2466 352 -2466 0 3
rlabel polysilicon 355 -2466 355 -2466 0 4
rlabel polysilicon 359 -2460 359 -2460 0 1
rlabel polysilicon 359 -2466 359 -2466 0 3
rlabel polysilicon 366 -2460 366 -2460 0 1
rlabel polysilicon 366 -2466 366 -2466 0 3
rlabel polysilicon 373 -2460 373 -2460 0 1
rlabel polysilicon 376 -2460 376 -2460 0 2
rlabel polysilicon 373 -2466 373 -2466 0 3
rlabel polysilicon 376 -2466 376 -2466 0 4
rlabel polysilicon 380 -2460 380 -2460 0 1
rlabel polysilicon 380 -2466 380 -2466 0 3
rlabel polysilicon 387 -2460 387 -2460 0 1
rlabel polysilicon 387 -2466 387 -2466 0 3
rlabel polysilicon 394 -2460 394 -2460 0 1
rlabel polysilicon 394 -2466 394 -2466 0 3
rlabel polysilicon 401 -2460 401 -2460 0 1
rlabel polysilicon 401 -2466 401 -2466 0 3
rlabel polysilicon 408 -2460 408 -2460 0 1
rlabel polysilicon 408 -2466 408 -2466 0 3
rlabel polysilicon 415 -2460 415 -2460 0 1
rlabel polysilicon 415 -2466 415 -2466 0 3
rlabel polysilicon 422 -2460 422 -2460 0 1
rlabel polysilicon 422 -2466 422 -2466 0 3
rlabel polysilicon 429 -2460 429 -2460 0 1
rlabel polysilicon 429 -2466 429 -2466 0 3
rlabel polysilicon 439 -2460 439 -2460 0 2
rlabel polysilicon 436 -2466 436 -2466 0 3
rlabel polysilicon 439 -2466 439 -2466 0 4
rlabel polysilicon 443 -2460 443 -2460 0 1
rlabel polysilicon 446 -2460 446 -2460 0 2
rlabel polysilicon 443 -2466 443 -2466 0 3
rlabel polysilicon 446 -2466 446 -2466 0 4
rlabel polysilicon 450 -2460 450 -2460 0 1
rlabel polysilicon 450 -2466 450 -2466 0 3
rlabel polysilicon 457 -2460 457 -2460 0 1
rlabel polysilicon 457 -2466 457 -2466 0 3
rlabel polysilicon 464 -2460 464 -2460 0 1
rlabel polysilicon 467 -2460 467 -2460 0 2
rlabel polysilicon 467 -2466 467 -2466 0 4
rlabel polysilicon 471 -2460 471 -2460 0 1
rlabel polysilicon 471 -2466 471 -2466 0 3
rlabel polysilicon 478 -2460 478 -2460 0 1
rlabel polysilicon 478 -2466 478 -2466 0 3
rlabel polysilicon 485 -2460 485 -2460 0 1
rlabel polysilicon 485 -2466 485 -2466 0 3
rlabel polysilicon 492 -2460 492 -2460 0 1
rlabel polysilicon 492 -2466 492 -2466 0 3
rlabel polysilicon 499 -2460 499 -2460 0 1
rlabel polysilicon 499 -2466 499 -2466 0 3
rlabel polysilicon 506 -2460 506 -2460 0 1
rlabel polysilicon 506 -2466 506 -2466 0 3
rlabel polysilicon 513 -2460 513 -2460 0 1
rlabel polysilicon 516 -2460 516 -2460 0 2
rlabel polysilicon 513 -2466 513 -2466 0 3
rlabel polysilicon 520 -2460 520 -2460 0 1
rlabel polysilicon 520 -2466 520 -2466 0 3
rlabel polysilicon 527 -2460 527 -2460 0 1
rlabel polysilicon 527 -2466 527 -2466 0 3
rlabel polysilicon 534 -2460 534 -2460 0 1
rlabel polysilicon 534 -2466 534 -2466 0 3
rlabel polysilicon 541 -2460 541 -2460 0 1
rlabel polysilicon 541 -2466 541 -2466 0 3
rlabel polysilicon 548 -2460 548 -2460 0 1
rlabel polysilicon 548 -2466 548 -2466 0 3
rlabel polysilicon 555 -2460 555 -2460 0 1
rlabel polysilicon 555 -2466 555 -2466 0 3
rlabel polysilicon 562 -2460 562 -2460 0 1
rlabel polysilicon 562 -2466 562 -2466 0 3
rlabel polysilicon 565 -2466 565 -2466 0 4
rlabel polysilicon 569 -2460 569 -2460 0 1
rlabel polysilicon 572 -2460 572 -2460 0 2
rlabel polysilicon 569 -2466 569 -2466 0 3
rlabel polysilicon 572 -2466 572 -2466 0 4
rlabel polysilicon 576 -2460 576 -2460 0 1
rlabel polysilicon 576 -2466 576 -2466 0 3
rlabel polysilicon 583 -2460 583 -2460 0 1
rlabel polysilicon 583 -2466 583 -2466 0 3
rlabel polysilicon 590 -2460 590 -2460 0 1
rlabel polysilicon 590 -2466 590 -2466 0 3
rlabel polysilicon 597 -2460 597 -2460 0 1
rlabel polysilicon 597 -2466 597 -2466 0 3
rlabel polysilicon 604 -2460 604 -2460 0 1
rlabel polysilicon 604 -2466 604 -2466 0 3
rlabel polysilicon 611 -2460 611 -2460 0 1
rlabel polysilicon 614 -2460 614 -2460 0 2
rlabel polysilicon 611 -2466 611 -2466 0 3
rlabel polysilicon 618 -2460 618 -2460 0 1
rlabel polysilicon 618 -2466 618 -2466 0 3
rlabel polysilicon 625 -2460 625 -2460 0 1
rlabel polysilicon 625 -2466 625 -2466 0 3
rlabel polysilicon 632 -2460 632 -2460 0 1
rlabel polysilicon 632 -2466 632 -2466 0 3
rlabel polysilicon 639 -2460 639 -2460 0 1
rlabel polysilicon 639 -2466 639 -2466 0 3
rlabel polysilicon 646 -2460 646 -2460 0 1
rlabel polysilicon 646 -2466 646 -2466 0 3
rlabel polysilicon 653 -2460 653 -2460 0 1
rlabel polysilicon 653 -2466 653 -2466 0 3
rlabel polysilicon 660 -2460 660 -2460 0 1
rlabel polysilicon 663 -2460 663 -2460 0 2
rlabel polysilicon 660 -2466 660 -2466 0 3
rlabel polysilicon 667 -2460 667 -2460 0 1
rlabel polysilicon 667 -2466 667 -2466 0 3
rlabel polysilicon 674 -2460 674 -2460 0 1
rlabel polysilicon 674 -2466 674 -2466 0 3
rlabel polysilicon 677 -2466 677 -2466 0 4
rlabel polysilicon 681 -2460 681 -2460 0 1
rlabel polysilicon 681 -2466 681 -2466 0 3
rlabel polysilicon 688 -2460 688 -2460 0 1
rlabel polysilicon 688 -2466 688 -2466 0 3
rlabel polysilicon 695 -2460 695 -2460 0 1
rlabel polysilicon 695 -2466 695 -2466 0 3
rlabel polysilicon 702 -2460 702 -2460 0 1
rlabel polysilicon 702 -2466 702 -2466 0 3
rlabel polysilicon 709 -2460 709 -2460 0 1
rlabel polysilicon 709 -2466 709 -2466 0 3
rlabel polysilicon 716 -2460 716 -2460 0 1
rlabel polysilicon 716 -2466 716 -2466 0 3
rlabel polysilicon 723 -2460 723 -2460 0 1
rlabel polysilicon 726 -2460 726 -2460 0 2
rlabel polysilicon 723 -2466 723 -2466 0 3
rlabel polysilicon 730 -2460 730 -2460 0 1
rlabel polysilicon 730 -2466 730 -2466 0 3
rlabel polysilicon 737 -2460 737 -2460 0 1
rlabel polysilicon 737 -2466 737 -2466 0 3
rlabel polysilicon 744 -2460 744 -2460 0 1
rlabel polysilicon 744 -2466 744 -2466 0 3
rlabel polysilicon 751 -2460 751 -2460 0 1
rlabel polysilicon 751 -2466 751 -2466 0 3
rlabel polysilicon 758 -2460 758 -2460 0 1
rlabel polysilicon 758 -2466 758 -2466 0 3
rlabel polysilicon 765 -2460 765 -2460 0 1
rlabel polysilicon 765 -2466 765 -2466 0 3
rlabel polysilicon 772 -2460 772 -2460 0 1
rlabel polysilicon 772 -2466 772 -2466 0 3
rlabel polysilicon 779 -2460 779 -2460 0 1
rlabel polysilicon 779 -2466 779 -2466 0 3
rlabel polysilicon 786 -2460 786 -2460 0 1
rlabel polysilicon 786 -2466 786 -2466 0 3
rlabel polysilicon 796 -2460 796 -2460 0 2
rlabel polysilicon 793 -2466 793 -2466 0 3
rlabel polysilicon 800 -2460 800 -2460 0 1
rlabel polysilicon 800 -2466 800 -2466 0 3
rlabel polysilicon 807 -2460 807 -2460 0 1
rlabel polysilicon 807 -2466 807 -2466 0 3
rlabel polysilicon 814 -2460 814 -2460 0 1
rlabel polysilicon 814 -2466 814 -2466 0 3
rlabel polysilicon 821 -2460 821 -2460 0 1
rlabel polysilicon 821 -2466 821 -2466 0 3
rlabel polysilicon 828 -2460 828 -2460 0 1
rlabel polysilicon 828 -2466 828 -2466 0 3
rlabel polysilicon 835 -2460 835 -2460 0 1
rlabel polysilicon 835 -2466 835 -2466 0 3
rlabel polysilicon 842 -2460 842 -2460 0 1
rlabel polysilicon 842 -2466 842 -2466 0 3
rlabel polysilicon 849 -2460 849 -2460 0 1
rlabel polysilicon 849 -2466 849 -2466 0 3
rlabel polysilicon 856 -2460 856 -2460 0 1
rlabel polysilicon 856 -2466 856 -2466 0 3
rlabel polysilicon 863 -2460 863 -2460 0 1
rlabel polysilicon 863 -2466 863 -2466 0 3
rlabel polysilicon 870 -2460 870 -2460 0 1
rlabel polysilicon 870 -2466 870 -2466 0 3
rlabel polysilicon 877 -2460 877 -2460 0 1
rlabel polysilicon 877 -2466 877 -2466 0 3
rlabel polysilicon 884 -2460 884 -2460 0 1
rlabel polysilicon 884 -2466 884 -2466 0 3
rlabel polysilicon 891 -2460 891 -2460 0 1
rlabel polysilicon 891 -2466 891 -2466 0 3
rlabel polysilicon 898 -2460 898 -2460 0 1
rlabel polysilicon 898 -2466 898 -2466 0 3
rlabel polysilicon 905 -2460 905 -2460 0 1
rlabel polysilicon 908 -2460 908 -2460 0 2
rlabel polysilicon 905 -2466 905 -2466 0 3
rlabel polysilicon 912 -2460 912 -2460 0 1
rlabel polysilicon 912 -2466 912 -2466 0 3
rlabel polysilicon 919 -2460 919 -2460 0 1
rlabel polysilicon 919 -2466 919 -2466 0 3
rlabel polysilicon 926 -2460 926 -2460 0 1
rlabel polysilicon 926 -2466 926 -2466 0 3
rlabel polysilicon 933 -2460 933 -2460 0 1
rlabel polysilicon 933 -2466 933 -2466 0 3
rlabel polysilicon 940 -2460 940 -2460 0 1
rlabel polysilicon 943 -2460 943 -2460 0 2
rlabel polysilicon 943 -2466 943 -2466 0 4
rlabel polysilicon 947 -2460 947 -2460 0 1
rlabel polysilicon 947 -2466 947 -2466 0 3
rlabel polysilicon 954 -2460 954 -2460 0 1
rlabel polysilicon 954 -2466 954 -2466 0 3
rlabel polysilicon 961 -2460 961 -2460 0 1
rlabel polysilicon 961 -2466 961 -2466 0 3
rlabel polysilicon 968 -2460 968 -2460 0 1
rlabel polysilicon 968 -2466 968 -2466 0 3
rlabel polysilicon 975 -2460 975 -2460 0 1
rlabel polysilicon 975 -2466 975 -2466 0 3
rlabel polysilicon 982 -2460 982 -2460 0 1
rlabel polysilicon 982 -2466 982 -2466 0 3
rlabel polysilicon 989 -2460 989 -2460 0 1
rlabel polysilicon 989 -2466 989 -2466 0 3
rlabel polysilicon 996 -2460 996 -2460 0 1
rlabel polysilicon 996 -2466 996 -2466 0 3
rlabel polysilicon 1003 -2460 1003 -2460 0 1
rlabel polysilicon 1003 -2466 1003 -2466 0 3
rlabel polysilicon 1010 -2460 1010 -2460 0 1
rlabel polysilicon 1013 -2460 1013 -2460 0 2
rlabel polysilicon 1013 -2466 1013 -2466 0 4
rlabel polysilicon 1017 -2460 1017 -2460 0 1
rlabel polysilicon 1017 -2466 1017 -2466 0 3
rlabel polysilicon 1024 -2460 1024 -2460 0 1
rlabel polysilicon 1024 -2466 1024 -2466 0 3
rlabel polysilicon 1031 -2460 1031 -2460 0 1
rlabel polysilicon 1031 -2466 1031 -2466 0 3
rlabel polysilicon 1059 -2460 1059 -2460 0 1
rlabel polysilicon 1059 -2466 1059 -2466 0 3
rlabel polysilicon 1066 -2460 1066 -2460 0 1
rlabel polysilicon 1066 -2466 1066 -2466 0 3
rlabel polysilicon 1073 -2460 1073 -2460 0 1
rlabel polysilicon 1073 -2466 1073 -2466 0 3
rlabel polysilicon 1080 -2460 1080 -2460 0 1
rlabel polysilicon 1080 -2466 1080 -2466 0 3
rlabel polysilicon 1087 -2460 1087 -2460 0 1
rlabel polysilicon 1087 -2466 1087 -2466 0 3
rlabel polysilicon 1094 -2460 1094 -2460 0 1
rlabel polysilicon 1094 -2466 1094 -2466 0 3
rlabel polysilicon 1101 -2460 1101 -2460 0 1
rlabel polysilicon 1104 -2460 1104 -2460 0 2
rlabel polysilicon 1101 -2466 1101 -2466 0 3
rlabel polysilicon 1104 -2466 1104 -2466 0 4
rlabel polysilicon 1108 -2460 1108 -2460 0 1
rlabel polysilicon 1108 -2466 1108 -2466 0 3
rlabel polysilicon 1129 -2460 1129 -2460 0 1
rlabel polysilicon 1129 -2466 1129 -2466 0 3
rlabel polysilicon 1192 -2460 1192 -2460 0 1
rlabel polysilicon 1192 -2466 1192 -2466 0 3
rlabel polysilicon 128 -2543 128 -2543 0 1
rlabel polysilicon 128 -2549 128 -2549 0 3
rlabel polysilicon 135 -2543 135 -2543 0 1
rlabel polysilicon 135 -2549 135 -2549 0 3
rlabel polysilicon 226 -2543 226 -2543 0 1
rlabel polysilicon 226 -2549 226 -2549 0 3
rlabel polysilicon 233 -2543 233 -2543 0 1
rlabel polysilicon 233 -2549 233 -2549 0 3
rlabel polysilicon 247 -2543 247 -2543 0 1
rlabel polysilicon 247 -2549 247 -2549 0 3
rlabel polysilicon 254 -2543 254 -2543 0 1
rlabel polysilicon 254 -2549 254 -2549 0 3
rlabel polysilicon 261 -2543 261 -2543 0 1
rlabel polysilicon 261 -2549 261 -2549 0 3
rlabel polysilicon 268 -2543 268 -2543 0 1
rlabel polysilicon 268 -2549 268 -2549 0 3
rlabel polysilicon 278 -2543 278 -2543 0 2
rlabel polysilicon 275 -2549 275 -2549 0 3
rlabel polysilicon 282 -2543 282 -2543 0 1
rlabel polysilicon 282 -2549 282 -2549 0 3
rlabel polysilicon 289 -2543 289 -2543 0 1
rlabel polysilicon 289 -2549 289 -2549 0 3
rlabel polysilicon 296 -2543 296 -2543 0 1
rlabel polysilicon 296 -2549 296 -2549 0 3
rlabel polysilicon 303 -2543 303 -2543 0 1
rlabel polysilicon 303 -2549 303 -2549 0 3
rlabel polysilicon 310 -2543 310 -2543 0 1
rlabel polysilicon 310 -2549 310 -2549 0 3
rlabel polysilicon 317 -2543 317 -2543 0 1
rlabel polysilicon 317 -2549 317 -2549 0 3
rlabel polysilicon 327 -2543 327 -2543 0 2
rlabel polysilicon 324 -2549 324 -2549 0 3
rlabel polysilicon 331 -2543 331 -2543 0 1
rlabel polysilicon 331 -2549 331 -2549 0 3
rlabel polysilicon 338 -2543 338 -2543 0 1
rlabel polysilicon 338 -2549 338 -2549 0 3
rlabel polysilicon 345 -2543 345 -2543 0 1
rlabel polysilicon 345 -2549 345 -2549 0 3
rlabel polysilicon 352 -2543 352 -2543 0 1
rlabel polysilicon 352 -2549 352 -2549 0 3
rlabel polysilicon 359 -2543 359 -2543 0 1
rlabel polysilicon 359 -2549 359 -2549 0 3
rlabel polysilicon 366 -2543 366 -2543 0 1
rlabel polysilicon 366 -2549 366 -2549 0 3
rlabel polysilicon 373 -2543 373 -2543 0 1
rlabel polysilicon 373 -2549 373 -2549 0 3
rlabel polysilicon 380 -2543 380 -2543 0 1
rlabel polysilicon 380 -2549 380 -2549 0 3
rlabel polysilicon 387 -2543 387 -2543 0 1
rlabel polysilicon 390 -2543 390 -2543 0 2
rlabel polysilicon 387 -2549 387 -2549 0 3
rlabel polysilicon 394 -2543 394 -2543 0 1
rlabel polysilicon 394 -2549 394 -2549 0 3
rlabel polysilicon 401 -2543 401 -2543 0 1
rlabel polysilicon 401 -2549 401 -2549 0 3
rlabel polysilicon 408 -2543 408 -2543 0 1
rlabel polysilicon 408 -2549 408 -2549 0 3
rlabel polysilicon 415 -2543 415 -2543 0 1
rlabel polysilicon 415 -2549 415 -2549 0 3
rlabel polysilicon 422 -2543 422 -2543 0 1
rlabel polysilicon 422 -2549 422 -2549 0 3
rlabel polysilicon 429 -2543 429 -2543 0 1
rlabel polysilicon 429 -2549 429 -2549 0 3
rlabel polysilicon 436 -2543 436 -2543 0 1
rlabel polysilicon 436 -2549 436 -2549 0 3
rlabel polysilicon 443 -2543 443 -2543 0 1
rlabel polysilicon 443 -2549 443 -2549 0 3
rlabel polysilicon 450 -2543 450 -2543 0 1
rlabel polysilicon 450 -2549 450 -2549 0 3
rlabel polysilicon 457 -2543 457 -2543 0 1
rlabel polysilicon 460 -2543 460 -2543 0 2
rlabel polysilicon 460 -2549 460 -2549 0 4
rlabel polysilicon 464 -2543 464 -2543 0 1
rlabel polysilicon 464 -2549 464 -2549 0 3
rlabel polysilicon 471 -2543 471 -2543 0 1
rlabel polysilicon 474 -2543 474 -2543 0 2
rlabel polysilicon 478 -2543 478 -2543 0 1
rlabel polysilicon 478 -2549 478 -2549 0 3
rlabel polysilicon 485 -2543 485 -2543 0 1
rlabel polysilicon 485 -2549 485 -2549 0 3
rlabel polysilicon 488 -2549 488 -2549 0 4
rlabel polysilicon 492 -2543 492 -2543 0 1
rlabel polysilicon 492 -2549 492 -2549 0 3
rlabel polysilicon 499 -2543 499 -2543 0 1
rlabel polysilicon 499 -2549 499 -2549 0 3
rlabel polysilicon 506 -2543 506 -2543 0 1
rlabel polysilicon 509 -2543 509 -2543 0 2
rlabel polysilicon 506 -2549 506 -2549 0 3
rlabel polysilicon 513 -2543 513 -2543 0 1
rlabel polysilicon 513 -2549 513 -2549 0 3
rlabel polysilicon 520 -2543 520 -2543 0 1
rlabel polysilicon 523 -2543 523 -2543 0 2
rlabel polysilicon 523 -2549 523 -2549 0 4
rlabel polysilicon 530 -2543 530 -2543 0 2
rlabel polysilicon 527 -2549 527 -2549 0 3
rlabel polysilicon 530 -2549 530 -2549 0 4
rlabel polysilicon 534 -2543 534 -2543 0 1
rlabel polysilicon 534 -2549 534 -2549 0 3
rlabel polysilicon 544 -2543 544 -2543 0 2
rlabel polysilicon 541 -2549 541 -2549 0 3
rlabel polysilicon 548 -2543 548 -2543 0 1
rlabel polysilicon 551 -2543 551 -2543 0 2
rlabel polysilicon 548 -2549 548 -2549 0 3
rlabel polysilicon 555 -2543 555 -2543 0 1
rlabel polysilicon 555 -2549 555 -2549 0 3
rlabel polysilicon 562 -2543 562 -2543 0 1
rlabel polysilicon 562 -2549 562 -2549 0 3
rlabel polysilicon 569 -2543 569 -2543 0 1
rlabel polysilicon 572 -2543 572 -2543 0 2
rlabel polysilicon 569 -2549 569 -2549 0 3
rlabel polysilicon 576 -2543 576 -2543 0 1
rlabel polysilicon 576 -2549 576 -2549 0 3
rlabel polysilicon 583 -2543 583 -2543 0 1
rlabel polysilicon 586 -2543 586 -2543 0 2
rlabel polysilicon 590 -2543 590 -2543 0 1
rlabel polysilicon 590 -2549 590 -2549 0 3
rlabel polysilicon 593 -2549 593 -2549 0 4
rlabel polysilicon 597 -2543 597 -2543 0 1
rlabel polysilicon 597 -2549 597 -2549 0 3
rlabel polysilicon 604 -2543 604 -2543 0 1
rlabel polysilicon 604 -2549 604 -2549 0 3
rlabel polysilicon 611 -2543 611 -2543 0 1
rlabel polysilicon 611 -2549 611 -2549 0 3
rlabel polysilicon 618 -2543 618 -2543 0 1
rlabel polysilicon 621 -2549 621 -2549 0 4
rlabel polysilicon 625 -2543 625 -2543 0 1
rlabel polysilicon 625 -2549 625 -2549 0 3
rlabel polysilicon 632 -2543 632 -2543 0 1
rlabel polysilicon 632 -2549 632 -2549 0 3
rlabel polysilicon 639 -2543 639 -2543 0 1
rlabel polysilicon 639 -2549 639 -2549 0 3
rlabel polysilicon 646 -2543 646 -2543 0 1
rlabel polysilicon 646 -2549 646 -2549 0 3
rlabel polysilicon 653 -2543 653 -2543 0 1
rlabel polysilicon 653 -2549 653 -2549 0 3
rlabel polysilicon 660 -2543 660 -2543 0 1
rlabel polysilicon 660 -2549 660 -2549 0 3
rlabel polysilicon 667 -2543 667 -2543 0 1
rlabel polysilicon 667 -2549 667 -2549 0 3
rlabel polysilicon 674 -2543 674 -2543 0 1
rlabel polysilicon 674 -2549 674 -2549 0 3
rlabel polysilicon 681 -2543 681 -2543 0 1
rlabel polysilicon 684 -2543 684 -2543 0 2
rlabel polysilicon 681 -2549 681 -2549 0 3
rlabel polysilicon 684 -2549 684 -2549 0 4
rlabel polysilicon 691 -2543 691 -2543 0 2
rlabel polysilicon 688 -2549 688 -2549 0 3
rlabel polysilicon 691 -2549 691 -2549 0 4
rlabel polysilicon 695 -2543 695 -2543 0 1
rlabel polysilicon 695 -2549 695 -2549 0 3
rlabel polysilicon 702 -2543 702 -2543 0 1
rlabel polysilicon 702 -2549 702 -2549 0 3
rlabel polysilicon 709 -2543 709 -2543 0 1
rlabel polysilicon 709 -2549 709 -2549 0 3
rlabel polysilicon 716 -2543 716 -2543 0 1
rlabel polysilicon 716 -2549 716 -2549 0 3
rlabel polysilicon 723 -2543 723 -2543 0 1
rlabel polysilicon 723 -2549 723 -2549 0 3
rlabel polysilicon 730 -2543 730 -2543 0 1
rlabel polysilicon 730 -2549 730 -2549 0 3
rlabel polysilicon 737 -2543 737 -2543 0 1
rlabel polysilicon 740 -2543 740 -2543 0 2
rlabel polysilicon 744 -2543 744 -2543 0 1
rlabel polysilicon 744 -2549 744 -2549 0 3
rlabel polysilicon 747 -2549 747 -2549 0 4
rlabel polysilicon 751 -2543 751 -2543 0 1
rlabel polysilicon 751 -2549 751 -2549 0 3
rlabel polysilicon 758 -2543 758 -2543 0 1
rlabel polysilicon 758 -2549 758 -2549 0 3
rlabel polysilicon 765 -2543 765 -2543 0 1
rlabel polysilicon 765 -2549 765 -2549 0 3
rlabel polysilicon 772 -2543 772 -2543 0 1
rlabel polysilicon 772 -2549 772 -2549 0 3
rlabel polysilicon 779 -2543 779 -2543 0 1
rlabel polysilicon 779 -2549 779 -2549 0 3
rlabel polysilicon 786 -2543 786 -2543 0 1
rlabel polysilicon 786 -2549 786 -2549 0 3
rlabel polysilicon 793 -2543 793 -2543 0 1
rlabel polysilicon 793 -2549 793 -2549 0 3
rlabel polysilicon 800 -2543 800 -2543 0 1
rlabel polysilicon 800 -2549 800 -2549 0 3
rlabel polysilicon 807 -2543 807 -2543 0 1
rlabel polysilicon 810 -2543 810 -2543 0 2
rlabel polysilicon 807 -2549 807 -2549 0 3
rlabel polysilicon 828 -2543 828 -2543 0 1
rlabel polysilicon 828 -2549 828 -2549 0 3
rlabel polysilicon 863 -2543 863 -2543 0 1
rlabel polysilicon 866 -2543 866 -2543 0 2
rlabel polysilicon 866 -2549 866 -2549 0 4
rlabel polysilicon 870 -2543 870 -2543 0 1
rlabel polysilicon 870 -2549 870 -2549 0 3
rlabel polysilicon 912 -2543 912 -2543 0 1
rlabel polysilicon 912 -2549 912 -2549 0 3
rlabel polysilicon 926 -2543 926 -2543 0 1
rlabel polysilicon 926 -2549 926 -2549 0 3
rlabel polysilicon 933 -2543 933 -2543 0 1
rlabel polysilicon 933 -2549 933 -2549 0 3
rlabel polysilicon 947 -2543 947 -2543 0 1
rlabel polysilicon 947 -2549 947 -2549 0 3
rlabel polysilicon 954 -2543 954 -2543 0 1
rlabel polysilicon 954 -2549 954 -2549 0 3
rlabel polysilicon 975 -2543 975 -2543 0 1
rlabel polysilicon 975 -2549 975 -2549 0 3
rlabel polysilicon 1017 -2543 1017 -2543 0 1
rlabel polysilicon 1017 -2549 1017 -2549 0 3
rlabel polysilicon 1031 -2543 1031 -2543 0 1
rlabel polysilicon 1031 -2549 1031 -2549 0 3
rlabel polysilicon 1038 -2543 1038 -2543 0 1
rlabel polysilicon 1038 -2549 1038 -2549 0 3
rlabel polysilicon 1052 -2543 1052 -2543 0 1
rlabel polysilicon 1052 -2549 1052 -2549 0 3
rlabel polysilicon 1066 -2543 1066 -2543 0 1
rlabel polysilicon 1066 -2549 1066 -2549 0 3
rlabel polysilicon 1094 -2543 1094 -2543 0 1
rlabel polysilicon 1143 -2543 1143 -2543 0 1
rlabel polysilicon 1143 -2549 1143 -2549 0 3
rlabel polysilicon 1178 -2543 1178 -2543 0 1
rlabel polysilicon 1178 -2549 1178 -2549 0 3
rlabel polysilicon 1181 -2549 1181 -2549 0 4
rlabel polysilicon 1185 -2543 1185 -2543 0 1
rlabel polysilicon 1185 -2549 1185 -2549 0 3
rlabel polysilicon 131 -2588 131 -2588 0 2
rlabel polysilicon 131 -2594 131 -2594 0 4
rlabel polysilicon 135 -2588 135 -2588 0 1
rlabel polysilicon 135 -2594 135 -2594 0 3
rlabel polysilicon 254 -2588 254 -2588 0 1
rlabel polysilicon 257 -2588 257 -2588 0 2
rlabel polysilicon 324 -2588 324 -2588 0 1
rlabel polysilicon 324 -2594 324 -2594 0 3
rlabel polysilicon 331 -2588 331 -2588 0 1
rlabel polysilicon 331 -2594 331 -2594 0 3
rlabel polysilicon 338 -2588 338 -2588 0 1
rlabel polysilicon 338 -2594 338 -2594 0 3
rlabel polysilicon 348 -2594 348 -2594 0 4
rlabel polysilicon 366 -2588 366 -2588 0 1
rlabel polysilicon 366 -2594 366 -2594 0 3
rlabel polysilicon 373 -2588 373 -2588 0 1
rlabel polysilicon 373 -2594 373 -2594 0 3
rlabel polysilicon 383 -2588 383 -2588 0 2
rlabel polysilicon 380 -2594 380 -2594 0 3
rlabel polysilicon 383 -2594 383 -2594 0 4
rlabel polysilicon 443 -2588 443 -2588 0 1
rlabel polysilicon 443 -2594 443 -2594 0 3
rlabel polysilicon 450 -2588 450 -2588 0 1
rlabel polysilicon 450 -2594 450 -2594 0 3
rlabel polysilicon 471 -2588 471 -2588 0 1
rlabel polysilicon 471 -2594 471 -2594 0 3
rlabel polysilicon 492 -2588 492 -2588 0 1
rlabel polysilicon 492 -2594 492 -2594 0 3
rlabel polysilicon 499 -2588 499 -2588 0 1
rlabel polysilicon 499 -2594 499 -2594 0 3
rlabel polysilicon 506 -2588 506 -2588 0 1
rlabel polysilicon 506 -2594 506 -2594 0 3
rlabel polysilicon 513 -2588 513 -2588 0 1
rlabel polysilicon 513 -2594 513 -2594 0 3
rlabel polysilicon 516 -2594 516 -2594 0 4
rlabel polysilicon 527 -2588 527 -2588 0 1
rlabel polysilicon 530 -2588 530 -2588 0 2
rlabel polysilicon 534 -2588 534 -2588 0 1
rlabel polysilicon 534 -2594 534 -2594 0 3
rlabel polysilicon 541 -2588 541 -2588 0 1
rlabel polysilicon 544 -2588 544 -2588 0 2
rlabel polysilicon 544 -2594 544 -2594 0 4
rlabel polysilicon 551 -2588 551 -2588 0 2
rlabel polysilicon 548 -2594 548 -2594 0 3
rlabel polysilicon 551 -2594 551 -2594 0 4
rlabel polysilicon 555 -2588 555 -2588 0 1
rlabel polysilicon 555 -2594 555 -2594 0 3
rlabel polysilicon 562 -2588 562 -2588 0 1
rlabel polysilicon 565 -2588 565 -2588 0 2
rlabel polysilicon 565 -2594 565 -2594 0 4
rlabel polysilicon 569 -2588 569 -2588 0 1
rlabel polysilicon 569 -2594 569 -2594 0 3
rlabel polysilicon 576 -2588 576 -2588 0 1
rlabel polysilicon 576 -2594 576 -2594 0 3
rlabel polysilicon 597 -2588 597 -2588 0 1
rlabel polysilicon 600 -2588 600 -2588 0 2
rlabel polysilicon 600 -2594 600 -2594 0 4
rlabel polysilicon 646 -2588 646 -2588 0 1
rlabel polysilicon 649 -2588 649 -2588 0 2
rlabel polysilicon 649 -2594 649 -2594 0 4
rlabel polysilicon 663 -2588 663 -2588 0 2
rlabel polysilicon 660 -2594 660 -2594 0 3
rlabel polysilicon 663 -2594 663 -2594 0 4
rlabel polysilicon 667 -2588 667 -2588 0 1
rlabel polysilicon 667 -2594 667 -2594 0 3
rlabel polysilicon 677 -2588 677 -2588 0 2
rlabel polysilicon 674 -2594 674 -2594 0 3
rlabel polysilicon 681 -2588 681 -2588 0 1
rlabel polysilicon 681 -2594 681 -2594 0 3
rlabel polysilicon 684 -2594 684 -2594 0 4
rlabel polysilicon 691 -2588 691 -2588 0 2
rlabel polysilicon 709 -2588 709 -2588 0 1
rlabel polysilicon 712 -2588 712 -2588 0 2
rlabel polysilicon 709 -2594 709 -2594 0 3
rlabel polysilicon 716 -2588 716 -2588 0 1
rlabel polysilicon 716 -2594 716 -2594 0 3
rlabel polysilicon 723 -2588 723 -2588 0 1
rlabel polysilicon 723 -2594 723 -2594 0 3
rlabel polysilicon 730 -2588 730 -2588 0 1
rlabel polysilicon 730 -2594 730 -2594 0 3
rlabel polysilicon 751 -2588 751 -2588 0 1
rlabel polysilicon 751 -2594 751 -2594 0 3
rlabel polysilicon 810 -2588 810 -2588 0 2
rlabel polysilicon 807 -2594 807 -2594 0 3
rlabel polysilicon 810 -2594 810 -2594 0 4
rlabel polysilicon 814 -2588 814 -2588 0 1
rlabel polysilicon 814 -2594 814 -2594 0 3
rlabel polysilicon 884 -2588 884 -2588 0 1
rlabel polysilicon 887 -2588 887 -2588 0 2
rlabel polysilicon 884 -2594 884 -2594 0 3
rlabel polysilicon 898 -2588 898 -2588 0 1
rlabel polysilicon 898 -2594 898 -2594 0 3
rlabel polysilicon 954 -2588 954 -2588 0 1
rlabel polysilicon 954 -2594 954 -2594 0 3
rlabel polysilicon 964 -2588 964 -2588 0 2
rlabel polysilicon 961 -2594 961 -2594 0 3
rlabel polysilicon 964 -2594 964 -2594 0 4
rlabel polysilicon 968 -2588 968 -2588 0 1
rlabel polysilicon 968 -2594 968 -2594 0 3
rlabel polysilicon 1013 -2588 1013 -2588 0 2
rlabel polysilicon 1010 -2594 1010 -2594 0 3
rlabel polysilicon 1013 -2594 1013 -2594 0 4
rlabel polysilicon 1017 -2588 1017 -2588 0 1
rlabel polysilicon 1017 -2594 1017 -2594 0 3
rlabel polysilicon 1024 -2588 1024 -2588 0 1
rlabel polysilicon 1024 -2594 1024 -2594 0 3
rlabel polysilicon 1045 -2588 1045 -2588 0 1
rlabel polysilicon 1045 -2594 1045 -2594 0 3
rlabel polysilicon 1052 -2594 1052 -2594 0 3
rlabel polysilicon 1055 -2594 1055 -2594 0 4
rlabel polysilicon 1059 -2588 1059 -2588 0 1
rlabel polysilicon 1059 -2594 1059 -2594 0 3
rlabel metal2 215 1 215 1 0 net=1305
rlabel metal2 247 1 247 1 0 net=2815
rlabel metal2 562 1 562 1 0 net=8063
rlabel metal2 667 1 667 1 0 net=5721
rlabel metal2 800 1 800 1 0 net=8275
rlabel metal2 261 -1 261 -1 0 net=3607
rlabel metal2 275 -1 275 -1 0 net=4657
rlabel metal2 411 -1 411 -1 0 net=4351
rlabel metal2 576 -1 576 -1 0 net=4661
rlabel metal2 681 -1 681 -1 0 net=5079
rlabel metal2 338 -3 338 -3 0 net=7915
rlabel metal2 387 -3 387 -3 0 net=2123
rlabel metal2 586 -3 586 -3 0 net=4003
rlabel metal2 373 -5 373 -5 0 net=2915
rlabel metal2 415 -5 415 -5 0 net=4809
rlabel metal2 464 -5 464 -5 0 net=7263
rlabel metal2 604 -5 604 -5 0 net=7851
rlabel metal2 397 -7 397 -7 0 net=6643
rlabel metal2 425 -9 425 -9 0 net=3833
rlabel metal2 429 -11 429 -11 0 net=3669
rlabel metal2 467 -13 467 -13 0 net=6621
rlabel metal2 156 -24 156 -24 0 net=204
rlabel metal2 156 -24 156 -24 0 net=204
rlabel metal2 163 -24 163 -24 0 net=5017
rlabel metal2 292 -24 292 -24 0 net=7916
rlabel metal2 359 -24 359 -24 0 net=5097
rlabel metal2 478 -24 478 -24 0 net=7993
rlabel metal2 621 -24 621 -24 0 net=7071
rlabel metal2 800 -24 800 -24 0 net=1029
rlabel metal2 191 -26 191 -26 0 net=2817
rlabel metal2 254 -26 254 -26 0 net=2953
rlabel metal2 404 -26 404 -26 0 net=5025
rlabel metal2 464 -26 464 -26 0 net=4201
rlabel metal2 639 -26 639 -26 0 net=8065
rlabel metal2 702 -26 702 -26 0 net=5895
rlabel metal2 828 -26 828 -26 0 net=8277
rlabel metal2 215 -28 215 -28 0 net=4319
rlabel metal2 226 -28 226 -28 0 net=4659
rlabel metal2 282 -28 282 -28 0 net=4763
rlabel metal2 401 -28 401 -28 0 net=2211
rlabel metal2 436 -28 436 -28 0 net=3797
rlabel metal2 481 -28 481 -28 0 net=5655
rlabel metal2 667 -28 667 -28 0 net=5723
rlabel metal2 709 -28 709 -28 0 net=4005
rlabel metal2 765 -28 765 -28 0 net=7853
rlabel metal2 233 -30 233 -30 0 net=1307
rlabel metal2 247 -30 247 -30 0 net=3609
rlabel metal2 268 -30 268 -30 0 net=3775
rlabel metal2 408 -30 408 -30 0 net=4543
rlabel metal2 485 -30 485 -30 0 net=6645
rlabel metal2 527 -30 527 -30 0 net=7265
rlabel metal2 551 -30 551 -30 0 net=4589
rlabel metal2 639 -30 639 -30 0 net=5081
rlabel metal2 719 -30 719 -30 0 net=6627
rlabel metal2 261 -32 261 -32 0 net=2125
rlabel metal2 492 -32 492 -32 0 net=5595
rlabel metal2 555 -32 555 -32 0 net=5927
rlabel metal2 275 -34 275 -34 0 net=1447
rlabel metal2 366 -34 366 -34 0 net=1483
rlabel metal2 516 -34 516 -34 0 net=5771
rlabel metal2 653 -34 653 -34 0 net=4449
rlabel metal2 282 -36 282 -36 0 net=2263
rlabel metal2 499 -36 499 -36 0 net=6623
rlabel metal2 534 -36 534 -36 0 net=8231
rlabel metal2 296 -38 296 -38 0 net=3671
rlabel metal2 502 -38 502 -38 0 net=1911
rlabel metal2 548 -38 548 -38 0 net=7459
rlabel metal2 303 -40 303 -40 0 net=3233
rlabel metal2 429 -40 429 -40 0 net=7847
rlabel metal2 569 -40 569 -40 0 net=3835
rlabel metal2 310 -42 310 -42 0 net=6005
rlabel metal2 457 -42 457 -42 0 net=6935
rlabel metal2 576 -42 576 -42 0 net=4663
rlabel metal2 317 -44 317 -44 0 net=3339
rlabel metal2 583 -44 583 -44 0 net=2129
rlabel metal2 324 -46 324 -46 0 net=2917
rlabel metal2 380 -46 380 -46 0 net=6109
rlabel metal2 506 -46 506 -46 0 net=4353
rlabel metal2 593 -46 593 -46 0 net=6807
rlabel metal2 331 -48 331 -48 0 net=2301
rlabel metal2 457 -48 457 -48 0 net=3997
rlabel metal2 506 -48 506 -48 0 net=6797
rlabel metal2 345 -50 345 -50 0 net=238
rlabel metal2 373 -52 373 -52 0 net=4811
rlabel metal2 380 -54 380 -54 0 net=8185
rlabel metal2 387 -56 387 -56 0 net=3405
rlabel metal2 23 -67 23 -67 0 net=3955
rlabel metal2 415 -67 415 -67 0 net=7460
rlabel metal2 562 -67 562 -67 0 net=8187
rlabel metal2 723 -67 723 -67 0 net=7073
rlabel metal2 828 -67 828 -67 0 net=7855
rlabel metal2 877 -67 877 -67 0 net=6629
rlabel metal2 1500 -67 1500 -67 0 net=6315
rlabel metal2 30 -69 30 -69 0 net=2845
rlabel metal2 156 -69 156 -69 0 net=1145
rlabel metal2 303 -69 303 -69 0 net=3235
rlabel metal2 303 -69 303 -69 0 net=3235
rlabel metal2 313 -69 313 -69 0 net=778
rlabel metal2 422 -69 422 -69 0 net=6007
rlabel metal2 562 -69 562 -69 0 net=5083
rlabel metal2 663 -69 663 -69 0 net=7677
rlabel metal2 905 -69 905 -69 0 net=1031
rlabel metal2 37 -71 37 -71 0 net=2303
rlabel metal2 373 -71 373 -71 0 net=4813
rlabel metal2 478 -71 478 -71 0 net=5439
rlabel metal2 702 -71 702 -71 0 net=8233
rlabel metal2 849 -71 849 -71 0 net=8279
rlabel metal2 44 -73 44 -73 0 net=5959
rlabel metal2 170 -73 170 -73 0 net=3735
rlabel metal2 324 -73 324 -73 0 net=2919
rlabel metal2 394 -73 394 -73 0 net=4765
rlabel metal2 481 -73 481 -73 0 net=6110
rlabel metal2 499 -73 499 -73 0 net=4773
rlabel metal2 541 -73 541 -73 0 net=7266
rlabel metal2 604 -73 604 -73 0 net=7995
rlabel metal2 751 -73 751 -73 0 net=5897
rlabel metal2 51 -75 51 -75 0 net=1485
rlabel metal2 373 -75 373 -75 0 net=7849
rlabel metal2 471 -75 471 -75 0 net=4545
rlabel metal2 576 -75 576 -75 0 net=8017
rlabel metal2 75 -77 75 -77 0 net=3297
rlabel metal2 107 -77 107 -77 0 net=1581
rlabel metal2 121 -77 121 -77 0 net=1731
rlabel metal2 471 -77 471 -77 0 net=3083
rlabel metal2 576 -77 576 -77 0 net=4847
rlabel metal2 604 -77 604 -77 0 net=8091
rlabel metal2 758 -77 758 -77 0 net=4007
rlabel metal2 79 -79 79 -79 0 net=2269
rlabel metal2 429 -79 429 -79 0 net=3999
rlabel metal2 485 -79 485 -79 0 net=4665
rlabel metal2 618 -79 618 -79 0 net=7839
rlabel metal2 772 -79 772 -79 0 net=6809
rlabel metal2 86 -81 86 -81 0 net=544
rlabel metal2 93 -81 93 -81 0 net=1449
rlabel metal2 296 -81 296 -81 0 net=3673
rlabel metal2 436 -81 436 -81 0 net=3799
rlabel metal2 499 -81 499 -81 0 net=3259
rlabel metal2 618 -81 618 -81 0 net=5725
rlabel metal2 681 -81 681 -81 0 net=5929
rlabel metal2 114 -83 114 -83 0 net=2539
rlabel metal2 299 -83 299 -83 0 net=622
rlabel metal2 450 -83 450 -83 0 net=4591
rlabel metal2 632 -83 632 -83 0 net=5773
rlabel metal2 688 -83 688 -83 0 net=8067
rlabel metal2 128 -85 128 -85 0 net=1271
rlabel metal2 219 -85 219 -85 0 net=4321
rlabel metal2 352 -85 352 -85 0 net=4297
rlabel metal2 625 -85 625 -85 0 net=3837
rlabel metal2 646 -85 646 -85 0 net=2131
rlabel metal2 135 -87 135 -87 0 net=3341
rlabel metal2 352 -87 352 -87 0 net=5099
rlabel metal2 366 -87 366 -87 0 net=3407
rlabel metal2 404 -87 404 -87 0 net=6803
rlabel metal2 660 -87 660 -87 0 net=5657
rlabel metal2 142 -89 142 -89 0 net=5019
rlabel metal2 177 -89 177 -89 0 net=2443
rlabel metal2 359 -89 359 -89 0 net=7453
rlabel metal2 163 -91 163 -91 0 net=1903
rlabel metal2 338 -91 338 -91 0 net=3253
rlabel metal2 453 -91 453 -91 0 net=7231
rlabel metal2 184 -93 184 -93 0 net=2264
rlabel metal2 338 -93 338 -93 0 net=2577
rlabel metal2 506 -93 506 -93 0 net=6799
rlabel metal2 625 -93 625 -93 0 net=4451
rlabel metal2 660 -93 660 -93 0 net=8055
rlabel metal2 187 -95 187 -95 0 net=4660
rlabel metal2 254 -95 254 -95 0 net=2955
rlabel metal2 464 -95 464 -95 0 net=4203
rlabel metal2 513 -95 513 -95 0 net=6625
rlabel metal2 667 -95 667 -95 0 net=6245
rlabel metal2 149 -97 149 -97 0 net=5451
rlabel metal2 254 -97 254 -97 0 net=2127
rlabel metal2 268 -97 268 -97 0 net=3777
rlabel metal2 411 -97 411 -97 0 net=4367
rlabel metal2 520 -97 520 -97 0 net=6647
rlabel metal2 670 -97 670 -97 0 net=7199
rlabel metal2 149 -99 149 -99 0 net=3151
rlabel metal2 198 -99 198 -99 0 net=1309
rlabel metal2 247 -99 247 -99 0 net=3610
rlabel metal2 271 -99 271 -99 0 net=358
rlabel metal2 520 -99 520 -99 0 net=4175
rlabel metal2 191 -101 191 -101 0 net=2819
rlabel metal2 247 -101 247 -101 0 net=1679
rlabel metal2 527 -101 527 -101 0 net=1913
rlabel metal2 205 -103 205 -103 0 net=1321
rlabel metal2 530 -103 530 -103 0 net=5253
rlabel metal2 219 -105 219 -105 0 net=1589
rlabel metal2 569 -105 569 -105 0 net=6937
rlabel metal2 233 -107 233 -107 0 net=2551
rlabel metal2 345 -107 345 -107 0 net=2681
rlabel metal2 65 -109 65 -109 0 net=2209
rlabel metal2 443 -109 443 -109 0 net=5027
rlabel metal2 261 -111 261 -111 0 net=2213
rlabel metal2 439 -111 439 -111 0 net=3429
rlabel metal2 492 -111 492 -111 0 net=5597
rlabel metal2 282 -113 282 -113 0 net=1555
rlabel metal2 401 -115 401 -115 0 net=6089
rlabel metal2 492 -115 492 -115 0 net=4355
rlabel metal2 583 -117 583 -117 0 net=4929
rlabel metal2 16 -128 16 -128 0 net=4133
rlabel metal2 488 -128 488 -128 0 net=1914
rlabel metal2 793 -128 793 -128 0 net=5255
rlabel metal2 849 -128 849 -128 0 net=6811
rlabel metal2 940 -128 940 -128 0 net=6631
rlabel metal2 975 -128 975 -128 0 net=7625
rlabel metal2 1500 -128 1500 -128 0 net=6317
rlabel metal2 1500 -128 1500 -128 0 net=6317
rlabel metal2 9 -130 9 -130 0 net=2371
rlabel metal2 516 -130 516 -130 0 net=6626
rlabel metal2 604 -130 604 -130 0 net=2132
rlabel metal2 800 -130 800 -130 0 net=8235
rlabel metal2 947 -130 947 -130 0 net=1032
rlabel metal2 23 -132 23 -132 0 net=3957
rlabel metal2 23 -132 23 -132 0 net=3957
rlabel metal2 30 -132 30 -132 0 net=2846
rlabel metal2 58 -132 58 -132 0 net=3473
rlabel metal2 72 -132 72 -132 0 net=3691
rlabel metal2 86 -132 86 -132 0 net=3409
rlabel metal2 394 -132 394 -132 0 net=3067
rlabel metal2 30 -134 30 -134 0 net=1195
rlabel metal2 107 -134 107 -134 0 net=1583
rlabel metal2 117 -134 117 -134 0 net=926
rlabel metal2 537 -134 537 -134 0 net=7937
rlabel metal2 849 -134 849 -134 0 net=7411
rlabel metal2 44 -136 44 -136 0 net=5960
rlabel metal2 275 -136 275 -136 0 net=2541
rlabel metal2 541 -136 541 -136 0 net=4547
rlabel metal2 607 -136 607 -136 0 net=8315
rlabel metal2 51 -138 51 -138 0 net=1486
rlabel metal2 464 -138 464 -138 0 net=6090
rlabel metal2 611 -138 611 -138 0 net=6801
rlabel metal2 856 -138 856 -138 0 net=7679
rlabel metal2 51 -140 51 -140 0 net=5020
rlabel metal2 145 -140 145 -140 0 net=678
rlabel metal2 310 -140 310 -140 0 net=4283
rlabel metal2 443 -140 443 -140 0 net=3431
rlabel metal2 478 -140 478 -140 0 net=4767
rlabel metal2 632 -140 632 -140 0 net=3839
rlabel metal2 632 -140 632 -140 0 net=3839
rlabel metal2 646 -140 646 -140 0 net=6805
rlabel metal2 807 -140 807 -140 0 net=7201
rlabel metal2 58 -142 58 -142 0 net=2271
rlabel metal2 93 -142 93 -142 0 net=1451
rlabel metal2 289 -142 289 -142 0 net=2210
rlabel metal2 555 -142 555 -142 0 net=4299
rlabel metal2 79 -144 79 -144 0 net=1905
rlabel metal2 226 -144 226 -144 0 net=5452
rlabel metal2 327 -144 327 -144 0 net=5100
rlabel metal2 422 -144 422 -144 0 net=3675
rlabel metal2 513 -144 513 -144 0 net=4369
rlabel metal2 562 -144 562 -144 0 net=5085
rlabel metal2 779 -144 779 -144 0 net=7075
rlabel metal2 870 -144 870 -144 0 net=7857
rlabel metal2 121 -146 121 -146 0 net=1733
rlabel metal2 226 -146 226 -146 0 net=1495
rlabel metal2 422 -146 422 -146 0 net=3261
rlabel metal2 520 -146 520 -146 0 net=4177
rlabel metal2 646 -146 646 -146 0 net=5775
rlabel metal2 688 -146 688 -146 0 net=7233
rlabel metal2 779 -146 779 -146 0 net=5899
rlabel metal2 821 -146 821 -146 0 net=8019
rlabel metal2 89 -148 89 -148 0 net=4629
rlabel metal2 639 -148 639 -148 0 net=6649
rlabel metal2 877 -148 877 -148 0 net=8281
rlabel metal2 100 -150 100 -150 0 net=3299
rlabel metal2 131 -150 131 -150 0 net=2841
rlabel metal2 324 -150 324 -150 0 net=4877
rlabel metal2 429 -150 429 -150 0 net=4001
rlabel metal2 583 -150 583 -150 0 net=4931
rlabel metal2 653 -150 653 -150 0 net=6939
rlabel metal2 68 -152 68 -152 0 net=953
rlabel metal2 135 -152 135 -152 0 net=3343
rlabel metal2 443 -152 443 -152 0 net=8188
rlabel metal2 716 -152 716 -152 0 net=7841
rlabel metal2 135 -154 135 -154 0 net=3737
rlabel metal2 233 -154 233 -154 0 net=2553
rlabel metal2 485 -154 485 -154 0 net=4667
rlabel metal2 590 -154 590 -154 0 net=5599
rlabel metal2 719 -154 719 -154 0 net=6697
rlabel metal2 807 -154 807 -154 0 net=4515
rlabel metal2 142 -156 142 -156 0 net=226
rlabel metal2 194 -156 194 -156 0 net=1847
rlabel metal2 247 -156 247 -156 0 net=1681
rlabel metal2 415 -156 415 -156 0 net=4815
rlabel metal2 625 -156 625 -156 0 net=4453
rlabel metal2 660 -156 660 -156 0 net=4009
rlabel metal2 149 -158 149 -158 0 net=3152
rlabel metal2 247 -158 247 -158 0 net=2133
rlabel metal2 415 -158 415 -158 0 net=3085
rlabel metal2 485 -158 485 -158 0 net=4225
rlabel metal2 576 -158 576 -158 0 net=4849
rlabel metal2 667 -158 667 -158 0 net=6247
rlabel metal2 44 -160 44 -160 0 net=1201
rlabel metal2 152 -160 152 -160 0 net=1693
rlabel metal2 254 -160 254 -160 0 net=2128
rlabel metal2 387 -160 387 -160 0 net=3255
rlabel metal2 492 -160 492 -160 0 net=4357
rlabel metal2 663 -160 663 -160 0 net=5073
rlabel metal2 674 -160 674 -160 0 net=5659
rlabel metal2 163 -162 163 -162 0 net=2445
rlabel metal2 219 -162 219 -162 0 net=1591
rlabel metal2 271 -162 271 -162 0 net=2956
rlabel metal2 373 -162 373 -162 0 net=7850
rlabel metal2 457 -162 457 -162 0 net=3801
rlabel metal2 569 -162 569 -162 0 net=5029
rlabel metal2 688 -162 688 -162 0 net=5441
rlabel metal2 702 -162 702 -162 0 net=7455
rlabel metal2 170 -164 170 -164 0 net=1323
rlabel metal2 219 -164 219 -164 0 net=3523
rlabel metal2 317 -164 317 -164 0 net=5605
rlabel metal2 723 -164 723 -164 0 net=7997
rlabel metal2 177 -166 177 -166 0 net=1273
rlabel metal2 268 -166 268 -166 0 net=6123
rlabel metal2 730 -166 730 -166 0 net=5931
rlabel metal2 107 -168 107 -168 0 net=1943
rlabel metal2 282 -168 282 -168 0 net=1557
rlabel metal2 303 -168 303 -168 0 net=3237
rlabel metal2 457 -168 457 -168 0 net=5101
rlabel metal2 737 -168 737 -168 0 net=8057
rlabel metal2 198 -170 198 -170 0 net=1311
rlabel metal2 240 -170 240 -170 0 net=2821
rlabel metal2 303 -170 303 -170 0 net=2927
rlabel metal2 530 -170 530 -170 0 net=6101
rlabel metal2 744 -170 744 -170 0 net=8069
rlabel metal2 128 -172 128 -172 0 net=1645
rlabel metal2 331 -172 331 -172 0 net=4323
rlabel metal2 618 -172 618 -172 0 net=5727
rlabel metal2 751 -172 751 -172 0 net=8093
rlabel metal2 93 -174 93 -174 0 net=1963
rlabel metal2 334 -174 334 -174 0 net=5921
rlabel metal2 156 -176 156 -176 0 net=1147
rlabel metal2 436 -176 436 -176 0 net=6209
rlabel metal2 156 -178 156 -178 0 net=2203
rlabel metal2 436 -178 436 -178 0 net=3559
rlabel metal2 534 -178 534 -178 0 net=4775
rlabel metal2 450 -180 450 -180 0 net=4592
rlabel metal2 548 -180 548 -180 0 net=6009
rlabel metal2 408 -182 408 -182 0 net=3779
rlabel metal2 506 -182 506 -182 0 net=4205
rlabel metal2 103 -184 103 -184 0 net=4137
rlabel metal2 380 -186 380 -186 0 net=2921
rlabel metal2 338 -188 338 -188 0 net=2579
rlabel metal2 338 -190 338 -190 0 net=2683
rlabel metal2 37 -192 37 -192 0 net=2305
rlabel metal2 37 -194 37 -194 0 net=2215
rlabel metal2 261 -196 261 -196 0 net=1653
rlabel metal2 2 -207 2 -207 0 net=1197
rlabel metal2 37 -207 37 -207 0 net=2216
rlabel metal2 436 -207 436 -207 0 net=4816
rlabel metal2 604 -207 604 -207 0 net=6989
rlabel metal2 1150 -207 1150 -207 0 net=3745
rlabel metal2 1500 -207 1500 -207 0 net=6319
rlabel metal2 1500 -207 1500 -207 0 net=6319
rlabel metal2 16 -209 16 -209 0 net=4135
rlabel metal2 16 -209 16 -209 0 net=4135
rlabel metal2 37 -209 37 -209 0 net=7499
rlabel metal2 394 -209 394 -209 0 net=3069
rlabel metal2 439 -209 439 -209 0 net=6802
rlabel metal2 849 -209 849 -209 0 net=7413
rlabel metal2 44 -211 44 -211 0 net=1202
rlabel metal2 303 -211 303 -211 0 net=236
rlabel metal2 446 -211 446 -211 0 net=6806
rlabel metal2 835 -211 835 -211 0 net=7939
rlabel metal2 44 -213 44 -213 0 net=3475
rlabel metal2 72 -213 72 -213 0 net=3692
rlabel metal2 103 -213 103 -213 0 net=202
rlabel metal2 243 -213 243 -213 0 net=173
rlabel metal2 544 -213 544 -213 0 net=6650
rlabel metal2 863 -213 863 -213 0 net=8071
rlabel metal2 51 -215 51 -215 0 net=6233
rlabel metal2 1024 -215 1024 -215 0 net=7627
rlabel metal2 51 -217 51 -217 0 net=2219
rlabel metal2 107 -217 107 -217 0 net=1945
rlabel metal2 310 -217 310 -217 0 net=2843
rlabel metal2 453 -217 453 -217 0 net=6940
rlabel metal2 891 -217 891 -217 0 net=7203
rlabel metal2 65 -219 65 -219 0 net=1277
rlabel metal2 107 -219 107 -219 0 net=1543
rlabel metal2 464 -219 464 -219 0 net=3433
rlabel metal2 464 -219 464 -219 0 net=3433
rlabel metal2 471 -219 471 -219 0 net=3257
rlabel metal2 471 -219 471 -219 0 net=3257
rlabel metal2 485 -219 485 -219 0 net=6248
rlabel metal2 821 -219 821 -219 0 net=5257
rlabel metal2 870 -219 870 -219 0 net=8059
rlabel metal2 96 -221 96 -221 0 net=5809
rlabel metal2 912 -221 912 -221 0 net=8237
rlabel metal2 205 -223 205 -223 0 net=1312
rlabel metal2 282 -223 282 -223 0 net=2823
rlabel metal2 159 -225 159 -225 0 net=822
rlabel metal2 310 -225 310 -225 0 net=3133
rlabel metal2 362 -225 362 -225 0 net=5315
rlabel metal2 926 -225 926 -225 0 net=7859
rlabel metal2 198 -227 198 -227 0 net=1149
rlabel metal2 233 -227 233 -227 0 net=1848
rlabel metal2 415 -227 415 -227 0 net=3087
rlabel metal2 457 -227 457 -227 0 net=6043
rlabel metal2 947 -227 947 -227 0 net=8283
rlabel metal2 177 -229 177 -229 0 net=1275
rlabel metal2 233 -229 233 -229 0 net=3267
rlabel metal2 408 -229 408 -229 0 net=2923
rlabel metal2 425 -229 425 -229 0 net=5285
rlabel metal2 947 -229 947 -229 0 net=6307
rlabel metal2 54 -231 54 -231 0 net=6833
rlabel metal2 177 -233 177 -233 0 net=2869
rlabel metal2 320 -233 320 -233 0 net=8353
rlabel metal2 240 -235 240 -235 0 net=2111
rlabel metal2 429 -235 429 -235 0 net=2929
rlabel metal2 506 -235 506 -235 0 net=4139
rlabel metal2 607 -235 607 -235 0 net=7917
rlabel metal2 124 -237 124 -237 0 net=3903
rlabel metal2 513 -237 513 -237 0 net=8201
rlabel metal2 261 -239 261 -239 0 net=1655
rlabel metal2 261 -239 261 -239 0 net=1655
rlabel metal2 268 -239 268 -239 0 net=4002
rlabel metal2 579 -239 579 -239 0 net=8263
rlabel metal2 128 -241 128 -241 0 net=1647
rlabel metal2 373 -241 373 -241 0 net=3239
rlabel metal2 513 -241 513 -241 0 net=4207
rlabel metal2 607 -241 607 -241 0 net=8094
rlabel metal2 954 -241 954 -241 0 net=8021
rlabel metal2 26 -243 26 -243 0 net=6473
rlabel metal2 961 -243 961 -243 0 net=7681
rlabel metal2 128 -245 128 -245 0 net=2205
rlabel metal2 219 -245 219 -245 0 net=3525
rlabel metal2 408 -245 408 -245 0 net=4141
rlabel metal2 632 -245 632 -245 0 net=3841
rlabel metal2 632 -245 632 -245 0 net=3841
rlabel metal2 639 -245 639 -245 0 net=4933
rlabel metal2 919 -245 919 -245 0 net=8317
rlabel metal2 968 -245 968 -245 0 net=6632
rlabel metal2 170 -247 170 -247 0 net=1325
rlabel metal2 219 -247 219 -247 0 net=1497
rlabel metal2 401 -247 401 -247 0 net=4285
rlabel metal2 674 -247 674 -247 0 net=5031
rlabel metal2 800 -247 800 -247 0 net=6699
rlabel metal2 978 -247 978 -247 0 net=6991
rlabel metal2 40 -249 40 -249 0 net=4375
rlabel metal2 345 -249 345 -249 0 net=2307
rlabel metal2 492 -249 492 -249 0 net=3803
rlabel metal2 576 -249 576 -249 0 net=4359
rlabel metal2 688 -249 688 -249 0 net=5442
rlabel metal2 719 -249 719 -249 0 net=7137
rlabel metal2 86 -251 86 -251 0 net=3411
rlabel metal2 516 -251 516 -251 0 net=478
rlabel metal2 58 -253 58 -253 0 net=2273
rlabel metal2 163 -253 163 -253 0 net=2447
rlabel metal2 327 -253 327 -253 0 net=4497
rlabel metal2 695 -253 695 -253 0 net=5103
rlabel metal2 58 -255 58 -255 0 net=1559
rlabel metal2 345 -255 345 -255 0 net=2555
rlabel metal2 534 -255 534 -255 0 net=7998
rlabel metal2 23 -257 23 -257 0 net=3959
rlabel metal2 359 -257 359 -257 0 net=2543
rlabel metal2 534 -257 534 -257 0 net=3591
rlabel metal2 163 -259 163 -259 0 net=3263
rlabel metal2 576 -259 576 -259 0 net=7842
rlabel metal2 191 -261 191 -261 0 net=1694
rlabel metal2 618 -261 618 -261 0 net=4777
rlabel metal2 737 -261 737 -261 0 net=6103
rlabel metal2 33 -263 33 -263 0 net=1199
rlabel metal2 562 -263 562 -263 0 net=4227
rlabel metal2 625 -263 625 -263 0 net=4851
rlabel metal2 744 -263 744 -263 0 net=6211
rlabel metal2 541 -265 541 -265 0 net=4371
rlabel metal2 583 -265 583 -265 0 net=4669
rlabel metal2 758 -265 758 -265 0 net=7235
rlabel metal2 380 -267 380 -267 0 net=2580
rlabel metal2 611 -267 611 -267 0 net=4769
rlabel metal2 667 -267 667 -267 0 net=5075
rlabel metal2 884 -267 884 -267 0 net=6813
rlabel metal2 121 -269 121 -269 0 net=3301
rlabel metal2 527 -269 527 -269 0 net=4179
rlabel metal2 698 -269 698 -269 0 net=5563
rlabel metal2 121 -271 121 -271 0 net=3757
rlabel metal2 499 -271 499 -271 0 net=3561
rlabel metal2 541 -271 541 -271 0 net=7393
rlabel metal2 142 -273 142 -273 0 net=6093
rlabel metal2 114 -275 114 -275 0 net=1585
rlabel metal2 296 -275 296 -275 0 net=3345
rlabel metal2 702 -275 702 -275 0 net=6125
rlabel metal2 114 -277 114 -277 0 net=3739
rlabel metal2 296 -277 296 -277 0 net=3207
rlabel metal2 705 -277 705 -277 0 net=7456
rlabel metal2 135 -279 135 -279 0 net=2003
rlabel metal2 709 -279 709 -279 0 net=5601
rlabel metal2 352 -281 352 -281 0 net=4879
rlabel metal2 730 -281 730 -281 0 net=5923
rlabel metal2 93 -283 93 -283 0 net=1965
rlabel metal2 520 -283 520 -283 0 net=4631
rlabel metal2 758 -283 758 -283 0 net=7419
rlabel metal2 9 -285 9 -285 0 net=2372
rlabel metal2 478 -285 478 -285 0 net=3677
rlabel metal2 597 -285 597 -285 0 net=4549
rlabel metal2 765 -285 765 -285 0 net=5661
rlabel metal2 9 -287 9 -287 0 net=1907
rlabel metal2 184 -287 184 -287 0 net=1735
rlabel metal2 779 -287 779 -287 0 net=5901
rlabel metal2 184 -289 184 -289 0 net=2135
rlabel metal2 390 -289 390 -289 0 net=4975
rlabel metal2 779 -289 779 -289 0 net=4301
rlabel metal2 247 -291 247 -291 0 net=1453
rlabel metal2 450 -291 450 -291 0 net=3781
rlabel metal2 786 -291 786 -291 0 net=5933
rlabel metal2 254 -293 254 -293 0 net=1593
rlabel metal2 450 -293 450 -293 0 net=6010
rlabel metal2 856 -293 856 -293 0 net=7077
rlabel metal2 254 -295 254 -295 0 net=1683
rlabel metal2 646 -295 646 -295 0 net=5777
rlabel metal2 324 -297 324 -297 0 net=2684
rlabel metal2 569 -297 569 -297 0 net=4325
rlabel metal2 681 -297 681 -297 0 net=5607
rlabel metal2 68 -299 68 -299 0 net=2873
rlabel metal2 653 -299 653 -299 0 net=4455
rlabel metal2 723 -299 723 -299 0 net=5729
rlabel metal2 156 -301 156 -301 0 net=4555
rlabel metal2 653 -301 653 -301 0 net=4011
rlabel metal2 723 -301 723 -301 0 net=4517
rlabel metal2 149 -303 149 -303 0 net=3017
rlabel metal2 660 -303 660 -303 0 net=3419
rlabel metal2 772 -303 772 -303 0 net=5087
rlabel metal2 30 -305 30 -305 0 net=5021
rlabel metal2 54 -307 54 -307 0 net=1573
rlabel metal2 2 -318 2 -318 0 net=1198
rlabel metal2 65 -318 65 -318 0 net=2275
rlabel metal2 93 -318 93 -318 0 net=2448
rlabel metal2 264 -318 264 -318 0 net=1594
rlabel metal2 285 -318 285 -318 0 net=8321
rlabel metal2 1500 -318 1500 -318 0 net=6321
rlabel metal2 1500 -318 1500 -318 0 net=6321
rlabel metal2 2 -320 2 -320 0 net=3477
rlabel metal2 58 -320 58 -320 0 net=1561
rlabel metal2 310 -320 310 -320 0 net=1203
rlabel metal2 471 -320 471 -320 0 net=3258
rlabel metal2 586 -320 586 -320 0 net=7414
rlabel metal2 1101 -320 1101 -320 0 net=8061
rlabel metal2 1178 -320 1178 -320 0 net=3746
rlabel metal2 9 -322 9 -322 0 net=1909
rlabel metal2 37 -322 37 -322 0 net=262
rlabel metal2 604 -322 604 -322 0 net=4229
rlabel metal2 681 -322 681 -322 0 net=4457
rlabel metal2 681 -322 681 -322 0 net=4457
rlabel metal2 688 -322 688 -322 0 net=4499
rlabel metal2 688 -322 688 -322 0 net=4499
rlabel metal2 695 -322 695 -322 0 net=7809
rlabel metal2 1115 -322 1115 -322 0 net=8203
rlabel metal2 9 -324 9 -324 0 net=3269
rlabel metal2 317 -324 317 -324 0 net=3346
rlabel metal2 527 -324 527 -324 0 net=3563
rlabel metal2 702 -324 702 -324 0 net=6435
rlabel metal2 16 -326 16 -326 0 net=4136
rlabel metal2 93 -326 93 -326 0 net=2871
rlabel metal2 184 -326 184 -326 0 net=2136
rlabel metal2 702 -326 702 -326 0 net=4551
rlabel metal2 758 -326 758 -326 0 net=6094
rlabel metal2 912 -326 912 -326 0 net=6045
rlabel metal2 912 -326 912 -326 0 net=6045
rlabel metal2 961 -326 961 -326 0 net=8319
rlabel metal2 16 -328 16 -328 0 net=1925
rlabel metal2 327 -328 327 -328 0 net=1736
rlabel metal2 667 -328 667 -328 0 net=4881
rlabel metal2 842 -328 842 -328 0 net=5565
rlabel metal2 842 -328 842 -328 0 net=5565
rlabel metal2 856 -328 856 -328 0 net=5609
rlabel metal2 856 -328 856 -328 0 net=5609
rlabel metal2 863 -328 863 -328 0 net=5663
rlabel metal2 863 -328 863 -328 0 net=5663
rlabel metal2 884 -328 884 -328 0 net=5935
rlabel metal2 1031 -328 1031 -328 0 net=7395
rlabel metal2 1129 -328 1129 -328 0 net=8285
rlabel metal2 26 -330 26 -330 0 net=1200
rlabel metal2 198 -330 198 -330 0 net=1276
rlabel metal2 359 -330 359 -330 0 net=823
rlabel metal2 709 -330 709 -330 0 net=4519
rlabel metal2 891 -330 891 -330 0 net=5903
rlabel metal2 996 -330 996 -330 0 net=7079
rlabel metal2 1052 -330 1052 -330 0 net=7861
rlabel metal2 1136 -330 1136 -330 0 net=8355
rlabel metal2 37 -332 37 -332 0 net=6234
rlabel metal2 1087 -332 1087 -332 0 net=7941
rlabel metal2 44 -334 44 -334 0 net=467
rlabel metal2 61 -334 61 -334 0 net=1885
rlabel metal2 254 -334 254 -334 0 net=1685
rlabel metal2 394 -334 394 -334 0 net=2844
rlabel metal2 422 -334 422 -334 0 net=3782
rlabel metal2 485 -334 485 -334 0 net=3759
rlabel metal2 653 -334 653 -334 0 net=4013
rlabel metal2 765 -334 765 -334 0 net=4977
rlabel metal2 1024 -334 1024 -334 0 net=7237
rlabel metal2 1094 -334 1094 -334 0 net=8023
rlabel metal2 68 -336 68 -336 0 net=4632
rlabel metal2 786 -336 786 -336 0 net=5779
rlabel metal2 947 -336 947 -336 0 net=6309
rlabel metal2 72 -338 72 -338 0 net=1278
rlabel metal2 107 -338 107 -338 0 net=1545
rlabel metal2 121 -338 121 -338 0 net=4140
rlabel metal2 625 -338 625 -338 0 net=4771
rlabel metal2 786 -338 786 -338 0 net=5105
rlabel metal2 940 -338 940 -338 0 net=6213
rlabel metal2 982 -338 982 -338 0 net=6993
rlabel metal2 1045 -338 1045 -338 0 net=7629
rlabel metal2 75 -340 75 -340 0 net=8264
rlabel metal2 79 -342 79 -342 0 net=6953
rlabel metal2 1122 -342 1122 -342 0 net=8239
rlabel metal2 82 -344 82 -344 0 net=2824
rlabel metal2 1073 -344 1073 -344 0 net=7919
rlabel metal2 107 -346 107 -346 0 net=2005
rlabel metal2 156 -346 156 -346 0 net=3018
rlabel metal2 471 -346 471 -346 0 net=3413
rlabel metal2 499 -346 499 -346 0 net=4372
rlabel metal2 569 -346 569 -346 0 net=4557
rlabel metal2 814 -346 814 -346 0 net=5259
rlabel metal2 898 -346 898 -346 0 net=5925
rlabel metal2 968 -346 968 -346 0 net=6701
rlabel metal2 1017 -346 1017 -346 0 net=7205
rlabel metal2 163 -348 163 -348 0 net=3265
rlabel metal2 516 -348 516 -348 0 net=5867
rlabel metal2 954 -348 954 -348 0 net=6475
rlabel metal2 975 -348 975 -348 0 net=6835
rlabel metal2 1038 -348 1038 -348 0 net=7421
rlabel metal2 96 -350 96 -350 0 net=5975
rlabel metal2 1003 -350 1003 -350 0 net=7139
rlabel metal2 100 -352 100 -352 0 net=2221
rlabel metal2 177 -352 177 -352 0 net=3953
rlabel metal2 303 -352 303 -352 0 net=1947
rlabel metal2 331 -352 331 -352 0 net=3135
rlabel metal2 429 -352 429 -352 0 net=3905
rlabel metal2 555 -352 555 -352 0 net=4143
rlabel metal2 625 -352 625 -352 0 net=3843
rlabel metal2 653 -352 653 -352 0 net=4361
rlabel metal2 800 -352 800 -352 0 net=5077
rlabel metal2 926 -352 926 -352 0 net=6127
rlabel metal2 51 -354 51 -354 0 net=2665
rlabel metal2 114 -354 114 -354 0 net=3740
rlabel metal2 128 -354 128 -354 0 net=2207
rlabel metal2 191 -354 191 -354 0 net=1327
rlabel metal2 219 -354 219 -354 0 net=1499
rlabel metal2 282 -354 282 -354 0 net=3527
rlabel metal2 380 -354 380 -354 0 net=3303
rlabel metal2 509 -354 509 -354 0 net=4187
rlabel metal2 674 -354 674 -354 0 net=4303
rlabel metal2 800 -354 800 -354 0 net=5037
rlabel metal2 72 -356 72 -356 0 net=4633
rlabel metal2 128 -356 128 -356 0 net=4181
rlabel metal2 779 -356 779 -356 0 net=5089
rlabel metal2 919 -356 919 -356 0 net=6105
rlabel metal2 933 -356 933 -356 0 net=6815
rlabel metal2 142 -358 142 -358 0 net=1587
rlabel metal2 303 -358 303 -358 0 net=1967
rlabel metal2 366 -358 366 -358 0 net=2545
rlabel metal2 397 -358 397 -358 0 net=6990
rlabel metal2 86 -360 86 -360 0 net=2063
rlabel metal2 198 -360 198 -360 0 net=1151
rlabel metal2 212 -360 212 -360 0 net=1613
rlabel metal2 772 -360 772 -360 0 net=5023
rlabel metal2 849 -360 849 -360 0 net=5603
rlabel metal2 1010 -360 1010 -360 0 net=7683
rlabel metal2 149 -362 149 -362 0 net=1575
rlabel metal2 289 -362 289 -362 0 net=3961
rlabel metal2 366 -362 366 -362 0 net=2993
rlabel metal2 772 -362 772 -362 0 net=5033
rlabel metal2 828 -362 828 -362 0 net=5287
rlabel metal2 870 -362 870 -362 0 net=5811
rlabel metal2 1010 -362 1010 -362 0 net=8073
rlabel metal2 79 -364 79 -364 0 net=5403
rlabel metal2 149 -366 149 -366 0 net=1455
rlabel metal2 289 -366 289 -366 0 net=187
rlabel metal2 569 -366 569 -366 0 net=4934
rlabel metal2 247 -368 247 -368 0 net=1649
rlabel metal2 373 -368 373 -368 0 net=3679
rlabel metal2 583 -368 583 -368 0 net=6343
rlabel metal2 835 -368 835 -368 0 net=5317
rlabel metal2 23 -370 23 -370 0 net=5421
rlabel metal2 23 -372 23 -372 0 net=841
rlabel metal2 261 -372 261 -372 0 net=1657
rlabel metal2 387 -372 387 -372 0 net=7501
rlabel metal2 261 -374 261 -374 0 net=3240
rlabel metal2 513 -374 513 -374 0 net=4209
rlabel metal2 583 -374 583 -374 0 net=3421
rlabel metal2 751 -374 751 -374 0 net=5731
rlabel metal2 331 -376 331 -376 0 net=2173
rlabel metal2 737 -376 737 -376 0 net=4853
rlabel metal2 345 -378 345 -378 0 net=2557
rlabel metal2 401 -378 401 -378 0 net=2309
rlabel metal2 401 -378 401 -378 0 net=2309
rlabel metal2 408 -378 408 -378 0 net=6445
rlabel metal2 51 -380 51 -380 0 net=3401
rlabel metal2 415 -380 415 -380 0 net=2925
rlabel metal2 436 -380 436 -380 0 net=3071
rlabel metal2 296 -382 296 -382 0 net=3209
rlabel metal2 415 -382 415 -382 0 net=2913
rlabel metal2 124 -384 124 -384 0 net=1705
rlabel metal2 338 -384 338 -384 0 net=2875
rlabel metal2 450 -384 450 -384 0 net=2931
rlabel metal2 464 -384 464 -384 0 net=3435
rlabel metal2 506 -384 506 -384 0 net=4670
rlabel metal2 124 -386 124 -386 0 net=3163
rlabel metal2 338 -386 338 -386 0 net=3697
rlabel metal2 579 -386 579 -386 0 net=4647
rlabel metal2 324 -388 324 -388 0 net=3443
rlabel metal2 590 -388 590 -388 0 net=7557
rlabel metal2 240 -390 240 -390 0 net=2113
rlabel metal2 443 -390 443 -390 0 net=3089
rlabel metal2 464 -390 464 -390 0 net=4309
rlabel metal2 520 -390 520 -390 0 net=3593
rlabel metal2 611 -390 611 -390 0 net=4327
rlabel metal2 716 -390 716 -390 0 net=4779
rlabel metal2 58 -392 58 -392 0 net=2319
rlabel metal2 411 -392 411 -392 0 net=4581
rlabel metal2 170 -394 170 -394 0 net=4377
rlabel metal2 534 -394 534 -394 0 net=3805
rlabel metal2 639 -394 639 -394 0 net=4287
rlabel metal2 26 -396 26 -396 0 net=3709
rlabel metal2 254 -396 254 -396 0 net=2509
rlabel metal2 565 -396 565 -396 0 net=180
rlabel metal2 23 -407 23 -407 0 net=7502
rlabel metal2 1129 -407 1129 -407 0 net=7943
rlabel metal2 1500 -407 1500 -407 0 net=6323
rlabel metal2 1500 -407 1500 -407 0 net=6323
rlabel metal2 23 -409 23 -409 0 net=2685
rlabel metal2 331 -409 331 -409 0 net=2174
rlabel metal2 541 -409 541 -409 0 net=3565
rlabel metal2 541 -409 541 -409 0 net=3565
rlabel metal2 548 -409 548 -409 0 net=8062
rlabel metal2 1209 -409 1209 -409 0 net=6867
rlabel metal2 26 -411 26 -411 0 net=6128
rlabel metal2 1017 -411 1017 -411 0 net=6837
rlabel metal2 30 -413 30 -413 0 net=1910
rlabel metal2 75 -413 75 -413 0 net=3031
rlabel metal2 128 -413 128 -413 0 net=4182
rlabel metal2 408 -413 408 -413 0 net=2926
rlabel metal2 460 -413 460 -413 0 net=5812
rlabel metal2 975 -413 975 -413 0 net=5909
rlabel metal2 30 -415 30 -415 0 net=5926
rlabel metal2 1038 -415 1038 -415 0 net=7141
rlabel metal2 1136 -415 1136 -415 0 net=8025
rlabel metal2 40 -417 40 -417 0 net=3528
rlabel metal2 331 -417 331 -417 0 net=4363
rlabel metal2 663 -417 663 -417 0 net=8204
rlabel metal2 44 -419 44 -419 0 net=3954
rlabel metal2 201 -419 201 -419 0 net=1576
rlabel metal2 261 -419 261 -419 0 net=2558
rlabel metal2 401 -419 401 -419 0 net=2311
rlabel metal2 471 -419 471 -419 0 net=3415
rlabel metal2 551 -419 551 -419 0 net=5024
rlabel metal2 814 -419 814 -419 0 net=5261
rlabel metal2 870 -419 870 -419 0 net=5733
rlabel metal2 968 -419 968 -419 0 net=6477
rlabel metal2 1045 -419 1045 -419 0 net=7207
rlabel metal2 1143 -419 1143 -419 0 net=8241
rlabel metal2 2 -421 2 -421 0 net=3479
rlabel metal2 58 -421 58 -421 0 net=2277
rlabel metal2 79 -421 79 -421 0 net=5323
rlabel metal2 961 -421 961 -421 0 net=6447
rlabel metal2 1059 -421 1059 -421 0 net=7397
rlabel metal2 1150 -421 1150 -421 0 net=8287
rlabel metal2 9 -423 9 -423 0 net=3271
rlabel metal2 86 -423 86 -423 0 net=1359
rlabel metal2 198 -423 198 -423 0 net=1153
rlabel metal2 261 -423 261 -423 0 net=3681
rlabel metal2 401 -423 401 -423 0 net=4329
rlabel metal2 625 -423 625 -423 0 net=3845
rlabel metal2 670 -423 670 -423 0 net=6310
rlabel metal2 1066 -423 1066 -423 0 net=7423
rlabel metal2 1157 -423 1157 -423 0 net=8357
rlabel metal2 61 -425 61 -425 0 net=7697
rlabel metal2 65 -427 65 -427 0 net=4211
rlabel metal2 562 -427 562 -427 0 net=5318
rlabel metal2 898 -427 898 -427 0 net=5869
rlabel metal2 982 -427 982 -427 0 net=6703
rlabel metal2 1073 -427 1073 -427 0 net=7559
rlabel metal2 47 -429 47 -429 0 net=5283
rlabel metal2 884 -429 884 -429 0 net=5937
rlabel metal2 905 -429 905 -429 0 net=5905
rlabel metal2 1003 -429 1003 -429 0 net=6817
rlabel metal2 1080 -429 1080 -429 0 net=7685
rlabel metal2 86 -431 86 -431 0 net=1588
rlabel metal2 275 -431 275 -431 0 net=1563
rlabel metal2 411 -431 411 -431 0 net=4310
rlabel metal2 478 -431 478 -431 0 net=3266
rlabel metal2 520 -431 520 -431 0 net=3595
rlabel metal2 569 -431 569 -431 0 net=5604
rlabel metal2 1003 -431 1003 -431 0 net=8075
rlabel metal2 89 -433 89 -433 0 net=6099
rlabel metal2 89 -435 89 -435 0 net=5078
rlabel metal2 828 -435 828 -435 0 net=5405
rlabel metal2 989 -435 989 -435 0 net=6995
rlabel metal2 93 -437 93 -437 0 net=2872
rlabel metal2 138 -437 138 -437 0 net=8322
rlabel metal2 72 -439 72 -439 0 net=1331
rlabel metal2 100 -439 100 -439 0 net=2667
rlabel metal2 422 -439 422 -439 0 net=3137
rlabel metal2 478 -439 478 -439 0 net=4883
rlabel metal2 772 -439 772 -439 0 net=5035
rlabel metal2 835 -439 835 -439 0 net=5423
rlabel metal2 1122 -439 1122 -439 0 net=7921
rlabel metal2 33 -441 33 -441 0 net=4623
rlabel metal2 779 -441 779 -441 0 net=5091
rlabel metal2 849 -441 849 -441 0 net=5289
rlabel metal2 1031 -441 1031 -441 0 net=7081
rlabel metal2 100 -443 100 -443 0 net=2065
rlabel metal2 145 -443 145 -443 0 net=5171
rlabel metal2 863 -443 863 -443 0 net=5665
rlabel metal2 107 -445 107 -445 0 net=2007
rlabel metal2 142 -445 142 -445 0 net=2208
rlabel metal2 198 -445 198 -445 0 net=3444
rlabel metal2 590 -445 590 -445 0 net=672
rlabel metal2 698 -445 698 -445 0 net=6131
rlabel metal2 107 -447 107 -447 0 net=5303
rlabel metal2 156 -449 156 -449 0 net=3165
rlabel metal2 572 -449 572 -449 0 net=5269
rlabel metal2 163 -451 163 -451 0 net=2223
rlabel metal2 338 -451 338 -451 0 net=3699
rlabel metal2 576 -451 576 -451 0 net=3761
rlabel metal2 632 -451 632 -451 0 net=4189
rlabel metal2 705 -451 705 -451 0 net=8320
rlabel metal2 170 -453 170 -453 0 net=3711
rlabel metal2 593 -453 593 -453 0 net=3072
rlabel metal2 716 -453 716 -453 0 net=4583
rlabel metal2 793 -453 793 -453 0 net=6345
rlabel metal2 1101 -453 1101 -453 0 net=7811
rlabel metal2 149 -455 149 -455 0 net=1457
rlabel metal2 184 -455 184 -455 0 net=1205
rlabel metal2 338 -455 338 -455 0 net=3437
rlabel metal2 509 -455 509 -455 0 net=4772
rlabel metal2 800 -455 800 -455 0 net=5039
rlabel metal2 114 -457 114 -457 0 net=4635
rlabel metal2 814 -457 814 -457 0 net=6107
rlabel metal2 114 -459 114 -459 0 net=1811
rlabel metal2 310 -459 310 -459 0 net=1949
rlabel metal2 345 -459 345 -459 0 net=3211
rlabel metal2 856 -459 856 -459 0 net=5611
rlabel metal2 51 -461 51 -461 0 net=3403
rlabel metal2 296 -461 296 -461 0 net=1707
rlabel metal2 373 -461 373 -461 0 net=2933
rlabel metal2 457 -461 457 -461 0 net=3091
rlabel metal2 485 -461 485 -461 0 net=3305
rlabel metal2 520 -461 520 -461 0 net=3423
rlabel metal2 597 -461 597 -461 0 net=4145
rlabel metal2 642 -461 642 -461 0 net=5943
rlabel metal2 51 -463 51 -463 0 net=2547
rlabel metal2 422 -463 422 -463 0 net=4465
rlabel metal2 149 -465 149 -465 0 net=2321
rlabel metal2 268 -465 268 -465 0 net=1659
rlabel metal2 296 -465 296 -465 0 net=3929
rlabel metal2 425 -465 425 -465 0 net=6779
rlabel metal2 212 -467 212 -467 0 net=1615
rlabel metal2 366 -467 366 -467 0 net=2995
rlabel metal2 457 -467 457 -467 0 net=4153
rlabel metal2 597 -467 597 -467 0 net=8323
rlabel metal2 212 -469 212 -469 0 net=1887
rlabel metal2 366 -469 366 -469 0 net=3309
rlabel metal2 534 -469 534 -469 0 net=3807
rlabel metal2 600 -469 600 -469 0 net=4978
rlabel metal2 219 -471 219 -471 0 net=2115
rlabel metal2 380 -471 380 -471 0 net=6827
rlabel metal2 226 -473 226 -473 0 net=1501
rlabel metal2 303 -473 303 -473 0 net=1969
rlabel metal2 436 -473 436 -473 0 net=2877
rlabel metal2 604 -473 604 -473 0 net=4231
rlabel metal2 646 -473 646 -473 0 net=4289
rlabel metal2 16 -475 16 -475 0 net=1927
rlabel metal2 317 -475 317 -475 0 net=1961
rlabel metal2 611 -475 611 -475 0 net=7238
rlabel metal2 16 -477 16 -477 0 net=1651
rlabel metal2 352 -477 352 -477 0 net=3963
rlabel metal2 527 -477 527 -477 0 net=3907
rlabel metal2 614 -477 614 -477 0 net=6655
rlabel metal2 82 -479 82 -479 0 net=4183
rlabel metal2 681 -479 681 -479 0 net=4459
rlabel metal2 737 -479 737 -479 0 net=4649
rlabel metal2 912 -479 912 -479 0 net=6047
rlabel metal2 1024 -479 1024 -479 0 net=6955
rlabel metal2 159 -481 159 -481 0 net=5483
rlabel metal2 947 -481 947 -481 0 net=6215
rlabel metal2 191 -483 191 -483 0 net=1329
rlabel metal2 233 -483 233 -483 0 net=2473
rlabel metal2 499 -483 499 -483 0 net=4291
rlabel metal2 751 -483 751 -483 0 net=4855
rlabel metal2 891 -483 891 -483 0 net=5781
rlabel metal2 135 -485 135 -485 0 net=1547
rlabel metal2 254 -485 254 -485 0 net=2511
rlabel metal2 527 -485 527 -485 0 net=7019
rlabel metal2 135 -487 135 -487 0 net=5976
rlabel metal2 37 -489 37 -489 0 net=5831
rlabel metal2 37 -491 37 -491 0 net=455
rlabel metal2 163 -491 163 -491 0 net=1899
rlabel metal2 565 -491 565 -491 0 net=4509
rlabel metal2 842 -491 842 -491 0 net=5567
rlabel metal2 352 -493 352 -493 0 net=1687
rlabel metal2 618 -493 618 -493 0 net=4305
rlabel metal2 702 -493 702 -493 0 net=4553
rlabel metal2 786 -493 786 -493 0 net=5107
rlabel metal2 110 -495 110 -495 0 net=2237
rlabel metal2 415 -495 415 -495 0 net=2914
rlabel metal2 730 -495 730 -495 0 net=4559
rlabel metal2 415 -497 415 -497 0 net=6436
rlabel metal2 502 -499 502 -499 0 net=7323
rlabel metal2 688 -499 688 -499 0 net=4501
rlabel metal2 1094 -499 1094 -499 0 net=7631
rlabel metal2 9 -501 9 -501 0 net=1805
rlabel metal2 688 -501 688 -501 0 net=4015
rlabel metal2 1094 -501 1094 -501 0 net=7863
rlabel metal2 723 -503 723 -503 0 net=4781
rlabel metal2 1115 -503 1115 -503 0 net=4979
rlabel metal2 667 -505 667 -505 0 net=7931
rlabel metal2 660 -507 660 -507 0 net=4065
rlabel metal2 709 -507 709 -507 0 net=4521
rlabel metal2 443 -509 443 -509 0 net=4379
rlabel metal2 443 -511 443 -511 0 net=3019
rlabel metal2 660 -511 660 -511 0 net=8387
rlabel metal2 2 -522 2 -522 0 net=6100
rlabel metal2 1248 -522 1248 -522 0 net=8325
rlabel metal2 1395 -522 1395 -522 0 net=6869
rlabel metal2 1500 -522 1500 -522 0 net=6325
rlabel metal2 2 -524 2 -524 0 net=1641
rlabel metal2 600 -524 600 -524 0 net=7049
rlabel metal2 16 -526 16 -526 0 net=1652
rlabel metal2 261 -526 261 -526 0 net=3682
rlabel metal2 460 -526 460 -526 0 net=5324
rlabel metal2 1003 -526 1003 -526 0 net=8077
rlabel metal2 30 -528 30 -528 0 net=3809
rlabel metal2 635 -528 635 -528 0 net=4650
rlabel metal2 828 -528 828 -528 0 net=5173
rlabel metal2 940 -528 940 -528 0 net=5735
rlabel metal2 1087 -528 1087 -528 0 net=6957
rlabel metal2 1087 -528 1087 -528 0 net=6957
rlabel metal2 1094 -528 1094 -528 0 net=7865
rlabel metal2 33 -530 33 -530 0 net=705
rlabel metal2 75 -530 75 -530 0 net=2116
rlabel metal2 226 -530 226 -530 0 net=1330
rlabel metal2 425 -530 425 -530 0 net=413
rlabel metal2 639 -530 639 -530 0 net=3847
rlabel metal2 639 -530 639 -530 0 net=3847
rlabel metal2 660 -530 660 -530 0 net=6108
rlabel metal2 870 -530 870 -530 0 net=5291
rlabel metal2 1024 -530 1024 -530 0 net=6217
rlabel metal2 1150 -530 1150 -530 0 net=7425
rlabel metal2 1255 -530 1255 -530 0 net=8359
rlabel metal2 40 -532 40 -532 0 net=6838
rlabel metal2 1213 -532 1213 -532 0 net=7945
rlabel metal2 40 -534 40 -534 0 net=6780
rlabel metal2 1080 -534 1080 -534 0 net=6829
rlabel metal2 1157 -534 1157 -534 0 net=7561
rlabel metal2 1262 -534 1262 -534 0 net=8389
rlabel metal2 47 -536 47 -536 0 net=558
rlabel metal2 226 -536 226 -536 0 net=1661
rlabel metal2 317 -536 317 -536 0 net=1962
rlabel metal2 614 -536 614 -536 0 net=5036
rlabel metal2 954 -536 954 -536 0 net=5833
rlabel metal2 1136 -536 1136 -536 0 net=7209
rlabel metal2 1220 -536 1220 -536 0 net=8027
rlabel metal2 72 -538 72 -538 0 net=2474
rlabel metal2 240 -538 240 -538 0 net=1503
rlabel metal2 271 -538 271 -538 0 net=3212
rlabel metal2 912 -538 912 -538 0 net=5485
rlabel metal2 996 -538 996 -538 0 net=6049
rlabel metal2 1164 -538 1164 -538 0 net=7633
rlabel metal2 1227 -538 1227 -538 0 net=8243
rlabel metal2 110 -540 110 -540 0 net=3306
rlabel metal2 499 -540 499 -540 0 net=6855
rlabel metal2 1171 -540 1171 -540 0 net=7687
rlabel metal2 114 -542 114 -542 0 net=1813
rlabel metal2 331 -542 331 -542 0 net=4364
rlabel metal2 520 -542 520 -542 0 net=3425
rlabel metal2 530 -542 530 -542 0 net=4554
rlabel metal2 779 -542 779 -542 0 net=4585
rlabel metal2 842 -542 842 -542 0 net=5109
rlabel metal2 933 -542 933 -542 0 net=5667
rlabel metal2 1017 -542 1017 -542 0 net=6133
rlabel metal2 1108 -542 1108 -542 0 net=7021
rlabel metal2 1178 -542 1178 -542 0 net=7699
rlabel metal2 114 -544 114 -544 0 net=8209
rlabel metal2 117 -546 117 -546 0 net=4330
rlabel metal2 408 -546 408 -546 0 net=2669
rlabel metal2 502 -546 502 -546 0 net=4290
rlabel metal2 1122 -546 1122 -546 0 net=7083
rlabel metal2 1185 -546 1185 -546 0 net=7813
rlabel metal2 135 -548 135 -548 0 net=6448
rlabel metal2 1192 -548 1192 -548 0 net=7923
rlabel metal2 121 -550 121 -550 0 net=3033
rlabel metal2 142 -550 142 -550 0 net=5284
rlabel metal2 898 -550 898 -550 0 net=5939
rlabel metal2 1199 -550 1199 -550 0 net=7933
rlabel metal2 121 -552 121 -552 0 net=1117
rlabel metal2 275 -552 275 -552 0 net=1349
rlabel metal2 401 -552 401 -552 0 net=3713
rlabel metal2 611 -552 611 -552 0 net=6763
rlabel metal2 1234 -552 1234 -552 0 net=8289
rlabel metal2 44 -554 44 -554 0 net=3481
rlabel metal2 625 -554 625 -554 0 net=4233
rlabel metal2 765 -554 765 -554 0 net=4637
rlabel metal2 142 -556 142 -556 0 net=1873
rlabel metal2 212 -556 212 -556 0 net=1889
rlabel metal2 338 -556 338 -556 0 net=3438
rlabel metal2 443 -556 443 -556 0 net=3021
rlabel metal2 509 -556 509 -556 0 net=6941
rlabel metal2 849 -556 849 -556 0 net=5041
rlabel metal2 968 -556 968 -556 0 net=5907
rlabel metal2 1129 -556 1129 -556 0 net=7143
rlabel metal2 58 -558 58 -558 0 net=2278
rlabel metal2 450 -558 450 -558 0 net=2997
rlabel metal2 457 -558 457 -558 0 net=3701
rlabel metal2 625 -558 625 -558 0 net=8041
rlabel metal2 37 -560 37 -560 0 net=3717
rlabel metal2 138 -560 138 -560 0 net=1515
rlabel metal2 233 -560 233 -560 0 net=1951
rlabel metal2 338 -560 338 -560 0 net=2935
rlabel metal2 450 -560 450 -560 0 net=3417
rlabel metal2 534 -560 534 -560 0 net=6191
rlabel metal2 79 -562 79 -562 0 net=3273
rlabel metal2 548 -562 548 -562 0 net=3167
rlabel metal2 628 -562 628 -562 0 net=6507
rlabel metal2 1143 -562 1143 -562 0 net=7399
rlabel metal2 65 -564 65 -564 0 net=4213
rlabel metal2 660 -564 660 -564 0 net=5425
rlabel metal2 1031 -564 1031 -564 0 net=6347
rlabel metal2 65 -566 65 -566 0 net=1901
rlabel metal2 170 -566 170 -566 0 net=1459
rlabel metal2 345 -566 345 -566 0 net=1708
rlabel metal2 464 -566 464 -566 0 net=3139
rlabel metal2 663 -566 663 -566 0 net=4385
rlabel metal2 786 -566 786 -566 0 net=4561
rlabel metal2 835 -566 835 -566 0 net=5093
rlabel metal2 1031 -566 1031 -566 0 net=8255
rlabel metal2 5 -568 5 -568 0 net=2157
rlabel metal2 481 -568 481 -568 0 net=5406
rlabel metal2 1052 -568 1052 -568 0 net=6657
rlabel metal2 23 -570 23 -570 0 net=2687
rlabel metal2 485 -570 485 -570 0 net=2879
rlabel metal2 670 -570 670 -570 0 net=4980
rlabel metal2 23 -572 23 -572 0 net=1971
rlabel metal2 348 -572 348 -572 0 net=5547
rlabel metal2 1010 -572 1010 -572 0 net=6997
rlabel metal2 1059 -572 1059 -572 0 net=6819
rlabel metal2 79 -574 79 -574 0 net=2067
rlabel metal2 107 -574 107 -574 0 net=5587
rlabel metal2 989 -574 989 -574 0 net=5945
rlabel metal2 96 -576 96 -576 0 net=2261
rlabel metal2 107 -576 107 -576 0 net=1369
rlabel metal2 163 -576 163 -576 0 net=1207
rlabel metal2 191 -576 191 -576 0 net=1549
rlabel metal2 240 -576 240 -576 0 net=1617
rlabel metal2 324 -576 324 -576 0 net=3093
rlabel metal2 506 -576 506 -576 0 net=4671
rlabel metal2 863 -576 863 -576 0 net=5271
rlabel metal2 947 -576 947 -576 0 net=5783
rlabel metal2 19 -578 19 -578 0 net=1033
rlabel metal2 191 -578 191 -578 0 net=1155
rlabel metal2 247 -578 247 -578 0 net=3811
rlabel metal2 268 -578 268 -578 0 net=439
rlabel metal2 723 -578 723 -578 0 net=4783
rlabel metal2 884 -578 884 -578 0 net=5305
rlabel metal2 145 -580 145 -580 0 net=4466
rlabel metal2 800 -580 800 -580 0 net=4857
rlabel metal2 926 -580 926 -580 0 net=5613
rlabel metal2 170 -582 170 -582 0 net=1895
rlabel metal2 250 -582 250 -582 0 net=4431
rlabel metal2 856 -582 856 -582 0 net=5263
rlabel metal2 86 -584 86 -584 0 net=4749
rlabel metal2 86 -586 86 -586 0 net=3597
rlabel metal2 618 -586 618 -586 0 net=4307
rlabel metal2 177 -588 177 -588 0 net=1361
rlabel metal2 177 -588 177 -588 0 net=1361
rlabel metal2 205 -588 205 -588 0 net=1929
rlabel metal2 352 -588 352 -588 0 net=1688
rlabel metal2 506 -588 506 -588 0 net=5910
rlabel metal2 282 -590 282 -590 0 net=2225
rlabel metal2 674 -590 674 -590 0 net=7325
rlabel metal2 51 -592 51 -592 0 net=2549
rlabel metal2 303 -592 303 -592 0 net=1337
rlabel metal2 359 -592 359 -592 0 net=2239
rlabel metal2 436 -592 436 -592 0 net=3965
rlabel metal2 681 -592 681 -592 0 net=4293
rlabel metal2 765 -592 765 -592 0 net=6479
rlabel metal2 359 -594 359 -594 0 net=1565
rlabel metal2 418 -594 418 -594 0 net=2625
rlabel metal2 471 -594 471 -594 0 net=3119
rlabel metal2 590 -594 590 -594 0 net=4155
rlabel metal2 688 -594 688 -594 0 net=4017
rlabel metal2 730 -594 730 -594 0 net=4503
rlabel metal2 891 -594 891 -594 0 net=5569
rlabel metal2 89 -596 89 -596 0 net=4945
rlabel metal2 961 -596 961 -596 0 net=5871
rlabel metal2 289 -598 289 -598 0 net=3404
rlabel metal2 418 -598 418 -598 0 net=6587
rlabel metal2 289 -600 289 -600 0 net=2513
rlabel metal2 443 -600 443 -600 0 net=3489
rlabel metal2 646 -600 646 -600 0 net=4185
rlabel metal2 737 -600 737 -600 0 net=4511
rlabel metal2 863 -600 863 -600 0 net=4753
rlabel metal2 373 -602 373 -602 0 net=1981
rlabel metal2 653 -602 653 -602 0 net=4191
rlabel metal2 744 -602 744 -602 0 net=4523
rlabel metal2 394 -604 394 -604 0 net=2313
rlabel metal2 478 -604 478 -604 0 net=4885
rlabel metal2 653 -604 653 -604 0 net=4381
rlabel metal2 716 -604 716 -604 0 net=4461
rlabel metal2 44 -606 44 -606 0 net=4103
rlabel metal2 747 -606 747 -606 0 net=5847
rlabel metal2 149 -608 149 -608 0 net=2323
rlabel metal2 541 -608 541 -608 0 net=3567
rlabel metal2 576 -608 576 -608 0 net=3763
rlabel metal2 667 -608 667 -608 0 net=4067
rlabel metal2 695 -608 695 -608 0 net=6704
rlabel metal2 37 -610 37 -610 0 net=3573
rlabel metal2 632 -610 632 -610 0 net=4147
rlabel metal2 772 -610 772 -610 0 net=4625
rlabel metal2 149 -612 149 -612 0 net=1229
rlabel metal2 390 -612 390 -612 0 net=5977
rlabel metal2 366 -614 366 -614 0 net=3311
rlabel metal2 632 -614 632 -614 0 net=4073
rlabel metal2 702 -614 702 -614 0 net=7387
rlabel metal2 156 -616 156 -616 0 net=4089
rlabel metal2 772 -616 772 -616 0 net=3463
rlabel metal2 128 -618 128 -618 0 net=2009
rlabel metal2 296 -618 296 -618 0 net=3931
rlabel metal2 667 -618 667 -618 0 net=5801
rlabel metal2 9 -620 9 -620 0 net=1807
rlabel metal2 9 -622 9 -622 0 net=3909
rlabel metal2 93 -624 93 -624 0 net=1333
rlabel metal2 604 -624 604 -624 0 net=3623
rlabel metal2 51 -626 51 -626 0 net=1279
rlabel metal2 16 -637 16 -637 0 net=2373
rlabel metal2 16 -637 16 -637 0 net=2373
rlabel metal2 37 -637 37 -637 0 net=3095
rlabel metal2 383 -637 383 -637 0 net=4186
rlabel metal2 747 -637 747 -637 0 net=5668
rlabel metal2 1034 -637 1034 -637 0 net=8360
rlabel metal2 1472 -637 1472 -637 0 net=6871
rlabel metal2 2 -639 2 -639 0 net=1643
rlabel metal2 387 -639 387 -639 0 net=3418
rlabel metal2 506 -639 506 -639 0 net=3464
rlabel metal2 807 -639 807 -639 0 net=4513
rlabel metal2 1507 -639 1507 -639 0 net=6327
rlabel metal2 5 -641 5 -641 0 net=8191
rlabel metal2 44 -643 44 -643 0 net=4638
rlabel metal2 1206 -643 1206 -643 0 net=7635
rlabel metal2 44 -645 44 -645 0 net=1953
rlabel metal2 282 -645 282 -645 0 net=2550
rlabel metal2 387 -645 387 -645 0 net=3313
rlabel metal2 544 -645 544 -645 0 net=8097
rlabel metal2 47 -647 47 -647 0 net=2158
rlabel metal2 443 -647 443 -647 0 net=4214
rlabel metal2 614 -647 614 -647 0 net=4234
rlabel metal2 807 -647 807 -647 0 net=5265
rlabel metal2 940 -647 940 -647 0 net=5293
rlabel metal2 1101 -647 1101 -647 0 net=6349
rlabel metal2 1255 -647 1255 -647 0 net=7701
rlabel metal2 30 -649 30 -649 0 net=3810
rlabel metal2 429 -649 429 -649 0 net=2325
rlabel metal2 446 -649 446 -649 0 net=8127
rlabel metal2 30 -651 30 -651 0 net=3587
rlabel metal2 408 -651 408 -651 0 net=2241
rlabel metal2 471 -651 471 -651 0 net=3120
rlabel metal2 870 -651 870 -651 0 net=4785
rlabel metal2 1059 -651 1059 -651 0 net=5947
rlabel metal2 1150 -651 1150 -651 0 net=6831
rlabel metal2 1262 -651 1262 -651 0 net=7815
rlabel metal2 65 -653 65 -653 0 net=1902
rlabel metal2 100 -653 100 -653 0 net=2262
rlabel metal2 191 -653 191 -653 0 net=1157
rlabel metal2 191 -653 191 -653 0 net=1157
rlabel metal2 233 -653 233 -653 0 net=2415
rlabel metal2 415 -653 415 -653 0 net=5426
rlabel metal2 663 -653 663 -653 0 net=8078
rlabel metal2 1346 -653 1346 -653 0 net=8257
rlabel metal2 65 -655 65 -655 0 net=1897
rlabel metal2 261 -655 261 -655 0 net=1505
rlabel metal2 296 -655 296 -655 0 net=1809
rlabel metal2 870 -655 870 -655 0 net=6219
rlabel metal2 1150 -655 1150 -655 0 net=7023
rlabel metal2 1227 -655 1227 -655 0 net=7389
rlabel metal2 1353 -655 1353 -655 0 net=8291
rlabel metal2 23 -657 23 -657 0 net=1973
rlabel metal2 296 -657 296 -657 0 net=2315
rlabel metal2 401 -657 401 -657 0 net=3715
rlabel metal2 1157 -657 1157 -657 0 net=6857
rlabel metal2 1283 -657 1283 -657 0 net=7867
rlabel metal2 23 -659 23 -659 0 net=3605
rlabel metal2 345 -659 345 -659 0 net=2689
rlabel metal2 506 -659 506 -659 0 net=4157
rlabel metal2 688 -659 688 -659 0 net=4069
rlabel metal2 688 -659 688 -659 0 net=4069
rlabel metal2 730 -659 730 -659 0 net=4193
rlabel metal2 744 -659 744 -659 0 net=7617
rlabel metal2 9 -661 9 -661 0 net=3911
rlabel metal2 702 -661 702 -661 0 net=4091
rlabel metal2 744 -661 744 -661 0 net=5908
rlabel metal2 1052 -661 1052 -661 0 net=6999
rlabel metal2 1290 -661 1290 -661 0 net=7925
rlabel metal2 79 -663 79 -663 0 net=2069
rlabel metal2 415 -663 415 -663 0 net=2177
rlabel metal2 628 -663 628 -663 0 net=4308
rlabel metal2 1171 -663 1171 -663 0 net=7085
rlabel metal2 1304 -663 1304 -663 0 net=7947
rlabel metal2 79 -665 79 -665 0 net=1119
rlabel metal2 128 -665 128 -665 0 net=1335
rlabel metal2 219 -665 219 -665 0 net=1815
rlabel metal2 348 -665 348 -665 0 net=2137
rlabel metal2 436 -665 436 -665 0 net=2627
rlabel metal2 509 -665 509 -665 0 net=3274
rlabel metal2 548 -665 548 -665 0 net=3169
rlabel metal2 597 -665 597 -665 0 net=4887
rlabel metal2 940 -665 940 -665 0 net=6483
rlabel metal2 1248 -665 1248 -665 0 net=7563
rlabel metal2 1360 -665 1360 -665 0 net=8327
rlabel metal2 58 -667 58 -667 0 net=3719
rlabel metal2 614 -667 614 -667 0 net=6311
rlabel metal2 1171 -667 1171 -667 0 net=7401
rlabel metal2 1297 -667 1297 -667 0 net=7935
rlabel metal2 1367 -667 1367 -667 0 net=8391
rlabel metal2 58 -669 58 -669 0 net=2010
rlabel metal2 268 -669 268 -669 0 net=7603
rlabel metal2 61 -671 61 -671 0 net=4645
rlabel metal2 1311 -671 1311 -671 0 net=8029
rlabel metal2 86 -673 86 -673 0 net=3599
rlabel metal2 436 -673 436 -673 0 net=3625
rlabel metal2 628 -673 628 -673 0 net=7050
rlabel metal2 1318 -673 1318 -673 0 net=8043
rlabel metal2 86 -675 86 -675 0 net=1891
rlabel metal2 359 -675 359 -675 0 net=1567
rlabel metal2 604 -675 604 -675 0 net=4075
rlabel metal2 702 -675 702 -675 0 net=4463
rlabel metal2 842 -675 842 -675 0 net=6943
rlabel metal2 1325 -675 1325 -675 0 net=8211
rlabel metal2 93 -677 93 -677 0 net=4709
rlabel metal2 635 -677 635 -677 0 net=5736
rlabel metal2 1010 -677 1010 -677 0 net=5785
rlabel metal2 1073 -677 1073 -677 0 net=6051
rlabel metal2 1129 -677 1129 -677 0 net=6659
rlabel metal2 1332 -677 1332 -677 0 net=8245
rlabel metal2 19 -679 19 -679 0 net=4831
rlabel metal2 1080 -679 1080 -679 0 net=6135
rlabel metal2 1143 -679 1143 -679 0 net=6821
rlabel metal2 72 -681 72 -681 0 net=6145
rlabel metal2 1199 -681 1199 -681 0 net=7145
rlabel metal2 72 -683 72 -683 0 net=592
rlabel metal2 747 -683 747 -683 0 net=6192
rlabel metal2 1199 -683 1199 -683 0 net=7427
rlabel metal2 96 -685 96 -685 0 net=6633
rlabel metal2 100 -687 100 -687 0 net=2226
rlabel metal2 761 -687 761 -687 0 net=6249
rlabel metal2 1213 -687 1213 -687 0 net=7211
rlabel metal2 114 -689 114 -689 0 net=1982
rlabel metal2 380 -689 380 -689 0 net=3703
rlabel metal2 478 -689 478 -689 0 net=5863
rlabel metal2 1108 -689 1108 -689 0 net=6509
rlabel metal2 1220 -689 1220 -689 0 net=7327
rlabel metal2 114 -691 114 -691 0 net=5174
rlabel metal2 943 -691 943 -691 0 net=7688
rlabel metal2 121 -693 121 -693 0 net=1375
rlabel metal2 618 -693 618 -693 0 net=7107
rlabel metal2 128 -695 128 -695 0 net=1993
rlabel metal2 425 -695 425 -695 0 net=3935
rlabel metal2 765 -695 765 -695 0 net=6481
rlabel metal2 135 -697 135 -697 0 net=3034
rlabel metal2 247 -697 247 -697 0 net=3813
rlabel metal2 359 -697 359 -697 0 net=2999
rlabel metal2 513 -697 513 -697 0 net=2881
rlabel metal2 779 -697 779 -697 0 net=4387
rlabel metal2 856 -697 856 -697 0 net=4751
rlabel metal2 12 -699 12 -699 0 net=4613
rlabel metal2 877 -699 877 -699 0 net=4859
rlabel metal2 1066 -699 1066 -699 0 net=5979
rlabel metal2 1136 -699 1136 -699 0 net=6765
rlabel metal2 107 -701 107 -701 0 net=1371
rlabel metal2 310 -701 310 -701 0 net=3427
rlabel metal2 537 -701 537 -701 0 net=6071
rlabel metal2 849 -701 849 -701 0 net=4673
rlabel metal2 919 -701 919 -701 0 net=5615
rlabel metal2 1017 -701 1017 -701 0 net=5803
rlabel metal2 1087 -701 1087 -701 0 net=6959
rlabel metal2 107 -703 107 -703 0 net=1619
rlabel metal2 313 -703 313 -703 0 net=2655
rlabel metal2 485 -703 485 -703 0 net=3023
rlabel metal2 499 -703 499 -703 0 net=2671
rlabel metal2 653 -703 653 -703 0 net=4383
rlabel metal2 149 -705 149 -705 0 net=1231
rlabel metal2 177 -705 177 -705 0 net=1363
rlabel metal2 317 -705 317 -705 0 net=4149
rlabel metal2 835 -705 835 -705 0 net=4627
rlabel metal2 1024 -705 1024 -705 0 net=5835
rlabel metal2 149 -707 149 -707 0 net=1421
rlabel metal2 639 -707 639 -707 0 net=3849
rlabel metal2 667 -707 667 -707 0 net=5495
rlabel metal2 1038 -707 1038 -707 0 net=5873
rlabel metal2 103 -709 103 -709 0 net=5887
rlabel metal2 667 -709 667 -709 0 net=4105
rlabel metal2 716 -709 716 -709 0 net=4505
rlabel metal2 814 -709 814 -709 0 net=4525
rlabel metal2 849 -709 849 -709 0 net=4947
rlabel metal2 947 -709 947 -709 0 net=5307
rlabel metal2 177 -711 177 -711 0 net=1035
rlabel metal2 338 -711 338 -711 0 net=2937
rlabel metal2 565 -711 565 -711 0 net=8265
rlabel metal2 184 -713 184 -713 0 net=1517
rlabel metal2 338 -713 338 -713 0 net=3967
rlabel metal2 709 -713 709 -713 0 net=4019
rlabel metal2 786 -713 786 -713 0 net=4433
rlabel metal2 814 -713 814 -713 0 net=4563
rlabel metal2 954 -713 954 -713 0 net=5487
rlabel metal2 163 -715 163 -715 0 net=1209
rlabel metal2 355 -715 355 -715 0 net=4999
rlabel metal2 961 -715 961 -715 0 net=7247
rlabel metal2 142 -717 142 -717 0 net=1875
rlabel metal2 355 -717 355 -717 0 net=3702
rlabel metal2 492 -717 492 -717 0 net=3785
rlabel metal2 786 -717 786 -717 0 net=6589
rlabel metal2 142 -719 142 -719 0 net=1443
rlabel metal2 366 -719 366 -719 0 net=3933
rlabel metal2 758 -719 758 -719 0 net=4295
rlabel metal2 75 -721 75 -721 0 net=929
rlabel metal2 373 -721 373 -721 0 net=3141
rlabel metal2 632 -721 632 -721 0 net=6377
rlabel metal2 898 -721 898 -721 0 net=5043
rlabel metal2 964 -721 964 -721 0 net=8153
rlabel metal2 289 -723 289 -723 0 net=2515
rlabel metal2 646 -723 646 -723 0 net=3765
rlabel metal2 758 -723 758 -723 0 net=5940
rlabel metal2 226 -725 226 -725 0 net=1663
rlabel metal2 457 -725 457 -725 0 net=3575
rlabel metal2 590 -725 590 -725 0 net=3491
rlabel metal2 821 -725 821 -725 0 net=4057
rlabel metal2 905 -725 905 -725 0 net=5095
rlabel metal2 968 -725 968 -725 0 net=5549
rlabel metal2 226 -727 226 -727 0 net=1461
rlabel metal2 499 -727 499 -727 0 net=2713
rlabel metal2 555 -727 555 -727 0 net=3569
rlabel metal2 611 -727 611 -727 0 net=6449
rlabel metal2 205 -729 205 -729 0 net=1931
rlabel metal2 534 -729 534 -729 0 net=3281
rlabel metal2 569 -729 569 -729 0 net=3483
rlabel metal2 611 -729 611 -729 0 net=6139
rlabel metal2 205 -731 205 -731 0 net=1351
rlabel metal2 562 -731 562 -731 0 net=4955
rlabel metal2 863 -731 863 -731 0 net=4755
rlabel metal2 905 -731 905 -731 0 net=5571
rlabel metal2 982 -731 982 -731 0 net=5589
rlabel metal2 117 -733 117 -733 0 net=4447
rlabel metal2 275 -735 275 -735 0 net=1339
rlabel metal2 366 -735 366 -735 0 net=5243
rlabel metal2 198 -737 198 -737 0 net=1551
rlabel metal2 380 -737 380 -737 0 net=2227
rlabel metal2 863 -737 863 -737 0 net=5273
rlabel metal2 51 -739 51 -739 0 net=1281
rlabel metal2 828 -739 828 -739 0 net=4587
rlabel metal2 51 -741 51 -741 0 net=1529
rlabel metal2 117 -741 117 -741 0 net=8009
rlabel metal2 912 -741 912 -741 0 net=5111
rlabel metal2 884 -743 884 -743 0 net=5849
rlabel metal2 842 -745 842 -745 0 net=4117
rlabel metal2 2 -756 2 -756 0 net=3716
rlabel metal2 2 -758 2 -758 0 net=4827
rlabel metal2 614 -758 614 -758 0 net=4514
rlabel metal2 9 -760 9 -760 0 net=3968
rlabel metal2 369 -760 369 -760 0 net=344
rlabel metal2 1066 -760 1066 -760 0 net=7249
rlabel metal2 1437 -760 1437 -760 0 net=8129
rlabel metal2 9 -762 9 -762 0 net=4807
rlabel metal2 649 -762 649 -762 0 net=4646
rlabel metal2 1458 -762 1458 -762 0 net=8193
rlabel metal2 12 -764 12 -764 0 net=5112
rlabel metal2 1066 -764 1066 -764 0 net=6511
rlabel metal2 1472 -764 1472 -764 0 net=8259
rlabel metal2 23 -766 23 -766 0 net=3606
rlabel metal2 310 -766 310 -766 0 net=3428
rlabel metal2 747 -766 747 -766 0 net=6889
rlabel metal2 16 -768 16 -768 0 net=2375
rlabel metal2 47 -768 47 -768 0 net=2516
rlabel metal2 653 -768 653 -768 0 net=3850
rlabel metal2 775 -768 775 -768 0 net=8392
rlabel metal2 16 -770 16 -770 0 net=1519
rlabel metal2 226 -770 226 -770 0 net=1462
rlabel metal2 394 -770 394 -770 0 net=1569
rlabel metal2 443 -770 443 -770 0 net=2327
rlabel metal2 443 -770 443 -770 0 net=2327
rlabel metal2 471 -770 471 -770 0 net=2629
rlabel metal2 471 -770 471 -770 0 net=2629
rlabel metal2 478 -770 478 -770 0 net=2657
rlabel metal2 478 -770 478 -770 0 net=2657
rlabel metal2 485 -770 485 -770 0 net=3025
rlabel metal2 499 -770 499 -770 0 net=2715
rlabel metal2 499 -770 499 -770 0 net=2715
rlabel metal2 509 -770 509 -770 0 net=4860
rlabel metal2 1164 -770 1164 -770 0 net=6313
rlabel metal2 58 -772 58 -772 0 net=5590
rlabel metal2 58 -774 58 -774 0 net=1121
rlabel metal2 117 -774 117 -774 0 net=3934
rlabel metal2 884 -774 884 -774 0 net=6822
rlabel metal2 51 -776 51 -776 0 net=1531
rlabel metal2 121 -776 121 -776 0 net=1377
rlabel metal2 324 -776 324 -776 0 net=1644
rlabel metal2 485 -776 485 -776 0 net=2673
rlabel metal2 534 -776 534 -776 0 net=5836
rlabel metal2 51 -778 51 -778 0 net=2317
rlabel metal2 324 -778 324 -778 0 net=1849
rlabel metal2 520 -778 520 -778 0 net=59
rlabel metal2 537 -778 537 -778 0 net=1810
rlabel metal2 887 -778 887 -778 0 net=8328
rlabel metal2 61 -780 61 -780 0 net=4832
rlabel metal2 1164 -780 1164 -780 0 net=7329
rlabel metal2 1332 -780 1332 -780 0 net=7565
rlabel metal2 1444 -780 1444 -780 0 net=8247
rlabel metal2 65 -782 65 -782 0 net=1898
rlabel metal2 520 -782 520 -782 0 net=4077
rlabel metal2 611 -782 611 -782 0 net=4757
rlabel metal2 940 -782 940 -782 0 net=8030
rlabel metal2 65 -784 65 -784 0 net=4151
rlabel metal2 338 -784 338 -784 0 net=1703
rlabel metal2 394 -784 394 -784 0 net=2071
rlabel metal2 422 -784 422 -784 0 net=3485
rlabel metal2 583 -784 583 -784 0 net=3721
rlabel metal2 618 -784 618 -784 0 net=4464
rlabel metal2 723 -784 723 -784 0 net=4435
rlabel metal2 856 -784 856 -784 0 net=4615
rlabel metal2 943 -784 943 -784 0 net=6832
rlabel metal2 72 -786 72 -786 0 net=7936
rlabel metal2 72 -788 72 -788 0 net=1975
rlabel metal2 296 -788 296 -788 0 net=1853
rlabel metal2 800 -788 800 -788 0 net=4059
rlabel metal2 856 -788 856 -788 0 net=5001
rlabel metal2 968 -788 968 -788 0 net=5949
rlabel metal2 1150 -788 1150 -788 0 net=7025
rlabel metal2 1360 -788 1360 -788 0 net=7927
rlabel metal2 75 -790 75 -790 0 net=4752
rlabel metal2 1199 -790 1199 -790 0 net=7429
rlabel metal2 1409 -790 1409 -790 0 net=8045
rlabel metal2 100 -792 100 -792 0 net=8079
rlabel metal2 1430 -792 1430 -792 0 net=8099
rlabel metal2 100 -794 100 -794 0 net=3001
rlabel metal2 401 -794 401 -794 0 net=2139
rlabel metal2 464 -794 464 -794 0 net=3705
rlabel metal2 597 -794 597 -794 0 net=5096
rlabel metal2 1017 -794 1017 -794 0 net=5497
rlabel metal2 1101 -794 1101 -794 0 net=6137
rlabel metal2 1199 -794 1199 -794 0 net=6661
rlabel metal2 1248 -794 1248 -794 0 net=7001
rlabel metal2 1451 -794 1451 -794 0 net=8155
rlabel metal2 114 -796 114 -796 0 net=4045
rlabel metal2 1465 -796 1465 -796 0 net=8213
rlabel metal2 114 -798 114 -798 0 net=1507
rlabel metal2 408 -798 408 -798 0 net=2179
rlabel metal2 464 -798 464 -798 0 net=4296
rlabel metal2 1129 -798 1129 -798 0 net=6451
rlabel metal2 1234 -798 1234 -798 0 net=6945
rlabel metal2 1283 -798 1283 -798 0 net=7147
rlabel metal2 1479 -798 1479 -798 0 net=8293
rlabel metal2 121 -800 121 -800 0 net=1037
rlabel metal2 184 -800 184 -800 0 net=1553
rlabel metal2 425 -800 425 -800 0 net=6299
rlabel metal2 1171 -800 1171 -800 0 net=7403
rlabel metal2 1500 -800 1500 -800 0 net=6328
rlabel metal2 131 -802 131 -802 0 net=1336
rlabel metal2 177 -802 177 -802 0 net=1211
rlabel metal2 226 -802 226 -802 0 net=2229
rlabel metal2 523 -802 523 -802 0 net=4628
rlabel metal2 1017 -802 1017 -802 0 net=6859
rlabel metal2 1269 -802 1269 -802 0 net=7109
rlabel metal2 1514 -802 1514 -802 0 net=6873
rlabel metal2 107 -804 107 -804 0 net=1621
rlabel metal2 205 -804 205 -804 0 net=1353
rlabel metal2 380 -804 380 -804 0 net=3283
rlabel metal2 569 -804 569 -804 0 net=4957
rlabel metal2 891 -804 891 -804 0 net=6379
rlabel metal2 1192 -804 1192 -804 0 net=6635
rlabel metal2 107 -806 107 -806 0 net=1817
rlabel metal2 236 -806 236 -806 0 net=3641
rlabel metal2 289 -806 289 -806 0 net=1665
rlabel metal2 436 -806 436 -806 0 net=3627
rlabel metal2 618 -806 618 -806 0 net=4889
rlabel metal2 989 -806 989 -806 0 net=5787
rlabel metal2 1115 -806 1115 -806 0 net=6053
rlabel metal2 1227 -806 1227 -806 0 net=7087
rlabel metal2 30 -808 30 -808 0 net=3589
rlabel metal2 30 -810 30 -810 0 net=2243
rlabel metal2 467 -810 467 -810 0 net=7315
rlabel metal2 135 -812 135 -812 0 net=831
rlabel metal2 695 -812 695 -812 0 net=3937
rlabel metal2 779 -812 779 -812 0 net=6073
rlabel metal2 135 -814 135 -814 0 net=1877
rlabel metal2 205 -814 205 -814 0 net=3003
rlabel metal2 138 -816 138 -816 0 net=132
rlabel metal2 779 -816 779 -816 0 net=4389
rlabel metal2 814 -816 814 -816 0 net=4565
rlabel metal2 905 -816 905 -816 0 net=5573
rlabel metal2 1038 -816 1038 -816 0 net=8267
rlabel metal2 93 -818 93 -818 0 net=4711
rlabel metal2 905 -818 905 -818 0 net=5045
rlabel metal2 1038 -818 1038 -818 0 net=5865
rlabel metal2 93 -820 93 -820 0 net=4159
rlabel metal2 534 -820 534 -820 0 net=3367
rlabel metal2 632 -820 632 -820 0 net=3767
rlabel metal2 681 -820 681 -820 0 net=3913
rlabel metal2 730 -820 730 -820 0 net=4195
rlabel metal2 786 -820 786 -820 0 net=6591
rlabel metal2 142 -822 142 -822 0 net=1445
rlabel metal2 429 -822 429 -822 0 net=3601
rlabel metal2 688 -822 688 -822 0 net=4071
rlabel metal2 758 -822 758 -822 0 net=5501
rlabel metal2 1045 -822 1045 -822 0 net=5875
rlabel metal2 86 -824 86 -824 0 net=1893
rlabel metal2 436 -824 436 -824 0 net=5049
rlabel metal2 919 -824 919 -824 0 net=5617
rlabel metal2 1080 -824 1080 -824 0 net=6141
rlabel metal2 86 -826 86 -826 0 net=4021
rlabel metal2 758 -826 758 -826 0 net=5267
rlabel metal2 919 -826 919 -826 0 net=5295
rlabel metal2 1087 -826 1087 -826 0 net=6485
rlabel metal2 103 -828 103 -828 0 net=3439
rlabel metal2 163 -828 163 -828 0 net=8439
rlabel metal2 212 -830 212 -830 0 net=2435
rlabel metal2 450 -830 450 -830 0 net=4507
rlabel metal2 793 -830 793 -830 0 net=4527
rlabel metal2 947 -830 947 -830 0 net=5453
rlabel metal2 1136 -830 1136 -830 0 net=6351
rlabel metal2 1206 -830 1206 -830 0 net=6767
rlabel metal2 219 -832 219 -832 0 net=2011
rlabel metal2 492 -832 492 -832 0 net=3787
rlabel metal2 709 -832 709 -832 0 net=5550
rlabel metal2 1241 -832 1241 -832 0 net=6961
rlabel metal2 240 -834 240 -834 0 net=1365
rlabel metal2 331 -834 331 -834 0 net=3815
rlabel metal2 506 -834 506 -834 0 net=628
rlabel metal2 1024 -834 1024 -834 0 net=5981
rlabel metal2 1276 -834 1276 -834 0 net=7391
rlabel metal2 233 -836 233 -836 0 net=2417
rlabel metal2 254 -836 254 -836 0 net=1933
rlabel metal2 541 -836 541 -836 0 net=4786
rlabel metal2 1108 -836 1108 -836 0 net=6147
rlabel metal2 191 -838 191 -838 0 net=1158
rlabel metal2 261 -838 261 -838 0 net=1509
rlabel metal2 667 -838 667 -838 0 net=4107
rlabel metal2 912 -838 912 -838 0 net=5851
rlabel metal2 1143 -838 1143 -838 0 net=7213
rlabel metal2 191 -840 191 -840 0 net=1341
rlabel metal2 331 -840 331 -840 0 net=3143
rlabel metal2 541 -840 541 -840 0 net=965
rlabel metal2 863 -840 863 -840 0 net=5275
rlabel metal2 999 -840 999 -840 0 net=7407
rlabel metal2 128 -842 128 -842 0 net=1995
rlabel metal2 373 -842 373 -842 0 net=2939
rlabel metal2 544 -842 544 -842 0 net=2882
rlabel metal2 1157 -842 1157 -842 0 net=6251
rlabel metal2 37 -844 37 -844 0 net=3097
rlabel metal2 548 -844 548 -844 0 net=3171
rlabel metal2 600 -844 600 -844 0 net=4393
rlabel metal2 838 -844 838 -844 0 net=6577
rlabel metal2 128 -846 128 -846 0 net=6482
rlabel metal2 198 -848 198 -848 0 net=1283
rlabel metal2 268 -848 268 -848 0 net=2691
rlabel metal2 530 -848 530 -848 0 net=1
rlabel metal2 551 -848 551 -848 0 net=4448
rlabel metal2 1353 -848 1353 -848 0 net=7605
rlabel metal2 198 -850 198 -850 0 net=1373
rlabel metal2 345 -850 345 -850 0 net=2281
rlabel metal2 562 -850 562 -850 0 net=5941
rlabel metal2 1367 -850 1367 -850 0 net=7619
rlabel metal2 44 -852 44 -852 0 net=1955
rlabel metal2 562 -852 562 -852 0 net=3571
rlabel metal2 639 -852 639 -852 0 net=5889
rlabel metal2 1374 -852 1374 -852 0 net=7637
rlabel metal2 44 -854 44 -854 0 net=7335
rlabel metal2 737 -854 737 -854 0 net=4093
rlabel metal2 765 -854 765 -854 0 net=4588
rlabel metal2 1381 -854 1381 -854 0 net=7703
rlabel metal2 166 -856 166 -856 0 net=3445
rlabel metal2 646 -856 646 -856 0 net=3493
rlabel metal2 737 -856 737 -856 0 net=4675
rlabel metal2 933 -856 933 -856 0 net=5309
rlabel metal2 1388 -856 1388 -856 0 net=7817
rlabel metal2 457 -858 457 -858 0 net=3577
rlabel metal2 1395 -858 1395 -858 0 net=7869
rlabel metal2 457 -860 457 -860 0 net=4384
rlabel metal2 1402 -860 1402 -860 0 net=7949
rlabel metal2 569 -862 569 -862 0 net=3683
rlabel metal2 625 -864 625 -864 0 net=5837
rlabel metal2 40 -866 40 -866 0 net=5877
rlabel metal2 646 -866 646 -866 0 net=7033
rlabel metal2 653 -868 653 -868 0 net=6165
rlabel metal2 656 -870 656 -870 0 net=6220
rlabel metal2 660 -872 660 -872 0 net=5699
rlabel metal2 870 -872 870 -872 0 net=5245
rlabel metal2 149 -874 149 -874 0 net=1422
rlabel metal2 761 -874 761 -874 0 net=5807
rlabel metal2 149 -876 149 -876 0 net=1233
rlabel metal2 828 -876 828 -876 0 net=8011
rlabel metal2 156 -878 156 -878 0 net=3315
rlabel metal2 639 -878 639 -878 0 net=4761
rlabel metal2 975 -878 975 -878 0 net=5489
rlabel metal2 369 -880 369 -880 0 net=2039
rlabel metal2 1010 -880 1010 -880 0 net=5805
rlabel metal2 842 -882 842 -882 0 net=4119
rlabel metal2 842 -884 842 -884 0 net=4949
rlabel metal2 537 -886 537 -886 0 net=3307
rlabel metal2 23 -897 23 -897 0 net=2377
rlabel metal2 23 -897 23 -897 0 net=2377
rlabel metal2 40 -897 40 -897 0 net=1446
rlabel metal2 376 -897 376 -897 0 net=5942
rlabel metal2 1318 -897 1318 -897 0 net=6252
rlabel metal2 1503 -897 1503 -897 0 net=6874
rlabel metal2 44 -899 44 -899 0 net=6138
rlabel metal2 1178 -899 1178 -899 0 net=6947
rlabel metal2 1402 -899 1402 -899 0 net=7951
rlabel metal2 1402 -899 1402 -899 0 net=7951
rlabel metal2 51 -901 51 -901 0 net=2318
rlabel metal2 467 -901 467 -901 0 net=5498
rlabel metal2 1234 -901 1234 -901 0 net=7027
rlabel metal2 51 -903 51 -903 0 net=1855
rlabel metal2 334 -903 334 -903 0 net=1704
rlabel metal2 352 -903 352 -903 0 net=1935
rlabel metal2 387 -903 387 -903 0 net=2040
rlabel metal2 604 -903 604 -903 0 net=3723
rlabel metal2 604 -903 604 -903 0 net=3723
rlabel metal2 646 -903 646 -903 0 net=5866
rlabel metal2 1066 -903 1066 -903 0 net=6513
rlabel metal2 1073 -903 1073 -903 0 net=6369
rlabel metal2 30 -905 30 -905 0 net=2245
rlabel metal2 429 -905 429 -905 0 net=1894
rlabel metal2 443 -905 443 -905 0 net=2329
rlabel metal2 471 -905 471 -905 0 net=2631
rlabel metal2 471 -905 471 -905 0 net=2631
rlabel metal2 485 -905 485 -905 0 net=2675
rlabel metal2 485 -905 485 -905 0 net=2675
rlabel metal2 492 -905 492 -905 0 net=3816
rlabel metal2 656 -905 656 -905 0 net=4072
rlabel metal2 747 -905 747 -905 0 net=5268
rlabel metal2 761 -905 761 -905 0 net=6314
rlabel metal2 30 -907 30 -907 0 net=1623
rlabel metal2 184 -907 184 -907 0 net=1554
rlabel metal2 296 -907 296 -907 0 net=3590
rlabel metal2 1066 -907 1066 -907 0 net=6149
rlabel metal2 1297 -907 1297 -907 0 net=7639
rlabel metal2 16 -909 16 -909 0 net=1521
rlabel metal2 184 -909 184 -909 0 net=1343
rlabel metal2 198 -909 198 -909 0 net=1374
rlabel metal2 436 -909 436 -909 0 net=3027
rlabel metal2 534 -909 534 -909 0 net=3572
rlabel metal2 660 -909 660 -909 0 net=5876
rlabel metal2 1094 -909 1094 -909 0 net=7251
rlabel metal2 1374 -909 1374 -909 0 net=8131
rlabel metal2 58 -911 58 -911 0 net=1123
rlabel metal2 58 -911 58 -911 0 net=1123
rlabel metal2 65 -911 65 -911 0 net=4152
rlabel metal2 681 -911 681 -911 0 net=3789
rlabel metal2 681 -911 681 -911 0 net=3789
rlabel metal2 691 -911 691 -911 0 net=5806
rlabel metal2 1017 -911 1017 -911 0 net=6861
rlabel metal2 1437 -911 1437 -911 0 net=8441
rlabel metal2 65 -913 65 -913 0 net=1533
rlabel metal2 100 -913 100 -913 0 net=3002
rlabel metal2 495 -913 495 -913 0 net=4331
rlabel metal2 705 -913 705 -913 0 net=7330
rlabel metal2 79 -915 79 -915 0 net=4161
rlabel metal2 100 -915 100 -915 0 net=3005
rlabel metal2 212 -915 212 -915 0 net=2437
rlabel metal2 450 -915 450 -915 0 net=4508
rlabel metal2 639 -915 639 -915 0 net=6397
rlabel metal2 16 -917 16 -917 0 net=3821
rlabel metal2 114 -917 114 -917 0 net=1508
rlabel metal2 240 -917 240 -917 0 net=2419
rlabel metal2 499 -917 499 -917 0 net=2717
rlabel metal2 499 -917 499 -917 0 net=2717
rlabel metal2 509 -917 509 -917 0 net=3602
rlabel metal2 709 -917 709 -917 0 net=8046
rlabel metal2 9 -919 9 -919 0 net=4808
rlabel metal2 712 -919 712 -919 0 net=6074
rlabel metal2 9 -921 9 -921 0 net=1977
rlabel metal2 96 -921 96 -921 0 net=3129
rlabel metal2 338 -921 338 -921 0 net=4891
rlabel metal2 639 -921 639 -921 0 net=5227
rlabel metal2 1024 -921 1024 -921 0 net=5983
rlabel metal2 1024 -921 1024 -921 0 net=5983
rlabel metal2 1045 -921 1045 -921 0 net=6301
rlabel metal2 1143 -921 1143 -921 0 net=7215
rlabel metal2 72 -923 72 -923 0 net=3441
rlabel metal2 145 -923 145 -923 0 net=6091
rlabel metal2 1122 -923 1122 -923 0 net=6353
rlabel metal2 1143 -923 1143 -923 0 net=6663
rlabel metal2 1290 -923 1290 -923 0 net=7317
rlabel metal2 114 -925 114 -925 0 net=1379
rlabel metal2 352 -925 352 -925 0 net=1345
rlabel metal2 513 -925 513 -925 0 net=3099
rlabel metal2 534 -925 534 -925 0 net=3865
rlabel metal2 667 -925 667 -925 0 net=3495
rlabel metal2 730 -925 730 -925 0 net=4061
rlabel metal2 807 -925 807 -925 0 net=7928
rlabel metal2 142 -927 142 -927 0 net=8100
rlabel metal2 163 -929 163 -929 0 net=2230
rlabel metal2 310 -929 310 -929 0 net=1571
rlabel metal2 513 -929 513 -929 0 net=3769
rlabel metal2 754 -929 754 -929 0 net=7088
rlabel metal2 1290 -929 1290 -929 0 net=7607
rlabel metal2 1360 -929 1360 -929 0 net=8081
rlabel metal2 37 -931 37 -931 0 net=7089
rlabel metal2 1353 -931 1353 -931 0 net=8013
rlabel metal2 37 -933 37 -933 0 net=3317
rlabel metal2 163 -933 163 -933 0 net=2659
rlabel metal2 520 -933 520 -933 0 net=4079
rlabel metal2 758 -933 758 -933 0 net=7392
rlabel metal2 1416 -933 1416 -933 0 net=8215
rlabel metal2 2 -935 2 -935 0 net=4829
rlabel metal2 537 -935 537 -935 0 net=4046
rlabel metal2 2 -937 2 -937 0 net=3915
rlabel metal2 768 -937 768 -937 0 net=8248
rlabel metal2 131 -939 131 -939 0 net=4269
rlabel metal2 800 -939 800 -939 0 net=5051
rlabel metal2 898 -939 898 -939 0 net=4617
rlabel metal2 898 -939 898 -939 0 net=4617
rlabel metal2 908 -939 908 -939 0 net=7566
rlabel metal2 1444 -939 1444 -939 0 net=8261
rlabel metal2 156 -941 156 -941 0 net=2195
rlabel metal2 807 -941 807 -941 0 net=5003
rlabel metal2 891 -941 891 -941 0 net=5047
rlabel metal2 919 -941 919 -941 0 net=5297
rlabel metal2 919 -941 919 -941 0 net=5297
rlabel metal2 940 -941 940 -941 0 net=5503
rlabel metal2 975 -941 975 -941 0 net=5491
rlabel metal2 989 -941 989 -941 0 net=5789
rlabel metal2 1129 -941 1129 -941 0 net=6453
rlabel metal2 1199 -941 1199 -941 0 net=7003
rlabel metal2 1325 -941 1325 -941 0 net=7705
rlabel metal2 177 -943 177 -943 0 net=1213
rlabel metal2 380 -943 380 -943 0 net=3285
rlabel metal2 478 -943 478 -943 0 net=3578
rlabel metal2 943 -943 943 -943 0 net=6845
rlabel metal2 1248 -943 1248 -943 0 net=7149
rlabel metal2 1332 -943 1332 -943 0 net=7819
rlabel metal2 128 -945 128 -945 0 net=1001
rlabel metal2 191 -945 191 -945 0 net=1511
rlabel metal2 275 -945 275 -945 0 net=1997
rlabel metal2 415 -945 415 -945 0 net=6593
rlabel metal2 1283 -945 1283 -945 0 net=7431
rlabel metal2 1381 -945 1381 -945 0 net=8157
rlabel metal2 121 -947 121 -947 0 net=1039
rlabel metal2 198 -947 198 -947 0 net=2017
rlabel metal2 254 -947 254 -947 0 net=1285
rlabel metal2 373 -947 373 -947 0 net=2941
rlabel metal2 121 -949 121 -949 0 net=1235
rlabel metal2 205 -949 205 -949 0 net=1085
rlabel metal2 537 -949 537 -949 0 net=6054
rlabel metal2 1185 -949 1185 -949 0 net=6963
rlabel metal2 1388 -949 1388 -949 0 net=8195
rlabel metal2 149 -951 149 -951 0 net=1045
rlabel metal2 824 -951 824 -951 0 net=5574
rlabel metal2 975 -951 975 -951 0 net=5891
rlabel metal2 1010 -951 1010 -951 0 net=3969
rlabel metal2 212 -953 212 -953 0 net=1667
rlabel metal2 541 -953 541 -953 0 net=5808
rlabel metal2 1241 -953 1241 -953 0 net=7111
rlabel metal2 254 -955 254 -955 0 net=1851
rlabel metal2 541 -955 541 -955 0 net=3501
rlabel metal2 576 -955 576 -955 0 net=3707
rlabel metal2 677 -955 677 -955 0 net=7061
rlabel metal2 1269 -955 1269 -955 0 net=7405
rlabel metal2 261 -957 261 -957 0 net=1367
rlabel metal2 303 -957 303 -957 0 net=2073
rlabel metal2 544 -957 544 -957 0 net=3446
rlabel metal2 828 -957 828 -957 0 net=4762
rlabel metal2 926 -957 926 -957 0 net=5311
rlabel metal2 1059 -957 1059 -957 0 net=4121
rlabel metal2 44 -959 44 -959 0 net=3693
rlabel metal2 548 -959 548 -959 0 net=8423
rlabel metal2 289 -961 289 -961 0 net=2181
rlabel metal2 551 -961 551 -961 0 net=7985
rlabel metal2 324 -963 324 -963 0 net=2283
rlabel metal2 394 -963 394 -963 0 net=4109
rlabel metal2 828 -963 828 -963 0 net=8295
rlabel metal2 1311 -963 1311 -963 0 net=7409
rlabel metal2 247 -965 247 -965 0 net=1957
rlabel metal2 401 -965 401 -965 0 net=2141
rlabel metal2 555 -965 555 -965 0 net=3629
rlabel metal2 590 -965 590 -965 0 net=3369
rlabel metal2 831 -965 831 -965 0 net=5852
rlabel metal2 1059 -965 1059 -965 0 net=6143
rlabel metal2 1129 -965 1129 -965 0 net=6637
rlabel metal2 1339 -965 1339 -965 0 net=7871
rlabel metal2 86 -967 86 -967 0 net=4023
rlabel metal2 597 -967 597 -967 0 net=4676
rlabel metal2 838 -967 838 -967 0 net=8294
rlabel metal2 86 -969 86 -969 0 net=1819
rlabel metal2 219 -969 219 -969 0 net=2013
rlabel metal2 723 -969 723 -969 0 net=4437
rlabel metal2 849 -969 849 -969 0 net=3308
rlabel metal2 877 -969 877 -969 0 net=4959
rlabel metal2 933 -969 933 -969 0 net=5455
rlabel metal2 996 -969 996 -969 0 net=8379
rlabel metal2 107 -971 107 -971 0 net=1879
rlabel metal2 219 -971 219 -971 0 net=1177
rlabel metal2 625 -971 625 -971 0 net=5879
rlabel metal2 856 -971 856 -971 0 net=5507
rlabel metal2 968 -971 968 -971 0 net=5951
rlabel metal2 1003 -971 1003 -971 0 net=5839
rlabel metal2 1069 -971 1069 -971 0 net=1
rlabel metal2 1171 -971 1171 -971 0 net=6891
rlabel metal2 135 -973 135 -973 0 net=1021
rlabel metal2 583 -973 583 -973 0 net=3173
rlabel metal2 884 -973 884 -973 0 net=5277
rlabel metal2 947 -973 947 -973 0 net=5619
rlabel metal2 1003 -973 1003 -973 0 net=6167
rlabel metal2 1192 -973 1192 -973 0 net=7621
rlabel metal2 247 -975 247 -975 0 net=2895
rlabel metal2 331 -975 331 -975 0 net=3145
rlabel metal2 611 -975 611 -975 0 net=4759
rlabel metal2 1080 -975 1080 -975 0 net=6381
rlabel metal2 1213 -975 1213 -975 0 net=7035
rlabel metal2 1367 -975 1367 -975 0 net=8269
rlabel metal2 282 -977 282 -977 0 net=3643
rlabel metal2 611 -977 611 -977 0 net=3939
rlabel metal2 716 -977 716 -977 0 net=7337
rlabel metal2 282 -979 282 -979 0 net=3685
rlabel metal2 632 -979 632 -979 0 net=2737
rlabel metal2 863 -979 863 -979 0 net=5701
rlabel metal2 1087 -979 1087 -979 0 net=6487
rlabel metal2 1150 -979 1150 -979 0 net=6769
rlabel metal2 366 -981 366 -981 0 net=5381
rlabel metal2 835 -981 835 -981 0 net=7007
rlabel metal2 268 -983 268 -983 0 net=2693
rlabel metal2 422 -983 422 -983 0 net=3487
rlabel metal2 688 -983 688 -983 0 net=5319
rlabel metal2 1087 -983 1087 -983 0 net=6579
rlabel metal2 268 -985 268 -985 0 net=1355
rlabel metal2 422 -985 422 -985 0 net=4095
rlabel metal2 751 -985 751 -985 0 net=6667
rlabel metal2 317 -987 317 -987 0 net=3231
rlabel metal2 691 -987 691 -987 0 net=3611
rlabel metal2 744 -987 744 -987 0 net=6419
rlabel metal2 569 -989 569 -989 0 net=1493
rlabel metal2 786 -989 786 -989 0 net=4395
rlabel metal2 863 -989 863 -989 0 net=5247
rlabel metal2 653 -991 653 -991 0 net=5631
rlabel metal2 765 -993 765 -993 0 net=4197
rlabel metal2 786 -993 786 -993 0 net=4713
rlabel metal2 548 -995 548 -995 0 net=4533
rlabel metal2 793 -995 793 -995 0 net=4529
rlabel metal2 779 -997 779 -997 0 net=4391
rlabel metal2 779 -999 779 -999 0 net=4951
rlabel metal2 821 -1001 821 -1001 0 net=4567
rlabel metal2 821 -1003 821 -1003 0 net=5961
rlabel metal2 72 -1014 72 -1014 0 net=3442
rlabel metal2 796 -1014 796 -1014 0 net=5790
rlabel metal2 1150 -1014 1150 -1014 0 net=6771
rlabel metal2 1150 -1014 1150 -1014 0 net=6771
rlabel metal2 1164 -1014 1164 -1014 0 net=6847
rlabel metal2 72 -1016 72 -1016 0 net=2381
rlabel metal2 93 -1016 93 -1016 0 net=4760
rlabel metal2 989 -1016 989 -1016 0 net=7028
rlabel metal2 1276 -1016 1276 -1016 0 net=8297
rlabel metal2 93 -1018 93 -1018 0 net=1179
rlabel metal2 226 -1018 226 -1018 0 net=1214
rlabel metal2 310 -1018 310 -1018 0 net=1572
rlabel metal2 541 -1018 541 -1018 0 net=7410
rlabel metal2 1325 -1018 1325 -1018 0 net=7707
rlabel metal2 2 -1020 2 -1020 0 net=3917
rlabel metal2 548 -1020 548 -1020 0 net=4392
rlabel metal2 821 -1020 821 -1020 0 net=7216
rlabel metal2 1423 -1020 1423 -1020 0 net=8262
rlabel metal2 1451 -1020 1451 -1020 0 net=2943
rlabel metal2 2 -1022 2 -1022 0 net=1357
rlabel metal2 310 -1022 310 -1022 0 net=2969
rlabel metal2 908 -1022 908 -1022 0 net=7965
rlabel metal2 44 -1024 44 -1024 0 net=3695
rlabel metal2 240 -1024 240 -1024 0 net=3851
rlabel metal2 254 -1024 254 -1024 0 net=1852
rlabel metal2 705 -1024 705 -1024 0 net=7587
rlabel metal2 23 -1026 23 -1026 0 net=2379
rlabel metal2 96 -1026 96 -1026 0 net=3488
rlabel metal2 590 -1026 590 -1026 0 net=3371
rlabel metal2 691 -1026 691 -1026 0 net=5175
rlabel metal2 992 -1026 992 -1026 0 net=6144
rlabel metal2 1108 -1026 1108 -1026 0 net=6515
rlabel metal2 1255 -1026 1255 -1026 0 net=7253
rlabel metal2 1437 -1026 1437 -1026 0 net=8443
rlabel metal2 23 -1028 23 -1028 0 net=1131
rlabel metal2 107 -1028 107 -1028 0 net=1880
rlabel metal2 170 -1028 170 -1028 0 net=1523
rlabel metal2 170 -1028 170 -1028 0 net=1523
rlabel metal2 184 -1028 184 -1028 0 net=1344
rlabel metal2 345 -1028 345 -1028 0 net=1959
rlabel metal2 345 -1028 345 -1028 0 net=1959
rlabel metal2 376 -1028 376 -1028 0 net=1494
rlabel metal2 576 -1028 576 -1028 0 net=3630
rlabel metal2 600 -1028 600 -1028 0 net=6599
rlabel metal2 1283 -1028 1283 -1028 0 net=7433
rlabel metal2 37 -1030 37 -1030 0 net=3319
rlabel metal2 607 -1030 607 -1030 0 net=6092
rlabel metal2 1143 -1030 1143 -1030 0 net=6665
rlabel metal2 1297 -1030 1297 -1030 0 net=7641
rlabel metal2 37 -1032 37 -1032 0 net=1124
rlabel metal2 107 -1032 107 -1032 0 net=1003
rlabel metal2 184 -1032 184 -1032 0 net=1347
rlabel metal2 390 -1032 390 -1032 0 net=6150
rlabel metal2 1192 -1032 1192 -1032 0 net=7623
rlabel metal2 33 -1034 33 -1034 0 net=2095
rlabel metal2 201 -1034 201 -1034 0 net=3103
rlabel metal2 240 -1034 240 -1034 0 net=2643
rlabel metal2 842 -1034 842 -1034 0 net=4569
rlabel metal2 940 -1034 940 -1034 0 net=5505
rlabel metal2 1192 -1034 1192 -1034 0 net=7037
rlabel metal2 1304 -1034 1304 -1034 0 net=7319
rlabel metal2 58 -1036 58 -1036 0 net=2019
rlabel metal2 247 -1036 247 -1036 0 net=2897
rlabel metal2 593 -1036 593 -1036 0 net=6862
rlabel metal2 1332 -1036 1332 -1036 0 net=7821
rlabel metal2 79 -1038 79 -1038 0 net=4163
rlabel metal2 856 -1038 856 -1038 0 net=5048
rlabel metal2 940 -1038 940 -1038 0 net=5953
rlabel metal2 1052 -1038 1052 -1038 0 net=4123
rlabel metal2 86 -1040 86 -1040 0 net=1820
rlabel metal2 247 -1040 247 -1040 0 net=1287
rlabel metal2 394 -1040 394 -1040 0 net=4110
rlabel metal2 569 -1040 569 -1040 0 net=4271
rlabel metal2 702 -1040 702 -1040 0 net=3497
rlabel metal2 716 -1040 716 -1040 0 net=3612
rlabel metal2 758 -1040 758 -1040 0 net=3793
rlabel metal2 859 -1040 859 -1040 0 net=8216
rlabel metal2 114 -1042 114 -1042 0 net=1381
rlabel metal2 275 -1042 275 -1042 0 net=2749
rlabel metal2 415 -1042 415 -1042 0 net=6595
rlabel metal2 611 -1042 611 -1042 0 net=3940
rlabel metal2 719 -1042 719 -1042 0 net=6905
rlabel metal2 1339 -1042 1339 -1042 0 net=7873
rlabel metal2 114 -1044 114 -1044 0 net=4531
rlabel metal2 331 -1044 331 -1044 0 net=3385
rlabel metal2 733 -1044 733 -1044 0 net=5443
rlabel metal2 1136 -1044 1136 -1044 0 net=6455
rlabel metal2 1290 -1044 1290 -1044 0 net=7609
rlabel metal2 30 -1046 30 -1046 0 net=1625
rlabel metal2 408 -1046 408 -1046 0 net=2143
rlabel metal2 422 -1046 422 -1046 0 net=4097
rlabel metal2 422 -1046 422 -1046 0 net=4097
rlabel metal2 432 -1046 432 -1046 0 net=3708
rlabel metal2 663 -1046 663 -1046 0 net=8361
rlabel metal2 30 -1048 30 -1048 0 net=1107
rlabel metal2 142 -1048 142 -1048 0 net=1087
rlabel metal2 254 -1048 254 -1048 0 net=2739
rlabel metal2 660 -1048 660 -1048 0 net=4530
rlabel metal2 859 -1048 859 -1048 0 net=7367
rlabel metal2 156 -1050 156 -1050 0 net=2197
rlabel metal2 338 -1050 338 -1050 0 net=4893
rlabel metal2 667 -1050 667 -1050 0 net=4081
rlabel metal2 863 -1050 863 -1050 0 net=5249
rlabel metal2 996 -1050 996 -1050 0 net=5985
rlabel metal2 1171 -1050 1171 -1050 0 net=6893
rlabel metal2 1346 -1050 1346 -1050 0 net=7987
rlabel metal2 135 -1052 135 -1052 0 net=1023
rlabel metal2 205 -1052 205 -1052 0 net=2847
rlabel metal2 870 -1052 870 -1052 0 net=7952
rlabel metal2 121 -1054 121 -1054 0 net=1237
rlabel metal2 261 -1054 261 -1054 0 net=1368
rlabel metal2 408 -1054 408 -1054 0 net=3791
rlabel metal2 730 -1054 730 -1054 0 net=4063
rlabel metal2 936 -1054 936 -1054 0 net=6709
rlabel metal2 1311 -1054 1311 -1054 0 net=8425
rlabel metal2 121 -1056 121 -1056 0 net=1513
rlabel metal2 212 -1056 212 -1056 0 net=1669
rlabel metal2 338 -1056 338 -1056 0 net=1983
rlabel metal2 485 -1056 485 -1056 0 net=2677
rlabel metal2 562 -1056 562 -1056 0 net=3503
rlabel metal2 747 -1056 747 -1056 0 net=5004
rlabel metal2 954 -1056 954 -1056 0 net=5509
rlabel metal2 1178 -1056 1178 -1056 0 net=6949
rlabel metal2 1353 -1056 1353 -1056 0 net=8015
rlabel metal2 9 -1058 9 -1058 0 net=1979
rlabel metal2 359 -1058 359 -1058 0 net=1937
rlabel metal2 394 -1058 394 -1058 0 net=2121
rlabel metal2 793 -1058 793 -1058 0 net=7165
rlabel metal2 145 -1060 145 -1060 0 net=1067
rlabel metal2 359 -1060 359 -1060 0 net=1999
rlabel metal2 446 -1060 446 -1060 0 net=5341
rlabel metal2 1045 -1060 1045 -1060 0 net=6303
rlabel metal2 1185 -1060 1185 -1060 0 net=6965
rlabel metal2 1367 -1060 1367 -1060 0 net=8271
rlabel metal2 163 -1062 163 -1062 0 net=2661
rlabel metal2 460 -1062 460 -1062 0 net=6651
rlabel metal2 1374 -1062 1374 -1062 0 net=8133
rlabel metal2 166 -1064 166 -1064 0 net=6355
rlabel metal2 1199 -1064 1199 -1064 0 net=7005
rlabel metal2 1381 -1064 1381 -1064 0 net=8159
rlabel metal2 464 -1066 464 -1066 0 net=2331
rlabel metal2 933 -1066 933 -1066 0 net=5457
rlabel metal2 1073 -1066 1073 -1066 0 net=6371
rlabel metal2 1220 -1066 1220 -1066 0 net=7063
rlabel metal2 1388 -1066 1388 -1066 0 net=8197
rlabel metal2 9 -1068 9 -1068 0 net=6467
rlabel metal2 1227 -1068 1227 -1068 0 net=7091
rlabel metal2 1395 -1068 1395 -1068 0 net=8381
rlabel metal2 243 -1070 243 -1070 0 net=1991
rlabel metal2 478 -1070 478 -1070 0 net=4830
rlabel metal2 534 -1070 534 -1070 0 net=7267
rlabel metal2 429 -1072 429 -1072 0 net=2439
rlabel metal2 485 -1072 485 -1072 0 net=2485
rlabel metal2 933 -1072 933 -1072 0 net=7406
rlabel metal2 492 -1074 492 -1074 0 net=6971
rlabel metal2 355 -1076 355 -1076 0 net=2505
rlabel metal2 495 -1076 495 -1076 0 net=4311
rlabel metal2 947 -1076 947 -1076 0 net=5621
rlabel metal2 1080 -1076 1080 -1076 0 net=6383
rlabel metal2 499 -1078 499 -1078 0 net=2719
rlabel metal2 544 -1078 544 -1078 0 net=3321
rlabel metal2 828 -1078 828 -1078 0 net=6055
rlabel metal2 1241 -1078 1241 -1078 0 net=7113
rlabel metal2 471 -1080 471 -1080 0 net=2633
rlabel metal2 555 -1080 555 -1080 0 net=4025
rlabel metal2 877 -1080 877 -1080 0 net=4961
rlabel metal2 954 -1080 954 -1080 0 net=7779
rlabel metal2 443 -1082 443 -1082 0 net=2421
rlabel metal2 555 -1082 555 -1082 0 net=1403
rlabel metal2 957 -1082 957 -1082 0 net=6668
rlabel metal2 1248 -1082 1248 -1082 0 net=7151
rlabel metal2 443 -1084 443 -1084 0 net=6063
rlabel metal2 1248 -1084 1248 -1084 0 net=8083
rlabel metal2 562 -1086 562 -1086 0 net=2767
rlabel metal2 835 -1086 835 -1086 0 net=4397
rlabel metal2 975 -1086 975 -1086 0 net=5893
rlabel metal2 1115 -1086 1115 -1086 0 net=6489
rlabel metal2 1262 -1086 1262 -1086 0 net=7339
rlabel metal2 79 -1088 79 -1088 0 net=6617
rlabel metal2 611 -1090 611 -1090 0 net=4535
rlabel metal2 779 -1090 779 -1090 0 net=4953
rlabel metal2 1129 -1090 1129 -1090 0 net=6639
rlabel metal2 831 -1092 831 -1092 0 net=6793
rlabel metal2 628 -1094 628 -1094 0 net=6163
rlabel metal2 653 -1096 653 -1096 0 net=5633
rlabel metal2 1087 -1096 1087 -1096 0 net=6581
rlabel metal2 604 -1098 604 -1098 0 net=3725
rlabel metal2 670 -1098 670 -1098 0 net=6281
rlabel metal2 1206 -1098 1206 -1098 0 net=7009
rlabel metal2 674 -1100 674 -1100 0 net=7611
rlabel metal2 674 -1102 674 -1102 0 net=2983
rlabel metal2 751 -1102 751 -1102 0 net=4981
rlabel metal2 835 -1102 835 -1102 0 net=5493
rlabel metal2 1003 -1102 1003 -1102 0 net=6169
rlabel metal2 513 -1104 513 -1104 0 net=3771
rlabel metal2 751 -1104 751 -1104 0 net=6354
rlabel metal2 401 -1106 401 -1106 0 net=2015
rlabel metal2 639 -1106 639 -1106 0 net=5229
rlabel metal2 1003 -1106 1003 -1106 0 net=5963
rlabel metal2 1094 -1106 1094 -1106 0 net=6399
rlabel metal2 401 -1108 401 -1108 0 net=3287
rlabel metal2 457 -1108 457 -1108 0 net=3147
rlabel metal2 884 -1108 884 -1108 0 net=5279
rlabel metal2 450 -1110 450 -1110 0 net=4333
rlabel metal2 737 -1110 737 -1110 0 net=4439
rlabel metal2 912 -1110 912 -1110 0 net=5321
rlabel metal2 1031 -1110 1031 -1110 0 net=5841
rlabel metal2 1101 -1110 1101 -1110 0 net=6421
rlabel metal2 457 -1112 457 -1112 0 net=2741
rlabel metal2 604 -1112 604 -1112 0 net=4605
rlabel metal2 919 -1112 919 -1112 0 net=5299
rlabel metal2 625 -1114 625 -1114 0 net=3175
rlabel metal2 723 -1114 723 -1114 0 net=5383
rlabel metal2 282 -1116 282 -1116 0 net=3687
rlabel metal2 737 -1116 737 -1116 0 net=3225
rlabel metal2 849 -1116 849 -1116 0 net=5881
rlabel metal2 282 -1118 282 -1118 0 net=1471
rlabel metal2 849 -1118 849 -1118 0 net=3971
rlabel metal2 317 -1120 317 -1120 0 net=3232
rlabel metal2 898 -1120 898 -1120 0 net=4619
rlabel metal2 926 -1120 926 -1120 0 net=5313
rlabel metal2 100 -1122 100 -1122 0 net=3007
rlabel metal2 436 -1122 436 -1122 0 net=3029
rlabel metal2 961 -1122 961 -1122 0 net=5703
rlabel metal2 100 -1124 100 -1124 0 net=2075
rlabel metal2 387 -1124 387 -1124 0 net=2247
rlabel metal2 786 -1124 786 -1124 0 net=4715
rlabel metal2 975 -1124 975 -1124 0 net=5223
rlabel metal2 65 -1126 65 -1126 0 net=1535
rlabel metal2 667 -1126 667 -1126 0 net=3883
rlabel metal2 800 -1126 800 -1126 0 net=5053
rlabel metal2 51 -1128 51 -1128 0 net=1857
rlabel metal2 765 -1128 765 -1128 0 net=4199
rlabel metal2 16 -1130 16 -1130 0 net=3823
rlabel metal2 16 -1132 16 -1132 0 net=2183
rlabel metal2 51 -1134 51 -1134 0 net=3645
rlabel metal2 233 -1136 233 -1136 0 net=3131
rlabel metal2 506 -1136 506 -1136 0 net=3295
rlabel metal2 149 -1138 149 -1138 0 net=1047
rlabel metal2 128 -1140 128 -1140 0 net=1041
rlabel metal2 128 -1142 128 -1142 0 net=3867
rlabel metal2 527 -1144 527 -1144 0 net=3101
rlabel metal2 366 -1146 366 -1146 0 net=2695
rlabel metal2 324 -1148 324 -1148 0 net=2285
rlabel metal2 324 -1150 324 -1150 0 net=1821
rlabel metal2 9 -1161 9 -1161 0 net=1536
rlabel metal2 341 -1161 341 -1161 0 net=1960
rlabel metal2 352 -1161 352 -1161 0 net=378
rlabel metal2 670 -1161 670 -1161 0 net=4200
rlabel metal2 828 -1161 828 -1161 0 net=5300
rlabel metal2 1248 -1161 1248 -1161 0 net=8085
rlabel metal2 9 -1163 9 -1163 0 net=3783
rlabel metal2 667 -1163 667 -1163 0 net=3853
rlabel metal2 782 -1163 782 -1163 0 net=4026
rlabel metal2 828 -1163 828 -1163 0 net=4313
rlabel metal2 894 -1163 894 -1163 0 net=6384
rlabel metal2 12 -1165 12 -1165 0 net=2380
rlabel metal2 61 -1165 61 -1165 0 net=3320
rlabel metal2 674 -1165 674 -1165 0 net=2985
rlabel metal2 674 -1165 674 -1165 0 net=2985
rlabel metal2 719 -1165 719 -1165 0 net=5280
rlabel metal2 1248 -1165 1248 -1165 0 net=7589
rlabel metal2 23 -1167 23 -1167 0 net=1133
rlabel metal2 23 -1167 23 -1167 0 net=1133
rlabel metal2 30 -1167 30 -1167 0 net=3499
rlabel metal2 719 -1167 719 -1167 0 net=7610
rlabel metal2 33 -1169 33 -1169 0 net=3132
rlabel metal2 310 -1169 310 -1169 0 net=2971
rlabel metal2 408 -1169 408 -1169 0 net=3792
rlabel metal2 957 -1169 957 -1169 0 net=8016
rlabel metal2 37 -1171 37 -1171 0 net=3688
rlabel metal2 730 -1171 730 -1171 0 net=7624
rlabel metal2 1528 -1171 1528 -1171 0 net=8273
rlabel metal2 37 -1173 37 -1173 0 net=3795
rlabel metal2 772 -1173 772 -1173 0 net=4027
rlabel metal2 954 -1173 954 -1173 0 net=5231
rlabel metal2 989 -1173 989 -1173 0 net=5251
rlabel metal2 1055 -1173 1055 -1173 0 net=5551
rlabel metal2 40 -1175 40 -1175 0 net=6596
rlabel metal2 597 -1175 597 -1175 0 net=3149
rlabel metal2 702 -1175 702 -1175 0 net=6641
rlabel metal2 1367 -1175 1367 -1175 0 net=7167
rlabel metal2 1451 -1175 1451 -1175 0 net=7823
rlabel metal2 44 -1177 44 -1177 0 net=1181
rlabel metal2 103 -1177 103 -1177 0 net=4098
rlabel metal2 457 -1177 457 -1177 0 net=3102
rlabel metal2 625 -1177 625 -1177 0 net=5339
rlabel metal2 989 -1177 989 -1177 0 net=5385
rlabel metal2 1122 -1177 1122 -1177 0 net=6065
rlabel metal2 1171 -1177 1171 -1177 0 net=6305
rlabel metal2 51 -1179 51 -1179 0 net=3647
rlabel metal2 481 -1179 481 -1179 0 net=6164
rlabel metal2 1381 -1179 1381 -1179 0 net=7093
rlabel metal2 51 -1181 51 -1181 0 net=2097
rlabel metal2 184 -1181 184 -1181 0 net=1348
rlabel metal2 754 -1181 754 -1181 0 net=5506
rlabel metal2 1143 -1181 1143 -1181 0 net=6283
rlabel metal2 1251 -1181 1251 -1181 0 net=1
rlabel metal2 72 -1183 72 -1183 0 net=2383
rlabel metal2 72 -1183 72 -1183 0 net=2383
rlabel metal2 79 -1183 79 -1183 0 net=2076
rlabel metal2 107 -1183 107 -1183 0 net=1004
rlabel metal2 618 -1183 618 -1183 0 net=3347
rlabel metal2 758 -1183 758 -1183 0 net=4083
rlabel metal2 831 -1183 831 -1183 0 net=5894
rlabel metal2 1164 -1183 1164 -1183 0 net=6423
rlabel metal2 1297 -1183 1297 -1183 0 net=6907
rlabel metal2 1381 -1183 1381 -1183 0 net=7369
rlabel metal2 79 -1185 79 -1185 0 net=3337
rlabel metal2 408 -1185 408 -1185 0 net=2487
rlabel metal2 506 -1185 506 -1185 0 net=3296
rlabel metal2 863 -1185 863 -1185 0 net=4399
rlabel metal2 922 -1185 922 -1185 0 net=7064
rlabel metal2 1402 -1185 1402 -1185 0 net=7321
rlabel metal2 82 -1187 82 -1187 0 net=1992
rlabel metal2 485 -1187 485 -1187 0 net=2769
rlabel metal2 569 -1187 569 -1187 0 net=4273
rlabel metal2 835 -1187 835 -1187 0 net=5494
rlabel metal2 996 -1187 996 -1187 0 net=5987
rlabel metal2 1192 -1187 1192 -1187 0 net=7039
rlabel metal2 1374 -1187 1374 -1187 0 net=7341
rlabel metal2 86 -1189 86 -1189 0 net=1109
rlabel metal2 114 -1189 114 -1189 0 net=4532
rlabel metal2 509 -1189 509 -1189 0 net=2332
rlabel metal2 877 -1189 877 -1189 0 net=4571
rlabel metal2 1059 -1189 1059 -1189 0 net=6057
rlabel metal2 1192 -1189 1192 -1189 0 net=7115
rlabel metal2 1430 -1189 1430 -1189 0 net=7643
rlabel metal2 86 -1191 86 -1191 0 net=3529
rlabel metal2 205 -1191 205 -1191 0 net=2849
rlabel metal2 310 -1191 310 -1191 0 net=1737
rlabel metal2 723 -1191 723 -1191 0 net=5322
rlabel metal2 1136 -1191 1136 -1191 0 net=6171
rlabel metal2 1206 -1191 1206 -1191 0 net=6491
rlabel metal2 1262 -1191 1262 -1191 0 net=6619
rlabel metal2 1479 -1191 1479 -1191 0 net=8161
rlabel metal2 93 -1193 93 -1193 0 net=1915
rlabel metal2 730 -1193 730 -1193 0 net=5635
rlabel metal2 1157 -1193 1157 -1193 0 net=7889
rlabel metal2 1227 -1193 1227 -1193 0 net=6601
rlabel metal2 1262 -1193 1262 -1193 0 net=7709
rlabel metal2 100 -1195 100 -1195 0 net=5407
rlabel metal2 1080 -1195 1080 -1195 0 net=5843
rlabel metal2 1255 -1195 1255 -1195 0 net=8427
rlabel metal2 1360 -1195 1360 -1195 0 net=7011
rlabel metal2 114 -1197 114 -1197 0 net=2441
rlabel metal2 513 -1197 513 -1197 0 net=2016
rlabel metal2 611 -1197 611 -1197 0 net=4537
rlabel metal2 905 -1197 905 -1197 0 net=4621
rlabel metal2 940 -1197 940 -1197 0 net=5955
rlabel metal2 1311 -1197 1311 -1197 0 net=6951
rlabel metal2 1360 -1197 1360 -1197 0 net=7153
rlabel metal2 2 -1199 2 -1199 0 net=1358
rlabel metal2 541 -1199 541 -1199 0 net=3919
rlabel metal2 639 -1199 639 -1199 0 net=3177
rlabel metal2 653 -1199 653 -1199 0 net=3727
rlabel metal2 2 -1201 2 -1201 0 net=5225
rlabel metal2 1003 -1201 1003 -1201 0 net=5965
rlabel metal2 1220 -1201 1220 -1201 0 net=6469
rlabel metal2 1388 -1201 1388 -1201 0 net=8135
rlabel metal2 121 -1203 121 -1203 0 net=1514
rlabel metal2 541 -1203 541 -1203 0 net=1405
rlabel metal2 583 -1203 583 -1203 0 net=3825
rlabel metal2 786 -1203 786 -1203 0 net=3885
rlabel metal2 856 -1203 856 -1203 0 net=7874
rlabel metal2 1542 -1203 1542 -1203 0 net=8445
rlabel metal2 121 -1205 121 -1205 0 net=1383
rlabel metal2 282 -1205 282 -1205 0 net=1473
rlabel metal2 282 -1205 282 -1205 0 net=1473
rlabel metal2 289 -1205 289 -1205 0 net=1985
rlabel metal2 366 -1205 366 -1205 0 net=2287
rlabel metal2 394 -1205 394 -1205 0 net=2122
rlabel metal2 751 -1205 751 -1205 0 net=5675
rlabel metal2 1395 -1205 1395 -1205 0 net=7435
rlabel metal2 1507 -1205 1507 -1205 0 net=8299
rlabel metal2 131 -1207 131 -1207 0 net=106
rlabel metal2 936 -1207 936 -1207 0 net=6557
rlabel metal2 1276 -1207 1276 -1207 0 net=6653
rlabel metal2 166 -1209 166 -1209 0 net=3030
rlabel metal2 940 -1209 940 -1209 0 net=5055
rlabel metal2 975 -1209 975 -1209 0 net=5623
rlabel metal2 1150 -1209 1150 -1209 0 net=6773
rlabel metal2 177 -1211 177 -1211 0 net=1289
rlabel metal2 254 -1211 254 -1211 0 net=2740
rlabel metal2 961 -1211 961 -1211 0 net=5459
rlabel metal2 1150 -1211 1150 -1211 0 net=6357
rlabel metal2 16 -1213 16 -1213 0 net=2185
rlabel metal2 261 -1213 261 -1213 0 net=1671
rlabel metal2 362 -1213 362 -1213 0 net=5639
rlabel metal2 1178 -1213 1178 -1213 0 net=6895
rlabel metal2 16 -1215 16 -1215 0 net=2751
rlabel metal2 366 -1215 366 -1215 0 net=1939
rlabel metal2 394 -1215 394 -1215 0 net=2145
rlabel metal2 422 -1215 422 -1215 0 net=2389
rlabel metal2 520 -1215 520 -1215 0 net=2743
rlabel metal2 653 -1215 653 -1215 0 net=3227
rlabel metal2 765 -1215 765 -1215 0 net=4954
rlabel metal2 1318 -1215 1318 -1215 0 net=6973
rlabel metal2 65 -1217 65 -1217 0 net=1859
rlabel metal2 275 -1217 275 -1217 0 net=1463
rlabel metal2 436 -1217 436 -1217 0 net=2249
rlabel metal2 520 -1217 520 -1217 0 net=2944
rlabel metal2 65 -1219 65 -1219 0 net=2697
rlabel metal2 548 -1219 548 -1219 0 net=2679
rlabel metal2 590 -1219 590 -1219 0 net=6429
rlabel metal2 1535 -1219 1535 -1219 0 net=8383
rlabel metal2 170 -1221 170 -1221 0 net=1525
rlabel metal2 317 -1221 317 -1221 0 net=3009
rlabel metal2 527 -1221 527 -1221 0 net=6749
rlabel metal2 170 -1223 170 -1223 0 net=3817
rlabel metal2 373 -1223 373 -1223 0 net=2635
rlabel metal2 548 -1223 548 -1223 0 net=3183
rlabel metal2 628 -1223 628 -1223 0 net=5427
rlabel metal2 184 -1225 184 -1225 0 net=2621
rlabel metal2 590 -1225 590 -1225 0 net=3323
rlabel metal2 744 -1225 744 -1225 0 net=3773
rlabel metal2 191 -1227 191 -1227 0 net=1069
rlabel metal2 212 -1227 212 -1227 0 net=1980
rlabel metal2 555 -1227 555 -1227 0 net=6848
rlabel metal2 191 -1229 191 -1229 0 net=1049
rlabel metal2 240 -1229 240 -1229 0 net=2645
rlabel metal2 429 -1229 429 -1229 0 net=2423
rlabel metal2 604 -1229 604 -1229 0 net=6666
rlabel metal2 58 -1231 58 -1231 0 net=2021
rlabel metal2 338 -1231 338 -1231 0 net=4047
rlabel metal2 786 -1231 786 -1231 0 net=4165
rlabel metal2 859 -1231 859 -1231 0 net=7006
rlabel metal2 149 -1233 149 -1233 0 net=1043
rlabel metal2 380 -1233 380 -1233 0 net=2663
rlabel metal2 681 -1233 681 -1233 0 net=3373
rlabel metal2 796 -1233 796 -1233 0 net=5314
rlabel metal2 1199 -1233 1199 -1233 0 net=6401
rlabel metal2 1353 -1233 1353 -1233 0 net=7781
rlabel metal2 128 -1235 128 -1235 0 net=3869
rlabel metal2 768 -1235 768 -1235 0 net=6979
rlabel metal2 1409 -1235 1409 -1235 0 net=7255
rlabel metal2 149 -1237 149 -1237 0 net=1779
rlabel metal2 800 -1237 800 -1237 0 net=3973
rlabel metal2 898 -1237 898 -1237 0 net=4963
rlabel metal2 1010 -1237 1010 -1237 0 net=5511
rlabel metal2 1409 -1237 1409 -1237 0 net=7269
rlabel metal2 198 -1239 198 -1239 0 net=4235
rlabel metal2 401 -1239 401 -1239 0 net=3289
rlabel metal2 660 -1239 660 -1239 0 net=3241
rlabel metal2 814 -1239 814 -1239 0 net=4064
rlabel metal2 947 -1239 947 -1239 0 net=5177
rlabel metal2 1066 -1239 1066 -1239 0 net=5705
rlabel metal2 1416 -1239 1416 -1239 0 net=7613
rlabel metal2 212 -1241 212 -1241 0 net=2001
rlabel metal2 401 -1241 401 -1241 0 net=2899
rlabel metal2 632 -1241 632 -1241 0 net=4895
rlabel metal2 838 -1241 838 -1241 0 net=5791
rlabel metal2 1087 -1241 1087 -1241 0 net=5883
rlabel metal2 1465 -1241 1465 -1241 0 net=7967
rlabel metal2 219 -1243 219 -1243 0 net=3105
rlabel metal2 576 -1243 576 -1243 0 net=4717
rlabel metal2 968 -1243 968 -1243 0 net=5343
rlabel metal2 1514 -1243 1514 -1243 0 net=8363
rlabel metal2 142 -1245 142 -1245 0 net=1089
rlabel metal2 226 -1245 226 -1245 0 net=3696
rlabel metal2 450 -1245 450 -1245 0 net=4335
rlabel metal2 849 -1245 849 -1245 0 net=4441
rlabel metal2 912 -1245 912 -1245 0 net=4607
rlabel metal2 58 -1247 58 -1247 0 net=4651
rlabel metal2 926 -1247 926 -1247 0 net=4125
rlabel metal2 128 -1249 128 -1249 0 net=1055
rlabel metal2 226 -1249 226 -1249 0 net=1823
rlabel metal2 450 -1249 450 -1249 0 net=2721
rlabel metal2 632 -1249 632 -1249 0 net=3387
rlabel metal2 737 -1249 737 -1249 0 net=3015
rlabel metal2 296 -1251 296 -1251 0 net=2199
rlabel metal2 471 -1251 471 -1251 0 net=3505
rlabel metal2 779 -1251 779 -1251 0 net=4983
rlabel metal2 1024 -1251 1024 -1251 0 net=5445
rlabel metal2 163 -1253 163 -1253 0 net=6011
rlabel metal2 779 -1253 779 -1253 0 net=7715
rlabel metal2 156 -1255 156 -1255 0 net=1025
rlabel metal2 296 -1255 296 -1255 0 net=2507
rlabel metal2 534 -1255 534 -1255 0 net=1103
rlabel metal2 1038 -1255 1038 -1255 0 net=6373
rlabel metal2 135 -1257 135 -1257 0 net=1239
rlabel metal2 173 -1257 173 -1257 0 net=4033
rlabel metal2 1185 -1257 1185 -1257 0 net=6457
rlabel metal2 135 -1259 135 -1259 0 net=7131
rlabel metal2 492 -1259 492 -1259 0 net=2581
rlabel metal2 1213 -1259 1213 -1259 0 net=6517
rlabel metal2 320 -1261 320 -1261 0 net=3983
rlabel metal2 1234 -1261 1234 -1261 0 net=6583
rlabel metal2 324 -1263 324 -1263 0 net=1627
rlabel metal2 1241 -1263 1241 -1263 0 net=6711
rlabel metal2 331 -1265 331 -1265 0 net=4099
rlabel metal2 1290 -1265 1290 -1265 0 net=6795
rlabel metal2 443 -1267 443 -1267 0 net=2457
rlabel metal2 1304 -1267 1304 -1267 0 net=6967
rlabel metal2 1339 -1269 1339 -1269 0 net=7989
rlabel metal2 1521 -1271 1521 -1271 0 net=8199
rlabel metal2 891 -1273 891 -1273 0 net=2857
rlabel metal2 355 -1275 355 -1275 0 net=4593
rlabel metal2 2 -1286 2 -1286 0 net=5226
rlabel metal2 562 -1286 562 -1286 0 net=2680
rlabel metal2 649 -1286 649 -1286 0 net=7012
rlabel metal2 2 -1288 2 -1288 0 net=2637
rlabel metal2 478 -1288 478 -1288 0 net=6796
rlabel metal2 1409 -1288 1409 -1288 0 net=7271
rlabel metal2 1409 -1288 1409 -1288 0 net=7271
rlabel metal2 1451 -1288 1451 -1288 0 net=7825
rlabel metal2 1486 -1288 1486 -1288 0 net=8365
rlabel metal2 23 -1290 23 -1290 0 net=1135
rlabel metal2 23 -1290 23 -1290 0 net=1135
rlabel metal2 30 -1290 30 -1290 0 net=3500
rlabel metal2 765 -1290 765 -1290 0 net=6430
rlabel metal2 1451 -1290 1451 -1290 0 net=7969
rlabel metal2 1514 -1290 1514 -1290 0 net=8447
rlabel metal2 30 -1292 30 -1292 0 net=1183
rlabel metal2 61 -1292 61 -1292 0 net=6306
rlabel metal2 37 -1294 37 -1294 0 net=3796
rlabel metal2 527 -1294 527 -1294 0 net=1406
rlabel metal2 548 -1294 548 -1294 0 net=3728
rlabel metal2 37 -1296 37 -1296 0 net=2459
rlabel metal2 488 -1296 488 -1296 0 net=2664
rlabel metal2 509 -1296 509 -1296 0 net=5340
rlabel metal2 1052 -1296 1052 -1296 0 net=7094
rlabel metal2 1472 -1296 1472 -1296 0 net=8163
rlabel metal2 44 -1298 44 -1298 0 net=2023
rlabel metal2 268 -1298 268 -1298 0 net=1673
rlabel metal2 268 -1298 268 -1298 0 net=1673
rlabel metal2 282 -1298 282 -1298 0 net=1475
rlabel metal2 282 -1298 282 -1298 0 net=1475
rlabel metal2 338 -1298 338 -1298 0 net=2489
rlabel metal2 422 -1298 422 -1298 0 net=2391
rlabel metal2 467 -1298 467 -1298 0 net=2593
rlabel metal2 548 -1298 548 -1298 0 net=1749
rlabel metal2 782 -1298 782 -1298 0 net=8200
rlabel metal2 68 -1300 68 -1300 0 net=4896
rlabel metal2 835 -1300 835 -1300 0 net=6584
rlabel metal2 1241 -1300 1241 -1300 0 net=6713
rlabel metal2 1241 -1300 1241 -1300 0 net=6713
rlabel metal2 1346 -1300 1346 -1300 0 net=7169
rlabel metal2 1388 -1300 1388 -1300 0 net=8137
rlabel metal2 1479 -1300 1479 -1300 0 net=8301
rlabel metal2 100 -1302 100 -1302 0 net=2424
rlabel metal2 555 -1302 555 -1302 0 net=2987
rlabel metal2 719 -1302 719 -1302 0 net=136
rlabel metal2 100 -1304 100 -1304 0 net=1781
rlabel metal2 156 -1304 156 -1304 0 net=1241
rlabel metal2 156 -1304 156 -1304 0 net=1241
rlabel metal2 177 -1304 177 -1304 0 net=1290
rlabel metal2 345 -1304 345 -1304 0 net=2973
rlabel metal2 387 -1304 387 -1304 0 net=2289
rlabel metal2 562 -1304 562 -1304 0 net=4167
rlabel metal2 793 -1304 793 -1304 0 net=4034
rlabel metal2 1055 -1304 1055 -1304 0 net=8274
rlabel metal2 79 -1306 79 -1306 0 net=3338
rlabel metal2 401 -1306 401 -1306 0 net=2901
rlabel metal2 674 -1306 674 -1306 0 net=3375
rlabel metal2 723 -1306 723 -1306 0 net=5252
rlabel metal2 1094 -1306 1094 -1306 0 net=5967
rlabel metal2 1094 -1306 1094 -1306 0 net=5967
rlabel metal2 1171 -1306 1171 -1306 0 net=7322
rlabel metal2 1507 -1306 1507 -1306 0 net=8385
rlabel metal2 79 -1308 79 -1308 0 net=4236
rlabel metal2 233 -1308 233 -1308 0 net=1044
rlabel metal2 366 -1308 366 -1308 0 net=1941
rlabel metal2 366 -1308 366 -1308 0 net=1941
rlabel metal2 418 -1308 418 -1308 0 net=7575
rlabel metal2 1388 -1308 1388 -1308 0 net=7645
rlabel metal2 1528 -1308 1528 -1308 0 net=2859
rlabel metal2 82 -1310 82 -1310 0 net=1007
rlabel metal2 191 -1310 191 -1310 0 net=1051
rlabel metal2 191 -1310 191 -1310 0 net=1051
rlabel metal2 198 -1310 198 -1310 0 net=4249
rlabel metal2 632 -1310 632 -1310 0 net=3389
rlabel metal2 723 -1310 723 -1310 0 net=3635
rlabel metal2 772 -1310 772 -1310 0 net=4029
rlabel metal2 772 -1310 772 -1310 0 net=4029
rlabel metal2 779 -1310 779 -1310 0 net=4315
rlabel metal2 835 -1310 835 -1310 0 net=4337
rlabel metal2 880 -1310 880 -1310 0 net=8086
rlabel metal2 86 -1312 86 -1312 0 net=3530
rlabel metal2 345 -1312 345 -1312 0 net=1789
rlabel metal2 422 -1312 422 -1312 0 net=2723
rlabel metal2 481 -1312 481 -1312 0 net=4035
rlabel metal2 828 -1312 828 -1312 0 net=4237
rlabel metal2 922 -1312 922 -1312 0 net=6654
rlabel metal2 86 -1314 86 -1314 0 net=2647
rlabel metal2 450 -1314 450 -1314 0 net=2771
rlabel metal2 604 -1314 604 -1314 0 net=3213
rlabel metal2 933 -1314 933 -1314 0 net=7256
rlabel metal2 9 -1316 9 -1316 0 net=3784
rlabel metal2 737 -1316 737 -1316 0 net=3016
rlabel metal2 933 -1316 933 -1316 0 net=5233
rlabel metal2 975 -1316 975 -1316 0 net=5625
rlabel metal2 1101 -1316 1101 -1316 0 net=4609
rlabel metal2 9 -1318 9 -1318 0 net=2699
rlabel metal2 93 -1318 93 -1318 0 net=1917
rlabel metal2 212 -1318 212 -1318 0 net=2002
rlabel metal2 667 -1318 667 -1318 0 net=3855
rlabel metal2 744 -1318 744 -1318 0 net=4049
rlabel metal2 838 -1318 838 -1318 0 net=4400
rlabel metal2 898 -1318 898 -1318 0 net=4965
rlabel metal2 982 -1318 982 -1318 0 net=5409
rlabel metal2 1024 -1318 1024 -1318 0 net=5447
rlabel metal2 1101 -1318 1101 -1318 0 net=6519
rlabel metal2 1220 -1318 1220 -1318 0 net=6559
rlabel metal2 1220 -1318 1220 -1318 0 net=6559
rlabel metal2 1234 -1318 1234 -1318 0 net=7711
rlabel metal2 1339 -1318 1339 -1318 0 net=7991
rlabel metal2 93 -1320 93 -1320 0 net=3291
rlabel metal2 618 -1320 618 -1320 0 net=3349
rlabel metal2 688 -1320 688 -1320 0 net=3871
rlabel metal2 751 -1320 751 -1320 0 net=6952
rlabel metal2 1353 -1320 1353 -1320 0 net=7783
rlabel metal2 103 -1322 103 -1322 0 net=6620
rlabel metal2 110 -1324 110 -1324 0 net=2508
rlabel metal2 303 -1324 303 -1324 0 net=2851
rlabel metal2 765 -1324 765 -1324 0 net=3975
rlabel metal2 849 -1324 849 -1324 0 net=4443
rlabel metal2 961 -1324 961 -1324 0 net=5461
rlabel metal2 1038 -1324 1038 -1324 0 net=6375
rlabel metal2 1255 -1324 1255 -1324 0 net=8429
rlabel metal2 128 -1326 128 -1326 0 net=203
rlabel metal2 863 -1326 863 -1326 0 net=4127
rlabel metal2 940 -1326 940 -1326 0 net=5057
rlabel metal2 996 -1326 996 -1326 0 net=5429
rlabel metal2 1010 -1326 1010 -1326 0 net=5513
rlabel metal2 1087 -1326 1087 -1326 0 net=5885
rlabel metal2 1395 -1326 1395 -1326 0 net=7437
rlabel metal2 1416 -1326 1416 -1326 0 net=7615
rlabel metal2 107 -1328 107 -1328 0 net=1111
rlabel metal2 131 -1328 131 -1328 0 net=6642
rlabel metal2 712 -1328 712 -1328 0 net=6839
rlabel metal2 1311 -1328 1311 -1328 0 net=7155
rlabel metal2 1395 -1328 1395 -1328 0 net=7717
rlabel metal2 107 -1330 107 -1330 0 net=2442
rlabel metal2 215 -1330 215 -1330 0 net=1599
rlabel metal2 303 -1330 303 -1330 0 net=1629
rlabel metal2 352 -1330 352 -1330 0 net=3819
rlabel metal2 618 -1330 618 -1330 0 net=3179
rlabel metal2 730 -1330 730 -1330 0 net=5637
rlabel metal2 1143 -1330 1143 -1330 0 net=6285
rlabel metal2 1178 -1330 1178 -1330 0 net=6897
rlabel metal2 1332 -1330 1332 -1330 0 net=6471
rlabel metal2 16 -1332 16 -1332 0 net=2753
rlabel metal2 436 -1332 436 -1332 0 net=3011
rlabel metal2 639 -1332 639 -1332 0 net=4985
rlabel metal2 926 -1332 926 -1332 0 net=5387
rlabel metal2 1059 -1332 1059 -1332 0 net=6059
rlabel metal2 1157 -1332 1157 -1332 0 net=7891
rlabel metal2 16 -1334 16 -1334 0 net=1071
rlabel metal2 233 -1334 233 -1334 0 net=1739
rlabel metal2 436 -1334 436 -1334 0 net=2251
rlabel metal2 471 -1334 471 -1334 0 net=3507
rlabel metal2 786 -1334 786 -1334 0 net=4539
rlabel metal2 940 -1334 940 -1334 0 net=4861
rlabel metal2 989 -1334 989 -1334 0 net=6359
rlabel metal2 1164 -1334 1164 -1334 0 net=6425
rlabel metal2 1192 -1334 1192 -1334 0 net=7117
rlabel metal2 1360 -1334 1360 -1334 0 net=7343
rlabel metal2 51 -1336 51 -1336 0 net=2099
rlabel metal2 170 -1336 170 -1336 0 net=3535
rlabel metal2 457 -1336 457 -1336 0 net=3649
rlabel metal2 800 -1336 800 -1336 0 net=3887
rlabel metal2 842 -1336 842 -1336 0 net=4401
rlabel metal2 856 -1336 856 -1336 0 net=4573
rlabel metal2 947 -1336 947 -1336 0 net=5179
rlabel metal2 1122 -1336 1122 -1336 0 net=6067
rlabel metal2 1255 -1336 1255 -1336 0 net=6775
rlabel metal2 1374 -1336 1374 -1336 0 net=7371
rlabel metal2 51 -1338 51 -1338 0 net=1527
rlabel metal2 275 -1338 275 -1338 0 net=1465
rlabel metal2 317 -1338 317 -1338 0 net=6781
rlabel metal2 877 -1338 877 -1338 0 net=4594
rlabel metal2 905 -1338 905 -1338 0 net=4622
rlabel metal2 1003 -1338 1003 -1338 0 net=6111
rlabel metal2 1122 -1338 1122 -1338 0 net=6603
rlabel metal2 1248 -1338 1248 -1338 0 net=7591
rlabel metal2 65 -1340 65 -1340 0 net=4725
rlabel metal2 1080 -1340 1080 -1340 0 net=5845
rlabel metal2 1269 -1340 1269 -1340 0 net=6751
rlabel metal2 142 -1342 142 -1342 0 net=1057
rlabel metal2 184 -1342 184 -1342 0 net=2623
rlabel metal2 317 -1342 317 -1342 0 net=3353
rlabel metal2 695 -1342 695 -1342 0 net=3985
rlabel metal2 58 -1344 58 -1344 0 net=3541
rlabel metal2 884 -1344 884 -1344 0 net=4653
rlabel metal2 1073 -1344 1073 -1344 0 net=5793
rlabel metal2 1129 -1344 1129 -1344 0 net=5677
rlabel metal2 58 -1346 58 -1346 0 net=3921
rlabel metal2 884 -1346 884 -1346 0 net=5345
rlabel metal2 1066 -1346 1066 -1346 0 net=5707
rlabel metal2 1136 -1346 1136 -1346 0 net=6173
rlabel metal2 1227 -1346 1227 -1346 0 net=6975
rlabel metal2 135 -1348 135 -1348 0 net=7133
rlabel metal2 1136 -1348 1136 -1348 0 net=6981
rlabel metal2 1297 -1348 1297 -1348 0 net=6909
rlabel metal2 72 -1350 72 -1350 0 net=2385
rlabel metal2 142 -1350 142 -1350 0 net=1987
rlabel metal2 457 -1350 457 -1350 0 net=2583
rlabel metal2 495 -1350 495 -1350 0 net=547
rlabel metal2 891 -1350 891 -1350 0 net=4317
rlabel metal2 1045 -1350 1045 -1350 0 net=5641
rlabel metal2 1150 -1350 1150 -1350 0 net=6459
rlabel metal2 1199 -1350 1199 -1350 0 net=6493
rlabel metal2 1297 -1350 1297 -1350 0 net=7041
rlabel metal2 72 -1352 72 -1352 0 net=1091
rlabel metal2 226 -1352 226 -1352 0 net=1825
rlabel metal2 478 -1352 478 -1352 0 net=3639
rlabel metal2 1108 -1352 1108 -1352 0 net=5989
rlabel metal2 1304 -1352 1304 -1352 0 net=6969
rlabel metal2 121 -1354 121 -1354 0 net=1385
rlabel metal2 464 -1354 464 -1354 0 net=3150
rlabel metal2 625 -1354 625 -1354 0 net=3243
rlabel metal2 709 -1354 709 -1354 0 net=6013
rlabel metal2 1185 -1354 1185 -1354 0 net=5553
rlabel metal2 121 -1356 121 -1356 0 net=4101
rlabel metal2 492 -1356 492 -1356 0 net=115
rlabel metal2 523 -1356 523 -1356 0 net=5529
rlabel metal2 163 -1358 163 -1358 0 net=1027
rlabel metal2 205 -1358 205 -1358 0 net=2431
rlabel metal2 597 -1358 597 -1358 0 net=3035
rlabel metal2 1017 -1358 1017 -1358 0 net=5957
rlabel metal2 163 -1360 163 -1360 0 net=1595
rlabel metal2 506 -1360 506 -1360 0 net=7757
rlabel metal2 219 -1362 219 -1362 0 net=1105
rlabel metal2 611 -1362 611 -1362 0 net=3185
rlabel metal2 709 -1362 709 -1362 0 net=3774
rlabel metal2 226 -1364 226 -1364 0 net=3275
rlabel metal2 845 -1364 845 -1364 0 net=6039
rlabel metal2 240 -1366 240 -1366 0 net=2201
rlabel metal2 390 -1366 390 -1366 0 net=3979
rlabel metal2 551 -1366 551 -1366 0 net=3741
rlabel metal2 247 -1368 247 -1368 0 net=2187
rlabel metal2 506 -1368 506 -1368 0 net=2781
rlabel metal2 247 -1370 247 -1370 0 net=3827
rlabel metal2 590 -1370 590 -1370 0 net=3325
rlabel metal2 254 -1372 254 -1372 0 net=1861
rlabel metal2 380 -1372 380 -1372 0 net=2147
rlabel metal2 513 -1372 513 -1372 0 net=3107
rlabel metal2 590 -1372 590 -1372 0 net=3121
rlabel metal2 212 -1374 212 -1374 0 net=1319
rlabel metal2 261 -1374 261 -1374 0 net=1709
rlabel metal2 331 -1376 331 -1376 0 net=2791
rlabel metal2 394 -1378 394 -1378 0 net=3229
rlabel metal2 513 -1380 513 -1380 0 net=6402
rlabel metal2 516 -1382 516 -1382 0 net=6849
rlabel metal2 523 -1384 523 -1384 0 net=5061
rlabel metal2 576 -1386 576 -1386 0 net=4719
rlabel metal2 576 -1388 576 -1388 0 net=4275
rlabel metal2 758 -1390 758 -1390 0 net=4085
rlabel metal2 646 -1392 646 -1392 0 net=2745
rlabel metal2 646 -1394 646 -1394 0 net=5149
rlabel metal2 23 -1405 23 -1405 0 net=1137
rlabel metal2 23 -1405 23 -1405 0 net=1137
rlabel metal2 44 -1405 44 -1405 0 net=2024
rlabel metal2 684 -1405 684 -1405 0 net=3640
rlabel metal2 800 -1405 800 -1405 0 net=3888
rlabel metal2 842 -1405 842 -1405 0 net=7118
rlabel metal2 1528 -1405 1528 -1405 0 net=2861
rlabel metal2 1528 -1405 1528 -1405 0 net=2861
rlabel metal2 1535 -1405 1535 -1405 0 net=4611
rlabel metal2 1535 -1405 1535 -1405 0 net=4611
rlabel metal2 44 -1407 44 -1407 0 net=2101
rlabel metal2 121 -1407 121 -1407 0 net=4102
rlabel metal2 471 -1407 471 -1407 0 net=1826
rlabel metal2 520 -1407 520 -1407 0 net=3820
rlabel metal2 646 -1407 646 -1407 0 net=3986
rlabel metal2 1346 -1407 1346 -1407 0 net=7171
rlabel metal2 1346 -1407 1346 -1407 0 net=7171
rlabel metal2 1353 -1407 1353 -1407 0 net=7345
rlabel metal2 51 -1409 51 -1409 0 net=1528
rlabel metal2 478 -1409 478 -1409 0 net=5062
rlabel metal2 1241 -1409 1241 -1409 0 net=6715
rlabel metal2 1241 -1409 1241 -1409 0 net=6715
rlabel metal2 1311 -1409 1311 -1409 0 net=7157
rlabel metal2 51 -1411 51 -1411 0 net=165
rlabel metal2 320 -1411 320 -1411 0 net=2188
rlabel metal2 478 -1411 478 -1411 0 net=6061
rlabel metal2 1192 -1411 1192 -1411 0 net=7043
rlabel metal2 65 -1413 65 -1413 0 net=1600
rlabel metal2 366 -1413 366 -1413 0 net=1942
rlabel metal2 408 -1413 408 -1413 0 net=5471
rlabel metal2 499 -1413 499 -1413 0 net=2595
rlabel metal2 646 -1413 646 -1413 0 net=6041
rlabel metal2 1276 -1413 1276 -1413 0 net=6753
rlabel metal2 65 -1415 65 -1415 0 net=3013
rlabel metal2 712 -1415 712 -1415 0 net=4316
rlabel metal2 800 -1415 800 -1415 0 net=5958
rlabel metal2 82 -1417 82 -1417 0 net=2624
rlabel metal2 296 -1417 296 -1417 0 net=2491
rlabel metal2 390 -1417 390 -1417 0 net=53
rlabel metal2 562 -1417 562 -1417 0 net=4169
rlabel metal2 807 -1417 807 -1417 0 net=6783
rlabel metal2 68 -1419 68 -1419 0 net=1827
rlabel metal2 394 -1419 394 -1419 0 net=3230
rlabel metal2 842 -1419 842 -1419 0 net=4575
rlabel metal2 873 -1419 873 -1419 0 net=7712
rlabel metal2 1262 -1419 1262 -1419 0 net=6841
rlabel metal2 82 -1421 82 -1421 0 net=2405
rlabel metal2 184 -1421 184 -1421 0 net=1028
rlabel metal2 562 -1421 562 -1421 0 net=3187
rlabel metal2 723 -1421 723 -1421 0 net=3636
rlabel metal2 730 -1421 730 -1421 0 net=4339
rlabel metal2 856 -1421 856 -1421 0 net=5990
rlabel metal2 1234 -1421 1234 -1421 0 net=6679
rlabel metal2 93 -1423 93 -1423 0 net=3293
rlabel metal2 513 -1423 513 -1423 0 net=2903
rlabel metal2 569 -1423 569 -1423 0 net=3329
rlabel metal2 1003 -1423 1003 -1423 0 net=5531
rlabel metal2 1076 -1423 1076 -1423 0 net=6910
rlabel metal2 1332 -1423 1332 -1423 0 net=5678
rlabel metal2 37 -1425 37 -1425 0 net=2461
rlabel metal2 100 -1425 100 -1425 0 net=1782
rlabel metal2 464 -1425 464 -1425 0 net=6363
rlabel metal2 1164 -1425 1164 -1425 0 net=6175
rlabel metal2 37 -1427 37 -1427 0 net=1393
rlabel metal2 880 -1427 880 -1427 0 net=5234
rlabel metal2 950 -1427 950 -1427 0 net=7826
rlabel metal2 100 -1429 100 -1429 0 net=1320
rlabel metal2 268 -1429 268 -1429 0 net=1675
rlabel metal2 268 -1429 268 -1429 0 net=1675
rlabel metal2 275 -1429 275 -1429 0 net=3509
rlabel metal2 723 -1429 723 -1429 0 net=6376
rlabel metal2 1444 -1429 1444 -1429 0 net=7893
rlabel metal2 103 -1431 103 -1431 0 net=339
rlabel metal2 436 -1431 436 -1431 0 net=2253
rlabel metal2 481 -1431 481 -1431 0 net=6911
rlabel metal2 1416 -1431 1416 -1431 0 net=7759
rlabel metal2 114 -1433 114 -1433 0 net=1711
rlabel metal2 324 -1433 324 -1433 0 net=3537
rlabel metal2 436 -1433 436 -1433 0 net=3355
rlabel metal2 660 -1433 660 -1433 0 net=3873
rlabel metal2 768 -1433 768 -1433 0 net=4427
rlabel metal2 880 -1433 880 -1433 0 net=6970
rlabel metal2 1381 -1433 1381 -1433 0 net=7593
rlabel metal2 135 -1435 135 -1435 0 net=2387
rlabel metal2 261 -1435 261 -1435 0 net=1863
rlabel metal2 541 -1435 541 -1435 0 net=4403
rlabel metal2 884 -1435 884 -1435 0 net=5347
rlabel metal2 919 -1435 919 -1435 0 net=8386
rlabel metal2 79 -1437 79 -1437 0 net=8311
rlabel metal2 135 -1439 135 -1439 0 net=1689
rlabel metal2 184 -1439 184 -1439 0 net=1053
rlabel metal2 205 -1439 205 -1439 0 net=2433
rlabel metal2 555 -1439 555 -1439 0 net=2989
rlabel metal2 1178 -1439 1178 -1439 0 net=6427
rlabel metal2 1381 -1439 1381 -1439 0 net=7273
rlabel metal2 72 -1441 72 -1441 0 net=1093
rlabel metal2 219 -1441 219 -1441 0 net=1106
rlabel metal2 688 -1441 688 -1441 0 net=3543
rlabel metal2 744 -1441 744 -1441 0 net=4031
rlabel metal2 803 -1441 803 -1441 0 net=5763
rlabel metal2 1080 -1441 1080 -1441 0 net=5795
rlabel metal2 1213 -1441 1213 -1441 0 net=6561
rlabel metal2 1409 -1441 1409 -1441 0 net=8139
rlabel metal2 72 -1443 72 -1443 0 net=4721
rlabel metal2 772 -1443 772 -1443 0 net=4445
rlabel metal2 905 -1443 905 -1443 0 net=4655
rlabel metal2 1129 -1443 1129 -1443 0 net=7135
rlabel metal2 191 -1445 191 -1445 0 net=3109
rlabel metal2 653 -1445 653 -1445 0 net=3377
rlabel metal2 849 -1445 849 -1445 0 net=5515
rlabel metal2 1129 -1445 1129 -1445 0 net=6777
rlabel metal2 219 -1447 219 -1447 0 net=2479
rlabel metal2 583 -1447 583 -1447 0 net=3181
rlabel metal2 859 -1447 859 -1447 0 net=7843
rlabel metal2 233 -1449 233 -1449 0 net=1741
rlabel metal2 324 -1449 324 -1449 0 net=1751
rlabel metal2 884 -1449 884 -1449 0 net=5059
rlabel metal2 975 -1449 975 -1449 0 net=8448
rlabel metal2 177 -1451 177 -1451 0 net=1009
rlabel metal2 240 -1451 240 -1451 0 net=2202
rlabel metal2 978 -1451 978 -1451 0 net=5846
rlabel metal2 1514 -1451 1514 -1451 0 net=3399
rlabel metal2 177 -1453 177 -1453 0 net=3123
rlabel metal2 674 -1453 674 -1453 0 net=6729
rlabel metal2 1437 -1453 1437 -1453 0 net=6472
rlabel metal2 198 -1455 198 -1455 0 net=4251
rlabel metal2 898 -1455 898 -1455 0 net=4967
rlabel metal2 1006 -1455 1006 -1455 0 net=7616
rlabel metal2 16 -1457 16 -1457 0 net=1073
rlabel metal2 226 -1457 226 -1457 0 net=3277
rlabel metal2 905 -1457 905 -1457 0 net=4863
rlabel metal2 947 -1457 947 -1457 0 net=6759
rlabel metal2 1388 -1457 1388 -1457 0 net=7647
rlabel metal2 16 -1459 16 -1459 0 net=1185
rlabel metal2 226 -1459 226 -1459 0 net=1791
rlabel metal2 359 -1459 359 -1459 0 net=2393
rlabel metal2 485 -1459 485 -1459 0 net=3073
rlabel metal2 919 -1459 919 -1459 0 net=5151
rlabel metal2 1017 -1459 1017 -1459 0 net=5638
rlabel metal2 1136 -1459 1136 -1459 0 net=6983
rlabel metal2 1374 -1459 1374 -1459 0 net=7373
rlabel metal2 30 -1461 30 -1461 0 net=2783
rlabel metal2 877 -1461 877 -1461 0 net=5361
rlabel metal2 989 -1461 989 -1461 0 net=6361
rlabel metal2 1150 -1461 1150 -1461 0 net=6461
rlabel metal2 1220 -1461 1220 -1461 0 net=6977
rlabel metal2 107 -1463 107 -1463 0 net=5591
rlabel metal2 758 -1463 758 -1463 0 net=2746
rlabel metal2 926 -1463 926 -1463 0 net=5389
rlabel metal2 989 -1463 989 -1463 0 net=7438
rlabel metal2 107 -1465 107 -1465 0 net=1597
rlabel metal2 240 -1465 240 -1465 0 net=2585
rlabel metal2 488 -1465 488 -1465 0 net=7357
rlabel metal2 128 -1467 128 -1467 0 net=1113
rlabel metal2 247 -1467 247 -1467 0 net=3828
rlabel metal2 933 -1467 933 -1467 0 net=5753
rlabel metal2 1017 -1467 1017 -1467 0 net=5709
rlabel metal2 1087 -1467 1087 -1467 0 net=5969
rlabel metal2 1122 -1467 1122 -1467 0 net=6605
rlabel metal2 128 -1469 128 -1469 0 net=5679
rlabel metal2 940 -1469 940 -1469 0 net=5411
rlabel metal2 1020 -1469 1020 -1469 0 net=7992
rlabel metal2 79 -1471 79 -1471 0 net=4823
rlabel metal2 947 -1471 947 -1471 0 net=5643
rlabel metal2 1094 -1471 1094 -1471 0 net=6015
rlabel metal2 1150 -1471 1150 -1471 0 net=6899
rlabel metal2 1486 -1471 1486 -1471 0 net=8367
rlabel metal2 247 -1473 247 -1473 0 net=1387
rlabel metal2 331 -1473 331 -1473 0 net=2793
rlabel metal2 632 -1473 632 -1473 0 net=4341
rlabel metal2 1283 -1473 1283 -1473 0 net=6851
rlabel metal2 1479 -1473 1479 -1473 0 net=8303
rlabel metal2 282 -1475 282 -1475 0 net=1477
rlabel metal2 331 -1475 331 -1475 0 net=2725
rlabel metal2 443 -1475 443 -1475 0 net=1265
rlabel metal2 695 -1475 695 -1475 0 net=3579
rlabel metal2 1283 -1475 1283 -1475 0 net=8431
rlabel metal2 282 -1477 282 -1477 0 net=1631
rlabel metal2 345 -1477 345 -1477 0 net=5117
rlabel metal2 502 -1477 502 -1477 0 net=5165
rlabel metal2 954 -1477 954 -1477 0 net=5181
rlabel metal2 1024 -1477 1024 -1477 0 net=5463
rlabel metal2 1472 -1477 1472 -1477 0 net=8165
rlabel metal2 303 -1479 303 -1479 0 net=1467
rlabel metal2 352 -1479 352 -1479 0 net=2755
rlabel metal2 709 -1479 709 -1479 0 net=8107
rlabel metal2 9 -1481 9 -1481 0 net=2701
rlabel metal2 387 -1481 387 -1481 0 net=4467
rlabel metal2 450 -1481 450 -1481 0 net=2773
rlabel metal2 716 -1481 716 -1481 0 net=3743
rlabel metal2 1451 -1481 1451 -1481 0 net=7971
rlabel metal2 9 -1483 9 -1483 0 net=3391
rlabel metal2 758 -1483 758 -1483 0 net=3977
rlabel metal2 982 -1483 982 -1483 0 net=5431
rlabel metal2 1010 -1483 1010 -1483 0 net=6113
rlabel metal2 1430 -1483 1430 -1483 0 net=7785
rlabel metal2 54 -1485 54 -1485 0 net=7477
rlabel metal2 765 -1485 765 -1485 0 net=997
rlabel metal2 1024 -1485 1024 -1485 0 net=5627
rlabel metal2 1059 -1485 1059 -1485 0 net=6287
rlabel metal2 1395 -1485 1395 -1485 0 net=7719
rlabel metal2 58 -1487 58 -1487 0 net=3923
rlabel metal2 751 -1487 751 -1487 0 net=2853
rlabel metal2 1367 -1487 1367 -1487 0 net=7577
rlabel metal2 58 -1489 58 -1489 0 net=4051
rlabel metal2 1031 -1489 1031 -1489 0 net=5449
rlabel metal2 212 -1491 212 -1491 0 net=5399
rlabel metal2 471 -1491 471 -1491 0 net=6385
rlabel metal2 149 -1493 149 -1493 0 net=1919
rlabel metal2 310 -1493 310 -1493 0 net=1723
rlabel metal2 751 -1493 751 -1493 0 net=4087
rlabel metal2 1031 -1493 1031 -1493 0 net=6069
rlabel metal2 149 -1495 149 -1495 0 net=1059
rlabel metal2 387 -1495 387 -1495 0 net=2291
rlabel metal2 681 -1495 681 -1495 0 net=6437
rlabel metal2 401 -1497 401 -1497 0 net=6273
rlabel metal2 2 -1499 2 -1499 0 net=2639
rlabel metal2 415 -1499 415 -1499 0 net=7457
rlabel metal2 2 -1501 2 -1501 0 net=1989
rlabel metal2 373 -1501 373 -1501 0 net=2975
rlabel metal2 429 -1501 429 -1501 0 net=4318
rlabel metal2 1038 -1501 1038 -1501 0 net=5555
rlabel metal2 142 -1503 142 -1503 0 net=1243
rlabel metal2 373 -1503 373 -1503 0 net=2149
rlabel metal2 814 -1503 814 -1503 0 net=5886
rlabel metal2 86 -1505 86 -1505 0 net=2649
rlabel metal2 821 -1505 821 -1505 0 net=4129
rlabel metal2 891 -1505 891 -1505 0 net=4727
rlabel metal2 1101 -1505 1101 -1505 0 net=6521
rlabel metal2 86 -1507 86 -1507 0 net=3215
rlabel metal2 639 -1507 639 -1507 0 net=4987
rlabel metal2 1101 -1507 1101 -1507 0 net=6495
rlabel metal2 110 -1509 110 -1509 0 net=7065
rlabel metal2 156 -1511 156 -1511 0 net=4277
rlabel metal2 604 -1511 604 -1511 0 net=3245
rlabel metal2 639 -1511 639 -1511 0 net=3351
rlabel metal2 786 -1511 786 -1511 0 net=4541
rlabel metal2 534 -1513 534 -1513 0 net=3981
rlabel metal2 786 -1513 786 -1513 0 net=4239
rlabel metal2 534 -1515 534 -1515 0 net=3037
rlabel metal2 611 -1515 611 -1515 0 net=3327
rlabel metal2 817 -1515 817 -1515 0 net=6533
rlabel metal2 576 -1517 576 -1517 0 net=430
rlabel metal2 597 -1519 597 -1519 0 net=7735
rlabel metal2 611 -1521 611 -1521 0 net=3651
rlabel metal2 828 -1521 828 -1521 0 net=7051
rlabel metal2 702 -1523 702 -1523 0 net=3857
rlabel metal2 737 -1525 737 -1525 0 net=4037
rlabel metal2 394 -1527 394 -1527 0 net=4255
rlabel metal2 2 -1538 2 -1538 0 net=1990
rlabel metal2 142 -1538 142 -1538 0 net=1244
rlabel metal2 212 -1538 212 -1538 0 net=1920
rlabel metal2 471 -1538 471 -1538 0 net=3982
rlabel metal2 674 -1538 674 -1538 0 net=7136
rlabel metal2 1349 -1538 1349 -1538 0 net=4612
rlabel metal2 2 -1540 2 -1540 0 net=3511
rlabel metal2 303 -1540 303 -1540 0 net=1469
rlabel metal2 303 -1540 303 -1540 0 net=1469
rlabel metal2 345 -1540 345 -1540 0 net=5119
rlabel metal2 859 -1540 859 -1540 0 net=3400
rlabel metal2 9 -1542 9 -1542 0 net=3393
rlabel metal2 16 -1542 16 -1542 0 net=1187
rlabel metal2 16 -1542 16 -1542 0 net=1187
rlabel metal2 23 -1542 23 -1542 0 net=1139
rlabel metal2 23 -1542 23 -1542 0 net=1139
rlabel metal2 30 -1542 30 -1542 0 net=2784
rlabel metal2 474 -1542 474 -1542 0 net=664
rlabel metal2 838 -1542 838 -1542 0 net=6978
rlabel metal2 1325 -1542 1325 -1542 0 net=7579
rlabel metal2 9 -1544 9 -1544 0 net=2775
rlabel metal2 502 -1544 502 -1544 0 net=3328
rlabel metal2 639 -1544 639 -1544 0 net=3352
rlabel metal2 758 -1544 758 -1544 0 net=3978
rlabel metal2 782 -1544 782 -1544 0 net=5516
rlabel metal2 880 -1544 880 -1544 0 net=6522
rlabel metal2 1220 -1544 1220 -1544 0 net=6913
rlabel metal2 30 -1546 30 -1546 0 net=1691
rlabel metal2 142 -1546 142 -1546 0 net=4342
rlabel metal2 639 -1546 639 -1546 0 net=3379
rlabel metal2 667 -1546 667 -1546 0 net=4429
rlabel metal2 849 -1546 849 -1546 0 net=4989
rlabel metal2 947 -1546 947 -1546 0 net=5645
rlabel metal2 992 -1546 992 -1546 0 net=6428
rlabel metal2 44 -1548 44 -1548 0 net=2103
rlabel metal2 366 -1548 366 -1548 0 net=3539
rlabel metal2 653 -1548 653 -1548 0 net=3925
rlabel metal2 765 -1548 765 -1548 0 net=6386
rlabel metal2 1185 -1548 1185 -1548 0 net=6731
rlabel metal2 1297 -1548 1297 -1548 0 net=7359
rlabel metal2 44 -1550 44 -1550 0 net=3653
rlabel metal2 618 -1550 618 -1550 0 net=2795
rlabel metal2 677 -1550 677 -1550 0 net=279
rlabel metal2 51 -1552 51 -1552 0 net=1598
rlabel metal2 128 -1552 128 -1552 0 net=5681
rlabel metal2 397 -1552 397 -1552 0 net=3744
rlabel metal2 51 -1554 51 -1554 0 net=3189
rlabel metal2 579 -1554 579 -1554 0 net=4340
rlabel metal2 765 -1554 765 -1554 0 net=4821
rlabel metal2 996 -1554 996 -1554 0 net=5450
rlabel metal2 1122 -1554 1122 -1554 0 net=8140
rlabel metal2 54 -1556 54 -1556 0 net=4446
rlabel metal2 863 -1556 863 -1556 0 net=5153
rlabel metal2 947 -1556 947 -1556 0 net=5533
rlabel metal2 1010 -1556 1010 -1556 0 net=6115
rlabel metal2 1010 -1556 1010 -1556 0 net=6115
rlabel metal2 1073 -1556 1073 -1556 0 net=8166
rlabel metal2 65 -1558 65 -1558 0 net=3014
rlabel metal2 506 -1558 506 -1558 0 net=5593
rlabel metal2 919 -1558 919 -1558 0 net=5433
rlabel metal2 992 -1558 992 -1558 0 net=6023
rlabel metal2 1115 -1558 1115 -1558 0 net=6365
rlabel metal2 1150 -1558 1150 -1558 0 net=6901
rlabel metal2 1171 -1558 1171 -1558 0 net=6681
rlabel metal2 1374 -1558 1374 -1558 0 net=7787
rlabel metal2 65 -1560 65 -1560 0 net=4723
rlabel metal2 75 -1560 75 -1560 0 net=2434
rlabel metal2 534 -1560 534 -1560 0 net=3039
rlabel metal2 534 -1560 534 -1560 0 net=3039
rlabel metal2 583 -1560 583 -1560 0 net=3182
rlabel metal2 681 -1560 681 -1560 0 net=4656
rlabel metal2 1101 -1560 1101 -1560 0 net=6497
rlabel metal2 1150 -1560 1150 -1560 0 net=6535
rlabel metal2 1234 -1560 1234 -1560 0 net=7595
rlabel metal2 1451 -1560 1451 -1560 0 net=2863
rlabel metal2 58 -1562 58 -1562 0 net=4053
rlabel metal2 583 -1562 583 -1562 0 net=3279
rlabel metal2 600 -1562 600 -1562 0 net=4088
rlabel metal2 800 -1562 800 -1562 0 net=6201
rlabel metal2 1101 -1562 1101 -1562 0 net=6275
rlabel metal2 1192 -1562 1192 -1562 0 net=7045
rlabel metal2 1283 -1562 1283 -1562 0 net=8433
rlabel metal2 58 -1564 58 -1564 0 net=2151
rlabel metal2 394 -1564 394 -1564 0 net=8205
rlabel metal2 72 -1566 72 -1566 0 net=2388
rlabel metal2 373 -1566 373 -1566 0 net=2757
rlabel metal2 478 -1566 478 -1566 0 net=6062
rlabel metal2 982 -1566 982 -1566 0 net=5711
rlabel metal2 1059 -1566 1059 -1566 0 net=6289
rlabel metal2 1192 -1566 1192 -1566 0 net=6785
rlabel metal2 1283 -1566 1283 -1566 0 net=6755
rlabel metal2 1402 -1566 1402 -1566 0 net=8109
rlabel metal2 79 -1568 79 -1568 0 net=1713
rlabel metal2 135 -1568 135 -1568 0 net=1223
rlabel metal2 730 -1568 730 -1568 0 net=4257
rlabel metal2 800 -1568 800 -1568 0 net=4577
rlabel metal2 989 -1568 989 -1568 0 net=5737
rlabel metal2 1024 -1568 1024 -1568 0 net=5629
rlabel metal2 1311 -1568 1311 -1568 0 net=7845
rlabel metal2 82 -1570 82 -1570 0 net=3294
rlabel metal2 506 -1570 506 -1570 0 net=4825
rlabel metal2 898 -1570 898 -1570 0 net=4969
rlabel metal2 1059 -1570 1059 -1570 0 net=5813
rlabel metal2 103 -1572 103 -1572 0 net=1792
rlabel metal2 380 -1572 380 -1572 0 net=2651
rlabel metal2 492 -1572 492 -1572 0 net=2597
rlabel metal2 590 -1572 590 -1572 0 net=3859
rlabel metal2 716 -1572 716 -1572 0 net=4039
rlabel metal2 751 -1572 751 -1572 0 net=6070
rlabel metal2 107 -1574 107 -1574 0 net=1828
rlabel metal2 348 -1574 348 -1574 0 net=5133
rlabel metal2 394 -1574 394 -1574 0 net=3075
rlabel metal2 611 -1574 611 -1574 0 net=3875
rlabel metal2 681 -1574 681 -1574 0 net=3581
rlabel metal2 702 -1574 702 -1574 0 net=4241
rlabel metal2 793 -1574 793 -1574 0 net=5827
rlabel metal2 114 -1576 114 -1576 0 net=1865
rlabel metal2 338 -1576 338 -1576 0 net=2825
rlabel metal2 737 -1576 737 -1576 0 net=6176
rlabel metal2 145 -1578 145 -1578 0 net=4032
rlabel metal2 786 -1578 786 -1578 0 net=5669
rlabel metal2 870 -1578 870 -1578 0 net=5167
rlabel metal2 933 -1578 933 -1578 0 net=5755
rlabel metal2 1262 -1578 1262 -1578 0 net=7067
rlabel metal2 128 -1580 128 -1580 0 net=5465
rlabel metal2 996 -1580 996 -1580 0 net=7191
rlabel metal2 1255 -1580 1255 -1580 0 net=6761
rlabel metal2 149 -1582 149 -1582 0 net=1061
rlabel metal2 149 -1582 149 -1582 0 net=1061
rlabel metal2 156 -1582 156 -1582 0 net=4279
rlabel metal2 646 -1582 646 -1582 0 net=6042
rlabel metal2 898 -1582 898 -1582 0 net=5391
rlabel metal2 999 -1582 999 -1582 0 net=6778
rlabel metal2 156 -1584 156 -1584 0 net=1433
rlabel metal2 408 -1584 408 -1584 0 net=5473
rlabel metal2 814 -1584 814 -1584 0 net=5060
rlabel metal2 975 -1584 975 -1584 0 net=5557
rlabel metal2 1045 -1584 1045 -1584 0 net=5765
rlabel metal2 163 -1586 163 -1586 0 net=1115
rlabel metal2 884 -1586 884 -1586 0 net=5349
rlabel metal2 1038 -1586 1038 -1586 0 net=5971
rlabel metal2 1129 -1586 1129 -1586 0 net=6439
rlabel metal2 163 -1588 163 -1588 0 net=2641
rlabel metal2 429 -1588 429 -1588 0 net=2255
rlabel metal2 474 -1588 474 -1588 0 net=2777
rlabel metal2 555 -1588 555 -1588 0 net=7458
rlabel metal2 170 -1590 170 -1590 0 net=750
rlabel metal2 450 -1590 450 -1590 0 net=5401
rlabel metal2 817 -1590 817 -1590 0 net=7119
rlabel metal2 1045 -1590 1045 -1590 0 net=6017
rlabel metal2 1157 -1590 1157 -1590 0 net=6563
rlabel metal2 1367 -1590 1367 -1590 0 net=7761
rlabel metal2 170 -1592 170 -1592 0 net=1095
rlabel metal2 261 -1592 261 -1592 0 net=1725
rlabel metal2 352 -1592 352 -1592 0 net=2703
rlabel metal2 415 -1592 415 -1592 0 net=2977
rlabel metal2 499 -1592 499 -1592 0 net=5671
rlabel metal2 1094 -1592 1094 -1592 0 net=6843
rlabel metal2 100 -1594 100 -1594 0 net=2193
rlabel metal2 240 -1594 240 -1594 0 net=2587
rlabel metal2 331 -1594 331 -1594 0 net=2727
rlabel metal2 450 -1594 450 -1594 0 net=4707
rlabel metal2 1213 -1594 1213 -1594 0 net=7721
rlabel metal2 100 -1596 100 -1596 0 net=2407
rlabel metal2 177 -1596 177 -1596 0 net=3125
rlabel metal2 499 -1596 499 -1596 0 net=7655
rlabel metal2 93 -1598 93 -1598 0 net=2463
rlabel metal2 177 -1598 177 -1598 0 net=1005
rlabel metal2 621 -1598 621 -1598 0 net=4542
rlabel metal2 1052 -1598 1052 -1598 0 net=2855
rlabel metal2 93 -1600 93 -1600 0 net=2481
rlabel metal2 240 -1600 240 -1600 0 net=2293
rlabel metal2 457 -1600 457 -1600 0 net=2905
rlabel metal2 646 -1600 646 -1600 0 net=6362
rlabel metal2 1153 -1600 1153 -1600 0 net=1
rlabel metal2 1276 -1600 1276 -1600 0 net=7173
rlabel metal2 86 -1602 86 -1602 0 net=3217
rlabel metal2 660 -1602 660 -1602 0 net=3545
rlabel metal2 695 -1602 695 -1602 0 net=4171
rlabel metal2 912 -1602 912 -1602 0 net=5363
rlabel metal2 989 -1602 989 -1602 0 net=12
rlabel metal2 86 -1604 86 -1604 0 net=1633
rlabel metal2 296 -1604 296 -1604 0 net=2493
rlabel metal2 369 -1604 369 -1604 0 net=4215
rlabel metal2 471 -1604 471 -1604 0 net=4111
rlabel metal2 723 -1604 723 -1604 0 net=4131
rlabel metal2 968 -1604 968 -1604 0 net=2991
rlabel metal2 184 -1606 184 -1606 0 net=1054
rlabel metal2 684 -1606 684 -1606 0 net=8312
rlabel metal2 184 -1608 184 -1608 0 net=1011
rlabel metal2 282 -1608 282 -1608 0 net=1479
rlabel metal2 331 -1608 331 -1608 0 net=2571
rlabel metal2 740 -1608 740 -1608 0 net=6253
rlabel metal2 1136 -1608 1136 -1608 0 net=6463
rlabel metal2 191 -1610 191 -1610 0 net=3111
rlabel metal2 744 -1610 744 -1610 0 net=3471
rlabel metal2 1052 -1610 1052 -1610 0 net=7053
rlabel metal2 191 -1612 191 -1612 0 net=2957
rlabel metal2 709 -1612 709 -1612 0 net=7479
rlabel metal2 198 -1614 198 -1614 0 net=1075
rlabel metal2 289 -1614 289 -1614 0 net=2395
rlabel metal2 548 -1614 548 -1614 0 net=4253
rlabel metal2 779 -1614 779 -1614 0 net=5464
rlabel metal2 1164 -1614 1164 -1614 0 net=6607
rlabel metal2 198 -1616 198 -1616 0 net=1677
rlabel metal2 359 -1616 359 -1616 0 net=5469
rlabel metal2 821 -1616 821 -1616 0 net=4925
rlabel metal2 835 -1616 835 -1616 0 net=4729
rlabel metal2 905 -1616 905 -1616 0 net=4865
rlabel metal2 1178 -1616 1178 -1616 0 net=6717
rlabel metal2 219 -1618 219 -1618 0 net=1389
rlabel metal2 541 -1618 541 -1618 0 net=4405
rlabel metal2 828 -1618 828 -1618 0 net=6407
rlabel metal2 1227 -1618 1227 -1618 0 net=7347
rlabel metal2 226 -1620 226 -1620 0 net=2117
rlabel metal2 422 -1620 422 -1620 0 net=4469
rlabel metal2 548 -1620 548 -1620 0 net=3247
rlabel metal2 891 -1620 891 -1620 0 net=5183
rlabel metal2 1241 -1620 1241 -1620 0 net=6985
rlabel metal2 1353 -1620 1353 -1620 0 net=7275
rlabel metal2 233 -1622 233 -1622 0 net=1215
rlabel metal2 569 -1622 569 -1622 0 net=3331
rlabel metal2 905 -1622 905 -1622 0 net=5413
rlabel metal2 954 -1622 954 -1622 0 net=7158
rlabel metal2 1381 -1622 1381 -1622 0 net=7895
rlabel metal2 247 -1624 247 -1624 0 net=1267
rlabel metal2 877 -1624 877 -1624 0 net=4365
rlabel metal2 1304 -1624 1304 -1624 0 net=7375
rlabel metal2 296 -1626 296 -1626 0 net=3531
rlabel metal2 877 -1626 877 -1626 0 net=5796
rlabel metal2 1360 -1626 1360 -1626 0 net=7737
rlabel metal2 324 -1628 324 -1628 0 net=1753
rlabel metal2 436 -1628 436 -1628 0 net=3357
rlabel metal2 1206 -1628 1206 -1628 0 net=6853
rlabel metal2 1388 -1628 1388 -1628 0 net=7973
rlabel metal2 317 -1630 317 -1630 0 net=1743
rlabel metal2 1290 -1630 1290 -1630 0 net=7649
rlabel metal2 1437 -1630 1437 -1630 0 net=8305
rlabel metal2 37 -1632 37 -1632 0 net=1395
rlabel metal2 1423 -1632 1423 -1632 0 net=8369
rlabel metal2 37 -1634 37 -1634 0 net=5499
rlabel metal2 2 -1645 2 -1645 0 net=3512
rlabel metal2 446 -1645 446 -1645 0 net=380
rlabel metal2 488 -1645 488 -1645 0 net=6854
rlabel metal2 1283 -1645 1283 -1645 0 net=6756
rlabel metal2 1377 -1645 1377 -1645 0 net=2864
rlabel metal2 23 -1647 23 -1647 0 net=1141
rlabel metal2 23 -1647 23 -1647 0 net=1141
rlabel metal2 37 -1647 37 -1647 0 net=5500
rlabel metal2 429 -1647 429 -1647 0 net=2257
rlabel metal2 471 -1647 471 -1647 0 net=3394
rlabel metal2 621 -1647 621 -1647 0 net=4822
rlabel metal2 800 -1647 800 -1647 0 net=4579
rlabel metal2 800 -1647 800 -1647 0 net=4579
rlabel metal2 814 -1647 814 -1647 0 net=5739
rlabel metal2 1206 -1647 1206 -1647 0 net=7361
rlabel metal2 37 -1649 37 -1649 0 net=4217
rlabel metal2 429 -1649 429 -1649 0 net=2779
rlabel metal2 555 -1649 555 -1649 0 net=4430
rlabel metal2 709 -1649 709 -1649 0 net=4254
rlabel metal2 877 -1649 877 -1649 0 net=5646
rlabel metal2 1017 -1649 1017 -1649 0 net=6537
rlabel metal2 1283 -1649 1283 -1649 0 net=7763
rlabel metal2 51 -1651 51 -1651 0 net=3191
rlabel metal2 51 -1651 51 -1651 0 net=3191
rlabel metal2 65 -1651 65 -1651 0 net=4724
rlabel metal2 597 -1651 597 -1651 0 net=5155
rlabel metal2 877 -1651 877 -1651 0 net=7797
rlabel metal2 1367 -1651 1367 -1651 0 net=2856
rlabel metal2 65 -1653 65 -1653 0 net=1063
rlabel metal2 163 -1653 163 -1653 0 net=2642
rlabel metal2 436 -1653 436 -1653 0 net=1601
rlabel metal2 828 -1653 828 -1653 0 net=6844
rlabel metal2 1150 -1653 1150 -1653 0 net=6903
rlabel metal2 72 -1655 72 -1655 0 net=4826
rlabel metal2 513 -1655 513 -1655 0 net=3218
rlabel metal2 744 -1655 744 -1655 0 net=3472
rlabel metal2 817 -1655 817 -1655 0 net=7353
rlabel metal2 82 -1657 82 -1657 0 net=4280
rlabel metal2 635 -1657 635 -1657 0 net=5670
rlabel metal2 828 -1657 828 -1657 0 net=5467
rlabel metal2 1094 -1657 1094 -1657 0 net=7377
rlabel metal2 128 -1659 128 -1659 0 net=3540
rlabel metal2 653 -1659 653 -1659 0 net=3927
rlabel metal2 667 -1659 667 -1659 0 net=2797
rlabel metal2 709 -1659 709 -1659 0 net=4041
rlabel metal2 719 -1659 719 -1659 0 net=2992
rlabel metal2 1006 -1659 1006 -1659 0 net=7827
rlabel metal2 128 -1661 128 -1661 0 net=1225
rlabel metal2 149 -1661 149 -1661 0 net=1217
rlabel metal2 240 -1661 240 -1661 0 net=2294
rlabel metal2 387 -1661 387 -1661 0 net=2599
rlabel metal2 513 -1661 513 -1661 0 net=5005
rlabel metal2 555 -1661 555 -1661 0 net=3861
rlabel metal2 604 -1661 604 -1661 0 net=3333
rlabel metal2 723 -1661 723 -1661 0 net=4132
rlabel metal2 933 -1661 933 -1661 0 net=6203
rlabel metal2 9 -1663 9 -1663 0 net=2776
rlabel metal2 471 -1663 471 -1663 0 net=2077
rlabel metal2 751 -1663 751 -1663 0 net=8217
rlabel metal2 9 -1665 9 -1665 0 net=2483
rlabel metal2 121 -1665 121 -1665 0 net=2465
rlabel metal2 142 -1665 142 -1665 0 net=2295
rlabel metal2 240 -1665 240 -1665 0 net=1077
rlabel metal2 303 -1665 303 -1665 0 net=1470
rlabel metal2 359 -1665 359 -1665 0 net=5470
rlabel metal2 653 -1665 653 -1665 0 net=4113
rlabel metal2 751 -1665 751 -1665 0 net=4927
rlabel metal2 863 -1665 863 -1665 0 net=5185
rlabel metal2 968 -1665 968 -1665 0 net=5973
rlabel metal2 1080 -1665 1080 -1665 0 net=6733
rlabel metal2 93 -1667 93 -1667 0 net=3249
rlabel metal2 562 -1667 562 -1667 0 net=5766
rlabel metal2 114 -1669 114 -1669 0 net=1867
rlabel metal2 310 -1669 310 -1669 0 net=2588
rlabel metal2 527 -1669 527 -1669 0 net=4055
rlabel metal2 565 -1669 565 -1669 0 net=5594
rlabel metal2 821 -1669 821 -1669 0 net=5351
rlabel metal2 891 -1669 891 -1669 0 net=5535
rlabel metal2 1038 -1669 1038 -1669 0 net=6499
rlabel metal2 1255 -1669 1255 -1669 0 net=7651
rlabel metal2 79 -1671 79 -1671 0 net=1715
rlabel metal2 121 -1671 121 -1671 0 net=1435
rlabel metal2 163 -1671 163 -1671 0 net=1013
rlabel metal2 198 -1671 198 -1671 0 net=1678
rlabel metal2 310 -1671 310 -1671 0 net=2705
rlabel metal2 408 -1671 408 -1671 0 net=3113
rlabel metal2 590 -1671 590 -1671 0 net=3547
rlabel metal2 758 -1671 758 -1671 0 net=5402
rlabel metal2 845 -1671 845 -1671 0 net=7349
rlabel metal2 1290 -1671 1290 -1671 0 net=7789
rlabel metal2 58 -1673 58 -1673 0 net=2153
rlabel metal2 177 -1673 177 -1673 0 net=1006
rlabel metal2 604 -1673 604 -1673 0 net=3613
rlabel metal2 786 -1673 786 -1673 0 net=7229
rlabel metal2 58 -1675 58 -1675 0 net=4471
rlabel metal2 625 -1675 625 -1675 0 net=3381
rlabel metal2 758 -1675 758 -1675 0 net=5757
rlabel metal2 79 -1677 79 -1677 0 net=1744
rlabel metal2 345 -1677 345 -1677 0 net=2729
rlabel metal2 485 -1677 485 -1677 0 net=3127
rlabel metal2 765 -1677 765 -1677 0 net=5673
rlabel metal2 1031 -1677 1031 -1677 0 net=6565
rlabel metal2 110 -1679 110 -1679 0 net=6259
rlabel metal2 492 -1679 492 -1679 0 net=4695
rlabel metal2 660 -1679 660 -1679 0 net=4259
rlabel metal2 779 -1679 779 -1679 0 net=4731
rlabel metal2 880 -1679 880 -1679 0 net=6116
rlabel metal2 1157 -1679 1157 -1679 0 net=6987
rlabel metal2 110 -1681 110 -1681 0 net=1116
rlabel metal2 884 -1681 884 -1681 0 net=5415
rlabel metal2 926 -1681 926 -1681 0 net=7121
rlabel metal2 142 -1683 142 -1683 0 net=4173
rlabel metal2 730 -1683 730 -1683 0 net=4991
rlabel metal2 905 -1683 905 -1683 0 net=3513
rlabel metal2 177 -1685 177 -1685 0 net=3749
rlabel metal2 835 -1685 835 -1685 0 net=5169
rlabel metal2 926 -1685 926 -1685 0 net=6277
rlabel metal2 184 -1687 184 -1687 0 net=2865
rlabel metal2 506 -1687 506 -1687 0 net=7567
rlabel metal2 198 -1689 198 -1689 0 net=1253
rlabel metal2 961 -1689 961 -1689 0 net=5713
rlabel metal2 1010 -1689 1010 -1689 0 net=6683
rlabel metal2 205 -1691 205 -1691 0 net=2194
rlabel metal2 576 -1691 576 -1691 0 net=4407
rlabel metal2 842 -1691 842 -1691 0 net=7348
rlabel metal2 205 -1693 205 -1693 0 net=1727
rlabel metal2 268 -1693 268 -1693 0 net=2041
rlabel metal2 576 -1693 576 -1693 0 net=1831
rlabel metal2 1101 -1693 1101 -1693 0 net=6915
rlabel metal2 1227 -1693 1227 -1693 0 net=8207
rlabel metal2 219 -1695 219 -1695 0 net=1391
rlabel metal2 268 -1695 268 -1695 0 net=1397
rlabel metal2 359 -1695 359 -1695 0 net=2979
rlabel metal2 611 -1695 611 -1695 0 net=3877
rlabel metal2 849 -1695 849 -1695 0 net=5435
rlabel metal2 947 -1695 947 -1695 0 net=6019
rlabel metal2 1220 -1695 1220 -1695 0 net=7481
rlabel metal2 219 -1697 219 -1697 0 net=2883
rlabel metal2 870 -1697 870 -1697 0 net=7596
rlabel metal2 1248 -1697 1248 -1697 0 net=7047
rlabel metal2 254 -1699 254 -1699 0 net=1291
rlabel metal2 464 -1699 464 -1699 0 net=2653
rlabel metal2 611 -1699 611 -1699 0 net=5121
rlabel metal2 901 -1699 901 -1699 0 net=6757
rlabel metal2 289 -1701 289 -1701 0 net=2397
rlabel metal2 366 -1701 366 -1701 0 net=6263
rlabel metal2 856 -1701 856 -1701 0 net=5393
rlabel metal2 919 -1701 919 -1701 0 net=6255
rlabel metal2 1234 -1701 1234 -1701 0 net=7975
rlabel metal2 212 -1703 212 -1703 0 net=5682
rlabel metal2 394 -1703 394 -1703 0 net=3077
rlabel metal2 898 -1703 898 -1703 0 net=4366
rlabel metal2 954 -1703 954 -1703 0 net=6441
rlabel metal2 131 -1705 131 -1705 0 net=7095
rlabel metal2 212 -1707 212 -1707 0 net=2105
rlabel metal2 282 -1707 282 -1707 0 net=1481
rlabel metal2 296 -1707 296 -1707 0 net=3533
rlabel metal2 394 -1707 394 -1707 0 net=1755
rlabel metal2 478 -1707 478 -1707 0 net=3041
rlabel metal2 940 -1707 940 -1707 0 net=5559
rlabel metal2 982 -1707 982 -1707 0 net=6025
rlabel metal2 1087 -1707 1087 -1707 0 net=6787
rlabel metal2 75 -1709 75 -1709 0 net=1159
rlabel metal2 401 -1709 401 -1709 0 net=3359
rlabel metal2 975 -1709 975 -1709 0 net=6409
rlabel metal2 1192 -1709 1192 -1709 0 net=7069
rlabel metal2 75 -1711 75 -1711 0 net=4485
rlabel metal2 996 -1711 996 -1711 0 net=7193
rlabel metal2 1262 -1711 1262 -1711 0 net=7657
rlabel metal2 107 -1713 107 -1713 0 net=1423
rlabel metal2 282 -1713 282 -1713 0 net=2759
rlabel metal2 380 -1713 380 -1713 0 net=5135
rlabel metal2 996 -1713 996 -1713 0 net=6291
rlabel metal2 1332 -1713 1332 -1713 0 net=8111
rlabel metal2 72 -1715 72 -1715 0 net=3447
rlabel metal2 422 -1715 422 -1715 0 net=3280
rlabel metal2 1024 -1715 1024 -1715 0 net=4971
rlabel metal2 107 -1717 107 -1717 0 net=4708
rlabel metal2 502 -1717 502 -1717 0 net=6547
rlabel metal2 1045 -1717 1045 -1717 0 net=6609
rlabel metal2 1402 -1717 1402 -1717 0 net=8371
rlabel metal2 247 -1719 247 -1719 0 net=1269
rlabel metal2 534 -1719 534 -1719 0 net=5829
rlabel metal2 1052 -1719 1052 -1719 0 net=7055
rlabel metal2 1164 -1719 1164 -1719 0 net=7175
rlabel metal2 1423 -1719 1423 -1719 0 net=8307
rlabel metal2 145 -1721 145 -1721 0 net=3397
rlabel metal2 331 -1721 331 -1721 0 net=2573
rlabel metal2 793 -1721 793 -1721 0 net=7846
rlabel metal2 331 -1723 331 -1723 0 net=2495
rlabel metal2 810 -1723 810 -1723 0 net=6685
rlabel metal2 1066 -1723 1066 -1723 0 net=4867
rlabel metal2 338 -1725 338 -1725 0 net=2827
rlabel metal2 992 -1725 992 -1725 0 net=7875
rlabel metal2 30 -1727 30 -1727 0 net=1692
rlabel metal2 992 -1727 992 -1727 0 net=6762
rlabel metal2 16 -1729 16 -1729 0 net=1189
rlabel metal2 646 -1729 646 -1729 0 net=8141
rlabel metal2 16 -1731 16 -1731 0 net=2409
rlabel metal2 646 -1731 646 -1731 0 net=3583
rlabel metal2 1066 -1731 1066 -1731 0 net=6367
rlabel metal2 1276 -1731 1276 -1731 0 net=7739
rlabel metal2 100 -1733 100 -1733 0 net=2959
rlabel metal2 530 -1733 530 -1733 0 net=7029
rlabel metal2 191 -1735 191 -1735 0 net=1745
rlabel metal2 681 -1735 681 -1735 0 net=4243
rlabel metal2 716 -1735 716 -1735 0 net=4747
rlabel metal2 702 -1737 702 -1737 0 net=5475
rlabel metal2 1073 -1737 1073 -1737 0 net=6719
rlabel metal2 772 -1739 772 -1739 0 net=5630
rlabel metal2 1108 -1741 1108 -1741 0 net=6465
rlabel metal2 1178 -1741 1178 -1741 0 net=7897
rlabel metal2 1136 -1743 1136 -1743 0 net=7581
rlabel metal2 1374 -1743 1374 -1743 0 net=2265
rlabel metal2 618 -1745 618 -1745 0 net=8227
rlabel metal2 44 -1747 44 -1747 0 net=3655
rlabel metal2 1213 -1747 1213 -1747 0 net=7723
rlabel metal2 44 -1749 44 -1749 0 net=2119
rlabel metal2 1213 -1749 1213 -1749 0 net=6597
rlabel metal2 86 -1751 86 -1751 0 net=1635
rlabel metal2 1353 -1751 1353 -1751 0 net=7277
rlabel metal2 86 -1753 86 -1753 0 net=1097
rlabel metal2 1353 -1753 1353 -1753 0 net=8435
rlabel metal2 170 -1755 170 -1755 0 net=2907
rlabel metal2 912 -1755 912 -1755 0 net=5365
rlabel metal2 457 -1757 457 -1757 0 net=2517
rlabel metal2 912 -1757 912 -1757 0 net=5815
rlabel metal2 1059 -1759 1059 -1759 0 net=6403
rlabel metal2 2 -1770 2 -1770 0 net=3549
rlabel metal2 667 -1770 667 -1770 0 net=2798
rlabel metal2 877 -1770 877 -1770 0 net=6988
rlabel metal2 1164 -1770 1164 -1770 0 net=7177
rlabel metal2 1164 -1770 1164 -1770 0 net=7177
rlabel metal2 1255 -1770 1255 -1770 0 net=7653
rlabel metal2 1360 -1770 1360 -1770 0 net=4748
rlabel metal2 1377 -1770 1377 -1770 0 net=7278
rlabel metal2 1423 -1770 1423 -1770 0 net=8309
rlabel metal2 1423 -1770 1423 -1770 0 net=8309
rlabel metal2 19 -1772 19 -1772 0 net=5830
rlabel metal2 562 -1772 562 -1772 0 net=4056
rlabel metal2 667 -1772 667 -1772 0 net=4245
rlabel metal2 684 -1772 684 -1772 0 net=7230
rlabel metal2 793 -1772 793 -1772 0 net=5170
rlabel metal2 842 -1772 842 -1772 0 net=5187
rlabel metal2 887 -1772 887 -1772 0 net=5974
rlabel metal2 1003 -1772 1003 -1772 0 net=6368
rlabel metal2 1255 -1772 1255 -1772 0 net=7659
rlabel metal2 1367 -1772 1367 -1772 0 net=8372
rlabel metal2 61 -1774 61 -1774 0 net=8208
rlabel metal2 1346 -1774 1346 -1774 0 net=8219
rlabel metal2 1381 -1774 1381 -1774 0 net=2267
rlabel metal2 72 -1776 72 -1776 0 net=746
rlabel metal2 800 -1776 800 -1776 0 net=4580
rlabel metal2 814 -1776 814 -1776 0 net=5741
rlabel metal2 849 -1776 849 -1776 0 net=5437
rlabel metal2 898 -1776 898 -1776 0 net=7070
rlabel metal2 1339 -1776 1339 -1776 0 net=8143
rlabel metal2 1353 -1776 1353 -1776 0 net=8437
rlabel metal2 30 -1778 30 -1778 0 net=1191
rlabel metal2 75 -1778 75 -1778 0 net=4174
rlabel metal2 177 -1778 177 -1778 0 net=3751
rlabel metal2 177 -1778 177 -1778 0 net=3751
rlabel metal2 198 -1778 198 -1778 0 net=1255
rlabel metal2 198 -1778 198 -1778 0 net=1255
rlabel metal2 205 -1778 205 -1778 0 net=1729
rlabel metal2 205 -1778 205 -1778 0 net=1729
rlabel metal2 247 -1778 247 -1778 0 net=3398
rlabel metal2 898 -1778 898 -1778 0 net=5561
rlabel metal2 968 -1778 968 -1778 0 net=6405
rlabel metal2 1066 -1778 1066 -1778 0 net=6466
rlabel metal2 1332 -1778 1332 -1778 0 net=8113
rlabel metal2 1353 -1778 1353 -1778 0 net=8167
rlabel metal2 23 -1780 23 -1780 0 net=1143
rlabel metal2 89 -1780 89 -1780 0 net=2706
rlabel metal2 324 -1780 324 -1780 0 net=3534
rlabel metal2 373 -1780 373 -1780 0 net=1270
rlabel metal2 513 -1780 513 -1780 0 net=5007
rlabel metal2 793 -1780 793 -1780 0 net=2799
rlabel metal2 23 -1782 23 -1782 0 net=2051
rlabel metal2 635 -1782 635 -1782 0 net=7331
rlabel metal2 1234 -1782 1234 -1782 0 net=7977
rlabel metal2 51 -1784 51 -1784 0 net=3193
rlabel metal2 674 -1784 674 -1784 0 net=3335
rlabel metal2 674 -1784 674 -1784 0 net=3335
rlabel metal2 691 -1784 691 -1784 0 net=6758
rlabel metal2 1325 -1784 1325 -1784 0 net=8229
rlabel metal2 51 -1786 51 -1786 0 net=1437
rlabel metal2 138 -1786 138 -1786 0 net=60
rlabel metal2 436 -1786 436 -1786 0 net=1603
rlabel metal2 464 -1786 464 -1786 0 net=2654
rlabel metal2 513 -1786 513 -1786 0 net=3079
rlabel metal2 569 -1786 569 -1786 0 net=5137
rlabel metal2 849 -1786 849 -1786 0 net=5395
rlabel metal2 863 -1786 863 -1786 0 net=5537
rlabel metal2 908 -1786 908 -1786 0 net=6904
rlabel metal2 1178 -1786 1178 -1786 0 net=7899
rlabel metal2 58 -1788 58 -1788 0 net=4473
rlabel metal2 191 -1788 191 -1788 0 net=1747
rlabel metal2 380 -1788 380 -1788 0 net=3449
rlabel metal2 569 -1788 569 -1788 0 net=5674
rlabel metal2 800 -1788 800 -1788 0 net=6684
rlabel metal2 1129 -1788 1129 -1788 0 net=7097
rlabel metal2 1234 -1788 1234 -1788 0 net=4869
rlabel metal2 9 -1790 9 -1790 0 net=2484
rlabel metal2 82 -1790 82 -1790 0 net=5991
rlabel metal2 926 -1790 926 -1790 0 net=6279
rlabel metal2 1241 -1790 1241 -1790 0 net=7569
rlabel metal2 9 -1792 9 -1792 0 net=2155
rlabel metal2 191 -1792 191 -1792 0 net=1399
rlabel metal2 275 -1792 275 -1792 0 net=1424
rlabel metal2 716 -1792 716 -1792 0 net=6875
rlabel metal2 1136 -1792 1136 -1792 0 net=7583
rlabel metal2 37 -1794 37 -1794 0 net=4219
rlabel metal2 212 -1794 212 -1794 0 net=2107
rlabel metal2 289 -1794 289 -1794 0 net=1482
rlabel metal2 310 -1794 310 -1794 0 net=4793
rlabel metal2 436 -1794 436 -1794 0 net=2519
rlabel metal2 464 -1794 464 -1794 0 net=4409
rlabel metal2 719 -1794 719 -1794 0 net=6026
rlabel metal2 989 -1794 989 -1794 0 net=7013
rlabel metal2 107 -1796 107 -1796 0 net=46
rlabel metal2 415 -1796 415 -1796 0 net=3615
rlabel metal2 611 -1796 611 -1796 0 net=5123
rlabel metal2 810 -1796 810 -1796 0 net=8329
rlabel metal2 100 -1798 100 -1798 0 net=2961
rlabel metal2 114 -1798 114 -1798 0 net=1717
rlabel metal2 212 -1798 212 -1798 0 net=3631
rlabel metal2 380 -1798 380 -1798 0 net=2259
rlabel metal2 527 -1798 527 -1798 0 net=4928
rlabel metal2 765 -1798 765 -1798 0 net=4733
rlabel metal2 803 -1798 803 -1798 0 net=7541
rlabel metal2 1258 -1798 1258 -1798 0 net=1
rlabel metal2 100 -1800 100 -1800 0 net=2867
rlabel metal2 226 -1800 226 -1800 0 net=1637
rlabel metal2 296 -1800 296 -1800 0 net=1161
rlabel metal2 387 -1800 387 -1800 0 net=2601
rlabel metal2 527 -1800 527 -1800 0 net=5477
rlabel metal2 719 -1800 719 -1800 0 net=5468
rlabel metal2 856 -1800 856 -1800 0 net=5417
rlabel metal2 926 -1800 926 -1800 0 net=5715
rlabel metal2 989 -1800 989 -1800 0 net=7195
rlabel metal2 65 -1802 65 -1802 0 net=1065
rlabel metal2 247 -1802 247 -1802 0 net=1293
rlabel metal2 261 -1802 261 -1802 0 net=1392
rlabel metal2 534 -1802 534 -1802 0 net=4993
rlabel metal2 737 -1802 737 -1802 0 net=3128
rlabel metal2 779 -1802 779 -1802 0 net=7483
rlabel metal2 65 -1804 65 -1804 0 net=1099
rlabel metal2 114 -1804 114 -1804 0 net=1219
rlabel metal2 163 -1804 163 -1804 0 net=1015
rlabel metal2 233 -1804 233 -1804 0 net=2297
rlabel metal2 296 -1804 296 -1804 0 net=130
rlabel metal2 1094 -1804 1094 -1804 0 net=7379
rlabel metal2 135 -1806 135 -1806 0 net=2467
rlabel metal2 163 -1806 163 -1806 0 net=2909
rlabel metal2 233 -1806 233 -1806 0 net=2731
rlabel metal2 352 -1806 352 -1806 0 net=2829
rlabel metal2 485 -1806 485 -1806 0 net=5325
rlabel metal2 919 -1806 919 -1806 0 net=6257
rlabel metal2 37 -1808 37 -1808 0 net=3689
rlabel metal2 240 -1808 240 -1808 0 net=1079
rlabel metal2 324 -1808 324 -1808 0 net=1833
rlabel metal2 604 -1808 604 -1808 0 net=3657
rlabel metal2 695 -1808 695 -1808 0 net=4487
rlabel metal2 737 -1808 737 -1808 0 net=6539
rlabel metal2 1087 -1808 1087 -1808 0 net=6789
rlabel metal2 1122 -1808 1122 -1808 0 net=7057
rlabel metal2 44 -1810 44 -1810 0 net=2120
rlabel metal2 352 -1810 352 -1810 0 net=2079
rlabel metal2 488 -1810 488 -1810 0 net=4343
rlabel metal2 611 -1810 611 -1810 0 net=3585
rlabel metal2 702 -1810 702 -1810 0 net=4043
rlabel metal2 723 -1810 723 -1810 0 net=3603
rlabel metal2 940 -1810 940 -1810 0 net=5367
rlabel metal2 44 -1812 44 -1812 0 net=6261
rlabel metal2 492 -1812 492 -1812 0 net=4697
rlabel metal2 744 -1812 744 -1812 0 net=6265
rlabel metal2 996 -1812 996 -1812 0 net=6293
rlabel metal2 1006 -1812 1006 -1812 0 net=7048
rlabel metal2 93 -1814 93 -1814 0 net=3251
rlabel metal2 240 -1814 240 -1814 0 net=2575
rlabel metal2 530 -1814 530 -1814 0 net=1793
rlabel metal2 751 -1814 751 -1814 0 net=6075
rlabel metal2 975 -1814 975 -1814 0 net=6411
rlabel metal2 1073 -1814 1073 -1814 0 net=6721
rlabel metal2 1311 -1814 1311 -1814 0 net=7877
rlabel metal2 93 -1816 93 -1816 0 net=5647
rlabel metal2 450 -1816 450 -1816 0 net=2559
rlabel metal2 821 -1816 821 -1816 0 net=5353
rlabel metal2 870 -1816 870 -1816 0 net=8407
rlabel metal2 128 -1818 128 -1818 0 net=1227
rlabel metal2 506 -1818 506 -1818 0 net=6227
rlabel metal2 996 -1818 996 -1818 0 net=7123
rlabel metal2 1304 -1818 1304 -1818 0 net=7829
rlabel metal2 128 -1820 128 -1820 0 net=1829
rlabel metal2 597 -1820 597 -1820 0 net=5157
rlabel metal2 870 -1820 870 -1820 0 net=5817
rlabel metal2 919 -1820 919 -1820 0 net=6735
rlabel metal2 1115 -1820 1115 -1820 0 net=7031
rlabel metal2 1297 -1820 1297 -1820 0 net=7799
rlabel metal2 317 -1822 317 -1822 0 net=2399
rlabel metal2 478 -1822 478 -1822 0 net=3043
rlabel metal2 541 -1822 541 -1822 0 net=3115
rlabel metal2 555 -1822 555 -1822 0 net=3863
rlabel metal2 618 -1822 618 -1822 0 net=6549
rlabel metal2 1045 -1822 1045 -1822 0 net=6611
rlabel metal2 1290 -1822 1290 -1822 0 net=7791
rlabel metal2 282 -1824 282 -1824 0 net=2761
rlabel metal2 331 -1824 331 -1824 0 net=2497
rlabel metal2 432 -1824 432 -1824 0 net=6523
rlabel metal2 1052 -1824 1052 -1824 0 net=6687
rlabel metal2 1283 -1824 1283 -1824 0 net=7765
rlabel metal2 282 -1826 282 -1826 0 net=2981
rlabel metal2 387 -1826 387 -1826 0 net=4115
rlabel metal2 681 -1826 681 -1826 0 net=6925
rlabel metal2 219 -1828 219 -1828 0 net=2885
rlabel metal2 401 -1828 401 -1828 0 net=3361
rlabel metal2 555 -1828 555 -1828 0 net=3928
rlabel metal2 709 -1828 709 -1828 0 net=3515
rlabel metal2 933 -1828 933 -1828 0 net=6205
rlabel metal2 1031 -1828 1031 -1828 0 net=6567
rlabel metal2 1101 -1828 1101 -1828 0 net=6917
rlabel metal2 79 -1830 79 -1830 0 net=2453
rlabel metal2 303 -1830 303 -1830 0 net=1869
rlabel metal2 338 -1830 338 -1830 0 net=4833
rlabel metal2 558 -1830 558 -1830 0 net=5697
rlabel metal2 1010 -1830 1010 -1830 0 net=7363
rlabel metal2 16 -1832 16 -1832 0 net=2411
rlabel metal2 303 -1832 303 -1832 0 net=1757
rlabel metal2 401 -1832 401 -1832 0 net=2347
rlabel metal2 873 -1832 873 -1832 0 net=8251
rlabel metal2 1185 -1832 1185 -1832 0 net=7351
rlabel metal2 86 -1834 86 -1834 0 net=7289
rlabel metal2 338 -1836 338 -1836 0 net=4817
rlabel metal2 586 -1836 586 -1836 0 net=367
rlabel metal2 1031 -1836 1031 -1836 0 net=6501
rlabel metal2 1101 -1836 1101 -1836 0 net=4973
rlabel metal2 341 -1838 341 -1838 0 net=6598
rlabel metal2 394 -1840 394 -1840 0 net=8181
rlabel metal2 478 -1842 478 -1842 0 net=2043
rlabel metal2 583 -1842 583 -1842 0 net=3879
rlabel metal2 653 -1842 653 -1842 0 net=5759
rlabel metal2 901 -1842 901 -1842 0 net=8373
rlabel metal2 289 -1844 289 -1844 0 net=4595
rlabel metal2 625 -1844 625 -1844 0 net=3383
rlabel metal2 688 -1844 688 -1844 0 net=7239
rlabel metal2 1199 -1844 1199 -1844 0 net=7355
rlabel metal2 625 -1846 625 -1846 0 net=4261
rlabel metal2 716 -1846 716 -1846 0 net=4935
rlabel metal2 954 -1846 954 -1846 0 net=6443
rlabel metal2 639 -1848 639 -1848 0 net=2159
rlabel metal2 947 -1848 947 -1848 0 net=6021
rlabel metal2 1038 -1848 1038 -1848 0 net=7741
rlabel metal2 572 -1850 572 -1850 0 net=6027
rlabel metal2 1269 -1850 1269 -1850 0 net=7725
rlabel metal2 660 -1852 660 -1852 0 net=8337
rlabel metal2 772 -1854 772 -1854 0 net=7665
rlabel metal2 429 -1856 429 -1856 0 net=2780
rlabel metal2 2 -1867 2 -1867 0 net=3551
rlabel metal2 9 -1867 9 -1867 0 net=2156
rlabel metal2 432 -1867 432 -1867 0 net=1794
rlabel metal2 751 -1867 751 -1867 0 net=6918
rlabel metal2 1395 -1867 1395 -1867 0 net=8310
rlabel metal2 2 -1869 2 -1869 0 net=1439
rlabel metal2 100 -1869 100 -1869 0 net=2868
rlabel metal2 303 -1869 303 -1869 0 net=1759
rlabel metal2 303 -1869 303 -1869 0 net=1759
rlabel metal2 373 -1869 373 -1869 0 net=1748
rlabel metal2 565 -1869 565 -1869 0 net=5698
rlabel metal2 933 -1869 933 -1869 0 net=8438
rlabel metal2 9 -1871 9 -1871 0 net=2299
rlabel metal2 282 -1871 282 -1871 0 net=2982
rlabel metal2 471 -1871 471 -1871 0 net=1228
rlabel metal2 618 -1871 618 -1871 0 net=6550
rlabel metal2 775 -1871 775 -1871 0 net=6406
rlabel metal2 1062 -1871 1062 -1871 0 net=7654
rlabel metal2 19 -1873 19 -1873 0 net=476
rlabel metal2 100 -1873 100 -1873 0 net=1221
rlabel metal2 128 -1873 128 -1873 0 net=1830
rlabel metal2 968 -1873 968 -1873 0 net=6229
rlabel metal2 1234 -1873 1234 -1873 0 net=4871
rlabel metal2 26 -1875 26 -1875 0 net=1144
rlabel metal2 37 -1875 37 -1875 0 net=3690
rlabel metal2 401 -1875 401 -1875 0 net=2349
rlabel metal2 499 -1875 499 -1875 0 net=3864
rlabel metal2 618 -1875 618 -1875 0 net=2427
rlabel metal2 856 -1875 856 -1875 0 net=5419
rlabel metal2 912 -1875 912 -1875 0 net=5717
rlabel metal2 933 -1875 933 -1875 0 net=6295
rlabel metal2 1066 -1875 1066 -1875 0 net=7663
rlabel metal2 30 -1877 30 -1877 0 net=1605
rlabel metal2 502 -1877 502 -1877 0 net=8393
rlabel metal2 37 -1879 37 -1879 0 net=6444
rlabel metal2 44 -1881 44 -1881 0 net=6262
rlabel metal2 523 -1881 523 -1881 0 net=7352
rlabel metal2 44 -1883 44 -1883 0 net=3659
rlabel metal2 646 -1883 646 -1883 0 net=3384
rlabel metal2 681 -1883 681 -1883 0 net=113
rlabel metal2 51 -1885 51 -1885 0 net=3633
rlabel metal2 219 -1885 219 -1885 0 net=2455
rlabel metal2 527 -1885 527 -1885 0 net=5479
rlabel metal2 604 -1885 604 -1885 0 net=3941
rlabel metal2 1199 -1885 1199 -1885 0 net=7585
rlabel metal2 58 -1887 58 -1887 0 net=5575
rlabel metal2 884 -1887 884 -1887 0 net=2268
rlabel metal2 58 -1889 58 -1889 0 net=3081
rlabel metal2 555 -1889 555 -1889 0 net=4263
rlabel metal2 660 -1889 660 -1889 0 net=6280
rlabel metal2 1206 -1889 1206 -1889 0 net=7793
rlabel metal2 40 -1891 40 -1891 0 net=7473
rlabel metal2 1241 -1891 1241 -1891 0 net=7661
rlabel metal2 1297 -1891 1297 -1891 0 net=7979
rlabel metal2 61 -1893 61 -1893 0 net=1407
rlabel metal2 282 -1893 282 -1893 0 net=2401
rlabel metal2 513 -1893 513 -1893 0 net=3604
rlabel metal2 726 -1893 726 -1893 0 net=7245
rlabel metal2 1332 -1893 1332 -1893 0 net=8221
rlabel metal2 79 -1895 79 -1895 0 net=2413
rlabel metal2 219 -1895 219 -1895 0 net=2081
rlabel metal2 355 -1895 355 -1895 0 net=6543
rlabel metal2 996 -1895 996 -1895 0 net=7125
rlabel metal2 1122 -1895 1122 -1895 0 net=8253
rlabel metal2 79 -1897 79 -1897 0 net=1719
rlabel metal2 170 -1897 170 -1897 0 net=3252
rlabel metal2 688 -1897 688 -1897 0 net=6258
rlabel metal2 1255 -1897 1255 -1897 0 net=7831
rlabel metal2 89 -1899 89 -1899 0 net=4677
rlabel metal2 660 -1899 660 -1899 0 net=5063
rlabel metal2 691 -1899 691 -1899 0 net=7503
rlabel metal2 1311 -1899 1311 -1899 0 net=8115
rlabel metal2 121 -1901 121 -1901 0 net=4475
rlabel metal2 625 -1901 625 -1901 0 net=3517
rlabel metal2 737 -1901 737 -1901 0 net=6541
rlabel metal2 1003 -1901 1003 -1901 0 net=6613
rlabel metal2 1122 -1901 1122 -1901 0 net=7381
rlabel metal2 1339 -1901 1339 -1901 0 net=8331
rlabel metal2 121 -1903 121 -1903 0 net=3045
rlabel metal2 702 -1903 702 -1903 0 net=4044
rlabel metal2 737 -1903 737 -1903 0 net=5125
rlabel metal2 870 -1903 870 -1903 0 net=5819
rlabel metal2 926 -1903 926 -1903 0 net=6413
rlabel metal2 1038 -1903 1038 -1903 0 net=7743
rlabel metal2 1388 -1903 1388 -1903 0 net=8409
rlabel metal2 128 -1905 128 -1905 0 net=2831
rlabel metal2 506 -1905 506 -1905 0 net=7570
rlabel metal2 135 -1907 135 -1907 0 net=7032
rlabel metal2 1248 -1907 1248 -1907 0 net=7801
rlabel metal2 135 -1909 135 -1909 0 net=2469
rlabel metal2 170 -1909 170 -1909 0 net=8230
rlabel metal2 142 -1911 142 -1911 0 net=2025
rlabel metal2 338 -1911 338 -1911 0 net=4819
rlabel metal2 1038 -1911 1038 -1911 0 net=6877
rlabel metal2 1143 -1911 1143 -1911 0 net=7333
rlabel metal2 1374 -1911 1374 -1911 0 net=8375
rlabel metal2 149 -1913 149 -1913 0 net=4247
rlabel metal2 716 -1913 716 -1913 0 net=8005
rlabel metal2 205 -1915 205 -1915 0 net=1730
rlabel metal2 611 -1915 611 -1915 0 net=3586
rlabel metal2 716 -1915 716 -1915 0 net=4937
rlabel metal2 772 -1915 772 -1915 0 net=5355
rlabel metal2 870 -1915 870 -1915 0 net=5993
rlabel metal2 1059 -1915 1059 -1915 0 net=7015
rlabel metal2 1192 -1915 1192 -1915 0 net=7727
rlabel metal2 205 -1917 205 -1917 0 net=1871
rlabel metal2 338 -1917 338 -1917 0 net=1163
rlabel metal2 387 -1917 387 -1917 0 net=4116
rlabel metal2 744 -1917 744 -1917 0 net=5159
rlabel metal2 828 -1917 828 -1917 0 net=5539
rlabel metal2 891 -1917 891 -1917 0 net=6029
rlabel metal2 1108 -1917 1108 -1917 0 net=8339
rlabel metal2 93 -1919 93 -1919 0 net=5649
rlabel metal2 898 -1919 898 -1919 0 net=5562
rlabel metal2 1024 -1919 1024 -1919 0 net=6207
rlabel metal2 93 -1921 93 -1921 0 net=1257
rlabel metal2 233 -1921 233 -1921 0 net=2732
rlabel metal2 492 -1921 492 -1921 0 net=4835
rlabel metal2 751 -1921 751 -1921 0 net=7217
rlabel metal2 1129 -1921 1129 -1921 0 net=7901
rlabel metal2 198 -1923 198 -1923 0 net=5009
rlabel metal2 800 -1923 800 -1923 0 net=6022
rlabel metal2 1024 -1923 1024 -1923 0 net=6723
rlabel metal2 1276 -1923 1276 -1923 0 net=7879
rlabel metal2 1325 -1923 1325 -1923 0 net=8169
rlabel metal2 86 -1925 86 -1925 0 net=8189
rlabel metal2 86 -1927 86 -1927 0 net=2231
rlabel metal2 352 -1927 352 -1927 0 net=2335
rlabel metal2 408 -1927 408 -1927 0 net=1577
rlabel metal2 569 -1927 569 -1927 0 net=4345
rlabel metal2 611 -1927 611 -1927 0 net=6705
rlabel metal2 723 -1927 723 -1927 0 net=5199
rlabel metal2 800 -1927 800 -1927 0 net=5369
rlabel metal2 954 -1927 954 -1927 0 net=6525
rlabel metal2 1087 -1927 1087 -1927 0 net=7667
rlabel metal2 1318 -1927 1318 -1927 0 net=8145
rlabel metal2 138 -1929 138 -1929 0 net=6185
rlabel metal2 1346 -1929 1346 -1929 0 net=8183
rlabel metal2 233 -1931 233 -1931 0 net=3195
rlabel metal2 653 -1931 653 -1931 0 net=5761
rlabel metal2 940 -1931 940 -1931 0 net=6927
rlabel metal2 240 -1933 240 -1933 0 net=2576
rlabel metal2 754 -1933 754 -1933 0 net=5438
rlabel metal2 989 -1933 989 -1933 0 net=7197
rlabel metal2 240 -1935 240 -1935 0 net=2499
rlabel metal2 429 -1935 429 -1935 0 net=2449
rlabel metal2 989 -1935 989 -1935 0 net=6569
rlabel metal2 1115 -1935 1115 -1935 0 net=7291
rlabel metal2 191 -1937 191 -1937 0 net=1401
rlabel metal2 464 -1937 464 -1937 0 net=4411
rlabel metal2 520 -1937 520 -1937 0 net=2602
rlabel metal2 674 -1937 674 -1937 0 net=3336
rlabel metal2 758 -1937 758 -1937 0 net=4735
rlabel metal2 782 -1937 782 -1937 0 net=4974
rlabel metal2 1150 -1937 1150 -1937 0 net=7099
rlabel metal2 72 -1939 72 -1939 0 net=1193
rlabel metal2 247 -1939 247 -1939 0 net=1295
rlabel metal2 464 -1939 464 -1939 0 net=2801
rlabel metal2 807 -1939 807 -1939 0 net=8087
rlabel metal2 72 -1941 72 -1941 0 net=480
rlabel metal2 254 -1941 254 -1941 0 net=1081
rlabel metal2 254 -1941 254 -1941 0 net=1081
rlabel metal2 268 -1941 268 -1941 0 net=2109
rlabel metal2 485 -1941 485 -1941 0 net=5327
rlabel metal2 821 -1941 821 -1941 0 net=5397
rlabel metal2 1010 -1941 1010 -1941 0 net=7365
rlabel metal2 107 -1943 107 -1943 0 net=2963
rlabel metal2 268 -1943 268 -1943 0 net=1639
rlabel metal2 289 -1943 289 -1943 0 net=4597
rlabel metal2 765 -1943 765 -1943 0 net=5139
rlabel metal2 835 -1943 835 -1943 0 net=5743
rlabel metal2 1010 -1943 1010 -1943 0 net=6689
rlabel metal2 1101 -1943 1101 -1943 0 net=7241
rlabel metal2 16 -1945 16 -1945 0 net=3153
rlabel metal2 163 -1945 163 -1945 0 net=2911
rlabel metal2 296 -1945 296 -1945 0 net=3117
rlabel metal2 572 -1945 572 -1945 0 net=5517
rlabel metal2 835 -1945 835 -1945 0 net=5189
rlabel metal2 1052 -1945 1052 -1945 0 net=6791
rlabel metal2 1178 -1945 1178 -1945 0 net=7543
rlabel metal2 16 -1947 16 -1947 0 net=2053
rlabel metal2 163 -1947 163 -1947 0 net=5301
rlabel metal2 842 -1947 842 -1947 0 net=6077
rlabel metal2 1080 -1947 1080 -1947 0 net=7059
rlabel metal2 23 -1949 23 -1949 0 net=7356
rlabel metal2 229 -1951 229 -1951 0 net=1699
rlabel metal2 310 -1951 310 -1951 0 net=4795
rlabel metal2 579 -1951 579 -1951 0 net=4911
rlabel metal2 705 -1951 705 -1951 0 net=7461
rlabel metal2 1213 -1951 1213 -1951 0 net=7767
rlabel metal2 310 -1953 310 -1953 0 net=1835
rlabel metal2 331 -1953 331 -1953 0 net=3363
rlabel metal2 887 -1953 887 -1953 0 net=7929
rlabel metal2 65 -1955 65 -1955 0 net=1101
rlabel metal2 345 -1955 345 -1955 0 net=2945
rlabel metal2 548 -1955 548 -1955 0 net=3451
rlabel metal2 961 -1955 961 -1955 0 net=6267
rlabel metal2 1094 -1955 1094 -1955 0 net=7179
rlabel metal2 65 -1957 65 -1957 0 net=5141
rlabel metal2 317 -1957 317 -1957 0 net=2762
rlabel metal2 779 -1957 779 -1957 0 net=7485
rlabel metal2 317 -1959 317 -1959 0 net=2521
rlabel metal2 478 -1959 478 -1959 0 net=2045
rlabel metal2 681 -1959 681 -1959 0 net=4683
rlabel metal2 982 -1959 982 -1959 0 net=6503
rlabel metal2 359 -1961 359 -1961 0 net=2887
rlabel metal2 919 -1961 919 -1961 0 net=6737
rlabel metal2 359 -1963 359 -1963 0 net=2561
rlabel metal2 590 -1963 590 -1963 0 net=6177
rlabel metal2 177 -1965 177 -1965 0 net=3753
rlabel metal2 583 -1965 583 -1965 0 net=3881
rlabel metal2 177 -1967 177 -1967 0 net=1017
rlabel metal2 366 -1967 366 -1967 0 net=2161
rlabel metal2 184 -1969 184 -1969 0 net=1066
rlabel metal2 373 -1969 373 -1969 0 net=8031
rlabel metal2 68 -1971 68 -1971 0 net=1425
rlabel metal2 380 -1971 380 -1971 0 net=2260
rlabel metal2 583 -1971 583 -1971 0 net=7713
rlabel metal2 156 -1973 156 -1973 0 net=4221
rlabel metal2 415 -1973 415 -1973 0 net=3617
rlabel metal2 639 -1973 639 -1973 0 net=4417
rlabel metal2 436 -1975 436 -1975 0 net=2055
rlabel metal2 156 -1977 156 -1977 0 net=4489
rlabel metal2 695 -1979 695 -1979 0 net=4699
rlabel metal2 534 -1981 534 -1981 0 net=4995
rlabel metal2 411 -1983 411 -1983 0 net=1315
rlabel metal2 2 -1994 2 -1994 0 net=1440
rlabel metal2 51 -1994 51 -1994 0 net=3634
rlabel metal2 663 -1994 663 -1994 0 net=6542
rlabel metal2 1010 -1994 1010 -1994 0 net=6691
rlabel metal2 1010 -1994 1010 -1994 0 net=6691
rlabel metal2 1024 -1994 1024 -1994 0 net=6725
rlabel metal2 1024 -1994 1024 -1994 0 net=6725
rlabel metal2 1031 -1994 1031 -1994 0 net=6739
rlabel metal2 1031 -1994 1031 -1994 0 net=6739
rlabel metal2 1139 -1994 1139 -1994 0 net=8254
rlabel metal2 5 -1996 5 -1996 0 net=1194
rlabel metal2 205 -1996 205 -1996 0 net=1872
rlabel metal2 324 -1996 324 -1996 0 net=1102
rlabel metal2 408 -1996 408 -1996 0 net=7246
rlabel metal2 37 -1998 37 -1998 0 net=1165
rlabel metal2 408 -1998 408 -1998 0 net=2047
rlabel metal2 579 -1998 579 -1998 0 net=7100
rlabel metal2 1262 -1998 1262 -1998 0 net=8089
rlabel metal2 51 -2000 51 -2000 0 net=1409
rlabel metal2 268 -2000 268 -2000 0 net=1640
rlabel metal2 373 -2000 373 -2000 0 net=7689
rlabel metal2 1283 -2000 1283 -2000 0 net=8171
rlabel metal2 58 -2002 58 -2002 0 net=3082
rlabel metal2 502 -2002 502 -2002 0 net=8006
rlabel metal2 1325 -2002 1325 -2002 0 net=8411
rlabel metal2 58 -2004 58 -2004 0 net=2965
rlabel metal2 261 -2004 261 -2004 0 net=2337
rlabel metal2 411 -2004 411 -2004 0 net=7664
rlabel metal2 65 -2006 65 -2006 0 net=2912
rlabel metal2 334 -2006 334 -2006 0 net=7880
rlabel metal2 65 -2008 65 -2008 0 net=1761
rlabel metal2 338 -2008 338 -2008 0 net=1297
rlabel metal2 415 -2008 415 -2008 0 net=3553
rlabel metal2 614 -2008 614 -2008 0 net=7662
rlabel metal2 68 -2010 68 -2010 0 net=1539
rlabel metal2 373 -2010 373 -2010 0 net=3619
rlabel metal2 513 -2010 513 -2010 0 net=7930
rlabel metal2 72 -2012 72 -2012 0 net=7714
rlabel metal2 1290 -2012 1290 -2012 0 net=8223
rlabel metal2 72 -2014 72 -2014 0 net=3365
rlabel metal2 387 -2014 387 -2014 0 net=4797
rlabel metal2 513 -2014 513 -2014 0 net=3519
rlabel metal2 639 -2014 639 -2014 0 net=7060
rlabel metal2 1108 -2014 1108 -2014 0 net=8341
rlabel metal2 93 -2016 93 -2016 0 net=1259
rlabel metal2 268 -2016 268 -2016 0 net=2451
rlabel metal2 453 -2016 453 -2016 0 net=7953
rlabel metal2 93 -2018 93 -2018 0 net=4479
rlabel metal2 646 -2018 646 -2018 0 net=4679
rlabel metal2 691 -2018 691 -2018 0 net=7198
rlabel metal2 96 -2020 96 -2020 0 net=1222
rlabel metal2 107 -2020 107 -2020 0 net=3155
rlabel metal2 289 -2020 289 -2020 0 net=2057
rlabel metal2 478 -2020 478 -2020 0 net=1579
rlabel metal2 604 -2020 604 -2020 0 net=3943
rlabel metal2 646 -2020 646 -2020 0 net=4685
rlabel metal2 705 -2020 705 -2020 0 net=5356
rlabel metal2 782 -2020 782 -2020 0 net=5398
rlabel metal2 849 -2020 849 -2020 0 net=6296
rlabel metal2 947 -2020 947 -2020 0 net=7334
rlabel metal2 1213 -2020 1213 -2020 0 net=7769
rlabel metal2 100 -2022 100 -2022 0 net=2279
rlabel metal2 177 -2022 177 -2022 0 net=1018
rlabel metal2 415 -2022 415 -2022 0 net=4413
rlabel metal2 516 -2022 516 -2022 0 net=5140
rlabel metal2 807 -2022 807 -2022 0 net=6186
rlabel metal2 1059 -2022 1059 -2022 0 net=7017
rlabel metal2 1129 -2022 1129 -2022 0 net=7903
rlabel metal2 114 -2024 114 -2024 0 net=5143
rlabel metal2 114 -2024 114 -2024 0 net=5143
rlabel metal2 121 -2024 121 -2024 0 net=3047
rlabel metal2 499 -2024 499 -2024 0 net=4477
rlabel metal2 821 -2024 821 -2024 0 net=7586
rlabel metal2 1206 -2024 1206 -2024 0 net=7795
rlabel metal2 1227 -2024 1227 -2024 0 net=7833
rlabel metal2 23 -2026 23 -2026 0 net=2707
rlabel metal2 128 -2026 128 -2026 0 net=2833
rlabel metal2 726 -2026 726 -2026 0 net=6208
rlabel metal2 16 -2028 16 -2028 0 net=2054
rlabel metal2 131 -2028 131 -2028 0 net=6431
rlabel metal2 422 -2028 422 -2028 0 net=1402
rlabel metal2 520 -2028 520 -2028 0 net=3882
rlabel metal2 621 -2028 621 -2028 0 net=8190
rlabel metal2 16 -2030 16 -2030 0 net=2501
rlabel metal2 296 -2030 296 -2030 0 net=3118
rlabel metal2 520 -2030 520 -2030 0 net=4801
rlabel metal2 849 -2030 849 -2030 0 net=5577
rlabel metal2 877 -2030 877 -2030 0 net=5745
rlabel metal2 877 -2030 877 -2030 0 net=5745
rlabel metal2 884 -2030 884 -2030 0 net=5821
rlabel metal2 884 -2030 884 -2030 0 net=5821
rlabel metal2 912 -2030 912 -2030 0 net=5719
rlabel metal2 1129 -2030 1129 -2030 0 net=7463
rlabel metal2 1143 -2030 1143 -2030 0 net=7487
rlabel metal2 1199 -2030 1199 -2030 0 net=7745
rlabel metal2 23 -2032 23 -2032 0 net=4491
rlabel metal2 163 -2032 163 -2032 0 net=5302
rlabel metal2 296 -2032 296 -2032 0 net=1771
rlabel metal2 730 -2032 730 -2032 0 net=4997
rlabel metal2 737 -2032 737 -2032 0 net=5127
rlabel metal2 779 -2032 779 -2032 0 net=7535
rlabel metal2 1206 -2032 1206 -2032 0 net=8147
rlabel metal2 9 -2034 9 -2034 0 net=2300
rlabel metal2 166 -2034 166 -2034 0 net=4820
rlabel metal2 1059 -2034 1059 -2034 0 net=7181
rlabel metal2 1220 -2034 1220 -2034 0 net=7803
rlabel metal2 1318 -2034 1318 -2034 0 net=8395
rlabel metal2 9 -2036 9 -2036 0 net=8047
rlabel metal2 135 -2038 135 -2038 0 net=2471
rlabel metal2 173 -2038 173 -2038 0 net=2414
rlabel metal2 219 -2038 219 -2038 0 net=2083
rlabel metal2 303 -2038 303 -2038 0 net=1837
rlabel metal2 422 -2038 422 -2038 0 net=3755
rlabel metal2 527 -2038 527 -2038 0 net=3453
rlabel metal2 555 -2038 555 -2038 0 net=4265
rlabel metal2 716 -2038 716 -2038 0 net=4939
rlabel metal2 754 -2038 754 -2038 0 net=5762
rlabel metal2 933 -2038 933 -2038 0 net=6221
rlabel metal2 996 -2038 996 -2038 0 net=7383
rlabel metal2 1248 -2038 1248 -2038 0 net=8033
rlabel metal2 110 -2040 110 -2040 0 net=2733
rlabel metal2 219 -2040 219 -2040 0 net=1317
rlabel metal2 548 -2040 548 -2040 0 net=6389
rlabel metal2 842 -2040 842 -2040 0 net=6079
rlabel metal2 968 -2040 968 -2040 0 net=6231
rlabel metal2 1094 -2040 1094 -2040 0 net=7729
rlabel metal2 1269 -2040 1269 -2040 0 net=8117
rlabel metal2 135 -2042 135 -2042 0 net=2531
rlabel metal2 730 -2042 730 -2042 0 net=5371
rlabel metal2 828 -2042 828 -2042 0 net=5541
rlabel metal2 852 -2042 852 -2042 0 net=5420
rlabel metal2 971 -2042 971 -2042 0 net=7980
rlabel metal2 1311 -2042 1311 -2042 0 net=8377
rlabel metal2 142 -2044 142 -2044 0 net=2027
rlabel metal2 429 -2044 429 -2044 0 net=2609
rlabel metal2 856 -2044 856 -2044 0 net=6527
rlabel metal2 1017 -2044 1017 -2044 0 net=7669
rlabel metal2 1101 -2044 1101 -2044 0 net=7243
rlabel metal2 1297 -2044 1297 -2044 0 net=8333
rlabel metal2 142 -2046 142 -2046 0 net=2563
rlabel metal2 436 -2046 436 -2046 0 net=2351
rlabel metal2 485 -2046 485 -2046 0 net=4903
rlabel metal2 765 -2046 765 -2046 0 net=5651
rlabel metal2 870 -2046 870 -2046 0 net=5995
rlabel metal2 954 -2046 954 -2046 0 net=6571
rlabel metal2 1073 -2046 1073 -2046 0 net=7219
rlabel metal2 1101 -2046 1101 -2046 0 net=7293
rlabel metal2 30 -2048 30 -2048 0 net=1607
rlabel metal2 443 -2048 443 -2048 0 net=2110
rlabel metal2 457 -2048 457 -2048 0 net=2889
rlabel metal2 555 -2048 555 -2048 0 net=1125
rlabel metal2 590 -2048 590 -2048 0 net=4599
rlabel metal2 779 -2048 779 -2048 0 net=8184
rlabel metal2 30 -2050 30 -2050 0 net=2617
rlabel metal2 170 -2050 170 -2050 0 net=5853
rlabel metal2 457 -2050 457 -2050 0 net=2803
rlabel metal2 569 -2050 569 -2050 0 net=4347
rlabel metal2 786 -2050 786 -2050 0 net=5201
rlabel metal2 863 -2050 863 -2050 0 net=5683
rlabel metal2 1066 -2050 1066 -2050 0 net=7127
rlabel metal2 75 -2052 75 -2052 0 net=994
rlabel metal2 177 -2052 177 -2052 0 net=1019
rlabel metal2 744 -2052 744 -2052 0 net=5161
rlabel metal2 870 -2052 870 -2052 0 net=7307
rlabel metal2 191 -2054 191 -2054 0 net=2429
rlabel metal2 674 -2054 674 -2054 0 net=4913
rlabel metal2 891 -2054 891 -2054 0 net=6031
rlabel metal2 149 -2056 149 -2056 0 net=4248
rlabel metal2 674 -2056 674 -2056 0 net=4701
rlabel metal2 149 -2058 149 -2058 0 net=7475
rlabel metal2 198 -2060 198 -2060 0 net=5011
rlabel metal2 506 -2060 506 -2060 0 net=7105
rlabel metal2 184 -2062 184 -2062 0 net=1427
rlabel metal2 226 -2062 226 -2062 0 net=3063
rlabel metal2 184 -2064 184 -2064 0 net=1083
rlabel metal2 562 -2064 562 -2064 0 net=7531
rlabel metal2 229 -2066 229 -2066 0 net=1537
rlabel metal2 562 -2066 562 -2066 0 net=6545
rlabel metal2 233 -2068 233 -2068 0 net=3197
rlabel metal2 569 -2068 569 -2068 0 net=4837
rlabel metal2 695 -2068 695 -2068 0 net=5329
rlabel metal2 975 -2068 975 -2068 0 net=6505
rlabel metal2 86 -2070 86 -2070 0 net=2233
rlabel metal2 254 -2070 254 -2070 0 net=2403
rlabel metal2 576 -2070 576 -2070 0 net=5219
rlabel metal2 667 -2070 667 -2070 0 net=7366
rlabel metal2 86 -2072 86 -2072 0 net=3899
rlabel metal2 282 -2072 282 -2072 0 net=2947
rlabel metal2 576 -2072 576 -2072 0 net=6268
rlabel metal2 982 -2072 982 -2072 0 net=4873
rlabel metal2 345 -2074 345 -2074 0 net=2456
rlabel metal2 579 -2074 579 -2074 0 net=6235
rlabel metal2 1150 -2074 1150 -2074 0 net=7505
rlabel metal2 401 -2076 401 -2076 0 net=1411
rlabel metal2 751 -2076 751 -2076 0 net=4737
rlabel metal2 793 -2076 793 -2076 0 net=6615
rlabel metal2 1171 -2076 1171 -2076 0 net=7545
rlabel metal2 597 -2078 597 -2078 0 net=5481
rlabel metal2 835 -2078 835 -2078 0 net=5191
rlabel metal2 523 -2080 523 -2080 0 net=5113
rlabel metal2 688 -2080 688 -2080 0 net=5065
rlabel metal2 814 -2080 814 -2080 0 net=5519
rlabel metal2 926 -2080 926 -2080 0 net=6415
rlabel metal2 583 -2082 583 -2082 0 net=362
rlabel metal2 709 -2082 709 -2082 0 net=6707
rlabel metal2 380 -2084 380 -2084 0 net=4223
rlabel metal2 814 -2084 814 -2084 0 net=6792
rlabel metal2 44 -2086 44 -2086 0 net=3661
rlabel metal2 583 -2086 583 -2086 0 net=4419
rlabel metal2 919 -2086 919 -2086 0 net=6179
rlabel metal2 940 -2086 940 -2086 0 net=6929
rlabel metal2 2 -2088 2 -2088 0 net=3951
rlabel metal2 940 -2088 940 -2088 0 net=6879
rlabel metal2 44 -2090 44 -2090 0 net=1721
rlabel metal2 352 -2090 352 -2090 0 net=6151
rlabel metal2 968 -2090 968 -2090 0 net=6823
rlabel metal2 79 -2092 79 -2092 0 net=2523
rlabel metal2 275 -2094 275 -2094 0 net=1701
rlabel metal2 275 -2096 275 -2096 0 net=2163
rlabel metal2 317 -2098 317 -2098 0 net=7439
rlabel metal2 366 -2100 366 -2100 0 net=4921
rlabel metal2 702 -2102 702 -2102 0 net=3829
rlabel metal2 9 -2113 9 -2113 0 net=1722
rlabel metal2 51 -2113 51 -2113 0 net=1410
rlabel metal2 765 -2113 765 -2113 0 net=5653
rlabel metal2 793 -2113 793 -2113 0 net=6616
rlabel metal2 936 -2113 936 -2113 0 net=6506
rlabel metal2 989 -2113 989 -2113 0 net=6232
rlabel metal2 1115 -2113 1115 -2113 0 net=8090
rlabel metal2 9 -2115 9 -2115 0 net=2891
rlabel metal2 478 -2115 478 -2115 0 net=1580
rlabel metal2 695 -2115 695 -2115 0 net=5331
rlabel metal2 814 -2115 814 -2115 0 net=6032
rlabel metal2 961 -2115 961 -2115 0 net=6417
rlabel metal2 961 -2115 961 -2115 0 net=6417
rlabel metal2 968 -2115 968 -2115 0 net=7517
rlabel metal2 1118 -2115 1118 -2115 0 net=7796
rlabel metal2 1262 -2115 1262 -2115 0 net=8173
rlabel metal2 30 -2117 30 -2117 0 net=2619
rlabel metal2 51 -2117 51 -2117 0 net=4681
rlabel metal2 667 -2117 667 -2117 0 net=4941
rlabel metal2 765 -2117 765 -2117 0 net=5521
rlabel metal2 891 -2117 891 -2117 0 net=6931
rlabel metal2 1139 -2117 1139 -2117 0 net=7770
rlabel metal2 75 -2119 75 -2119 0 net=4224
rlabel metal2 814 -2119 814 -2119 0 net=5997
rlabel metal2 905 -2119 905 -2119 0 net=6573
rlabel metal2 985 -2119 985 -2119 0 net=8313
rlabel metal2 107 -2121 107 -2121 0 net=7244
rlabel metal2 1213 -2121 1213 -2121 0 net=7955
rlabel metal2 1276 -2121 1276 -2121 0 net=8225
rlabel metal2 107 -2123 107 -2123 0 net=3987
rlabel metal2 450 -2123 450 -2123 0 net=7018
rlabel metal2 1192 -2123 1192 -2123 0 net=7805
rlabel metal2 1241 -2123 1241 -2123 0 net=8049
rlabel metal2 1290 -2123 1290 -2123 0 net=8335
rlabel metal2 40 -2125 40 -2125 0 net=7981
rlabel metal2 1297 -2125 1297 -2125 0 net=8397
rlabel metal2 110 -2127 110 -2127 0 net=2452
rlabel metal2 320 -2127 320 -2127 0 net=933
rlabel metal2 488 -2127 488 -2127 0 net=6193
rlabel metal2 989 -2127 989 -2127 0 net=6693
rlabel metal2 1045 -2127 1045 -2127 0 net=7221
rlabel metal2 1206 -2127 1206 -2127 0 net=8149
rlabel metal2 131 -2129 131 -2129 0 net=2472
rlabel metal2 170 -2129 170 -2129 0 net=1020
rlabel metal2 184 -2129 184 -2129 0 net=1084
rlabel metal2 345 -2129 345 -2129 0 net=1127
rlabel metal2 579 -2129 579 -2129 0 net=2834
rlabel metal2 695 -2129 695 -2129 0 net=4875
rlabel metal2 992 -2129 992 -2129 0 net=8378
rlabel metal2 37 -2131 37 -2131 0 net=1167
rlabel metal2 191 -2131 191 -2131 0 net=2430
rlabel metal2 821 -2131 821 -2131 0 net=5579
rlabel metal2 856 -2131 856 -2131 0 net=6529
rlabel metal2 996 -2131 996 -2131 0 net=7385
rlabel metal2 1206 -2131 1206 -2131 0 net=7905
rlabel metal2 79 -2133 79 -2133 0 net=2525
rlabel metal2 191 -2133 191 -2133 0 net=1245
rlabel metal2 331 -2133 331 -2133 0 net=4373
rlabel metal2 996 -2133 996 -2133 0 net=6741
rlabel metal2 1080 -2133 1080 -2133 0 net=7441
rlabel metal2 79 -2135 79 -2135 0 net=3555
rlabel metal2 555 -2135 555 -2135 0 net=3952
rlabel metal2 660 -2135 660 -2135 0 net=5373
rlabel metal2 849 -2135 849 -2135 0 net=5823
rlabel metal2 940 -2135 940 -2135 0 net=6881
rlabel metal2 1031 -2135 1031 -2135 0 net=6825
rlabel metal2 138 -2137 138 -2137 0 net=3893
rlabel metal2 163 -2137 163 -2137 0 net=2361
rlabel metal2 1003 -2137 1003 -2137 0 net=5193
rlabel metal2 170 -2139 170 -2139 0 net=1795
rlabel metal2 628 -2139 628 -2139 0 net=8007
rlabel metal2 205 -2141 205 -2141 0 net=1261
rlabel metal2 219 -2141 219 -2141 0 net=1318
rlabel metal2 1003 -2141 1003 -2141 0 net=6727
rlabel metal2 1038 -2141 1038 -2141 0 net=7731
rlabel metal2 205 -2143 205 -2143 0 net=2235
rlabel metal2 247 -2143 247 -2143 0 net=3157
rlabel metal2 478 -2143 478 -2143 0 net=4481
rlabel metal2 649 -2143 649 -2143 0 net=4998
rlabel metal2 884 -2143 884 -2143 0 net=6153
rlabel metal2 1094 -2143 1094 -2143 0 net=7465
rlabel metal2 247 -2145 247 -2145 0 net=1695
rlabel metal2 317 -2145 317 -2145 0 net=1299
rlabel metal2 352 -2145 352 -2145 0 net=1702
rlabel metal2 450 -2145 450 -2145 0 net=427
rlabel metal2 1129 -2145 1129 -2145 0 net=7537
rlabel metal2 5 -2147 5 -2147 0 net=2425
rlabel metal2 373 -2147 373 -2147 0 net=3621
rlabel metal2 702 -2147 702 -2147 0 net=3831
rlabel metal2 1164 -2147 1164 -2147 0 net=7691
rlabel metal2 72 -2149 72 -2149 0 net=3366
rlabel metal2 394 -2149 394 -2149 0 net=6433
rlabel metal2 1185 -2149 1185 -2149 0 net=7747
rlabel metal2 72 -2151 72 -2151 0 net=7476
rlabel metal2 254 -2151 254 -2151 0 net=2404
rlabel metal2 394 -2151 394 -2151 0 net=3756
rlabel metal2 464 -2151 464 -2151 0 net=5013
rlabel metal2 730 -2151 730 -2151 0 net=2747
rlabel metal2 1199 -2151 1199 -2151 0 net=7835
rlabel metal2 2 -2153 2 -2153 0 net=3057
rlabel metal2 261 -2153 261 -2153 0 net=2339
rlabel metal2 310 -2153 310 -2153 0 net=2029
rlabel metal2 397 -2153 397 -2153 0 net=876
rlabel metal2 464 -2153 464 -2153 0 net=2333
rlabel metal2 541 -2153 541 -2153 0 net=4601
rlabel metal2 597 -2153 597 -2153 0 net=5115
rlabel metal2 744 -2153 744 -2153 0 net=6237
rlabel metal2 1227 -2153 1227 -2153 0 net=8035
rlabel metal2 65 -2155 65 -2155 0 net=1763
rlabel metal2 261 -2155 261 -2155 0 net=2165
rlabel metal2 296 -2155 296 -2155 0 net=1773
rlabel metal2 404 -2155 404 -2155 0 net=759
rlabel metal2 702 -2155 702 -2155 0 net=4915
rlabel metal2 768 -2155 768 -2155 0 net=1
rlabel metal2 1248 -2155 1248 -2155 0 net=8119
rlabel metal2 65 -2157 65 -2157 0 net=3901
rlabel metal2 275 -2157 275 -2157 0 net=1839
rlabel metal2 453 -2157 453 -2157 0 net=4478
rlabel metal2 1269 -2157 1269 -2157 0 net=8343
rlabel metal2 86 -2159 86 -2159 0 net=3065
rlabel metal2 240 -2159 240 -2159 0 net=2085
rlabel metal2 485 -2159 485 -2159 0 net=3455
rlabel metal2 548 -2159 548 -2159 0 net=6391
rlabel metal2 1304 -2159 1304 -2159 0 net=8413
rlabel metal2 198 -2161 198 -2161 0 net=1429
rlabel metal2 240 -2161 240 -2161 0 net=1609
rlabel metal2 443 -2161 443 -2161 0 net=5855
rlabel metal2 590 -2161 590 -2161 0 net=4905
rlabel metal2 723 -2161 723 -2161 0 net=5067
rlabel metal2 772 -2161 772 -2161 0 net=5129
rlabel metal2 198 -2163 198 -2163 0 net=4799
rlabel metal2 436 -2163 436 -2163 0 net=2353
rlabel metal2 499 -2163 499 -2163 0 net=6708
rlabel metal2 128 -2165 128 -2165 0 net=7695
rlabel metal2 114 -2167 114 -2167 0 net=5145
rlabel metal2 219 -2167 219 -2167 0 net=1487
rlabel metal2 576 -2167 576 -2167 0 net=5213
rlabel metal2 807 -2167 807 -2167 0 net=7521
rlabel metal2 296 -2169 296 -2169 0 net=6269
rlabel metal2 359 -2169 359 -2169 0 net=2475
rlabel metal2 324 -2171 324 -2171 0 net=1541
rlabel metal2 415 -2171 415 -2171 0 net=4415
rlabel metal2 499 -2171 499 -2171 0 net=3219
rlabel metal2 212 -2173 212 -2173 0 net=2735
rlabel metal2 502 -2173 502 -2173 0 net=5235
rlabel metal2 212 -2175 212 -2175 0 net=3049
rlabel metal2 520 -2175 520 -2175 0 net=4803
rlabel metal2 653 -2175 653 -2175 0 net=2835
rlabel metal2 324 -2177 324 -2177 0 net=1413
rlabel metal2 492 -2177 492 -2177 0 net=6181
rlabel metal2 401 -2179 401 -2179 0 net=6129
rlabel metal2 523 -2181 523 -2181 0 net=6337
rlabel metal2 576 -2183 576 -2183 0 net=4703
rlabel metal2 716 -2183 716 -2183 0 net=4739
rlabel metal2 758 -2183 758 -2183 0 net=5163
rlabel metal2 597 -2185 597 -2185 0 net=6669
rlabel metal2 621 -2185 621 -2185 0 net=5482
rlabel metal2 506 -2187 506 -2187 0 net=1538
rlabel metal2 632 -2187 632 -2187 0 net=5221
rlabel metal2 93 -2189 93 -2189 0 net=3465
rlabel metal2 611 -2189 611 -2189 0 net=4349
rlabel metal2 751 -2189 751 -2189 0 net=5203
rlabel metal2 828 -2189 828 -2189 0 net=5685
rlabel metal2 93 -2191 93 -2191 0 net=2949
rlabel metal2 583 -2191 583 -2191 0 net=4421
rlabel metal2 786 -2191 786 -2191 0 net=6329
rlabel metal2 117 -2193 117 -2193 0 net=4639
rlabel metal2 800 -2193 800 -2193 0 net=5543
rlabel metal2 863 -2193 863 -2193 0 net=6081
rlabel metal2 1136 -2193 1136 -2193 0 net=7533
rlabel metal2 282 -2195 282 -2195 0 net=3521
rlabel metal2 534 -2195 534 -2195 0 net=3199
rlabel metal2 842 -2195 842 -2195 0 net=5747
rlabel metal2 912 -2195 912 -2195 0 net=6223
rlabel metal2 1017 -2195 1017 -2195 0 net=7671
rlabel metal2 37 -2197 37 -2197 0 net=6117
rlabel metal2 933 -2197 933 -2197 0 net=5720
rlabel metal2 380 -2199 380 -2199 0 net=3663
rlabel metal2 534 -2199 534 -2199 0 net=4839
rlabel metal2 1017 -2199 1017 -2199 0 net=7183
rlabel metal2 1108 -2199 1108 -2199 0 net=7507
rlabel metal2 135 -2201 135 -2201 0 net=2533
rlabel metal2 520 -2201 520 -2201 0 net=7279
rlabel metal2 135 -2203 135 -2203 0 net=4922
rlabel metal2 569 -2203 569 -2203 0 net=3945
rlabel metal2 16 -2205 16 -2205 0 net=2503
rlabel metal2 562 -2205 562 -2205 0 net=6546
rlabel metal2 16 -2207 16 -2207 0 net=2805
rlabel metal2 562 -2207 562 -2207 0 net=4267
rlabel metal2 58 -2209 58 -2209 0 net=2967
rlabel metal2 604 -2209 604 -2209 0 net=4687
rlabel metal2 58 -2211 58 -2211 0 net=2565
rlabel metal2 152 -2211 152 -2211 0 net=7597
rlabel metal2 100 -2213 100 -2213 0 net=2280
rlabel metal2 100 -2215 100 -2215 0 net=2059
rlabel metal2 121 -2217 121 -2217 0 net=2709
rlabel metal2 289 -2217 289 -2217 0 net=2611
rlabel metal2 23 -2219 23 -2219 0 net=4493
rlabel metal2 23 -2221 23 -2221 0 net=387
rlabel metal2 121 -2221 121 -2221 0 net=2049
rlabel metal2 408 -2223 408 -2223 0 net=7106
rlabel metal2 1066 -2225 1066 -2225 0 net=7295
rlabel metal2 1101 -2227 1101 -2227 0 net=7489
rlabel metal2 1143 -2229 1143 -2229 0 net=7547
rlabel metal2 1073 -2231 1073 -2231 0 net=7129
rlabel metal2 870 -2233 870 -2233 0 net=7309
rlabel metal2 870 -2235 870 -2235 0 net=7257
rlabel metal2 5 -2246 5 -2246 0 net=2620
rlabel metal2 61 -2246 61 -2246 0 net=6182
rlabel metal2 516 -2246 516 -2246 0 net=108
rlabel metal2 747 -2246 747 -2246 0 net=7386
rlabel metal2 23 -2248 23 -2248 0 net=6130
rlabel metal2 1034 -2248 1034 -2248 0 net=8336
rlabel metal2 23 -2250 23 -2250 0 net=5207
rlabel metal2 408 -2250 408 -2250 0 net=2736
rlabel metal2 425 -2250 425 -2250 0 net=4350
rlabel metal2 761 -2250 761 -2250 0 net=3832
rlabel metal2 870 -2250 870 -2250 0 net=8008
rlabel metal2 33 -2252 33 -2252 0 net=4800
rlabel metal2 205 -2252 205 -2252 0 net=2236
rlabel metal2 387 -2252 387 -2252 0 net=1542
rlabel metal2 527 -2252 527 -2252 0 net=5116
rlabel metal2 810 -2252 810 -2252 0 net=6418
rlabel metal2 982 -2252 982 -2252 0 net=8226
rlabel metal2 9 -2254 9 -2254 0 net=2893
rlabel metal2 205 -2254 205 -2254 0 net=2031
rlabel metal2 387 -2254 387 -2254 0 net=5693
rlabel metal2 520 -2254 520 -2254 0 net=4268
rlabel metal2 579 -2254 579 -2254 0 net=6434
rlabel metal2 982 -2254 982 -2254 0 net=6187
rlabel metal2 1024 -2254 1024 -2254 0 net=7467
rlabel metal2 9 -2256 9 -2256 0 net=2477
rlabel metal2 411 -2256 411 -2256 0 net=2334
rlabel metal2 527 -2256 527 -2256 0 net=1783
rlabel metal2 961 -2256 961 -2256 0 net=7185
rlabel metal2 1094 -2256 1094 -2256 0 net=7599
rlabel metal2 37 -2258 37 -2258 0 net=4374
rlabel metal2 1017 -2258 1017 -2258 0 net=7443
rlabel metal2 1150 -2258 1150 -2258 0 net=7983
rlabel metal2 37 -2260 37 -2260 0 net=271
rlabel metal2 359 -2260 359 -2260 0 net=3457
rlabel metal2 530 -2260 530 -2260 0 net=5222
rlabel metal2 933 -2260 933 -2260 0 net=7281
rlabel metal2 1080 -2260 1080 -2260 0 net=8399
rlabel metal2 40 -2262 40 -2262 0 net=2426
rlabel metal2 464 -2262 464 -2262 0 net=5825
rlabel metal2 856 -2262 856 -2262 0 net=6883
rlabel metal2 1059 -2262 1059 -2262 0 net=7523
rlabel metal2 40 -2264 40 -2264 0 net=6919
rlabel metal2 975 -2264 975 -2264 0 net=8345
rlabel metal2 44 -2266 44 -2266 0 net=2535
rlabel metal2 485 -2266 485 -2266 0 net=3665
rlabel metal2 548 -2266 548 -2266 0 net=5857
rlabel metal2 695 -2266 695 -2266 0 net=4876
rlabel metal2 870 -2266 870 -2266 0 net=6339
rlabel metal2 1122 -2266 1122 -2266 0 net=7807
rlabel metal2 79 -2268 79 -2268 0 net=3557
rlabel metal2 548 -2268 548 -2268 0 net=4689
rlabel metal2 625 -2268 625 -2268 0 net=4805
rlabel metal2 674 -2268 674 -2268 0 net=5215
rlabel metal2 873 -2268 873 -2268 0 net=6826
rlabel metal2 1192 -2268 1192 -2268 0 net=8051
rlabel metal2 16 -2270 16 -2270 0 net=2807
rlabel metal2 86 -2270 86 -2270 0 net=3066
rlabel metal2 306 -2270 306 -2270 0 net=5357
rlabel metal2 492 -2270 492 -2270 0 net=2603
rlabel metal2 1129 -2270 1129 -2270 0 net=7539
rlabel metal2 16 -2272 16 -2272 0 net=1301
rlabel metal2 320 -2272 320 -2272 0 net=7227
rlabel metal2 86 -2274 86 -2274 0 net=5069
rlabel metal2 737 -2274 737 -2274 0 net=6239
rlabel metal2 772 -2274 772 -2274 0 net=5545
rlabel metal2 96 -2276 96 -2276 0 net=296
rlabel metal2 628 -2276 628 -2276 0 net=6865
rlabel metal2 100 -2278 100 -2278 0 net=2060
rlabel metal2 117 -2278 117 -2278 0 net=7696
rlabel metal2 100 -2280 100 -2280 0 net=1129
rlabel metal2 352 -2280 352 -2280 0 net=4483
rlabel metal2 513 -2280 513 -2280 0 net=7771
rlabel metal2 1178 -2280 1178 -2280 0 net=8151
rlabel metal2 114 -2282 114 -2282 0 net=1247
rlabel metal2 240 -2282 240 -2282 0 net=1611
rlabel metal2 558 -2282 558 -2282 0 net=3622
rlabel metal2 695 -2282 695 -2282 0 net=5333
rlabel metal2 800 -2282 800 -2282 0 net=5999
rlabel metal2 121 -2284 121 -2284 0 net=2050
rlabel metal2 793 -2284 793 -2284 0 net=5915
rlabel metal2 814 -2284 814 -2284 0 net=6119
rlabel metal2 121 -2286 121 -2286 0 net=2785
rlabel metal2 555 -2286 555 -2286 0 net=6387
rlabel metal2 877 -2286 877 -2286 0 net=6393
rlabel metal2 149 -2288 149 -2288 0 net=5130
rlabel metal2 947 -2288 947 -2288 0 net=7223
rlabel metal2 149 -2290 149 -2290 0 net=4416
rlabel metal2 450 -2290 450 -2290 0 net=3201
rlabel metal2 593 -2290 593 -2290 0 net=5654
rlabel metal2 919 -2290 919 -2290 0 net=6695
rlabel metal2 1045 -2290 1045 -2290 0 net=8415
rlabel metal2 152 -2292 152 -2292 0 net=559
rlabel metal2 989 -2292 989 -2292 0 net=7297
rlabel metal2 156 -2294 156 -2294 0 net=3895
rlabel metal2 331 -2294 331 -2294 0 net=6271
rlabel metal2 1066 -2294 1066 -2294 0 net=7693
rlabel metal2 2 -2296 2 -2296 0 net=3059
rlabel metal2 341 -2296 341 -2296 0 net=2968
rlabel metal2 562 -2296 562 -2296 0 net=5375
rlabel metal2 677 -2296 677 -2296 0 net=7534
rlabel metal2 2 -2298 2 -2298 0 net=5281
rlabel metal2 569 -2298 569 -2298 0 net=3947
rlabel metal2 604 -2298 604 -2298 0 net=4917
rlabel metal2 786 -2298 786 -2298 0 net=6331
rlabel metal2 107 -2300 107 -2300 0 net=3989
rlabel metal2 471 -2300 471 -2300 0 net=3159
rlabel metal2 611 -2300 611 -2300 0 net=4423
rlabel metal2 635 -2300 635 -2300 0 net=5164
rlabel metal2 807 -2300 807 -2300 0 net=6728
rlabel metal2 107 -2302 107 -2302 0 net=5147
rlabel metal2 156 -2302 156 -2302 0 net=1169
rlabel metal2 191 -2302 191 -2302 0 net=2613
rlabel metal2 380 -2302 380 -2302 0 net=4705
rlabel metal2 611 -2302 611 -2302 0 net=4641
rlabel metal2 639 -2302 639 -2302 0 net=5015
rlabel metal2 758 -2302 758 -2302 0 net=7130
rlabel metal2 75 -2304 75 -2304 0 net=28
rlabel metal2 646 -2304 646 -2304 0 net=7305
rlabel metal2 128 -2306 128 -2306 0 net=1441
rlabel metal2 471 -2306 471 -2306 0 net=3467
rlabel metal2 576 -2306 576 -2306 0 net=1251
rlabel metal2 51 -2308 51 -2308 0 net=4682
rlabel metal2 499 -2308 499 -2308 0 net=3221
rlabel metal2 597 -2308 597 -2308 0 net=6671
rlabel metal2 660 -2308 660 -2308 0 net=8314
rlabel metal2 51 -2310 51 -2310 0 net=488
rlabel metal2 163 -2310 163 -2310 0 net=2363
rlabel metal2 338 -2310 338 -2310 0 net=7999
rlabel metal2 138 -2312 138 -2312 0 net=7571
rlabel metal2 163 -2314 163 -2314 0 net=2589
rlabel metal2 499 -2314 499 -2314 0 net=4841
rlabel metal2 590 -2314 590 -2314 0 net=4907
rlabel metal2 702 -2314 702 -2314 0 net=5205
rlabel metal2 1003 -2314 1003 -2314 0 net=7907
rlabel metal2 177 -2316 177 -2316 0 net=2527
rlabel metal2 534 -2316 534 -2316 0 net=6083
rlabel metal2 1206 -2316 1206 -2316 0 net=8121
rlabel metal2 170 -2318 170 -2318 0 net=1797
rlabel metal2 184 -2318 184 -2318 0 net=1263
rlabel metal2 254 -2318 254 -2318 0 net=1765
rlabel metal2 590 -2318 590 -2318 0 net=7881
rlabel metal2 1248 -2318 1248 -2318 0 net=5195
rlabel metal2 93 -2320 93 -2320 0 net=2951
rlabel metal2 261 -2320 261 -2320 0 net=2167
rlabel metal2 709 -2320 709 -2320 0 net=4741
rlabel metal2 751 -2320 751 -2320 0 net=5749
rlabel metal2 863 -2320 863 -2320 0 net=6531
rlabel metal2 65 -2322 65 -2322 0 net=3902
rlabel metal2 170 -2322 170 -2322 0 net=5767
rlabel metal2 397 -2322 397 -2322 0 net=6297
rlabel metal2 954 -2322 954 -2322 0 net=7509
rlabel metal2 30 -2324 30 -2324 0 net=5911
rlabel metal2 219 -2324 219 -2324 0 net=1489
rlabel metal2 261 -2324 261 -2324 0 net=4897
rlabel metal2 716 -2324 716 -2324 0 net=5523
rlabel metal2 1108 -2324 1108 -2324 0 net=7749
rlabel metal2 30 -2326 30 -2326 0 net=5131
rlabel metal2 1185 -2326 1185 -2326 0 net=8037
rlabel metal2 135 -2328 135 -2328 0 net=5797
rlabel metal2 891 -2328 891 -2328 0 net=6933
rlabel metal2 135 -2330 135 -2330 0 net=2504
rlabel metal2 397 -2330 397 -2330 0 net=2748
rlabel metal2 891 -2330 891 -2330 0 net=6743
rlabel metal2 219 -2332 219 -2332 0 net=1415
rlabel metal2 366 -2332 366 -2332 0 net=4603
rlabel metal2 730 -2332 730 -2332 0 net=5581
rlabel metal2 996 -2332 996 -2332 0 net=7311
rlabel metal2 226 -2334 226 -2334 0 net=1431
rlabel metal2 821 -2334 821 -2334 0 net=6155
rlabel metal2 1073 -2334 1073 -2334 0 net=7549
rlabel metal2 142 -2336 142 -2336 0 net=2711
rlabel metal2 233 -2336 233 -2336 0 net=2341
rlabel metal2 282 -2336 282 -2336 0 net=3522
rlabel metal2 779 -2336 779 -2336 0 net=5237
rlabel metal2 1143 -2336 1143 -2336 0 net=7837
rlabel metal2 142 -2338 142 -2338 0 net=5687
rlabel metal2 268 -2340 268 -2340 0 net=1775
rlabel metal2 324 -2340 324 -2340 0 net=2355
rlabel metal2 541 -2340 541 -2340 0 net=2837
rlabel metal2 779 -2340 779 -2340 0 net=6225
rlabel metal2 275 -2342 275 -2342 0 net=1841
rlabel metal2 443 -2342 443 -2342 0 net=4787
rlabel metal2 621 -2342 621 -2342 0 net=8101
rlabel metal2 275 -2344 275 -2344 0 net=4495
rlabel metal2 653 -2344 653 -2344 0 net=4943
rlabel metal2 828 -2344 828 -2344 0 net=6195
rlabel metal2 912 -2344 912 -2344 0 net=7259
rlabel metal2 72 -2346 72 -2346 0 net=7511
rlabel metal2 898 -2346 898 -2346 0 net=6575
rlabel metal2 72 -2348 72 -2348 0 net=1697
rlabel metal2 282 -2348 282 -2348 0 net=5209
rlabel metal2 436 -2348 436 -2348 0 net=7525
rlabel metal2 58 -2350 58 -2350 0 net=2567
rlabel metal2 905 -2350 905 -2350 0 net=7519
rlabel metal2 58 -2352 58 -2352 0 net=7415
rlabel metal2 1038 -2352 1038 -2352 0 net=7733
rlabel metal2 212 -2354 212 -2354 0 net=3051
rlabel metal2 1038 -2354 1038 -2354 0 net=7491
rlabel metal2 212 -2356 212 -2356 0 net=2087
rlabel metal2 1101 -2356 1101 -2356 0 net=7673
rlabel metal2 1157 -2358 1157 -2358 0 net=7957
rlabel metal2 1213 -2360 1213 -2360 0 net=8175
rlabel metal2 9 -2371 9 -2371 0 net=2478
rlabel metal2 394 -2371 394 -2371 0 net=7228
rlabel metal2 23 -2373 23 -2373 0 net=5208
rlabel metal2 352 -2373 352 -2373 0 net=4484
rlabel metal2 446 -2373 446 -2373 0 net=6226
rlabel metal2 796 -2373 796 -2373 0 net=7510
rlabel metal2 1031 -2373 1031 -2373 0 net=7551
rlabel metal2 1104 -2373 1104 -2373 0 net=7734
rlabel metal2 30 -2375 30 -2375 0 net=5132
rlabel metal2 303 -2375 303 -2375 0 net=6298
rlabel metal2 849 -2375 849 -2375 0 net=6696
rlabel metal2 954 -2375 954 -2375 0 net=8417
rlabel metal2 1073 -2375 1073 -2375 0 net=8103
rlabel metal2 37 -2377 37 -2377 0 net=3896
rlabel metal2 303 -2377 303 -2377 0 net=6033
rlabel metal2 464 -2377 464 -2377 0 net=5826
rlabel metal2 779 -2377 779 -2377 0 net=7417
rlabel metal2 1034 -2377 1034 -2377 0 net=8152
rlabel metal2 40 -2379 40 -2379 0 net=6272
rlabel metal2 1010 -2379 1010 -2379 0 net=7524
rlabel metal2 54 -2381 54 -2381 0 net=2952
rlabel metal2 310 -2381 310 -2381 0 net=1843
rlabel metal2 310 -2381 310 -2381 0 net=1843
rlabel metal2 320 -2381 320 -2381 0 net=1432
rlabel metal2 807 -2381 807 -2381 0 net=7838
rlabel metal2 61 -2383 61 -2383 0 net=3160
rlabel metal2 576 -2383 576 -2383 0 net=7520
rlabel metal2 908 -2383 908 -2383 0 net=1252
rlabel metal2 65 -2385 65 -2385 0 net=5913
rlabel metal2 65 -2385 65 -2385 0 net=5913
rlabel metal2 72 -2385 72 -2385 0 net=1698
rlabel metal2 520 -2385 520 -2385 0 net=1612
rlabel metal2 842 -2385 842 -2385 0 net=7751
rlabel metal2 72 -2387 72 -2387 0 net=5769
rlabel metal2 184 -2387 184 -2387 0 net=1264
rlabel metal2 338 -2387 338 -2387 0 net=4789
rlabel metal2 485 -2387 485 -2387 0 net=3667
rlabel metal2 898 -2387 898 -2387 0 net=6576
rlabel metal2 1059 -2387 1059 -2387 0 net=8401
rlabel metal2 79 -2389 79 -2389 0 net=2809
rlabel metal2 163 -2389 163 -2389 0 net=2591
rlabel metal2 359 -2389 359 -2389 0 net=3459
rlabel metal2 366 -2389 366 -2389 0 net=4604
rlabel metal2 520 -2389 520 -2389 0 net=3729
rlabel metal2 614 -2389 614 -2389 0 net=6532
rlabel metal2 898 -2389 898 -2389 0 net=7959
rlabel metal2 44 -2391 44 -2391 0 net=2537
rlabel metal2 86 -2391 86 -2391 0 net=5071
rlabel metal2 394 -2391 394 -2391 0 net=3469
rlabel metal2 516 -2391 516 -2391 0 net=7306
rlabel metal2 86 -2393 86 -2393 0 net=5211
rlabel metal2 359 -2393 359 -2393 0 net=5359
rlabel metal2 422 -2393 422 -2393 0 net=5858
rlabel metal2 723 -2393 723 -2393 0 net=5546
rlabel metal2 786 -2393 786 -2393 0 net=7101
rlabel metal2 905 -2393 905 -2393 0 net=7540
rlabel metal2 93 -2395 93 -2395 0 net=6863
rlabel metal2 450 -2395 450 -2395 0 net=3203
rlabel metal2 919 -2395 919 -2395 0 net=7313
rlabel metal2 1080 -2395 1080 -2395 0 net=7883
rlabel metal2 93 -2397 93 -2397 0 net=3395
rlabel metal2 450 -2397 450 -2397 0 net=6341
rlabel metal2 884 -2397 884 -2397 0 net=5239
rlabel metal2 100 -2399 100 -2399 0 net=1130
rlabel metal2 751 -2399 751 -2399 0 net=5751
rlabel metal2 765 -2399 765 -2399 0 net=5799
rlabel metal2 870 -2399 870 -2399 0 net=7261
rlabel metal2 940 -2399 940 -2399 0 net=7808
rlabel metal2 100 -2401 100 -2401 0 net=5689
rlabel metal2 184 -2401 184 -2401 0 net=5377
rlabel metal2 569 -2401 569 -2401 0 net=4806
rlabel metal2 635 -2401 635 -2401 0 net=5206
rlabel metal2 709 -2401 709 -2401 0 net=4743
rlabel metal2 912 -2401 912 -2401 0 net=8001
rlabel metal2 107 -2403 107 -2403 0 net=5148
rlabel metal2 198 -2403 198 -2403 0 net=2894
rlabel metal2 457 -2403 457 -2403 0 net=3991
rlabel metal2 548 -2403 548 -2403 0 net=4691
rlabel metal2 590 -2403 590 -2403 0 net=4944
rlabel metal2 660 -2403 660 -2403 0 net=6934
rlabel metal2 107 -2405 107 -2405 0 net=4909
rlabel metal2 611 -2405 611 -2405 0 net=4643
rlabel metal2 663 -2405 663 -2405 0 net=7694
rlabel metal2 58 -2407 58 -2407 0 net=4923
rlabel metal2 646 -2407 646 -2407 0 net=6673
rlabel metal2 751 -2407 751 -2407 0 net=6745
rlabel metal2 961 -2407 961 -2407 0 net=7187
rlabel metal2 58 -2409 58 -2409 0 net=2569
rlabel metal2 261 -2409 261 -2409 0 net=4899
rlabel metal2 646 -2409 646 -2409 0 net=7283
rlabel metal2 1066 -2409 1066 -2409 0 net=7773
rlabel metal2 114 -2411 114 -2411 0 net=1249
rlabel metal2 114 -2411 114 -2411 0 net=1249
rlabel metal2 121 -2411 121 -2411 0 net=2787
rlabel metal2 261 -2411 261 -2411 0 net=3223
rlabel metal2 555 -2411 555 -2411 0 net=5583
rlabel metal2 765 -2411 765 -2411 0 net=8347
rlabel metal2 1129 -2411 1129 -2411 0 net=5197
rlabel metal2 124 -2413 124 -2413 0 net=6866
rlabel metal2 128 -2415 128 -2415 0 net=1442
rlabel metal2 198 -2415 198 -2415 0 net=2712
rlabel metal2 247 -2415 247 -2415 0 net=2357
rlabel metal2 415 -2415 415 -2415 0 net=3558
rlabel metal2 667 -2415 667 -2415 0 net=7513
rlabel metal2 709 -2415 709 -2415 0 net=7299
rlabel metal2 128 -2417 128 -2417 0 net=944
rlabel metal2 142 -2417 142 -2417 0 net=7447
rlabel metal2 387 -2417 387 -2417 0 net=5695
rlabel metal2 667 -2417 667 -2417 0 net=6197
rlabel metal2 877 -2417 877 -2417 0 net=6395
rlabel metal2 989 -2417 989 -2417 0 net=8053
rlabel metal2 131 -2419 131 -2419 0 net=6183
rlabel metal2 558 -2419 558 -2419 0 net=5016
rlabel metal2 674 -2419 674 -2419 0 net=5217
rlabel metal2 1192 -2419 1192 -2419 0 net=8123
rlabel metal2 135 -2421 135 -2421 0 net=5859
rlabel metal2 135 -2421 135 -2421 0 net=5859
rlabel metal2 226 -2421 226 -2421 0 net=3061
rlabel metal2 380 -2421 380 -2421 0 net=4706
rlabel metal2 681 -2421 681 -2421 0 net=6388
rlabel metal2 726 -2421 726 -2421 0 net=1313
rlabel metal2 51 -2423 51 -2423 0 net=6585
rlabel metal2 387 -2423 387 -2423 0 net=3053
rlabel metal2 439 -2423 439 -2423 0 net=662
rlabel metal2 772 -2423 772 -2423 0 net=6885
rlabel metal2 877 -2423 877 -2423 0 net=7445
rlabel metal2 275 -2425 275 -2425 0 net=4496
rlabel metal2 814 -2425 814 -2425 0 net=6121
rlabel metal2 1017 -2425 1017 -2425 0 net=8177
rlabel metal2 212 -2427 212 -2427 0 net=2089
rlabel metal2 282 -2427 282 -2427 0 net=2169
rlabel metal2 415 -2427 415 -2427 0 net=1921
rlabel metal2 471 -2427 471 -2427 0 net=4919
rlabel metal2 611 -2427 611 -2427 0 net=3747
rlabel metal2 212 -2429 212 -2429 0 net=1491
rlabel metal2 289 -2429 289 -2429 0 net=2365
rlabel metal2 331 -2429 331 -2429 0 net=1767
rlabel metal2 401 -2429 401 -2429 0 net=3161
rlabel metal2 579 -2429 579 -2429 0 net=1881
rlabel metal2 814 -2429 814 -2429 0 net=7601
rlabel metal2 177 -2431 177 -2431 0 net=1799
rlabel metal2 289 -2431 289 -2431 0 net=3897
rlabel metal2 373 -2431 373 -2431 0 net=931
rlabel metal2 856 -2431 856 -2431 0 net=7493
rlabel metal2 156 -2433 156 -2433 0 net=1171
rlabel metal2 317 -2433 317 -2433 0 net=2529
rlabel metal2 429 -2433 429 -2433 0 net=6085
rlabel metal2 604 -2433 604 -2433 0 net=7573
rlabel metal2 156 -2435 156 -2435 0 net=2343
rlabel metal2 345 -2435 345 -2435 0 net=2189
rlabel metal2 478 -2435 478 -2435 0 net=5282
rlabel metal2 618 -2435 618 -2435 0 net=4425
rlabel metal2 688 -2435 688 -2435 0 net=6921
rlabel metal2 982 -2435 982 -2435 0 net=6189
rlabel metal2 233 -2437 233 -2437 0 net=1785
rlabel metal2 534 -2437 534 -2437 0 net=7159
rlabel metal2 639 -2437 639 -2437 0 net=6241
rlabel metal2 926 -2437 926 -2437 0 net=7909
rlabel metal2 457 -2439 457 -2439 0 net=2605
rlabel metal2 499 -2439 499 -2439 0 net=4843
rlabel metal2 527 -2439 527 -2439 0 net=5335
rlabel metal2 737 -2439 737 -2439 0 net=6551
rlabel metal2 982 -2439 982 -2439 0 net=7675
rlabel metal2 478 -2441 478 -2441 0 net=3949
rlabel metal2 618 -2441 618 -2441 0 net=5525
rlabel metal2 821 -2441 821 -2441 0 net=6157
rlabel metal2 1094 -2441 1094 -2441 0 net=2175
rlabel metal2 268 -2443 268 -2443 0 net=1777
rlabel metal2 632 -2443 632 -2443 0 net=6001
rlabel metal2 821 -2443 821 -2443 0 net=7527
rlabel metal2 205 -2445 205 -2445 0 net=2033
rlabel metal2 492 -2445 492 -2445 0 net=5917
rlabel metal2 205 -2447 205 -2447 0 net=1417
rlabel metal2 499 -2447 499 -2447 0 net=8249
rlabel metal2 695 -2447 695 -2447 0 net=7984
rlabel metal2 191 -2449 191 -2449 0 net=2615
rlabel metal2 541 -2449 541 -2449 0 net=2839
rlabel metal2 16 -2451 16 -2451 0 net=1303
rlabel metal2 443 -2451 443 -2451 0 net=3889
rlabel metal2 716 -2451 716 -2451 0 net=6333
rlabel metal2 835 -2453 835 -2453 0 net=7469
rlabel metal2 947 -2455 947 -2455 0 net=7225
rlabel metal2 947 -2457 947 -2457 0 net=8039
rlabel metal2 58 -2468 58 -2468 0 net=2570
rlabel metal2 471 -2468 471 -2468 0 net=4920
rlabel metal2 530 -2468 530 -2468 0 net=1778
rlabel metal2 625 -2468 625 -2468 0 net=5696
rlabel metal2 961 -2468 961 -2468 0 net=1314
rlabel metal2 1108 -2468 1108 -2468 0 net=7189
rlabel metal2 1185 -2468 1185 -2468 0 net=8125
rlabel metal2 65 -2470 65 -2470 0 net=5914
rlabel metal2 366 -2470 366 -2470 0 net=5072
rlabel metal2 625 -2470 625 -2470 0 net=7529
rlabel metal2 828 -2470 828 -2470 0 net=7262
rlabel metal2 1013 -2470 1013 -2470 0 net=5198
rlabel metal2 72 -2472 72 -2472 0 net=5770
rlabel metal2 135 -2472 135 -2472 0 net=5861
rlabel metal2 135 -2472 135 -2472 0 net=5861
rlabel metal2 149 -2472 149 -2472 0 net=2811
rlabel metal2 366 -2472 366 -2472 0 net=7574
rlabel metal2 639 -2472 639 -2472 0 net=6243
rlabel metal2 674 -2472 674 -2472 0 net=5752
rlabel metal2 793 -2472 793 -2472 0 net=5800
rlabel metal2 828 -2472 828 -2472 0 net=7495
rlabel metal2 863 -2472 863 -2472 0 net=3205
rlabel metal2 1024 -2472 1024 -2472 0 net=7226
rlabel metal2 79 -2474 79 -2474 0 net=2538
rlabel metal2 478 -2474 478 -2474 0 net=3950
rlabel metal2 723 -2474 723 -2474 0 net=8040
rlabel metal2 1038 -2474 1038 -2474 0 net=8105
rlabel metal2 1087 -2474 1087 -2474 0 net=6190
rlabel metal2 86 -2476 86 -2476 0 net=5212
rlabel metal2 191 -2476 191 -2476 0 net=1304
rlabel metal2 740 -2476 740 -2476 0 net=7446
rlabel metal2 926 -2476 926 -2476 0 net=7911
rlabel metal2 1052 -2476 1052 -2476 0 net=8403
rlabel metal2 1094 -2476 1094 -2476 0 net=2176
rlabel metal2 1094 -2476 1094 -2476 0 net=2176
rlabel metal2 107 -2478 107 -2478 0 net=4910
rlabel metal2 492 -2478 492 -2478 0 net=5919
rlabel metal2 618 -2478 618 -2478 0 net=5527
rlabel metal2 758 -2478 758 -2478 0 net=7753
rlabel metal2 863 -2478 863 -2478 0 net=7676
rlabel metal2 124 -2480 124 -2480 0 net=3062
rlabel metal2 247 -2480 247 -2480 0 net=2359
rlabel metal2 499 -2480 499 -2480 0 net=8250
rlabel metal2 639 -2480 639 -2480 0 net=7103
rlabel metal2 800 -2480 800 -2480 0 net=2840
rlabel metal2 926 -2480 926 -2480 0 net=5241
rlabel metal2 173 -2482 173 -2482 0 net=2217
rlabel metal2 254 -2482 254 -2482 0 net=2789
rlabel metal2 254 -2482 254 -2482 0 net=2789
rlabel metal2 278 -2482 278 -2482 0 net=5360
rlabel metal2 373 -2482 373 -2482 0 net=575
rlabel metal2 446 -2482 446 -2482 0 net=3668
rlabel metal2 201 -2484 201 -2484 0 net=6087
rlabel metal2 282 -2484 282 -2484 0 net=2171
rlabel metal2 499 -2484 499 -2484 0 net=6675
rlabel metal2 772 -2484 772 -2484 0 net=6887
rlabel metal2 800 -2484 800 -2484 0 net=8003
rlabel metal2 212 -2486 212 -2486 0 net=1492
rlabel metal2 565 -2486 565 -2486 0 net=5218
rlabel metal2 219 -2488 219 -2488 0 net=2616
rlabel metal2 359 -2488 359 -2488 0 net=2763
rlabel metal2 380 -2488 380 -2488 0 net=6586
rlabel metal2 730 -2488 730 -2488 0 net=1883
rlabel metal2 807 -2488 807 -2488 0 net=8054
rlabel metal2 205 -2490 205 -2490 0 net=1419
rlabel metal2 390 -2490 390 -2490 0 net=25
rlabel metal2 520 -2490 520 -2490 0 net=3731
rlabel metal2 730 -2490 730 -2490 0 net=6747
rlabel metal2 772 -2490 772 -2490 0 net=7471
rlabel metal2 912 -2490 912 -2490 0 net=8419
rlabel metal2 975 -2490 975 -2490 0 net=6159
rlabel metal2 93 -2492 93 -2492 0 net=3396
rlabel metal2 544 -2492 544 -2492 0 net=605
rlabel metal2 597 -2492 597 -2492 0 net=4924
rlabel metal2 954 -2492 954 -2492 0 net=8179
rlabel metal2 114 -2494 114 -2494 0 net=1250
rlabel metal2 597 -2494 597 -2494 0 net=6553
rlabel metal2 1017 -2494 1017 -2494 0 net=7553
rlabel metal2 282 -2496 282 -2496 0 net=2191
rlabel metal2 373 -2496 373 -2496 0 net=7161
rlabel metal2 548 -2496 548 -2496 0 net=6184
rlabel metal2 1031 -2496 1031 -2496 0 net=7775
rlabel metal2 289 -2498 289 -2498 0 net=3898
rlabel metal2 646 -2498 646 -2498 0 net=7285
rlabel metal2 1066 -2498 1066 -2498 0 net=7885
rlabel metal2 233 -2500 233 -2500 0 net=1787
rlabel metal2 296 -2500 296 -2500 0 net=2592
rlabel metal2 170 -2502 170 -2502 0 net=8095
rlabel metal2 296 -2502 296 -2502 0 net=6035
rlabel metal2 317 -2502 317 -2502 0 net=2530
rlabel metal2 443 -2502 443 -2502 0 net=5585
rlabel metal2 569 -2502 569 -2502 0 net=7418
rlabel metal2 100 -2504 100 -2504 0 net=5691
rlabel metal2 327 -2504 327 -2504 0 net=3162
rlabel metal2 415 -2504 415 -2504 0 net=1923
rlabel metal2 541 -2504 541 -2504 0 net=3891
rlabel metal2 653 -2504 653 -2504 0 net=4644
rlabel metal2 240 -2506 240 -2506 0 net=1801
rlabel metal2 422 -2506 422 -2506 0 net=6864
rlabel metal2 653 -2506 653 -2506 0 net=7515
rlabel metal2 275 -2508 275 -2508 0 net=2091
rlabel metal2 331 -2508 331 -2508 0 net=1769
rlabel metal2 509 -2508 509 -2508 0 net=3748
rlabel metal2 128 -2510 128 -2510 0 net=3637
rlabel metal2 338 -2510 338 -2510 0 net=4791
rlabel metal2 338 -2510 338 -2510 0 net=4791
rlabel metal2 345 -2510 345 -2510 0 net=3993
rlabel metal2 513 -2510 513 -2510 0 net=7301
rlabel metal2 121 -2512 121 -2512 0 net=6095
rlabel metal2 310 -2512 310 -2512 0 net=1845
rlabel metal2 429 -2512 429 -2512 0 net=6086
rlabel metal2 667 -2512 667 -2512 0 net=6199
rlabel metal2 702 -2512 702 -2512 0 net=6335
rlabel metal2 184 -2514 184 -2514 0 net=5379
rlabel metal2 408 -2514 408 -2514 0 net=3461
rlabel metal2 436 -2514 436 -2514 0 net=13
rlabel metal2 268 -2516 268 -2516 0 net=2035
rlabel metal2 450 -2516 450 -2516 0 net=6342
rlabel metal2 485 -2516 485 -2516 0 net=7602
rlabel metal2 142 -2518 142 -2518 0 net=7449
rlabel metal2 387 -2518 387 -2518 0 net=3055
rlabel metal2 527 -2518 527 -2518 0 net=5337
rlabel metal2 177 -2520 177 -2520 0 net=1173
rlabel metal2 548 -2520 548 -2520 0 net=7314
rlabel metal2 387 -2522 387 -2522 0 net=3470
rlabel metal2 555 -2522 555 -2522 0 net=6923
rlabel metal2 324 -2524 324 -2524 0 net=2367
rlabel metal2 569 -2524 569 -2524 0 net=4426
rlabel metal2 576 -2526 576 -2526 0 net=4693
rlabel metal2 681 -2526 681 -2526 0 net=6396
rlabel metal2 457 -2528 457 -2528 0 net=2607
rlabel metal2 590 -2528 590 -2528 0 net=4901
rlabel metal2 884 -2528 884 -2528 0 net=4745
rlabel metal2 422 -2530 422 -2530 0 net=2061
rlabel metal2 590 -2530 590 -2530 0 net=6122
rlabel metal2 632 -2532 632 -2532 0 net=6003
rlabel metal2 562 -2534 562 -2534 0 net=4281
rlabel metal2 660 -2534 660 -2534 0 net=8349
rlabel metal2 506 -2536 506 -2536 0 net=4845
rlabel metal2 765 -2536 765 -2536 0 net=7961
rlabel metal2 261 -2538 261 -2538 0 net=3224
rlabel metal2 156 -2540 156 -2540 0 net=2345
rlabel metal2 131 -2551 131 -2551 0 net=5862
rlabel metal2 226 -2551 226 -2551 0 net=6088
rlabel metal2 261 -2551 261 -2551 0 net=2346
rlabel metal2 380 -2551 380 -2551 0 net=1420
rlabel metal2 530 -2551 530 -2551 0 net=6336
rlabel metal2 716 -2551 716 -2551 0 net=6004
rlabel metal2 814 -2551 814 -2551 0 net=7497
rlabel metal2 866 -2551 866 -2551 0 net=5242
rlabel metal2 933 -2551 933 -2551 0 net=4746
rlabel metal2 968 -2551 968 -2551 0 net=6161
rlabel metal2 1013 -2551 1013 -2551 0 net=8106
rlabel metal2 1045 -2551 1045 -2551 0 net=8405
rlabel metal2 1059 -2551 1059 -2551 0 net=7887
rlabel metal2 1143 -2551 1143 -2551 0 net=7190
rlabel metal2 1181 -2551 1181 -2551 0 net=8126
rlabel metal2 128 -2553 128 -2553 0 net=6097
rlabel metal2 233 -2553 233 -2553 0 net=8096
rlabel metal2 282 -2553 282 -2553 0 net=2192
rlabel metal2 394 -2553 394 -2553 0 net=2369
rlabel metal2 478 -2553 478 -2553 0 net=2172
rlabel metal2 681 -2553 681 -2553 0 net=7472
rlabel metal2 870 -2553 870 -2553 0 net=3206
rlabel metal2 898 -2553 898 -2553 0 net=8421
rlabel metal2 1017 -2553 1017 -2553 0 net=7555
rlabel metal2 1017 -2553 1017 -2553 0 net=7555
rlabel metal2 1024 -2553 1024 -2553 0 net=7777
rlabel metal2 247 -2555 247 -2555 0 net=2218
rlabel metal2 331 -2555 331 -2555 0 net=3638
rlabel metal2 492 -2555 492 -2555 0 net=2360
rlabel metal2 688 -2555 688 -2555 0 net=6748
rlabel metal2 744 -2555 744 -2555 0 net=6888
rlabel metal2 884 -2555 884 -2555 0 net=8180
rlabel metal2 254 -2557 254 -2557 0 net=2790
rlabel metal2 254 -2557 254 -2557 0 net=2790
rlabel metal2 268 -2557 268 -2557 0 net=7451
rlabel metal2 345 -2557 345 -2557 0 net=3995
rlabel metal2 401 -2557 401 -2557 0 net=1846
rlabel metal2 551 -2557 551 -2557 0 net=7516
rlabel metal2 663 -2557 663 -2557 0 net=4694
rlabel metal2 681 -2557 681 -2557 0 net=4902
rlabel metal2 947 -2557 947 -2557 0 net=7913
rlabel metal2 289 -2559 289 -2559 0 net=1788
rlabel metal2 415 -2559 415 -2559 0 net=1803
rlabel metal2 499 -2559 499 -2559 0 net=6677
rlabel metal2 499 -2559 499 -2559 0 net=6677
rlabel metal2 506 -2559 506 -2559 0 net=3892
rlabel metal2 621 -2559 621 -2559 0 net=8004
rlabel metal2 303 -2561 303 -2561 0 net=5692
rlabel metal2 600 -2561 600 -2561 0 net=6244
rlabel metal2 660 -2561 660 -2561 0 net=8351
rlabel metal2 691 -2561 691 -2561 0 net=756
rlabel metal2 691 -2561 691 -2561 0 net=756
rlabel metal2 716 -2561 716 -2561 0 net=7755
rlabel metal2 310 -2563 310 -2563 0 net=5380
rlabel metal2 723 -2563 723 -2563 0 net=5528
rlabel metal2 317 -2565 317 -2565 0 net=2093
rlabel metal2 359 -2565 359 -2565 0 net=2765
rlabel metal2 523 -2565 523 -2565 0 net=863
rlabel metal2 565 -2565 565 -2565 0 net=7104
rlabel metal2 723 -2565 723 -2565 0 net=7963
rlabel metal2 429 -2567 429 -2567 0 net=3462
rlabel metal2 527 -2567 527 -2567 0 net=6924
rlabel metal2 569 -2567 569 -2567 0 net=6200
rlabel metal2 730 -2567 730 -2567 0 net=7287
rlabel metal2 436 -2569 436 -2569 0 net=3056
rlabel metal2 576 -2569 576 -2569 0 net=2608
rlabel metal2 632 -2569 632 -2569 0 net=4282
rlabel metal2 747 -2569 747 -2569 0 net=1884
rlabel metal2 443 -2571 443 -2571 0 net=5586
rlabel metal2 513 -2571 513 -2571 0 net=7303
rlabel metal2 576 -2571 576 -2571 0 net=6555
rlabel metal2 695 -2571 695 -2571 0 net=3733
rlabel metal2 338 -2573 338 -2573 0 net=4792
rlabel metal2 530 -2573 530 -2573 0 net=4846
rlabel metal2 296 -2575 296 -2575 0 net=6037
rlabel metal2 373 -2575 373 -2575 0 net=7163
rlabel metal2 450 -2575 450 -2575 0 net=1175
rlabel metal2 352 -2577 352 -2577 0 net=2813
rlabel metal2 464 -2577 464 -2577 0 net=1770
rlabel metal2 373 -2579 373 -2579 0 net=2062
rlabel metal2 534 -2579 534 -2579 0 net=1924
rlabel metal2 408 -2581 408 -2581 0 net=2037
rlabel metal2 541 -2581 541 -2581 0 net=5338
rlabel metal2 562 -2583 562 -2583 0 net=7530
rlabel metal2 604 -2585 604 -2585 0 net=5920
rlabel metal2 131 -2596 131 -2596 0 net=6098
rlabel metal2 324 -2596 324 -2596 0 net=7452
rlabel metal2 443 -2596 443 -2596 0 net=7164
rlabel metal2 534 -2596 534 -2596 0 net=2038
rlabel metal2 674 -2596 674 -2596 0 net=7964
rlabel metal2 751 -2596 751 -2596 0 net=3734
rlabel metal2 810 -2596 810 -2596 0 net=7498
rlabel metal2 884 -2596 884 -2596 0 net=8422
rlabel metal2 954 -2596 954 -2596 0 net=7914
rlabel metal2 1010 -2596 1010 -2596 0 net=7556
rlabel metal2 1045 -2596 1045 -2596 0 net=8406
rlabel metal2 1055 -2596 1055 -2596 0 net=7888
rlabel metal2 331 -2598 331 -2598 0 net=2094
rlabel metal2 366 -2598 366 -2598 0 net=3996
rlabel metal2 450 -2598 450 -2598 0 net=2814
rlabel metal2 548 -2598 548 -2598 0 net=6556
rlabel metal2 660 -2598 660 -2598 0 net=8352
rlabel metal2 684 -2598 684 -2598 0 net=7756
rlabel metal2 961 -2598 961 -2598 0 net=6162
rlabel metal2 1013 -2598 1013 -2598 0 net=7778
rlabel metal2 338 -2600 338 -2600 0 net=6038
rlabel metal2 471 -2600 471 -2600 0 net=2370
rlabel metal2 555 -2600 555 -2600 0 net=7304
rlabel metal2 709 -2600 709 -2600 0 net=7288
rlabel metal2 492 -2602 492 -2602 0 net=1804
rlabel metal2 569 -2602 569 -2602 0 net=1176
rlabel metal2 499 -2604 499 -2604 0 net=6678
rlabel metal2 506 -2606 506 -2606 0 net=2766
<< end >>
