magic
tech scmos
timestamp 1555071776 
<< pdiffusion >>
rect 1 -8 7 -2
rect 8 -8 14 -2
rect 15 -8 21 -2
rect 50 -8 53 -2
rect 57 -8 63 -2
rect 64 -8 70 -2
rect 71 -8 77 -2
rect 78 -8 84 -2
rect 85 -8 88 -2
rect 92 -8 98 -2
rect 99 -8 102 -2
rect 106 -8 112 -2
rect 1 -25 7 -19
rect 8 -25 14 -19
rect 64 -25 70 -19
rect 71 -25 77 -19
rect 78 -25 84 -19
rect 85 -25 91 -19
rect 92 -25 95 -19
rect 99 -25 102 -19
rect 106 -25 112 -19
rect 113 -25 119 -19
rect 120 -25 123 -19
rect 1 -44 7 -38
rect 43 -44 49 -38
rect 50 -44 53 -38
rect 57 -44 60 -38
rect 64 -44 70 -38
rect 71 -44 77 -38
rect 78 -44 84 -38
rect 85 -44 91 -38
rect 92 -44 98 -38
rect 99 -44 102 -38
rect 106 -44 109 -38
rect 113 -44 116 -38
rect 1 -65 7 -59
rect 29 -65 32 -59
rect 36 -65 39 -59
rect 43 -65 49 -59
rect 50 -65 56 -59
rect 57 -65 60 -59
rect 64 -65 67 -59
rect 71 -65 74 -59
rect 78 -65 84 -59
rect 85 -65 91 -59
rect 92 -65 98 -59
rect 99 -65 102 -59
rect 106 -65 109 -59
rect 113 -65 119 -59
rect 22 -82 28 -76
rect 36 -82 42 -76
rect 43 -82 46 -76
rect 57 -82 63 -76
rect 64 -82 70 -76
rect 71 -82 74 -76
rect 78 -82 81 -76
rect 85 -82 91 -76
rect 92 -82 95 -76
rect 99 -82 102 -76
rect 106 -82 109 -76
rect 113 -82 119 -76
rect 120 -82 126 -76
rect 127 -82 130 -76
rect 134 -82 140 -76
rect 8 -103 11 -97
rect 15 -103 21 -97
rect 22 -103 28 -97
rect 29 -103 32 -97
rect 36 -103 42 -97
rect 43 -103 49 -97
rect 50 -103 53 -97
rect 57 -103 60 -97
rect 64 -103 67 -97
rect 71 -103 77 -97
rect 78 -103 84 -97
rect 85 -103 91 -97
rect 92 -103 98 -97
rect 99 -103 102 -97
rect 106 -103 109 -97
rect 113 -103 119 -97
rect 120 -103 123 -97
rect 127 -103 130 -97
rect 134 -103 137 -97
rect 141 -103 144 -97
rect 148 -103 151 -97
rect 155 -103 158 -97
rect 29 -130 32 -124
rect 36 -130 39 -124
rect 43 -130 46 -124
rect 50 -130 56 -124
rect 57 -130 63 -124
rect 64 -130 70 -124
rect 71 -130 74 -124
rect 78 -130 81 -124
rect 85 -130 91 -124
rect 92 -130 95 -124
rect 99 -130 105 -124
rect 106 -130 112 -124
rect 113 -130 119 -124
rect 120 -130 126 -124
rect 127 -130 130 -124
rect 134 -130 137 -124
rect 141 -130 144 -124
rect 148 -130 154 -124
rect 155 -130 158 -124
rect 162 -130 165 -124
rect 169 -130 172 -124
rect 176 -130 179 -124
rect 183 -130 189 -124
rect 190 -130 193 -124
rect 8 -161 11 -155
rect 15 -161 18 -155
rect 22 -161 25 -155
rect 29 -161 32 -155
rect 36 -161 39 -155
rect 43 -161 46 -155
rect 50 -161 56 -155
rect 57 -161 63 -155
rect 64 -161 70 -155
rect 71 -161 77 -155
rect 78 -161 81 -155
rect 85 -161 91 -155
rect 92 -161 95 -155
rect 99 -161 105 -155
rect 106 -161 109 -155
rect 113 -161 119 -155
rect 120 -161 126 -155
rect 127 -161 130 -155
rect 134 -161 140 -155
rect 141 -161 144 -155
rect 148 -161 151 -155
rect 155 -161 158 -155
rect 162 -161 165 -155
rect 169 -161 172 -155
rect 176 -161 179 -155
rect 183 -161 189 -155
rect 29 -194 32 -188
rect 36 -194 42 -188
rect 43 -194 49 -188
rect 50 -194 53 -188
rect 57 -194 60 -188
rect 64 -194 70 -188
rect 71 -194 77 -188
rect 78 -194 84 -188
rect 85 -194 91 -188
rect 92 -194 95 -188
rect 99 -194 105 -188
rect 106 -194 109 -188
rect 113 -194 119 -188
rect 120 -194 123 -188
rect 127 -194 133 -188
rect 134 -194 137 -188
rect 141 -194 144 -188
rect 148 -194 151 -188
rect 155 -194 158 -188
rect 162 -194 165 -188
rect 169 -194 172 -188
rect 176 -194 179 -188
rect 183 -194 189 -188
rect 190 -194 193 -188
rect 43 -217 49 -211
rect 50 -217 53 -211
rect 57 -217 63 -211
rect 71 -217 74 -211
rect 78 -217 84 -211
rect 85 -217 88 -211
rect 92 -217 95 -211
rect 99 -217 105 -211
rect 106 -217 109 -211
rect 113 -217 119 -211
rect 120 -217 123 -211
rect 127 -217 133 -211
rect 134 -217 140 -211
rect 141 -217 147 -211
rect 148 -217 151 -211
rect 155 -217 158 -211
rect 29 -242 32 -236
rect 36 -242 39 -236
rect 43 -242 46 -236
rect 50 -242 56 -236
rect 57 -242 63 -236
rect 64 -242 67 -236
rect 71 -242 77 -236
rect 78 -242 84 -236
rect 85 -242 91 -236
rect 92 -242 98 -236
rect 99 -242 105 -236
rect 106 -242 109 -236
rect 113 -242 116 -236
rect 120 -242 123 -236
rect 127 -242 130 -236
rect 134 -242 137 -236
rect 141 -242 144 -236
rect 50 -263 53 -257
rect 57 -263 63 -257
rect 64 -263 67 -257
rect 71 -263 74 -257
rect 78 -263 84 -257
rect 85 -263 91 -257
rect 92 -263 98 -257
rect 99 -263 105 -257
rect 106 -263 109 -257
rect 113 -263 116 -257
rect 120 -263 123 -257
rect 134 -263 140 -257
rect 134 -278 137 -272
rect 141 -278 147 -272
<< polysilicon >>
rect 51 -3 52 -1
rect 51 -9 52 -7
rect 58 -9 59 -7
rect 61 -9 62 -7
rect 65 -3 66 -1
rect 72 -9 73 -7
rect 79 -3 80 -1
rect 79 -9 80 -7
rect 86 -3 87 -1
rect 86 -9 87 -7
rect 93 -3 94 -1
rect 100 -3 101 -1
rect 100 -9 101 -7
rect 107 -9 108 -7
rect 110 -9 111 -7
rect 9 -26 10 -24
rect 12 -26 13 -24
rect 65 -20 66 -18
rect 68 -26 69 -24
rect 75 -20 76 -18
rect 72 -26 73 -24
rect 75 -26 76 -24
rect 82 -26 83 -24
rect 86 -20 87 -18
rect 89 -20 90 -18
rect 93 -20 94 -18
rect 93 -26 94 -24
rect 100 -20 101 -18
rect 100 -26 101 -24
rect 110 -26 111 -24
rect 114 -26 115 -24
rect 121 -20 122 -18
rect 121 -26 122 -24
rect 47 -39 48 -37
rect 51 -39 52 -37
rect 51 -45 52 -43
rect 58 -39 59 -37
rect 58 -45 59 -43
rect 68 -39 69 -37
rect 72 -39 73 -37
rect 75 -39 76 -37
rect 72 -45 73 -43
rect 82 -39 83 -37
rect 79 -45 80 -43
rect 82 -45 83 -43
rect 86 -39 87 -37
rect 89 -39 90 -37
rect 86 -45 87 -43
rect 96 -39 97 -37
rect 93 -45 94 -43
rect 96 -45 97 -43
rect 100 -39 101 -37
rect 100 -45 101 -43
rect 107 -39 108 -37
rect 107 -45 108 -43
rect 114 -39 115 -37
rect 114 -45 115 -43
rect 30 -60 31 -58
rect 30 -66 31 -64
rect 37 -60 38 -58
rect 37 -66 38 -64
rect 44 -60 45 -58
rect 47 -66 48 -64
rect 51 -60 52 -58
rect 54 -60 55 -58
rect 58 -60 59 -58
rect 58 -66 59 -64
rect 65 -60 66 -58
rect 65 -66 66 -64
rect 72 -60 73 -58
rect 72 -66 73 -64
rect 79 -60 80 -58
rect 82 -66 83 -64
rect 89 -60 90 -58
rect 86 -66 87 -64
rect 89 -66 90 -64
rect 96 -60 97 -58
rect 96 -66 97 -64
rect 100 -60 101 -58
rect 100 -66 101 -64
rect 107 -60 108 -58
rect 107 -66 108 -64
rect 114 -60 115 -58
rect 117 -60 118 -58
rect 117 -66 118 -64
rect 23 -83 24 -81
rect 26 -83 27 -81
rect 40 -77 41 -75
rect 40 -83 41 -81
rect 44 -77 45 -75
rect 44 -83 45 -81
rect 61 -77 62 -75
rect 58 -83 59 -81
rect 61 -83 62 -81
rect 65 -77 66 -75
rect 68 -77 69 -75
rect 65 -83 66 -81
rect 68 -83 69 -81
rect 72 -77 73 -75
rect 72 -83 73 -81
rect 79 -77 80 -75
rect 79 -83 80 -81
rect 86 -83 87 -81
rect 89 -83 90 -81
rect 93 -77 94 -75
rect 93 -83 94 -81
rect 100 -77 101 -75
rect 100 -83 101 -81
rect 107 -77 108 -75
rect 107 -83 108 -81
rect 114 -77 115 -75
rect 124 -77 125 -75
rect 124 -83 125 -81
rect 128 -77 129 -75
rect 128 -83 129 -81
rect 135 -83 136 -81
rect 9 -98 10 -96
rect 9 -104 10 -102
rect 16 -104 17 -102
rect 26 -104 27 -102
rect 30 -98 31 -96
rect 30 -104 31 -102
rect 40 -104 41 -102
rect 47 -104 48 -102
rect 51 -98 52 -96
rect 51 -104 52 -102
rect 58 -98 59 -96
rect 58 -104 59 -102
rect 65 -98 66 -96
rect 65 -104 66 -102
rect 72 -98 73 -96
rect 75 -98 76 -96
rect 72 -104 73 -102
rect 75 -104 76 -102
rect 79 -98 80 -96
rect 79 -104 80 -102
rect 82 -104 83 -102
rect 86 -98 87 -96
rect 89 -98 90 -96
rect 86 -104 87 -102
rect 89 -104 90 -102
rect 96 -98 97 -96
rect 93 -104 94 -102
rect 96 -104 97 -102
rect 100 -98 101 -96
rect 100 -104 101 -102
rect 107 -98 108 -96
rect 107 -104 108 -102
rect 114 -98 115 -96
rect 117 -104 118 -102
rect 121 -98 122 -96
rect 121 -104 122 -102
rect 128 -98 129 -96
rect 128 -104 129 -102
rect 135 -98 136 -96
rect 135 -104 136 -102
rect 142 -98 143 -96
rect 142 -104 143 -102
rect 149 -98 150 -96
rect 149 -104 150 -102
rect 156 -98 157 -96
rect 156 -104 157 -102
rect 30 -125 31 -123
rect 30 -131 31 -129
rect 37 -125 38 -123
rect 37 -131 38 -129
rect 44 -125 45 -123
rect 44 -131 45 -129
rect 51 -131 52 -129
rect 54 -131 55 -129
rect 61 -125 62 -123
rect 58 -131 59 -129
rect 61 -131 62 -129
rect 65 -125 66 -123
rect 65 -131 66 -129
rect 68 -131 69 -129
rect 72 -125 73 -123
rect 72 -131 73 -129
rect 79 -125 80 -123
rect 79 -131 80 -129
rect 86 -125 87 -123
rect 89 -125 90 -123
rect 86 -131 87 -129
rect 89 -131 90 -129
rect 93 -125 94 -123
rect 93 -131 94 -129
rect 103 -125 104 -123
rect 107 -125 108 -123
rect 110 -125 111 -123
rect 107 -131 108 -129
rect 110 -131 111 -129
rect 114 -125 115 -123
rect 117 -131 118 -129
rect 121 -125 122 -123
rect 124 -125 125 -123
rect 128 -125 129 -123
rect 128 -131 129 -129
rect 135 -125 136 -123
rect 135 -131 136 -129
rect 142 -125 143 -123
rect 142 -131 143 -129
rect 152 -125 153 -123
rect 149 -131 150 -129
rect 156 -125 157 -123
rect 156 -131 157 -129
rect 163 -125 164 -123
rect 163 -131 164 -129
rect 170 -125 171 -123
rect 170 -131 171 -129
rect 177 -125 178 -123
rect 177 -131 178 -129
rect 187 -125 188 -123
rect 184 -131 185 -129
rect 191 -125 192 -123
rect 191 -131 192 -129
rect 9 -156 10 -154
rect 9 -162 10 -160
rect 16 -156 17 -154
rect 16 -162 17 -160
rect 23 -156 24 -154
rect 23 -162 24 -160
rect 30 -156 31 -154
rect 30 -162 31 -160
rect 37 -156 38 -154
rect 37 -162 38 -160
rect 44 -156 45 -154
rect 44 -162 45 -160
rect 51 -156 52 -154
rect 54 -156 55 -154
rect 51 -162 52 -160
rect 61 -156 62 -154
rect 58 -162 59 -160
rect 61 -162 62 -160
rect 68 -156 69 -154
rect 65 -162 66 -160
rect 72 -156 73 -154
rect 72 -162 73 -160
rect 75 -162 76 -160
rect 79 -156 80 -154
rect 79 -162 80 -160
rect 86 -156 87 -154
rect 86 -162 87 -160
rect 93 -156 94 -154
rect 93 -162 94 -160
rect 100 -156 101 -154
rect 103 -162 104 -160
rect 107 -156 108 -154
rect 107 -162 108 -160
rect 114 -156 115 -154
rect 117 -162 118 -160
rect 121 -156 122 -154
rect 124 -156 125 -154
rect 121 -162 122 -160
rect 124 -162 125 -160
rect 128 -156 129 -154
rect 128 -162 129 -160
rect 135 -162 136 -160
rect 142 -156 143 -154
rect 142 -162 143 -160
rect 149 -156 150 -154
rect 149 -162 150 -160
rect 156 -156 157 -154
rect 156 -162 157 -160
rect 163 -156 164 -154
rect 163 -162 164 -160
rect 170 -156 171 -154
rect 170 -162 171 -160
rect 177 -156 178 -154
rect 177 -162 178 -160
rect 184 -156 185 -154
rect 184 -162 185 -160
rect 187 -162 188 -160
rect 30 -189 31 -187
rect 30 -195 31 -193
rect 37 -189 38 -187
rect 44 -189 45 -187
rect 47 -195 48 -193
rect 51 -189 52 -187
rect 51 -195 52 -193
rect 58 -189 59 -187
rect 58 -195 59 -193
rect 65 -189 66 -187
rect 68 -195 69 -193
rect 72 -189 73 -187
rect 75 -189 76 -187
rect 72 -195 73 -193
rect 79 -189 80 -187
rect 82 -189 83 -187
rect 86 -189 87 -187
rect 86 -195 87 -193
rect 93 -189 94 -187
rect 93 -195 94 -193
rect 100 -189 101 -187
rect 100 -195 101 -193
rect 103 -195 104 -193
rect 107 -189 108 -187
rect 107 -195 108 -193
rect 114 -189 115 -187
rect 117 -189 118 -187
rect 121 -189 122 -187
rect 121 -195 122 -193
rect 128 -189 129 -187
rect 131 -189 132 -187
rect 135 -189 136 -187
rect 135 -195 136 -193
rect 142 -189 143 -187
rect 142 -195 143 -193
rect 149 -189 150 -187
rect 149 -195 150 -193
rect 156 -189 157 -187
rect 156 -195 157 -193
rect 163 -189 164 -187
rect 163 -195 164 -193
rect 170 -189 171 -187
rect 170 -195 171 -193
rect 177 -189 178 -187
rect 177 -195 178 -193
rect 187 -189 188 -187
rect 191 -189 192 -187
rect 191 -195 192 -193
rect 44 -218 45 -216
rect 51 -212 52 -210
rect 51 -218 52 -216
rect 61 -212 62 -210
rect 72 -212 73 -210
rect 72 -218 73 -216
rect 82 -212 83 -210
rect 86 -212 87 -210
rect 86 -218 87 -216
rect 93 -212 94 -210
rect 93 -218 94 -216
rect 100 -218 101 -216
rect 103 -218 104 -216
rect 107 -212 108 -210
rect 107 -218 108 -216
rect 114 -212 115 -210
rect 117 -212 118 -210
rect 121 -212 122 -210
rect 121 -218 122 -216
rect 128 -212 129 -210
rect 128 -218 129 -216
rect 131 -218 132 -216
rect 138 -212 139 -210
rect 138 -218 139 -216
rect 142 -218 143 -216
rect 149 -212 150 -210
rect 149 -218 150 -216
rect 156 -212 157 -210
rect 156 -218 157 -216
rect 30 -237 31 -235
rect 30 -243 31 -241
rect 37 -237 38 -235
rect 37 -243 38 -241
rect 44 -237 45 -235
rect 44 -243 45 -241
rect 51 -237 52 -235
rect 54 -237 55 -235
rect 54 -243 55 -241
rect 58 -237 59 -235
rect 61 -237 62 -235
rect 65 -237 66 -235
rect 65 -243 66 -241
rect 75 -237 76 -235
rect 72 -243 73 -241
rect 75 -243 76 -241
rect 79 -237 80 -235
rect 82 -237 83 -235
rect 82 -243 83 -241
rect 86 -237 87 -235
rect 89 -237 90 -235
rect 86 -243 87 -241
rect 89 -243 90 -241
rect 93 -237 94 -235
rect 93 -243 94 -241
rect 103 -237 104 -235
rect 100 -243 101 -241
rect 107 -237 108 -235
rect 107 -243 108 -241
rect 114 -237 115 -235
rect 114 -243 115 -241
rect 121 -237 122 -235
rect 121 -243 122 -241
rect 128 -237 129 -235
rect 128 -243 129 -241
rect 135 -237 136 -235
rect 135 -243 136 -241
rect 142 -237 143 -235
rect 142 -243 143 -241
rect 51 -258 52 -256
rect 51 -264 52 -262
rect 61 -258 62 -256
rect 58 -264 59 -262
rect 65 -258 66 -256
rect 65 -264 66 -262
rect 72 -258 73 -256
rect 72 -264 73 -262
rect 79 -258 80 -256
rect 82 -264 83 -262
rect 86 -264 87 -262
rect 89 -264 90 -262
rect 96 -258 97 -256
rect 96 -264 97 -262
rect 103 -264 104 -262
rect 107 -258 108 -256
rect 107 -264 108 -262
rect 114 -258 115 -256
rect 114 -264 115 -262
rect 121 -258 122 -256
rect 121 -264 122 -262
rect 138 -258 139 -256
rect 138 -264 139 -262
rect 135 -273 136 -271
rect 135 -279 136 -277
rect 145 -279 146 -277
<< metal1 >>
rect 51 0 66 1
rect 79 0 87 1
rect 93 0 101 1
rect 51 -11 62 -10
rect 65 -11 73 -10
rect 79 -11 111 -10
rect 58 -13 76 -12
rect 89 -13 101 -12
rect 107 -13 122 -12
rect 86 -15 101 -14
rect 86 -17 94 -16
rect 9 -28 13 -27
rect 58 -28 90 -27
rect 107 -28 111 -27
rect 114 -28 122 -27
rect 68 -30 76 -29
rect 82 -30 101 -29
rect 47 -32 76 -31
rect 86 -32 115 -31
rect 51 -34 69 -33
rect 72 -34 83 -33
rect 96 -34 101 -33
rect 72 -36 94 -35
rect 37 -47 45 -46
rect 51 -47 83 -46
rect 89 -47 115 -46
rect 30 -49 52 -48
rect 54 -49 66 -48
rect 79 -49 118 -48
rect 72 -51 80 -50
rect 96 -51 108 -50
rect 58 -53 97 -52
rect 100 -53 108 -52
rect 58 -55 94 -54
rect 100 -55 115 -54
rect 72 -57 87 -56
rect 30 -68 48 -67
rect 58 -68 87 -67
rect 93 -68 125 -67
rect 37 -70 62 -69
rect 65 -70 69 -69
rect 72 -70 83 -69
rect 96 -70 108 -69
rect 117 -70 129 -69
rect 40 -72 45 -71
rect 65 -72 73 -71
rect 79 -72 101 -71
rect 107 -72 115 -71
rect 89 -74 101 -73
rect 9 -85 24 -84
rect 26 -85 41 -84
rect 51 -85 97 -84
rect 100 -85 122 -84
rect 128 -85 143 -84
rect 30 -87 45 -86
rect 58 -87 69 -86
rect 75 -87 129 -86
rect 79 -89 90 -88
rect 107 -89 125 -88
rect 58 -91 80 -90
rect 86 -91 101 -90
rect 114 -91 150 -90
rect 65 -93 90 -92
rect 93 -93 108 -92
rect 61 -95 66 -94
rect 86 -95 157 -94
rect 9 -106 17 -105
rect 26 -106 73 -105
rect 82 -106 122 -105
rect 124 -106 171 -105
rect 187 -106 192 -105
rect 30 -108 41 -107
rect 44 -108 62 -107
rect 65 -108 73 -107
rect 86 -108 101 -107
rect 103 -108 150 -107
rect 30 -110 111 -109
rect 117 -110 136 -109
rect 142 -110 178 -109
rect 37 -112 80 -111
rect 93 -112 108 -111
rect 114 -112 143 -111
rect 47 -114 59 -113
rect 75 -114 94 -113
rect 121 -114 164 -113
rect 51 -116 90 -115
rect 135 -116 157 -115
rect 65 -118 90 -117
rect 152 -118 157 -117
rect 79 -120 97 -119
rect 86 -122 108 -121
rect 23 -133 45 -132
rect 61 -133 94 -132
rect 110 -133 178 -132
rect 16 -135 62 -134
rect 68 -135 73 -134
rect 79 -135 90 -134
rect 107 -135 178 -134
rect 30 -137 52 -136
rect 68 -137 80 -136
rect 100 -137 108 -136
rect 117 -137 136 -136
rect 149 -137 171 -136
rect 9 -139 52 -138
rect 72 -139 87 -138
rect 121 -139 164 -138
rect 30 -141 59 -140
rect 124 -141 150 -140
rect 156 -141 171 -140
rect 44 -143 66 -142
rect 114 -143 157 -142
rect 128 -145 185 -144
rect 86 -147 129 -146
rect 142 -147 164 -146
rect 184 -147 192 -146
rect 37 -149 143 -148
rect 37 -151 55 -150
rect 54 -153 94 -152
rect 9 -164 73 -163
rect 75 -164 188 -163
rect 23 -166 52 -165
rect 61 -166 108 -165
rect 128 -166 192 -165
rect 30 -168 66 -167
rect 79 -168 108 -167
rect 128 -168 164 -167
rect 30 -170 83 -169
rect 103 -170 122 -169
rect 131 -170 164 -169
rect 37 -172 59 -171
rect 117 -172 122 -171
rect 135 -172 171 -171
rect 16 -174 38 -173
rect 44 -174 87 -173
rect 117 -174 150 -173
rect 156 -174 185 -173
rect 44 -176 125 -175
rect 149 -176 178 -175
rect 51 -178 73 -177
rect 75 -178 87 -177
rect 114 -178 157 -177
rect 170 -178 188 -177
rect 58 -180 94 -179
rect 142 -180 178 -179
rect 65 -182 136 -181
rect 79 -184 143 -183
rect 93 -186 101 -185
rect 30 -197 62 -196
rect 68 -197 108 -196
rect 117 -197 164 -196
rect 58 -199 73 -198
rect 86 -199 178 -198
rect 51 -201 73 -200
rect 82 -201 87 -200
rect 100 -201 122 -200
rect 128 -201 171 -200
rect 47 -203 52 -202
rect 93 -203 122 -202
rect 138 -203 150 -202
rect 93 -205 115 -204
rect 142 -205 150 -204
rect 103 -207 192 -206
rect 107 -209 136 -208
rect 30 -220 59 -219
rect 61 -220 94 -219
rect 103 -220 136 -219
rect 138 -220 150 -219
rect 44 -222 52 -221
rect 54 -222 101 -221
rect 103 -222 108 -221
rect 121 -222 132 -221
rect 142 -222 157 -221
rect 37 -224 52 -223
rect 65 -224 83 -223
rect 89 -224 115 -223
rect 128 -224 143 -223
rect 44 -226 94 -225
rect 75 -228 108 -227
rect 79 -230 122 -229
rect 86 -232 129 -231
rect 72 -234 87 -233
rect 30 -245 62 -244
rect 79 -245 115 -244
rect 138 -245 143 -244
rect 37 -247 76 -246
rect 86 -247 129 -246
rect 44 -249 73 -248
rect 89 -249 122 -248
rect 51 -251 97 -250
rect 121 -251 136 -250
rect 54 -253 83 -252
rect 93 -253 115 -252
rect 72 -255 101 -254
rect 51 -266 59 -265
rect 65 -266 90 -265
rect 96 -266 122 -265
rect 135 -266 139 -265
rect 72 -268 83 -267
rect 86 -268 108 -267
rect 103 -270 115 -269
rect 135 -281 146 -280
<< m2contact >>
rect 51 0 52 1
rect 65 0 66 1
rect 79 0 80 1
rect 86 0 87 1
rect 93 0 94 1
rect 100 0 101 1
rect 51 -11 52 -10
rect 61 -11 62 -10
rect 65 -11 66 -10
rect 72 -11 73 -10
rect 79 -11 80 -10
rect 110 -11 111 -10
rect 58 -13 59 -12
rect 75 -13 76 -12
rect 89 -13 90 -12
rect 100 -13 101 -12
rect 107 -13 108 -12
rect 121 -13 122 -12
rect 86 -15 87 -14
rect 100 -15 101 -14
rect 86 -17 87 -16
rect 93 -17 94 -16
rect 9 -28 10 -27
rect 12 -28 13 -27
rect 58 -28 59 -27
rect 89 -28 90 -27
rect 107 -28 108 -27
rect 110 -28 111 -27
rect 114 -28 115 -27
rect 121 -28 122 -27
rect 68 -30 69 -29
rect 75 -30 76 -29
rect 82 -30 83 -29
rect 100 -30 101 -29
rect 47 -32 48 -31
rect 75 -32 76 -31
rect 86 -32 87 -31
rect 114 -32 115 -31
rect 51 -34 52 -33
rect 68 -34 69 -33
rect 72 -34 73 -33
rect 82 -34 83 -33
rect 96 -34 97 -33
rect 100 -34 101 -33
rect 72 -36 73 -35
rect 93 -36 94 -35
rect 37 -47 38 -46
rect 44 -47 45 -46
rect 51 -47 52 -46
rect 82 -47 83 -46
rect 89 -47 90 -46
rect 114 -47 115 -46
rect 30 -49 31 -48
rect 51 -49 52 -48
rect 54 -49 55 -48
rect 65 -49 66 -48
rect 79 -49 80 -48
rect 117 -49 118 -48
rect 72 -51 73 -50
rect 79 -51 80 -50
rect 96 -51 97 -50
rect 107 -51 108 -50
rect 58 -53 59 -52
rect 96 -53 97 -52
rect 100 -53 101 -52
rect 107 -53 108 -52
rect 58 -55 59 -54
rect 93 -55 94 -54
rect 100 -55 101 -54
rect 114 -55 115 -54
rect 72 -57 73 -56
rect 86 -57 87 -56
rect 30 -68 31 -67
rect 47 -68 48 -67
rect 58 -68 59 -67
rect 86 -68 87 -67
rect 93 -68 94 -67
rect 124 -68 125 -67
rect 37 -70 38 -69
rect 61 -70 62 -69
rect 65 -70 66 -69
rect 68 -70 69 -69
rect 72 -70 73 -69
rect 82 -70 83 -69
rect 96 -70 97 -69
rect 107 -70 108 -69
rect 117 -70 118 -69
rect 128 -70 129 -69
rect 40 -72 41 -71
rect 44 -72 45 -71
rect 65 -72 66 -71
rect 72 -72 73 -71
rect 79 -72 80 -71
rect 100 -72 101 -71
rect 107 -72 108 -71
rect 114 -72 115 -71
rect 89 -74 90 -73
rect 100 -74 101 -73
rect 9 -85 10 -84
rect 23 -85 24 -84
rect 26 -85 27 -84
rect 40 -85 41 -84
rect 51 -85 52 -84
rect 96 -85 97 -84
rect 100 -85 101 -84
rect 121 -85 122 -84
rect 128 -85 129 -84
rect 142 -85 143 -84
rect 30 -87 31 -86
rect 44 -87 45 -86
rect 58 -87 59 -86
rect 68 -87 69 -86
rect 75 -87 76 -86
rect 128 -87 129 -86
rect 79 -89 80 -88
rect 89 -89 90 -88
rect 107 -89 108 -88
rect 124 -89 125 -88
rect 58 -91 59 -90
rect 79 -91 80 -90
rect 86 -91 87 -90
rect 100 -91 101 -90
rect 114 -91 115 -90
rect 149 -91 150 -90
rect 65 -93 66 -92
rect 89 -93 90 -92
rect 93 -93 94 -92
rect 107 -93 108 -92
rect 61 -95 62 -94
rect 65 -95 66 -94
rect 86 -95 87 -94
rect 156 -95 157 -94
rect 9 -106 10 -105
rect 16 -106 17 -105
rect 26 -106 27 -105
rect 72 -106 73 -105
rect 82 -106 83 -105
rect 121 -106 122 -105
rect 124 -106 125 -105
rect 170 -106 171 -105
rect 187 -106 188 -105
rect 191 -106 192 -105
rect 30 -108 31 -107
rect 40 -108 41 -107
rect 44 -108 45 -107
rect 61 -108 62 -107
rect 65 -108 66 -107
rect 72 -108 73 -107
rect 86 -108 87 -107
rect 100 -108 101 -107
rect 103 -108 104 -107
rect 149 -108 150 -107
rect 30 -110 31 -109
rect 110 -110 111 -109
rect 117 -110 118 -109
rect 135 -110 136 -109
rect 142 -110 143 -109
rect 177 -110 178 -109
rect 37 -112 38 -111
rect 79 -112 80 -111
rect 93 -112 94 -111
rect 107 -112 108 -111
rect 114 -112 115 -111
rect 142 -112 143 -111
rect 47 -114 48 -113
rect 58 -114 59 -113
rect 75 -114 76 -113
rect 93 -114 94 -113
rect 121 -114 122 -113
rect 163 -114 164 -113
rect 51 -116 52 -115
rect 89 -116 90 -115
rect 135 -116 136 -115
rect 156 -116 157 -115
rect 65 -118 66 -117
rect 89 -118 90 -117
rect 152 -118 153 -117
rect 156 -118 157 -117
rect 79 -120 80 -119
rect 96 -120 97 -119
rect 86 -122 87 -121
rect 107 -122 108 -121
rect 23 -133 24 -132
rect 44 -133 45 -132
rect 61 -133 62 -132
rect 93 -133 94 -132
rect 110 -133 111 -132
rect 177 -133 178 -132
rect 16 -135 17 -134
rect 61 -135 62 -134
rect 68 -135 69 -134
rect 72 -135 73 -134
rect 79 -135 80 -134
rect 89 -135 90 -134
rect 107 -135 108 -134
rect 177 -135 178 -134
rect 30 -137 31 -136
rect 51 -137 52 -136
rect 68 -137 69 -136
rect 79 -137 80 -136
rect 100 -137 101 -136
rect 107 -137 108 -136
rect 117 -137 118 -136
rect 135 -137 136 -136
rect 149 -137 150 -136
rect 170 -137 171 -136
rect 9 -139 10 -138
rect 51 -139 52 -138
rect 72 -139 73 -138
rect 86 -139 87 -138
rect 121 -139 122 -138
rect 163 -139 164 -138
rect 30 -141 31 -140
rect 58 -141 59 -140
rect 124 -141 125 -140
rect 149 -141 150 -140
rect 156 -141 157 -140
rect 170 -141 171 -140
rect 44 -143 45 -142
rect 65 -143 66 -142
rect 114 -143 115 -142
rect 156 -143 157 -142
rect 128 -145 129 -144
rect 184 -145 185 -144
rect 86 -147 87 -146
rect 128 -147 129 -146
rect 142 -147 143 -146
rect 163 -147 164 -146
rect 184 -147 185 -146
rect 191 -147 192 -146
rect 37 -149 38 -148
rect 142 -149 143 -148
rect 37 -151 38 -150
rect 54 -151 55 -150
rect 54 -153 55 -152
rect 93 -153 94 -152
rect 9 -164 10 -163
rect 72 -164 73 -163
rect 75 -164 76 -163
rect 187 -164 188 -163
rect 23 -166 24 -165
rect 51 -166 52 -165
rect 61 -166 62 -165
rect 107 -166 108 -165
rect 128 -166 129 -165
rect 191 -166 192 -165
rect 30 -168 31 -167
rect 65 -168 66 -167
rect 79 -168 80 -167
rect 107 -168 108 -167
rect 128 -168 129 -167
rect 163 -168 164 -167
rect 30 -170 31 -169
rect 82 -170 83 -169
rect 103 -170 104 -169
rect 121 -170 122 -169
rect 131 -170 132 -169
rect 163 -170 164 -169
rect 37 -172 38 -171
rect 58 -172 59 -171
rect 117 -172 118 -171
rect 121 -172 122 -171
rect 135 -172 136 -171
rect 170 -172 171 -171
rect 16 -174 17 -173
rect 37 -174 38 -173
rect 44 -174 45 -173
rect 86 -174 87 -173
rect 117 -174 118 -173
rect 149 -174 150 -173
rect 156 -174 157 -173
rect 184 -174 185 -173
rect 44 -176 45 -175
rect 124 -176 125 -175
rect 149 -176 150 -175
rect 177 -176 178 -175
rect 51 -178 52 -177
rect 72 -178 73 -177
rect 75 -178 76 -177
rect 86 -178 87 -177
rect 114 -178 115 -177
rect 156 -178 157 -177
rect 170 -178 171 -177
rect 187 -178 188 -177
rect 58 -180 59 -179
rect 93 -180 94 -179
rect 142 -180 143 -179
rect 177 -180 178 -179
rect 65 -182 66 -181
rect 135 -182 136 -181
rect 79 -184 80 -183
rect 142 -184 143 -183
rect 93 -186 94 -185
rect 100 -186 101 -185
rect 30 -197 31 -196
rect 61 -197 62 -196
rect 68 -197 69 -196
rect 107 -197 108 -196
rect 117 -197 118 -196
rect 163 -197 164 -196
rect 58 -199 59 -198
rect 72 -199 73 -198
rect 86 -199 87 -198
rect 177 -199 178 -198
rect 51 -201 52 -200
rect 72 -201 73 -200
rect 82 -201 83 -200
rect 86 -201 87 -200
rect 100 -201 101 -200
rect 121 -201 122 -200
rect 128 -201 129 -200
rect 170 -201 171 -200
rect 47 -203 48 -202
rect 51 -203 52 -202
rect 93 -203 94 -202
rect 121 -203 122 -202
rect 138 -203 139 -202
rect 149 -203 150 -202
rect 93 -205 94 -204
rect 114 -205 115 -204
rect 142 -205 143 -204
rect 149 -205 150 -204
rect 103 -207 104 -206
rect 191 -207 192 -206
rect 107 -209 108 -208
rect 135 -209 136 -208
rect 30 -220 31 -219
rect 58 -220 59 -219
rect 61 -220 62 -219
rect 93 -220 94 -219
rect 103 -220 104 -219
rect 135 -220 136 -219
rect 138 -220 139 -219
rect 149 -220 150 -219
rect 44 -222 45 -221
rect 51 -222 52 -221
rect 54 -222 55 -221
rect 100 -222 101 -221
rect 103 -222 104 -221
rect 107 -222 108 -221
rect 121 -222 122 -221
rect 131 -222 132 -221
rect 142 -222 143 -221
rect 156 -222 157 -221
rect 37 -224 38 -223
rect 51 -224 52 -223
rect 65 -224 66 -223
rect 82 -224 83 -223
rect 89 -224 90 -223
rect 114 -224 115 -223
rect 128 -224 129 -223
rect 142 -224 143 -223
rect 44 -226 45 -225
rect 93 -226 94 -225
rect 75 -228 76 -227
rect 107 -228 108 -227
rect 79 -230 80 -229
rect 121 -230 122 -229
rect 86 -232 87 -231
rect 128 -232 129 -231
rect 72 -234 73 -233
rect 86 -234 87 -233
rect 30 -245 31 -244
rect 61 -245 62 -244
rect 79 -245 80 -244
rect 114 -245 115 -244
rect 138 -245 139 -244
rect 142 -245 143 -244
rect 37 -247 38 -246
rect 75 -247 76 -246
rect 86 -247 87 -246
rect 128 -247 129 -246
rect 44 -249 45 -248
rect 72 -249 73 -248
rect 89 -249 90 -248
rect 121 -249 122 -248
rect 51 -251 52 -250
rect 96 -251 97 -250
rect 121 -251 122 -250
rect 135 -251 136 -250
rect 54 -253 55 -252
rect 82 -253 83 -252
rect 93 -253 94 -252
rect 114 -253 115 -252
rect 72 -255 73 -254
rect 100 -255 101 -254
rect 51 -266 52 -265
rect 58 -266 59 -265
rect 65 -266 66 -265
rect 89 -266 90 -265
rect 96 -266 97 -265
rect 121 -266 122 -265
rect 135 -266 136 -265
rect 138 -266 139 -265
rect 72 -268 73 -267
rect 82 -268 83 -267
rect 86 -268 87 -267
rect 107 -268 108 -267
rect 103 -270 104 -269
rect 114 -270 115 -269
rect 135 -281 136 -280
rect 145 -281 146 -280
<< metal2 >>
rect 51 -1 52 1
rect 65 -1 66 1
rect 79 -1 80 1
rect 86 -1 87 1
rect 93 -1 94 1
rect 100 -1 101 1
rect 51 -11 52 -9
rect 61 -11 62 -9
rect 65 -18 66 -10
rect 72 -11 73 -9
rect 79 -11 80 -9
rect 110 -11 111 -9
rect 58 -13 59 -9
rect 75 -18 76 -12
rect 89 -18 90 -12
rect 100 -13 101 -9
rect 107 -13 108 -9
rect 121 -18 122 -12
rect 86 -15 87 -9
rect 100 -18 101 -14
rect 86 -18 87 -16
rect 93 -18 94 -16
rect 9 -28 10 -26
rect 12 -28 13 -26
rect 58 -37 59 -27
rect 89 -37 90 -27
rect 107 -37 108 -27
rect 110 -28 111 -26
rect 114 -28 115 -26
rect 121 -28 122 -26
rect 68 -30 69 -26
rect 75 -30 76 -26
rect 82 -30 83 -26
rect 100 -30 101 -26
rect 47 -37 48 -31
rect 75 -37 76 -31
rect 86 -37 87 -31
rect 114 -37 115 -31
rect 51 -37 52 -33
rect 68 -37 69 -33
rect 72 -34 73 -26
rect 82 -37 83 -33
rect 96 -37 97 -33
rect 100 -37 101 -33
rect 72 -37 73 -35
rect 93 -36 94 -26
rect 37 -58 38 -46
rect 44 -58 45 -46
rect 51 -47 52 -45
rect 82 -47 83 -45
rect 89 -58 90 -46
rect 114 -47 115 -45
rect 30 -58 31 -48
rect 51 -58 52 -48
rect 54 -58 55 -48
rect 65 -58 66 -48
rect 79 -49 80 -45
rect 117 -58 118 -48
rect 72 -51 73 -45
rect 79 -58 80 -50
rect 96 -51 97 -45
rect 107 -51 108 -45
rect 58 -53 59 -45
rect 96 -58 97 -52
rect 100 -53 101 -45
rect 107 -58 108 -52
rect 58 -58 59 -54
rect 93 -55 94 -45
rect 100 -58 101 -54
rect 114 -58 115 -54
rect 72 -58 73 -56
rect 86 -57 87 -45
rect 30 -68 31 -66
rect 47 -68 48 -66
rect 58 -68 59 -66
rect 86 -68 87 -66
rect 93 -75 94 -67
rect 124 -75 125 -67
rect 37 -70 38 -66
rect 61 -75 62 -69
rect 65 -70 66 -66
rect 68 -75 69 -69
rect 72 -70 73 -66
rect 82 -70 83 -66
rect 96 -70 97 -66
rect 107 -70 108 -66
rect 117 -70 118 -66
rect 128 -75 129 -69
rect 40 -75 41 -71
rect 44 -75 45 -71
rect 65 -75 66 -71
rect 72 -75 73 -71
rect 79 -75 80 -71
rect 100 -72 101 -66
rect 107 -75 108 -71
rect 114 -75 115 -71
rect 89 -74 90 -66
rect 100 -75 101 -73
rect 9 -96 10 -84
rect 23 -85 24 -83
rect 26 -85 27 -83
rect 40 -85 41 -83
rect 51 -96 52 -84
rect 96 -96 97 -84
rect 100 -85 101 -83
rect 121 -96 122 -84
rect 128 -85 129 -83
rect 142 -96 143 -84
rect 30 -96 31 -86
rect 44 -87 45 -83
rect 58 -87 59 -83
rect 68 -87 69 -83
rect 72 -87 73 -83
rect 72 -96 73 -86
rect 72 -87 73 -83
rect 72 -96 73 -86
rect 75 -96 76 -86
rect 128 -96 129 -86
rect 135 -87 136 -83
rect 135 -96 136 -86
rect 135 -87 136 -83
rect 135 -96 136 -86
rect 79 -89 80 -83
rect 89 -89 90 -83
rect 107 -89 108 -83
rect 124 -89 125 -83
rect 58 -96 59 -90
rect 79 -96 80 -90
rect 86 -91 87 -83
rect 100 -96 101 -90
rect 114 -96 115 -90
rect 149 -96 150 -90
rect 65 -93 66 -83
rect 89 -96 90 -92
rect 93 -93 94 -83
rect 107 -96 108 -92
rect 61 -95 62 -83
rect 65 -96 66 -94
rect 86 -96 87 -94
rect 156 -96 157 -94
rect 9 -106 10 -104
rect 16 -106 17 -104
rect 26 -106 27 -104
rect 72 -106 73 -104
rect 82 -106 83 -104
rect 121 -106 122 -104
rect 124 -123 125 -105
rect 170 -123 171 -105
rect 187 -123 188 -105
rect 191 -123 192 -105
rect 30 -108 31 -104
rect 40 -108 41 -104
rect 44 -123 45 -107
rect 61 -123 62 -107
rect 65 -108 66 -104
rect 72 -123 73 -107
rect 86 -108 87 -104
rect 100 -108 101 -104
rect 103 -123 104 -107
rect 149 -108 150 -104
rect 30 -123 31 -109
rect 110 -123 111 -109
rect 117 -110 118 -104
rect 135 -110 136 -104
rect 142 -110 143 -104
rect 177 -123 178 -109
rect 37 -123 38 -111
rect 79 -112 80 -104
rect 93 -112 94 -104
rect 107 -112 108 -104
rect 114 -123 115 -111
rect 142 -123 143 -111
rect 47 -114 48 -104
rect 58 -114 59 -104
rect 75 -114 76 -104
rect 93 -123 94 -113
rect 121 -123 122 -113
rect 163 -123 164 -113
rect 51 -116 52 -104
rect 89 -116 90 -104
rect 128 -116 129 -104
rect 128 -123 129 -115
rect 128 -116 129 -104
rect 128 -123 129 -115
rect 135 -123 136 -115
rect 156 -116 157 -104
rect 65 -123 66 -117
rect 89 -123 90 -117
rect 152 -123 153 -117
rect 156 -123 157 -117
rect 79 -123 80 -119
rect 96 -120 97 -104
rect 86 -123 87 -121
rect 107 -123 108 -121
rect 23 -154 24 -132
rect 44 -133 45 -131
rect 61 -133 62 -131
rect 93 -133 94 -131
rect 110 -133 111 -131
rect 177 -133 178 -131
rect 16 -154 17 -134
rect 61 -154 62 -134
rect 68 -135 69 -131
rect 72 -135 73 -131
rect 79 -135 80 -131
rect 89 -135 90 -131
rect 107 -135 108 -131
rect 177 -154 178 -134
rect 30 -137 31 -131
rect 51 -137 52 -131
rect 68 -154 69 -136
rect 79 -154 80 -136
rect 100 -154 101 -136
rect 107 -154 108 -136
rect 117 -137 118 -131
rect 135 -137 136 -131
rect 149 -137 150 -131
rect 170 -137 171 -131
rect 9 -154 10 -138
rect 51 -154 52 -138
rect 72 -154 73 -138
rect 86 -139 87 -131
rect 121 -154 122 -138
rect 163 -139 164 -131
rect 30 -154 31 -140
rect 58 -141 59 -131
rect 124 -154 125 -140
rect 149 -154 150 -140
rect 156 -141 157 -131
rect 170 -154 171 -140
rect 44 -154 45 -142
rect 65 -143 66 -131
rect 114 -154 115 -142
rect 156 -154 157 -142
rect 128 -145 129 -131
rect 184 -145 185 -131
rect 86 -154 87 -146
rect 128 -154 129 -146
rect 142 -147 143 -131
rect 163 -154 164 -146
rect 184 -154 185 -146
rect 191 -147 192 -131
rect 37 -149 38 -131
rect 142 -154 143 -148
rect 37 -154 38 -150
rect 54 -151 55 -131
rect 54 -154 55 -152
rect 93 -154 94 -152
rect 9 -164 10 -162
rect 72 -164 73 -162
rect 75 -164 76 -162
rect 187 -164 188 -162
rect 23 -166 24 -162
rect 51 -166 52 -162
rect 61 -166 62 -162
rect 107 -166 108 -162
rect 128 -166 129 -162
rect 191 -187 192 -165
rect 30 -168 31 -162
rect 65 -168 66 -162
rect 79 -168 80 -162
rect 107 -187 108 -167
rect 128 -187 129 -167
rect 163 -168 164 -162
rect 30 -187 31 -169
rect 82 -187 83 -169
rect 103 -170 104 -162
rect 121 -170 122 -162
rect 131 -187 132 -169
rect 163 -187 164 -169
rect 37 -172 38 -162
rect 58 -172 59 -162
rect 117 -172 118 -162
rect 121 -187 122 -171
rect 135 -172 136 -162
rect 170 -172 171 -162
rect 16 -174 17 -162
rect 37 -187 38 -173
rect 44 -174 45 -162
rect 86 -174 87 -162
rect 117 -187 118 -173
rect 149 -174 150 -162
rect 156 -174 157 -162
rect 184 -174 185 -162
rect 44 -187 45 -175
rect 124 -176 125 -162
rect 149 -187 150 -175
rect 177 -176 178 -162
rect 51 -187 52 -177
rect 72 -187 73 -177
rect 75 -187 76 -177
rect 86 -187 87 -177
rect 114 -187 115 -177
rect 156 -187 157 -177
rect 170 -187 171 -177
rect 187 -187 188 -177
rect 58 -187 59 -179
rect 93 -180 94 -162
rect 142 -180 143 -162
rect 177 -187 178 -179
rect 65 -187 66 -181
rect 135 -187 136 -181
rect 79 -187 80 -183
rect 142 -187 143 -183
rect 93 -187 94 -185
rect 100 -187 101 -185
rect 30 -197 31 -195
rect 61 -210 62 -196
rect 68 -197 69 -195
rect 107 -197 108 -195
rect 117 -210 118 -196
rect 163 -197 164 -195
rect 58 -199 59 -195
rect 72 -199 73 -195
rect 86 -199 87 -195
rect 177 -199 178 -195
rect 51 -201 52 -195
rect 72 -210 73 -200
rect 82 -210 83 -200
rect 86 -210 87 -200
rect 100 -201 101 -195
rect 121 -201 122 -195
rect 128 -210 129 -200
rect 170 -201 171 -195
rect 47 -203 48 -195
rect 51 -210 52 -202
rect 93 -203 94 -195
rect 121 -210 122 -202
rect 138 -210 139 -202
rect 149 -203 150 -195
rect 156 -203 157 -195
rect 156 -210 157 -202
rect 156 -203 157 -195
rect 156 -210 157 -202
rect 93 -210 94 -204
rect 114 -210 115 -204
rect 142 -205 143 -195
rect 149 -210 150 -204
rect 103 -207 104 -195
rect 191 -207 192 -195
rect 107 -210 108 -208
rect 135 -209 136 -195
rect 30 -235 31 -219
rect 58 -235 59 -219
rect 61 -235 62 -219
rect 93 -220 94 -218
rect 103 -220 104 -218
rect 135 -235 136 -219
rect 138 -220 139 -218
rect 149 -220 150 -218
rect 44 -222 45 -218
rect 51 -222 52 -218
rect 54 -235 55 -221
rect 100 -222 101 -218
rect 103 -235 104 -221
rect 107 -222 108 -218
rect 121 -222 122 -218
rect 131 -222 132 -218
rect 142 -222 143 -218
rect 156 -222 157 -218
rect 37 -235 38 -223
rect 51 -235 52 -223
rect 65 -235 66 -223
rect 82 -235 83 -223
rect 89 -235 90 -223
rect 114 -235 115 -223
rect 128 -224 129 -218
rect 142 -235 143 -223
rect 44 -235 45 -225
rect 93 -235 94 -225
rect 75 -235 76 -227
rect 107 -235 108 -227
rect 79 -235 80 -229
rect 121 -235 122 -229
rect 86 -232 87 -218
rect 128 -235 129 -231
rect 72 -234 73 -218
rect 86 -235 87 -233
rect 30 -245 31 -243
rect 61 -256 62 -244
rect 65 -245 66 -243
rect 65 -256 66 -244
rect 65 -245 66 -243
rect 65 -256 66 -244
rect 79 -256 80 -244
rect 114 -245 115 -243
rect 138 -256 139 -244
rect 142 -245 143 -243
rect 37 -247 38 -243
rect 75 -247 76 -243
rect 86 -247 87 -243
rect 128 -247 129 -243
rect 44 -249 45 -243
rect 72 -249 73 -243
rect 89 -249 90 -243
rect 121 -249 122 -243
rect 51 -256 52 -250
rect 96 -256 97 -250
rect 107 -251 108 -243
rect 107 -256 108 -250
rect 107 -251 108 -243
rect 107 -256 108 -250
rect 121 -256 122 -250
rect 135 -251 136 -243
rect 54 -253 55 -243
rect 82 -253 83 -243
rect 93 -253 94 -243
rect 114 -256 115 -252
rect 72 -256 73 -254
rect 100 -255 101 -243
rect 51 -266 52 -264
rect 58 -266 59 -264
rect 65 -266 66 -264
rect 89 -266 90 -264
rect 96 -266 97 -264
rect 121 -266 122 -264
rect 135 -271 136 -265
rect 138 -266 139 -264
rect 72 -268 73 -264
rect 82 -268 83 -264
rect 86 -268 87 -264
rect 107 -268 108 -264
rect 103 -270 104 -264
rect 114 -270 115 -264
rect 135 -281 136 -279
rect 145 -281 146 -279
<< labels >>
rlabel pdiffusion 3 -6 3 -6 0 cellNo=35
rlabel pdiffusion 10 -6 10 -6 0 cellNo=48
rlabel pdiffusion 17 -6 17 -6 0 cellNo=69
rlabel pdiffusion 52 -6 52 -6 0 feedthrough
rlabel pdiffusion 59 -6 59 -6 0 cellNo=30
rlabel pdiffusion 66 -6 66 -6 0 cellNo=34
rlabel pdiffusion 73 -6 73 -6 0 cellNo=95
rlabel pdiffusion 80 -6 80 -6 0 cellNo=40
rlabel pdiffusion 87 -6 87 -6 0 feedthrough
rlabel pdiffusion 94 -6 94 -6 0 cellNo=97
rlabel pdiffusion 101 -6 101 -6 0 feedthrough
rlabel pdiffusion 108 -6 108 -6 0 cellNo=51
rlabel pdiffusion 3 -23 3 -23 0 cellNo=41
rlabel pdiffusion 10 -23 10 -23 0 cellNo=15
rlabel pdiffusion 66 -23 66 -23 0 cellNo=18
rlabel pdiffusion 73 -23 73 -23 0 cellNo=5
rlabel pdiffusion 80 -23 80 -23 0 cellNo=68
rlabel pdiffusion 87 -23 87 -23 0 cellNo=71
rlabel pdiffusion 94 -23 94 -23 0 feedthrough
rlabel pdiffusion 101 -23 101 -23 0 feedthrough
rlabel pdiffusion 108 -23 108 -23 0 cellNo=17
rlabel pdiffusion 115 -23 115 -23 0 cellNo=63
rlabel pdiffusion 122 -23 122 -23 0 feedthrough
rlabel pdiffusion 3 -42 3 -42 0 cellNo=75
rlabel pdiffusion 45 -42 45 -42 0 cellNo=12
rlabel pdiffusion 52 -42 52 -42 0 feedthrough
rlabel pdiffusion 59 -42 59 -42 0 feedthrough
rlabel pdiffusion 66 -42 66 -42 0 cellNo=27
rlabel pdiffusion 73 -42 73 -42 0 cellNo=33
rlabel pdiffusion 80 -42 80 -42 0 cellNo=98
rlabel pdiffusion 87 -42 87 -42 0 cellNo=26
rlabel pdiffusion 94 -42 94 -42 0 cellNo=37
rlabel pdiffusion 101 -42 101 -42 0 feedthrough
rlabel pdiffusion 108 -42 108 -42 0 feedthrough
rlabel pdiffusion 115 -42 115 -42 0 feedthrough
rlabel pdiffusion 3 -63 3 -63 0 cellNo=92
rlabel pdiffusion 31 -63 31 -63 0 feedthrough
rlabel pdiffusion 38 -63 38 -63 0 feedthrough
rlabel pdiffusion 45 -63 45 -63 0 cellNo=60
rlabel pdiffusion 52 -63 52 -63 0 cellNo=32
rlabel pdiffusion 59 -63 59 -63 0 feedthrough
rlabel pdiffusion 66 -63 66 -63 0 feedthrough
rlabel pdiffusion 73 -63 73 -63 0 feedthrough
rlabel pdiffusion 80 -63 80 -63 0 cellNo=85
rlabel pdiffusion 87 -63 87 -63 0 cellNo=4
rlabel pdiffusion 94 -63 94 -63 0 cellNo=16
rlabel pdiffusion 101 -63 101 -63 0 feedthrough
rlabel pdiffusion 108 -63 108 -63 0 feedthrough
rlabel pdiffusion 115 -63 115 -63 0 cellNo=61
rlabel pdiffusion 24 -80 24 -80 0 cellNo=59
rlabel pdiffusion 38 -80 38 -80 0 cellNo=9
rlabel pdiffusion 45 -80 45 -80 0 feedthrough
rlabel pdiffusion 59 -80 59 -80 0 cellNo=43
rlabel pdiffusion 66 -80 66 -80 0 cellNo=55
rlabel pdiffusion 73 -80 73 -80 0 feedthrough
rlabel pdiffusion 80 -80 80 -80 0 feedthrough
rlabel pdiffusion 87 -80 87 -80 0 cellNo=42
rlabel pdiffusion 94 -80 94 -80 0 feedthrough
rlabel pdiffusion 101 -80 101 -80 0 feedthrough
rlabel pdiffusion 108 -80 108 -80 0 feedthrough
rlabel pdiffusion 115 -80 115 -80 0 cellNo=19
rlabel pdiffusion 122 -80 122 -80 0 cellNo=58
rlabel pdiffusion 129 -80 129 -80 0 feedthrough
rlabel pdiffusion 136 -80 136 -80 0 cellNo=90
rlabel pdiffusion 10 -101 10 -101 0 feedthrough
rlabel pdiffusion 17 -101 17 -101 0 cellNo=96
rlabel pdiffusion 24 -101 24 -101 0 cellNo=8
rlabel pdiffusion 31 -101 31 -101 0 feedthrough
rlabel pdiffusion 38 -101 38 -101 0 cellNo=2
rlabel pdiffusion 45 -101 45 -101 0 cellNo=45
rlabel pdiffusion 52 -101 52 -101 0 feedthrough
rlabel pdiffusion 59 -101 59 -101 0 feedthrough
rlabel pdiffusion 66 -101 66 -101 0 feedthrough
rlabel pdiffusion 73 -101 73 -101 0 cellNo=100
rlabel pdiffusion 80 -101 80 -101 0 cellNo=39
rlabel pdiffusion 87 -101 87 -101 0 cellNo=44
rlabel pdiffusion 94 -101 94 -101 0 cellNo=52
rlabel pdiffusion 101 -101 101 -101 0 feedthrough
rlabel pdiffusion 108 -101 108 -101 0 feedthrough
rlabel pdiffusion 115 -101 115 -101 0 cellNo=99
rlabel pdiffusion 122 -101 122 -101 0 feedthrough
rlabel pdiffusion 129 -101 129 -101 0 feedthrough
rlabel pdiffusion 136 -101 136 -101 0 feedthrough
rlabel pdiffusion 143 -101 143 -101 0 feedthrough
rlabel pdiffusion 150 -101 150 -101 0 feedthrough
rlabel pdiffusion 157 -101 157 -101 0 feedthrough
rlabel pdiffusion 31 -128 31 -128 0 feedthrough
rlabel pdiffusion 38 -128 38 -128 0 feedthrough
rlabel pdiffusion 45 -128 45 -128 0 feedthrough
rlabel pdiffusion 52 -128 52 -128 0 cellNo=83
rlabel pdiffusion 59 -128 59 -128 0 cellNo=67
rlabel pdiffusion 66 -128 66 -128 0 cellNo=94
rlabel pdiffusion 73 -128 73 -128 0 feedthrough
rlabel pdiffusion 80 -128 80 -128 0 feedthrough
rlabel pdiffusion 87 -128 87 -128 0 cellNo=84
rlabel pdiffusion 94 -128 94 -128 0 feedthrough
rlabel pdiffusion 101 -128 101 -128 0 cellNo=89
rlabel pdiffusion 108 -128 108 -128 0 cellNo=14
rlabel pdiffusion 115 -128 115 -128 0 cellNo=3
rlabel pdiffusion 122 -128 122 -128 0 cellNo=25
rlabel pdiffusion 129 -128 129 -128 0 feedthrough
rlabel pdiffusion 136 -128 136 -128 0 feedthrough
rlabel pdiffusion 143 -128 143 -128 0 feedthrough
rlabel pdiffusion 150 -128 150 -128 0 cellNo=72
rlabel pdiffusion 157 -128 157 -128 0 feedthrough
rlabel pdiffusion 164 -128 164 -128 0 feedthrough
rlabel pdiffusion 171 -128 171 -128 0 feedthrough
rlabel pdiffusion 178 -128 178 -128 0 feedthrough
rlabel pdiffusion 185 -128 185 -128 0 cellNo=56
rlabel pdiffusion 192 -128 192 -128 0 feedthrough
rlabel pdiffusion 10 -159 10 -159 0 feedthrough
rlabel pdiffusion 17 -159 17 -159 0 feedthrough
rlabel pdiffusion 24 -159 24 -159 0 feedthrough
rlabel pdiffusion 31 -159 31 -159 0 feedthrough
rlabel pdiffusion 38 -159 38 -159 0 feedthrough
rlabel pdiffusion 45 -159 45 -159 0 feedthrough
rlabel pdiffusion 52 -159 52 -159 0 cellNo=36
rlabel pdiffusion 59 -159 59 -159 0 cellNo=38
rlabel pdiffusion 66 -159 66 -159 0 cellNo=28
rlabel pdiffusion 73 -159 73 -159 0 cellNo=88
rlabel pdiffusion 80 -159 80 -159 0 feedthrough
rlabel pdiffusion 87 -159 87 -159 0 cellNo=29
rlabel pdiffusion 94 -159 94 -159 0 feedthrough
rlabel pdiffusion 101 -159 101 -159 0 cellNo=91
rlabel pdiffusion 108 -159 108 -159 0 feedthrough
rlabel pdiffusion 115 -159 115 -159 0 cellNo=78
rlabel pdiffusion 122 -159 122 -159 0 cellNo=87
rlabel pdiffusion 129 -159 129 -159 0 feedthrough
rlabel pdiffusion 136 -159 136 -159 0 cellNo=21
rlabel pdiffusion 143 -159 143 -159 0 feedthrough
rlabel pdiffusion 150 -159 150 -159 0 feedthrough
rlabel pdiffusion 157 -159 157 -159 0 feedthrough
rlabel pdiffusion 164 -159 164 -159 0 feedthrough
rlabel pdiffusion 171 -159 171 -159 0 feedthrough
rlabel pdiffusion 178 -159 178 -159 0 feedthrough
rlabel pdiffusion 185 -159 185 -159 0 cellNo=7
rlabel pdiffusion 31 -192 31 -192 0 feedthrough
rlabel pdiffusion 38 -192 38 -192 0 cellNo=80
rlabel pdiffusion 45 -192 45 -192 0 cellNo=46
rlabel pdiffusion 52 -192 52 -192 0 feedthrough
rlabel pdiffusion 59 -192 59 -192 0 feedthrough
rlabel pdiffusion 66 -192 66 -192 0 cellNo=22
rlabel pdiffusion 73 -192 73 -192 0 cellNo=74
rlabel pdiffusion 80 -192 80 -192 0 cellNo=47
rlabel pdiffusion 87 -192 87 -192 0 cellNo=66
rlabel pdiffusion 94 -192 94 -192 0 feedthrough
rlabel pdiffusion 101 -192 101 -192 0 cellNo=70
rlabel pdiffusion 108 -192 108 -192 0 feedthrough
rlabel pdiffusion 115 -192 115 -192 0 cellNo=64
rlabel pdiffusion 122 -192 122 -192 0 feedthrough
rlabel pdiffusion 129 -192 129 -192 0 cellNo=54
rlabel pdiffusion 136 -192 136 -192 0 feedthrough
rlabel pdiffusion 143 -192 143 -192 0 feedthrough
rlabel pdiffusion 150 -192 150 -192 0 feedthrough
rlabel pdiffusion 157 -192 157 -192 0 feedthrough
rlabel pdiffusion 164 -192 164 -192 0 feedthrough
rlabel pdiffusion 171 -192 171 -192 0 feedthrough
rlabel pdiffusion 178 -192 178 -192 0 feedthrough
rlabel pdiffusion 185 -192 185 -192 0 cellNo=62
rlabel pdiffusion 192 -192 192 -192 0 feedthrough
rlabel pdiffusion 45 -215 45 -215 0 cellNo=57
rlabel pdiffusion 52 -215 52 -215 0 feedthrough
rlabel pdiffusion 59 -215 59 -215 0 cellNo=31
rlabel pdiffusion 73 -215 73 -215 0 feedthrough
rlabel pdiffusion 80 -215 80 -215 0 cellNo=49
rlabel pdiffusion 87 -215 87 -215 0 feedthrough
rlabel pdiffusion 94 -215 94 -215 0 feedthrough
rlabel pdiffusion 101 -215 101 -215 0 cellNo=86
rlabel pdiffusion 108 -215 108 -215 0 feedthrough
rlabel pdiffusion 115 -215 115 -215 0 cellNo=24
rlabel pdiffusion 122 -215 122 -215 0 feedthrough
rlabel pdiffusion 129 -215 129 -215 0 cellNo=1
rlabel pdiffusion 136 -215 136 -215 0 cellNo=53
rlabel pdiffusion 143 -215 143 -215 0 cellNo=20
rlabel pdiffusion 150 -215 150 -215 0 feedthrough
rlabel pdiffusion 157 -215 157 -215 0 feedthrough
rlabel pdiffusion 31 -240 31 -240 0 feedthrough
rlabel pdiffusion 38 -240 38 -240 0 feedthrough
rlabel pdiffusion 45 -240 45 -240 0 feedthrough
rlabel pdiffusion 52 -240 52 -240 0 cellNo=10
rlabel pdiffusion 59 -240 59 -240 0 cellNo=50
rlabel pdiffusion 66 -240 66 -240 0 feedthrough
rlabel pdiffusion 73 -240 73 -240 0 cellNo=82
rlabel pdiffusion 80 -240 80 -240 0 cellNo=76
rlabel pdiffusion 87 -240 87 -240 0 cellNo=13
rlabel pdiffusion 94 -240 94 -240 0 cellNo=11
rlabel pdiffusion 101 -240 101 -240 0 cellNo=81
rlabel pdiffusion 108 -240 108 -240 0 feedthrough
rlabel pdiffusion 115 -240 115 -240 0 feedthrough
rlabel pdiffusion 122 -240 122 -240 0 feedthrough
rlabel pdiffusion 129 -240 129 -240 0 feedthrough
rlabel pdiffusion 136 -240 136 -240 0 feedthrough
rlabel pdiffusion 143 -240 143 -240 0 feedthrough
rlabel pdiffusion 52 -261 52 -261 0 feedthrough
rlabel pdiffusion 59 -261 59 -261 0 cellNo=79
rlabel pdiffusion 66 -261 66 -261 0 feedthrough
rlabel pdiffusion 73 -261 73 -261 0 feedthrough
rlabel pdiffusion 80 -261 80 -261 0 cellNo=65
rlabel pdiffusion 87 -261 87 -261 0 cellNo=93
rlabel pdiffusion 94 -261 94 -261 0 cellNo=23
rlabel pdiffusion 101 -261 101 -261 0 cellNo=73
rlabel pdiffusion 108 -261 108 -261 0 feedthrough
rlabel pdiffusion 115 -261 115 -261 0 feedthrough
rlabel pdiffusion 122 -261 122 -261 0 feedthrough
rlabel pdiffusion 136 -261 136 -261 0 cellNo=6
rlabel pdiffusion 136 -276 136 -276 0 feedthrough
rlabel pdiffusion 143 -276 143 -276 0 cellNo=77
rlabel polysilicon 51 -2 51 -2 0 1
rlabel polysilicon 51 -8 51 -8 0 3
rlabel polysilicon 58 -8 58 -8 0 3
rlabel polysilicon 61 -8 61 -8 0 4
rlabel polysilicon 65 -2 65 -2 0 1
rlabel polysilicon 72 -8 72 -8 0 3
rlabel polysilicon 79 -2 79 -2 0 1
rlabel polysilicon 79 -8 79 -8 0 3
rlabel polysilicon 86 -2 86 -2 0 1
rlabel polysilicon 86 -8 86 -8 0 3
rlabel polysilicon 93 -2 93 -2 0 1
rlabel polysilicon 100 -2 100 -2 0 1
rlabel polysilicon 100 -8 100 -8 0 3
rlabel polysilicon 107 -8 107 -8 0 3
rlabel polysilicon 110 -8 110 -8 0 4
rlabel polysilicon 9 -25 9 -25 0 3
rlabel polysilicon 12 -25 12 -25 0 4
rlabel polysilicon 65 -19 65 -19 0 1
rlabel polysilicon 68 -25 68 -25 0 4
rlabel polysilicon 75 -19 75 -19 0 2
rlabel polysilicon 72 -25 72 -25 0 3
rlabel polysilicon 75 -25 75 -25 0 4
rlabel polysilicon 82 -25 82 -25 0 4
rlabel polysilicon 86 -19 86 -19 0 1
rlabel polysilicon 89 -19 89 -19 0 2
rlabel polysilicon 93 -19 93 -19 0 1
rlabel polysilicon 93 -25 93 -25 0 3
rlabel polysilicon 100 -19 100 -19 0 1
rlabel polysilicon 100 -25 100 -25 0 3
rlabel polysilicon 110 -25 110 -25 0 4
rlabel polysilicon 114 -25 114 -25 0 3
rlabel polysilicon 121 -19 121 -19 0 1
rlabel polysilicon 121 -25 121 -25 0 3
rlabel polysilicon 47 -38 47 -38 0 2
rlabel polysilicon 51 -38 51 -38 0 1
rlabel polysilicon 51 -44 51 -44 0 3
rlabel polysilicon 58 -38 58 -38 0 1
rlabel polysilicon 58 -44 58 -44 0 3
rlabel polysilicon 68 -38 68 -38 0 2
rlabel polysilicon 72 -38 72 -38 0 1
rlabel polysilicon 75 -38 75 -38 0 2
rlabel polysilicon 72 -44 72 -44 0 3
rlabel polysilicon 82 -38 82 -38 0 2
rlabel polysilicon 79 -44 79 -44 0 3
rlabel polysilicon 82 -44 82 -44 0 4
rlabel polysilicon 86 -38 86 -38 0 1
rlabel polysilicon 89 -38 89 -38 0 2
rlabel polysilicon 86 -44 86 -44 0 3
rlabel polysilicon 96 -38 96 -38 0 2
rlabel polysilicon 93 -44 93 -44 0 3
rlabel polysilicon 96 -44 96 -44 0 4
rlabel polysilicon 100 -38 100 -38 0 1
rlabel polysilicon 100 -44 100 -44 0 3
rlabel polysilicon 107 -38 107 -38 0 1
rlabel polysilicon 107 -44 107 -44 0 3
rlabel polysilicon 114 -38 114 -38 0 1
rlabel polysilicon 114 -44 114 -44 0 3
rlabel polysilicon 30 -59 30 -59 0 1
rlabel polysilicon 30 -65 30 -65 0 3
rlabel polysilicon 37 -59 37 -59 0 1
rlabel polysilicon 37 -65 37 -65 0 3
rlabel polysilicon 44 -59 44 -59 0 1
rlabel polysilicon 47 -65 47 -65 0 4
rlabel polysilicon 51 -59 51 -59 0 1
rlabel polysilicon 54 -59 54 -59 0 2
rlabel polysilicon 58 -59 58 -59 0 1
rlabel polysilicon 58 -65 58 -65 0 3
rlabel polysilicon 65 -59 65 -59 0 1
rlabel polysilicon 65 -65 65 -65 0 3
rlabel polysilicon 72 -59 72 -59 0 1
rlabel polysilicon 72 -65 72 -65 0 3
rlabel polysilicon 79 -59 79 -59 0 1
rlabel polysilicon 82 -65 82 -65 0 4
rlabel polysilicon 89 -59 89 -59 0 2
rlabel polysilicon 86 -65 86 -65 0 3
rlabel polysilicon 89 -65 89 -65 0 4
rlabel polysilicon 96 -59 96 -59 0 2
rlabel polysilicon 96 -65 96 -65 0 4
rlabel polysilicon 100 -59 100 -59 0 1
rlabel polysilicon 100 -65 100 -65 0 3
rlabel polysilicon 107 -59 107 -59 0 1
rlabel polysilicon 107 -65 107 -65 0 3
rlabel polysilicon 114 -59 114 -59 0 1
rlabel polysilicon 117 -59 117 -59 0 2
rlabel polysilicon 117 -65 117 -65 0 4
rlabel polysilicon 23 -82 23 -82 0 3
rlabel polysilicon 26 -82 26 -82 0 4
rlabel polysilicon 40 -76 40 -76 0 2
rlabel polysilicon 40 -82 40 -82 0 4
rlabel polysilicon 44 -76 44 -76 0 1
rlabel polysilicon 44 -82 44 -82 0 3
rlabel polysilicon 61 -76 61 -76 0 2
rlabel polysilicon 58 -82 58 -82 0 3
rlabel polysilicon 61 -82 61 -82 0 4
rlabel polysilicon 65 -76 65 -76 0 1
rlabel polysilicon 68 -76 68 -76 0 2
rlabel polysilicon 65 -82 65 -82 0 3
rlabel polysilicon 68 -82 68 -82 0 4
rlabel polysilicon 72 -76 72 -76 0 1
rlabel polysilicon 72 -82 72 -82 0 3
rlabel polysilicon 79 -76 79 -76 0 1
rlabel polysilicon 79 -82 79 -82 0 3
rlabel polysilicon 86 -82 86 -82 0 3
rlabel polysilicon 89 -82 89 -82 0 4
rlabel polysilicon 93 -76 93 -76 0 1
rlabel polysilicon 93 -82 93 -82 0 3
rlabel polysilicon 100 -76 100 -76 0 1
rlabel polysilicon 100 -82 100 -82 0 3
rlabel polysilicon 107 -76 107 -76 0 1
rlabel polysilicon 107 -82 107 -82 0 3
rlabel polysilicon 114 -76 114 -76 0 1
rlabel polysilicon 124 -76 124 -76 0 2
rlabel polysilicon 124 -82 124 -82 0 4
rlabel polysilicon 128 -76 128 -76 0 1
rlabel polysilicon 128 -82 128 -82 0 3
rlabel polysilicon 135 -82 135 -82 0 3
rlabel polysilicon 9 -97 9 -97 0 1
rlabel polysilicon 9 -103 9 -103 0 3
rlabel polysilicon 16 -103 16 -103 0 3
rlabel polysilicon 26 -103 26 -103 0 4
rlabel polysilicon 30 -97 30 -97 0 1
rlabel polysilicon 30 -103 30 -103 0 3
rlabel polysilicon 40 -103 40 -103 0 4
rlabel polysilicon 47 -103 47 -103 0 4
rlabel polysilicon 51 -97 51 -97 0 1
rlabel polysilicon 51 -103 51 -103 0 3
rlabel polysilicon 58 -97 58 -97 0 1
rlabel polysilicon 58 -103 58 -103 0 3
rlabel polysilicon 65 -97 65 -97 0 1
rlabel polysilicon 65 -103 65 -103 0 3
rlabel polysilicon 72 -97 72 -97 0 1
rlabel polysilicon 75 -97 75 -97 0 2
rlabel polysilicon 72 -103 72 -103 0 3
rlabel polysilicon 75 -103 75 -103 0 4
rlabel polysilicon 79 -97 79 -97 0 1
rlabel polysilicon 79 -103 79 -103 0 3
rlabel polysilicon 82 -103 82 -103 0 4
rlabel polysilicon 86 -97 86 -97 0 1
rlabel polysilicon 89 -97 89 -97 0 2
rlabel polysilicon 86 -103 86 -103 0 3
rlabel polysilicon 89 -103 89 -103 0 4
rlabel polysilicon 96 -97 96 -97 0 2
rlabel polysilicon 93 -103 93 -103 0 3
rlabel polysilicon 96 -103 96 -103 0 4
rlabel polysilicon 100 -97 100 -97 0 1
rlabel polysilicon 100 -103 100 -103 0 3
rlabel polysilicon 107 -97 107 -97 0 1
rlabel polysilicon 107 -103 107 -103 0 3
rlabel polysilicon 114 -97 114 -97 0 1
rlabel polysilicon 117 -103 117 -103 0 4
rlabel polysilicon 121 -97 121 -97 0 1
rlabel polysilicon 121 -103 121 -103 0 3
rlabel polysilicon 128 -97 128 -97 0 1
rlabel polysilicon 128 -103 128 -103 0 3
rlabel polysilicon 135 -97 135 -97 0 1
rlabel polysilicon 135 -103 135 -103 0 3
rlabel polysilicon 142 -97 142 -97 0 1
rlabel polysilicon 142 -103 142 -103 0 3
rlabel polysilicon 149 -97 149 -97 0 1
rlabel polysilicon 149 -103 149 -103 0 3
rlabel polysilicon 156 -97 156 -97 0 1
rlabel polysilicon 156 -103 156 -103 0 3
rlabel polysilicon 30 -124 30 -124 0 1
rlabel polysilicon 30 -130 30 -130 0 3
rlabel polysilicon 37 -124 37 -124 0 1
rlabel polysilicon 37 -130 37 -130 0 3
rlabel polysilicon 44 -124 44 -124 0 1
rlabel polysilicon 44 -130 44 -130 0 3
rlabel polysilicon 51 -130 51 -130 0 3
rlabel polysilicon 54 -130 54 -130 0 4
rlabel polysilicon 61 -124 61 -124 0 2
rlabel polysilicon 58 -130 58 -130 0 3
rlabel polysilicon 61 -130 61 -130 0 4
rlabel polysilicon 65 -124 65 -124 0 1
rlabel polysilicon 65 -130 65 -130 0 3
rlabel polysilicon 68 -130 68 -130 0 4
rlabel polysilicon 72 -124 72 -124 0 1
rlabel polysilicon 72 -130 72 -130 0 3
rlabel polysilicon 79 -124 79 -124 0 1
rlabel polysilicon 79 -130 79 -130 0 3
rlabel polysilicon 86 -124 86 -124 0 1
rlabel polysilicon 89 -124 89 -124 0 2
rlabel polysilicon 86 -130 86 -130 0 3
rlabel polysilicon 89 -130 89 -130 0 4
rlabel polysilicon 93 -124 93 -124 0 1
rlabel polysilicon 93 -130 93 -130 0 3
rlabel polysilicon 103 -124 103 -124 0 2
rlabel polysilicon 107 -124 107 -124 0 1
rlabel polysilicon 110 -124 110 -124 0 2
rlabel polysilicon 107 -130 107 -130 0 3
rlabel polysilicon 110 -130 110 -130 0 4
rlabel polysilicon 114 -124 114 -124 0 1
rlabel polysilicon 117 -130 117 -130 0 4
rlabel polysilicon 121 -124 121 -124 0 1
rlabel polysilicon 124 -124 124 -124 0 2
rlabel polysilicon 128 -124 128 -124 0 1
rlabel polysilicon 128 -130 128 -130 0 3
rlabel polysilicon 135 -124 135 -124 0 1
rlabel polysilicon 135 -130 135 -130 0 3
rlabel polysilicon 142 -124 142 -124 0 1
rlabel polysilicon 142 -130 142 -130 0 3
rlabel polysilicon 152 -124 152 -124 0 2
rlabel polysilicon 149 -130 149 -130 0 3
rlabel polysilicon 156 -124 156 -124 0 1
rlabel polysilicon 156 -130 156 -130 0 3
rlabel polysilicon 163 -124 163 -124 0 1
rlabel polysilicon 163 -130 163 -130 0 3
rlabel polysilicon 170 -124 170 -124 0 1
rlabel polysilicon 170 -130 170 -130 0 3
rlabel polysilicon 177 -124 177 -124 0 1
rlabel polysilicon 177 -130 177 -130 0 3
rlabel polysilicon 187 -124 187 -124 0 2
rlabel polysilicon 184 -130 184 -130 0 3
rlabel polysilicon 191 -124 191 -124 0 1
rlabel polysilicon 191 -130 191 -130 0 3
rlabel polysilicon 9 -155 9 -155 0 1
rlabel polysilicon 9 -161 9 -161 0 3
rlabel polysilicon 16 -155 16 -155 0 1
rlabel polysilicon 16 -161 16 -161 0 3
rlabel polysilicon 23 -155 23 -155 0 1
rlabel polysilicon 23 -161 23 -161 0 3
rlabel polysilicon 30 -155 30 -155 0 1
rlabel polysilicon 30 -161 30 -161 0 3
rlabel polysilicon 37 -155 37 -155 0 1
rlabel polysilicon 37 -161 37 -161 0 3
rlabel polysilicon 44 -155 44 -155 0 1
rlabel polysilicon 44 -161 44 -161 0 3
rlabel polysilicon 51 -155 51 -155 0 1
rlabel polysilicon 54 -155 54 -155 0 2
rlabel polysilicon 51 -161 51 -161 0 3
rlabel polysilicon 61 -155 61 -155 0 2
rlabel polysilicon 58 -161 58 -161 0 3
rlabel polysilicon 61 -161 61 -161 0 4
rlabel polysilicon 68 -155 68 -155 0 2
rlabel polysilicon 65 -161 65 -161 0 3
rlabel polysilicon 72 -155 72 -155 0 1
rlabel polysilicon 72 -161 72 -161 0 3
rlabel polysilicon 75 -161 75 -161 0 4
rlabel polysilicon 79 -155 79 -155 0 1
rlabel polysilicon 79 -161 79 -161 0 3
rlabel polysilicon 86 -155 86 -155 0 1
rlabel polysilicon 86 -161 86 -161 0 3
rlabel polysilicon 93 -155 93 -155 0 1
rlabel polysilicon 93 -161 93 -161 0 3
rlabel polysilicon 100 -155 100 -155 0 1
rlabel polysilicon 103 -161 103 -161 0 4
rlabel polysilicon 107 -155 107 -155 0 1
rlabel polysilicon 107 -161 107 -161 0 3
rlabel polysilicon 114 -155 114 -155 0 1
rlabel polysilicon 117 -161 117 -161 0 4
rlabel polysilicon 121 -155 121 -155 0 1
rlabel polysilicon 124 -155 124 -155 0 2
rlabel polysilicon 121 -161 121 -161 0 3
rlabel polysilicon 124 -161 124 -161 0 4
rlabel polysilicon 128 -155 128 -155 0 1
rlabel polysilicon 128 -161 128 -161 0 3
rlabel polysilicon 135 -161 135 -161 0 3
rlabel polysilicon 142 -155 142 -155 0 1
rlabel polysilicon 142 -161 142 -161 0 3
rlabel polysilicon 149 -155 149 -155 0 1
rlabel polysilicon 149 -161 149 -161 0 3
rlabel polysilicon 156 -155 156 -155 0 1
rlabel polysilicon 156 -161 156 -161 0 3
rlabel polysilicon 163 -155 163 -155 0 1
rlabel polysilicon 163 -161 163 -161 0 3
rlabel polysilicon 170 -155 170 -155 0 1
rlabel polysilicon 170 -161 170 -161 0 3
rlabel polysilicon 177 -155 177 -155 0 1
rlabel polysilicon 177 -161 177 -161 0 3
rlabel polysilicon 184 -155 184 -155 0 1
rlabel polysilicon 184 -161 184 -161 0 3
rlabel polysilicon 187 -161 187 -161 0 4
rlabel polysilicon 30 -188 30 -188 0 1
rlabel polysilicon 30 -194 30 -194 0 3
rlabel polysilicon 37 -188 37 -188 0 1
rlabel polysilicon 44 -188 44 -188 0 1
rlabel polysilicon 47 -194 47 -194 0 4
rlabel polysilicon 51 -188 51 -188 0 1
rlabel polysilicon 51 -194 51 -194 0 3
rlabel polysilicon 58 -188 58 -188 0 1
rlabel polysilicon 58 -194 58 -194 0 3
rlabel polysilicon 65 -188 65 -188 0 1
rlabel polysilicon 68 -194 68 -194 0 4
rlabel polysilicon 72 -188 72 -188 0 1
rlabel polysilicon 75 -188 75 -188 0 2
rlabel polysilicon 72 -194 72 -194 0 3
rlabel polysilicon 79 -188 79 -188 0 1
rlabel polysilicon 82 -188 82 -188 0 2
rlabel polysilicon 86 -188 86 -188 0 1
rlabel polysilicon 86 -194 86 -194 0 3
rlabel polysilicon 93 -188 93 -188 0 1
rlabel polysilicon 93 -194 93 -194 0 3
rlabel polysilicon 100 -188 100 -188 0 1
rlabel polysilicon 100 -194 100 -194 0 3
rlabel polysilicon 103 -194 103 -194 0 4
rlabel polysilicon 107 -188 107 -188 0 1
rlabel polysilicon 107 -194 107 -194 0 3
rlabel polysilicon 114 -188 114 -188 0 1
rlabel polysilicon 117 -188 117 -188 0 2
rlabel polysilicon 121 -188 121 -188 0 1
rlabel polysilicon 121 -194 121 -194 0 3
rlabel polysilicon 128 -188 128 -188 0 1
rlabel polysilicon 131 -188 131 -188 0 2
rlabel polysilicon 135 -188 135 -188 0 1
rlabel polysilicon 135 -194 135 -194 0 3
rlabel polysilicon 142 -188 142 -188 0 1
rlabel polysilicon 142 -194 142 -194 0 3
rlabel polysilicon 149 -188 149 -188 0 1
rlabel polysilicon 149 -194 149 -194 0 3
rlabel polysilicon 156 -188 156 -188 0 1
rlabel polysilicon 156 -194 156 -194 0 3
rlabel polysilicon 163 -188 163 -188 0 1
rlabel polysilicon 163 -194 163 -194 0 3
rlabel polysilicon 170 -188 170 -188 0 1
rlabel polysilicon 170 -194 170 -194 0 3
rlabel polysilicon 177 -188 177 -188 0 1
rlabel polysilicon 177 -194 177 -194 0 3
rlabel polysilicon 187 -188 187 -188 0 2
rlabel polysilicon 191 -188 191 -188 0 1
rlabel polysilicon 191 -194 191 -194 0 3
rlabel polysilicon 44 -217 44 -217 0 3
rlabel polysilicon 51 -211 51 -211 0 1
rlabel polysilicon 51 -217 51 -217 0 3
rlabel polysilicon 61 -211 61 -211 0 2
rlabel polysilicon 72 -211 72 -211 0 1
rlabel polysilicon 72 -217 72 -217 0 3
rlabel polysilicon 82 -211 82 -211 0 2
rlabel polysilicon 86 -211 86 -211 0 1
rlabel polysilicon 86 -217 86 -217 0 3
rlabel polysilicon 93 -211 93 -211 0 1
rlabel polysilicon 93 -217 93 -217 0 3
rlabel polysilicon 100 -217 100 -217 0 3
rlabel polysilicon 103 -217 103 -217 0 4
rlabel polysilicon 107 -211 107 -211 0 1
rlabel polysilicon 107 -217 107 -217 0 3
rlabel polysilicon 114 -211 114 -211 0 1
rlabel polysilicon 117 -211 117 -211 0 2
rlabel polysilicon 121 -211 121 -211 0 1
rlabel polysilicon 121 -217 121 -217 0 3
rlabel polysilicon 128 -211 128 -211 0 1
rlabel polysilicon 128 -217 128 -217 0 3
rlabel polysilicon 131 -217 131 -217 0 4
rlabel polysilicon 138 -211 138 -211 0 2
rlabel polysilicon 138 -217 138 -217 0 4
rlabel polysilicon 142 -217 142 -217 0 3
rlabel polysilicon 149 -211 149 -211 0 1
rlabel polysilicon 149 -217 149 -217 0 3
rlabel polysilicon 156 -211 156 -211 0 1
rlabel polysilicon 156 -217 156 -217 0 3
rlabel polysilicon 30 -236 30 -236 0 1
rlabel polysilicon 30 -242 30 -242 0 3
rlabel polysilicon 37 -236 37 -236 0 1
rlabel polysilicon 37 -242 37 -242 0 3
rlabel polysilicon 44 -236 44 -236 0 1
rlabel polysilicon 44 -242 44 -242 0 3
rlabel polysilicon 51 -236 51 -236 0 1
rlabel polysilicon 54 -236 54 -236 0 2
rlabel polysilicon 54 -242 54 -242 0 4
rlabel polysilicon 58 -236 58 -236 0 1
rlabel polysilicon 61 -236 61 -236 0 2
rlabel polysilicon 65 -236 65 -236 0 1
rlabel polysilicon 65 -242 65 -242 0 3
rlabel polysilicon 75 -236 75 -236 0 2
rlabel polysilicon 72 -242 72 -242 0 3
rlabel polysilicon 75 -242 75 -242 0 4
rlabel polysilicon 79 -236 79 -236 0 1
rlabel polysilicon 82 -236 82 -236 0 2
rlabel polysilicon 82 -242 82 -242 0 4
rlabel polysilicon 86 -236 86 -236 0 1
rlabel polysilicon 89 -236 89 -236 0 2
rlabel polysilicon 86 -242 86 -242 0 3
rlabel polysilicon 89 -242 89 -242 0 4
rlabel polysilicon 93 -236 93 -236 0 1
rlabel polysilicon 93 -242 93 -242 0 3
rlabel polysilicon 103 -236 103 -236 0 2
rlabel polysilicon 100 -242 100 -242 0 3
rlabel polysilicon 107 -236 107 -236 0 1
rlabel polysilicon 107 -242 107 -242 0 3
rlabel polysilicon 114 -236 114 -236 0 1
rlabel polysilicon 114 -242 114 -242 0 3
rlabel polysilicon 121 -236 121 -236 0 1
rlabel polysilicon 121 -242 121 -242 0 3
rlabel polysilicon 128 -236 128 -236 0 1
rlabel polysilicon 128 -242 128 -242 0 3
rlabel polysilicon 135 -236 135 -236 0 1
rlabel polysilicon 135 -242 135 -242 0 3
rlabel polysilicon 142 -236 142 -236 0 1
rlabel polysilicon 142 -242 142 -242 0 3
rlabel polysilicon 51 -257 51 -257 0 1
rlabel polysilicon 51 -263 51 -263 0 3
rlabel polysilicon 61 -257 61 -257 0 2
rlabel polysilicon 58 -263 58 -263 0 3
rlabel polysilicon 65 -257 65 -257 0 1
rlabel polysilicon 65 -263 65 -263 0 3
rlabel polysilicon 72 -257 72 -257 0 1
rlabel polysilicon 72 -263 72 -263 0 3
rlabel polysilicon 79 -257 79 -257 0 1
rlabel polysilicon 82 -263 82 -263 0 4
rlabel polysilicon 86 -263 86 -263 0 3
rlabel polysilicon 89 -263 89 -263 0 4
rlabel polysilicon 96 -257 96 -257 0 2
rlabel polysilicon 96 -263 96 -263 0 4
rlabel polysilicon 103 -263 103 -263 0 4
rlabel polysilicon 107 -257 107 -257 0 1
rlabel polysilicon 107 -263 107 -263 0 3
rlabel polysilicon 114 -257 114 -257 0 1
rlabel polysilicon 114 -263 114 -263 0 3
rlabel polysilicon 121 -257 121 -257 0 1
rlabel polysilicon 121 -263 121 -263 0 3
rlabel polysilicon 138 -257 138 -257 0 2
rlabel polysilicon 138 -263 138 -263 0 4
rlabel polysilicon 135 -272 135 -272 0 1
rlabel polysilicon 135 -278 135 -278 0 3
rlabel polysilicon 145 -278 145 -278 0 4
rlabel metal2 51 1 51 1 0 net=307
rlabel metal2 79 1 79 1 0 net=135
rlabel metal2 93 1 93 1 0 net=237
rlabel metal2 51 -10 51 -10 0 net=308
rlabel metal2 65 -10 65 -10 0 net=66
rlabel metal2 79 -10 79 -10 0 net=51
rlabel metal2 58 -12 58 -12 0 net=6
rlabel metal2 89 -12 89 -12 0 net=238
rlabel metal2 107 -12 107 -12 0 net=217
rlabel metal2 86 -14 86 -14 0 net=137
rlabel metal2 86 -16 86 -16 0 net=117
rlabel metal2 9 -27 9 -27 0 net=23
rlabel metal2 58 -27 58 -27 0 net=163
rlabel metal2 107 -27 107 -27 0 net=221
rlabel metal2 114 -27 114 -27 0 net=218
rlabel metal2 68 -29 68 -29 0 net=46
rlabel metal2 82 -29 82 -29 0 net=138
rlabel metal2 47 -31 47 -31 0 net=64
rlabel metal2 86 -31 86 -31 0 net=263
rlabel metal2 51 -33 51 -33 0 net=285
rlabel metal2 72 -33 72 -33 0 net=93
rlabel metal2 96 -33 96 -33 0 net=201
rlabel metal2 72 -35 72 -35 0 net=118
rlabel metal2 37 -46 37 -46 0 net=291
rlabel metal2 51 -46 51 -46 0 net=286
rlabel metal2 89 -46 89 -46 0 net=264
rlabel metal2 30 -48 30 -48 0 net=171
rlabel metal2 54 -48 54 -48 0 net=133
rlabel metal2 79 -48 79 -48 0 net=20
rlabel metal2 72 -50 72 -50 0 net=70
rlabel metal2 96 -50 96 -50 0 net=222
rlabel metal2 58 -52 58 -52 0 net=164
rlabel metal2 100 -52 100 -52 0 net=203
rlabel metal2 58 -54 58 -54 0 net=107
rlabel metal2 100 -54 100 -54 0 net=113
rlabel metal2 72 -56 72 -56 0 net=267
rlabel metal2 30 -67 30 -67 0 net=172
rlabel metal2 58 -67 58 -67 0 net=108
rlabel metal2 93 -67 93 -67 0 net=109
rlabel metal2 37 -69 37 -69 0 net=292
rlabel metal2 65 -69 65 -69 0 net=134
rlabel metal2 72 -69 72 -69 0 net=268
rlabel metal2 96 -69 96 -69 0 net=204
rlabel metal2 117 -69 117 -69 0 net=309
rlabel metal2 40 -71 40 -71 0 net=141
rlabel metal2 65 -71 65 -71 0 net=125
rlabel metal2 79 -71 79 -71 0 net=115
rlabel metal2 107 -71 107 -71 0 net=273
rlabel metal2 89 -73 89 -73 0 net=189
rlabel metal2 9 -84 9 -84 0 net=213
rlabel metal2 26 -84 26 -84 0 net=53
rlabel metal2 51 -84 51 -84 0 net=275
rlabel metal2 100 -84 100 -84 0 net=191
rlabel metal2 128 -84 128 -84 0 net=311
rlabel metal2 30 -86 30 -86 0 net=143
rlabel metal2 58 -86 58 -86 0 net=74
rlabel metal2 72 -86 72 -86 0 net=126
rlabel metal2 72 -86 72 -86 0 net=126
rlabel metal2 75 -86 75 -86 0 net=247
rlabel metal2 135 -86 135 -86 0 net=269
rlabel metal2 135 -86 135 -86 0 net=269
rlabel metal2 79 -88 79 -88 0 net=116
rlabel metal2 107 -88 107 -88 0 net=274
rlabel metal2 58 -90 58 -90 0 net=123
rlabel metal2 86 -90 86 -90 0 net=103
rlabel metal2 114 -90 114 -90 0 net=169
rlabel metal2 65 -92 65 -92 0 net=14
rlabel metal2 93 -92 93 -92 0 net=111
rlabel metal2 61 -94 61 -94 0 net=119
rlabel metal2 86 -94 86 -94 0 net=253
rlabel metal2 9 -105 9 -105 0 net=214
rlabel metal2 26 -105 26 -105 0 net=96
rlabel metal2 82 -105 82 -105 0 net=192
rlabel metal2 124 -105 124 -105 0 net=299
rlabel metal2 187 -105 187 -105 0 net=293
rlabel metal2 30 -107 30 -107 0 net=144
rlabel metal2 44 -107 44 -107 0 net=227
rlabel metal2 65 -107 65 -107 0 net=121
rlabel metal2 86 -107 86 -107 0 net=104
rlabel metal2 103 -107 103 -107 0 net=170
rlabel metal2 30 -109 30 -109 0 net=225
rlabel metal2 117 -109 117 -109 0 net=270
rlabel metal2 142 -109 142 -109 0 net=313
rlabel metal2 37 -111 37 -111 0 net=193
rlabel metal2 93 -111 93 -111 0 net=112
rlabel metal2 114 -111 114 -111 0 net=257
rlabel metal2 47 -113 47 -113 0 net=124
rlabel metal2 75 -113 75 -113 0 net=199
rlabel metal2 121 -113 121 -113 0 net=295
rlabel metal2 51 -115 51 -115 0 net=276
rlabel metal2 128 -115 128 -115 0 net=249
rlabel metal2 128 -115 128 -115 0 net=249
rlabel metal2 135 -115 135 -115 0 net=255
rlabel metal2 65 -117 65 -117 0 net=3
rlabel metal2 152 -117 152 -117 0 net=279
rlabel metal2 79 -119 79 -119 0 net=251
rlabel metal2 86 -121 86 -121 0 net=35
rlabel metal2 23 -132 23 -132 0 net=229
rlabel metal2 61 -132 61 -132 0 net=200
rlabel metal2 110 -132 110 -132 0 net=314
rlabel metal2 16 -134 16 -134 0 net=235
rlabel metal2 68 -134 68 -134 0 net=122
rlabel metal2 79 -134 79 -134 0 net=252
rlabel metal2 107 -134 107 -134 0 net=243
rlabel metal2 30 -136 30 -136 0 net=226
rlabel metal2 68 -136 68 -136 0 net=145
rlabel metal2 100 -136 100 -136 0 net=159
rlabel metal2 117 -136 117 -136 0 net=256
rlabel metal2 149 -136 149 -136 0 net=300
rlabel metal2 9 -138 9 -138 0 net=297
rlabel metal2 72 -138 72 -138 0 net=94
rlabel metal2 121 -138 121 -138 0 net=296
rlabel metal2 30 -140 30 -140 0 net=127
rlabel metal2 124 -140 124 -140 0 net=219
rlabel metal2 156 -140 156 -140 0 net=281
rlabel metal2 44 -142 44 -142 0 net=105
rlabel metal2 114 -142 114 -142 0 net=233
rlabel metal2 128 -144 128 -144 0 net=250
rlabel metal2 86 -146 86 -146 0 net=165
rlabel metal2 142 -146 142 -146 0 net=259
rlabel metal2 184 -146 184 -146 0 net=294
rlabel metal2 37 -148 37 -148 0 net=195
rlabel metal2 37 -150 37 -150 0 net=177
rlabel metal2 54 -152 54 -152 0 net=155
rlabel metal2 9 -163 9 -163 0 net=298
rlabel metal2 75 -163 75 -163 0 net=69
rlabel metal2 23 -165 23 -165 0 net=230
rlabel metal2 61 -165 61 -165 0 net=160
rlabel metal2 128 -165 128 -165 0 net=167
rlabel metal2 30 -167 30 -167 0 net=128
rlabel metal2 79 -167 79 -167 0 net=147
rlabel metal2 128 -167 128 -167 0 net=260
rlabel metal2 30 -169 30 -169 0 net=149
rlabel metal2 103 -169 103 -169 0 net=32
rlabel metal2 131 -169 131 -169 0 net=265
rlabel metal2 37 -171 37 -171 0 net=178
rlabel metal2 117 -171 117 -171 0 net=161
rlabel metal2 135 -171 135 -171 0 net=282
rlabel metal2 16 -173 16 -173 0 net=236
rlabel metal2 44 -173 44 -173 0 net=106
rlabel metal2 117 -173 117 -173 0 net=220
rlabel metal2 156 -173 156 -173 0 net=234
rlabel metal2 44 -175 44 -175 0 net=73
rlabel metal2 149 -175 149 -175 0 net=245
rlabel metal2 51 -177 51 -177 0 net=301
rlabel metal2 75 -177 75 -177 0 net=50
rlabel metal2 114 -177 114 -177 0 net=209
rlabel metal2 170 -177 170 -177 0 net=271
rlabel metal2 58 -179 58 -179 0 net=157
rlabel metal2 142 -179 142 -179 0 net=197
rlabel metal2 65 -181 65 -181 0 net=179
rlabel metal2 79 -183 79 -183 0 net=183
rlabel metal2 93 -185 93 -185 0 net=151
rlabel metal2 30 -196 30 -196 0 net=150
rlabel metal2 68 -196 68 -196 0 net=148
rlabel metal2 117 -196 117 -196 0 net=266
rlabel metal2 58 -198 58 -198 0 net=158
rlabel metal2 86 -198 86 -198 0 net=198
rlabel metal2 51 -200 51 -200 0 net=303
rlabel metal2 82 -200 82 -200 0 net=239
rlabel metal2 100 -200 100 -200 0 net=162
rlabel metal2 128 -200 128 -200 0 net=272
rlabel metal2 47 -202 47 -202 0 net=139
rlabel metal2 93 -202 93 -202 0 net=153
rlabel metal2 138 -202 138 -202 0 net=246
rlabel metal2 156 -202 156 -202 0 net=211
rlabel metal2 156 -202 156 -202 0 net=211
rlabel metal2 93 -204 93 -204 0 net=283
rlabel metal2 142 -204 142 -204 0 net=185
rlabel metal2 103 -206 103 -206 0 net=168
rlabel metal2 107 -208 107 -208 0 net=181
rlabel metal2 30 -219 30 -219 0 net=129
rlabel metal2 61 -219 61 -219 0 net=284
rlabel metal2 103 -219 103 -219 0 net=287
rlabel metal2 138 -219 138 -219 0 net=186
rlabel metal2 44 -221 44 -221 0 net=140
rlabel metal2 54 -221 54 -221 0 net=55
rlabel metal2 103 -221 103 -221 0 net=182
rlabel metal2 121 -221 121 -221 0 net=154
rlabel metal2 142 -221 142 -221 0 net=212
rlabel metal2 37 -223 37 -223 0 net=305
rlabel metal2 65 -223 65 -223 0 net=173
rlabel metal2 89 -223 89 -223 0 net=215
rlabel metal2 128 -223 128 -223 0 net=261
rlabel metal2 44 -225 44 -225 0 net=277
rlabel metal2 75 -227 75 -227 0 net=205
rlabel metal2 79 -229 79 -229 0 net=223
rlabel metal2 86 -231 86 -231 0 net=241
rlabel metal2 72 -233 72 -233 0 net=304
rlabel metal2 30 -244 30 -244 0 net=130
rlabel metal2 65 -244 65 -244 0 net=175
rlabel metal2 65 -244 65 -244 0 net=175
rlabel metal2 79 -244 79 -244 0 net=216
rlabel metal2 138 -244 138 -244 0 net=262
rlabel metal2 37 -246 37 -246 0 net=306
rlabel metal2 86 -246 86 -246 0 net=242
rlabel metal2 44 -248 44 -248 0 net=278
rlabel metal2 89 -248 89 -248 0 net=224
rlabel metal2 51 -250 51 -250 0 net=187
rlabel metal2 107 -250 107 -250 0 net=207
rlabel metal2 107 -250 107 -250 0 net=207
rlabel metal2 121 -250 121 -250 0 net=289
rlabel metal2 54 -252 54 -252 0 net=83
rlabel metal2 93 -252 93 -252 0 net=131
rlabel metal2 72 -254 72 -254 0 net=101
rlabel metal2 51 -265 51 -265 0 net=188
rlabel metal2 65 -265 65 -265 0 net=176
rlabel metal2 96 -265 96 -265 0 net=290
rlabel metal2 135 -265 135 -265 0 net=231
rlabel metal2 72 -267 72 -267 0 net=102
rlabel metal2 86 -267 86 -267 0 net=208
rlabel metal2 103 -269 103 -269 0 net=132
rlabel metal2 135 -280 135 -280 0 net=232
<< end >>
